module basic_5000_50000_5000_200_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_130,In_1508);
xor U1 (N_1,In_2227,In_1955);
nand U2 (N_2,In_279,In_4676);
and U3 (N_3,In_3201,In_2124);
xor U4 (N_4,In_3995,In_2776);
nand U5 (N_5,In_1430,In_446);
xnor U6 (N_6,In_276,In_1422);
nand U7 (N_7,In_1342,In_490);
or U8 (N_8,In_986,In_2995);
or U9 (N_9,In_3750,In_2720);
or U10 (N_10,In_2994,In_3179);
or U11 (N_11,In_4385,In_1299);
or U12 (N_12,In_1116,In_2166);
nand U13 (N_13,In_3968,In_4023);
nor U14 (N_14,In_3161,In_2877);
or U15 (N_15,In_2749,In_2358);
and U16 (N_16,In_843,In_4192);
and U17 (N_17,In_4048,In_4378);
nand U18 (N_18,In_4167,In_2694);
nand U19 (N_19,In_235,In_1914);
and U20 (N_20,In_3707,In_4829);
nand U21 (N_21,In_2182,In_2319);
nand U22 (N_22,In_3277,In_2099);
nand U23 (N_23,In_18,In_49);
xnor U24 (N_24,In_4819,In_567);
and U25 (N_25,In_4109,In_3236);
and U26 (N_26,In_4517,In_4802);
and U27 (N_27,In_2086,In_2512);
or U28 (N_28,In_4103,In_3785);
or U29 (N_29,In_2596,In_1573);
xor U30 (N_30,In_1080,In_1418);
nand U31 (N_31,In_4709,In_1306);
and U32 (N_32,In_4081,In_444);
or U33 (N_33,In_4939,In_4730);
nand U34 (N_34,In_932,In_1839);
nand U35 (N_35,In_2217,In_4163);
or U36 (N_36,In_1200,In_4738);
nor U37 (N_37,In_2249,In_2208);
xnor U38 (N_38,In_3193,In_2944);
nand U39 (N_39,In_437,In_3931);
nand U40 (N_40,In_4274,In_4373);
nand U41 (N_41,In_281,In_3418);
or U42 (N_42,In_1178,In_4690);
xnor U43 (N_43,In_2882,In_3478);
xnor U44 (N_44,In_1603,In_1691);
nor U45 (N_45,In_55,In_439);
or U46 (N_46,In_1474,In_2379);
nand U47 (N_47,In_3199,In_4439);
nor U48 (N_48,In_1131,In_1888);
nor U49 (N_49,In_1582,In_773);
nand U50 (N_50,In_54,In_2840);
or U51 (N_51,In_1627,In_3532);
and U52 (N_52,In_1722,In_4796);
nor U53 (N_53,In_4040,In_1468);
or U54 (N_54,In_3318,In_4025);
nand U55 (N_55,In_497,In_4407);
or U56 (N_56,In_2525,In_3229);
nor U57 (N_57,In_2946,In_2583);
nand U58 (N_58,In_318,In_777);
nand U59 (N_59,In_1331,In_1000);
nand U60 (N_60,In_4967,In_3259);
xor U61 (N_61,In_325,In_103);
nor U62 (N_62,In_4985,In_1668);
or U63 (N_63,In_3767,In_1847);
nor U64 (N_64,In_1919,In_2385);
and U65 (N_65,In_1526,In_2355);
nor U66 (N_66,In_2120,In_227);
or U67 (N_67,In_1545,In_1031);
or U68 (N_68,In_1742,In_1317);
nor U69 (N_69,In_1107,In_2743);
or U70 (N_70,In_4760,In_4897);
nor U71 (N_71,In_1,In_3149);
and U72 (N_72,In_2490,In_4297);
xor U73 (N_73,In_2365,In_4506);
nor U74 (N_74,In_2737,In_2572);
nor U75 (N_75,In_1216,In_4642);
xor U76 (N_76,In_3728,In_4762);
and U77 (N_77,In_1989,In_2346);
and U78 (N_78,In_3312,In_2387);
or U79 (N_79,In_1466,In_2054);
or U80 (N_80,In_4994,In_3598);
or U81 (N_81,In_3485,In_26);
nand U82 (N_82,In_3714,In_3925);
nand U83 (N_83,In_3594,In_913);
nor U84 (N_84,In_1171,In_1821);
nor U85 (N_85,In_2618,In_2243);
nor U86 (N_86,In_4448,In_1601);
or U87 (N_87,In_4839,In_3586);
or U88 (N_88,In_2560,In_1834);
xnor U89 (N_89,In_4504,In_2866);
xor U90 (N_90,In_1053,In_2218);
xor U91 (N_91,In_3031,In_4921);
xnor U92 (N_92,In_2106,In_4085);
nand U93 (N_93,In_4152,In_3194);
nor U94 (N_94,In_4367,In_4420);
nor U95 (N_95,In_2517,In_1992);
and U96 (N_96,In_3162,In_725);
nand U97 (N_97,In_2532,In_4126);
nand U98 (N_98,In_3512,In_4519);
nand U99 (N_99,In_4004,In_2260);
xnor U100 (N_100,In_1854,In_2050);
xor U101 (N_101,In_300,In_2303);
xnor U102 (N_102,In_745,In_1935);
nor U103 (N_103,In_381,In_3319);
and U104 (N_104,In_826,In_3295);
nand U105 (N_105,In_4923,In_2757);
or U106 (N_106,In_2949,In_2812);
and U107 (N_107,In_476,In_2536);
nor U108 (N_108,In_1251,In_2666);
and U109 (N_109,In_1309,In_2224);
xor U110 (N_110,In_2448,In_2085);
or U111 (N_111,In_1666,In_2261);
and U112 (N_112,In_895,In_1607);
nor U113 (N_113,In_3231,In_268);
nor U114 (N_114,In_2063,In_2003);
or U115 (N_115,In_2384,In_3939);
and U116 (N_116,In_4983,In_4371);
and U117 (N_117,In_1684,In_2349);
nand U118 (N_118,In_1260,In_2065);
xor U119 (N_119,In_1767,In_3487);
nand U120 (N_120,In_4368,In_574);
and U121 (N_121,In_4454,In_3847);
xnor U122 (N_122,In_1170,In_2804);
nand U123 (N_123,In_1502,In_3751);
nor U124 (N_124,In_3207,In_271);
nor U125 (N_125,In_1290,In_4238);
or U126 (N_126,In_2912,In_4336);
nor U127 (N_127,In_1762,In_731);
nor U128 (N_128,In_4075,In_186);
nand U129 (N_129,In_880,In_833);
and U130 (N_130,In_2991,In_438);
nor U131 (N_131,In_4694,In_3286);
nand U132 (N_132,In_921,In_1010);
nand U133 (N_133,In_564,In_4876);
nor U134 (N_134,In_2865,In_4785);
xnor U135 (N_135,In_3365,In_1752);
nand U136 (N_136,In_1305,In_4417);
and U137 (N_137,In_3906,In_1493);
nor U138 (N_138,In_188,In_150);
nand U139 (N_139,In_1275,In_1106);
or U140 (N_140,In_1122,In_2441);
xor U141 (N_141,In_1494,In_2011);
nand U142 (N_142,In_4810,In_2271);
xnor U143 (N_143,In_781,In_2640);
nand U144 (N_144,In_1584,In_1467);
or U145 (N_145,In_4107,In_3469);
and U146 (N_146,In_1934,In_1844);
nor U147 (N_147,In_1091,In_2699);
and U148 (N_148,In_3007,In_1209);
and U149 (N_149,In_825,In_3926);
and U150 (N_150,In_4953,In_3025);
nor U151 (N_151,In_4665,In_478);
or U152 (N_152,In_1268,In_1723);
nand U153 (N_153,In_3701,In_798);
or U154 (N_154,In_3035,In_1866);
nor U155 (N_155,In_233,In_1193);
or U156 (N_156,In_4571,In_2102);
or U157 (N_157,In_4383,In_3611);
or U158 (N_158,In_1105,In_2623);
and U159 (N_159,In_4815,In_716);
and U160 (N_160,In_86,In_4707);
nand U161 (N_161,In_549,In_1486);
and U162 (N_162,In_4550,In_3816);
nand U163 (N_163,In_2678,In_3185);
xor U164 (N_164,In_2969,In_4283);
nor U165 (N_165,In_1337,In_297);
xor U166 (N_166,In_3501,In_3629);
and U167 (N_167,In_3648,In_4596);
nor U168 (N_168,In_583,In_962);
or U169 (N_169,In_2849,In_3516);
xnor U170 (N_170,In_4035,In_3972);
and U171 (N_171,In_3895,In_3668);
nor U172 (N_172,In_4534,In_754);
and U173 (N_173,In_4380,In_3104);
and U174 (N_174,In_2133,In_2191);
and U175 (N_175,In_1294,In_2343);
nand U176 (N_176,In_4943,In_4364);
nor U177 (N_177,In_1123,In_170);
nand U178 (N_178,In_4930,In_3517);
nand U179 (N_179,In_695,In_1232);
nand U180 (N_180,In_4271,In_3248);
and U181 (N_181,In_3637,In_4604);
xor U182 (N_182,In_2404,In_1527);
nand U183 (N_183,In_1375,In_917);
and U184 (N_184,In_1349,In_4486);
xnor U185 (N_185,In_2450,In_1033);
nor U186 (N_186,In_3669,In_3923);
nand U187 (N_187,In_4240,In_3155);
nor U188 (N_188,In_1744,In_3698);
or U189 (N_189,In_1581,In_3003);
and U190 (N_190,In_1340,In_3950);
nor U191 (N_191,In_2164,In_2126);
nand U192 (N_192,In_263,In_1089);
and U193 (N_193,In_4732,In_1956);
and U194 (N_194,In_116,In_3122);
nor U195 (N_195,In_4119,In_2281);
nor U196 (N_196,In_3994,In_1524);
xnor U197 (N_197,In_232,In_2884);
and U198 (N_198,In_2277,In_900);
nor U199 (N_199,In_1827,In_3342);
or U200 (N_200,In_3190,In_3435);
and U201 (N_201,In_4901,In_1185);
or U202 (N_202,In_2683,In_3971);
nand U203 (N_203,In_4833,In_4352);
nand U204 (N_204,In_2864,In_1730);
or U205 (N_205,In_2819,In_265);
nand U206 (N_206,In_4761,In_3301);
xor U207 (N_207,In_3726,In_4354);
nand U208 (N_208,In_2619,In_4675);
and U209 (N_209,In_3406,In_3244);
nor U210 (N_210,In_1499,In_1871);
and U211 (N_211,In_3840,In_1617);
xor U212 (N_212,In_1085,In_2007);
nor U213 (N_213,In_3583,In_2432);
xor U214 (N_214,In_925,In_3324);
or U215 (N_215,In_2053,In_1954);
nand U216 (N_216,In_3183,In_2792);
nand U217 (N_217,In_3173,In_4501);
nand U218 (N_218,In_4659,In_4422);
nor U219 (N_219,In_977,In_2297);
xnor U220 (N_220,In_4266,In_3504);
and U221 (N_221,In_4703,In_3924);
or U222 (N_222,In_3993,In_4891);
nor U223 (N_223,In_1168,In_2199);
and U224 (N_224,In_4357,In_1417);
or U225 (N_225,In_3294,In_4058);
nor U226 (N_226,In_4115,In_4838);
nand U227 (N_227,In_3720,In_4700);
nand U228 (N_228,In_4072,In_231);
and U229 (N_229,In_4453,In_3903);
and U230 (N_230,In_4197,In_2809);
or U231 (N_231,In_723,In_1024);
or U232 (N_232,In_3030,In_4108);
nand U233 (N_233,In_3021,In_2984);
nand U234 (N_234,In_1857,In_1565);
xnor U235 (N_235,In_4055,In_3097);
xor U236 (N_236,In_1343,In_4818);
xnor U237 (N_237,In_1728,In_587);
nand U238 (N_238,In_377,In_316);
and U239 (N_239,In_378,In_1945);
nor U240 (N_240,In_3609,In_4854);
nand U241 (N_241,In_264,In_4456);
nand U242 (N_242,In_68,In_34);
xnor U243 (N_243,In_1177,In_3266);
xnor U244 (N_244,In_197,In_1921);
nand U245 (N_245,In_2424,In_3397);
or U246 (N_246,In_3800,In_3940);
or U247 (N_247,In_4595,In_1917);
or U248 (N_248,In_3797,In_1246);
or U249 (N_249,In_4823,In_152);
xor U250 (N_250,In_685,In_3577);
xnor U251 (N_251,In_2301,In_537);
or U252 (N_252,In_660,In_4711);
nand U253 (N_253,In_4840,In_2515);
and U254 (N_254,In_3922,In_2159);
nand U255 (N_255,In_342,In_1427);
nand U256 (N_256,In_2276,In_3380);
xor U257 (N_257,In_2713,In_2751);
xnor U258 (N_258,In_1274,In_1987);
and U259 (N_259,In_4621,In_99);
nand U260 (N_260,In_4104,In_205);
nand U261 (N_261,In_3716,N_148);
xnor U262 (N_262,In_693,In_4204);
or U263 (N_263,In_3588,In_410);
xnor U264 (N_264,In_4544,In_3929);
nand U265 (N_265,N_179,In_1735);
and U266 (N_266,In_1883,In_960);
and U267 (N_267,In_2937,In_1994);
xnor U268 (N_268,In_217,In_4117);
and U269 (N_269,In_230,In_74);
and U270 (N_270,In_1555,In_4080);
and U271 (N_271,In_3001,In_273);
nor U272 (N_272,In_4019,In_3006);
nor U273 (N_273,In_3886,In_1937);
nor U274 (N_274,In_330,In_3690);
and U275 (N_275,In_935,In_1140);
nor U276 (N_276,In_4122,In_4050);
xor U277 (N_277,In_3537,N_29);
xnor U278 (N_278,In_807,In_2556);
or U279 (N_279,In_2674,In_1947);
xnor U280 (N_280,In_4977,In_3742);
xnor U281 (N_281,In_4490,In_795);
xor U282 (N_282,N_32,In_3676);
and U283 (N_283,N_141,In_2451);
nand U284 (N_284,In_4415,In_2562);
xnor U285 (N_285,In_1488,In_275);
nand U286 (N_286,In_3565,In_598);
and U287 (N_287,In_4817,In_529);
xor U288 (N_288,In_3325,N_70);
or U289 (N_289,In_2136,In_3269);
nand U290 (N_290,In_2643,In_3362);
and U291 (N_291,In_3459,In_4687);
and U292 (N_292,In_3234,In_2844);
xor U293 (N_293,In_3002,In_4386);
xor U294 (N_294,In_1428,In_319);
nor U295 (N_295,In_3808,In_1498);
xor U296 (N_296,In_3761,In_3531);
nand U297 (N_297,In_841,In_661);
and U298 (N_298,In_1591,In_538);
or U299 (N_299,In_1678,In_4461);
nand U300 (N_300,In_765,In_2847);
nor U301 (N_301,In_688,In_1461);
and U302 (N_302,In_404,In_2048);
xnor U303 (N_303,In_1538,In_3297);
nor U304 (N_304,In_2103,In_3889);
nand U305 (N_305,In_4405,In_3921);
and U306 (N_306,In_3076,N_127);
xnor U307 (N_307,In_3946,In_128);
or U308 (N_308,In_1137,In_1230);
or U309 (N_309,In_2073,In_2466);
and U310 (N_310,In_4426,In_2993);
nor U311 (N_311,In_3261,In_4451);
nor U312 (N_312,In_3715,In_4160);
nand U313 (N_313,In_1109,In_1166);
nor U314 (N_314,In_4601,In_3635);
nand U315 (N_315,In_3029,In_3096);
and U316 (N_316,In_2597,In_1070);
or U317 (N_317,In_4173,In_1902);
nor U318 (N_318,In_1640,In_568);
xnor U319 (N_319,In_4264,In_3412);
nand U320 (N_320,In_4531,In_2222);
and U321 (N_321,In_4775,In_3752);
xnor U322 (N_322,In_1289,In_3053);
nor U323 (N_323,In_274,In_4963);
xnor U324 (N_324,In_3382,In_4844);
xnor U325 (N_325,In_1506,In_1151);
xor U326 (N_326,In_2704,In_2843);
or U327 (N_327,In_4344,In_4555);
xor U328 (N_328,In_818,In_1923);
nor U329 (N_329,In_4398,In_968);
nor U330 (N_330,In_345,N_215);
and U331 (N_331,In_3191,In_4106);
and U332 (N_332,In_3832,N_200);
and U333 (N_333,In_3178,In_4217);
or U334 (N_334,In_1062,In_4671);
nor U335 (N_335,In_4443,In_3340);
or U336 (N_336,In_261,N_111);
xnor U337 (N_337,In_1890,In_1804);
and U338 (N_338,In_4482,In_3528);
and U339 (N_339,In_4165,In_1088);
or U340 (N_340,In_3468,In_3477);
nor U341 (N_341,In_1361,In_1279);
xnor U342 (N_342,In_4828,In_1835);
nand U343 (N_343,In_3361,In_2338);
nand U344 (N_344,In_67,In_701);
xnor U345 (N_345,In_3456,In_1451);
or U346 (N_346,In_4056,In_4276);
and U347 (N_347,In_737,In_3333);
xnor U348 (N_348,In_4583,In_1240);
and U349 (N_349,In_4199,In_1720);
xor U350 (N_350,In_2397,In_2921);
xnor U351 (N_351,In_1759,In_2446);
nand U352 (N_352,In_3270,In_2661);
xor U353 (N_353,N_4,In_3147);
or U354 (N_354,In_1570,In_4776);
and U355 (N_355,In_4885,In_4142);
xor U356 (N_356,In_2571,In_1783);
nor U357 (N_357,In_4651,In_2582);
nor U358 (N_358,N_56,In_1985);
and U359 (N_359,In_2922,In_1977);
xor U360 (N_360,In_3275,In_4693);
and U361 (N_361,In_4114,In_28);
nand U362 (N_362,In_2600,In_2433);
nand U363 (N_363,In_458,In_1030);
xor U364 (N_364,In_2098,In_1798);
xnor U365 (N_365,In_2286,N_236);
or U366 (N_366,In_1163,In_2101);
nand U367 (N_367,N_171,In_1731);
xnor U368 (N_368,N_206,In_2235);
or U369 (N_369,In_3084,In_4189);
nand U370 (N_370,In_1434,In_2726);
nor U371 (N_371,In_4580,N_97);
and U372 (N_372,N_175,In_1159);
nor U373 (N_373,In_1132,In_1906);
or U374 (N_374,In_1415,In_3536);
or U375 (N_375,In_2669,In_2284);
and U376 (N_376,In_361,In_1761);
or U377 (N_377,In_2603,In_4273);
and U378 (N_378,In_2593,In_3127);
nand U379 (N_379,In_391,In_2851);
and U380 (N_380,In_4610,In_2196);
nand U381 (N_381,In_4944,In_1393);
or U382 (N_382,In_4881,In_2302);
xor U383 (N_383,In_4585,In_647);
nand U384 (N_384,In_3257,In_4300);
and U385 (N_385,N_98,In_3136);
xor U386 (N_386,In_610,In_1850);
nand U387 (N_387,In_4090,In_1768);
nand U388 (N_388,In_1266,In_4812);
nor U389 (N_389,In_4771,In_4190);
or U390 (N_390,In_3640,In_4622);
nand U391 (N_391,In_3449,In_3225);
and U392 (N_392,In_4299,In_748);
or U393 (N_393,In_4589,In_3055);
xor U394 (N_394,In_1374,N_82);
nor U395 (N_395,In_2421,In_2900);
or U396 (N_396,In_4617,In_2841);
xor U397 (N_397,In_4475,In_2814);
nor U398 (N_398,In_4379,In_3241);
and U399 (N_399,In_4597,In_3163);
or U400 (N_400,In_4993,In_3421);
xnor U401 (N_401,In_2317,In_1776);
nand U402 (N_402,In_738,In_496);
xnor U403 (N_403,In_30,In_2692);
or U404 (N_404,In_4030,In_3796);
nor U405 (N_405,In_3189,In_1069);
nand U406 (N_406,In_1512,N_115);
or U407 (N_407,In_1843,In_4800);
nand U408 (N_408,In_4070,N_102);
nand U409 (N_409,In_1223,N_201);
xnor U410 (N_410,In_3633,In_1135);
or U411 (N_411,N_186,In_1881);
and U412 (N_412,In_3144,In_834);
and U413 (N_413,In_617,In_3059);
or U414 (N_414,N_17,In_4302);
nor U415 (N_415,In_3011,In_842);
xor U416 (N_416,In_4867,In_1420);
or U417 (N_417,In_2916,In_590);
nor U418 (N_418,In_1625,In_1050);
nand U419 (N_419,In_2251,In_4442);
xnor U420 (N_420,In_3102,In_3486);
nor U421 (N_421,In_2676,In_1805);
or U422 (N_422,In_332,In_2188);
and U423 (N_423,In_62,In_2893);
or U424 (N_424,In_3441,In_1702);
or U425 (N_425,In_2725,N_249);
xnor U426 (N_426,In_4479,N_225);
or U427 (N_427,In_1202,In_618);
nor U428 (N_428,In_2585,In_956);
or U429 (N_429,In_4646,In_1929);
nand U430 (N_430,In_1865,In_1121);
xnor U431 (N_431,In_4015,In_2783);
and U432 (N_432,In_4399,In_4057);
or U433 (N_433,In_113,In_3483);
xor U434 (N_434,N_85,In_206);
nand U435 (N_435,In_770,In_2483);
nand U436 (N_436,In_1283,In_1118);
nor U437 (N_437,In_4971,In_222);
and U438 (N_438,In_1087,In_721);
nor U439 (N_439,In_83,In_46);
and U440 (N_440,In_266,In_2953);
nor U441 (N_441,In_2568,N_131);
nor U442 (N_442,In_472,In_1351);
and U443 (N_443,In_4492,In_4612);
xor U444 (N_444,In_2735,In_4384);
or U445 (N_445,In_3187,N_244);
nand U446 (N_446,In_4547,In_1300);
xor U447 (N_447,In_3019,In_4212);
and U448 (N_448,In_2129,N_34);
nor U449 (N_449,In_4991,In_577);
xnor U450 (N_450,In_3065,In_4934);
or U451 (N_451,In_741,In_3466);
or U452 (N_452,In_4598,In_3520);
or U453 (N_453,In_1450,In_4491);
and U454 (N_454,In_1282,In_4633);
nor U455 (N_455,In_489,N_139);
or U456 (N_456,In_1602,In_3978);
xnor U457 (N_457,In_41,In_4673);
or U458 (N_458,In_3192,In_461);
or U459 (N_459,In_2779,In_1739);
or U460 (N_460,In_3222,In_2455);
and U461 (N_461,In_4446,In_2083);
xor U462 (N_462,In_3892,In_3167);
nand U463 (N_463,In_4602,In_4314);
or U464 (N_464,In_899,N_213);
and U465 (N_465,In_4868,In_1846);
xor U466 (N_466,In_2702,In_4086);
and U467 (N_467,In_794,In_2059);
and U468 (N_468,In_1515,In_4554);
or U469 (N_469,In_4347,In_3729);
nor U470 (N_470,In_310,In_696);
and U471 (N_471,In_124,In_2340);
nor U472 (N_472,In_3708,In_4100);
xor U473 (N_473,In_4409,In_623);
nor U474 (N_474,In_2219,In_1704);
and U475 (N_475,In_3949,In_555);
and U476 (N_476,In_3237,In_1732);
nand U477 (N_477,In_1808,N_33);
xnor U478 (N_478,In_1622,In_4756);
nor U479 (N_479,In_2706,In_3928);
and U480 (N_480,In_397,N_109);
xor U481 (N_481,In_1242,In_561);
nor U482 (N_482,In_845,In_3589);
or U483 (N_483,In_335,In_59);
nor U484 (N_484,In_3581,In_2748);
or U485 (N_485,N_217,N_147);
nor U486 (N_486,In_884,In_4681);
nand U487 (N_487,In_485,In_2823);
or U488 (N_488,In_1599,In_2428);
xnor U489 (N_489,In_2604,In_625);
nor U490 (N_490,In_1423,In_4712);
nand U491 (N_491,In_2764,In_578);
xnor U492 (N_492,N_247,In_190);
xor U493 (N_493,In_2153,In_3743);
or U494 (N_494,In_4870,In_4431);
and U495 (N_495,In_2256,In_573);
and U496 (N_496,In_3366,In_905);
or U497 (N_497,In_4986,In_3592);
xor U498 (N_498,In_1476,In_2128);
and U499 (N_499,In_180,In_3314);
or U500 (N_500,In_3659,In_2904);
xor U501 (N_501,In_644,In_237);
or U502 (N_502,In_3492,In_1635);
nor U503 (N_503,N_153,N_137);
nand U504 (N_504,N_461,In_3845);
xor U505 (N_505,In_2056,In_4942);
nand U506 (N_506,In_1411,In_1608);
and U507 (N_507,N_205,In_1891);
xor U508 (N_508,In_3680,N_255);
nor U509 (N_509,In_2097,In_3371);
xnor U510 (N_510,N_157,In_3665);
xor U511 (N_511,In_1519,In_1303);
or U512 (N_512,In_4722,In_3211);
and U513 (N_513,In_1687,In_2724);
or U514 (N_514,In_430,N_110);
and U515 (N_515,In_2906,In_3563);
or U516 (N_516,N_421,In_4306);
or U517 (N_517,In_1714,In_1692);
or U518 (N_518,In_1483,In_2440);
xor U519 (N_519,In_2506,In_2482);
nand U520 (N_520,In_4852,In_2550);
or U521 (N_521,N_425,In_4037);
or U522 (N_522,In_828,In_2067);
nor U523 (N_523,In_2519,In_4961);
xor U524 (N_524,In_4503,In_4396);
nand U525 (N_525,In_4495,N_112);
nand U526 (N_526,In_3447,In_1447);
xor U527 (N_527,In_4801,In_2878);
xor U528 (N_528,In_1416,In_2345);
xor U529 (N_529,In_4112,In_112);
nand U530 (N_530,In_2143,In_3175);
xnor U531 (N_531,In_4905,N_466);
nand U532 (N_532,In_1165,In_73);
nor U533 (N_533,In_3881,In_2853);
nand U534 (N_534,In_2013,In_1345);
nor U535 (N_535,N_152,In_1455);
or U536 (N_536,In_1385,In_77);
xor U537 (N_537,In_4325,In_3541);
nand U538 (N_538,In_504,In_289);
or U539 (N_539,N_92,In_1071);
and U540 (N_540,In_3116,In_2452);
or U541 (N_541,In_1661,In_2967);
nand U542 (N_542,In_4261,In_1381);
nand U543 (N_543,In_1364,N_370);
and U544 (N_544,In_3781,In_3628);
nor U545 (N_545,N_362,In_2614);
and U546 (N_546,In_3529,In_2335);
xor U547 (N_547,N_192,In_3488);
nand U548 (N_548,In_1205,In_1550);
nand U549 (N_549,In_1931,In_4728);
xor U550 (N_550,In_1976,In_492);
nor U551 (N_551,N_260,In_2119);
nand U552 (N_552,In_1228,N_301);
xor U553 (N_553,In_4795,In_1243);
xnor U554 (N_554,In_2610,N_410);
or U555 (N_555,In_3126,In_683);
nand U556 (N_556,In_2653,In_3268);
or U557 (N_557,In_2104,N_181);
or U558 (N_558,In_4444,N_391);
xor U559 (N_559,In_2832,In_949);
nand U560 (N_560,In_76,In_4726);
nand U561 (N_561,In_2088,N_395);
and U562 (N_562,In_363,In_3176);
nor U563 (N_563,In_941,N_83);
nand U564 (N_564,In_4882,In_1669);
xor U565 (N_565,In_4937,In_3717);
nand U566 (N_566,In_105,In_3775);
and U567 (N_567,In_431,In_3219);
and U568 (N_568,In_182,In_1459);
nor U569 (N_569,In_350,In_3860);
nand U570 (N_570,In_985,In_2531);
nand U571 (N_571,In_1997,In_2584);
or U572 (N_572,In_4960,In_2631);
nand U573 (N_573,In_3534,In_728);
and U574 (N_574,In_2563,In_2732);
xnor U575 (N_575,In_1514,In_3841);
or U576 (N_576,In_609,N_316);
and U577 (N_577,In_865,In_2662);
and U578 (N_578,In_1660,In_885);
or U579 (N_579,In_2500,N_145);
nand U580 (N_580,In_4680,In_3613);
and U581 (N_581,In_2107,In_1112);
nor U582 (N_582,In_1067,In_1549);
or U583 (N_583,N_79,In_983);
and U584 (N_584,In_4592,In_3283);
and U585 (N_585,In_589,In_4270);
or U586 (N_586,In_2739,In_3137);
nor U587 (N_587,In_3792,N_135);
nand U588 (N_588,In_3885,In_2839);
and U589 (N_589,In_402,In_3580);
nor U590 (N_590,In_1966,In_3415);
and U591 (N_591,In_1480,In_1249);
nor U592 (N_592,In_322,In_69);
xnor U593 (N_593,In_2348,In_4753);
nand U594 (N_594,In_3322,In_4790);
nor U595 (N_595,In_4661,In_2366);
nand U596 (N_596,In_401,In_2318);
and U597 (N_597,In_1536,In_4510);
nor U598 (N_598,In_671,In_3696);
nor U599 (N_599,In_873,In_2649);
nand U600 (N_600,In_2760,In_3471);
xor U601 (N_601,In_2797,In_4186);
nand U602 (N_602,In_1039,In_2105);
and U603 (N_603,In_3139,In_3658);
xnor U604 (N_604,In_514,In_3671);
xnor U605 (N_605,In_3455,In_2232);
xor U606 (N_606,In_3113,In_3771);
and U607 (N_607,In_3854,In_2288);
nor U608 (N_608,N_400,In_4140);
nand U609 (N_609,In_4539,In_1736);
nand U610 (N_610,In_3706,In_495);
and U611 (N_611,In_2237,In_1706);
nor U612 (N_612,In_4335,In_4226);
and U613 (N_613,In_2770,In_4470);
nand U614 (N_614,In_846,In_1950);
xnor U615 (N_615,In_3616,In_4850);
and U616 (N_616,In_3082,In_4908);
nor U617 (N_617,N_487,In_4424);
and U618 (N_618,In_3393,N_27);
nor U619 (N_619,In_2486,In_2872);
xnor U620 (N_620,In_4154,In_3779);
or U621 (N_621,In_1542,In_1988);
nor U622 (N_622,In_449,In_4704);
or U623 (N_623,In_425,In_2989);
and U624 (N_624,In_955,In_2688);
nand U625 (N_625,In_4193,In_768);
or U626 (N_626,In_3081,In_772);
xor U627 (N_627,In_3794,In_2579);
and U628 (N_628,In_2507,In_3141);
nand U629 (N_629,In_3484,In_1452);
nand U630 (N_630,In_861,In_1196);
xor U631 (N_631,In_382,In_2156);
xor U632 (N_632,In_3042,In_1245);
xor U633 (N_633,In_3355,In_3846);
nand U634 (N_634,In_1990,In_211);
nor U635 (N_635,In_1566,In_2753);
and U636 (N_636,In_4759,In_4176);
nand U637 (N_637,In_3016,In_3036);
xnor U638 (N_638,N_259,In_763);
xor U639 (N_639,In_4806,In_2274);
nand U640 (N_640,In_3230,In_1855);
nor U641 (N_641,In_3905,In_635);
and U642 (N_642,In_3443,In_70);
xor U643 (N_643,In_1115,In_1445);
nand U644 (N_644,In_898,In_3734);
nand U645 (N_645,In_4845,In_3777);
or U646 (N_646,N_170,In_122);
nor U647 (N_647,In_3280,In_2311);
and U648 (N_648,In_1191,In_3754);
xor U649 (N_649,In_5,N_440);
nand U650 (N_650,In_4014,In_4627);
and U651 (N_651,In_1119,In_2030);
xor U652 (N_652,In_870,In_506);
xnor U653 (N_653,In_1878,In_32);
nor U654 (N_654,N_21,In_3975);
nand U655 (N_655,In_2295,In_1236);
xor U656 (N_656,In_511,In_3884);
nor U657 (N_657,N_158,In_3212);
nand U658 (N_658,In_2738,In_4235);
nand U659 (N_659,In_4082,In_930);
nor U660 (N_660,In_3411,N_3);
and U661 (N_661,In_2412,N_354);
or U662 (N_662,In_575,In_700);
xor U663 (N_663,In_2495,In_560);
or U664 (N_664,In_84,In_1983);
xnor U665 (N_665,In_185,N_420);
nor U666 (N_666,N_458,In_1758);
and U667 (N_667,In_23,In_280);
xor U668 (N_668,In_2833,In_3046);
nor U669 (N_669,In_4318,In_106);
or U670 (N_670,In_1108,In_4928);
and U671 (N_671,In_926,In_4996);
xnor U672 (N_672,In_3839,In_3111);
nand U673 (N_673,In_2716,In_1104);
nor U674 (N_674,In_2194,N_309);
and U675 (N_675,In_2091,In_3769);
nor U676 (N_676,In_3666,In_1296);
xnor U677 (N_677,In_2342,In_2200);
nor U678 (N_678,In_427,In_3883);
and U679 (N_679,In_2975,In_247);
nor U680 (N_680,In_3871,In_707);
xnor U681 (N_681,In_3265,In_600);
or U682 (N_682,N_241,In_570);
or U683 (N_683,In_1049,In_3156);
xnor U684 (N_684,In_2496,In_2836);
nand U685 (N_685,In_4032,N_392);
or U686 (N_686,In_1095,In_1101);
and U687 (N_687,N_130,In_2331);
or U688 (N_688,In_4628,In_970);
and U689 (N_689,N_185,In_4696);
xor U690 (N_690,In_220,In_2628);
or U691 (N_691,In_3224,In_3562);
and U692 (N_692,N_396,In_2493);
nor U693 (N_693,In_286,In_894);
nor U694 (N_694,In_2031,In_2869);
nor U695 (N_695,In_2670,In_4515);
nand U696 (N_696,In_2,In_4564);
nand U697 (N_697,In_1414,In_4254);
xnor U698 (N_698,In_2821,In_4195);
xnor U699 (N_699,In_2259,In_3251);
xor U700 (N_700,In_1490,In_920);
nor U701 (N_701,In_3085,In_1713);
xnor U702 (N_702,In_2035,In_2959);
and U703 (N_703,N_286,In_2411);
xnor U704 (N_704,In_1754,In_2229);
and U705 (N_705,In_1726,In_3758);
or U706 (N_706,In_1378,In_973);
nor U707 (N_707,In_1586,N_336);
nor U708 (N_708,In_1153,In_4654);
xor U709 (N_709,In_938,In_3851);
and U710 (N_710,In_1329,In_4747);
nor U711 (N_711,In_2971,In_221);
nand U712 (N_712,In_2489,In_4618);
nor U713 (N_713,In_2715,In_4557);
or U714 (N_714,In_1585,In_320);
and U715 (N_715,N_113,In_705);
xor U716 (N_716,N_194,In_3413);
nor U717 (N_717,In_2272,In_200);
nor U718 (N_718,In_1578,N_220);
nor U719 (N_719,In_4536,In_3083);
xor U720 (N_720,In_3866,In_3656);
xor U721 (N_721,N_101,In_4808);
and U722 (N_722,In_3159,In_2491);
or U723 (N_723,In_910,In_958);
nand U724 (N_724,In_3546,N_402);
nand U725 (N_725,N_231,In_374);
nor U726 (N_726,In_415,In_1598);
xor U727 (N_727,In_3506,In_4484);
and U728 (N_728,N_457,In_1148);
and U729 (N_729,In_2296,In_2216);
nor U730 (N_730,In_4686,In_2405);
nor U731 (N_731,In_1576,In_2762);
xor U732 (N_732,In_4907,In_3735);
and U733 (N_733,In_1833,In_3732);
and U734 (N_734,In_3444,In_24);
nor U735 (N_735,N_372,In_1457);
nor U736 (N_736,N_472,In_650);
nor U737 (N_737,In_42,In_407);
nor U738 (N_738,In_2238,In_2837);
nand U739 (N_739,In_4246,In_2150);
xnor U740 (N_740,N_118,In_2807);
xor U741 (N_741,In_764,In_4774);
nand U742 (N_742,In_4549,In_1740);
or U743 (N_743,In_2508,In_1352);
nor U744 (N_744,In_358,In_3688);
or U745 (N_745,In_2072,In_2001);
and U746 (N_746,In_3317,In_697);
or U747 (N_747,N_405,In_3465);
and U748 (N_748,In_752,In_682);
nand U749 (N_749,In_4174,In_3585);
nor U750 (N_750,In_4381,In_904);
nor U751 (N_751,In_2747,In_278);
nand U752 (N_752,In_2282,In_4649);
or U753 (N_753,In_3497,In_2827);
or U754 (N_754,In_3374,In_3595);
xor U755 (N_755,In_2205,In_1253);
xnor U756 (N_756,In_4206,In_4750);
and U757 (N_757,In_4421,In_3684);
xnor U758 (N_758,In_2045,In_4029);
nor U759 (N_759,N_559,In_451);
nor U760 (N_760,In_3419,In_724);
and U761 (N_761,In_1145,In_852);
xnor U762 (N_762,In_3174,In_178);
nand U763 (N_763,In_2589,In_991);
nor U764 (N_764,In_1077,In_2817);
or U765 (N_765,In_2790,In_4865);
nor U766 (N_766,In_4435,In_3605);
xor U767 (N_767,In_4211,In_2978);
or U768 (N_768,In_4169,In_3938);
nor U769 (N_769,In_1973,In_2524);
nor U770 (N_770,N_654,N_657);
nand U771 (N_771,In_1633,In_409);
or U772 (N_772,In_3855,In_3305);
nand U773 (N_773,In_889,In_3302);
or U774 (N_774,In_1717,In_1207);
nand U775 (N_775,N_504,N_12);
and U776 (N_776,N_547,In_4600);
or U777 (N_777,In_857,In_288);
nor U778 (N_778,In_927,In_1897);
nand U779 (N_779,In_3810,In_4258);
xnor U780 (N_780,In_2633,In_855);
xor U781 (N_781,In_3438,In_4856);
nor U782 (N_782,In_4219,In_2210);
and U783 (N_783,In_2874,In_251);
and U784 (N_784,In_4408,In_3642);
and U785 (N_785,N_696,In_1036);
or U786 (N_786,In_448,In_4031);
and U787 (N_787,In_2816,In_3772);
and U788 (N_788,In_4562,In_2268);
or U789 (N_789,In_144,In_4053);
and U790 (N_790,In_1880,In_3203);
nor U791 (N_791,N_723,N_417);
or U792 (N_792,In_1120,In_787);
and U793 (N_793,In_2039,In_2997);
or U794 (N_794,In_3952,In_1583);
xnor U795 (N_795,In_192,N_532);
xnor U796 (N_796,In_1321,In_1386);
xnor U797 (N_797,In_3762,In_4280);
nand U798 (N_798,In_3112,In_699);
or U799 (N_799,In_2990,In_676);
nor U800 (N_800,In_2968,In_1082);
xor U801 (N_801,In_1750,In_1297);
xnor U802 (N_802,N_24,In_2198);
nand U803 (N_803,In_3327,In_4241);
or U804 (N_804,In_799,In_213);
nand U805 (N_805,In_4691,In_4441);
xor U806 (N_806,In_4780,N_353);
nand U807 (N_807,In_3326,In_2019);
nor U808 (N_808,In_1792,In_634);
nand U809 (N_809,In_523,In_3409);
xor U810 (N_810,In_4419,In_3332);
or U811 (N_811,In_1656,In_380);
and U812 (N_812,In_4578,In_4500);
nor U813 (N_813,In_1868,N_544);
or U814 (N_814,In_2467,In_2068);
and U815 (N_815,In_4215,In_3394);
and U816 (N_816,In_4180,In_972);
nor U817 (N_817,In_4360,N_228);
or U818 (N_818,In_1712,N_534);
nand U819 (N_819,In_940,In_2066);
nand U820 (N_820,In_2768,N_341);
nand U821 (N_821,In_524,In_229);
xnor U822 (N_822,In_2530,In_4629);
nor U823 (N_823,In_201,In_4948);
xnor U824 (N_824,In_4874,In_4740);
nand U825 (N_825,In_1370,In_513);
nor U826 (N_826,In_4932,In_1020);
xor U827 (N_827,In_1905,In_1454);
xor U828 (N_828,In_2523,N_611);
and U829 (N_829,N_183,In_4432);
and U830 (N_830,In_4287,In_1092);
or U831 (N_831,In_110,In_2665);
xor U832 (N_832,In_2012,In_3338);
nand U833 (N_833,In_4764,In_3651);
and U834 (N_834,In_1190,In_1637);
and U835 (N_835,In_902,In_1649);
and U836 (N_836,In_1763,In_2828);
xnor U837 (N_837,In_3947,In_1680);
nand U838 (N_838,In_872,In_1859);
or U839 (N_839,In_2168,In_3618);
xor U840 (N_840,In_2701,In_3867);
xor U841 (N_841,N_748,N_271);
nor U842 (N_842,N_590,N_367);
or U843 (N_843,In_2236,In_1980);
nand U844 (N_844,In_3216,In_3223);
nor U845 (N_845,In_2020,In_980);
and U846 (N_846,N_625,In_1961);
nand U847 (N_847,In_3600,In_4038);
or U848 (N_848,In_2055,In_718);
or U849 (N_849,In_1167,In_353);
or U850 (N_850,In_1594,In_2474);
and U851 (N_851,In_3639,N_50);
nand U852 (N_852,In_3724,In_3760);
or U853 (N_853,In_1060,In_204);
and U854 (N_854,In_2587,In_616);
or U855 (N_855,In_1657,In_1628);
xor U856 (N_856,N_269,In_4846);
nand U857 (N_857,In_1225,In_4331);
xor U858 (N_858,In_372,In_1356);
xor U859 (N_859,In_2145,In_4305);
or U860 (N_860,In_2176,In_2648);
or U861 (N_861,In_1063,N_677);
nand U862 (N_862,In_4717,In_491);
or U863 (N_863,In_3143,In_1965);
and U864 (N_864,In_3835,In_1828);
xor U865 (N_865,In_670,In_3508);
nor U866 (N_866,In_659,In_4791);
and U867 (N_867,N_253,In_3252);
nand U868 (N_868,In_3457,In_3258);
nand U869 (N_869,In_4896,In_2336);
and U870 (N_870,In_3709,In_1802);
xor U871 (N_871,In_4637,N_278);
xnor U872 (N_872,In_3607,In_2986);
and U873 (N_873,In_3335,In_4509);
xnor U874 (N_874,In_791,In_2551);
xnor U875 (N_875,N_393,In_2044);
or U876 (N_876,In_4565,In_4296);
and U877 (N_877,N_239,In_816);
nand U878 (N_878,N_562,In_3786);
and U879 (N_879,In_2423,In_592);
and U880 (N_880,In_3285,In_269);
nand U881 (N_881,In_3507,In_835);
xor U882 (N_882,N_62,In_4540);
nand U883 (N_883,In_4445,In_4231);
xnor U884 (N_884,In_4834,In_483);
and U885 (N_885,In_469,In_4736);
nand U886 (N_886,In_4350,In_3791);
nand U887 (N_887,In_1860,In_1478);
nor U888 (N_888,In_2540,In_822);
or U889 (N_889,In_3292,In_1051);
xor U890 (N_890,In_2557,In_92);
nand U891 (N_891,In_1034,In_1948);
nor U892 (N_892,In_1575,In_2657);
nand U893 (N_893,In_2650,In_1967);
nor U894 (N_894,In_3290,In_3996);
nor U895 (N_895,In_1007,In_686);
or U896 (N_896,In_4135,In_102);
nor U897 (N_897,N_52,N_427);
xor U898 (N_898,In_4118,In_4389);
nor U899 (N_899,In_2856,In_4358);
nand U900 (N_900,In_4895,In_2686);
xor U901 (N_901,In_3099,In_2534);
or U902 (N_902,In_527,In_562);
xor U903 (N_903,In_4518,In_3549);
xnor U904 (N_904,In_2520,In_2171);
nor U905 (N_905,In_4918,N_295);
nor U906 (N_906,In_4458,In_2009);
xor U907 (N_907,In_4999,In_2914);
and U908 (N_908,In_1286,In_719);
nor U909 (N_909,In_1548,In_3138);
nor U910 (N_910,In_743,In_3856);
nand U911 (N_911,In_2449,In_4835);
or U912 (N_912,In_2356,In_3559);
nand U913 (N_913,In_4634,In_760);
or U914 (N_914,In_1567,In_3819);
xnor U915 (N_915,In_3617,In_3250);
nor U916 (N_916,In_1589,In_3664);
and U917 (N_917,N_477,In_950);
xnor U918 (N_918,In_3308,In_2860);
xnor U919 (N_919,In_3217,N_550);
or U920 (N_920,N_602,In_1809);
or U921 (N_921,In_343,In_4579);
xnor U922 (N_922,In_858,In_1975);
and U923 (N_923,In_936,In_80);
nor U924 (N_924,In_493,In_4767);
xor U925 (N_925,In_2416,In_1125);
or U926 (N_926,In_3678,In_1256);
or U927 (N_927,In_3347,In_678);
and U928 (N_928,In_224,In_1682);
xnor U929 (N_929,In_1943,In_164);
xor U930 (N_930,In_4758,In_3661);
xor U931 (N_931,In_4041,In_1397);
nor U932 (N_932,In_3299,In_907);
xnor U933 (N_933,In_4033,N_707);
nor U934 (N_934,In_887,In_3132);
and U935 (N_935,In_1743,In_1690);
xor U936 (N_936,In_4682,In_3417);
or U937 (N_937,In_2209,N_630);
xor U938 (N_938,In_1748,In_3255);
xor U939 (N_939,N_432,N_223);
nand U940 (N_940,In_61,In_2388);
nand U941 (N_941,In_252,N_735);
nand U942 (N_942,N_711,In_4949);
and U943 (N_943,In_1870,N_533);
xor U944 (N_944,In_1577,In_2677);
or U945 (N_945,N_612,In_675);
or U946 (N_946,In_2766,In_2987);
or U947 (N_947,In_3437,In_601);
or U948 (N_948,N_488,In_3602);
xnor U949 (N_949,In_3496,In_4433);
nand U950 (N_950,In_3276,N_203);
or U951 (N_951,In_1227,N_256);
and U952 (N_952,In_1876,In_207);
and U953 (N_953,In_771,In_4772);
or U954 (N_954,In_435,In_756);
xor U955 (N_955,In_1426,In_988);
and U956 (N_956,N_519,In_3392);
and U957 (N_957,N_413,In_4468);
nand U958 (N_958,In_223,In_2857);
xnor U959 (N_959,In_2383,In_3513);
nand U960 (N_960,In_3249,In_2413);
and U961 (N_961,In_3514,In_3899);
xor U962 (N_962,In_4706,In_4613);
xnor U963 (N_963,In_1658,N_328);
and U964 (N_964,In_2875,N_23);
and U965 (N_965,In_3168,In_3426);
or U966 (N_966,In_4912,In_154);
and U967 (N_967,In_2786,N_383);
and U968 (N_968,In_1288,In_1936);
and U969 (N_969,N_15,In_1693);
and U970 (N_970,In_136,In_3755);
nand U971 (N_971,N_198,In_1102);
or U972 (N_972,In_1449,In_3948);
and U973 (N_973,In_3215,In_4990);
nor U974 (N_974,In_2542,In_3089);
and U975 (N_975,In_944,N_250);
and U976 (N_976,In_2292,In_639);
and U977 (N_977,N_745,In_886);
nor U978 (N_978,In_4872,In_4260);
xnor U979 (N_979,In_3930,N_378);
or U980 (N_980,In_2811,In_1262);
nor U981 (N_981,In_3721,In_4312);
and U982 (N_982,In_412,In_4428);
nor U983 (N_983,In_2613,In_1141);
xor U984 (N_984,In_1711,In_4060);
and U985 (N_985,In_1563,In_4369);
nor U986 (N_986,In_2158,In_1530);
xor U987 (N_987,N_208,In_2970);
nand U988 (N_988,N_166,N_668);
nand U989 (N_989,In_1534,In_4811);
nor U990 (N_990,In_4572,In_769);
nor U991 (N_991,N_510,In_3452);
nand U992 (N_992,In_4851,In_107);
nand U993 (N_993,In_1293,In_658);
or U994 (N_994,In_912,In_867);
xnor U995 (N_995,In_1647,N_469);
xor U996 (N_996,In_4803,N_484);
and U997 (N_997,In_1579,In_3238);
or U998 (N_998,In_3873,In_3645);
xnor U999 (N_999,In_2607,In_2703);
nor U1000 (N_1000,In_1473,In_1214);
xnor U1001 (N_1001,In_3677,In_2956);
nor U1002 (N_1002,In_732,In_928);
and U1003 (N_1003,In_3364,In_4269);
xnor U1004 (N_1004,In_3103,N_990);
nand U1005 (N_1005,In_3783,In_3172);
nand U1006 (N_1006,N_140,In_4127);
and U1007 (N_1007,In_305,In_1932);
or U1008 (N_1008,In_2246,In_2769);
and U1009 (N_1009,In_2403,In_4866);
nor U1010 (N_1010,In_711,N_867);
and U1011 (N_1011,In_3653,In_3766);
xor U1012 (N_1012,In_863,In_2754);
xnor U1013 (N_1013,In_4914,In_167);
and U1014 (N_1014,In_1619,In_3125);
nor U1015 (N_1015,In_4825,In_3430);
and U1016 (N_1016,In_641,In_3603);
nand U1017 (N_1017,N_246,In_2920);
xor U1018 (N_1018,In_3756,In_4615);
or U1019 (N_1019,In_2599,N_926);
and U1020 (N_1020,In_994,In_640);
or U1021 (N_1021,N_233,In_2498);
xor U1022 (N_1022,In_3288,N_522);
xnor U1023 (N_1023,In_2468,N_717);
xnor U1024 (N_1024,In_4313,In_82);
and U1025 (N_1025,N_37,In_2925);
xnor U1026 (N_1026,In_706,In_3197);
and U1027 (N_1027,In_727,In_3008);
xnor U1028 (N_1028,N_73,In_1683);
and U1029 (N_1029,N_42,N_25);
and U1030 (N_1030,In_569,In_57);
nand U1031 (N_1031,N_965,In_789);
and U1032 (N_1032,In_421,N_296);
nand U1033 (N_1033,In_2609,In_2016);
nor U1034 (N_1034,In_877,N_731);
xor U1035 (N_1035,N_305,In_357);
xor U1036 (N_1036,In_160,In_2736);
or U1037 (N_1037,N_585,In_4607);
or U1038 (N_1038,N_188,In_508);
nand U1039 (N_1039,In_1117,In_1963);
xor U1040 (N_1040,In_1822,In_3321);
or U1041 (N_1041,In_2655,In_3383);
and U1042 (N_1042,In_420,In_2095);
nor U1043 (N_1043,In_2265,In_3699);
xnor U1044 (N_1044,N_890,In_291);
nor U1045 (N_1045,In_4282,In_4301);
nand U1046 (N_1046,In_2503,N_714);
xor U1047 (N_1047,N_627,In_1696);
xor U1048 (N_1048,In_3829,In_4087);
or U1049 (N_1049,In_1634,In_4830);
xnor U1050 (N_1050,In_1667,In_1316);
and U1051 (N_1051,In_2658,In_4185);
nor U1052 (N_1052,In_3330,N_207);
or U1053 (N_1053,N_950,In_1755);
xnor U1054 (N_1054,In_1968,In_759);
xor U1055 (N_1055,In_3853,In_1043);
nor U1056 (N_1056,In_3408,In_3509);
nor U1057 (N_1057,In_1244,In_2436);
or U1058 (N_1058,N_841,In_4341);
xnor U1059 (N_1059,In_2203,In_4789);
xnor U1060 (N_1060,N_416,In_1765);
or U1061 (N_1061,In_1161,In_2697);
and U1062 (N_1062,In_4976,N_938);
nand U1063 (N_1063,N_360,In_3169);
and U1064 (N_1064,In_2698,In_3646);
nand U1065 (N_1065,N_507,N_960);
or U1066 (N_1066,In_2394,In_4765);
xor U1067 (N_1067,In_2533,N_783);
xor U1068 (N_1068,In_3557,In_307);
xnor U1069 (N_1069,In_3120,In_1332);
and U1070 (N_1070,In_4130,N_512);
xor U1071 (N_1071,N_914,In_4769);
nand U1072 (N_1072,In_4366,In_892);
nand U1073 (N_1073,In_1221,In_2273);
and U1074 (N_1074,In_3511,In_1675);
nor U1075 (N_1075,In_2146,In_4702);
or U1076 (N_1076,In_2820,N_227);
and U1077 (N_1077,N_872,In_2731);
and U1078 (N_1078,In_2636,In_4599);
nor U1079 (N_1079,N_332,In_847);
or U1080 (N_1080,N_937,N_397);
nand U1081 (N_1081,In_4172,In_4998);
nor U1082 (N_1082,In_3606,N_121);
nand U1083 (N_1083,N_476,In_4209);
or U1084 (N_1084,In_2125,In_4877);
or U1085 (N_1085,In_540,N_688);
or U1086 (N_1086,In_979,In_183);
nand U1087 (N_1087,In_4098,In_2439);
nand U1088 (N_1088,In_3119,In_293);
or U1089 (N_1089,In_4847,In_1872);
or U1090 (N_1090,N_613,In_3587);
and U1091 (N_1091,In_1624,N_156);
or U1092 (N_1092,N_825,N_775);
and U1093 (N_1093,In_2214,In_3253);
nand U1094 (N_1094,In_81,In_4097);
nand U1095 (N_1095,In_1390,N_59);
nand U1096 (N_1096,In_792,In_2131);
nor U1097 (N_1097,In_606,N_573);
or U1098 (N_1098,In_4843,In_1005);
nor U1099 (N_1099,In_3850,In_3154);
nor U1100 (N_1100,In_996,In_4430);
xor U1101 (N_1101,In_243,In_2901);
nor U1102 (N_1102,In_2339,In_14);
nor U1103 (N_1103,In_4848,In_2891);
nand U1104 (N_1104,In_1784,N_248);
and U1105 (N_1105,In_1694,In_1172);
xor U1106 (N_1106,In_3110,In_2504);
xor U1107 (N_1107,In_3747,In_1265);
and U1108 (N_1108,In_2492,In_4516);
and U1109 (N_1109,N_609,N_282);
xor U1110 (N_1110,In_4489,In_142);
xor U1111 (N_1111,In_4593,In_3737);
xor U1112 (N_1112,N_746,In_4524);
or U1113 (N_1113,In_3121,In_2149);
and U1114 (N_1114,In_4862,In_4134);
nand U1115 (N_1115,In_976,In_630);
xor U1116 (N_1116,In_677,In_4695);
or U1117 (N_1117,In_627,In_4899);
and U1118 (N_1118,In_25,In_2710);
and U1119 (N_1119,N_483,In_2714);
xor U1120 (N_1120,In_1285,In_4224);
and U1121 (N_1121,In_3378,In_3573);
xor U1122 (N_1122,In_3227,In_3911);
nor U1123 (N_1123,In_3311,N_321);
or U1124 (N_1124,In_2240,In_2248);
xnor U1125 (N_1125,In_2673,N_0);
nor U1126 (N_1126,In_2481,In_1993);
or U1127 (N_1127,N_403,In_1124);
nand U1128 (N_1128,In_2316,N_523);
nor U1129 (N_1129,In_4992,N_842);
xnor U1130 (N_1130,In_1312,In_1898);
xnor U1131 (N_1131,In_984,In_3339);
nand U1132 (N_1132,In_3878,In_3558);
nand U1133 (N_1133,In_169,In_2911);
xor U1134 (N_1134,In_4755,In_1176);
or U1135 (N_1135,In_1057,In_761);
nor U1136 (N_1136,In_434,In_4251);
xor U1137 (N_1137,In_4625,In_1188);
xnor U1138 (N_1138,In_1778,In_3641);
nand U1139 (N_1139,N_319,In_146);
xnor U1140 (N_1140,In_1926,In_830);
nor U1141 (N_1141,N_373,N_802);
nor U1142 (N_1142,In_4664,In_1097);
xor U1143 (N_1143,In_4437,N_693);
or U1144 (N_1144,In_2808,In_1032);
xnor U1145 (N_1145,In_3391,In_4965);
nor U1146 (N_1146,N_406,In_4626);
and U1147 (N_1147,N_230,N_634);
xnor U1148 (N_1148,In_2220,In_1795);
nor U1149 (N_1149,N_338,N_411);
and U1150 (N_1150,N_49,In_2269);
nand U1151 (N_1151,In_2926,N_193);
or U1152 (N_1152,In_3186,In_4792);
or U1153 (N_1153,In_2800,N_214);
xor U1154 (N_1154,In_4362,In_4513);
nand U1155 (N_1155,In_3177,In_2859);
xor U1156 (N_1156,In_1477,N_969);
nor U1157 (N_1157,In_4272,N_940);
nand U1158 (N_1158,In_668,In_3390);
nand U1159 (N_1159,In_2154,In_1354);
nand U1160 (N_1160,In_2708,In_552);
or U1161 (N_1161,N_312,In_1023);
xor U1162 (N_1162,In_680,N_434);
nand U1163 (N_1163,In_3180,In_2115);
nor U1164 (N_1164,N_368,In_1212);
xor U1165 (N_1165,In_4718,In_2641);
nor U1166 (N_1166,In_4012,In_2873);
xor U1167 (N_1167,In_1796,In_2695);
nor U1168 (N_1168,In_747,N_105);
nor U1169 (N_1169,N_790,In_466);
nor U1170 (N_1170,N_889,In_893);
nand U1171 (N_1171,In_3912,In_2730);
xor U1172 (N_1172,In_4447,In_2791);
nand U1173 (N_1173,In_1916,In_517);
xor U1174 (N_1174,In_1681,In_2036);
nor U1175 (N_1175,N_540,In_488);
nand U1176 (N_1176,N_238,N_252);
or U1177 (N_1177,N_245,In_1469);
or U1178 (N_1178,In_4917,In_1424);
and U1179 (N_1179,N_822,In_4624);
and U1180 (N_1180,In_4317,In_1884);
or U1181 (N_1181,In_1688,In_4363);
and U1182 (N_1182,In_815,In_4981);
xnor U1183 (N_1183,In_3117,In_3263);
xor U1184 (N_1184,In_3359,N_587);
nor U1185 (N_1185,In_3129,In_4807);
xor U1186 (N_1186,In_238,In_1041);
xor U1187 (N_1187,In_4275,In_2141);
and U1188 (N_1188,In_3480,In_240);
nor U1189 (N_1189,In_3959,N_84);
nor U1190 (N_1190,N_935,N_329);
xnor U1191 (N_1191,In_4263,In_3964);
or U1192 (N_1192,In_965,In_1981);
or U1193 (N_1193,In_1817,In_2283);
nor U1194 (N_1194,In_3054,In_4933);
and U1195 (N_1195,In_4670,In_505);
xor U1196 (N_1196,In_2559,In_1823);
nand U1197 (N_1197,In_915,In_2337);
nand U1198 (N_1198,In_2000,In_862);
xor U1199 (N_1199,In_2139,N_191);
and U1200 (N_1200,In_4546,In_4465);
nor U1201 (N_1201,In_413,In_4387);
or U1202 (N_1202,In_1838,In_1002);
nand U1203 (N_1203,In_1780,In_3146);
and U1204 (N_1204,In_4911,N_430);
nand U1205 (N_1205,N_428,In_4071);
and U1206 (N_1206,In_4375,In_4884);
or U1207 (N_1207,In_746,In_2979);
xnor U1208 (N_1208,In_3385,In_3966);
and U1209 (N_1209,In_2425,N_431);
and U1210 (N_1210,In_565,In_3287);
or U1211 (N_1211,In_4859,In_1487);
nor U1212 (N_1212,In_1652,In_1460);
xor U1213 (N_1213,In_1747,In_2479);
and U1214 (N_1214,In_1642,In_4410);
and U1215 (N_1215,In_3164,In_2306);
xor U1216 (N_1216,In_4793,In_2008);
or U1217 (N_1217,In_2962,In_3068);
nand U1218 (N_1218,In_3551,N_641);
xnor U1219 (N_1219,In_694,In_2612);
or U1220 (N_1220,In_4093,In_4225);
or U1221 (N_1221,In_166,N_975);
xor U1222 (N_1222,In_1136,N_196);
xnor U1223 (N_1223,In_3291,In_2165);
nor U1224 (N_1224,In_3503,N_631);
nor U1225 (N_1225,In_2707,In_2620);
or U1226 (N_1226,N_564,In_3260);
nand U1227 (N_1227,In_1852,In_2427);
xnor U1228 (N_1228,In_1544,In_4768);
xor U1229 (N_1229,In_1009,N_911);
nor U1230 (N_1230,N_970,N_44);
nor U1231 (N_1231,N_715,In_4778);
xor U1232 (N_1232,In_3428,In_4416);
nor U1233 (N_1233,In_4020,N_20);
and U1234 (N_1234,In_387,In_2996);
nor U1235 (N_1235,In_3822,N_904);
xor U1236 (N_1236,In_2522,In_2313);
xnor U1237 (N_1237,In_2892,In_3813);
or U1238 (N_1238,In_3556,In_2061);
nor U1239 (N_1239,In_632,In_2096);
and U1240 (N_1240,In_1775,In_465);
and U1241 (N_1241,N_579,In_3621);
xor U1242 (N_1242,In_3463,In_262);
and U1243 (N_1243,In_4481,In_395);
nor U1244 (N_1244,N_349,In_416);
nor U1245 (N_1245,N_603,In_2367);
or U1246 (N_1246,In_3601,In_4656);
xnor U1247 (N_1247,N_756,In_4639);
nand U1248 (N_1248,In_4017,In_3615);
nand U1249 (N_1249,In_168,N_351);
xor U1250 (N_1250,In_2151,In_4303);
nand U1251 (N_1251,In_2010,N_806);
xnor U1252 (N_1252,In_2976,In_171);
and U1253 (N_1253,In_3343,In_2478);
and U1254 (N_1254,N_674,In_4345);
xor U1255 (N_1255,In_3027,In_751);
nand U1256 (N_1256,In_4523,In_1073);
nor U1257 (N_1257,In_1014,In_1893);
xnor U1258 (N_1258,N_734,In_4824);
xnor U1259 (N_1259,In_4290,In_4683);
xnor U1260 (N_1260,In_1401,In_2985);
nand U1261 (N_1261,In_547,N_720);
or U1262 (N_1262,In_1887,N_40);
nor U1263 (N_1263,In_1862,In_3498);
nor U1264 (N_1264,In_1746,N_1047);
or U1265 (N_1265,N_71,N_925);
and U1266 (N_1266,In_2573,In_118);
nor U1267 (N_1267,In_805,In_2880);
xnor U1268 (N_1268,In_4873,N_414);
or U1269 (N_1269,In_4577,N_267);
xor U1270 (N_1270,In_1389,In_1663);
xor U1271 (N_1271,In_3262,N_649);
xnor U1272 (N_1272,N_1191,In_4091);
nand U1273 (N_1273,In_17,In_1673);
xor U1274 (N_1274,In_964,In_2767);
xnor U1275 (N_1275,In_1699,In_2049);
nor U1276 (N_1276,N_623,N_636);
xnor U1277 (N_1277,In_208,In_3281);
xnor U1278 (N_1278,In_2927,In_3865);
nand U1279 (N_1279,In_3909,In_1518);
or U1280 (N_1280,In_2879,In_2163);
nand U1281 (N_1281,In_2687,N_887);
and U1282 (N_1282,N_584,In_784);
or U1283 (N_1283,In_4734,N_69);
nor U1284 (N_1284,N_608,N_758);
or U1285 (N_1285,In_4376,In_4202);
nor U1286 (N_1286,In_736,N_672);
nand U1287 (N_1287,In_1995,N_169);
nand U1288 (N_1288,N_551,N_1005);
or U1289 (N_1289,N_670,In_2905);
or U1290 (N_1290,In_740,In_3933);
xnor U1291 (N_1291,N_1110,In_2135);
and U1292 (N_1292,In_4343,In_3233);
or U1293 (N_1293,In_3282,N_730);
nor U1294 (N_1294,In_4052,N_322);
nor U1295 (N_1295,In_546,In_3404);
xnor U1296 (N_1296,In_836,In_111);
and U1297 (N_1297,N_275,In_2420);
or U1298 (N_1298,In_1653,In_4647);
and U1299 (N_1299,N_1086,N_182);
and U1300 (N_1300,In_1547,In_4631);
nand U1301 (N_1301,In_75,N_1221);
nand U1302 (N_1302,In_1960,N_997);
and U1303 (N_1303,In_1925,In_366);
and U1304 (N_1304,In_3697,N_452);
xnor U1305 (N_1305,In_897,In_475);
and U1306 (N_1306,In_1368,N_807);
and U1307 (N_1307,In_3576,In_3916);
xor U1308 (N_1308,N_262,N_471);
and U1309 (N_1309,In_4092,In_1484);
xnor U1310 (N_1310,N_834,In_762);
or U1311 (N_1311,In_4746,In_4046);
nand U1312 (N_1312,N_398,In_4927);
xnor U1313 (N_1313,In_3833,In_4556);
xnor U1314 (N_1314,In_3553,In_1875);
nor U1315 (N_1315,N_190,In_3182);
and U1316 (N_1316,N_1192,N_299);
xor U1317 (N_1317,In_249,In_2734);
or U1318 (N_1318,N_1121,In_1363);
or U1319 (N_1319,In_1505,In_1751);
nor U1320 (N_1320,In_4964,In_4418);
or U1321 (N_1321,In_3753,N_779);
or U1322 (N_1322,N_478,In_2681);
or U1323 (N_1323,In_4507,In_643);
nand U1324 (N_1324,In_615,In_3118);
xor U1325 (N_1325,N_460,N_195);
xnor U1326 (N_1326,N_816,In_3181);
or U1327 (N_1327,In_1338,In_3861);
or U1328 (N_1328,In_3830,N_930);
nand U1329 (N_1329,N_264,N_982);
nand U1330 (N_1330,N_902,In_4660);
nor U1331 (N_1331,In_4178,In_2950);
nand U1332 (N_1332,In_1892,In_876);
or U1333 (N_1333,In_2002,In_1419);
and U1334 (N_1334,N_1101,N_785);
or U1335 (N_1335,In_4904,In_4220);
or U1336 (N_1336,N_1232,In_952);
nor U1337 (N_1337,N_780,In_139);
nor U1338 (N_1338,In_3377,In_3547);
xnor U1339 (N_1339,In_1431,In_4584);
xnor U1340 (N_1340,In_3400,In_2077);
xor U1341 (N_1341,In_4770,In_4752);
or U1342 (N_1342,In_875,In_2477);
nor U1343 (N_1343,In_2850,N_426);
nor U1344 (N_1344,In_2813,N_907);
xor U1345 (N_1345,In_4128,In_3872);
nand U1346 (N_1346,In_285,N_419);
nor U1347 (N_1347,In_3369,In_4205);
or U1348 (N_1348,In_2958,In_4406);
nand U1349 (N_1349,In_3045,In_1384);
and U1350 (N_1350,In_3436,N_306);
xnor U1351 (N_1351,In_1218,In_2429);
nor U1352 (N_1352,N_1237,In_2954);
xnor U1353 (N_1353,In_1407,In_4786);
xnor U1354 (N_1354,N_772,In_4645);
nand U1355 (N_1355,In_16,N_451);
nor U1356 (N_1356,N_122,N_356);
nor U1357 (N_1357,N_496,In_1219);
nand U1358 (N_1358,In_3572,In_1719);
nand U1359 (N_1359,In_3274,In_2484);
xnor U1360 (N_1360,N_1069,In_2069);
nor U1361 (N_1361,In_1233,In_4662);
xnor U1362 (N_1362,N_382,N_859);
nor U1363 (N_1363,N_273,In_4105);
nor U1364 (N_1364,N_959,In_1529);
nand U1365 (N_1365,In_866,In_1741);
and U1366 (N_1366,In_2308,In_1774);
and U1367 (N_1367,In_2947,In_1074);
and U1368 (N_1368,N_1236,In_4879);
nand U1369 (N_1369,In_3434,In_3405);
xor U1370 (N_1370,In_4658,In_4591);
or U1371 (N_1371,In_3032,In_4200);
or U1372 (N_1372,In_4278,N_531);
and U1373 (N_1373,In_3012,N_582);
nor U1374 (N_1374,In_633,In_2863);
xnor U1375 (N_1375,In_539,In_2417);
and U1376 (N_1376,In_2122,In_3718);
nor U1377 (N_1377,In_4065,In_3402);
nor U1378 (N_1378,In_3608,In_2538);
nand U1379 (N_1379,N_1091,In_254);
nand U1380 (N_1380,N_284,N_683);
xor U1381 (N_1381,N_784,In_3619);
xnor U1382 (N_1382,N_1152,In_3062);
nor U1383 (N_1383,In_282,N_1081);
and U1384 (N_1384,In_4187,In_2369);
nand U1385 (N_1385,N_894,N_280);
nand U1386 (N_1386,In_2917,In_3555);
nand U1387 (N_1387,In_3898,In_2838);
or U1388 (N_1388,In_443,N_265);
xnor U1389 (N_1389,In_2555,In_4459);
nand U1390 (N_1390,N_347,In_4374);
xnor U1391 (N_1391,N_543,In_2090);
nand U1392 (N_1392,In_1456,N_437);
nor U1393 (N_1393,N_1073,In_3738);
and U1394 (N_1394,In_3228,In_548);
and U1395 (N_1395,In_2459,In_908);
or U1396 (N_1396,In_1257,In_4805);
and U1397 (N_1397,In_333,N_918);
and U1398 (N_1398,In_1021,In_2750);
and U1399 (N_1399,N_1,N_560);
nor U1400 (N_1400,In_4155,N_1027);
or U1401 (N_1401,In_4744,In_4779);
nand U1402 (N_1402,N_1082,In_3095);
and U1403 (N_1403,In_2183,N_1033);
nand U1404 (N_1404,N_854,In_1851);
nor U1405 (N_1405,In_3424,N_103);
xor U1406 (N_1406,In_1472,In_4440);
nor U1407 (N_1407,In_4558,In_1605);
nor U1408 (N_1408,In_3953,In_2454);
nor U1409 (N_1409,In_3893,N_178);
or U1410 (N_1410,In_742,In_3000);
nand U1411 (N_1411,In_1215,In_2646);
and U1412 (N_1412,In_1564,In_4400);
nand U1413 (N_1413,N_651,N_818);
and U1414 (N_1414,N_787,N_1049);
nand U1415 (N_1415,In_2437,In_780);
nand U1416 (N_1416,In_2189,In_3368);
or U1417 (N_1417,In_4724,N_375);
or U1418 (N_1418,In_298,N_1200);
nand U1419 (N_1419,N_877,In_3448);
nor U1420 (N_1420,In_1376,N_288);
nor U1421 (N_1421,In_4679,In_1503);
or U1422 (N_1422,In_4311,In_1371);
nand U1423 (N_1423,In_12,In_4794);
nor U1424 (N_1424,In_556,In_1734);
and U1425 (N_1425,N_408,N_956);
or U1426 (N_1426,In_2982,In_535);
nor U1427 (N_1427,In_3674,In_2294);
and U1428 (N_1428,In_3079,In_1500);
nor U1429 (N_1429,N_404,In_3679);
nor U1430 (N_1430,In_4855,In_896);
xor U1431 (N_1431,In_3446,In_4837);
or U1432 (N_1432,N_90,N_1063);
and U1433 (N_1433,In_2988,N_1088);
nor U1434 (N_1434,In_2553,In_3801);
and U1435 (N_1435,N_873,In_1910);
nand U1436 (N_1436,In_371,In_3702);
and U1437 (N_1437,In_4337,N_1100);
nand U1438 (N_1438,N_762,In_4957);
and U1439 (N_1439,N_1019,In_3759);
nor U1440 (N_1440,In_2569,In_2193);
nor U1441 (N_1441,In_4945,N_1039);
nand U1442 (N_1442,In_1928,In_426);
xor U1443 (N_1443,In_2868,N_628);
nand U1444 (N_1444,In_4733,In_2462);
and U1445 (N_1445,In_4954,In_2410);
and U1446 (N_1446,In_2963,In_3917);
and U1447 (N_1447,N_1064,In_922);
xor U1448 (N_1448,In_1504,N_924);
and U1449 (N_1449,In_317,In_1173);
or U1450 (N_1450,In_2453,N_949);
or U1451 (N_1451,In_4528,In_3569);
and U1452 (N_1452,In_4950,In_2576);
nand U1453 (N_1453,In_326,In_348);
nand U1454 (N_1454,N_661,In_4672);
or U1455 (N_1455,N_598,In_1099);
xor U1456 (N_1456,In_3479,In_3981);
or U1457 (N_1457,In_3522,N_511);
nand U1458 (N_1458,In_2431,N_912);
or U1459 (N_1459,In_2605,In_3918);
and U1460 (N_1460,In_1064,In_2280);
xor U1461 (N_1461,In_1410,N_99);
and U1462 (N_1462,In_1263,N_621);
nand U1463 (N_1463,In_482,In_4878);
and U1464 (N_1464,N_750,In_4751);
or U1465 (N_1465,In_1836,N_1004);
or U1466 (N_1466,In_467,In_844);
nand U1467 (N_1467,In_1169,In_1471);
nand U1468 (N_1468,In_1927,In_3705);
nor U1469 (N_1469,In_2601,In_2239);
or U1470 (N_1470,N_376,In_545);
and U1471 (N_1471,In_3982,In_2321);
xor U1472 (N_1472,N_1035,In_1856);
or U1473 (N_1473,In_2399,In_2632);
and U1474 (N_1474,In_4059,In_1616);
nor U1475 (N_1475,In_4982,In_1773);
xnor U1476 (N_1476,N_68,In_2566);
and U1477 (N_1477,In_2177,In_4857);
and U1478 (N_1478,In_2434,In_1631);
nor U1479 (N_1479,In_3157,N_985);
nand U1480 (N_1480,N_713,In_203);
or U1481 (N_1481,N_642,N_453);
and U1482 (N_1482,In_3037,N_1111);
nor U1483 (N_1483,In_767,N_43);
xor U1484 (N_1484,N_1099,In_810);
or U1485 (N_1485,In_4663,In_1737);
or U1486 (N_1486,In_1158,In_541);
xor U1487 (N_1487,N_998,In_1147);
or U1488 (N_1488,N_1015,In_4763);
nand U1489 (N_1489,N_589,N_39);
xor U1490 (N_1490,In_586,In_4883);
nand U1491 (N_1491,In_1922,In_101);
xnor U1492 (N_1492,In_3337,In_464);
and U1493 (N_1493,In_648,N_922);
nand U1494 (N_1494,In_1831,In_4894);
and U1495 (N_1495,N_423,In_3358);
nand U1496 (N_1496,In_3837,In_3877);
and U1497 (N_1497,In_1019,In_1553);
xor U1498 (N_1498,N_987,In_4002);
nand U1499 (N_1499,N_687,In_1829);
nor U1500 (N_1500,In_4956,N_708);
nor U1501 (N_1501,In_4916,In_2795);
or U1502 (N_1502,N_1008,In_2741);
nor U1503 (N_1503,In_4913,In_4820);
nor U1504 (N_1504,In_2826,In_2347);
nor U1505 (N_1505,In_500,In_3869);
and U1506 (N_1506,In_2414,In_2247);
or U1507 (N_1507,In_390,In_3894);
nand U1508 (N_1508,In_709,N_882);
and U1509 (N_1509,In_15,In_373);
or U1510 (N_1510,In_187,N_1458);
or U1511 (N_1511,In_91,In_2334);
or U1512 (N_1512,In_613,In_1531);
xnor U1513 (N_1513,In_4094,In_974);
and U1514 (N_1514,In_3130,In_4413);
or U1515 (N_1515,In_2300,In_2718);
nor U1516 (N_1516,In_4051,N_695);
and U1517 (N_1517,In_4078,In_3060);
and U1518 (N_1518,In_812,In_1972);
nor U1519 (N_1519,In_1791,In_3474);
xor U1520 (N_1520,N_1087,In_4799);
nor U1521 (N_1521,In_1951,In_2004);
nand U1522 (N_1522,In_43,In_819);
nand U1523 (N_1523,N_348,In_63);
and U1524 (N_1524,In_808,In_64);
xnor U1525 (N_1525,N_962,N_1007);
nor U1526 (N_1526,In_2910,N_991);
xor U1527 (N_1527,N_1296,In_2037);
nand U1528 (N_1528,In_2398,In_4244);
nor U1529 (N_1529,N_1480,In_1592);
or U1530 (N_1530,In_1877,N_528);
and U1531 (N_1531,In_1770,In_2588);
and U1532 (N_1532,In_1348,In_1677);
or U1533 (N_1533,N_388,N_1363);
xnor U1534 (N_1534,In_1513,In_4480);
xor U1535 (N_1535,N_1057,In_2543);
nand U1536 (N_1536,In_3805,In_1405);
nand U1537 (N_1537,In_3955,N_549);
and U1538 (N_1538,N_1135,In_734);
and U1539 (N_1539,In_3218,In_708);
nand U1540 (N_1540,In_1826,In_344);
nand U1541 (N_1541,In_530,In_4924);
or U1542 (N_1542,In_4110,In_1830);
nor U1543 (N_1543,In_389,N_219);
or U1544 (N_1544,N_888,N_1465);
nor U1545 (N_1545,In_4227,In_4958);
xor U1546 (N_1546,N_662,In_3153);
nor U1547 (N_1547,In_838,N_744);
and U1548 (N_1548,In_3956,N_617);
or U1549 (N_1549,In_2581,In_961);
or U1550 (N_1550,In_2332,In_1819);
nand U1551 (N_1551,In_4922,In_2896);
nor U1552 (N_1552,In_419,In_572);
nor U1553 (N_1553,In_422,In_2664);
xor U1554 (N_1554,In_4388,In_809);
nand U1555 (N_1555,N_503,In_499);
nor U1556 (N_1556,N_1123,In_3566);
nand U1557 (N_1557,In_1991,In_1793);
or U1558 (N_1558,N_1256,In_1800);
nand U1559 (N_1559,In_4414,In_4520);
and U1560 (N_1560,In_456,In_4113);
xor U1561 (N_1561,N_739,In_2190);
xnor U1562 (N_1562,In_595,In_4201);
and U1563 (N_1563,In_631,In_2829);
xnor U1564 (N_1564,N_1290,N_574);
nand U1565 (N_1565,In_1096,N_1056);
xnor U1566 (N_1566,In_4449,N_72);
xor U1567 (N_1567,N_899,In_3831);
or U1568 (N_1568,In_4043,In_4608);
and U1569 (N_1569,In_4088,In_133);
and U1570 (N_1570,In_2181,N_718);
and U1571 (N_1571,In_2806,In_39);
and U1572 (N_1572,In_3256,N_303);
nand U1573 (N_1573,In_2908,N_1468);
or U1574 (N_1574,In_4814,In_3763);
and U1575 (N_1575,In_2645,N_1305);
xor U1576 (N_1576,In_1698,In_4455);
xor U1577 (N_1577,N_1387,In_3491);
nand U1578 (N_1578,N_934,In_800);
nand U1579 (N_1579,In_4640,In_162);
or U1580 (N_1580,In_3579,In_2527);
nor U1581 (N_1581,In_4946,In_947);
nor U1582 (N_1582,In_1336,In_3989);
nor U1583 (N_1583,N_1369,In_241);
nand U1584 (N_1584,N_868,N_947);
nand U1585 (N_1585,N_1077,N_222);
and U1586 (N_1586,In_145,N_981);
or U1587 (N_1587,In_2870,In_2871);
nand U1588 (N_1588,In_3071,In_4242);
xnor U1589 (N_1589,In_4731,In_4603);
nor U1590 (N_1590,In_929,In_174);
xnor U1591 (N_1591,In_4973,N_885);
or U1592 (N_1592,In_1199,In_1412);
nor U1593 (N_1593,In_2682,N_1445);
nand U1594 (N_1594,In_3093,In_1953);
and U1595 (N_1595,In_3582,In_817);
nand U1596 (N_1596,In_356,In_1098);
and U1597 (N_1597,In_4213,N_939);
xor U1598 (N_1598,In_53,N_958);
or U1599 (N_1599,In_4892,In_1046);
or U1600 (N_1600,In_4692,In_2027);
nor U1601 (N_1601,N_385,In_2014);
and U1602 (N_1602,N_875,N_401);
and U1603 (N_1603,In_1129,N_1247);
nand U1604 (N_1604,N_330,In_4164);
xnor U1605 (N_1605,N_619,In_3733);
xnor U1606 (N_1606,N_747,In_3150);
nand U1607 (N_1607,In_4889,In_1323);
and U1608 (N_1608,In_399,N_726);
xor U1609 (N_1609,In_1915,N_1125);
nor U1610 (N_1610,In_779,In_1440);
or U1611 (N_1611,N_1432,In_4816);
and U1612 (N_1612,In_79,In_2071);
xor U1613 (N_1613,In_2518,In_4462);
or U1614 (N_1614,In_3703,In_4714);
and U1615 (N_1615,N_1479,In_656);
nand U1616 (N_1616,N_548,N_133);
xor U1617 (N_1617,In_1267,In_2855);
or U1618 (N_1618,In_58,In_1248);
or U1619 (N_1619,In_2696,In_1204);
xnor U1620 (N_1620,N_851,In_4587);
and U1621 (N_1621,N_1395,In_3795);
nand U1622 (N_1622,N_847,In_4322);
nand U1623 (N_1623,N_855,In_2371);
nor U1624 (N_1624,In_503,In_2876);
and U1625 (N_1625,In_104,In_2835);
xnor U1626 (N_1626,N_1228,In_52);
xor U1627 (N_1627,In_3963,In_1322);
and U1628 (N_1628,In_2565,In_355);
nand U1629 (N_1629,In_4748,In_1558);
nand U1630 (N_1630,In_3828,In_2211);
xor U1631 (N_1631,N_705,N_1180);
xnor U1632 (N_1632,In_3991,N_943);
or U1633 (N_1633,In_2267,In_827);
and U1634 (N_1634,In_664,In_1485);
and U1635 (N_1635,In_4938,In_2204);
nor U1636 (N_1636,In_2660,In_502);
nor U1637 (N_1637,In_1816,In_2390);
and U1638 (N_1638,N_817,N_684);
or U1639 (N_1639,In_3812,In_3407);
nand U1640 (N_1640,In_4477,In_4545);
and U1641 (N_1641,N_542,N_164);
or U1642 (N_1642,N_1267,N_563);
nand U1643 (N_1643,In_4887,In_3954);
and U1644 (N_1644,In_1886,N_1373);
or U1645 (N_1645,In_2472,In_2480);
xor U1646 (N_1646,In_4787,In_2642);
nor U1647 (N_1647,In_295,N_1277);
and U1648 (N_1648,In_673,In_4968);
nor U1649 (N_1649,In_3500,N_283);
nand U1650 (N_1650,In_2081,In_2638);
or U1651 (N_1651,In_3379,In_2861);
or U1652 (N_1652,N_467,In_40);
or U1653 (N_1653,In_48,In_4089);
and U1654 (N_1654,In_4980,In_1081);
or U1655 (N_1655,In_2127,In_257);
nand U1656 (N_1656,N_197,In_3962);
and U1657 (N_1657,In_126,N_1020);
xor U1658 (N_1658,In_906,In_2184);
or U1659 (N_1659,N_737,In_978);
nor U1660 (N_1660,N_1052,In_2207);
nor U1661 (N_1661,In_2201,In_94);
xor U1662 (N_1662,N_664,In_1150);
and U1663 (N_1663,N_839,In_2017);
nand U1664 (N_1664,In_1429,N_1217);
or U1665 (N_1665,N_381,In_1481);
xnor U1666 (N_1666,In_4138,In_1971);
xnor U1667 (N_1667,N_274,N_1150);
xor U1668 (N_1668,In_3458,In_234);
nand U1669 (N_1669,In_4027,N_897);
or U1670 (N_1670,In_2078,In_1641);
xnor U1671 (N_1671,N_13,N_1367);
nor U1672 (N_1672,In_4228,In_3687);
or U1673 (N_1673,N_132,N_1476);
and U1674 (N_1674,In_4001,In_4720);
xor U1675 (N_1675,In_4674,N_643);
or U1676 (N_1676,N_1276,N_1219);
or U1677 (N_1677,In_3040,In_4436);
nand U1678 (N_1678,In_2285,N_315);
or U1679 (N_1679,In_2178,In_2965);
xor U1680 (N_1680,N_258,In_710);
or U1681 (N_1681,In_259,In_4609);
and U1682 (N_1682,In_2575,N_921);
xor U1683 (N_1683,In_2680,N_710);
nor U1684 (N_1684,In_408,In_3973);
nand U1685 (N_1685,In_3440,In_97);
and U1686 (N_1686,In_4013,In_2395);
and U1687 (N_1687,In_4784,N_1454);
xor U1688 (N_1688,In_129,In_1341);
xnor U1689 (N_1689,In_4131,In_383);
xnor U1690 (N_1690,In_2616,In_735);
nor U1691 (N_1691,In_4781,In_957);
and U1692 (N_1692,In_4643,N_1204);
nor U1693 (N_1693,In_971,N_782);
nor U1694 (N_1694,N_864,In_161);
nor U1695 (N_1695,N_754,In_1462);
and U1696 (N_1696,N_1157,In_3757);
nand U1697 (N_1697,In_2234,In_4022);
nand U1698 (N_1698,In_1465,In_1788);
or U1699 (N_1699,N_450,In_3976);
and U1700 (N_1700,N_876,N_1261);
nor U1701 (N_1701,In_4450,In_2042);
nand U1702 (N_1702,In_4194,N_1356);
xnor U1703 (N_1703,In_3824,In_198);
xnor U1704 (N_1704,In_1786,In_1911);
and U1705 (N_1705,N_1326,In_3396);
xor U1706 (N_1706,In_1192,In_3242);
nand U1707 (N_1707,N_163,In_1373);
and U1708 (N_1708,N_498,In_1254);
and U1709 (N_1709,N_1462,In_2611);
xor U1710 (N_1710,In_4425,In_4245);
or U1711 (N_1711,N_1120,N_1411);
xnor U1712 (N_1712,N_456,In_1738);
or U1713 (N_1713,In_4699,N_254);
xnor U1714 (N_1714,N_1271,In_3958);
nor U1715 (N_1715,In_202,In_2514);
nor U1716 (N_1716,In_2463,In_629);
nor U1717 (N_1717,N_1324,In_990);
and U1718 (N_1718,In_3145,N_1079);
nand U1719 (N_1719,In_3550,N_1364);
xor U1720 (N_1720,In_117,In_1045);
and U1721 (N_1721,N_495,In_749);
and U1722 (N_1722,In_2712,In_2287);
xnor U1723 (N_1723,N_325,In_801);
xor U1724 (N_1724,In_337,N_1097);
xor U1725 (N_1725,In_755,In_2360);
and U1726 (N_1726,N_1083,In_3965);
or U1727 (N_1727,In_1239,N_565);
nor U1728 (N_1728,N_1440,In_2476);
and U1729 (N_1729,In_607,In_4502);
nand U1730 (N_1730,In_4150,In_2117);
or U1731 (N_1731,In_3148,In_2270);
nor U1732 (N_1732,N_270,In_3719);
nand U1733 (N_1733,N_765,In_1557);
and U1734 (N_1734,In_4708,In_3578);
and U1735 (N_1735,In_4392,In_4974);
nand U1736 (N_1736,In_3823,In_2516);
or U1737 (N_1737,In_4062,In_2961);
nor U1738 (N_1738,In_1335,In_255);
or U1739 (N_1739,In_722,In_236);
nor U1740 (N_1740,In_1018,N_1456);
nand U1741 (N_1741,In_1613,In_4713);
nand U1742 (N_1742,In_3309,N_9);
and U1743 (N_1743,In_151,In_3739);
nor U1744 (N_1744,In_2460,N_1147);
or U1745 (N_1745,N_1330,In_3202);
xnor U1746 (N_1746,In_3533,In_2915);
nand U1747 (N_1747,In_4320,In_1194);
nand U1748 (N_1748,In_669,In_1644);
nand U1749 (N_1749,N_789,In_1208);
nor U1750 (N_1750,In_89,In_1909);
or U1751 (N_1751,In_3074,In_2801);
or U1752 (N_1752,In_158,In_3198);
or U1753 (N_1753,N_1422,In_1213);
nor U1754 (N_1754,N_1122,In_1387);
nor U1755 (N_1755,N_1318,In_2545);
or U1756 (N_1756,In_1964,In_2157);
nor U1757 (N_1757,In_3388,In_2326);
nor U1758 (N_1758,In_4496,In_1287);
xnor U1759 (N_1759,N_202,In_4342);
nor U1760 (N_1760,N_229,In_2033);
and U1761 (N_1761,N_94,N_1670);
and U1762 (N_1762,In_3243,N_1584);
nor U1763 (N_1763,In_2509,In_1655);
or U1764 (N_1764,N_1573,In_3429);
nor U1765 (N_1765,In_4864,In_3834);
nor U1766 (N_1766,N_1078,In_2594);
nor U1767 (N_1767,In_153,In_3864);
xor U1768 (N_1768,N_435,N_880);
or U1769 (N_1769,N_1613,N_1029);
and U1770 (N_1770,In_804,In_611);
xor U1771 (N_1771,In_4141,N_1225);
xnor U1772 (N_1772,In_1815,In_3272);
nand U1773 (N_1773,In_2029,In_1333);
xor U1774 (N_1774,In_2262,In_1707);
nand U1775 (N_1775,N_1569,In_3510);
and U1776 (N_1776,In_3597,In_1298);
nor U1777 (N_1777,N_294,In_4735);
nor U1778 (N_1778,In_1432,In_3356);
nand U1779 (N_1779,In_181,N_1663);
or U1780 (N_1780,In_2162,In_4581);
nor U1781 (N_1781,N_1710,In_690);
or U1782 (N_1782,N_1529,In_209);
xnor U1783 (N_1783,In_2966,N_1176);
xnor U1784 (N_1784,In_2883,In_3535);
nand U1785 (N_1785,N_399,In_4588);
nor U1786 (N_1786,In_4697,In_869);
and U1787 (N_1787,N_285,N_1708);
nand U1788 (N_1788,N_704,In_3773);
nand U1789 (N_1789,N_1715,N_974);
nor U1790 (N_1790,In_3570,N_1346);
nand U1791 (N_1791,In_2858,In_3821);
and U1792 (N_1792,N_1443,N_1341);
and U1793 (N_1793,N_1144,In_1142);
or U1794 (N_1794,N_886,In_1840);
nand U1795 (N_1795,In_351,In_4970);
xor U1796 (N_1796,N_732,N_1317);
nor U1797 (N_1797,N_1350,In_368);
xor U1798 (N_1798,In_3010,In_1646);
or U1799 (N_1799,In_3736,In_3540);
nor U1800 (N_1800,N_308,In_2142);
and U1801 (N_1801,In_2245,In_1686);
xnor U1802 (N_1802,N_1104,In_4920);
nand U1803 (N_1803,In_4401,N_1704);
or U1804 (N_1804,In_1409,In_4903);
and U1805 (N_1805,In_4230,In_3681);
and U1806 (N_1806,In_1276,N_1674);
and U1807 (N_1807,In_2574,In_1394);
xnor U1808 (N_1808,N_1664,N_682);
nor U1809 (N_1809,N_93,In_3058);
or U1810 (N_1810,In_3662,In_3649);
nor U1811 (N_1811,N_1351,In_4310);
xnor U1812 (N_1812,In_806,In_245);
nor U1813 (N_1813,In_3350,In_369);
xor U1814 (N_1814,N_722,N_1066);
and U1815 (N_1815,N_629,In_4586);
and U1816 (N_1816,N_1419,N_1705);
or U1817 (N_1817,N_1473,N_866);
and U1818 (N_1818,In_4162,In_2307);
and U1819 (N_1819,In_4655,N_903);
and U1820 (N_1820,In_1523,In_4505);
nor U1821 (N_1821,In_214,In_3005);
xnor U1822 (N_1822,N_1061,In_739);
nor U1823 (N_1823,N_1024,In_871);
nand U1824 (N_1824,In_159,N_143);
nand U1825 (N_1825,In_1537,N_999);
or U1826 (N_1826,In_4208,N_377);
nand U1827 (N_1827,N_920,In_7);
or U1828 (N_1828,In_445,In_4067);
or U1829 (N_1829,In_797,In_933);
and U1830 (N_1830,N_1382,N_1545);
nand U1831 (N_1831,In_2155,In_3647);
xor U1832 (N_1832,N_1489,In_454);
nand U1833 (N_1833,In_38,In_823);
nand U1834 (N_1834,N_48,In_3420);
nand U1835 (N_1835,In_3453,N_1178);
and U1836 (N_1836,N_1340,N_685);
nand U1837 (N_1837,N_438,In_1013);
nor U1838 (N_1838,In_1217,N_1484);
or U1839 (N_1839,In_1044,N_689);
and U1840 (N_1840,In_3710,In_3807);
nor U1841 (N_1841,In_3208,In_2886);
nand U1842 (N_1842,In_1224,In_4548);
and U1843 (N_1843,In_2418,N_333);
nand U1844 (N_1844,In_2624,N_1702);
nor U1845 (N_1845,N_1493,N_1628);
xor U1846 (N_1846,In_2152,In_3691);
xnor U1847 (N_1847,In_2537,N_320);
nand U1848 (N_1848,N_517,In_3713);
xnor U1849 (N_1849,In_4561,N_1734);
nor U1850 (N_1850,In_2690,In_959);
nor U1851 (N_1851,N_1726,N_1474);
xor U1852 (N_1852,In_2320,In_2137);
nand U1853 (N_1853,N_1140,In_2175);
or U1854 (N_1854,In_1015,N_1092);
or U1855 (N_1855,In_4955,In_637);
nand U1856 (N_1856,In_2727,In_4021);
xor U1857 (N_1857,N_334,In_2443);
xnor U1858 (N_1858,N_1719,In_1404);
or U1859 (N_1859,N_1263,In_2197);
and U1860 (N_1860,N_1423,In_4068);
nor U1861 (N_1861,N_554,N_1060);
nand U1862 (N_1862,N_1530,In_1201);
or U1863 (N_1863,In_2407,N_874);
nand U1864 (N_1864,N_961,In_4749);
or U1865 (N_1865,N_337,In_132);
xnor U1866 (N_1866,N_1441,N_218);
or U1867 (N_1867,In_3700,In_284);
nor U1868 (N_1868,N_232,In_4391);
xnor U1869 (N_1869,In_2445,N_251);
and U1870 (N_1870,In_753,In_2185);
xor U1871 (N_1871,In_652,N_1212);
and U1872 (N_1872,N_1642,In_2470);
nand U1873 (N_1873,N_1000,In_1235);
or U1874 (N_1874,In_788,In_1360);
or U1875 (N_1875,N_1610,N_697);
nand U1876 (N_1876,N_1618,N_455);
nor U1877 (N_1877,In_3289,In_2668);
nor U1878 (N_1878,In_22,N_1074);
nor U1879 (N_1879,In_424,In_521);
nor U1880 (N_1880,In_339,In_1402);
or U1881 (N_1881,In_1709,In_3626);
xor U1882 (N_1882,In_3870,N_1500);
nor U1883 (N_1883,In_2907,N_1535);
or U1884 (N_1884,N_1355,In_4267);
xor U1885 (N_1885,N_1321,N_449);
nand U1886 (N_1886,In_1568,N_443);
nor U1887 (N_1887,In_1128,N_136);
or U1888 (N_1888,In_2341,In_4404);
nand U1889 (N_1889,In_2544,In_4024);
and U1890 (N_1890,N_709,In_824);
xnor U1891 (N_1891,In_4207,In_1521);
and U1892 (N_1892,In_4076,N_19);
nand U1893 (N_1893,In_2794,In_1400);
nor U1894 (N_1894,N_1372,In_4039);
nor U1895 (N_1895,In_3015,In_2393);
xor U1896 (N_1896,In_2830,In_811);
xor U1897 (N_1897,In_2948,In_1516);
and U1898 (N_1898,In_2344,N_1392);
xor U1899 (N_1899,In_4149,N_1154);
or U1900 (N_1900,N_941,In_486);
and U1901 (N_1901,In_1339,In_4255);
nor U1902 (N_1902,In_582,N_10);
xor U1903 (N_1903,In_2380,N_1130);
or U1904 (N_1904,N_527,In_1532);
xor U1905 (N_1905,N_1510,In_1841);
xor U1906 (N_1906,N_2,In_2252);
or U1907 (N_1907,N_1711,In_4652);
or U1908 (N_1908,In_2312,N_266);
xor U1909 (N_1909,In_793,In_4972);
or U1910 (N_1910,In_2006,In_4248);
and U1911 (N_1911,N_64,N_520);
nand U1912 (N_1912,In_3539,In_216);
nand U1913 (N_1913,N_1665,N_429);
xnor U1914 (N_1914,In_100,In_2510);
nand U1915 (N_1915,In_942,In_1552);
and U1916 (N_1916,In_1247,N_1397);
nand U1917 (N_1917,In_3915,In_2062);
or U1918 (N_1918,N_1331,N_849);
xnor U1919 (N_1919,In_1079,N_78);
and U1920 (N_1920,In_4338,N_54);
and U1921 (N_1921,In_1858,In_923);
or U1922 (N_1922,In_2564,N_1170);
xor U1923 (N_1923,In_2799,N_1537);
or U1924 (N_1924,In_3033,In_4809);
nor U1925 (N_1925,In_1725,In_2202);
nor U1926 (N_1926,In_1229,N_871);
nor U1927 (N_1927,N_1524,In_2469);
xnor U1928 (N_1928,In_1181,In_4471);
nand U1929 (N_1929,In_3530,In_975);
xor U1930 (N_1930,In_4011,N_811);
nor U1931 (N_1931,N_1028,In_4403);
and U1932 (N_1932,In_296,N_835);
nor U1933 (N_1933,In_3900,In_1025);
nor U1934 (N_1934,N_1709,In_1052);
nand U1935 (N_1935,N_638,In_4849);
and U1936 (N_1936,N_669,N_759);
nor U1937 (N_1937,N_1687,N_569);
or U1938 (N_1938,In_1790,In_1942);
and U1939 (N_1939,In_604,In_88);
xnor U1940 (N_1940,In_1610,N_1173);
nor U1941 (N_1941,N_1379,N_1718);
nand U1942 (N_1942,In_175,N_1262);
nand U1943 (N_1943,N_633,N_1444);
nor U1944 (N_1944,In_3205,In_258);
nor U1945 (N_1945,In_1497,In_2831);
or U1946 (N_1946,N_594,N_1388);
or U1947 (N_1947,N_1103,In_1029);
nand U1948 (N_1948,N_415,In_4182);
nor U1949 (N_1949,In_2501,N_513);
nand U1950 (N_1950,In_2689,N_1025);
or U1951 (N_1951,In_3109,In_3694);
nor U1952 (N_1952,In_2919,In_1437);
and U1953 (N_1953,In_4184,In_4827);
or U1954 (N_1954,In_2773,N_1699);
nand U1955 (N_1955,In_3868,N_314);
or U1956 (N_1956,In_3331,N_1637);
nor U1957 (N_1957,N_1002,N_1084);
nor U1958 (N_1958,In_147,N_1427);
nor U1959 (N_1959,N_1332,N_1488);
and U1960 (N_1960,In_3373,In_2130);
nor U1961 (N_1961,In_3460,In_4902);
xnor U1962 (N_1962,In_1632,In_2043);
and U1963 (N_1963,In_1957,N_1311);
and U1964 (N_1964,N_1582,In_1885);
xnor U1965 (N_1965,In_3357,N_808);
or U1966 (N_1966,In_4308,In_3882);
nor U1967 (N_1967,In_19,In_998);
nor U1968 (N_1968,In_2654,N_1466);
xnor U1969 (N_1969,In_1130,N_1189);
or U1970 (N_1970,In_3107,In_848);
nor U1971 (N_1971,N_1329,N_908);
xor U1972 (N_1972,N_576,N_698);
and U1973 (N_1973,In_3907,N_394);
and U1974 (N_1974,In_1671,In_484);
nand U1975 (N_1975,In_4216,In_2521);
nand U1976 (N_1976,In_2409,In_3034);
xor U1977 (N_1977,In_2093,In_3351);
nor U1978 (N_1978,In_1753,N_424);
xnor U1979 (N_1979,In_4095,In_919);
nor U1980 (N_1980,N_1216,In_1769);
and U1981 (N_1981,N_63,In_4288);
nand U1982 (N_1982,N_606,In_851);
nand U1983 (N_1983,N_993,N_1309);
nor U1984 (N_1984,N_692,In_992);
nand U1985 (N_1985,N_733,In_4223);
nor U1986 (N_1986,In_4332,In_3061);
or U1987 (N_1987,In_1952,In_2999);
or U1988 (N_1988,In_2685,In_2461);
nor U1989 (N_1989,N_1713,N_1697);
nand U1990 (N_1990,In_1517,In_2805);
and U1991 (N_1991,N_843,In_4330);
xnor U1992 (N_1992,In_1849,In_901);
xor U1993 (N_1993,In_4636,In_36);
or U1994 (N_1994,N_712,In_375);
and U1995 (N_1995,In_1197,In_2606);
nand U1996 (N_1996,In_782,In_155);
and U1997 (N_1997,In_951,N_869);
and U1998 (N_1998,N_1273,N_1021);
and U1999 (N_1999,N_971,N_1010);
and U2000 (N_2000,N_5,In_2885);
xor U2001 (N_2001,In_3316,In_423);
xnor U2002 (N_2002,N_1617,N_1787);
nor U2003 (N_2003,N_1467,In_1377);
nand U2004 (N_2004,In_553,N_1587);
and U2005 (N_2005,N_1068,N_1620);
and U2006 (N_2006,N_18,N_176);
nand U2007 (N_2007,In_4295,In_4614);
nor U2008 (N_2008,N_1910,In_4723);
nand U2009 (N_2009,N_475,In_432);
nor U2010 (N_2010,N_1730,In_1206);
and U2011 (N_2011,In_4423,N_1365);
nand U2012 (N_2012,In_4522,In_1004);
nand U2013 (N_2013,In_4452,N_1720);
or U2014 (N_2014,In_3904,In_4284);
or U2015 (N_2015,In_4133,In_3643);
and U2016 (N_2016,In_4265,N_1789);
nor U2017 (N_2017,In_2535,N_1956);
or U2018 (N_2018,N_159,In_2174);
or U2019 (N_2019,N_767,In_2924);
xnor U2020 (N_2020,In_1442,N_946);
or U2021 (N_2021,N_1193,In_2170);
xnor U2022 (N_2022,In_4151,In_4293);
or U2023 (N_2023,In_1837,In_1083);
nor U2024 (N_2024,In_3548,N_1418);
nand U2025 (N_2025,In_4009,In_2570);
and U2026 (N_2026,N_1538,In_726);
nand U2027 (N_2027,In_2651,In_3986);
and U2028 (N_2028,In_4286,In_405);
and U2029 (N_2029,In_4576,In_3788);
xnor U2030 (N_2030,N_1421,In_4018);
nor U2031 (N_2031,In_4853,In_3220);
nand U2032 (N_2032,In_704,N_1881);
or U2033 (N_2033,In_195,N_1732);
nor U2034 (N_2034,In_2233,In_3814);
nand U2035 (N_2035,N_1149,In_4210);
xnor U2036 (N_2036,In_2322,N_1565);
xor U2037 (N_2037,In_4648,In_1433);
nand U2038 (N_2038,In_3596,In_1326);
nand U2039 (N_2039,N_1371,In_352);
nand U2040 (N_2040,N_578,N_1391);
and U2041 (N_2041,In_1944,In_4315);
xnor U2042 (N_2042,In_1222,In_3372);
or U2043 (N_2043,N_1594,In_1978);
xnor U2044 (N_2044,In_4677,In_4268);
nor U2045 (N_2045,In_667,In_3568);
xnor U2046 (N_2046,N_1878,In_4007);
xor U2047 (N_2047,N_778,In_681);
nand U2048 (N_2048,N_1017,In_1705);
xnor U2049 (N_2049,N_1447,In_1066);
nand U2050 (N_2050,In_156,N_1794);
xor U2051 (N_2051,N_290,In_4689);
nand U2052 (N_2052,In_4797,In_2475);
or U2053 (N_2053,N_1724,N_1126);
xnor U2054 (N_2054,N_538,In_3999);
nor U2055 (N_2055,N_509,In_4429);
or U2056 (N_2056,In_596,In_2064);
xnor U2057 (N_2057,N_1716,In_4079);
and U2058 (N_2058,N_1823,In_1156);
nor U2059 (N_2059,In_859,In_65);
or U2060 (N_2060,In_4871,In_3346);
nand U2061 (N_2061,N_1835,N_505);
nand U2062 (N_2062,In_2824,N_1522);
nor U2063 (N_2063,N_716,In_744);
nor U2064 (N_2064,In_1996,In_4650);
nor U2065 (N_2065,N_1568,N_1376);
or U2066 (N_2066,N_1205,N_162);
nand U2067 (N_2067,N_1666,N_898);
and U2068 (N_2068,In_4120,In_340);
or U2069 (N_2069,In_542,In_3375);
or U2070 (N_2070,In_3389,In_1027);
and U2071 (N_2071,N_1127,N_514);
and U2072 (N_2072,N_1668,N_1314);
nor U2073 (N_2073,In_3887,N_819);
nor U2074 (N_2074,In_1969,In_1522);
xor U2075 (N_2075,In_2396,N_865);
or U2076 (N_2076,N_441,N_1765);
and U2077 (N_2077,In_3306,In_3908);
or U2078 (N_2078,In_4281,N_593);
nor U2079 (N_2079,In_2094,In_4754);
nand U2080 (N_2080,In_2442,In_2084);
nor U2081 (N_2081,N_1541,In_2761);
or U2082 (N_2082,N_1478,N_1051);
nor U2083 (N_2083,In_3977,In_1510);
nor U2084 (N_2084,N_1399,In_4798);
nor U2085 (N_2085,N_1023,N_331);
nand U2086 (N_2086,In_750,In_3213);
nand U2087 (N_2087,N_126,In_3914);
or U2088 (N_2088,In_3564,In_494);
or U2089 (N_2089,In_3675,N_812);
xnor U2090 (N_2090,In_1495,In_1543);
xor U2091 (N_2091,N_1775,In_2293);
or U2092 (N_2092,In_3935,In_963);
or U2093 (N_2093,In_1258,In_2353);
and U2094 (N_2094,In_981,In_691);
xor U2095 (N_2095,N_1293,N_1743);
nand U2096 (N_2096,In_1912,In_1528);
nand U2097 (N_2097,N_1160,In_323);
nand U2098 (N_2098,In_924,N_1093);
and U2099 (N_2099,N_801,In_4563);
or U2100 (N_2100,N_1335,In_3475);
or U2101 (N_2101,N_893,N_650);
or U2102 (N_2102,N_1935,In_1149);
nor U2103 (N_2103,N_482,In_2473);
and U2104 (N_2104,In_966,In_531);
and U2105 (N_2105,N_422,N_74);
or U2106 (N_2106,In_3970,In_3445);
and U2107 (N_2107,N_1624,In_2526);
or U2108 (N_2108,In_522,In_3293);
xor U2109 (N_2109,N_358,In_429);
xnor U2110 (N_2110,In_3844,N_116);
xnor U2111 (N_2111,In_191,N_1424);
nand U2112 (N_2112,N_361,N_1675);
xor U2113 (N_2113,N_493,In_4721);
and U2114 (N_2114,In_1396,N_485);
xnor U2115 (N_2115,In_31,N_1768);
nand U2116 (N_2116,N_1779,In_1325);
xnor U2117 (N_2117,N_830,In_3473);
xnor U2118 (N_2118,N_1143,In_3880);
nor U2119 (N_2119,N_749,N_1851);
nor U2120 (N_2120,In_614,In_2298);
nand U2121 (N_2121,In_33,In_4678);
nor U2122 (N_2122,In_3741,N_1544);
or U2123 (N_2123,N_1873,In_4926);
nor U2124 (N_2124,N_1991,In_1574);
nand U2125 (N_2125,In_452,N_1655);
and U2126 (N_2126,In_9,In_2057);
or U2127 (N_2127,In_2179,In_4334);
xor U2128 (N_2128,In_1882,In_450);
nand U2129 (N_2129,N_1942,In_1042);
and U2130 (N_2130,N_1133,In_4434);
nor U2131 (N_2131,In_2972,N_409);
and U2132 (N_2132,N_1600,N_1059);
xor U2133 (N_2133,In_1038,N_699);
and U2134 (N_2134,In_879,N_1893);
xor U2135 (N_2135,N_454,In_2022);
xnor U2136 (N_2136,N_439,N_691);
xor U2137 (N_2137,In_1869,N_614);
xnor U2138 (N_2138,In_3135,In_820);
nand U2139 (N_2139,N_462,N_1377);
nand U2140 (N_2140,N_963,N_829);
nor U2141 (N_2141,In_4668,N_1689);
and U2142 (N_2142,In_2709,In_4253);
nor U2143 (N_2143,In_4402,In_3300);
nand U2144 (N_2144,N_224,In_403);
nor U2145 (N_2145,In_1501,In_2250);
nand U2146 (N_2146,In_4066,In_2729);
xor U2147 (N_2147,In_4893,N_508);
and U2148 (N_2148,In_783,N_1174);
and U2149 (N_2149,In_51,In_2899);
nand U2150 (N_2150,N_1515,N_55);
and U2151 (N_2151,In_2980,N_1889);
nor U2152 (N_2152,N_1707,N_277);
and U2153 (N_2153,In_3784,In_311);
xnor U2154 (N_2154,N_1673,In_2382);
nand U2155 (N_2155,In_4989,N_1245);
or U2156 (N_2156,N_1862,In_1580);
nand U2157 (N_2157,N_279,N_1137);
nand U2158 (N_2158,In_2147,In_27);
nand U2159 (N_2159,In_2264,N_11);
nand U2160 (N_2160,In_874,N_1869);
nor U2161 (N_2161,In_1674,N_966);
nor U2162 (N_2162,N_856,N_1536);
nand U2163 (N_2163,N_1605,In_543);
xor U2164 (N_2164,In_839,In_2241);
or U2165 (N_2165,N_933,In_4005);
nor U2166 (N_2166,In_4566,N_317);
xor U2167 (N_2167,In_1255,N_1162);
or U2168 (N_2168,N_1721,In_654);
nor U2169 (N_2169,N_1660,N_1990);
xnor U2170 (N_2170,In_3336,In_3634);
nand U2171 (N_2171,In_4397,N_1250);
nor U2172 (N_2172,In_1721,In_3158);
or U2173 (N_2173,In_3041,In_4132);
nand U2174 (N_2174,N_1795,In_4249);
and U2175 (N_2175,In_3745,N_1109);
nand U2176 (N_2176,In_1022,In_2082);
and U2177 (N_2177,In_774,In_2659);
xnor U2178 (N_2178,In_3100,In_4483);
and U2179 (N_2179,In_645,In_2595);
xnor U2180 (N_2180,In_2787,In_3009);
xor U2181 (N_2181,In_4569,N_1280);
and U2182 (N_2182,In_4129,N_1849);
and U2183 (N_2183,N_1227,In_1382);
and U2184 (N_2184,In_1718,In_2263);
or U2185 (N_2185,N_984,In_1061);
xnor U2186 (N_2186,N_1616,In_1621);
nand U2187 (N_2187,In_2629,In_314);
xnor U2188 (N_2188,In_3264,In_3827);
or U2189 (N_2189,N_1799,N_1988);
and U2190 (N_2190,N_1353,In_2089);
nand U2191 (N_2191,N_1264,In_2793);
and U2192 (N_2192,In_3200,N_1791);
nand U2193 (N_2193,In_1463,In_1845);
and U2194 (N_2194,N_1701,In_2598);
nor U2195 (N_2195,In_3307,In_4757);
nand U2196 (N_2196,In_1448,In_4995);
xor U2197 (N_2197,N_992,N_1409);
or U2198 (N_2198,N_1685,N_663);
nor U2199 (N_2199,In_1264,In_287);
or U2200 (N_2200,N_1759,N_1425);
and U2201 (N_2201,N_1603,In_1380);
nand U2202 (N_2202,N_1442,In_3932);
nand U2203 (N_2203,N_1901,In_969);
nor U2204 (N_2204,N_1776,In_418);
or U2205 (N_2205,In_226,In_1040);
xor U2206 (N_2206,In_459,In_2577);
or U2207 (N_2207,In_4233,N_463);
or U2208 (N_2208,N_480,In_1689);
or U2209 (N_2209,N_289,In_1047);
nand U2210 (N_2210,In_1492,In_6);
nor U2211 (N_2211,In_4966,In_4727);
nor U2212 (N_2212,In_4574,N_1076);
or U2213 (N_2213,N_1001,N_1645);
or U2214 (N_2214,N_1923,In_1620);
nand U2215 (N_2215,In_324,In_649);
or U2216 (N_2216,N_1184,N_268);
and U2217 (N_2217,N_226,N_1780);
and U2218 (N_2218,In_1273,In_2798);
nor U2219 (N_2219,N_1338,In_143);
nand U2220 (N_2220,N_1548,In_2528);
nand U2221 (N_2221,In_945,In_1643);
or U2222 (N_2222,In_785,N_1815);
nand U2223 (N_2223,In_2627,In_1383);
or U2224 (N_2224,N_1096,In_1065);
nor U2225 (N_2225,N_878,N_1837);
xor U2226 (N_2226,In_2539,In_3538);
nand U2227 (N_2227,N_1022,In_3672);
nor U2228 (N_2228,N_1735,N_1906);
or U2229 (N_2229,In_1593,N_929);
nand U2230 (N_2230,In_3188,N_1850);
nand U2231 (N_2231,N_1268,In_4984);
or U2232 (N_2232,In_4000,In_1346);
or U2233 (N_2233,In_3644,In_4909);
nor U2234 (N_2234,In_2758,N_489);
or U2235 (N_2235,N_46,In_277);
xnor U2236 (N_2236,In_2324,N_1009);
or U2237 (N_2237,N_1816,In_346);
nand U2238 (N_2238,In_193,N_1611);
nor U2239 (N_2239,In_3160,N_901);
nor U2240 (N_2240,In_4010,N_1623);
nand U2241 (N_2241,N_1972,In_4236);
nand U2242 (N_2242,N_1985,In_4145);
and U2243 (N_2243,N_666,In_2788);
xnor U2244 (N_2244,In_1662,In_4321);
or U2245 (N_2245,In_4537,In_1011);
nor U2246 (N_2246,In_2075,In_1372);
nor U2247 (N_2247,In_3310,In_3818);
nand U2248 (N_2248,N_1667,N_1134);
or U2249 (N_2249,N_1811,In_457);
nand U2250 (N_2250,In_215,N_2123);
xnor U2251 (N_2251,In_400,N_824);
or U2252 (N_2252,N_2187,N_724);
xor U2253 (N_2253,In_2464,N_1984);
nor U2254 (N_2254,N_2234,In_3590);
and U2255 (N_2255,N_2153,In_4716);
xor U2256 (N_2256,N_1983,N_1576);
nor U2257 (N_2257,N_1857,N_442);
nor U2258 (N_2258,N_1297,In_481);
or U2259 (N_2259,In_347,N_555);
nand U2260 (N_2260,In_244,In_3432);
nand U2261 (N_2261,N_986,In_1453);
and U2262 (N_2262,N_813,N_1880);
xor U2263 (N_2263,In_832,In_4952);
xnor U2264 (N_2264,In_470,N_1578);
nand U2265 (N_2265,In_3820,N_1528);
xor U2266 (N_2266,N_1533,In_1533);
nor U2267 (N_2267,In_3490,In_1679);
nand U2268 (N_2268,In_2386,N_2232);
nand U2269 (N_2269,N_1997,In_989);
xnor U2270 (N_2270,N_1847,In_1399);
and U2271 (N_2271,In_4725,N_2173);
xor U2272 (N_2272,N_1041,N_1951);
nor U2273 (N_2273,N_1343,N_1328);
nor U2274 (N_2274,N_2008,N_1358);
and U2275 (N_2275,N_2219,In_396);
nand U2276 (N_2276,N_916,N_1295);
nand U2277 (N_2277,In_2377,N_1195);
or U2278 (N_2278,In_1595,N_1824);
or U2279 (N_2279,N_1453,N_2048);
and U2280 (N_2280,N_1949,In_3064);
nand U2281 (N_2281,In_4214,In_4832);
nand U2282 (N_2282,N_1661,N_1599);
xnor U2283 (N_2283,N_2087,N_365);
or U2284 (N_2284,In_1259,N_1339);
xor U2285 (N_2285,N_1532,In_173);
xor U2286 (N_2286,In_2894,N_541);
or U2287 (N_2287,In_2144,In_2026);
xnor U2288 (N_2288,N_2097,N_1451);
xnor U2289 (N_2289,In_157,In_1832);
and U2290 (N_2290,N_675,N_146);
nand U2291 (N_2291,N_2070,In_2100);
or U2292 (N_2292,N_2143,In_2778);
xnor U2293 (N_2293,N_1491,N_1897);
or U2294 (N_2294,N_828,In_2362);
xnor U2295 (N_2295,N_852,In_3044);
xor U2296 (N_2296,N_1690,In_1220);
or U2297 (N_2297,In_367,In_3303);
xor U2298 (N_2298,In_4685,In_4054);
xnor U2299 (N_2299,In_1651,In_1874);
or U2300 (N_2300,N_76,In_3727);
and U2301 (N_2301,N_1106,In_3489);
nand U2302 (N_2302,In_3184,In_3961);
or U2303 (N_2303,N_2222,In_4466);
nand U2304 (N_2304,In_3020,N_1769);
and U2305 (N_2305,In_4620,N_1040);
or U2306 (N_2306,In_1853,In_4532);
or U2307 (N_2307,N_1527,N_815);
and U2308 (N_2308,N_1531,In_3663);
nand U2309 (N_2309,N_2177,N_2184);
xor U2310 (N_2310,In_4842,N_1773);
xnor U2311 (N_2311,N_2108,In_2608);
xnor U2312 (N_2312,In_4042,In_2630);
or U2313 (N_2313,N_327,In_2672);
and U2314 (N_2314,N_525,N_2171);
and U2315 (N_2315,In_864,In_2693);
nor U2316 (N_2316,N_2146,In_306);
and U2317 (N_2317,N_556,In_3849);
xor U2318 (N_2318,In_3328,In_2230);
xnor U2319 (N_2319,N_1113,In_878);
xor U2320 (N_2320,In_440,In_3632);
nand U2321 (N_2321,In_398,In_3544);
and U2322 (N_2322,N_1498,In_2511);
or U2323 (N_2323,N_721,N_1782);
and U2324 (N_2324,In_163,N_1551);
nand U2325 (N_2325,In_3599,N_2026);
and U2326 (N_2326,In_3091,N_1016);
xor U2327 (N_2327,N_1762,N_1833);
nand U2328 (N_2328,N_1828,In_3957);
nor U2329 (N_2329,N_1175,In_3614);
or U2330 (N_2330,N_114,In_3725);
xnor U2331 (N_2331,In_1665,N_2055);
or U2332 (N_2332,N_1928,N_599);
nor U2333 (N_2333,N_1598,In_3685);
xnor U2334 (N_2334,In_4323,N_1284);
xnor U2335 (N_2335,N_1654,In_3066);
and U2336 (N_2336,In_1562,In_1160);
or U2337 (N_2337,In_646,In_2435);
and U2338 (N_2338,In_20,In_2549);
and U2339 (N_2339,In_2392,In_3874);
and U2340 (N_2340,N_490,N_2032);
nand U2341 (N_2341,N_1754,N_2061);
xor U2342 (N_2342,In_1152,N_1609);
nor U2343 (N_2343,N_1146,In_3214);
and U2344 (N_2344,In_3105,N_1867);
nand U2345 (N_2345,N_1970,In_651);
xor U2346 (N_2346,In_684,In_2023);
nor U2347 (N_2347,N_1543,N_2229);
or U2348 (N_2348,N_1316,N_2021);
nor U2349 (N_2349,In_123,In_3693);
and U2350 (N_2350,N_2084,N_1258);
or U2351 (N_2351,In_394,N_1738);
and U2352 (N_2352,In_2047,N_831);
nand U2353 (N_2353,N_1472,N_1336);
and U2354 (N_2354,In_3670,N_89);
nor U2355 (N_2355,N_1511,In_2763);
and U2356 (N_2356,N_725,N_1575);
xor U2357 (N_2357,N_1981,N_844);
and U2358 (N_2358,In_1211,N_1403);
xor U2359 (N_2359,N_2192,In_1970);
nand U2360 (N_2360,In_4298,In_1035);
nor U2361 (N_2361,In_3843,N_1207);
nand U2362 (N_2362,In_4382,N_2172);
nor U2363 (N_2363,N_2038,In_2936);
and U2364 (N_2364,N_2201,In_2275);
or U2365 (N_2365,In_4831,In_3094);
or U2366 (N_2366,N_2209,N_1481);
and U2367 (N_2367,N_906,In_2803);
or U2368 (N_2368,In_3422,In_1017);
nand U2369 (N_2369,N_1393,In_2626);
xnor U2370 (N_2370,N_371,In_3353);
nand U2371 (N_2371,N_2122,N_1574);
xnor U2372 (N_2372,N_1220,N_1477);
or U2373 (N_2373,N_2121,In_4237);
xnor U2374 (N_2374,In_1496,N_129);
and U2375 (N_2375,In_239,In_4541);
or U2376 (N_2376,N_558,In_4788);
nand U2377 (N_2377,In_228,In_4123);
or U2378 (N_2378,In_3695,In_3571);
or U2379 (N_2379,N_2024,In_283);
nand U2380 (N_2380,N_45,N_1546);
or U2381 (N_2381,N_1877,In_2058);
nor U2382 (N_2382,N_2004,In_4705);
xnor U2383 (N_2383,In_90,In_3862);
nor U2384 (N_2384,N_2202,In_2774);
xnor U2385 (N_2385,In_2076,N_1888);
and U2386 (N_2386,N_976,In_672);
nand U2387 (N_2387,N_736,In_4259);
nand U2388 (N_2388,In_776,In_2561);
or U2389 (N_2389,In_137,In_1231);
nor U2390 (N_2390,N_1745,In_3790);
nor U2391 (N_2391,In_2359,In_2034);
and U2392 (N_2392,N_1883,N_1459);
nand U2393 (N_2393,In_4567,In_1639);
and U2394 (N_2394,N_2203,N_776);
and U2395 (N_2395,In_1113,N_2248);
nand U2396 (N_2396,N_2088,N_648);
nor U2397 (N_2397,N_2134,N_1234);
or U2398 (N_2398,N_928,In_1250);
nor U2399 (N_2399,In_2881,N_793);
nand U2400 (N_2400,In_4841,In_2586);
nand U2401 (N_2401,N_1672,In_2110);
or U2402 (N_2402,N_1875,In_3481);
nor U2403 (N_2403,In_2079,N_359);
xor U2404 (N_2404,In_4821,In_359);
nor U2405 (N_2405,N_1941,N_1764);
or U2406 (N_2406,N_53,In_3273);
nand U2407 (N_2407,N_1252,N_753);
xnor U2408 (N_2408,In_1587,N_1072);
nor U2409 (N_2409,In_3890,In_4525);
nand U2410 (N_2410,N_1119,In_95);
nor U2411 (N_2411,In_3838,N_2112);
xor U2412 (N_2412,In_2333,In_1491);
and U2413 (N_2413,N_858,In_4351);
xnor U2414 (N_2414,N_702,In_148);
and U2415 (N_2415,In_4969,N_1408);
xnor U2416 (N_2416,In_1330,N_1118);
xnor U2417 (N_2417,N_1523,In_2266);
xnor U2418 (N_2418,In_720,N_905);
xnor U2419 (N_2419,N_1727,In_4869);
nand U2420 (N_2420,N_2168,In_11);
nor U2421 (N_2421,In_2255,In_47);
or U2422 (N_2422,N_676,N_1512);
and U2423 (N_2423,N_1308,In_2244);
or U2424 (N_2424,In_1006,In_3521);
nor U2425 (N_2425,N_1037,In_365);
and U2426 (N_2426,N_2116,In_4359);
xnor U2427 (N_2427,N_1918,N_2170);
or U2428 (N_2428,In_4729,In_1174);
xnor U2429 (N_2429,In_4063,N_1402);
nand U2430 (N_2430,In_3848,N_570);
nor U2431 (N_2431,In_2074,N_1139);
and U2432 (N_2432,N_1344,In_3802);
and U2433 (N_2433,In_1155,N_1361);
xnor U2434 (N_2434,N_1567,In_4632);
nand U2435 (N_2435,In_1889,In_520);
nor U2436 (N_2436,In_3543,In_4560);
nand U2437 (N_2437,N_1525,In_3013);
xnor U2438 (N_2438,N_2120,In_4377);
or U2439 (N_2439,In_860,In_3240);
xor U2440 (N_2440,N_626,N_1313);
nor U2441 (N_2441,In_4527,In_1614);
nand U2442 (N_2442,N_2125,In_2974);
or U2443 (N_2443,N_964,N_1583);
xor U2444 (N_2444,In_3090,In_1093);
nor U2445 (N_2445,N_1846,In_3806);
or U2446 (N_2446,N_1766,N_515);
or U2447 (N_2447,In_1787,In_3913);
or U2448 (N_2448,In_4978,N_1706);
and U2449 (N_2449,In_4188,In_4003);
or U2450 (N_2450,In_3323,In_4073);
nand U2451 (N_2451,In_1962,In_4979);
or U2452 (N_2452,In_4498,In_2494);
and U2453 (N_2453,In_308,N_616);
or U2454 (N_2454,N_1579,In_3123);
and U2455 (N_2455,N_1429,In_4183);
and U2456 (N_2456,N_680,In_3278);
or U2457 (N_2457,N_1171,N_1644);
nor U2458 (N_2458,N_1534,N_2011);
nor U2459 (N_2459,N_343,In_1597);
and U2460 (N_2460,In_2242,In_3768);
nor U2461 (N_2461,N_1763,In_292);
nand U2462 (N_2462,N_363,N_1181);
or U2463 (N_2463,In_2558,In_1058);
nor U2464 (N_2464,N_1978,In_4257);
or U2465 (N_2465,In_3654,N_357);
or U2466 (N_2466,In_4745,N_927);
xor U2467 (N_2467,In_4941,N_1166);
nand U2468 (N_2468,N_1265,N_134);
nor U2469 (N_2469,N_180,In_309);
nor U2470 (N_2470,N_957,N_281);
nand U2471 (N_2471,In_3863,In_4638);
or U2472 (N_2472,N_117,In_2060);
xnor U2473 (N_2473,In_453,In_3780);
xnor U2474 (N_2474,In_4096,N_1861);
or U2475 (N_2475,In_1733,N_1937);
or U2476 (N_2476,N_128,N_521);
nand U2477 (N_2477,N_1963,In_3047);
and U2478 (N_2478,In_4196,In_2114);
nand U2479 (N_2479,In_2401,In_2123);
and U2480 (N_2480,In_593,In_2932);
xor U2481 (N_2481,In_1551,In_1278);
or U2482 (N_2482,N_1571,N_2179);
or U2483 (N_2483,N_2092,N_1416);
xnor U2484 (N_2484,In_3,N_30);
and U2485 (N_2485,In_2087,N_120);
nor U2486 (N_2486,N_2195,In_2897);
xor U2487 (N_2487,N_1882,N_436);
or U2488 (N_2488,N_1231,N_660);
nor U2489 (N_2489,In_72,In_4139);
nor U2490 (N_2490,In_2957,N_38);
xnor U2491 (N_2491,N_2137,In_2918);
nor U2492 (N_2492,N_936,N_1018);
nor U2493 (N_2493,In_3980,In_3960);
xnor U2494 (N_2494,In_4348,In_3067);
or U2495 (N_2495,In_2108,In_1636);
xnor U2496 (N_2496,N_123,N_1482);
nor U2497 (N_2497,N_1299,In_455);
xor U2498 (N_2498,In_689,In_638);
nand U2499 (N_2499,In_584,In_362);
xor U2500 (N_2500,In_1779,N_1368);
and U2501 (N_2501,N_1053,N_2188);
nor U2502 (N_2502,In_2939,In_4743);
nor U2503 (N_2503,In_679,N_1044);
nand U2504 (N_2504,In_1810,In_4739);
nor U2505 (N_2505,N_1517,N_639);
or U2506 (N_2506,N_814,In_914);
xor U2507 (N_2507,In_2505,In_557);
nand U2508 (N_2508,N_1916,In_4783);
or U2509 (N_2509,N_7,In_149);
nand U2510 (N_2510,In_1037,N_187);
nand U2511 (N_2511,N_596,N_87);
and U2512 (N_2512,In_2329,In_4573);
xnor U2513 (N_2513,N_1407,In_999);
nor U2514 (N_2514,In_1319,N_2326);
or U2515 (N_2515,In_4158,In_2228);
nor U2516 (N_2516,N_1912,In_4175);
and U2517 (N_2517,In_918,In_3523);
nand U2518 (N_2518,In_1907,In_4667);
and U2519 (N_2519,In_2740,N_770);
or U2520 (N_2520,N_840,N_2364);
nand U2521 (N_2521,In_2929,N_1412);
nor U2522 (N_2522,In_1710,N_1504);
or U2523 (N_2523,N_1805,N_2243);
and U2524 (N_2524,N_795,N_1404);
xor U2525 (N_2525,N_2066,In_1439);
and U2526 (N_2526,In_714,N_2271);
nand U2527 (N_2527,In_3927,N_572);
or U2528 (N_2528,N_2311,N_2225);
or U2529 (N_2529,N_1542,In_1084);
nand U2530 (N_2530,In_1899,N_755);
and U2531 (N_2531,In_2169,In_997);
nand U2532 (N_2532,N_1975,N_2036);
nand U2533 (N_2533,In_3689,In_2028);
or U2534 (N_2534,In_715,In_354);
nor U2535 (N_2535,N_212,N_1834);
nand U2536 (N_2536,In_3088,N_979);
nand U2537 (N_2537,In_1238,N_104);
and U2538 (N_2538,In_3984,In_1701);
nand U2539 (N_2539,N_1807,In_4530);
xnor U2540 (N_2540,N_791,In_3815);
nor U2541 (N_2541,In_1825,In_4940);
nor U2542 (N_2542,N_1908,In_1727);
or U2543 (N_2543,In_1820,In_4890);
xnor U2544 (N_2544,In_3271,N_1159);
nand U2545 (N_2545,In_1930,In_2887);
or U2546 (N_2546,N_2279,In_3842);
and U2547 (N_2547,In_612,N_2389);
nand U2548 (N_2548,N_978,In_4594);
or U2549 (N_2549,N_138,In_4045);
nor U2550 (N_2550,In_2290,N_1483);
xor U2551 (N_2551,N_2082,N_1638);
and U2552 (N_2552,N_2212,In_802);
nor U2553 (N_2553,N_2175,N_1439);
xnor U2554 (N_2554,N_464,N_1647);
nand U2555 (N_2555,N_1114,N_761);
and U2556 (N_2556,In_510,In_642);
nand U2557 (N_2557,N_2373,N_1757);
or U2558 (N_2558,In_1507,N_1736);
nor U2559 (N_2559,In_2258,N_1959);
nor U2560 (N_2560,In_4474,In_2041);
and U2561 (N_2561,In_2415,N_1809);
nand U2562 (N_2562,N_1677,In_3296);
nor U2563 (N_2563,N_2199,In_4997);
nand U2564 (N_2564,N_1911,N_1555);
and U2565 (N_2565,In_3017,In_4116);
xor U2566 (N_2566,In_1127,N_2020);
or U2567 (N_2567,N_1325,In_3901);
or U2568 (N_2568,N_2469,N_1210);
nor U2569 (N_2569,In_1398,N_1994);
nand U2570 (N_2570,N_1526,In_3246);
and U2571 (N_2571,N_2305,In_1359);
nor U2572 (N_2572,N_2297,In_3836);
and U2573 (N_2573,In_1026,N_2400);
and U2574 (N_2574,In_3502,In_2140);
and U2575 (N_2575,In_3367,N_1345);
nand U2576 (N_2576,In_172,N_2359);
nor U2577 (N_2577,In_3667,In_3825);
or U2578 (N_2578,In_3442,In_3023);
nand U2579 (N_2579,N_2460,N_95);
xnor U2580 (N_2580,In_4836,N_1046);
nand U2581 (N_2581,N_1728,In_87);
and U2582 (N_2582,N_2069,In_3552);
xnor U2583 (N_2583,N_2244,In_1794);
xnor U2584 (N_2584,In_3134,N_1552);
and U2585 (N_2585,In_2622,N_2292);
or U2586 (N_2586,N_2390,N_862);
and U2587 (N_2587,N_2075,N_1892);
or U2588 (N_2588,In_4239,N_1930);
xor U2589 (N_2589,N_1860,In_2992);
nor U2590 (N_2590,In_3204,N_892);
or U2591 (N_2591,N_1071,N_1804);
and U2592 (N_2592,N_1496,N_799);
and U2593 (N_2593,In_4243,N_2482);
xnor U2594 (N_2594,N_1686,N_1169);
nand U2595 (N_2595,In_813,In_1162);
nand U2596 (N_2596,N_1235,In_1848);
xnor U2597 (N_2597,N_686,N_2287);
or U2598 (N_2598,In_516,In_1365);
nand U2599 (N_2599,N_1291,N_2019);
and U2600 (N_2600,N_2342,In_3746);
or U2601 (N_2601,In_3545,In_622);
and U2602 (N_2602,N_2266,N_2007);
xnor U2603 (N_2603,N_2031,In_3461);
nand U2604 (N_2604,N_1848,N_302);
or U2605 (N_2605,N_374,N_2058);
and U2606 (N_2606,In_4333,N_1786);
and U2607 (N_2607,N_788,In_4121);
and U2608 (N_2608,N_2130,In_1571);
nor U2609 (N_2609,In_2635,N_1890);
and U2610 (N_2610,In_1630,N_1627);
nor U2611 (N_2611,N_16,N_2430);
nor U2612 (N_2612,In_2952,In_1369);
and U2613 (N_2613,N_106,N_1622);
nand U2614 (N_2614,N_2299,In_2771);
nand U2615 (N_2615,In_3087,In_3979);
or U2616 (N_2616,N_1819,N_2028);
xor U2617 (N_2617,N_1566,In_1559);
xor U2618 (N_2618,In_1867,In_1284);
and U2619 (N_2619,N_1187,In_2602);
nand U2620 (N_2620,N_459,In_3431);
nor U2621 (N_2621,N_80,N_2034);
nand U2622 (N_2622,N_1286,N_2300);
and U2623 (N_2623,In_1252,In_140);
or U2624 (N_2624,N_2027,N_1383);
and U2625 (N_2625,In_1362,In_2309);
nor U2626 (N_2626,N_646,N_2003);
nand U2627 (N_2627,N_2246,In_3166);
nor U2628 (N_2628,In_665,N_1843);
xor U2629 (N_2629,N_1945,N_1370);
and U2630 (N_2630,N_2491,N_635);
or U2631 (N_2631,In_2350,N_2218);
or U2632 (N_2632,In_916,N_304);
and U2633 (N_2633,In_327,In_3774);
and U2634 (N_2634,N_615,In_4353);
nand U2635 (N_2635,N_1774,N_2466);
and U2636 (N_2636,In_349,In_1569);
nor U2637 (N_2637,In_1475,In_1781);
and U2638 (N_2638,In_3969,N_1158);
nor U2639 (N_2639,N_2072,In_619);
xor U2640 (N_2640,N_2458,In_3495);
and U2641 (N_2641,In_4457,In_4156);
nand U2642 (N_2642,In_1958,N_861);
xnor U2643 (N_2643,In_4861,In_2024);
nand U2644 (N_2644,N_1298,In_2721);
or U2645 (N_2645,N_2254,N_479);
or U2646 (N_2646,N_2423,N_1254);
xnor U2647 (N_2647,In_3114,N_760);
or U2648 (N_2648,N_2207,In_218);
and U2649 (N_2649,N_2039,In_2981);
and U2650 (N_2650,N_2298,In_4084);
or U2651 (N_2651,In_3401,N_2411);
or U2652 (N_2652,In_2113,In_551);
nand U2653 (N_2653,In_1366,N_1400);
nand U2654 (N_2654,N_1490,N_1054);
xor U2655 (N_2655,In_1182,N_1651);
nand U2656 (N_2656,N_1741,In_3348);
xor U2657 (N_2657,In_937,N_1606);
nand U2658 (N_2658,N_1006,N_1940);
nand U2659 (N_2659,N_2059,N_177);
or U2660 (N_2660,In_4804,In_4719);
or U2661 (N_2661,N_1430,In_3499);
nor U2662 (N_2662,In_509,N_1281);
nor U2663 (N_2663,In_3195,In_127);
and U2664 (N_2664,N_771,N_2280);
nor U2665 (N_2665,In_3857,N_1865);
xnor U2666 (N_2666,N_1067,N_2221);
nor U2667 (N_2667,N_2169,In_2684);
or U2668 (N_2668,N_1694,N_1438);
nand U2669 (N_2669,In_1520,In_1924);
and U2670 (N_2670,N_1253,N_836);
xor U2671 (N_2671,In_3936,N_1825);
xnor U2672 (N_2672,In_1075,N_1750);
or U2673 (N_2673,N_1859,N_1751);
xnor U2674 (N_2674,N_1681,N_1095);
nor U2675 (N_2675,In_3730,N_1043);
nor U2676 (N_2676,In_3567,In_501);
and U2677 (N_2677,N_1896,N_1306);
xor U2678 (N_2678,N_2481,In_13);
nor U2679 (N_2679,In_3942,N_1128);
nor U2680 (N_2680,N_1632,N_2356);
nor U2681 (N_2681,N_2223,In_597);
nor U2682 (N_2682,N_1772,In_2679);
xor U2683 (N_2683,In_993,In_1441);
and U2684 (N_2684,N_2321,In_2744);
xnor U2685 (N_2685,N_2099,N_1539);
and U2686 (N_2686,In_3363,In_837);
nor U2687 (N_2687,In_1344,In_512);
xor U2688 (N_2688,In_2458,In_733);
xor U2689 (N_2689,In_1261,N_2457);
nor U2690 (N_2690,N_2377,N_768);
nand U2691 (N_2691,N_1924,N_2407);
and U2692 (N_2692,N_536,N_2319);
nand U2693 (N_2693,In_2780,In_376);
or U2694 (N_2694,N_848,In_2021);
and U2695 (N_2695,In_2374,In_1749);
nand U2696 (N_2696,In_3026,N_1831);
and U2697 (N_2697,In_364,N_1211);
nand U2698 (N_2698,N_2413,In_487);
nand U2699 (N_2699,In_2913,N_1748);
nor U2700 (N_2700,N_1222,N_1031);
xnor U2701 (N_2701,In_4411,N_1785);
nand U2702 (N_2702,N_2410,N_1996);
nand U2703 (N_2703,In_3439,N_1657);
or U2704 (N_2704,In_4016,N_2374);
and U2705 (N_2705,N_2348,In_4074);
nand U2706 (N_2706,N_1954,N_1758);
nand U2707 (N_2707,N_884,N_1993);
nand U2708 (N_2708,In_2471,N_242);
nor U2709 (N_2709,In_882,In_3770);
nand U2710 (N_2710,N_2239,N_1151);
nand U2711 (N_2711,N_2439,N_1045);
or U2712 (N_2712,In_2499,N_1475);
nand U2713 (N_2713,N_2056,N_1695);
and U2714 (N_2714,In_4124,In_4232);
nor U2715 (N_2715,N_2490,In_2314);
xnor U2716 (N_2716,N_786,N_1494);
and U2717 (N_2717,In_4611,N_1957);
nor U2718 (N_2718,In_4782,N_1767);
xnor U2719 (N_2719,In_2818,N_2353);
xnor U2720 (N_2720,In_2781,N_537);
nand U2721 (N_2721,N_1394,In_393);
nor U2722 (N_2722,N_199,In_786);
nor U2723 (N_2723,N_2419,N_119);
or U2724 (N_2724,In_953,In_1623);
nor U2725 (N_2725,N_2000,N_1987);
nor U2726 (N_2726,N_2235,In_2363);
nor U2727 (N_2727,In_108,In_3519);
or U2728 (N_2728,In_3764,N_1703);
or U2729 (N_2729,N_1469,N_1375);
or U2730 (N_2730,N_1560,In_121);
nand U2731 (N_2731,In_1353,N_2303);
and U2732 (N_2732,In_3170,N_2424);
nor U2733 (N_2733,In_1203,In_392);
or U2734 (N_2734,In_2852,In_3593);
nor U2735 (N_2735,N_2205,In_1814);
nor U2736 (N_2736,In_1435,In_1164);
xnor U2737 (N_2737,N_1971,N_1601);
and U2738 (N_2738,N_1898,In_3945);
or U2739 (N_2739,N_2450,N_2333);
nor U2740 (N_2740,In_2279,In_1716);
nor U2741 (N_2741,In_2815,N_860);
nor U2742 (N_2742,In_2323,N_124);
nor U2743 (N_2743,In_2485,N_2037);
nand U2744 (N_2744,N_2210,In_50);
nand U2745 (N_2745,In_1590,N_2098);
nor U2746 (N_2746,N_1943,N_2161);
xor U2747 (N_2747,N_307,N_2492);
nand U2748 (N_2748,In_35,In_594);
or U2749 (N_2749,In_4915,N_2290);
nor U2750 (N_2750,In_1012,N_2516);
nand U2751 (N_2751,In_4356,N_2142);
and U2752 (N_2752,N_2393,N_2535);
and U2753 (N_2753,N_1832,N_1300);
nand U2754 (N_2754,In_4438,N_6);
nand U2755 (N_2755,N_2045,N_1508);
nand U2756 (N_2756,In_3386,In_528);
or U2757 (N_2757,In_1421,In_4467);
xor U2758 (N_2758,N_2461,N_2071);
or U2759 (N_2759,N_2141,In_1908);
or U2760 (N_2760,N_2023,N_1899);
nand U2761 (N_2761,In_2928,N_2160);
nand U2762 (N_2762,N_1913,In_4146);
or U2763 (N_2763,N_763,N_2436);
and U2764 (N_2764,In_2846,In_995);
nor U2765 (N_2765,N_2642,In_3142);
xor U2766 (N_2766,N_1597,In_3943);
nor U2767 (N_2767,In_4148,N_2570);
nor U2768 (N_2768,N_577,In_2895);
and U2769 (N_2769,N_2268,In_1358);
nand U2770 (N_2770,N_932,In_471);
nor U2771 (N_2771,In_2789,N_2204);
nor U2772 (N_2772,N_1255,N_1520);
and U2773 (N_2773,N_2543,In_4773);
nor U2774 (N_2774,N_1492,N_751);
nand U2775 (N_2775,N_2513,N_1357);
and U2776 (N_2776,In_302,In_3052);
xor U2777 (N_2777,N_1777,In_1350);
xor U2778 (N_2778,In_4494,N_1360);
and U2779 (N_2779,N_2567,N_1855);
xor U2780 (N_2780,In_1615,N_1319);
xnor U2781 (N_2781,In_56,In_853);
or U2782 (N_2782,N_313,In_1745);
and U2783 (N_2783,In_4221,In_1307);
nand U2784 (N_2784,N_2245,In_4568);
nor U2785 (N_2785,In_1664,N_1722);
nor U2786 (N_2786,N_2267,N_2600);
nand U2787 (N_2787,N_1521,N_1198);
and U2788 (N_2788,In_2591,N_2402);
or U2789 (N_2789,N_1214,N_2181);
or U2790 (N_2790,N_407,N_1389);
xnor U2791 (N_2791,N_1977,N_1938);
nand U2792 (N_2792,In_460,In_3902);
and U2793 (N_2793,N_2166,In_2941);
nand U2794 (N_2794,In_4737,N_1460);
and U2795 (N_2795,In_1406,N_2046);
xnor U2796 (N_2796,In_2756,In_1933);
nand U2797 (N_2797,N_2534,In_2225);
xnor U2798 (N_2798,N_535,In_1146);
and U2799 (N_2799,N_637,In_1324);
or U2800 (N_2800,In_3376,N_2051);
nand U2801 (N_2801,N_2694,N_2262);
and U2802 (N_2802,N_2346,N_2736);
nor U2803 (N_2803,In_379,In_3398);
xnor U2804 (N_2804,N_2506,N_2663);
nor U2805 (N_2805,In_2923,N_2676);
xor U2806 (N_2806,In_3660,In_2226);
or U2807 (N_2807,In_1086,N_2231);
or U2808 (N_2808,In_2118,In_1357);
and U2809 (N_2809,In_2854,N_827);
nand U2810 (N_2810,N_2434,N_2240);
nand U2811 (N_2811,In_3748,In_3622);
nor U2812 (N_2812,N_1590,N_51);
or U2813 (N_2813,In_803,N_1968);
and U2814 (N_2814,N_2073,N_2733);
or U2815 (N_2815,N_2208,In_2742);
or U2816 (N_2816,In_2092,In_3077);
or U2817 (N_2817,In_4047,In_4533);
and U2818 (N_2818,N_2257,In_2278);
nand U2819 (N_2819,N_665,In_2955);
and U2820 (N_2820,In_1626,In_3267);
nor U2821 (N_2821,In_4635,N_2504);
nor U2822 (N_2822,N_529,In_1540);
xor U2823 (N_2823,N_2697,N_2323);
and U2824 (N_2824,In_4346,N_2277);
or U2825 (N_2825,N_1885,In_2552);
nand U2826 (N_2826,N_2584,N_1683);
xor U2827 (N_2827,In_1179,In_246);
nand U2828 (N_2828,In_1133,In_4526);
nor U2829 (N_2829,N_955,N_954);
or U2830 (N_2830,N_994,N_2718);
and U2831 (N_2831,In_2376,In_4822);
and U2832 (N_2832,N_1461,N_287);
nand U2833 (N_2833,In_4028,N_499);
and U2834 (N_2834,In_2402,In_1055);
and U2835 (N_2835,N_1955,In_3852);
nand U2836 (N_2836,N_545,N_752);
nand U2837 (N_2837,In_331,N_2585);
nor U2838 (N_2838,N_1505,N_671);
or U2839 (N_2839,In_967,In_1183);
xor U2840 (N_2840,In_1103,N_2387);
and U2841 (N_2841,N_1662,In_98);
and U2842 (N_2842,In_1184,N_2728);
and U2843 (N_2843,In_4616,N_820);
nor U2844 (N_2844,N_2217,In_3712);
nor U2845 (N_2845,In_3934,N_1148);
or U2846 (N_2846,In_3254,N_2451);
nor U2847 (N_2847,In_4168,In_294);
or U2848 (N_2848,In_4329,In_1863);
nand U2849 (N_2849,N_2128,In_3638);
and U2850 (N_2850,In_3464,N_96);
or U2851 (N_2851,N_210,N_2309);
nor U2852 (N_2852,In_360,In_1392);
nand U2853 (N_2853,In_591,N_2550);
and U2854 (N_2854,In_462,In_939);
nand U2855 (N_2855,N_1354,In_2070);
or U2856 (N_2856,In_4064,N_1450);
nor U2857 (N_2857,N_1808,N_2514);
xor U2858 (N_2858,N_1829,N_618);
or U2859 (N_2859,In_1154,N_1812);
nor U2860 (N_2860,N_2155,In_109);
nand U2861 (N_2861,In_2765,In_4250);
nand U2862 (N_2862,In_608,In_1304);
or U2863 (N_2863,N_2639,N_1471);
nand U2864 (N_2864,N_311,N_2260);
or U2865 (N_2865,N_796,N_1756);
nand U2866 (N_2866,In_1438,N_2644);
and U2867 (N_2867,In_558,In_3723);
nand U2868 (N_2868,N_2592,In_1766);
xnor U2869 (N_2869,N_263,In_3985);
and U2870 (N_2870,N_2569,In_3210);
or U2871 (N_2871,In_2253,N_1420);
nor U2872 (N_2872,N_2555,N_2532);
nor U2873 (N_2873,N_2672,In_370);
nand U2874 (N_2874,N_2395,In_1676);
xor U2875 (N_2875,N_2165,In_1556);
nand U2876 (N_2876,N_2727,In_1801);
and U2877 (N_2877,In_4657,N_1944);
nand U2878 (N_2878,N_910,In_4222);
and U2879 (N_2879,N_1209,N_2713);
nand U2880 (N_2880,In_550,N_1304);
or U2881 (N_2881,In_1072,In_1938);
and U2882 (N_2882,In_4349,N_968);
or U2883 (N_2883,N_1925,N_324);
and U2884 (N_2884,N_1684,In_441);
or U2885 (N_2885,In_4512,N_2633);
nor U2886 (N_2886,In_1901,N_2183);
xor U2887 (N_2887,N_2151,In_4590);
nor U2888 (N_2888,N_530,N_1969);
or U2889 (N_2889,N_2327,In_3069);
nand U2890 (N_2890,N_473,In_1611);
and U2891 (N_2891,In_4962,N_2660);
or U2892 (N_2892,In_4630,N_972);
or U2893 (N_2893,In_2541,In_4340);
or U2894 (N_2894,N_2606,In_4170);
nor U2895 (N_2895,In_2160,N_1248);
nor U2896 (N_2896,N_2304,In_1999);
or U2897 (N_2897,N_2507,N_2746);
nor U2898 (N_2898,In_3804,In_8);
nor U2899 (N_2899,N_1723,N_1241);
or U2900 (N_2900,N_1032,In_4551);
xnor U2901 (N_2901,In_1195,N_2502);
or U2902 (N_2902,In_85,N_2433);
or U2903 (N_2903,N_2398,N_2706);
nand U2904 (N_2904,In_3888,In_2647);
and U2905 (N_2905,N_652,N_2399);
nor U2906 (N_2906,N_2626,N_1836);
or U2907 (N_2907,N_1866,N_1398);
nor U2908 (N_2908,In_3711,N_1636);
and U2909 (N_2909,N_2632,N_1487);
or U2910 (N_2910,N_2101,In_2310);
nand U2911 (N_2911,In_3749,N_2089);
or U2912 (N_2912,In_3070,N_913);
nor U2913 (N_2913,In_2951,In_2221);
nor U2914 (N_2914,In_4641,In_2289);
xnor U2915 (N_2915,N_653,In_2015);
nand U2916 (N_2916,In_2719,In_3778);
or U2917 (N_2917,N_2687,N_2392);
xnor U2918 (N_2918,N_2521,N_1136);
nand U2919 (N_2919,N_853,In_1291);
nand U2920 (N_2920,In_2051,In_3612);
or U2921 (N_2921,In_2547,N_863);
and U2922 (N_2922,N_2337,N_794);
nand U2923 (N_2923,In_477,N_165);
or U2924 (N_2924,In_2621,N_1658);
nor U2925 (N_2925,In_4292,N_2224);
nand U2926 (N_2926,In_4316,In_2942);
nand U2927 (N_2927,In_2497,N_2558);
and U2928 (N_2928,N_2629,In_1715);
xor U2929 (N_2929,N_2196,N_1581);
nand U2930 (N_2930,In_1090,N_2310);
nand U2931 (N_2931,In_119,In_1318);
or U2932 (N_2932,In_4653,N_931);
or U2933 (N_2933,In_3987,N_2612);
or U2934 (N_2934,N_681,N_1070);
or U2935 (N_2935,N_1714,N_2462);
and U2936 (N_2936,N_2361,N_2261);
nand U2937 (N_2937,In_312,In_3284);
and U2938 (N_2938,In_2834,In_1464);
nor U2939 (N_2939,N_1115,N_524);
or U2940 (N_2940,N_1939,N_1879);
xnor U2941 (N_2941,N_2705,N_2623);
or U2942 (N_2942,In_2746,In_507);
nor U2943 (N_2943,N_624,N_1036);
or U2944 (N_2944,N_2508,N_1729);
or U2945 (N_2945,N_667,N_1186);
or U2946 (N_2946,N_2501,N_2247);
or U2947 (N_2947,N_1842,N_2313);
nand U2948 (N_2948,N_2150,N_491);
nor U2949 (N_2949,N_1156,In_4906);
and U2950 (N_2950,N_1315,N_1749);
nand U2951 (N_2951,In_3304,In_2430);
nor U2952 (N_2952,In_3050,In_2109);
xnor U2953 (N_2953,In_2112,N_1696);
or U2954 (N_2954,In_3018,N_2673);
or U2955 (N_2955,N_1818,N_2132);
nand U2956 (N_2956,N_1249,N_1839);
and U2957 (N_2957,N_2695,In_3809);
nand U2958 (N_2958,In_480,N_2522);
or U2959 (N_2959,N_2255,N_2489);
or U2960 (N_2960,In_692,N_2599);
nor U2961 (N_2961,N_1448,In_3206);
xor U2962 (N_2962,In_1777,In_854);
or U2963 (N_2963,N_909,In_2745);
nand U2964 (N_2964,N_125,N_1549);
nand U2965 (N_2965,N_694,N_1907);
nor U2966 (N_2966,N_1827,In_1347);
xnor U2967 (N_2967,N_2397,N_2408);
or U2968 (N_2968,In_620,N_1737);
and U2969 (N_2969,In_45,N_1519);
or U2970 (N_2970,N_2573,N_1386);
or U2971 (N_2971,N_2422,N_448);
nor U2972 (N_2972,N_1589,N_2325);
or U2973 (N_2973,N_2580,N_2162);
nor U2974 (N_2974,N_2478,In_3470);
nand U2975 (N_2975,N_1755,N_2100);
nor U2976 (N_2976,N_2372,N_1926);
nand U2977 (N_2977,N_1915,N_2167);
or U2978 (N_2978,In_3941,N_2264);
xor U2979 (N_2979,N_622,N_1887);
nand U2980 (N_2980,N_2732,In_599);
and U2981 (N_2981,N_2636,In_566);
xnor U2982 (N_2982,N_1814,In_4463);
or U2983 (N_2983,In_954,N_2724);
nand U2984 (N_2984,In_2438,N_1625);
nor U2985 (N_2985,N_1348,N_1650);
and U2986 (N_2986,N_2029,N_891);
nand U2987 (N_2987,N_2517,N_2611);
and U2988 (N_2988,In_260,N_2509);
or U2989 (N_2989,In_2973,N_2646);
xnor U2990 (N_2990,N_2485,N_298);
xor U2991 (N_2991,N_1614,In_2752);
nand U2992 (N_2992,N_2381,N_1962);
or U2993 (N_2993,N_2140,N_2678);
xnor U2994 (N_2994,In_1764,N_2539);
xor U2995 (N_2995,In_2231,N_1856);
nor U2996 (N_2996,N_526,N_2735);
nand U2997 (N_2997,In_1138,N_1844);
nand U2998 (N_2998,N_673,N_2044);
and U2999 (N_2999,In_1638,N_1952);
xnor U3000 (N_3000,N_1048,N_769);
nand U3001 (N_3001,N_2013,In_588);
and U3002 (N_3002,N_610,N_2093);
xnor U3003 (N_3003,N_2936,N_1362);
xnor U3004 (N_3004,N_2384,In_3988);
xnor U3005 (N_3005,N_1615,N_2869);
or U3006 (N_3006,N_951,N_486);
nand U3007 (N_3007,In_796,N_2725);
or U3008 (N_3008,In_4464,N_2933);
and U3009 (N_3009,In_1986,In_1812);
nand U3010 (N_3010,N_75,N_2669);
nor U3011 (N_3011,N_1992,N_1810);
or U3012 (N_3012,In_3024,N_1800);
nand U3013 (N_3013,N_2409,N_2800);
nor U3014 (N_3014,N_2537,N_1269);
or U3015 (N_3015,N_2016,N_2388);
or U3016 (N_3016,In_1998,In_2381);
and U3017 (N_3017,N_2793,In_4372);
or U3018 (N_3018,N_2030,N_1347);
nor U3019 (N_3019,In_2040,N_2357);
xor U3020 (N_3020,In_498,In_219);
or U3021 (N_3021,In_4898,N_2014);
or U3022 (N_3022,N_335,N_1608);
nand U3023 (N_3023,N_1038,N_1591);
nand U3024 (N_3024,N_2703,N_823);
nand U3025 (N_3025,In_1979,In_2785);
xnor U3026 (N_3026,N_2180,N_2553);
nor U3027 (N_3027,N_2919,In_2212);
nand U3028 (N_3028,In_3636,N_1507);
or U3029 (N_3029,In_4925,N_2288);
nand U3030 (N_3030,In_4326,N_1671);
or U3031 (N_3031,N_944,N_470);
xor U3032 (N_3032,N_474,In_2934);
xnor U3033 (N_3033,N_2542,N_2743);
or U3034 (N_3034,N_2892,In_1708);
xnor U3035 (N_3035,N_2830,N_870);
nand U3036 (N_3036,In_2772,N_658);
and U3037 (N_3037,N_1301,N_2658);
nand U3038 (N_3038,In_3403,In_636);
nand U3039 (N_3039,N_2683,N_2899);
or U3040 (N_3040,In_212,N_1693);
nand U3041 (N_3041,N_2428,In_2529);
xor U3042 (N_3042,In_2327,N_1243);
nand U3043 (N_3043,N_1342,N_2740);
nand U3044 (N_3044,N_919,N_291);
or U3045 (N_3045,N_2117,In_4262);
and U3046 (N_3046,In_4553,N_2749);
or U3047 (N_3047,In_10,In_4684);
nor U3048 (N_3048,N_977,N_1639);
nor U3049 (N_3049,N_1561,N_2315);
nand U3050 (N_3050,In_3124,N_1310);
nand U3051 (N_3051,N_2613,N_340);
and U3052 (N_3052,N_2769,In_1111);
xor U3053 (N_3053,N_1630,In_1388);
nor U3054 (N_3054,N_2867,N_379);
xnor U3055 (N_3055,N_2854,N_36);
nand U3056 (N_3056,N_2614,In_2656);
and U3057 (N_3057,N_2417,N_2991);
nand U3058 (N_3058,N_1260,N_2744);
nor U3059 (N_3059,N_1931,In_3704);
nor U3060 (N_3060,In_603,N_2194);
and U3061 (N_3061,N_2976,In_2206);
nor U3062 (N_3062,N_2576,N_172);
and U3063 (N_3063,In_554,In_4860);
and U3064 (N_3064,In_473,In_1918);
xor U3065 (N_3065,In_1903,N_2649);
and U3066 (N_3066,N_2242,In_2784);
xor U3067 (N_3067,In_2213,In_3782);
nand U3068 (N_3068,In_2617,N_2035);
nand U3069 (N_3069,In_1269,N_2847);
xnor U3070 (N_3070,In_2733,N_1381);
or U3071 (N_3071,N_2775,In_1703);
nand U3072 (N_3072,In_3108,In_4198);
xor U3073 (N_3073,In_3467,N_797);
nand U3074 (N_3074,In_1984,N_2365);
xor U3075 (N_3075,N_2563,In_2930);
nor U3076 (N_3076,N_1124,In_3798);
nor U3077 (N_3077,N_261,N_2812);
and U3078 (N_3078,In_4880,N_2383);
xor U3079 (N_3079,In_2637,N_2909);
and U3080 (N_3080,N_881,N_2843);
or U3081 (N_3081,N_2418,In_4069);
nor U3082 (N_3082,N_2961,In_2325);
xnor U3083 (N_3083,In_1028,In_96);
nor U3084 (N_3084,N_2281,N_1129);
and U3085 (N_3085,N_47,N_2017);
nand U3086 (N_3086,N_1172,In_4473);
nand U3087 (N_3087,In_3765,In_982);
or U3088 (N_3088,N_2883,In_184);
nor U3089 (N_3089,N_2688,N_1858);
nor U3090 (N_3090,N_433,N_1244);
nand U3091 (N_3091,In_3731,N_690);
nand U3092 (N_3092,N_2662,N_2983);
or U3093 (N_3093,In_3591,N_2741);
or U3094 (N_3094,N_2578,N_1307);
or U3095 (N_3095,In_4355,In_2354);
nor U3096 (N_3096,In_2052,N_2096);
and U3097 (N_3097,In_4959,N_1801);
nor U3098 (N_3098,In_655,N_1903);
or U3099 (N_3099,In_2796,N_2330);
or U3100 (N_3100,N_2868,N_953);
or U3101 (N_3101,N_2890,N_2872);
nand U3102 (N_3102,In_2254,N_2090);
and U3103 (N_3103,N_2404,N_468);
or U3104 (N_3104,In_120,N_1116);
or U3105 (N_3105,In_571,In_2111);
and U3106 (N_3106,N_2159,N_2602);
or U3107 (N_3107,N_1965,N_701);
or U3108 (N_3108,N_2370,N_1826);
nor U3109 (N_3109,N_2875,N_240);
and U3110 (N_3110,N_2693,N_221);
or U3111 (N_3111,N_2973,In_1328);
nand U3112 (N_3112,N_1283,N_58);
or U3113 (N_3113,N_2900,N_2541);
nor U3114 (N_3114,N_2463,N_2604);
nand U3115 (N_3115,N_2982,In_2192);
or U3116 (N_3116,N_2289,In_3937);
or U3117 (N_3117,In_2400,In_2148);
and U3118 (N_3118,In_3315,In_3891);
nor U3119 (N_3119,In_4102,In_1311);
or U3120 (N_3120,In_4252,In_3151);
and U3121 (N_3121,In_3196,In_225);
xor U3122 (N_3122,N_2076,In_3627);
xnor U3123 (N_3123,N_2734,N_2894);
nand U3124 (N_3124,N_2929,N_1999);
and U3125 (N_3125,N_2827,N_1405);
nor U3126 (N_3126,N_2911,N_2078);
and U3127 (N_3127,N_1251,N_1927);
nand U3128 (N_3128,In_1629,N_2596);
and U3129 (N_3129,N_2974,In_329);
and U3130 (N_3130,N_2057,N_1557);
and U3131 (N_3131,N_465,N_2956);
xor U3132 (N_3132,N_1366,In_2305);
or U3133 (N_3133,N_2286,N_2498);
or U3134 (N_3134,N_980,N_2109);
nand U3135 (N_3135,N_1929,In_2005);
nor U3136 (N_3136,In_1789,N_2671);
and U3137 (N_3137,In_2132,N_2849);
and U3138 (N_3138,N_2448,N_809);
nand U3139 (N_3139,N_57,In_3057);
xnor U3140 (N_3140,In_4936,N_276);
or U3141 (N_3141,N_2568,N_2730);
xnor U3142 (N_3142,In_4144,N_2942);
nand U3143 (N_3143,In_3655,N_719);
and U3144 (N_3144,In_1391,N_1003);
xnor U3145 (N_3145,N_1238,In_2422);
or U3146 (N_3146,N_2213,N_1868);
and U3147 (N_3147,N_2429,N_2085);
nand U3148 (N_3148,In_1157,N_2475);
and U3149 (N_3149,In_4008,N_2102);
nor U3150 (N_3150,N_1246,N_1982);
xor U3151 (N_3151,N_2928,In_758);
or U3152 (N_3152,N_2786,N_2700);
and U3153 (N_3153,N_2302,In_2700);
and U3154 (N_3154,In_4171,In_78);
or U3155 (N_3155,N_1449,N_2086);
xor U3156 (N_3156,In_1941,In_1334);
and U3157 (N_3157,N_1760,In_1187);
nand U3158 (N_3158,N_2593,N_1669);
nand U3159 (N_3159,N_2104,N_2012);
xnor U3160 (N_3160,N_2339,In_1797);
nand U3161 (N_3161,In_868,N_2193);
xor U3162 (N_3162,N_2598,N_2396);
and U3163 (N_3163,In_4858,N_1289);
or U3164 (N_3164,In_3896,N_1062);
nor U3165 (N_3165,N_2062,N_2064);
nand U3166 (N_3166,N_2296,N_1161);
nand U3167 (N_3167,In_2567,In_2378);
nor U3168 (N_3168,N_350,In_1697);
or U3169 (N_3169,N_2220,In_2018);
nor U3170 (N_3170,N_2420,N_2380);
xor U3171 (N_3171,In_4034,N_1894);
nand U3172 (N_3172,N_2684,In_657);
nor U3173 (N_3173,N_742,In_2663);
nand U3174 (N_3174,In_2025,In_2304);
and U3175 (N_3175,In_4161,N_989);
or U3176 (N_3176,In_2639,In_2406);
xor U3177 (N_3177,In_4698,N_1163);
nand U3178 (N_3178,N_2722,N_369);
nand U3179 (N_3179,In_2375,N_318);
and U3180 (N_3180,In_1588,N_1821);
nor U3181 (N_3181,In_2592,In_1425);
and U3182 (N_3182,In_4487,N_2001);
nand U3183 (N_3183,In_301,N_2316);
or U3184 (N_3184,N_500,N_1793);
nand U3185 (N_3185,N_1633,N_1739);
nor U3186 (N_3186,In_2848,N_575);
and U3187 (N_3187,N_2903,N_2647);
xnor U3188 (N_3188,N_1188,N_2908);
xnor U3189 (N_3189,In_2890,In_2370);
or U3190 (N_3190,In_3686,N_2355);
xor U3191 (N_3191,N_1012,N_1327);
and U3192 (N_3192,In_3919,In_4485);
nand U3193 (N_3193,N_2344,N_506);
xnor U3194 (N_3194,N_2552,In_3098);
nor U3195 (N_3195,In_1470,In_4036);
xnor U3196 (N_3196,In_2935,N_1226);
or U3197 (N_3197,N_2813,In_2408);
or U3198 (N_3198,N_2345,N_2520);
xnor U3199 (N_3199,N_216,N_86);
xor U3200 (N_3200,N_151,In_515);
nand U3201 (N_3201,N_2681,N_2318);
and U3202 (N_3202,In_4304,In_125);
xor U3203 (N_3203,N_1359,In_4777);
and U3204 (N_3204,N_1509,N_2762);
or U3205 (N_3205,N_2627,N_2906);
or U3206 (N_3206,In_2038,In_3560);
nand U3207 (N_3207,N_2937,In_4307);
and U3208 (N_3208,N_2625,N_2369);
or U3209 (N_3209,N_2797,In_4644);
or U3210 (N_3210,In_3992,N_1435);
or U3211 (N_3211,N_2452,N_1648);
and U3212 (N_3212,In_702,In_1600);
nor U3213 (N_3213,N_2617,In_3983);
xnor U3214 (N_3214,In_3038,N_2360);
nor U3215 (N_3215,In_934,N_2792);
nand U3216 (N_3216,In_4508,In_2299);
and U3217 (N_3217,N_2807,N_1646);
and U3218 (N_3218,In_3063,N_2285);
nor U3219 (N_3219,N_2895,In_0);
xor U3220 (N_3220,N_1717,In_44);
nor U3221 (N_3221,N_444,In_4427);
and U3222 (N_3222,In_71,N_1986);
nand U3223 (N_3223,N_2441,In_544);
or U3224 (N_3224,N_1312,N_777);
nor U3225 (N_3225,N_2006,In_1560);
or U3226 (N_3226,In_1511,N_2574);
nand U3227 (N_3227,N_1145,In_3247);
xnor U3228 (N_3228,N_1634,In_3086);
or U3229 (N_3229,In_3239,N_2914);
and U3230 (N_3230,N_2464,N_2594);
nand U3231 (N_3231,N_2331,In_165);
nand U3232 (N_3232,In_1479,In_1920);
and U3233 (N_3233,N_204,In_1314);
and U3234 (N_3234,N_2845,N_168);
or U3235 (N_3235,N_300,N_1934);
nor U3236 (N_3236,N_1513,N_1680);
nor U3237 (N_3237,N_1486,In_2943);
nor U3238 (N_3238,N_1577,N_620);
nand U3239 (N_3239,In_2590,In_3625);
or U3240 (N_3240,In_1094,N_1058);
or U3241 (N_3241,In_4535,In_21);
xor U3242 (N_3242,In_1180,N_2670);
nand U3243 (N_3243,In_1001,N_2079);
nand U3244 (N_3244,N_1933,In_1554);
xor U3245 (N_3245,In_888,N_364);
nand U3246 (N_3246,N_2338,N_2178);
nor U3247 (N_3247,In_2977,N_2549);
nor U3248 (N_3248,In_2487,N_2144);
nand U3249 (N_3249,N_2871,In_2328);
xnor U3250 (N_3250,N_2546,N_2293);
nand U3251 (N_3251,N_2497,In_4951);
and U3252 (N_3252,N_2852,N_1495);
nand U3253 (N_3253,N_2857,N_292);
nor U3254 (N_3254,N_3024,N_3091);
nand U3255 (N_3255,N_2702,N_2877);
xor U3256 (N_3256,N_3115,In_1367);
or U3257 (N_3257,N_3215,In_1100);
or U3258 (N_3258,N_2790,N_2562);
and U3259 (N_3259,N_2715,In_1403);
xor U3260 (N_3260,In_2372,In_428);
and U3261 (N_3261,N_2616,N_2547);
nand U3262 (N_3262,In_3433,In_3078);
or U3263 (N_3263,N_2105,N_1288);
and U3264 (N_3264,N_1497,N_2737);
or U3265 (N_3265,N_3200,N_2955);
nand U3266 (N_3266,In_414,In_1310);
nand U3267 (N_3267,N_3058,In_3910);
xnor U3268 (N_3268,N_2620,N_2328);
and U3269 (N_3269,N_2503,In_4886);
or U3270 (N_3270,N_2468,In_563);
nor U3271 (N_3271,N_1790,N_2477);
or U3272 (N_3272,N_1678,N_3243);
or U3273 (N_3273,N_2886,N_2862);
nand U3274 (N_3274,N_3052,N_2002);
xnor U3275 (N_3275,In_850,In_3630);
and U3276 (N_3276,N_2912,N_2499);
or U3277 (N_3277,N_2941,N_1433);
nand U3278 (N_3278,N_2136,N_2696);
or U3279 (N_3279,N_2094,N_1279);
nand U3280 (N_3280,N_2851,N_2362);
or U3281 (N_3281,N_3009,N_518);
nand U3282 (N_3282,In_3518,N_1626);
nor U3283 (N_3283,N_2897,N_3189);
and U3284 (N_3284,In_1572,In_1408);
nor U3285 (N_3285,N_2653,N_2295);
nor U3286 (N_3286,N_2554,N_2779);
and U3287 (N_3287,N_2766,N_3241);
nand U3288 (N_3288,N_2445,In_3584);
xnor U3289 (N_3289,N_1550,N_2227);
and U3290 (N_3290,N_2804,N_386);
xor U3291 (N_3291,In_1799,N_1275);
nor U3292 (N_3292,N_800,N_3067);
or U3293 (N_3293,N_568,In_2134);
nor U3294 (N_3294,N_2747,In_2898);
and U3295 (N_3295,N_1385,N_1034);
and U3296 (N_3296,N_2719,N_2440);
and U3297 (N_3297,N_2065,N_2938);
or U3298 (N_3298,N_2918,N_2915);
nand U3299 (N_3299,N_492,N_418);
or U3300 (N_3300,N_1112,In_3352);
and U3301 (N_3301,N_1201,N_447);
nor U3302 (N_3302,In_4875,N_516);
xor U3303 (N_3303,In_2945,N_2421);
or U3304 (N_3304,N_2018,In_4412);
and U3305 (N_3305,In_1008,N_3222);
nand U3306 (N_3306,N_1239,In_757);
and U3307 (N_3307,In_1237,In_4234);
nor U3308 (N_3308,In_463,N_2921);
and U3309 (N_3309,N_3233,In_3811);
nor U3310 (N_3310,N_561,N_2828);
or U3311 (N_3311,N_3192,N_3087);
nor U3312 (N_3312,N_896,N_3013);
and U3313 (N_3313,N_3114,In_525);
nor U3314 (N_3314,N_2211,N_2880);
and U3315 (N_3315,N_3197,N_1909);
or U3316 (N_3316,N_1853,N_1203);
nor U3317 (N_3317,N_3127,In_3423);
nor U3318 (N_3318,N_3026,N_857);
nor U3319 (N_3319,N_1917,N_2953);
nor U3320 (N_3320,In_2502,N_3171);
nor U3321 (N_3321,N_2950,N_1976);
and U3322 (N_3322,N_3216,N_2655);
and U3323 (N_3323,N_2352,In_1048);
nor U3324 (N_3324,N_2126,In_4061);
nor U3325 (N_3325,N_3025,N_2538);
or U3326 (N_3326,N_1886,In_3354);
nand U3327 (N_3327,In_2675,In_328);
nor U3328 (N_3328,In_3526,N_2157);
and U3329 (N_3329,N_2838,In_4701);
nand U3330 (N_3330,In_1126,N_3193);
nand U3331 (N_3331,N_832,In_3128);
nand U3332 (N_3332,In_911,N_1292);
nor U3333 (N_3333,N_2969,In_1446);
and U3334 (N_3334,N_3146,In_3974);
and U3335 (N_3335,In_3493,In_1302);
and U3336 (N_3336,N_2848,In_4229);
or U3337 (N_3337,In_3056,N_1089);
xnor U3338 (N_3338,N_2720,N_3232);
nand U3339 (N_3339,N_1778,N_310);
nor U3340 (N_3340,N_2505,In_2802);
or U3341 (N_3341,N_2233,N_2835);
or U3342 (N_3342,N_3061,N_3226);
nand U3343 (N_3343,In_4688,In_3344);
or U3344 (N_3344,N_1904,In_4863);
nand U3345 (N_3345,N_2726,N_91);
xnor U3346 (N_3346,N_1050,N_3248);
xor U3347 (N_3347,N_1864,In_3245);
xor U3348 (N_3348,In_1612,N_2885);
or U3349 (N_3349,N_945,N_592);
nor U3350 (N_3350,In_3624,In_653);
or U3351 (N_3351,N_272,N_1213);
xor U3352 (N_3352,N_3105,N_3030);
nand U3353 (N_3353,N_3074,In_579);
or U3354 (N_3354,In_29,N_2878);
nor U3355 (N_3355,In_341,N_2113);
xnor U3356 (N_3356,N_35,N_3198);
or U3357 (N_3357,N_2476,N_211);
nand U3358 (N_3358,N_2947,N_1980);
and U3359 (N_3359,N_3039,N_3028);
nor U3360 (N_3360,In_1068,N_3214);
or U3361 (N_3361,In_3049,In_2964);
nor U3362 (N_3362,N_2837,N_1384);
and U3363 (N_3363,N_821,N_3230);
and U3364 (N_3364,In_1186,N_2772);
nor U3365 (N_3365,N_2946,N_3130);
nor U3366 (N_3366,N_3143,N_2040);
xnor U3367 (N_3367,In_2046,N_2832);
and U3368 (N_3368,N_2752,N_2787);
or U3369 (N_3369,In_2938,N_2751);
nand U3370 (N_3370,N_3167,In_4710);
or U3371 (N_3371,In_138,In_3515);
xnor U3372 (N_3372,N_2597,In_3221);
xor U3373 (N_3373,N_3079,N_2818);
xnor U3374 (N_3374,N_729,N_3213);
nor U3375 (N_3375,In_4177,N_1102);
nand U3376 (N_3376,N_243,N_2932);
nor U3377 (N_3377,N_2701,N_1691);
nor U3378 (N_3378,N_1218,N_2795);
nand U3379 (N_3379,In_3235,N_2889);
nand U3380 (N_3380,In_3092,In_2444);
nor U3381 (N_3381,N_3040,N_604);
nor U3382 (N_3382,N_2565,N_2052);
or U3383 (N_3383,N_2650,N_2774);
or U3384 (N_3384,In_1606,N_1653);
and U3385 (N_3385,In_4370,N_2651);
nor U3386 (N_3386,In_334,In_3657);
nand U3387 (N_3387,N_2449,In_4552);
and U3388 (N_3388,N_1870,N_3031);
nor U3389 (N_3389,N_645,N_1905);
and U3390 (N_3390,N_3047,N_1796);
nand U3391 (N_3391,N_1230,In_199);
or U3392 (N_3392,N_2314,In_386);
and U3393 (N_3393,N_2518,N_2252);
or U3394 (N_3394,N_3068,N_3076);
or U3395 (N_3395,N_2926,In_1949);
or U3396 (N_3396,In_3226,N_3033);
or U3397 (N_3397,N_3048,In_3789);
xnor U3398 (N_3398,N_923,N_2987);
or U3399 (N_3399,N_2794,N_2118);
and U3400 (N_3400,N_2391,In_4044);
nor U3401 (N_3401,In_4361,In_2116);
xnor U3402 (N_3402,N_3154,In_1895);
nand U3403 (N_3403,In_840,N_2363);
nand U3404 (N_3404,N_1640,In_943);
and U3405 (N_3405,In_4256,N_3207);
xnor U3406 (N_3406,N_3053,In_4247);
nand U3407 (N_3407,In_2548,N_387);
xnor U3408 (N_3408,N_805,N_2934);
nor U3409 (N_3409,N_1242,In_1695);
nor U3410 (N_3410,In_3022,In_3462);
and U3411 (N_3411,N_2891,N_1876);
or U3412 (N_3412,N_2095,N_1485);
nor U3413 (N_3413,N_150,N_952);
and U3414 (N_3414,N_3139,N_557);
xnor U3415 (N_3415,N_1413,N_2853);
xnor U3416 (N_3416,N_2879,N_2158);
nor U3417 (N_3417,N_2540,N_2068);
xnor U3418 (N_3418,N_2256,N_1979);
nor U3419 (N_3419,In_3476,N_2643);
nand U3420 (N_3420,In_1134,N_3110);
and U3421 (N_3421,N_2060,N_2814);
nand U3422 (N_3422,N_3085,N_2138);
or U3423 (N_3423,N_850,N_2858);
and U3424 (N_3424,N_1874,N_3070);
and U3425 (N_3425,N_1075,N_2556);
nor U3426 (N_3426,In_1650,N_1464);
xnor U3427 (N_3427,N_2025,N_3044);
and U3428 (N_3428,In_4285,N_3132);
nand U3429 (N_3429,N_2416,N_1080);
or U3430 (N_3430,N_160,In_2291);
or U3431 (N_3431,In_3320,N_2711);
xnor U3432 (N_3432,N_2587,N_3051);
nor U3433 (N_3433,N_2819,N_3072);
xnor U3434 (N_3434,N_2945,In_411);
or U3435 (N_3435,N_2707,N_2742);
nor U3436 (N_3436,N_2107,N_2981);
xor U3437 (N_3437,In_666,N_3049);
nand U3438 (N_3438,N_607,In_3951);
xor U3439 (N_3439,In_321,In_3620);
xor U3440 (N_3440,N_2385,N_2511);
xor U3441 (N_3441,In_3561,N_161);
nor U3442 (N_3442,In_1395,N_1958);
nor U3443 (N_3443,N_3095,N_1179);
or U3444 (N_3444,N_1333,N_3180);
nand U3445 (N_3445,N_1215,N_3206);
nor U3446 (N_3446,N_3151,N_2042);
nor U3447 (N_3447,N_3060,In_1144);
nand U3448 (N_3448,N_595,N_3157);
xor U3449 (N_3449,N_1564,N_2607);
or U3450 (N_3450,N_2951,N_2896);
or U3451 (N_3451,In_2722,N_3138);
and U3452 (N_3452,In_3574,N_2916);
or U3453 (N_3453,N_3220,N_1895);
nor U3454 (N_3454,In_4666,N_88);
nor U3455 (N_3455,In_4111,N_948);
nor U3456 (N_3456,N_366,N_3184);
nor U3457 (N_3457,N_2755,In_3673);
nand U3458 (N_3458,In_3722,In_4395);
nor U3459 (N_3459,N_1556,N_1747);
nand U3460 (N_3460,N_2531,N_2760);
or U3461 (N_3461,In_2667,N_3029);
nor U3462 (N_3462,N_2856,N_2675);
or U3463 (N_3463,In_3395,In_1939);
and U3464 (N_3464,N_2579,In_712);
and U3465 (N_3465,N_1964,In_4179);
or U3466 (N_3466,In_4559,N_1950);
nor U3467 (N_3467,N_3125,N_3234);
or U3468 (N_3468,N_1725,N_3147);
nand U3469 (N_3469,In_2167,N_1588);
and U3470 (N_3470,N_3187,N_2577);
nor U3471 (N_3471,N_1643,N_2618);
and U3472 (N_3472,N_2986,N_2601);
and U3473 (N_3473,N_2200,In_532);
and U3474 (N_3474,N_2110,N_257);
nor U3475 (N_3475,N_326,In_775);
nor U3476 (N_3476,In_2121,N_3010);
xnor U3477 (N_3477,N_1788,N_3249);
nand U3478 (N_3478,N_3131,N_3149);
xnor U3479 (N_3479,N_142,N_3185);
nand U3480 (N_3480,N_1771,N_3050);
nand U3481 (N_3481,In_1059,In_433);
xnor U3482 (N_3482,In_3876,In_3072);
or U3483 (N_3483,N_3032,In_4125);
nand U3484 (N_3484,N_3103,N_3065);
or U3485 (N_3485,N_1921,In_1864);
xnor U3486 (N_3486,N_3223,In_2457);
xnor U3487 (N_3487,N_3111,N_1011);
and U3488 (N_3488,N_2667,In_3370);
nand U3489 (N_3489,N_3218,N_2425);
and U3490 (N_3490,N_3086,N_445);
nor U3491 (N_3491,N_3042,N_2750);
xor U3492 (N_3492,N_605,In_2161);
nor U3493 (N_3493,N_1446,N_1085);
xor U3494 (N_3494,N_2731,N_2548);
or U3495 (N_3495,N_3117,N_2343);
or U3496 (N_3496,N_600,In_3387);
nand U3497 (N_3497,N_2957,N_1922);
nor U3498 (N_3498,N_2806,In_3329);
or U3499 (N_3499,In_1946,N_2047);
nor U3500 (N_3500,In_4476,N_3121);
and U3501 (N_3501,In_4291,N_2948);
nor U3502 (N_3502,N_1414,N_1559);
xor U3503 (N_3503,N_3316,N_2789);
or U3504 (N_3504,In_2357,In_4136);
xor U3505 (N_3505,N_2820,N_678);
or U3506 (N_3506,N_3484,N_22);
and U3507 (N_3507,N_1631,In_2315);
and U3508 (N_3508,N_743,N_3311);
or U3509 (N_3509,In_2759,N_3357);
nand U3510 (N_3510,N_2010,In_3028);
nor U3511 (N_3511,In_829,N_3078);
and U3512 (N_3512,N_3471,N_2763);
and U3513 (N_3513,N_3036,N_1822);
and U3514 (N_3514,N_3203,N_2041);
and U3515 (N_3515,N_3169,N_2654);
or U3516 (N_3516,N_2777,N_2284);
and U3517 (N_3517,In_674,N_2291);
nand U3518 (N_3518,In_1189,In_3793);
and U3519 (N_3519,N_3257,In_1444);
and U3520 (N_3520,N_2332,N_1914);
nand U3521 (N_3521,N_3430,N_3064);
or U3522 (N_3522,N_2811,N_2834);
or U3523 (N_3523,N_3400,N_3442);
nand U3524 (N_3524,N_3258,N_2691);
nor U3525 (N_3525,N_3463,N_942);
and U3526 (N_3526,N_3108,N_100);
or U3527 (N_3527,N_2971,In_2172);
and U3528 (N_3528,N_3439,N_3186);
nor U3529 (N_3529,N_1194,N_323);
nor U3530 (N_3530,In_304,N_2635);
nor U3531 (N_3531,In_1280,N_167);
xnor U3532 (N_3532,N_3035,N_2336);
nand U3533 (N_3533,N_3205,In_1904);
nor U3534 (N_3534,N_1989,N_1117);
and U3535 (N_3535,N_2998,N_846);
nor U3536 (N_3536,In_1648,N_2566);
xor U3537 (N_3537,N_3148,In_4181);
and U3538 (N_3538,N_2312,In_1313);
and U3539 (N_3539,N_2191,N_355);
nand U3540 (N_3540,In_3482,In_3039);
and U3541 (N_3541,N_3354,N_1783);
nor U3542 (N_3542,In_66,In_1272);
or U3543 (N_3543,N_3116,N_1401);
nand U3544 (N_3544,N_1740,In_3575);
nand U3545 (N_3545,N_77,In_4497);
nand U3546 (N_3546,N_3279,In_1413);
and U3547 (N_3547,In_1226,N_3374);
or U3548 (N_3548,N_3302,N_1619);
and U3549 (N_3549,In_3115,In_250);
nand U3550 (N_3550,N_2164,N_2823);
nand U3551 (N_3551,N_2283,N_2486);
xor U3552 (N_3552,N_2081,N_3487);
xnor U3553 (N_3553,N_3202,N_3159);
or U3554 (N_3554,N_2622,In_2330);
nor U3555 (N_3555,N_1752,In_703);
and U3556 (N_3556,N_2805,In_3967);
xnor U3557 (N_3557,In_2352,In_253);
or U3558 (N_3558,N_3097,In_3165);
xnor U3559 (N_3559,N_2721,In_602);
and U3560 (N_3560,In_2810,N_1731);
and U3561 (N_3561,N_189,N_3272);
nand U3562 (N_3562,In_4166,N_3290);
or U3563 (N_3563,In_729,N_2674);
nor U3564 (N_3564,N_2778,N_3080);
nor U3565 (N_3565,N_3280,N_3000);
or U3566 (N_3566,In_4919,N_2459);
xor U3567 (N_3567,N_1197,In_4339);
or U3568 (N_3568,N_3307,N_2152);
and U3569 (N_3569,N_2860,In_4083);
xor U3570 (N_3570,In_2173,N_184);
or U3571 (N_3571,N_1700,In_4543);
nor U3572 (N_3572,N_1142,In_4289);
and U3573 (N_3573,N_1781,N_3066);
nand U3574 (N_3574,N_2197,N_1098);
nand U3575 (N_3575,N_1995,N_3433);
or U3576 (N_3576,In_299,In_2822);
nor U3577 (N_3577,In_3004,In_1458);
xnor U3578 (N_3578,In_2723,N_2802);
xnor U3579 (N_3579,N_3045,N_3317);
nor U3580 (N_3580,In_447,N_2905);
and U3581 (N_3581,N_14,N_2995);
nor U3582 (N_3582,In_1320,N_2236);
and U3583 (N_3583,N_2583,N_1784);
nand U3584 (N_3584,N_1742,N_3451);
and U3585 (N_3585,N_2859,N_741);
xor U3586 (N_3586,N_591,In_2909);
nand U3587 (N_3587,In_1315,In_3341);
nand U3588 (N_3588,N_3429,N_2708);
nor U3589 (N_3589,N_1202,N_2308);
nand U3590 (N_3590,N_2238,N_2443);
or U3591 (N_3591,In_2373,In_2465);
nor U3592 (N_3592,N_3112,N_2992);
nor U3593 (N_3593,In_60,N_2949);
nand U3594 (N_3594,In_2195,N_2329);
xor U3595 (N_3595,N_2444,In_3623);
or U3596 (N_3596,In_4813,N_497);
nor U3597 (N_3597,In_4499,N_3395);
and U3598 (N_3598,N_2131,N_2182);
nor U3599 (N_3599,N_2913,N_3164);
nand U3600 (N_3600,N_1501,N_3150);
or U3601 (N_3601,N_2533,N_3351);
and U3602 (N_3602,N_3371,In_1482);
nand U3603 (N_3603,In_134,N_2237);
or U3604 (N_3604,In_2902,In_2644);
xnor U3605 (N_3605,N_2488,N_1798);
nor U3606 (N_3606,N_3289,N_3450);
or U3607 (N_3607,N_2944,N_2307);
xor U3608 (N_3608,N_3436,In_3997);
xor U3609 (N_3609,N_3104,N_2382);
nor U3610 (N_3610,N_1406,N_2870);
nor U3611 (N_3611,In_519,N_632);
xor U3612 (N_3612,N_2529,In_1308);
nand U3613 (N_3613,N_1891,N_2967);
xor U3614 (N_3614,N_2371,N_3160);
or U3615 (N_3615,N_3470,N_3347);
nor U3616 (N_3616,N_481,N_2865);
and U3617 (N_3617,N_1168,N_2776);
nand U3618 (N_3618,N_2640,N_2278);
nand U3619 (N_3619,In_1355,N_1902);
xor U3620 (N_3620,N_2925,N_1428);
and U3621 (N_3621,N_3144,In_242);
nand U3622 (N_3622,In_3554,N_1744);
and U3623 (N_3623,In_4669,N_3447);
xnor U3624 (N_3624,N_3285,N_1946);
nand U3625 (N_3625,N_3360,N_967);
and U3626 (N_3626,In_1327,In_4538);
and U3627 (N_3627,In_2364,N_3444);
and U3628 (N_3628,N_3333,In_663);
nand U3629 (N_3629,In_1489,N_3293);
xor U3630 (N_3630,N_2349,N_3263);
nand U3631 (N_3631,N_2274,In_3171);
xor U3632 (N_3632,N_3396,N_3002);
xor U3633 (N_3633,N_1746,N_3012);
nor U3634 (N_3634,N_1165,N_3262);
or U3635 (N_3635,N_2758,N_1013);
xnor U3636 (N_3636,In_4529,In_336);
and U3637 (N_3637,N_3454,N_1884);
xnor U3638 (N_3638,N_2582,N_3096);
or U3639 (N_3639,In_1054,In_1807);
and U3640 (N_3640,In_37,N_3004);
and U3641 (N_3641,N_2844,In_1604);
nand U3642 (N_3642,N_995,N_2907);
and U3643 (N_3643,N_2206,N_1229);
and U3644 (N_3644,N_3092,In_1509);
nor U3645 (N_3645,N_2759,In_2705);
xnor U3646 (N_3646,N_2712,N_3364);
or U3647 (N_3647,N_3346,N_1294);
and U3648 (N_3648,N_2952,N_2405);
and U3649 (N_3649,N_3445,N_2770);
xor U3650 (N_3650,N_3124,N_2641);
nand U3651 (N_3651,In_1782,N_173);
or U3652 (N_3652,In_4026,N_706);
nor U3653 (N_3653,N_3034,N_3310);
nand U3654 (N_3654,N_1094,N_2609);
xnor U3655 (N_3655,N_3342,In_4935);
nor U3656 (N_3656,In_135,N_810);
nor U3657 (N_3657,N_2864,N_3287);
nor U3658 (N_3658,In_3740,In_3450);
or U3659 (N_3659,In_210,N_2586);
nor U3660 (N_3660,N_3282,N_3069);
and U3661 (N_3661,N_1656,N_2426);
and U3662 (N_3662,In_4900,N_2519);
nor U3663 (N_3663,N_3422,In_856);
or U3664 (N_3664,N_3084,N_2512);
or U3665 (N_3665,In_2554,N_2431);
nor U3666 (N_3666,N_3382,N_1936);
xor U3667 (N_3667,In_1824,N_3499);
or U3668 (N_3668,In_2671,N_2590);
and U3669 (N_3669,N_2661,N_3410);
nor U3670 (N_3670,N_988,N_2127);
or U3671 (N_3671,N_3473,N_1974);
xor U3672 (N_3672,N_1797,In_883);
nor U3673 (N_3673,N_3402,N_2704);
xor U3674 (N_3674,N_3417,N_2545);
nor U3675 (N_3675,N_2495,N_2659);
nand U3676 (N_3676,N_1322,N_2881);
nor U3677 (N_3677,In_338,In_1896);
nor U3678 (N_3678,In_1974,N_3412);
and U3679 (N_3679,N_826,N_67);
nand U3680 (N_3680,N_1132,In_3683);
or U3681 (N_3681,N_3281,In_3505);
xor U3682 (N_3682,In_4493,N_2473);
or U3683 (N_3683,N_3468,N_2634);
or U3684 (N_3684,N_3120,N_3355);
nand U3685 (N_3685,N_346,In_2717);
nand U3686 (N_3686,N_3380,N_1820);
nor U3687 (N_3687,N_389,N_2833);
and U3688 (N_3688,In_1525,N_2685);
nor U3689 (N_3689,N_446,N_2988);
xor U3690 (N_3690,N_2269,N_3062);
and U3691 (N_3691,In_849,N_1390);
nand U3692 (N_3692,N_2989,N_2985);
and U3693 (N_3693,N_3179,In_2032);
and U3694 (N_3694,In_1618,In_3140);
nand U3695 (N_3695,N_2975,N_339);
and U3696 (N_3696,N_1602,In_4049);
xor U3697 (N_3697,N_3403,N_2251);
nand U3698 (N_3698,N_2528,N_2334);
nor U3699 (N_3699,N_2560,N_1065);
nor U3700 (N_3700,N_2494,N_2067);
and U3701 (N_3701,N_1090,N_3253);
xnor U3702 (N_3702,N_3330,In_3527);
xor U3703 (N_3703,N_2677,In_4947);
nand U3704 (N_3704,N_3340,In_1210);
nand U3705 (N_3705,In_194,N_838);
xnor U3706 (N_3706,N_3152,N_2761);
nand U3707 (N_3707,N_3259,N_644);
xnor U3708 (N_3708,In_385,N_1679);
nand U3709 (N_3709,In_3133,N_3250);
and U3710 (N_3710,N_345,N_804);
nand U3711 (N_3711,N_2782,N_3405);
or U3712 (N_3712,In_890,N_154);
nand U3713 (N_3713,In_4542,N_2366);
nand U3714 (N_3714,In_4741,In_2777);
nor U3715 (N_3715,N_2999,N_1641);
xor U3716 (N_3716,N_2980,N_1410);
xor U3717 (N_3717,N_2005,N_3486);
and U3718 (N_3718,N_2917,N_792);
nand U3719 (N_3719,N_2111,N_3434);
nor U3720 (N_3720,N_1270,N_1592);
and U3721 (N_3721,N_3392,N_2043);
or U3722 (N_3722,N_2993,N_2631);
nand U3723 (N_3723,N_1334,N_1572);
and U3724 (N_3724,N_2645,In_4390);
nor U3725 (N_3725,In_3152,N_3390);
xnor U3726 (N_3726,N_915,N_3498);
nor U3727 (N_3727,N_2765,N_2163);
and U3728 (N_3728,N_917,N_1055);
nor U3729 (N_3729,In_3787,N_2525);
nand U3730 (N_3730,N_1652,N_3305);
xnor U3731 (N_3731,In_417,N_1107);
and U3732 (N_3732,N_3136,In_814);
or U3733 (N_3733,N_2324,N_1185);
nand U3734 (N_3734,N_2888,N_3321);
nand U3735 (N_3735,N_2922,N_3268);
nand U3736 (N_3736,N_2275,N_3122);
and U3737 (N_3737,N_3407,N_2294);
nand U3738 (N_3738,In_1443,In_3232);
xor U3739 (N_3739,In_3542,N_2764);
nand U3740 (N_3740,N_3217,N_1105);
or U3741 (N_3741,N_3251,N_2863);
and U3742 (N_3742,N_108,N_1108);
nor U3743 (N_3743,N_2526,N_2347);
and U3744 (N_3744,N_3326,N_2709);
and U3745 (N_3745,In_4279,N_3155);
and U3746 (N_3746,N_3239,N_2575);
xor U3747 (N_3747,N_3387,N_3386);
or U3748 (N_3748,N_3014,In_4099);
nand U3749 (N_3749,N_2358,N_3465);
and U3750 (N_3750,In_1659,In_4006);
or U3751 (N_3751,N_3318,N_3441);
nand U3752 (N_3752,In_1757,N_1282);
and U3753 (N_3753,N_2447,N_3432);
and U3754 (N_3754,N_3274,N_1153);
xnor U3755 (N_3755,N_1593,In_626);
xnor U3756 (N_3756,In_4619,N_3704);
xnor U3757 (N_3757,N_3093,In_4570);
nor U3758 (N_3758,N_3539,N_3501);
and U3759 (N_3759,N_3277,N_3021);
nand U3760 (N_3760,In_2691,In_2138);
nand U3761 (N_3761,N_3722,N_757);
xnor U3762 (N_3762,N_3082,In_3776);
nor U3763 (N_3763,In_1535,N_3379);
nor U3764 (N_3764,N_2176,In_315);
xor U3765 (N_3765,N_3601,N_1932);
nor U3766 (N_3766,N_2958,N_2927);
nand U3767 (N_3767,In_1959,In_2257);
or U3768 (N_3768,N_2972,In_4623);
xor U3769 (N_3769,In_1729,N_2437);
and U3770 (N_3770,N_1919,In_526);
nand U3771 (N_3771,N_2846,In_2903);
or U3772 (N_3772,N_3332,N_3134);
nand U3773 (N_3773,N_3548,In_3990);
or U3774 (N_3774,In_821,In_891);
or U3775 (N_3775,N_1463,N_3329);
nand U3776 (N_3776,In_270,In_2728);
nand U3777 (N_3777,N_2401,In_698);
or U3778 (N_3778,N_2698,N_237);
nand U3779 (N_3779,N_2530,N_3715);
nand U3780 (N_3780,N_3691,N_3208);
nand U3781 (N_3781,N_1323,N_2147);
and U3782 (N_3782,N_3638,N_2840);
nand U3783 (N_3783,N_1806,N_3663);
and U3784 (N_3784,N_659,In_2223);
and U3785 (N_3785,N_2855,N_2306);
or U3786 (N_3786,N_149,N_3622);
nor U3787 (N_3787,In_4,N_3352);
nand U3788 (N_3788,N_3480,N_3338);
or U3789 (N_3789,In_4469,N_3313);
nor U3790 (N_3790,In_1685,In_2513);
or U3791 (N_3791,In_406,In_3209);
and U3792 (N_3792,N_3619,N_3341);
nor U3793 (N_3793,N_3176,N_3071);
nand U3794 (N_3794,N_1792,In_2180);
or U3795 (N_3795,N_3515,N_3135);
nor U3796 (N_3796,In_1234,N_3518);
nor U3797 (N_3797,N_3038,N_3531);
or U3798 (N_3798,In_4394,N_1688);
nand U3799 (N_3799,N_3276,N_1177);
or U3800 (N_3800,N_3635,N_2510);
nor U3801 (N_3801,N_3568,In_141);
xor U3802 (N_3802,N_879,N_2801);
nand U3803 (N_3803,N_3699,N_647);
nor U3804 (N_3804,In_946,N_3394);
or U3805 (N_3805,N_3481,N_2902);
and U3806 (N_3806,In_1700,N_1540);
nor U3807 (N_3807,N_2412,N_3654);
nor U3808 (N_3808,N_1138,N_3741);
or U3809 (N_3809,In_4488,N_3544);
and U3810 (N_3810,N_3497,N_3644);
nor U3811 (N_3811,N_2564,N_3181);
nor U3812 (N_3812,N_3008,N_2272);
nand U3813 (N_3813,In_3349,In_2389);
or U3814 (N_3814,N_297,In_533);
and U3815 (N_3815,N_1953,In_442);
nor U3816 (N_3816,N_3413,N_1961);
nor U3817 (N_3817,N_3046,N_2884);
nand U3818 (N_3818,N_3609,N_3648);
and U3819 (N_3819,N_3735,N_3331);
or U3820 (N_3820,N_1240,N_3631);
or U3821 (N_3821,N_2964,N_3275);
xor U3822 (N_3822,N_3594,N_1960);
and U3823 (N_3823,N_3746,N_174);
or U3824 (N_3824,N_2263,N_3001);
and U3825 (N_3825,N_1761,N_2114);
nand U3826 (N_3826,N_2966,In_2546);
and U3827 (N_3827,N_2816,N_3557);
and U3828 (N_3828,In_1281,In_4715);
or U3829 (N_3829,N_3269,N_3677);
nand U3830 (N_3830,N_3636,N_3408);
or U3831 (N_3831,N_3016,In_4478);
nand U3832 (N_3832,N_3560,In_2187);
or U3833 (N_3833,N_3409,In_4826);
and U3834 (N_3834,In_2867,N_3679);
nand U3835 (N_3835,N_3629,N_3455);
or U3836 (N_3836,N_597,N_3252);
or U3837 (N_3837,N_3511,N_3724);
or U3838 (N_3838,N_3572,N_3264);
nand U3839 (N_3839,N_3553,N_2637);
nand U3840 (N_3840,N_3423,N_2063);
or U3841 (N_3841,N_2438,In_256);
and U3842 (N_3842,N_3419,N_3689);
nand U3843 (N_3843,In_3524,N_2403);
nor U3844 (N_3844,N_3145,In_1771);
xnor U3845 (N_3845,In_2862,N_3106);
xor U3846 (N_3846,N_3694,N_344);
or U3847 (N_3847,N_2230,In_4931);
and U3848 (N_3848,N_3323,In_628);
nor U3849 (N_3849,N_3656,N_2621);
nand U3850 (N_3850,N_3547,N_3415);
and U3851 (N_3851,N_2831,N_3504);
and U3852 (N_3852,In_3334,In_3610);
xnor U3853 (N_3853,N_3492,N_3496);
nand U3854 (N_3854,In_1143,N_3165);
nand U3855 (N_3855,N_3489,In_3998);
nand U3856 (N_3856,N_3449,In_479);
xor U3857 (N_3857,N_3668,N_3438);
or U3858 (N_3858,In_177,N_3312);
and U3859 (N_3859,N_2615,In_468);
nand U3860 (N_3860,N_3461,N_2186);
or U3861 (N_3861,N_1518,N_3646);
nand U3862 (N_3862,N_2679,N_2103);
and U3863 (N_3863,In_4888,N_1585);
or U3864 (N_3864,N_2515,N_3173);
xor U3865 (N_3865,N_2557,N_3495);
nand U3866 (N_3866,In_4328,N_1553);
nor U3867 (N_3867,N_3284,N_3657);
or U3868 (N_3868,N_3491,N_3569);
nand U3869 (N_3869,N_1141,N_2930);
xor U3870 (N_3870,N_2836,In_518);
xor U3871 (N_3871,N_766,N_2994);
or U3872 (N_3872,N_3054,N_1182);
and U3873 (N_3873,N_3551,N_3582);
nand U3874 (N_3874,N_3687,In_1175);
or U3875 (N_3875,N_3098,N_3191);
xor U3876 (N_3876,In_384,N_2500);
nand U3877 (N_3877,N_3027,N_2496);
nor U3878 (N_3878,N_728,N_3140);
xnor U3879 (N_3879,In_4975,N_3005);
nor U3880 (N_3880,N_2561,N_3037);
and U3881 (N_3881,In_3631,N_2799);
xnor U3882 (N_3882,N_798,N_2785);
nand U3883 (N_3883,N_2692,N_3600);
xor U3884 (N_3884,In_1803,N_3315);
xor U3885 (N_3885,N_3260,N_2873);
and U3886 (N_3886,N_1841,N_3303);
and U3887 (N_3887,In_474,N_3188);
nand U3888 (N_3888,N_3599,N_2608);
xor U3889 (N_3889,N_3425,N_1502);
nand U3890 (N_3890,N_3261,N_3328);
nand U3891 (N_3891,N_2716,N_3651);
nand U3892 (N_3892,In_2652,N_3210);
nand U3893 (N_3893,N_3596,N_3376);
nor U3894 (N_3894,N_1948,N_3726);
nand U3895 (N_3895,N_3711,N_3562);
and U3896 (N_3896,N_1554,N_1155);
or U3897 (N_3897,N_2454,N_2990);
xnor U3898 (N_3898,In_2782,N_2265);
xnor U3899 (N_3899,N_1374,N_3665);
nand U3900 (N_3900,N_384,N_2962);
and U3901 (N_3901,N_3525,N_2572);
nor U3902 (N_3902,N_3119,N_3077);
nand U3903 (N_3903,N_3219,N_1285);
nor U3904 (N_3904,N_3649,N_2053);
and U3905 (N_3905,N_3542,In_4191);
xor U3906 (N_3906,N_390,N_3242);
nor U3907 (N_3907,N_1871,In_3494);
or U3908 (N_3908,N_2376,N_2091);
or U3909 (N_3909,N_1455,N_2729);
nor U3910 (N_3910,In_4159,N_2427);
nand U3911 (N_3911,N_2757,N_3482);
xnor U3912 (N_3912,N_2320,In_3525);
xor U3913 (N_3913,In_3451,N_2484);
nand U3914 (N_3914,N_3614,N_3081);
nor U3915 (N_3915,N_3398,N_2595);
nor U3916 (N_3916,N_3624,N_1863);
nor U3917 (N_3917,N_3411,N_3178);
nand U3918 (N_3918,N_1183,N_3306);
or U3919 (N_3919,N_3607,N_2652);
nor U3920 (N_3920,N_3059,N_3267);
xnor U3921 (N_3921,N_3123,N_2619);
or U3922 (N_3922,In_4218,N_1196);
nor U3923 (N_3923,N_2630,N_3304);
and U3924 (N_3924,In_3920,N_3254);
nand U3925 (N_3925,N_2083,N_2185);
nand U3926 (N_3926,N_3490,In_2080);
xor U3927 (N_3927,In_4521,N_3593);
or U3928 (N_3928,N_3359,N_3721);
and U3929 (N_3929,N_2753,N_3336);
or U3930 (N_3930,N_3418,N_2841);
xor U3931 (N_3931,N_1257,N_3195);
nor U3932 (N_3932,In_1913,In_605);
or U3933 (N_3933,In_2578,N_3585);
or U3934 (N_3934,N_3448,N_2135);
nor U3935 (N_3935,N_700,N_3478);
or U3936 (N_3936,N_764,In_2215);
nor U3937 (N_3937,N_3427,N_3350);
xnor U3938 (N_3938,N_3559,N_2803);
nor U3939 (N_3939,In_1900,N_2768);
xnor U3940 (N_3940,N_3113,N_3391);
nand U3941 (N_3941,N_3416,N_2783);
and U3942 (N_3942,N_3137,N_3345);
and U3943 (N_3943,N_2559,In_2361);
nand U3944 (N_3944,N_3650,N_3642);
and U3945 (N_3945,N_3550,N_3435);
nand U3946 (N_3946,In_303,N_3453);
and U3947 (N_3947,In_1198,N_1596);
and U3948 (N_3948,In_987,N_2022);
nand U3949 (N_3949,In_3410,N_3475);
or U3950 (N_3950,N_2920,N_3041);
nand U3951 (N_3951,N_2771,N_1320);
nor U3952 (N_3952,N_2638,In_1003);
xnor U3953 (N_3953,N_293,N_3697);
xor U3954 (N_3954,N_8,N_973);
or U3955 (N_3955,N_1302,N_3592);
nor U3956 (N_3956,N_3385,In_687);
nor U3957 (N_3957,In_3897,N_3196);
xor U3958 (N_3958,N_60,N_2571);
or U3959 (N_3959,N_2351,N_3710);
nor U3960 (N_3960,N_2270,In_248);
or U3961 (N_3961,N_3094,N_845);
and U3962 (N_3962,N_155,N_2432);
and U3963 (N_3963,N_3023,N_656);
or U3964 (N_3964,N_3603,N_3623);
xor U3965 (N_3965,In_3826,N_2710);
xnor U3966 (N_3966,N_3404,In_3425);
nand U3967 (N_3967,N_3535,In_1114);
nor U3968 (N_3968,N_3549,N_2415);
nor U3969 (N_3969,N_3723,N_1753);
and U3970 (N_3970,In_1894,N_2258);
xor U3971 (N_3971,In_3859,N_3707);
nor U3972 (N_3972,N_3503,N_3090);
or U3973 (N_3973,N_3381,In_1670);
and U3974 (N_3974,N_1629,N_1431);
or U3975 (N_3975,N_2756,N_1682);
and U3976 (N_3976,N_1030,N_3460);
and U3977 (N_3977,N_3373,N_3361);
and U3978 (N_3978,In_3279,N_1452);
xnor U3979 (N_3979,N_1233,N_3685);
or U3980 (N_3980,N_2784,N_2826);
nor U3981 (N_3981,N_3634,In_1672);
or U3982 (N_3982,N_3597,N_2714);
xor U3983 (N_3983,N_2189,N_3716);
and U3984 (N_3984,In_4514,N_1854);
or U3985 (N_3985,In_3384,N_1164);
and U3986 (N_3986,N_2241,N_583);
nor U3987 (N_3987,In_1813,N_3565);
and U3988 (N_3988,N_3632,N_601);
or U3989 (N_3989,N_2442,N_3667);
xor U3990 (N_3990,N_1817,In_3106);
nor U3991 (N_3991,N_1337,N_3397);
nand U3992 (N_3992,N_2226,N_3324);
and U3993 (N_3993,N_2780,In_1270);
nor U3994 (N_3994,N_2465,N_3183);
nand U3995 (N_3995,N_3502,N_2904);
nor U3996 (N_3996,N_3719,In_1940);
xnor U3997 (N_3997,N_2997,N_3567);
and U3998 (N_3998,N_2487,N_2317);
xor U3999 (N_3999,N_552,In_2711);
xnor U4000 (N_4000,N_3999,N_3906);
nor U4001 (N_4001,N_2588,N_2250);
and U4002 (N_4002,N_3291,In_1756);
or U4003 (N_4003,N_3730,In_730);
nand U4004 (N_4004,N_2523,N_3772);
or U4005 (N_4005,In_580,N_3399);
nand U4006 (N_4006,N_2215,In_2842);
nor U4007 (N_4007,N_3924,N_3944);
xnor U4008 (N_4008,N_2190,N_2322);
xor U4009 (N_4009,N_3583,N_3991);
nor U4010 (N_4010,N_3506,N_3866);
or U4011 (N_4011,N_3740,N_895);
xor U4012 (N_4012,N_502,N_3246);
xnor U4013 (N_4013,In_3075,In_576);
nand U4014 (N_4014,N_1131,N_3334);
or U4015 (N_4015,N_2876,N_3309);
and U4016 (N_4016,N_3414,N_3428);
or U4017 (N_4017,N_3314,N_2874);
xor U4018 (N_4018,N_2471,N_3467);
xor U4019 (N_4019,N_2798,N_2453);
xor U4020 (N_4020,N_3692,N_3575);
xor U4021 (N_4021,N_2074,N_3356);
and U4022 (N_4022,In_4157,N_2822);
or U4023 (N_4023,N_2850,N_65);
nor U4024 (N_4024,N_3245,N_3773);
xnor U4025 (N_4025,N_3043,N_1457);
nand U4026 (N_4026,N_1426,N_3375);
or U4027 (N_4027,N_3778,N_3885);
xor U4028 (N_4028,N_3853,N_107);
nor U4029 (N_4029,N_3940,N_3292);
or U4030 (N_4030,N_2686,N_3970);
nand U4031 (N_4031,N_3494,In_585);
and U4032 (N_4032,N_3640,In_3604);
and U4033 (N_4033,N_3814,In_1436);
and U4034 (N_4034,N_3949,In_2580);
and U4035 (N_4035,N_3680,N_3424);
nor U4036 (N_4036,N_1580,N_1612);
nand U4037 (N_4037,N_996,N_2754);
nand U4038 (N_4038,N_3891,N_2773);
xor U4039 (N_4039,N_3661,N_3020);
nor U4040 (N_4040,N_3990,N_3523);
or U4041 (N_4041,In_559,In_1760);
or U4042 (N_4042,N_3766,N_2796);
nor U4043 (N_4043,In_1379,In_1982);
nand U4044 (N_4044,N_3325,N_3876);
nand U4045 (N_4045,N_3750,N_3804);
or U4046 (N_4046,N_703,In_1292);
nand U4047 (N_4047,N_1506,N_2259);
nand U4048 (N_4048,N_2341,N_3878);
nand U4049 (N_4049,In_2634,N_3788);
nor U4050 (N_4050,N_3670,N_3946);
and U4051 (N_4051,N_3862,N_3744);
xor U4052 (N_4052,In_3381,N_3581);
nand U4053 (N_4053,N_3833,N_3231);
and U4054 (N_4054,N_1206,N_3118);
xor U4055 (N_4055,N_61,N_3658);
nor U4056 (N_4056,N_3172,N_3591);
and U4057 (N_4057,N_3856,N_2133);
or U4058 (N_4058,N_2589,N_3922);
nand U4059 (N_4059,N_3908,N_2968);
nand U4060 (N_4060,N_2480,N_580);
nand U4061 (N_4061,N_3666,N_1259);
nand U4062 (N_4062,N_3962,N_2723);
xnor U4063 (N_4063,N_3863,N_1570);
and U4064 (N_4064,N_2910,N_3483);
xnor U4065 (N_4065,N_1998,In_1724);
xor U4066 (N_4066,N_2340,N_2824);
nor U4067 (N_4067,N_3993,In_3652);
and U4068 (N_4068,In_196,N_983);
nor U4069 (N_4069,N_3011,N_3532);
or U4070 (N_4070,N_3761,In_2488);
nand U4071 (N_4071,N_1973,N_1223);
xnor U4072 (N_4072,N_738,N_3673);
nor U4073 (N_4073,N_2815,N_3851);
and U4074 (N_4074,In_2426,N_3696);
xnor U4075 (N_4075,N_3764,N_3500);
or U4076 (N_4076,N_3739,N_781);
and U4077 (N_4077,N_2648,In_790);
and U4078 (N_4078,N_3824,In_1078);
nand U4079 (N_4079,N_1604,N_3763);
xor U4080 (N_4080,N_3365,N_1698);
nand U4081 (N_4081,N_3227,N_2455);
xor U4082 (N_4082,N_3300,In_4327);
and U4083 (N_4083,N_234,N_2781);
or U4084 (N_4084,N_3779,N_3446);
and U4085 (N_4085,N_2603,N_3703);
nor U4086 (N_4086,In_1609,N_2978);
nand U4087 (N_4087,In_3073,In_189);
xnor U4088 (N_4088,N_3479,N_2970);
nor U4089 (N_4089,N_3839,N_3821);
and U4090 (N_4090,N_3780,N_1272);
nand U4091 (N_4091,N_2738,N_3298);
nand U4092 (N_4092,N_3664,N_1274);
and U4093 (N_4093,N_2893,In_1139);
nor U4094 (N_4094,N_3288,N_3626);
xor U4095 (N_4095,N_3015,N_3835);
xor U4096 (N_4096,N_2148,In_2447);
nand U4097 (N_4097,N_3630,N_3945);
nor U4098 (N_4098,In_3298,N_803);
or U4099 (N_4099,In_1654,N_3709);
nand U4100 (N_4100,N_3343,N_3605);
or U4101 (N_4101,N_2954,N_2817);
or U4102 (N_4102,N_2129,N_3327);
and U4103 (N_4103,N_3997,N_2657);
and U4104 (N_4104,N_3228,N_3948);
or U4105 (N_4105,N_1586,N_3488);
nand U4106 (N_4106,N_3832,N_3579);
nor U4107 (N_4107,N_3793,N_3530);
nand U4108 (N_4108,N_3984,N_3366);
nor U4109 (N_4109,N_3756,N_3297);
or U4110 (N_4110,N_3783,N_3571);
and U4111 (N_4111,N_3225,N_2959);
or U4112 (N_4112,N_2791,N_3753);
nand U4113 (N_4113,N_1635,N_3923);
and U4114 (N_4114,N_740,N_2788);
nor U4115 (N_4115,N_3903,N_3170);
nor U4116 (N_4116,In_4324,N_3564);
nand U4117 (N_4117,N_3212,N_640);
and U4118 (N_4118,N_2301,N_2456);
nand U4119 (N_4119,In_388,In_534);
and U4120 (N_4120,N_3823,N_3803);
and U4121 (N_4121,N_3925,N_3971);
and U4122 (N_4122,N_3714,N_3611);
nand U4123 (N_4123,N_3684,N_900);
or U4124 (N_4124,In_1076,N_1470);
nor U4125 (N_4125,N_3007,N_3980);
or U4126 (N_4126,In_2933,N_3860);
nand U4127 (N_4127,In_4766,In_4472);
nand U4128 (N_4128,N_2354,N_3896);
or U4129 (N_4129,N_3819,N_3608);
xnor U4130 (N_4130,In_4511,N_3526);
or U4131 (N_4131,N_3563,N_2479);
nand U4132 (N_4132,N_3156,N_3474);
xor U4133 (N_4133,N_81,N_1967);
and U4134 (N_4134,N_3337,N_3588);
nor U4135 (N_4135,N_3682,N_3844);
or U4136 (N_4136,N_2739,N_3998);
nand U4137 (N_4137,N_2963,N_546);
and U4138 (N_4138,N_3899,N_352);
or U4139 (N_4139,N_3941,N_2977);
or U4140 (N_4140,In_2755,N_3859);
or U4141 (N_4141,N_3892,N_3926);
or U4142 (N_4142,N_3982,N_3976);
and U4143 (N_4143,N_3826,N_3538);
nand U4144 (N_4144,In_4988,N_2536);
nand U4145 (N_4145,N_3377,N_883);
nand U4146 (N_4146,N_3247,N_66);
xor U4147 (N_4147,N_3319,N_679);
nand U4148 (N_4148,In_1596,N_3871);
nor U4149 (N_4149,N_3916,N_1840);
nand U4150 (N_4150,N_3517,N_3075);
nand U4151 (N_4151,N_3905,N_3848);
nor U4152 (N_4152,In_3399,N_3485);
xnor U4153 (N_4153,N_3615,N_2809);
nand U4154 (N_4154,N_3701,In_3879);
xnor U4155 (N_4155,N_3956,N_3362);
and U4156 (N_4156,In_2960,N_1966);
or U4157 (N_4157,In_4575,N_3299);
nand U4158 (N_4158,In_1772,N_2943);
or U4159 (N_4159,In_3692,N_3917);
and U4160 (N_4160,N_3929,N_3987);
nor U4161 (N_4161,N_3224,N_3963);
nor U4162 (N_4162,N_3769,N_539);
and U4163 (N_4163,N_3979,N_1303);
or U4164 (N_4164,N_3637,N_3974);
nor U4165 (N_4165,In_4929,N_3919);
or U4166 (N_4166,N_3939,N_3883);
nand U4167 (N_4167,N_3100,N_3736);
and U4168 (N_4168,N_3977,N_3602);
xor U4169 (N_4169,N_774,N_3728);
and U4170 (N_4170,N_2115,In_3101);
nor U4171 (N_4171,N_3469,In_4910);
nand U4172 (N_4172,In_2351,N_3864);
nor U4173 (N_4173,N_3477,N_655);
or U4174 (N_4174,N_3109,N_2810);
nor U4175 (N_4175,N_3690,N_3706);
nor U4176 (N_4176,N_3785,N_1712);
nor U4177 (N_4177,In_4365,N_3850);
xor U4178 (N_4178,N_3529,N_3505);
nand U4179 (N_4179,In_114,N_3828);
nor U4180 (N_4180,N_3126,N_3796);
nand U4181 (N_4181,N_3759,N_3570);
and U4182 (N_4182,N_3792,N_3545);
or U4183 (N_4183,N_2821,In_3360);
or U4184 (N_4184,N_3683,N_3063);
or U4185 (N_4185,N_3055,N_2984);
nand U4186 (N_4186,N_553,N_2350);
and U4187 (N_4187,N_3513,N_3909);
or U4188 (N_4188,N_3762,N_3236);
and U4189 (N_4189,N_1190,N_3627);
or U4190 (N_4190,N_2665,N_3367);
xor U4191 (N_4191,N_3652,N_2474);
nor U4192 (N_4192,N_3729,N_2898);
or U4193 (N_4193,N_3003,N_2825);
xnor U4194 (N_4194,N_3508,In_436);
nor U4195 (N_4195,N_3431,N_3786);
nand U4196 (N_4196,N_3443,In_1541);
nor U4197 (N_4197,In_2825,In_3043);
and U4198 (N_4198,N_2996,In_4987);
nand U4199 (N_4199,In_3014,N_26);
nand U4200 (N_4200,N_3774,N_1621);
xnor U4201 (N_4201,In_4143,In_3817);
nand U4202 (N_4202,N_3872,N_3017);
or U4203 (N_4203,In_1861,N_3493);
and U4204 (N_4204,N_3587,N_3808);
nor U4205 (N_4205,N_3363,N_3755);
nor U4206 (N_4206,N_3590,N_3958);
xnor U4207 (N_4207,N_3519,N_3388);
and U4208 (N_4208,In_2419,N_1224);
or U4209 (N_4209,In_1879,N_3737);
nand U4210 (N_4210,N_2551,N_3934);
and U4211 (N_4211,N_1830,N_3889);
nor U4212 (N_4212,In_1241,N_3286);
xor U4213 (N_4213,N_3947,N_3921);
nand U4214 (N_4214,N_1199,N_3464);
and U4215 (N_4215,N_3880,N_1208);
nand U4216 (N_4216,N_1434,N_3528);
nand U4217 (N_4217,N_3022,N_3128);
nand U4218 (N_4218,N_3742,N_3801);
or U4219 (N_4219,N_3904,N_2253);
xor U4220 (N_4220,N_3641,N_3320);
nor U4221 (N_4221,N_2472,N_3854);
xor U4222 (N_4222,N_3731,N_3595);
or U4223 (N_4223,N_3915,N_3552);
or U4224 (N_4224,In_93,N_3695);
nor U4225 (N_4225,N_3957,N_3073);
nor U4226 (N_4226,N_3985,N_2273);
nor U4227 (N_4227,N_3758,N_3784);
nand U4228 (N_4228,In_1295,N_2249);
nand U4229 (N_4229,N_2077,N_2174);
or U4230 (N_4230,In_536,N_2049);
xor U4231 (N_4231,N_3426,In_2889);
nand U4232 (N_4232,N_3527,N_2394);
xor U4233 (N_4233,In_3803,N_3265);
xor U4234 (N_4234,N_3782,N_3700);
and U4235 (N_4235,In_3427,N_3561);
xnor U4236 (N_4236,N_3865,N_3466);
nand U4237 (N_4237,N_3886,N_3368);
xor U4238 (N_4238,N_1558,N_3830);
and U4239 (N_4239,N_3747,N_2829);
xnor U4240 (N_4240,N_3512,N_3943);
nor U4241 (N_4241,In_4101,In_1277);
nor U4242 (N_4242,N_2406,N_3456);
nor U4243 (N_4243,N_3770,N_2467);
and U4244 (N_4244,N_3767,N_3937);
nand U4245 (N_4245,N_588,N_1514);
and U4246 (N_4246,In_717,In_1645);
and U4247 (N_4247,N_380,N_3760);
nor U4248 (N_4248,N_2214,N_3838);
and U4249 (N_4249,N_3791,N_3842);
xor U4250 (N_4250,N_3083,N_3089);
xor U4251 (N_4251,N_4025,N_3541);
or U4252 (N_4252,N_4157,N_3734);
xor U4253 (N_4253,N_4178,N_2228);
xnor U4254 (N_4254,In_581,N_3831);
xnor U4255 (N_4255,N_3867,N_4014);
xnor U4256 (N_4256,N_3175,N_4056);
xor U4257 (N_4257,N_4105,N_4104);
nand U4258 (N_4258,N_3221,N_3161);
xor U4259 (N_4259,N_4180,N_3672);
nor U4260 (N_4260,N_4159,N_4082);
nand U4261 (N_4261,N_4218,N_1852);
xor U4262 (N_4262,In_3080,N_3882);
nand U4263 (N_4263,N_3777,N_837);
and U4264 (N_4264,N_2446,N_2368);
xor U4265 (N_4265,N_4030,N_3358);
and U4266 (N_4266,N_4068,N_4013);
nand U4267 (N_4267,N_3705,N_4215);
xnor U4268 (N_4268,N_3166,N_3510);
xor U4269 (N_4269,N_3806,N_4031);
nor U4270 (N_4270,N_3845,N_4156);
or U4271 (N_4271,In_1546,N_28);
xnor U4272 (N_4272,N_3676,N_4016);
xnor U4273 (N_4273,N_1415,N_3353);
nand U4274 (N_4274,In_2983,N_4073);
nand U4275 (N_4275,N_581,N_1499);
nand U4276 (N_4276,N_1947,N_4120);
nand U4277 (N_4277,N_3322,N_4048);
xnor U4278 (N_4278,N_2717,In_2940);
nor U4279 (N_4279,N_4080,N_1595);
and U4280 (N_4280,N_2610,N_4119);
nor U4281 (N_4281,N_4233,N_3674);
nor U4282 (N_4282,N_3524,In_4077);
nand U4283 (N_4283,N_1838,N_3836);
or U4284 (N_4284,N_4221,N_1349);
or U4285 (N_4285,N_4111,N_4000);
nor U4286 (N_4286,N_4147,N_4152);
and U4287 (N_4287,N_4245,N_2666);
nand U4288 (N_4288,N_3757,N_2628);
nand U4289 (N_4289,N_4179,N_2664);
and U4290 (N_4290,In_3414,N_4219);
xor U4291 (N_4291,N_3344,N_4187);
xnor U4292 (N_4292,N_3847,N_4063);
nand U4293 (N_4293,N_2145,N_4032);
xnor U4294 (N_4294,N_3610,N_4039);
and U4295 (N_4295,N_1770,N_4019);
xnor U4296 (N_4296,N_3516,N_3554);
nor U4297 (N_4297,N_4130,N_3574);
or U4298 (N_4298,N_3255,N_3789);
nand U4299 (N_4299,N_3900,N_4064);
nand U4300 (N_4300,N_4198,N_4185);
nor U4301 (N_4301,N_4024,N_3975);
nor U4302 (N_4302,N_1733,N_4070);
nand U4303 (N_4303,N_4239,N_4047);
and U4304 (N_4304,N_3911,N_1803);
and U4305 (N_4305,In_176,N_494);
and U4306 (N_4306,N_4043,N_4226);
xor U4307 (N_4307,N_3702,N_3809);
nand U4308 (N_4308,N_3308,N_3056);
nand U4309 (N_4309,N_4225,N_3389);
nand U4310 (N_4310,N_2965,N_3846);
nand U4311 (N_4311,N_2367,N_3986);
xor U4312 (N_4312,N_3712,N_3653);
xnor U4313 (N_4313,N_2689,N_586);
or U4314 (N_4314,N_3969,N_3520);
nand U4315 (N_4315,N_3238,N_3827);
and U4316 (N_4316,N_4011,N_4055);
nor U4317 (N_4317,N_4247,N_4141);
or U4318 (N_4318,N_4075,N_2581);
and U4319 (N_4319,N_3910,N_4136);
and U4320 (N_4320,N_4089,N_4217);
and U4321 (N_4321,N_3018,N_4134);
or U4322 (N_4322,N_3812,N_3678);
nand U4323 (N_4323,N_4126,N_4027);
and U4324 (N_4324,In_115,N_1607);
xor U4325 (N_4325,N_3509,N_4057);
nor U4326 (N_4326,N_3820,N_2901);
nand U4327 (N_4327,N_1676,N_1437);
nand U4328 (N_4328,N_2414,In_1811);
or U4329 (N_4329,N_2656,N_4172);
and U4330 (N_4330,N_4087,In_624);
or U4331 (N_4331,N_3967,N_1167);
or U4332 (N_4332,N_4238,N_2378);
nand U4333 (N_4333,In_4294,N_3912);
or U4334 (N_4334,N_4022,N_3476);
nor U4335 (N_4335,N_3966,N_4021);
nand U4336 (N_4336,N_3981,N_3273);
and U4337 (N_4337,N_4138,N_3618);
nor U4338 (N_4338,N_1417,N_3874);
and U4339 (N_4339,N_3718,N_4200);
nand U4340 (N_4340,N_342,N_3142);
nor U4341 (N_4341,N_4145,N_2216);
nand U4342 (N_4342,N_3717,N_4206);
or U4343 (N_4343,In_1842,N_3813);
and U4344 (N_4344,In_1806,N_3625);
nand U4345 (N_4345,N_3894,N_3266);
nor U4346 (N_4346,N_4093,N_4175);
xnor U4347 (N_4347,N_3877,N_4220);
nor U4348 (N_4348,N_3182,N_3875);
nand U4349 (N_4349,In_2998,In_881);
or U4350 (N_4350,N_4208,N_4094);
or U4351 (N_4351,N_4090,N_3931);
nor U4352 (N_4352,N_567,N_4069);
and U4353 (N_4353,N_3537,N_2050);
nor U4354 (N_4354,N_3961,N_3805);
nor U4355 (N_4355,N_3177,N_3861);
nand U4356 (N_4356,N_3959,N_4146);
nand U4357 (N_4357,N_3887,N_3163);
xnor U4358 (N_4358,In_948,In_3416);
and U4359 (N_4359,N_4081,N_3995);
or U4360 (N_4360,N_3713,N_3606);
xor U4361 (N_4361,N_3749,N_3339);
nor U4362 (N_4362,N_3158,N_4211);
or U4363 (N_4363,N_3514,N_2154);
nand U4364 (N_4364,N_3816,N_3781);
xor U4365 (N_4365,N_4121,N_3522);
nand U4366 (N_4366,N_3153,In_179);
nand U4367 (N_4367,N_4045,N_3727);
nor U4368 (N_4368,N_2699,N_3655);
or U4369 (N_4369,N_3914,N_4041);
and U4370 (N_4370,N_3586,N_412);
and U4371 (N_4371,N_2054,N_3589);
and U4372 (N_4372,N_4097,N_4052);
and U4373 (N_4373,N_4106,N_4113);
xnor U4374 (N_4374,In_2845,N_4015);
and U4375 (N_4375,N_4053,N_4139);
nor U4376 (N_4376,N_4199,N_4046);
nand U4377 (N_4377,N_3613,In_1110);
or U4378 (N_4378,N_3099,N_4148);
xnor U4379 (N_4379,N_4065,N_3204);
xor U4380 (N_4380,N_3229,N_1266);
and U4381 (N_4381,N_4129,N_3199);
and U4382 (N_4382,In_3944,N_4029);
xnor U4383 (N_4383,N_3754,N_3988);
nor U4384 (N_4384,N_3401,N_3840);
nand U4385 (N_4385,In_4460,N_4223);
nand U4386 (N_4386,N_4210,N_3837);
or U4387 (N_4387,N_3301,N_3973);
or U4388 (N_4388,N_3459,N_4083);
and U4389 (N_4389,N_3645,N_3420);
xnor U4390 (N_4390,N_3660,In_3682);
and U4391 (N_4391,N_3393,N_4051);
xnor U4392 (N_4392,In_3051,In_909);
xor U4393 (N_4393,N_4244,N_3771);
nor U4394 (N_4394,N_3879,N_4209);
and U4395 (N_4395,N_3129,In_4153);
nor U4396 (N_4396,N_4164,N_4192);
xor U4397 (N_4397,In_4582,N_3953);
or U4398 (N_4398,N_2861,N_2119);
and U4399 (N_4399,N_3598,N_41);
or U4400 (N_4400,N_1503,N_3732);
nor U4401 (N_4401,N_3669,N_3462);
and U4402 (N_4402,N_4229,N_4143);
nor U4403 (N_4403,N_3536,N_3647);
xor U4404 (N_4404,N_4132,N_3932);
nor U4405 (N_4405,In_3744,In_1539);
and U4406 (N_4406,N_2931,N_1659);
and U4407 (N_4407,N_3534,N_4144);
nand U4408 (N_4408,N_4067,N_4099);
and U4409 (N_4409,N_3873,In_1271);
nor U4410 (N_4410,N_4074,N_3901);
xor U4411 (N_4411,N_3802,N_3372);
nand U4412 (N_4412,N_4140,N_4118);
xor U4413 (N_4413,N_3720,N_3576);
nor U4414 (N_4414,N_3457,In_3345);
nand U4415 (N_4415,N_2198,N_4033);
and U4416 (N_4416,N_2124,N_3918);
xnor U4417 (N_4417,N_2375,N_4177);
or U4418 (N_4418,N_3643,N_4040);
nor U4419 (N_4419,N_4214,N_4004);
xor U4420 (N_4420,N_3989,N_3628);
nor U4421 (N_4421,N_2682,N_3843);
xor U4422 (N_4422,N_3951,N_3295);
nand U4423 (N_4423,In_1785,N_4084);
nand U4424 (N_4424,In_4277,N_4190);
and U4425 (N_4425,N_3348,N_4028);
nand U4426 (N_4426,N_2282,N_3440);
nand U4427 (N_4427,N_3810,N_4103);
and U4428 (N_4428,N_3211,N_4194);
xnor U4429 (N_4429,N_4249,N_3633);
or U4430 (N_4430,N_3797,N_3868);
nor U4431 (N_4431,N_3890,N_3458);
and U4432 (N_4432,In_1016,In_3650);
and U4433 (N_4433,In_267,N_4008);
xnor U4434 (N_4434,N_4037,N_2808);
nor U4435 (N_4435,N_4154,In_4742);
or U4436 (N_4436,N_3708,N_3190);
nor U4437 (N_4437,N_2470,N_3964);
and U4438 (N_4438,N_1920,In_131);
and U4439 (N_4439,N_3751,N_4163);
xor U4440 (N_4440,N_3936,In_2888);
nand U4441 (N_4441,N_3671,N_4241);
xnor U4442 (N_4442,N_3927,N_4231);
and U4443 (N_4443,N_3996,N_3620);
and U4444 (N_4444,N_3546,N_4191);
or U4445 (N_4445,In_290,N_2923);
nor U4446 (N_4446,N_3738,N_571);
xnor U4447 (N_4447,N_4079,N_4034);
xnor U4448 (N_4448,N_4171,N_4169);
xor U4449 (N_4449,N_3384,In_1561);
nor U4450 (N_4450,N_3834,N_1563);
xor U4451 (N_4451,N_3107,In_4605);
nor U4452 (N_4452,N_3870,N_2940);
or U4453 (N_4453,N_4213,N_4151);
and U4454 (N_4454,N_3913,N_4222);
xnor U4455 (N_4455,N_4124,N_3938);
or U4456 (N_4456,N_4009,N_209);
xnor U4457 (N_4457,N_3621,N_3270);
xnor U4458 (N_4458,N_4062,N_3209);
nor U4459 (N_4459,N_4110,N_3693);
nor U4460 (N_4460,N_4243,In_3131);
xor U4461 (N_4461,N_4224,N_3725);
nand U4462 (N_4462,N_3168,N_2939);
nand U4463 (N_4463,In_4137,N_4150);
nor U4464 (N_4464,N_4205,N_3577);
and U4465 (N_4465,N_3688,N_3950);
and U4466 (N_4466,N_4212,In_621);
or U4467 (N_4467,N_4060,N_3194);
nand U4468 (N_4468,In_662,In_2615);
nor U4469 (N_4469,N_4189,N_4168);
and U4470 (N_4470,In_903,N_2335);
nor U4471 (N_4471,N_4193,N_1692);
or U4472 (N_4472,N_4042,N_3807);
nor U4473 (N_4473,N_3799,N_4230);
nand U4474 (N_4474,N_3675,N_3825);
and U4475 (N_4475,N_2839,N_3849);
or U4476 (N_4476,N_4100,N_4115);
or U4477 (N_4477,N_4125,N_4137);
nor U4478 (N_4478,N_4161,N_4086);
xor U4479 (N_4479,In_2186,N_4149);
nor U4480 (N_4480,N_4162,N_4195);
xnor U4481 (N_4481,N_3815,N_235);
nor U4482 (N_4482,N_3617,N_4173);
nand U4483 (N_4483,N_3765,N_2935);
and U4484 (N_4484,N_2524,N_4101);
nand U4485 (N_4485,N_3141,N_4122);
or U4486 (N_4486,N_3869,N_2745);
nand U4487 (N_4487,N_3556,N_3942);
nor U4488 (N_4488,In_3472,N_2591);
or U4489 (N_4489,N_4092,In_272);
xor U4490 (N_4490,N_4088,N_3822);
or U4491 (N_4491,N_501,N_3580);
nand U4492 (N_4492,N_4174,N_3768);
or U4493 (N_4493,In_4606,In_3313);
nand U4494 (N_4494,N_4228,In_3799);
or U4495 (N_4495,N_4182,N_1378);
and U4496 (N_4496,N_4114,N_3558);
nand U4497 (N_4497,N_3841,N_3256);
xor U4498 (N_4498,N_4098,N_3698);
nand U4499 (N_4499,N_3920,N_3133);
or U4500 (N_4500,N_4496,In_766);
nor U4501 (N_4501,N_4452,N_4440);
xor U4502 (N_4502,N_4361,N_4476);
or U4503 (N_4503,N_4326,N_4197);
nor U4504 (N_4504,N_3533,N_3573);
nand U4505 (N_4505,N_3930,N_3829);
xnor U4506 (N_4506,N_3244,N_4409);
xor U4507 (N_4507,N_4320,N_2106);
or U4508 (N_4508,N_4422,N_4256);
xor U4509 (N_4509,N_4232,N_1802);
xnor U4510 (N_4510,N_3335,N_4253);
or U4511 (N_4511,N_4466,In_1818);
and U4512 (N_4512,N_3057,N_4324);
nand U4513 (N_4513,N_2668,N_4072);
nor U4514 (N_4514,N_3743,N_4417);
xor U4515 (N_4515,N_1547,N_4313);
nor U4516 (N_4516,N_4300,N_4419);
nand U4517 (N_4517,N_4304,N_4462);
or U4518 (N_4518,N_4376,N_4349);
or U4519 (N_4519,N_31,N_3795);
nor U4520 (N_4520,N_4434,N_3935);
or U4521 (N_4521,N_4380,In_2456);
nand U4522 (N_4522,N_4456,N_4006);
nor U4523 (N_4523,N_4494,N_4003);
nand U4524 (N_4524,N_4095,N_4330);
or U4525 (N_4525,N_3965,N_4420);
and U4526 (N_4526,N_4390,N_3811);
nor U4527 (N_4527,N_4316,N_4254);
nand U4528 (N_4528,N_4305,N_4428);
or U4529 (N_4529,N_4309,N_4468);
xnor U4530 (N_4530,N_3787,N_4007);
xor U4531 (N_4531,N_3893,N_4275);
nand U4532 (N_4532,N_3162,N_3521);
nor U4533 (N_4533,N_4360,N_4471);
xnor U4534 (N_4534,N_4435,N_3283);
and U4535 (N_4535,N_4281,N_4319);
nand U4536 (N_4536,N_4259,N_2544);
and U4537 (N_4537,N_4176,N_4481);
nor U4538 (N_4538,N_4050,N_4289);
and U4539 (N_4539,N_4499,N_4017);
or U4540 (N_4540,N_4354,N_4166);
xor U4541 (N_4541,In_1056,N_4477);
and U4542 (N_4542,N_3174,N_3378);
xor U4543 (N_4543,N_4448,N_3240);
nor U4544 (N_4544,N_3296,N_4425);
or U4545 (N_4545,N_1287,N_4450);
or U4546 (N_4546,N_4387,N_3955);
or U4547 (N_4547,N_4290,N_4285);
xnor U4548 (N_4548,N_3349,N_4272);
and U4549 (N_4549,N_4077,N_4498);
or U4550 (N_4550,N_4299,N_3604);
or U4551 (N_4551,N_3960,N_4381);
nor U4552 (N_4552,N_3555,N_3994);
nand U4553 (N_4553,N_1872,N_4475);
nor U4554 (N_4554,N_2690,N_4342);
nor U4555 (N_4555,N_4373,N_4268);
or U4556 (N_4556,N_4356,N_4474);
nor U4557 (N_4557,N_4372,N_3566);
nand U4558 (N_4558,N_4375,N_4283);
nand U4559 (N_4559,N_3983,N_4461);
xor U4560 (N_4560,N_3472,N_4418);
or U4561 (N_4561,N_4485,N_3800);
or U4562 (N_4562,N_4398,N_4273);
nand U4563 (N_4563,N_4407,N_3662);
xnor U4564 (N_4564,N_4394,N_4287);
and U4565 (N_4565,N_4374,N_4447);
and U4566 (N_4566,N_4066,N_1026);
nor U4567 (N_4567,N_4405,N_4449);
xnor U4568 (N_4568,N_773,N_4339);
nand U4569 (N_4569,N_3968,N_4085);
or U4570 (N_4570,N_4061,N_4196);
or U4571 (N_4571,N_4391,N_4023);
nor U4572 (N_4572,N_3540,N_4184);
xnor U4573 (N_4573,N_4363,N_2015);
nor U4574 (N_4574,N_4001,N_2033);
nand U4575 (N_4575,N_4167,N_3681);
and U4576 (N_4576,N_4453,N_3578);
xor U4577 (N_4577,N_4492,N_4020);
and U4578 (N_4578,N_4250,In_713);
or U4579 (N_4579,N_4260,N_4385);
or U4580 (N_4580,N_4463,N_4411);
nand U4581 (N_4581,N_4329,N_4044);
nand U4582 (N_4582,N_4446,N_4227);
and U4583 (N_4583,N_2527,N_3790);
nand U4584 (N_4584,N_4333,N_4059);
nand U4585 (N_4585,N_4302,N_2748);
or U4586 (N_4586,N_4408,N_4382);
and U4587 (N_4587,N_3006,N_4251);
nand U4588 (N_4588,N_4237,N_4142);
nor U4589 (N_4589,N_4345,N_3659);
xnor U4590 (N_4590,N_4403,In_2931);
xnor U4591 (N_4591,N_4441,In_1873);
or U4592 (N_4592,N_4383,N_3102);
nand U4593 (N_4593,N_2080,N_4308);
or U4594 (N_4594,N_4038,N_4341);
or U4595 (N_4595,N_3406,N_4160);
and U4596 (N_4596,N_3933,N_4005);
xor U4597 (N_4597,N_4340,In_4393);
or U4598 (N_4598,N_4423,N_4467);
xnor U4599 (N_4599,N_4311,N_4413);
or U4600 (N_4600,N_144,N_3437);
and U4601 (N_4601,N_4303,N_1436);
nor U4602 (N_4602,N_4343,N_4002);
nand U4603 (N_4603,N_1649,N_4076);
or U4604 (N_4604,N_4116,N_4128);
xor U4605 (N_4605,N_3612,N_4306);
xor U4606 (N_4606,N_3383,N_4433);
and U4607 (N_4607,N_4344,N_4410);
nand U4608 (N_4608,N_4264,N_3271);
nand U4609 (N_4609,In_4203,N_3897);
xnor U4610 (N_4610,N_3775,N_3745);
xnor U4611 (N_4611,N_4203,N_4202);
or U4612 (N_4612,N_4258,N_4183);
or U4613 (N_4613,N_3992,N_4386);
and U4614 (N_4614,In_3858,N_4439);
xor U4615 (N_4615,N_3507,N_4277);
nand U4616 (N_4616,N_4350,N_2924);
xnor U4617 (N_4617,N_4271,N_4135);
nor U4618 (N_4618,N_2493,N_833);
and U4619 (N_4619,N_3733,N_4323);
nand U4620 (N_4620,N_1380,N_3895);
nor U4621 (N_4621,N_4480,N_3884);
nand U4622 (N_4622,N_4388,N_4487);
nor U4623 (N_4623,N_3421,N_1516);
nor U4624 (N_4624,N_1845,N_4416);
xnor U4625 (N_4625,N_4133,N_4310);
and U4626 (N_4626,N_4378,In_4319);
xnor U4627 (N_4627,N_3817,N_4401);
and U4628 (N_4628,N_4443,In_2625);
xnor U4629 (N_4629,N_3978,N_4454);
nand U4630 (N_4630,N_4325,N_4207);
nand U4631 (N_4631,N_4488,N_3776);
xnor U4632 (N_4632,N_4445,N_4318);
or U4633 (N_4633,N_3752,N_4370);
nand U4634 (N_4634,N_3294,N_4400);
or U4635 (N_4635,N_3954,N_2276);
nor U4636 (N_4636,N_3237,N_4109);
xor U4637 (N_4637,N_3748,N_3907);
nor U4638 (N_4638,N_4357,N_4314);
or U4639 (N_4639,N_4131,N_4444);
nor U4640 (N_4640,N_4054,N_2680);
nand U4641 (N_4641,N_4483,N_4397);
xor U4642 (N_4642,N_4255,N_4336);
nand U4643 (N_4643,N_4108,N_2009);
and U4644 (N_4644,N_4071,N_3972);
and U4645 (N_4645,N_3369,N_2379);
xor U4646 (N_4646,N_3855,N_3798);
xnor U4647 (N_4647,N_4406,N_3686);
xor U4648 (N_4648,N_4248,N_1278);
nand U4649 (N_4649,N_4035,N_4235);
xor U4650 (N_4650,N_4186,In_831);
and U4651 (N_4651,N_4412,N_4489);
nand U4652 (N_4652,N_4497,N_4430);
nor U4653 (N_4653,N_3818,N_4276);
nand U4654 (N_4654,N_4392,N_4355);
xor U4655 (N_4655,N_4460,N_4379);
nor U4656 (N_4656,N_4393,N_4246);
nor U4657 (N_4657,N_4389,N_4337);
nor U4658 (N_4658,N_3898,N_4335);
nand U4659 (N_4659,N_4096,N_4451);
or U4660 (N_4660,N_4295,N_4091);
nor U4661 (N_4661,N_3858,N_4490);
nor U4662 (N_4662,N_3278,N_4181);
xor U4663 (N_4663,N_2139,N_4493);
and U4664 (N_4664,N_4297,N_4424);
nor U4665 (N_4665,N_3452,N_4464);
or U4666 (N_4666,N_1813,N_4365);
nor U4667 (N_4667,N_3952,N_4322);
xor U4668 (N_4668,N_4472,N_4455);
and U4669 (N_4669,N_4155,In_2775);
xor U4670 (N_4670,N_2979,N_4236);
xor U4671 (N_4671,N_566,N_2156);
nand U4672 (N_4672,N_4296,N_4367);
nand U4673 (N_4673,N_4482,N_4352);
or U4674 (N_4674,N_3928,N_4058);
and U4675 (N_4675,N_4078,N_4284);
or U4676 (N_4676,N_2624,N_1396);
and U4677 (N_4677,N_4036,N_4368);
xor U4678 (N_4678,N_4112,N_4123);
xor U4679 (N_4679,N_4384,N_2882);
xnor U4680 (N_4680,In_931,N_4404);
nor U4681 (N_4681,N_4470,N_4267);
or U4682 (N_4682,N_4312,In_4147);
nand U4683 (N_4683,N_4286,N_4458);
and U4684 (N_4684,N_4331,N_4315);
and U4685 (N_4685,N_4421,N_4399);
or U4686 (N_4686,N_4240,N_4469);
or U4687 (N_4687,In_1301,N_4321);
and U4688 (N_4688,N_4351,N_4457);
nor U4689 (N_4689,N_4263,N_4334);
xnor U4690 (N_4690,N_4479,N_4338);
xnor U4691 (N_4691,N_4280,N_2483);
xnor U4692 (N_4692,N_4436,N_1352);
nand U4693 (N_4693,N_4442,N_4465);
nand U4694 (N_4694,N_3616,N_4327);
nand U4695 (N_4695,N_3888,N_4362);
nand U4696 (N_4696,N_3902,N_4204);
and U4697 (N_4697,N_4294,N_4117);
xnor U4698 (N_4698,N_4364,N_4288);
xnor U4699 (N_4699,N_3235,N_4158);
nor U4700 (N_4700,N_4396,N_4366);
xnor U4701 (N_4701,N_4346,N_3857);
or U4702 (N_4702,N_4307,N_2605);
nand U4703 (N_4703,N_4358,N_4270);
nand U4704 (N_4704,N_2149,N_3019);
nand U4705 (N_4705,N_4026,N_4153);
xor U4706 (N_4706,In_2368,N_4415);
or U4707 (N_4707,N_4301,N_4495);
xnor U4708 (N_4708,N_4216,N_3584);
nor U4709 (N_4709,N_2842,N_4353);
xor U4710 (N_4710,N_4459,N_4347);
or U4711 (N_4711,N_2887,N_1042);
or U4712 (N_4712,N_1562,N_4427);
and U4713 (N_4713,N_4473,N_4107);
nor U4714 (N_4714,N_4201,N_4429);
nand U4715 (N_4715,N_4348,N_4274);
xor U4716 (N_4716,N_4165,N_4328);
and U4717 (N_4717,N_4377,N_3852);
xor U4718 (N_4718,N_4491,N_3881);
or U4719 (N_4719,In_3048,N_4188);
nand U4720 (N_4720,N_4359,N_4414);
nand U4721 (N_4721,In_2391,N_4486);
and U4722 (N_4722,N_4269,N_4282);
xor U4723 (N_4723,N_4170,N_4371);
nor U4724 (N_4724,N_4332,N_4298);
and U4725 (N_4725,N_3101,N_4292);
and U4726 (N_4726,N_2767,N_2386);
nand U4727 (N_4727,N_2866,N_2435);
or U4728 (N_4728,In_3875,N_4402);
or U4729 (N_4729,N_4478,N_3794);
xor U4730 (N_4730,N_4261,N_4010);
or U4731 (N_4731,In_313,N_4426);
or U4732 (N_4732,N_4438,N_4252);
nand U4733 (N_4733,N_4432,N_727);
nand U4734 (N_4734,N_4395,N_4279);
or U4735 (N_4735,N_4369,N_3088);
nand U4736 (N_4736,N_3639,N_4012);
nand U4737 (N_4737,N_4102,In_3454);
xor U4738 (N_4738,N_4293,N_4431);
nand U4739 (N_4739,N_2960,N_4265);
nand U4740 (N_4740,N_1014,N_3201);
nor U4741 (N_4741,N_4257,N_4049);
xor U4742 (N_4742,N_4266,N_4317);
nor U4743 (N_4743,N_4127,In_778);
nand U4744 (N_4744,N_4262,N_1900);
xnor U4745 (N_4745,N_4018,N_3543);
or U4746 (N_4746,N_3370,N_4242);
xor U4747 (N_4747,N_4437,N_4484);
and U4748 (N_4748,In_4309,N_4278);
or U4749 (N_4749,N_4234,N_4291);
nor U4750 (N_4750,N_4706,N_4707);
or U4751 (N_4751,N_4630,N_4743);
and U4752 (N_4752,N_4702,N_4580);
and U4753 (N_4753,N_4593,N_4744);
or U4754 (N_4754,N_4546,N_4604);
xnor U4755 (N_4755,N_4688,N_4620);
or U4756 (N_4756,N_4575,N_4747);
or U4757 (N_4757,N_4663,N_4689);
nand U4758 (N_4758,N_4590,N_4556);
nor U4759 (N_4759,N_4699,N_4548);
nor U4760 (N_4760,N_4729,N_4660);
xor U4761 (N_4761,N_4700,N_4724);
and U4762 (N_4762,N_4639,N_4540);
xor U4763 (N_4763,N_4661,N_4645);
xor U4764 (N_4764,N_4682,N_4643);
and U4765 (N_4765,N_4693,N_4587);
xnor U4766 (N_4766,N_4670,N_4683);
xnor U4767 (N_4767,N_4500,N_4579);
or U4768 (N_4768,N_4685,N_4603);
or U4769 (N_4769,N_4710,N_4654);
or U4770 (N_4770,N_4733,N_4674);
or U4771 (N_4771,N_4607,N_4749);
xnor U4772 (N_4772,N_4555,N_4505);
nand U4773 (N_4773,N_4602,N_4647);
nor U4774 (N_4774,N_4718,N_4713);
nor U4775 (N_4775,N_4610,N_4629);
nand U4776 (N_4776,N_4574,N_4671);
nand U4777 (N_4777,N_4684,N_4739);
xnor U4778 (N_4778,N_4646,N_4734);
xor U4779 (N_4779,N_4737,N_4519);
or U4780 (N_4780,N_4565,N_4518);
and U4781 (N_4781,N_4513,N_4592);
xnor U4782 (N_4782,N_4619,N_4581);
or U4783 (N_4783,N_4637,N_4668);
or U4784 (N_4784,N_4732,N_4633);
nor U4785 (N_4785,N_4680,N_4676);
nor U4786 (N_4786,N_4551,N_4615);
nand U4787 (N_4787,N_4686,N_4711);
and U4788 (N_4788,N_4667,N_4554);
or U4789 (N_4789,N_4532,N_4503);
or U4790 (N_4790,N_4501,N_4605);
nand U4791 (N_4791,N_4648,N_4677);
xor U4792 (N_4792,N_4698,N_4588);
nor U4793 (N_4793,N_4578,N_4678);
xnor U4794 (N_4794,N_4552,N_4535);
xnor U4795 (N_4795,N_4502,N_4527);
nor U4796 (N_4796,N_4658,N_4517);
nor U4797 (N_4797,N_4509,N_4721);
or U4798 (N_4798,N_4632,N_4664);
nor U4799 (N_4799,N_4617,N_4599);
nand U4800 (N_4800,N_4563,N_4566);
xor U4801 (N_4801,N_4609,N_4511);
nor U4802 (N_4802,N_4585,N_4708);
and U4803 (N_4803,N_4672,N_4735);
xor U4804 (N_4804,N_4690,N_4745);
or U4805 (N_4805,N_4720,N_4545);
nor U4806 (N_4806,N_4717,N_4507);
xor U4807 (N_4807,N_4725,N_4601);
and U4808 (N_4808,N_4742,N_4570);
or U4809 (N_4809,N_4543,N_4714);
nand U4810 (N_4810,N_4538,N_4561);
xor U4811 (N_4811,N_4723,N_4541);
xor U4812 (N_4812,N_4697,N_4653);
and U4813 (N_4813,N_4560,N_4529);
xnor U4814 (N_4814,N_4526,N_4564);
and U4815 (N_4815,N_4569,N_4525);
or U4816 (N_4816,N_4726,N_4638);
and U4817 (N_4817,N_4596,N_4696);
xnor U4818 (N_4818,N_4536,N_4608);
nand U4819 (N_4819,N_4673,N_4523);
xnor U4820 (N_4820,N_4627,N_4651);
or U4821 (N_4821,N_4624,N_4571);
or U4822 (N_4822,N_4597,N_4675);
xor U4823 (N_4823,N_4572,N_4542);
nand U4824 (N_4824,N_4524,N_4635);
nor U4825 (N_4825,N_4665,N_4649);
nor U4826 (N_4826,N_4692,N_4515);
and U4827 (N_4827,N_4681,N_4650);
xnor U4828 (N_4828,N_4600,N_4642);
nand U4829 (N_4829,N_4634,N_4631);
nand U4830 (N_4830,N_4531,N_4589);
nand U4831 (N_4831,N_4528,N_4738);
xor U4832 (N_4832,N_4741,N_4618);
nand U4833 (N_4833,N_4557,N_4598);
xor U4834 (N_4834,N_4662,N_4623);
nor U4835 (N_4835,N_4736,N_4652);
nor U4836 (N_4836,N_4533,N_4577);
or U4837 (N_4837,N_4521,N_4594);
xor U4838 (N_4838,N_4730,N_4612);
or U4839 (N_4839,N_4613,N_4576);
nor U4840 (N_4840,N_4614,N_4512);
nand U4841 (N_4841,N_4728,N_4704);
and U4842 (N_4842,N_4636,N_4558);
nand U4843 (N_4843,N_4562,N_4659);
nand U4844 (N_4844,N_4616,N_4703);
and U4845 (N_4845,N_4727,N_4705);
and U4846 (N_4846,N_4559,N_4621);
nand U4847 (N_4847,N_4657,N_4606);
or U4848 (N_4848,N_4506,N_4716);
or U4849 (N_4849,N_4591,N_4626);
or U4850 (N_4850,N_4573,N_4530);
nand U4851 (N_4851,N_4539,N_4567);
or U4852 (N_4852,N_4520,N_4625);
and U4853 (N_4853,N_4719,N_4687);
xor U4854 (N_4854,N_4611,N_4722);
nand U4855 (N_4855,N_4516,N_4504);
nand U4856 (N_4856,N_4709,N_4731);
or U4857 (N_4857,N_4514,N_4655);
and U4858 (N_4858,N_4669,N_4534);
nor U4859 (N_4859,N_4522,N_4508);
and U4860 (N_4860,N_4746,N_4666);
nor U4861 (N_4861,N_4701,N_4694);
xor U4862 (N_4862,N_4691,N_4656);
or U4863 (N_4863,N_4549,N_4583);
xnor U4864 (N_4864,N_4641,N_4510);
or U4865 (N_4865,N_4537,N_4553);
nor U4866 (N_4866,N_4740,N_4712);
nor U4867 (N_4867,N_4584,N_4640);
or U4868 (N_4868,N_4644,N_4544);
or U4869 (N_4869,N_4582,N_4547);
and U4870 (N_4870,N_4622,N_4628);
xnor U4871 (N_4871,N_4695,N_4568);
nand U4872 (N_4872,N_4550,N_4595);
and U4873 (N_4873,N_4679,N_4748);
nand U4874 (N_4874,N_4715,N_4586);
or U4875 (N_4875,N_4648,N_4632);
or U4876 (N_4876,N_4676,N_4649);
or U4877 (N_4877,N_4609,N_4620);
or U4878 (N_4878,N_4513,N_4509);
xor U4879 (N_4879,N_4746,N_4526);
nor U4880 (N_4880,N_4646,N_4578);
nor U4881 (N_4881,N_4679,N_4715);
nand U4882 (N_4882,N_4584,N_4566);
nor U4883 (N_4883,N_4607,N_4582);
or U4884 (N_4884,N_4728,N_4530);
nor U4885 (N_4885,N_4740,N_4503);
nand U4886 (N_4886,N_4526,N_4739);
nor U4887 (N_4887,N_4686,N_4588);
or U4888 (N_4888,N_4596,N_4512);
or U4889 (N_4889,N_4516,N_4500);
nor U4890 (N_4890,N_4515,N_4526);
nand U4891 (N_4891,N_4648,N_4622);
and U4892 (N_4892,N_4557,N_4735);
xor U4893 (N_4893,N_4622,N_4515);
or U4894 (N_4894,N_4737,N_4738);
nor U4895 (N_4895,N_4621,N_4576);
and U4896 (N_4896,N_4537,N_4608);
xnor U4897 (N_4897,N_4529,N_4718);
and U4898 (N_4898,N_4529,N_4538);
nor U4899 (N_4899,N_4705,N_4626);
and U4900 (N_4900,N_4542,N_4651);
nor U4901 (N_4901,N_4571,N_4589);
xnor U4902 (N_4902,N_4523,N_4712);
nand U4903 (N_4903,N_4549,N_4633);
nand U4904 (N_4904,N_4651,N_4571);
nand U4905 (N_4905,N_4699,N_4575);
or U4906 (N_4906,N_4598,N_4640);
nand U4907 (N_4907,N_4573,N_4717);
and U4908 (N_4908,N_4738,N_4515);
nand U4909 (N_4909,N_4515,N_4568);
or U4910 (N_4910,N_4734,N_4718);
xnor U4911 (N_4911,N_4523,N_4728);
or U4912 (N_4912,N_4555,N_4686);
nor U4913 (N_4913,N_4749,N_4509);
xor U4914 (N_4914,N_4649,N_4721);
or U4915 (N_4915,N_4626,N_4515);
nand U4916 (N_4916,N_4706,N_4638);
xor U4917 (N_4917,N_4699,N_4710);
and U4918 (N_4918,N_4624,N_4711);
nor U4919 (N_4919,N_4679,N_4737);
xor U4920 (N_4920,N_4672,N_4698);
nor U4921 (N_4921,N_4585,N_4566);
and U4922 (N_4922,N_4627,N_4622);
xnor U4923 (N_4923,N_4645,N_4654);
nor U4924 (N_4924,N_4567,N_4538);
or U4925 (N_4925,N_4722,N_4587);
nor U4926 (N_4926,N_4571,N_4693);
nor U4927 (N_4927,N_4679,N_4682);
nand U4928 (N_4928,N_4543,N_4747);
and U4929 (N_4929,N_4576,N_4699);
or U4930 (N_4930,N_4674,N_4706);
nor U4931 (N_4931,N_4749,N_4520);
or U4932 (N_4932,N_4538,N_4703);
nor U4933 (N_4933,N_4506,N_4722);
nand U4934 (N_4934,N_4605,N_4510);
nand U4935 (N_4935,N_4529,N_4540);
and U4936 (N_4936,N_4528,N_4675);
xnor U4937 (N_4937,N_4549,N_4642);
and U4938 (N_4938,N_4541,N_4593);
nand U4939 (N_4939,N_4654,N_4517);
xor U4940 (N_4940,N_4615,N_4629);
xnor U4941 (N_4941,N_4547,N_4721);
xor U4942 (N_4942,N_4727,N_4534);
and U4943 (N_4943,N_4632,N_4671);
and U4944 (N_4944,N_4621,N_4517);
xor U4945 (N_4945,N_4710,N_4646);
nand U4946 (N_4946,N_4671,N_4643);
nor U4947 (N_4947,N_4609,N_4722);
nor U4948 (N_4948,N_4749,N_4724);
nor U4949 (N_4949,N_4603,N_4508);
xor U4950 (N_4950,N_4575,N_4530);
or U4951 (N_4951,N_4555,N_4586);
and U4952 (N_4952,N_4538,N_4722);
nor U4953 (N_4953,N_4669,N_4542);
and U4954 (N_4954,N_4522,N_4616);
or U4955 (N_4955,N_4578,N_4618);
or U4956 (N_4956,N_4702,N_4584);
or U4957 (N_4957,N_4657,N_4565);
and U4958 (N_4958,N_4614,N_4576);
nand U4959 (N_4959,N_4590,N_4711);
nor U4960 (N_4960,N_4743,N_4513);
xnor U4961 (N_4961,N_4565,N_4670);
xor U4962 (N_4962,N_4720,N_4647);
and U4963 (N_4963,N_4698,N_4718);
or U4964 (N_4964,N_4665,N_4617);
nor U4965 (N_4965,N_4677,N_4558);
and U4966 (N_4966,N_4606,N_4504);
xor U4967 (N_4967,N_4726,N_4690);
xnor U4968 (N_4968,N_4636,N_4749);
or U4969 (N_4969,N_4539,N_4613);
and U4970 (N_4970,N_4581,N_4501);
nor U4971 (N_4971,N_4674,N_4572);
xnor U4972 (N_4972,N_4608,N_4566);
or U4973 (N_4973,N_4699,N_4640);
and U4974 (N_4974,N_4639,N_4708);
nand U4975 (N_4975,N_4635,N_4592);
xor U4976 (N_4976,N_4526,N_4548);
nand U4977 (N_4977,N_4582,N_4548);
or U4978 (N_4978,N_4646,N_4523);
xnor U4979 (N_4979,N_4623,N_4609);
or U4980 (N_4980,N_4639,N_4655);
nor U4981 (N_4981,N_4655,N_4694);
xnor U4982 (N_4982,N_4622,N_4581);
nor U4983 (N_4983,N_4521,N_4647);
and U4984 (N_4984,N_4639,N_4515);
nor U4985 (N_4985,N_4551,N_4743);
xnor U4986 (N_4986,N_4619,N_4698);
xnor U4987 (N_4987,N_4508,N_4696);
xor U4988 (N_4988,N_4511,N_4613);
or U4989 (N_4989,N_4686,N_4717);
nor U4990 (N_4990,N_4518,N_4719);
xor U4991 (N_4991,N_4544,N_4558);
or U4992 (N_4992,N_4549,N_4579);
or U4993 (N_4993,N_4630,N_4520);
xnor U4994 (N_4994,N_4600,N_4611);
nor U4995 (N_4995,N_4513,N_4608);
nand U4996 (N_4996,N_4529,N_4661);
nor U4997 (N_4997,N_4690,N_4584);
nor U4998 (N_4998,N_4623,N_4550);
nor U4999 (N_4999,N_4696,N_4643);
or U5000 (N_5000,N_4889,N_4757);
xor U5001 (N_5001,N_4840,N_4756);
or U5002 (N_5002,N_4919,N_4763);
and U5003 (N_5003,N_4807,N_4761);
nand U5004 (N_5004,N_4862,N_4943);
nand U5005 (N_5005,N_4881,N_4957);
or U5006 (N_5006,N_4900,N_4989);
nand U5007 (N_5007,N_4818,N_4879);
nand U5008 (N_5008,N_4959,N_4805);
or U5009 (N_5009,N_4876,N_4750);
or U5010 (N_5010,N_4833,N_4874);
nand U5011 (N_5011,N_4983,N_4988);
and U5012 (N_5012,N_4754,N_4854);
and U5013 (N_5013,N_4952,N_4872);
and U5014 (N_5014,N_4991,N_4997);
nor U5015 (N_5015,N_4917,N_4838);
nand U5016 (N_5016,N_4877,N_4963);
nand U5017 (N_5017,N_4961,N_4871);
xor U5018 (N_5018,N_4998,N_4973);
nor U5019 (N_5019,N_4985,N_4899);
nand U5020 (N_5020,N_4849,N_4767);
nand U5021 (N_5021,N_4846,N_4867);
nand U5022 (N_5022,N_4822,N_4759);
xor U5023 (N_5023,N_4792,N_4853);
and U5024 (N_5024,N_4918,N_4855);
nand U5025 (N_5025,N_4824,N_4935);
xor U5026 (N_5026,N_4994,N_4987);
and U5027 (N_5027,N_4844,N_4930);
and U5028 (N_5028,N_4773,N_4888);
and U5029 (N_5029,N_4884,N_4825);
nor U5030 (N_5030,N_4982,N_4808);
nand U5031 (N_5031,N_4778,N_4771);
and U5032 (N_5032,N_4770,N_4954);
nor U5033 (N_5033,N_4772,N_4895);
nor U5034 (N_5034,N_4951,N_4751);
nor U5035 (N_5035,N_4910,N_4978);
nor U5036 (N_5036,N_4891,N_4921);
or U5037 (N_5037,N_4835,N_4933);
xnor U5038 (N_5038,N_4827,N_4828);
and U5039 (N_5039,N_4892,N_4839);
or U5040 (N_5040,N_4836,N_4782);
nand U5041 (N_5041,N_4793,N_4992);
nand U5042 (N_5042,N_4896,N_4811);
nor U5043 (N_5043,N_4866,N_4944);
xor U5044 (N_5044,N_4789,N_4799);
and U5045 (N_5045,N_4995,N_4848);
or U5046 (N_5046,N_4863,N_4801);
nand U5047 (N_5047,N_4769,N_4931);
and U5048 (N_5048,N_4832,N_4803);
nor U5049 (N_5049,N_4834,N_4893);
and U5050 (N_5050,N_4785,N_4981);
and U5051 (N_5051,N_4858,N_4870);
xor U5052 (N_5052,N_4783,N_4764);
nand U5053 (N_5053,N_4967,N_4928);
or U5054 (N_5054,N_4837,N_4906);
nor U5055 (N_5055,N_4986,N_4962);
nand U5056 (N_5056,N_4907,N_4851);
and U5057 (N_5057,N_4925,N_4913);
xnor U5058 (N_5058,N_4950,N_4760);
nand U5059 (N_5059,N_4817,N_4816);
or U5060 (N_5060,N_4923,N_4868);
or U5061 (N_5061,N_4775,N_4904);
xor U5062 (N_5062,N_4777,N_4860);
or U5063 (N_5063,N_4940,N_4886);
or U5064 (N_5064,N_4797,N_4971);
or U5065 (N_5065,N_4937,N_4946);
or U5066 (N_5066,N_4765,N_4762);
or U5067 (N_5067,N_4847,N_4780);
nor U5068 (N_5068,N_4831,N_4829);
xor U5069 (N_5069,N_4806,N_4953);
nor U5070 (N_5070,N_4955,N_4947);
or U5071 (N_5071,N_4794,N_4972);
nor U5072 (N_5072,N_4830,N_4880);
and U5073 (N_5073,N_4905,N_4968);
xor U5074 (N_5074,N_4878,N_4914);
xnor U5075 (N_5075,N_4915,N_4796);
or U5076 (N_5076,N_4788,N_4993);
nor U5077 (N_5077,N_4970,N_4768);
nor U5078 (N_5078,N_4800,N_4890);
xor U5079 (N_5079,N_4857,N_4755);
or U5080 (N_5080,N_4934,N_4938);
and U5081 (N_5081,N_4976,N_4814);
nor U5082 (N_5082,N_4980,N_4786);
nand U5083 (N_5083,N_4927,N_4936);
and U5084 (N_5084,N_4826,N_4873);
xor U5085 (N_5085,N_4926,N_4861);
and U5086 (N_5086,N_4865,N_4843);
and U5087 (N_5087,N_4798,N_4969);
xor U5088 (N_5088,N_4795,N_4804);
nor U5089 (N_5089,N_4903,N_4902);
and U5090 (N_5090,N_4945,N_4956);
xnor U5091 (N_5091,N_4932,N_4856);
nand U5092 (N_5092,N_4965,N_4887);
xnor U5093 (N_5093,N_4820,N_4990);
nand U5094 (N_5094,N_4841,N_4999);
and U5095 (N_5095,N_4875,N_4920);
nand U5096 (N_5096,N_4964,N_4779);
and U5097 (N_5097,N_4885,N_4821);
nor U5098 (N_5098,N_4996,N_4901);
and U5099 (N_5099,N_4984,N_4960);
and U5100 (N_5100,N_4758,N_4802);
and U5101 (N_5101,N_4897,N_4894);
nor U5102 (N_5102,N_4974,N_4784);
and U5103 (N_5103,N_4883,N_4823);
or U5104 (N_5104,N_4909,N_4809);
or U5105 (N_5105,N_4939,N_4924);
xor U5106 (N_5106,N_4958,N_4941);
or U5107 (N_5107,N_4977,N_4776);
or U5108 (N_5108,N_4752,N_4864);
nor U5109 (N_5109,N_4813,N_4898);
xnor U5110 (N_5110,N_4753,N_4787);
xnor U5111 (N_5111,N_4791,N_4774);
and U5112 (N_5112,N_4852,N_4766);
xor U5113 (N_5113,N_4916,N_4949);
nand U5114 (N_5114,N_4869,N_4790);
xnor U5115 (N_5115,N_4912,N_4911);
nor U5116 (N_5116,N_4845,N_4819);
or U5117 (N_5117,N_4850,N_4882);
nor U5118 (N_5118,N_4812,N_4929);
and U5119 (N_5119,N_4948,N_4975);
or U5120 (N_5120,N_4815,N_4842);
nand U5121 (N_5121,N_4979,N_4922);
nor U5122 (N_5122,N_4781,N_4908);
or U5123 (N_5123,N_4942,N_4859);
nand U5124 (N_5124,N_4966,N_4810);
nand U5125 (N_5125,N_4789,N_4917);
nor U5126 (N_5126,N_4833,N_4753);
nand U5127 (N_5127,N_4829,N_4842);
and U5128 (N_5128,N_4776,N_4997);
or U5129 (N_5129,N_4773,N_4862);
nor U5130 (N_5130,N_4755,N_4875);
nand U5131 (N_5131,N_4758,N_4861);
xor U5132 (N_5132,N_4906,N_4989);
nor U5133 (N_5133,N_4941,N_4954);
and U5134 (N_5134,N_4822,N_4818);
and U5135 (N_5135,N_4867,N_4961);
nand U5136 (N_5136,N_4801,N_4823);
nor U5137 (N_5137,N_4799,N_4982);
or U5138 (N_5138,N_4831,N_4845);
or U5139 (N_5139,N_4963,N_4828);
and U5140 (N_5140,N_4940,N_4961);
nand U5141 (N_5141,N_4778,N_4886);
xor U5142 (N_5142,N_4927,N_4876);
nand U5143 (N_5143,N_4996,N_4919);
nand U5144 (N_5144,N_4942,N_4770);
or U5145 (N_5145,N_4933,N_4808);
or U5146 (N_5146,N_4829,N_4930);
and U5147 (N_5147,N_4973,N_4791);
xnor U5148 (N_5148,N_4910,N_4827);
nand U5149 (N_5149,N_4772,N_4927);
xnor U5150 (N_5150,N_4756,N_4772);
and U5151 (N_5151,N_4987,N_4864);
nor U5152 (N_5152,N_4823,N_4968);
or U5153 (N_5153,N_4803,N_4973);
xor U5154 (N_5154,N_4934,N_4777);
nor U5155 (N_5155,N_4905,N_4754);
nand U5156 (N_5156,N_4820,N_4962);
or U5157 (N_5157,N_4908,N_4950);
xor U5158 (N_5158,N_4755,N_4761);
nand U5159 (N_5159,N_4797,N_4860);
nand U5160 (N_5160,N_4955,N_4879);
nand U5161 (N_5161,N_4887,N_4898);
and U5162 (N_5162,N_4914,N_4924);
and U5163 (N_5163,N_4809,N_4854);
nand U5164 (N_5164,N_4995,N_4974);
nand U5165 (N_5165,N_4818,N_4906);
nand U5166 (N_5166,N_4947,N_4800);
nand U5167 (N_5167,N_4892,N_4773);
or U5168 (N_5168,N_4877,N_4884);
and U5169 (N_5169,N_4943,N_4863);
or U5170 (N_5170,N_4995,N_4868);
nand U5171 (N_5171,N_4916,N_4914);
or U5172 (N_5172,N_4833,N_4900);
or U5173 (N_5173,N_4814,N_4865);
nand U5174 (N_5174,N_4858,N_4881);
nand U5175 (N_5175,N_4971,N_4902);
nand U5176 (N_5176,N_4772,N_4812);
or U5177 (N_5177,N_4796,N_4847);
xnor U5178 (N_5178,N_4899,N_4969);
or U5179 (N_5179,N_4891,N_4903);
and U5180 (N_5180,N_4874,N_4774);
nand U5181 (N_5181,N_4880,N_4961);
or U5182 (N_5182,N_4931,N_4870);
xnor U5183 (N_5183,N_4792,N_4764);
or U5184 (N_5184,N_4873,N_4908);
xor U5185 (N_5185,N_4876,N_4766);
or U5186 (N_5186,N_4960,N_4793);
and U5187 (N_5187,N_4851,N_4884);
nor U5188 (N_5188,N_4803,N_4996);
or U5189 (N_5189,N_4812,N_4932);
xor U5190 (N_5190,N_4770,N_4927);
xnor U5191 (N_5191,N_4842,N_4773);
nor U5192 (N_5192,N_4941,N_4797);
nand U5193 (N_5193,N_4809,N_4837);
xnor U5194 (N_5194,N_4853,N_4786);
nand U5195 (N_5195,N_4824,N_4838);
nand U5196 (N_5196,N_4761,N_4871);
nor U5197 (N_5197,N_4822,N_4779);
and U5198 (N_5198,N_4785,N_4984);
xor U5199 (N_5199,N_4917,N_4776);
or U5200 (N_5200,N_4865,N_4953);
or U5201 (N_5201,N_4923,N_4925);
or U5202 (N_5202,N_4752,N_4917);
and U5203 (N_5203,N_4843,N_4756);
or U5204 (N_5204,N_4780,N_4925);
or U5205 (N_5205,N_4824,N_4885);
and U5206 (N_5206,N_4984,N_4963);
and U5207 (N_5207,N_4896,N_4838);
nor U5208 (N_5208,N_4807,N_4942);
xor U5209 (N_5209,N_4905,N_4801);
and U5210 (N_5210,N_4878,N_4803);
nand U5211 (N_5211,N_4948,N_4843);
and U5212 (N_5212,N_4878,N_4825);
xor U5213 (N_5213,N_4994,N_4818);
and U5214 (N_5214,N_4830,N_4981);
nor U5215 (N_5215,N_4985,N_4890);
and U5216 (N_5216,N_4763,N_4872);
and U5217 (N_5217,N_4879,N_4904);
or U5218 (N_5218,N_4904,N_4816);
or U5219 (N_5219,N_4796,N_4835);
nand U5220 (N_5220,N_4958,N_4808);
or U5221 (N_5221,N_4917,N_4844);
or U5222 (N_5222,N_4895,N_4996);
xnor U5223 (N_5223,N_4949,N_4945);
or U5224 (N_5224,N_4798,N_4982);
nor U5225 (N_5225,N_4835,N_4829);
xor U5226 (N_5226,N_4868,N_4976);
xnor U5227 (N_5227,N_4831,N_4850);
or U5228 (N_5228,N_4937,N_4823);
nor U5229 (N_5229,N_4960,N_4921);
and U5230 (N_5230,N_4817,N_4978);
nand U5231 (N_5231,N_4837,N_4882);
xor U5232 (N_5232,N_4790,N_4793);
and U5233 (N_5233,N_4751,N_4886);
xnor U5234 (N_5234,N_4905,N_4872);
or U5235 (N_5235,N_4952,N_4835);
nor U5236 (N_5236,N_4832,N_4926);
or U5237 (N_5237,N_4807,N_4991);
and U5238 (N_5238,N_4799,N_4808);
and U5239 (N_5239,N_4983,N_4760);
xnor U5240 (N_5240,N_4937,N_4985);
nor U5241 (N_5241,N_4975,N_4937);
nand U5242 (N_5242,N_4820,N_4771);
or U5243 (N_5243,N_4849,N_4838);
and U5244 (N_5244,N_4896,N_4927);
and U5245 (N_5245,N_4846,N_4833);
xor U5246 (N_5246,N_4947,N_4824);
nor U5247 (N_5247,N_4881,N_4959);
nor U5248 (N_5248,N_4989,N_4876);
or U5249 (N_5249,N_4914,N_4873);
nor U5250 (N_5250,N_5078,N_5177);
and U5251 (N_5251,N_5108,N_5170);
nand U5252 (N_5252,N_5071,N_5091);
nor U5253 (N_5253,N_5193,N_5190);
or U5254 (N_5254,N_5129,N_5068);
or U5255 (N_5255,N_5223,N_5070);
and U5256 (N_5256,N_5030,N_5124);
xor U5257 (N_5257,N_5013,N_5132);
nor U5258 (N_5258,N_5086,N_5183);
nand U5259 (N_5259,N_5230,N_5060);
xnor U5260 (N_5260,N_5225,N_5148);
and U5261 (N_5261,N_5189,N_5167);
nand U5262 (N_5262,N_5113,N_5044);
xnor U5263 (N_5263,N_5202,N_5231);
nor U5264 (N_5264,N_5110,N_5056);
nor U5265 (N_5265,N_5150,N_5112);
nor U5266 (N_5266,N_5248,N_5180);
xnor U5267 (N_5267,N_5215,N_5235);
or U5268 (N_5268,N_5119,N_5239);
nand U5269 (N_5269,N_5023,N_5053);
nand U5270 (N_5270,N_5050,N_5125);
xor U5271 (N_5271,N_5214,N_5169);
and U5272 (N_5272,N_5038,N_5222);
and U5273 (N_5273,N_5079,N_5227);
and U5274 (N_5274,N_5122,N_5047);
nand U5275 (N_5275,N_5057,N_5074);
nand U5276 (N_5276,N_5166,N_5090);
nor U5277 (N_5277,N_5022,N_5042);
or U5278 (N_5278,N_5096,N_5158);
and U5279 (N_5279,N_5121,N_5012);
xnor U5280 (N_5280,N_5191,N_5218);
nand U5281 (N_5281,N_5186,N_5024);
xnor U5282 (N_5282,N_5233,N_5116);
nor U5283 (N_5283,N_5049,N_5104);
xnor U5284 (N_5284,N_5137,N_5051);
xor U5285 (N_5285,N_5246,N_5175);
or U5286 (N_5286,N_5066,N_5199);
and U5287 (N_5287,N_5092,N_5004);
nand U5288 (N_5288,N_5000,N_5134);
and U5289 (N_5289,N_5195,N_5018);
or U5290 (N_5290,N_5021,N_5102);
xnor U5291 (N_5291,N_5232,N_5153);
xor U5292 (N_5292,N_5217,N_5123);
or U5293 (N_5293,N_5156,N_5001);
and U5294 (N_5294,N_5184,N_5015);
nor U5295 (N_5295,N_5093,N_5131);
xor U5296 (N_5296,N_5085,N_5016);
nor U5297 (N_5297,N_5160,N_5052);
nand U5298 (N_5298,N_5025,N_5087);
xnor U5299 (N_5299,N_5036,N_5236);
nor U5300 (N_5300,N_5145,N_5094);
nor U5301 (N_5301,N_5157,N_5194);
nor U5302 (N_5302,N_5243,N_5172);
xnor U5303 (N_5303,N_5142,N_5206);
xor U5304 (N_5304,N_5221,N_5063);
xor U5305 (N_5305,N_5029,N_5247);
nor U5306 (N_5306,N_5084,N_5076);
and U5307 (N_5307,N_5234,N_5045);
or U5308 (N_5308,N_5212,N_5118);
nand U5309 (N_5309,N_5146,N_5220);
and U5310 (N_5310,N_5139,N_5111);
xnor U5311 (N_5311,N_5115,N_5017);
or U5312 (N_5312,N_5127,N_5174);
nand U5313 (N_5313,N_5228,N_5097);
or U5314 (N_5314,N_5171,N_5155);
nor U5315 (N_5315,N_5041,N_5002);
nor U5316 (N_5316,N_5198,N_5046);
and U5317 (N_5317,N_5072,N_5006);
nor U5318 (N_5318,N_5126,N_5027);
nor U5319 (N_5319,N_5120,N_5229);
or U5320 (N_5320,N_5031,N_5009);
nor U5321 (N_5321,N_5178,N_5182);
nand U5322 (N_5322,N_5179,N_5192);
nor U5323 (N_5323,N_5138,N_5208);
nand U5324 (N_5324,N_5117,N_5007);
nor U5325 (N_5325,N_5241,N_5034);
or U5326 (N_5326,N_5224,N_5210);
and U5327 (N_5327,N_5082,N_5065);
nand U5328 (N_5328,N_5154,N_5054);
or U5329 (N_5329,N_5032,N_5205);
and U5330 (N_5330,N_5095,N_5187);
nand U5331 (N_5331,N_5083,N_5033);
nand U5332 (N_5332,N_5249,N_5037);
nand U5333 (N_5333,N_5061,N_5073);
nand U5334 (N_5334,N_5008,N_5176);
xnor U5335 (N_5335,N_5014,N_5081);
xor U5336 (N_5336,N_5005,N_5055);
xnor U5337 (N_5337,N_5003,N_5238);
and U5338 (N_5338,N_5028,N_5162);
nor U5339 (N_5339,N_5040,N_5106);
nor U5340 (N_5340,N_5088,N_5020);
nand U5341 (N_5341,N_5140,N_5089);
nor U5342 (N_5342,N_5062,N_5011);
nor U5343 (N_5343,N_5147,N_5219);
nand U5344 (N_5344,N_5144,N_5101);
nor U5345 (N_5345,N_5105,N_5188);
or U5346 (N_5346,N_5237,N_5135);
or U5347 (N_5347,N_5075,N_5173);
and U5348 (N_5348,N_5240,N_5098);
or U5349 (N_5349,N_5185,N_5161);
nor U5350 (N_5350,N_5245,N_5204);
xor U5351 (N_5351,N_5039,N_5059);
xnor U5352 (N_5352,N_5067,N_5143);
nand U5353 (N_5353,N_5181,N_5130);
or U5354 (N_5354,N_5058,N_5149);
xnor U5355 (N_5355,N_5010,N_5026);
or U5356 (N_5356,N_5168,N_5209);
xnor U5357 (N_5357,N_5035,N_5080);
and U5358 (N_5358,N_5216,N_5207);
xnor U5359 (N_5359,N_5200,N_5099);
or U5360 (N_5360,N_5114,N_5165);
nor U5361 (N_5361,N_5109,N_5048);
nand U5362 (N_5362,N_5043,N_5201);
xnor U5363 (N_5363,N_5164,N_5128);
nand U5364 (N_5364,N_5163,N_5069);
or U5365 (N_5365,N_5244,N_5197);
and U5366 (N_5366,N_5213,N_5019);
nand U5367 (N_5367,N_5103,N_5141);
and U5368 (N_5368,N_5159,N_5107);
nand U5369 (N_5369,N_5196,N_5077);
nor U5370 (N_5370,N_5100,N_5136);
xor U5371 (N_5371,N_5064,N_5133);
or U5372 (N_5372,N_5152,N_5211);
nand U5373 (N_5373,N_5151,N_5203);
xnor U5374 (N_5374,N_5242,N_5226);
nor U5375 (N_5375,N_5200,N_5177);
nand U5376 (N_5376,N_5234,N_5018);
xnor U5377 (N_5377,N_5132,N_5039);
and U5378 (N_5378,N_5171,N_5152);
or U5379 (N_5379,N_5166,N_5031);
xor U5380 (N_5380,N_5168,N_5038);
xnor U5381 (N_5381,N_5072,N_5073);
and U5382 (N_5382,N_5219,N_5047);
or U5383 (N_5383,N_5192,N_5232);
nand U5384 (N_5384,N_5012,N_5230);
or U5385 (N_5385,N_5006,N_5166);
nor U5386 (N_5386,N_5120,N_5145);
nor U5387 (N_5387,N_5083,N_5005);
and U5388 (N_5388,N_5147,N_5211);
nor U5389 (N_5389,N_5201,N_5247);
nand U5390 (N_5390,N_5077,N_5192);
or U5391 (N_5391,N_5088,N_5187);
and U5392 (N_5392,N_5111,N_5231);
and U5393 (N_5393,N_5240,N_5108);
nand U5394 (N_5394,N_5229,N_5160);
and U5395 (N_5395,N_5203,N_5178);
xor U5396 (N_5396,N_5005,N_5039);
and U5397 (N_5397,N_5083,N_5088);
xor U5398 (N_5398,N_5070,N_5170);
nor U5399 (N_5399,N_5069,N_5037);
and U5400 (N_5400,N_5042,N_5152);
or U5401 (N_5401,N_5099,N_5146);
or U5402 (N_5402,N_5162,N_5174);
or U5403 (N_5403,N_5190,N_5239);
and U5404 (N_5404,N_5144,N_5049);
nor U5405 (N_5405,N_5206,N_5246);
nand U5406 (N_5406,N_5141,N_5161);
or U5407 (N_5407,N_5180,N_5102);
nand U5408 (N_5408,N_5218,N_5000);
or U5409 (N_5409,N_5054,N_5206);
and U5410 (N_5410,N_5197,N_5039);
xnor U5411 (N_5411,N_5075,N_5020);
and U5412 (N_5412,N_5217,N_5108);
or U5413 (N_5413,N_5223,N_5063);
xnor U5414 (N_5414,N_5041,N_5134);
or U5415 (N_5415,N_5082,N_5145);
nand U5416 (N_5416,N_5205,N_5104);
nand U5417 (N_5417,N_5064,N_5173);
nor U5418 (N_5418,N_5090,N_5005);
xor U5419 (N_5419,N_5005,N_5129);
or U5420 (N_5420,N_5209,N_5009);
xor U5421 (N_5421,N_5016,N_5206);
xor U5422 (N_5422,N_5004,N_5098);
nand U5423 (N_5423,N_5036,N_5209);
nor U5424 (N_5424,N_5157,N_5196);
nor U5425 (N_5425,N_5009,N_5029);
and U5426 (N_5426,N_5123,N_5247);
xor U5427 (N_5427,N_5065,N_5078);
or U5428 (N_5428,N_5035,N_5124);
or U5429 (N_5429,N_5248,N_5124);
nand U5430 (N_5430,N_5233,N_5226);
or U5431 (N_5431,N_5004,N_5075);
or U5432 (N_5432,N_5239,N_5071);
and U5433 (N_5433,N_5171,N_5187);
nand U5434 (N_5434,N_5057,N_5175);
and U5435 (N_5435,N_5046,N_5197);
and U5436 (N_5436,N_5141,N_5239);
or U5437 (N_5437,N_5153,N_5233);
nand U5438 (N_5438,N_5170,N_5232);
xor U5439 (N_5439,N_5095,N_5210);
xnor U5440 (N_5440,N_5079,N_5177);
xnor U5441 (N_5441,N_5087,N_5148);
and U5442 (N_5442,N_5170,N_5157);
xor U5443 (N_5443,N_5224,N_5103);
nand U5444 (N_5444,N_5023,N_5098);
and U5445 (N_5445,N_5157,N_5068);
or U5446 (N_5446,N_5137,N_5083);
nand U5447 (N_5447,N_5012,N_5005);
nor U5448 (N_5448,N_5176,N_5109);
and U5449 (N_5449,N_5186,N_5100);
and U5450 (N_5450,N_5249,N_5230);
xnor U5451 (N_5451,N_5148,N_5025);
xnor U5452 (N_5452,N_5186,N_5011);
nand U5453 (N_5453,N_5153,N_5127);
nand U5454 (N_5454,N_5065,N_5249);
nor U5455 (N_5455,N_5118,N_5130);
xnor U5456 (N_5456,N_5095,N_5216);
and U5457 (N_5457,N_5088,N_5081);
and U5458 (N_5458,N_5063,N_5210);
and U5459 (N_5459,N_5127,N_5232);
nor U5460 (N_5460,N_5233,N_5234);
xnor U5461 (N_5461,N_5244,N_5247);
nand U5462 (N_5462,N_5214,N_5235);
or U5463 (N_5463,N_5217,N_5063);
or U5464 (N_5464,N_5166,N_5059);
nand U5465 (N_5465,N_5235,N_5144);
xor U5466 (N_5466,N_5075,N_5198);
or U5467 (N_5467,N_5037,N_5108);
or U5468 (N_5468,N_5233,N_5214);
and U5469 (N_5469,N_5122,N_5147);
nand U5470 (N_5470,N_5068,N_5008);
and U5471 (N_5471,N_5191,N_5024);
or U5472 (N_5472,N_5012,N_5175);
nor U5473 (N_5473,N_5032,N_5012);
xor U5474 (N_5474,N_5224,N_5050);
xor U5475 (N_5475,N_5009,N_5068);
xor U5476 (N_5476,N_5124,N_5119);
xnor U5477 (N_5477,N_5085,N_5183);
xnor U5478 (N_5478,N_5005,N_5028);
xnor U5479 (N_5479,N_5058,N_5089);
and U5480 (N_5480,N_5146,N_5232);
or U5481 (N_5481,N_5080,N_5169);
and U5482 (N_5482,N_5219,N_5096);
or U5483 (N_5483,N_5102,N_5026);
nor U5484 (N_5484,N_5020,N_5033);
or U5485 (N_5485,N_5134,N_5107);
nand U5486 (N_5486,N_5136,N_5067);
and U5487 (N_5487,N_5224,N_5186);
xor U5488 (N_5488,N_5211,N_5171);
or U5489 (N_5489,N_5088,N_5203);
nor U5490 (N_5490,N_5234,N_5054);
nand U5491 (N_5491,N_5142,N_5119);
or U5492 (N_5492,N_5197,N_5037);
and U5493 (N_5493,N_5018,N_5039);
nand U5494 (N_5494,N_5040,N_5084);
or U5495 (N_5495,N_5115,N_5049);
or U5496 (N_5496,N_5111,N_5103);
xnor U5497 (N_5497,N_5224,N_5174);
nor U5498 (N_5498,N_5078,N_5224);
xor U5499 (N_5499,N_5114,N_5237);
nor U5500 (N_5500,N_5275,N_5279);
or U5501 (N_5501,N_5254,N_5396);
or U5502 (N_5502,N_5337,N_5259);
nor U5503 (N_5503,N_5319,N_5305);
nand U5504 (N_5504,N_5497,N_5310);
and U5505 (N_5505,N_5386,N_5339);
nor U5506 (N_5506,N_5426,N_5495);
and U5507 (N_5507,N_5300,N_5354);
or U5508 (N_5508,N_5288,N_5493);
xor U5509 (N_5509,N_5312,N_5353);
nand U5510 (N_5510,N_5447,N_5309);
and U5511 (N_5511,N_5324,N_5410);
or U5512 (N_5512,N_5494,N_5462);
or U5513 (N_5513,N_5315,N_5482);
xnor U5514 (N_5514,N_5468,N_5280);
nand U5515 (N_5515,N_5367,N_5424);
and U5516 (N_5516,N_5393,N_5477);
nand U5517 (N_5517,N_5350,N_5451);
and U5518 (N_5518,N_5401,N_5377);
or U5519 (N_5519,N_5290,N_5457);
xor U5520 (N_5520,N_5433,N_5306);
nand U5521 (N_5521,N_5258,N_5438);
or U5522 (N_5522,N_5422,N_5327);
nand U5523 (N_5523,N_5371,N_5281);
xnor U5524 (N_5524,N_5478,N_5403);
nor U5525 (N_5525,N_5454,N_5325);
xor U5526 (N_5526,N_5277,N_5360);
nor U5527 (N_5527,N_5363,N_5434);
nand U5528 (N_5528,N_5471,N_5348);
and U5529 (N_5529,N_5296,N_5423);
xnor U5530 (N_5530,N_5498,N_5404);
and U5531 (N_5531,N_5358,N_5256);
nor U5532 (N_5532,N_5336,N_5452);
nor U5533 (N_5533,N_5450,N_5342);
nor U5534 (N_5534,N_5407,N_5481);
or U5535 (N_5535,N_5460,N_5449);
and U5536 (N_5536,N_5344,N_5318);
or U5537 (N_5537,N_5408,N_5340);
and U5538 (N_5538,N_5472,N_5464);
or U5539 (N_5539,N_5267,N_5427);
nor U5540 (N_5540,N_5429,N_5417);
xnor U5541 (N_5541,N_5459,N_5330);
nand U5542 (N_5542,N_5383,N_5307);
xnor U5543 (N_5543,N_5262,N_5268);
xor U5544 (N_5544,N_5485,N_5334);
and U5545 (N_5545,N_5323,N_5376);
xnor U5546 (N_5546,N_5356,N_5320);
and U5547 (N_5547,N_5291,N_5373);
xor U5548 (N_5548,N_5313,N_5278);
or U5549 (N_5549,N_5338,N_5402);
xnor U5550 (N_5550,N_5366,N_5390);
xnor U5551 (N_5551,N_5251,N_5499);
xnor U5552 (N_5552,N_5436,N_5444);
xor U5553 (N_5553,N_5435,N_5297);
nand U5554 (N_5554,N_5362,N_5431);
nor U5555 (N_5555,N_5412,N_5441);
or U5556 (N_5556,N_5321,N_5394);
or U5557 (N_5557,N_5368,N_5491);
or U5558 (N_5558,N_5492,N_5475);
nand U5559 (N_5559,N_5474,N_5385);
xnor U5560 (N_5560,N_5289,N_5314);
nor U5561 (N_5561,N_5341,N_5374);
or U5562 (N_5562,N_5298,N_5398);
xor U5563 (N_5563,N_5440,N_5382);
and U5564 (N_5564,N_5399,N_5286);
nand U5565 (N_5565,N_5442,N_5389);
nor U5566 (N_5566,N_5272,N_5253);
xnor U5567 (N_5567,N_5489,N_5260);
xor U5568 (N_5568,N_5445,N_5295);
or U5569 (N_5569,N_5261,N_5328);
and U5570 (N_5570,N_5479,N_5448);
nand U5571 (N_5571,N_5416,N_5483);
nand U5572 (N_5572,N_5317,N_5443);
xnor U5573 (N_5573,N_5496,N_5488);
xor U5574 (N_5574,N_5409,N_5357);
or U5575 (N_5575,N_5364,N_5486);
xnor U5576 (N_5576,N_5331,N_5484);
and U5577 (N_5577,N_5400,N_5273);
nand U5578 (N_5578,N_5301,N_5351);
and U5579 (N_5579,N_5250,N_5395);
nand U5580 (N_5580,N_5255,N_5276);
nor U5581 (N_5581,N_5284,N_5470);
xor U5582 (N_5582,N_5487,N_5421);
nor U5583 (N_5583,N_5473,N_5269);
nor U5584 (N_5584,N_5264,N_5302);
or U5585 (N_5585,N_5391,N_5332);
nand U5586 (N_5586,N_5308,N_5425);
nand U5587 (N_5587,N_5480,N_5359);
or U5588 (N_5588,N_5405,N_5432);
and U5589 (N_5589,N_5304,N_5428);
nor U5590 (N_5590,N_5456,N_5490);
and U5591 (N_5591,N_5420,N_5387);
nor U5592 (N_5592,N_5397,N_5257);
nand U5593 (N_5593,N_5369,N_5384);
nor U5594 (N_5594,N_5379,N_5372);
and U5595 (N_5595,N_5437,N_5287);
nand U5596 (N_5596,N_5476,N_5316);
nor U5597 (N_5597,N_5292,N_5329);
and U5598 (N_5598,N_5365,N_5430);
xnor U5599 (N_5599,N_5346,N_5263);
xor U5600 (N_5600,N_5455,N_5411);
and U5601 (N_5601,N_5271,N_5461);
nand U5602 (N_5602,N_5355,N_5465);
nand U5603 (N_5603,N_5375,N_5333);
xor U5604 (N_5604,N_5406,N_5446);
or U5605 (N_5605,N_5335,N_5311);
or U5606 (N_5606,N_5293,N_5352);
nor U5607 (N_5607,N_5299,N_5467);
and U5608 (N_5608,N_5345,N_5294);
nor U5609 (N_5609,N_5326,N_5285);
and U5610 (N_5610,N_5361,N_5347);
xor U5611 (N_5611,N_5414,N_5270);
nor U5612 (N_5612,N_5439,N_5392);
xor U5613 (N_5613,N_5458,N_5282);
or U5614 (N_5614,N_5418,N_5303);
nor U5615 (N_5615,N_5388,N_5415);
nand U5616 (N_5616,N_5419,N_5370);
nand U5617 (N_5617,N_5252,N_5378);
and U5618 (N_5618,N_5274,N_5469);
xor U5619 (N_5619,N_5343,N_5463);
and U5620 (N_5620,N_5265,N_5413);
or U5621 (N_5621,N_5380,N_5322);
or U5622 (N_5622,N_5349,N_5283);
xor U5623 (N_5623,N_5453,N_5266);
nand U5624 (N_5624,N_5466,N_5381);
and U5625 (N_5625,N_5426,N_5283);
or U5626 (N_5626,N_5327,N_5485);
or U5627 (N_5627,N_5453,N_5495);
or U5628 (N_5628,N_5368,N_5363);
nor U5629 (N_5629,N_5455,N_5452);
xnor U5630 (N_5630,N_5289,N_5285);
nor U5631 (N_5631,N_5467,N_5322);
nor U5632 (N_5632,N_5368,N_5492);
nor U5633 (N_5633,N_5370,N_5315);
nand U5634 (N_5634,N_5329,N_5387);
nand U5635 (N_5635,N_5402,N_5345);
nor U5636 (N_5636,N_5277,N_5455);
and U5637 (N_5637,N_5284,N_5391);
or U5638 (N_5638,N_5395,N_5493);
or U5639 (N_5639,N_5395,N_5368);
and U5640 (N_5640,N_5414,N_5410);
or U5641 (N_5641,N_5335,N_5262);
nand U5642 (N_5642,N_5457,N_5464);
xor U5643 (N_5643,N_5317,N_5305);
nand U5644 (N_5644,N_5441,N_5273);
nand U5645 (N_5645,N_5483,N_5358);
nor U5646 (N_5646,N_5261,N_5435);
or U5647 (N_5647,N_5394,N_5332);
nand U5648 (N_5648,N_5290,N_5454);
or U5649 (N_5649,N_5376,N_5293);
or U5650 (N_5650,N_5367,N_5472);
xnor U5651 (N_5651,N_5373,N_5412);
xor U5652 (N_5652,N_5478,N_5434);
xor U5653 (N_5653,N_5417,N_5284);
xor U5654 (N_5654,N_5365,N_5358);
xnor U5655 (N_5655,N_5315,N_5473);
nor U5656 (N_5656,N_5308,N_5387);
or U5657 (N_5657,N_5477,N_5478);
or U5658 (N_5658,N_5462,N_5490);
or U5659 (N_5659,N_5441,N_5461);
and U5660 (N_5660,N_5251,N_5372);
nor U5661 (N_5661,N_5450,N_5440);
xnor U5662 (N_5662,N_5421,N_5269);
and U5663 (N_5663,N_5365,N_5439);
and U5664 (N_5664,N_5288,N_5254);
nor U5665 (N_5665,N_5353,N_5414);
and U5666 (N_5666,N_5497,N_5334);
or U5667 (N_5667,N_5455,N_5364);
xnor U5668 (N_5668,N_5431,N_5383);
nand U5669 (N_5669,N_5299,N_5341);
or U5670 (N_5670,N_5477,N_5318);
nor U5671 (N_5671,N_5317,N_5358);
and U5672 (N_5672,N_5483,N_5331);
xnor U5673 (N_5673,N_5296,N_5304);
xnor U5674 (N_5674,N_5435,N_5301);
nor U5675 (N_5675,N_5454,N_5402);
nand U5676 (N_5676,N_5364,N_5317);
nand U5677 (N_5677,N_5351,N_5330);
and U5678 (N_5678,N_5292,N_5424);
xor U5679 (N_5679,N_5415,N_5328);
nor U5680 (N_5680,N_5473,N_5382);
or U5681 (N_5681,N_5352,N_5484);
xor U5682 (N_5682,N_5477,N_5305);
xnor U5683 (N_5683,N_5419,N_5402);
xor U5684 (N_5684,N_5265,N_5479);
or U5685 (N_5685,N_5477,N_5452);
nor U5686 (N_5686,N_5298,N_5281);
nand U5687 (N_5687,N_5459,N_5341);
and U5688 (N_5688,N_5434,N_5442);
nor U5689 (N_5689,N_5483,N_5295);
nand U5690 (N_5690,N_5415,N_5417);
nand U5691 (N_5691,N_5395,N_5358);
nor U5692 (N_5692,N_5255,N_5275);
nand U5693 (N_5693,N_5475,N_5288);
nand U5694 (N_5694,N_5379,N_5296);
xor U5695 (N_5695,N_5408,N_5362);
nor U5696 (N_5696,N_5269,N_5440);
nor U5697 (N_5697,N_5285,N_5258);
and U5698 (N_5698,N_5348,N_5381);
nand U5699 (N_5699,N_5471,N_5276);
nand U5700 (N_5700,N_5298,N_5406);
or U5701 (N_5701,N_5347,N_5277);
xor U5702 (N_5702,N_5267,N_5467);
xor U5703 (N_5703,N_5470,N_5332);
nand U5704 (N_5704,N_5310,N_5258);
xor U5705 (N_5705,N_5430,N_5289);
nand U5706 (N_5706,N_5273,N_5446);
or U5707 (N_5707,N_5427,N_5370);
nor U5708 (N_5708,N_5332,N_5376);
and U5709 (N_5709,N_5290,N_5301);
xnor U5710 (N_5710,N_5320,N_5398);
or U5711 (N_5711,N_5301,N_5307);
xnor U5712 (N_5712,N_5422,N_5266);
or U5713 (N_5713,N_5496,N_5331);
nor U5714 (N_5714,N_5496,N_5295);
nor U5715 (N_5715,N_5374,N_5495);
and U5716 (N_5716,N_5252,N_5275);
nor U5717 (N_5717,N_5353,N_5326);
nor U5718 (N_5718,N_5300,N_5269);
xnor U5719 (N_5719,N_5335,N_5477);
nand U5720 (N_5720,N_5297,N_5392);
xor U5721 (N_5721,N_5278,N_5403);
and U5722 (N_5722,N_5251,N_5490);
nor U5723 (N_5723,N_5485,N_5354);
and U5724 (N_5724,N_5476,N_5307);
or U5725 (N_5725,N_5356,N_5305);
or U5726 (N_5726,N_5330,N_5294);
nand U5727 (N_5727,N_5466,N_5391);
and U5728 (N_5728,N_5265,N_5389);
and U5729 (N_5729,N_5398,N_5270);
or U5730 (N_5730,N_5330,N_5436);
nor U5731 (N_5731,N_5396,N_5338);
nand U5732 (N_5732,N_5367,N_5295);
and U5733 (N_5733,N_5415,N_5498);
nand U5734 (N_5734,N_5388,N_5310);
nor U5735 (N_5735,N_5420,N_5294);
nand U5736 (N_5736,N_5331,N_5292);
or U5737 (N_5737,N_5280,N_5278);
or U5738 (N_5738,N_5273,N_5494);
xor U5739 (N_5739,N_5398,N_5413);
nor U5740 (N_5740,N_5414,N_5406);
xnor U5741 (N_5741,N_5402,N_5335);
nor U5742 (N_5742,N_5442,N_5301);
nand U5743 (N_5743,N_5391,N_5323);
nand U5744 (N_5744,N_5339,N_5435);
xnor U5745 (N_5745,N_5255,N_5391);
or U5746 (N_5746,N_5318,N_5263);
or U5747 (N_5747,N_5388,N_5371);
xnor U5748 (N_5748,N_5384,N_5336);
nor U5749 (N_5749,N_5439,N_5333);
xnor U5750 (N_5750,N_5714,N_5553);
and U5751 (N_5751,N_5634,N_5696);
nor U5752 (N_5752,N_5551,N_5718);
nand U5753 (N_5753,N_5512,N_5618);
or U5754 (N_5754,N_5691,N_5531);
nand U5755 (N_5755,N_5568,N_5626);
nand U5756 (N_5756,N_5728,N_5511);
xnor U5757 (N_5757,N_5645,N_5736);
nand U5758 (N_5758,N_5679,N_5532);
nor U5759 (N_5759,N_5555,N_5589);
nor U5760 (N_5760,N_5621,N_5707);
or U5761 (N_5761,N_5600,N_5726);
nand U5762 (N_5762,N_5594,N_5574);
and U5763 (N_5763,N_5620,N_5617);
xor U5764 (N_5764,N_5748,N_5693);
xor U5765 (N_5765,N_5543,N_5677);
xnor U5766 (N_5766,N_5662,N_5722);
xor U5767 (N_5767,N_5702,N_5501);
xnor U5768 (N_5768,N_5710,N_5742);
nand U5769 (N_5769,N_5533,N_5519);
or U5770 (N_5770,N_5647,N_5689);
xnor U5771 (N_5771,N_5661,N_5639);
and U5772 (N_5772,N_5643,N_5578);
nor U5773 (N_5773,N_5672,N_5526);
nor U5774 (N_5774,N_5516,N_5703);
nand U5775 (N_5775,N_5561,N_5562);
xnor U5776 (N_5776,N_5541,N_5690);
nor U5777 (N_5777,N_5597,N_5652);
and U5778 (N_5778,N_5517,N_5573);
xnor U5779 (N_5779,N_5687,N_5566);
nand U5780 (N_5780,N_5613,N_5666);
nand U5781 (N_5781,N_5507,N_5536);
or U5782 (N_5782,N_5596,N_5683);
and U5783 (N_5783,N_5510,N_5524);
nand U5784 (N_5784,N_5500,N_5659);
nand U5785 (N_5785,N_5513,N_5725);
nand U5786 (N_5786,N_5583,N_5654);
nand U5787 (N_5787,N_5640,N_5641);
or U5788 (N_5788,N_5546,N_5591);
or U5789 (N_5789,N_5623,N_5658);
nor U5790 (N_5790,N_5684,N_5747);
or U5791 (N_5791,N_5603,N_5646);
and U5792 (N_5792,N_5530,N_5625);
or U5793 (N_5793,N_5638,N_5649);
nand U5794 (N_5794,N_5657,N_5651);
and U5795 (N_5795,N_5538,N_5539);
or U5796 (N_5796,N_5615,N_5540);
nand U5797 (N_5797,N_5550,N_5673);
nand U5798 (N_5798,N_5609,N_5616);
nand U5799 (N_5799,N_5695,N_5588);
and U5800 (N_5800,N_5542,N_5636);
or U5801 (N_5801,N_5586,N_5572);
and U5802 (N_5802,N_5685,N_5579);
nor U5803 (N_5803,N_5614,N_5544);
xor U5804 (N_5804,N_5624,N_5606);
xnor U5805 (N_5805,N_5669,N_5528);
nor U5806 (N_5806,N_5733,N_5744);
xor U5807 (N_5807,N_5664,N_5629);
xnor U5808 (N_5808,N_5719,N_5506);
xnor U5809 (N_5809,N_5502,N_5522);
xnor U5810 (N_5810,N_5523,N_5598);
or U5811 (N_5811,N_5503,N_5716);
nand U5812 (N_5812,N_5642,N_5631);
nor U5813 (N_5813,N_5715,N_5653);
xor U5814 (N_5814,N_5701,N_5682);
xnor U5815 (N_5815,N_5717,N_5515);
nand U5816 (N_5816,N_5705,N_5565);
nand U5817 (N_5817,N_5739,N_5721);
nand U5818 (N_5818,N_5724,N_5674);
nor U5819 (N_5819,N_5698,N_5569);
nor U5820 (N_5820,N_5697,N_5730);
nand U5821 (N_5821,N_5537,N_5548);
xnor U5822 (N_5822,N_5559,N_5729);
xnor U5823 (N_5823,N_5560,N_5552);
nor U5824 (N_5824,N_5590,N_5732);
nand U5825 (N_5825,N_5740,N_5650);
or U5826 (N_5826,N_5608,N_5708);
xor U5827 (N_5827,N_5602,N_5668);
or U5828 (N_5828,N_5709,N_5700);
xnor U5829 (N_5829,N_5720,N_5656);
nor U5830 (N_5830,N_5675,N_5581);
or U5831 (N_5831,N_5622,N_5681);
nand U5832 (N_5832,N_5592,N_5655);
nand U5833 (N_5833,N_5593,N_5694);
nor U5834 (N_5834,N_5670,N_5706);
xnor U5835 (N_5835,N_5627,N_5580);
xnor U5836 (N_5836,N_5712,N_5564);
nand U5837 (N_5837,N_5563,N_5619);
nand U5838 (N_5838,N_5630,N_5723);
nand U5839 (N_5839,N_5663,N_5727);
nor U5840 (N_5840,N_5612,N_5686);
and U5841 (N_5841,N_5514,N_5678);
xnor U5842 (N_5842,N_5676,N_5688);
or U5843 (N_5843,N_5504,N_5534);
and U5844 (N_5844,N_5577,N_5680);
nand U5845 (N_5845,N_5529,N_5518);
and U5846 (N_5846,N_5505,N_5509);
nand U5847 (N_5847,N_5637,N_5587);
nand U5848 (N_5848,N_5704,N_5545);
nor U5849 (N_5849,N_5575,N_5667);
nand U5850 (N_5850,N_5521,N_5508);
nand U5851 (N_5851,N_5599,N_5628);
or U5852 (N_5852,N_5749,N_5601);
nor U5853 (N_5853,N_5660,N_5644);
nand U5854 (N_5854,N_5610,N_5731);
xor U5855 (N_5855,N_5713,N_5633);
and U5856 (N_5856,N_5554,N_5605);
nand U5857 (N_5857,N_5585,N_5527);
nand U5858 (N_5858,N_5607,N_5635);
nor U5859 (N_5859,N_5671,N_5525);
nand U5860 (N_5860,N_5558,N_5632);
or U5861 (N_5861,N_5571,N_5584);
xor U5862 (N_5862,N_5738,N_5711);
xnor U5863 (N_5863,N_5604,N_5570);
nor U5864 (N_5864,N_5743,N_5741);
nor U5865 (N_5865,N_5576,N_5734);
and U5866 (N_5866,N_5557,N_5699);
and U5867 (N_5867,N_5737,N_5746);
nor U5868 (N_5868,N_5535,N_5582);
nor U5869 (N_5869,N_5692,N_5556);
nand U5870 (N_5870,N_5547,N_5735);
nand U5871 (N_5871,N_5549,N_5648);
nor U5872 (N_5872,N_5595,N_5520);
nand U5873 (N_5873,N_5745,N_5611);
nor U5874 (N_5874,N_5665,N_5567);
nor U5875 (N_5875,N_5597,N_5629);
xnor U5876 (N_5876,N_5615,N_5566);
and U5877 (N_5877,N_5584,N_5658);
or U5878 (N_5878,N_5612,N_5673);
nor U5879 (N_5879,N_5670,N_5565);
nor U5880 (N_5880,N_5622,N_5706);
or U5881 (N_5881,N_5513,N_5522);
xor U5882 (N_5882,N_5591,N_5515);
xnor U5883 (N_5883,N_5639,N_5720);
or U5884 (N_5884,N_5504,N_5562);
and U5885 (N_5885,N_5657,N_5658);
and U5886 (N_5886,N_5695,N_5736);
xnor U5887 (N_5887,N_5684,N_5634);
xor U5888 (N_5888,N_5713,N_5562);
or U5889 (N_5889,N_5732,N_5676);
or U5890 (N_5890,N_5517,N_5680);
or U5891 (N_5891,N_5538,N_5624);
or U5892 (N_5892,N_5699,N_5562);
nor U5893 (N_5893,N_5699,N_5573);
nand U5894 (N_5894,N_5730,N_5748);
nand U5895 (N_5895,N_5531,N_5574);
or U5896 (N_5896,N_5690,N_5503);
nor U5897 (N_5897,N_5630,N_5721);
nand U5898 (N_5898,N_5657,N_5587);
and U5899 (N_5899,N_5651,N_5571);
nor U5900 (N_5900,N_5727,N_5636);
nor U5901 (N_5901,N_5571,N_5626);
and U5902 (N_5902,N_5600,N_5637);
nand U5903 (N_5903,N_5659,N_5640);
nor U5904 (N_5904,N_5624,N_5586);
and U5905 (N_5905,N_5579,N_5714);
nand U5906 (N_5906,N_5530,N_5703);
or U5907 (N_5907,N_5605,N_5641);
nand U5908 (N_5908,N_5713,N_5531);
nand U5909 (N_5909,N_5742,N_5749);
nand U5910 (N_5910,N_5622,N_5606);
xnor U5911 (N_5911,N_5620,N_5706);
and U5912 (N_5912,N_5605,N_5505);
xnor U5913 (N_5913,N_5655,N_5610);
or U5914 (N_5914,N_5664,N_5643);
xor U5915 (N_5915,N_5731,N_5521);
nand U5916 (N_5916,N_5726,N_5727);
nor U5917 (N_5917,N_5596,N_5720);
xor U5918 (N_5918,N_5682,N_5704);
or U5919 (N_5919,N_5634,N_5542);
nor U5920 (N_5920,N_5632,N_5590);
and U5921 (N_5921,N_5612,N_5620);
and U5922 (N_5922,N_5620,N_5711);
or U5923 (N_5923,N_5675,N_5707);
and U5924 (N_5924,N_5737,N_5568);
nand U5925 (N_5925,N_5544,N_5509);
or U5926 (N_5926,N_5689,N_5590);
xor U5927 (N_5927,N_5678,N_5740);
nand U5928 (N_5928,N_5733,N_5648);
nand U5929 (N_5929,N_5658,N_5659);
or U5930 (N_5930,N_5501,N_5599);
and U5931 (N_5931,N_5606,N_5543);
nor U5932 (N_5932,N_5648,N_5538);
and U5933 (N_5933,N_5553,N_5584);
and U5934 (N_5934,N_5644,N_5656);
nand U5935 (N_5935,N_5614,N_5511);
and U5936 (N_5936,N_5637,N_5655);
or U5937 (N_5937,N_5638,N_5583);
nand U5938 (N_5938,N_5682,N_5727);
xnor U5939 (N_5939,N_5520,N_5560);
and U5940 (N_5940,N_5507,N_5607);
nand U5941 (N_5941,N_5651,N_5524);
xnor U5942 (N_5942,N_5578,N_5616);
nand U5943 (N_5943,N_5518,N_5642);
nand U5944 (N_5944,N_5599,N_5741);
nor U5945 (N_5945,N_5554,N_5642);
nand U5946 (N_5946,N_5667,N_5556);
and U5947 (N_5947,N_5695,N_5729);
and U5948 (N_5948,N_5506,N_5643);
and U5949 (N_5949,N_5716,N_5681);
or U5950 (N_5950,N_5673,N_5667);
and U5951 (N_5951,N_5693,N_5504);
xor U5952 (N_5952,N_5732,N_5602);
nand U5953 (N_5953,N_5605,N_5663);
xnor U5954 (N_5954,N_5543,N_5634);
nand U5955 (N_5955,N_5645,N_5663);
nand U5956 (N_5956,N_5540,N_5578);
xor U5957 (N_5957,N_5684,N_5512);
xor U5958 (N_5958,N_5616,N_5614);
and U5959 (N_5959,N_5744,N_5515);
and U5960 (N_5960,N_5549,N_5716);
xor U5961 (N_5961,N_5734,N_5556);
or U5962 (N_5962,N_5623,N_5644);
nand U5963 (N_5963,N_5642,N_5592);
xor U5964 (N_5964,N_5611,N_5721);
and U5965 (N_5965,N_5607,N_5566);
nand U5966 (N_5966,N_5730,N_5620);
and U5967 (N_5967,N_5600,N_5534);
and U5968 (N_5968,N_5601,N_5635);
nor U5969 (N_5969,N_5580,N_5632);
or U5970 (N_5970,N_5669,N_5594);
xnor U5971 (N_5971,N_5646,N_5641);
xnor U5972 (N_5972,N_5578,N_5713);
and U5973 (N_5973,N_5681,N_5566);
or U5974 (N_5974,N_5661,N_5700);
xor U5975 (N_5975,N_5501,N_5608);
and U5976 (N_5976,N_5679,N_5717);
nand U5977 (N_5977,N_5586,N_5590);
nand U5978 (N_5978,N_5662,N_5619);
and U5979 (N_5979,N_5592,N_5605);
and U5980 (N_5980,N_5554,N_5549);
nand U5981 (N_5981,N_5550,N_5508);
nand U5982 (N_5982,N_5690,N_5673);
and U5983 (N_5983,N_5514,N_5661);
and U5984 (N_5984,N_5740,N_5713);
nand U5985 (N_5985,N_5728,N_5615);
or U5986 (N_5986,N_5736,N_5687);
and U5987 (N_5987,N_5561,N_5672);
nand U5988 (N_5988,N_5602,N_5589);
and U5989 (N_5989,N_5737,N_5655);
xnor U5990 (N_5990,N_5553,N_5504);
or U5991 (N_5991,N_5605,N_5744);
and U5992 (N_5992,N_5635,N_5671);
nor U5993 (N_5993,N_5555,N_5682);
or U5994 (N_5994,N_5677,N_5576);
and U5995 (N_5995,N_5650,N_5668);
xor U5996 (N_5996,N_5656,N_5548);
and U5997 (N_5997,N_5657,N_5635);
nand U5998 (N_5998,N_5569,N_5735);
or U5999 (N_5999,N_5559,N_5539);
or U6000 (N_6000,N_5758,N_5948);
and U6001 (N_6001,N_5932,N_5945);
xnor U6002 (N_6002,N_5844,N_5913);
or U6003 (N_6003,N_5806,N_5953);
nand U6004 (N_6004,N_5996,N_5841);
nor U6005 (N_6005,N_5918,N_5791);
xor U6006 (N_6006,N_5797,N_5830);
nand U6007 (N_6007,N_5760,N_5924);
nand U6008 (N_6008,N_5979,N_5891);
or U6009 (N_6009,N_5973,N_5802);
nor U6010 (N_6010,N_5867,N_5951);
nand U6011 (N_6011,N_5858,N_5870);
xnor U6012 (N_6012,N_5818,N_5795);
nor U6013 (N_6013,N_5845,N_5936);
nor U6014 (N_6014,N_5976,N_5880);
nor U6015 (N_6015,N_5974,N_5952);
xor U6016 (N_6016,N_5782,N_5939);
nor U6017 (N_6017,N_5804,N_5846);
nand U6018 (N_6018,N_5832,N_5761);
nor U6019 (N_6019,N_5889,N_5912);
or U6020 (N_6020,N_5834,N_5815);
nor U6021 (N_6021,N_5772,N_5800);
nor U6022 (N_6022,N_5878,N_5957);
or U6023 (N_6023,N_5768,N_5794);
nor U6024 (N_6024,N_5927,N_5935);
nand U6025 (N_6025,N_5993,N_5781);
nand U6026 (N_6026,N_5971,N_5915);
or U6027 (N_6027,N_5970,N_5926);
and U6028 (N_6028,N_5963,N_5958);
nor U6029 (N_6029,N_5868,N_5986);
nor U6030 (N_6030,N_5966,N_5871);
xnor U6031 (N_6031,N_5967,N_5810);
nand U6032 (N_6032,N_5763,N_5774);
xnor U6033 (N_6033,N_5849,N_5903);
or U6034 (N_6034,N_5929,N_5798);
or U6035 (N_6035,N_5778,N_5854);
or U6036 (N_6036,N_5920,N_5765);
xor U6037 (N_6037,N_5848,N_5754);
nor U6038 (N_6038,N_5999,N_5808);
nand U6039 (N_6039,N_5792,N_5885);
nand U6040 (N_6040,N_5817,N_5931);
and U6041 (N_6041,N_5910,N_5998);
nor U6042 (N_6042,N_5786,N_5865);
nor U6043 (N_6043,N_5907,N_5762);
xor U6044 (N_6044,N_5828,N_5895);
xnor U6045 (N_6045,N_5975,N_5984);
nand U6046 (N_6046,N_5886,N_5835);
nor U6047 (N_6047,N_5964,N_5888);
nor U6048 (N_6048,N_5839,N_5937);
nand U6049 (N_6049,N_5938,N_5807);
and U6050 (N_6050,N_5960,N_5972);
xor U6051 (N_6051,N_5803,N_5823);
nor U6052 (N_6052,N_5850,N_5801);
and U6053 (N_6053,N_5842,N_5836);
xnor U6054 (N_6054,N_5769,N_5900);
nor U6055 (N_6055,N_5940,N_5847);
or U6056 (N_6056,N_5787,N_5862);
xor U6057 (N_6057,N_5969,N_5827);
xor U6058 (N_6058,N_5876,N_5946);
xnor U6059 (N_6059,N_5879,N_5959);
nor U6060 (N_6060,N_5991,N_5892);
and U6061 (N_6061,N_5904,N_5997);
nand U6062 (N_6062,N_5829,N_5825);
xnor U6063 (N_6063,N_5954,N_5866);
xnor U6064 (N_6064,N_5788,N_5987);
nand U6065 (N_6065,N_5775,N_5923);
xor U6066 (N_6066,N_5942,N_5881);
or U6067 (N_6067,N_5864,N_5752);
nand U6068 (N_6068,N_5983,N_5820);
nand U6069 (N_6069,N_5988,N_5790);
or U6070 (N_6070,N_5980,N_5965);
nor U6071 (N_6071,N_5899,N_5783);
nand U6072 (N_6072,N_5811,N_5950);
or U6073 (N_6073,N_5821,N_5919);
or U6074 (N_6074,N_5793,N_5838);
xnor U6075 (N_6075,N_5921,N_5814);
nand U6076 (N_6076,N_5859,N_5776);
xor U6077 (N_6077,N_5757,N_5855);
or U6078 (N_6078,N_5977,N_5833);
and U6079 (N_6079,N_5861,N_5962);
and U6080 (N_6080,N_5785,N_5956);
xnor U6081 (N_6081,N_5819,N_5943);
xnor U6082 (N_6082,N_5796,N_5887);
nand U6083 (N_6083,N_5750,N_5771);
and U6084 (N_6084,N_5994,N_5989);
or U6085 (N_6085,N_5933,N_5961);
nor U6086 (N_6086,N_5934,N_5930);
nand U6087 (N_6087,N_5767,N_5902);
nand U6088 (N_6088,N_5857,N_5789);
nand U6089 (N_6089,N_5826,N_5822);
nand U6090 (N_6090,N_5853,N_5756);
and U6091 (N_6091,N_5851,N_5824);
or U6092 (N_6092,N_5909,N_5856);
or U6093 (N_6093,N_5914,N_5869);
xnor U6094 (N_6094,N_5917,N_5908);
and U6095 (N_6095,N_5901,N_5884);
or U6096 (N_6096,N_5894,N_5906);
nand U6097 (N_6097,N_5816,N_5982);
xnor U6098 (N_6098,N_5922,N_5773);
and U6099 (N_6099,N_5766,N_5944);
or U6100 (N_6100,N_5770,N_5751);
xor U6101 (N_6101,N_5837,N_5759);
or U6102 (N_6102,N_5947,N_5777);
nand U6103 (N_6103,N_5882,N_5978);
nand U6104 (N_6104,N_5784,N_5755);
nand U6105 (N_6105,N_5928,N_5753);
or U6106 (N_6106,N_5896,N_5872);
or U6107 (N_6107,N_5893,N_5877);
nor U6108 (N_6108,N_5898,N_5831);
nor U6109 (N_6109,N_5843,N_5874);
or U6110 (N_6110,N_5941,N_5985);
and U6111 (N_6111,N_5990,N_5873);
or U6112 (N_6112,N_5955,N_5905);
nor U6113 (N_6113,N_5968,N_5949);
or U6114 (N_6114,N_5779,N_5799);
nand U6115 (N_6115,N_5981,N_5992);
xor U6116 (N_6116,N_5812,N_5863);
xor U6117 (N_6117,N_5860,N_5925);
or U6118 (N_6118,N_5852,N_5764);
nor U6119 (N_6119,N_5911,N_5875);
and U6120 (N_6120,N_5809,N_5840);
nor U6121 (N_6121,N_5883,N_5897);
nand U6122 (N_6122,N_5916,N_5995);
xor U6123 (N_6123,N_5780,N_5805);
xnor U6124 (N_6124,N_5813,N_5890);
or U6125 (N_6125,N_5936,N_5906);
or U6126 (N_6126,N_5931,N_5911);
nand U6127 (N_6127,N_5820,N_5787);
nand U6128 (N_6128,N_5769,N_5841);
nor U6129 (N_6129,N_5750,N_5855);
nand U6130 (N_6130,N_5966,N_5949);
and U6131 (N_6131,N_5822,N_5775);
nor U6132 (N_6132,N_5981,N_5766);
nor U6133 (N_6133,N_5984,N_5832);
or U6134 (N_6134,N_5861,N_5967);
and U6135 (N_6135,N_5757,N_5802);
or U6136 (N_6136,N_5948,N_5931);
and U6137 (N_6137,N_5987,N_5930);
nand U6138 (N_6138,N_5939,N_5997);
nand U6139 (N_6139,N_5769,N_5829);
nand U6140 (N_6140,N_5884,N_5863);
or U6141 (N_6141,N_5876,N_5993);
xnor U6142 (N_6142,N_5803,N_5910);
and U6143 (N_6143,N_5772,N_5786);
and U6144 (N_6144,N_5775,N_5964);
or U6145 (N_6145,N_5997,N_5774);
nand U6146 (N_6146,N_5846,N_5982);
or U6147 (N_6147,N_5789,N_5780);
or U6148 (N_6148,N_5968,N_5778);
nand U6149 (N_6149,N_5822,N_5907);
nand U6150 (N_6150,N_5888,N_5773);
or U6151 (N_6151,N_5840,N_5974);
nor U6152 (N_6152,N_5870,N_5981);
and U6153 (N_6153,N_5968,N_5805);
nor U6154 (N_6154,N_5870,N_5963);
nand U6155 (N_6155,N_5981,N_5984);
xnor U6156 (N_6156,N_5907,N_5939);
xnor U6157 (N_6157,N_5886,N_5991);
and U6158 (N_6158,N_5826,N_5789);
or U6159 (N_6159,N_5761,N_5799);
or U6160 (N_6160,N_5790,N_5917);
nor U6161 (N_6161,N_5965,N_5976);
nand U6162 (N_6162,N_5767,N_5848);
nor U6163 (N_6163,N_5878,N_5782);
nand U6164 (N_6164,N_5758,N_5810);
xnor U6165 (N_6165,N_5790,N_5825);
and U6166 (N_6166,N_5804,N_5821);
or U6167 (N_6167,N_5761,N_5864);
and U6168 (N_6168,N_5950,N_5802);
and U6169 (N_6169,N_5877,N_5929);
nand U6170 (N_6170,N_5899,N_5910);
or U6171 (N_6171,N_5969,N_5825);
and U6172 (N_6172,N_5979,N_5804);
or U6173 (N_6173,N_5759,N_5835);
and U6174 (N_6174,N_5856,N_5828);
nand U6175 (N_6175,N_5843,N_5955);
xor U6176 (N_6176,N_5960,N_5939);
or U6177 (N_6177,N_5879,N_5784);
or U6178 (N_6178,N_5887,N_5922);
nor U6179 (N_6179,N_5858,N_5938);
or U6180 (N_6180,N_5848,N_5840);
nand U6181 (N_6181,N_5879,N_5910);
nor U6182 (N_6182,N_5791,N_5878);
nor U6183 (N_6183,N_5845,N_5860);
nor U6184 (N_6184,N_5811,N_5923);
and U6185 (N_6185,N_5913,N_5823);
xor U6186 (N_6186,N_5951,N_5782);
xnor U6187 (N_6187,N_5858,N_5759);
or U6188 (N_6188,N_5932,N_5816);
nand U6189 (N_6189,N_5821,N_5965);
or U6190 (N_6190,N_5802,N_5883);
xor U6191 (N_6191,N_5794,N_5862);
nand U6192 (N_6192,N_5820,N_5760);
xnor U6193 (N_6193,N_5888,N_5916);
or U6194 (N_6194,N_5917,N_5909);
or U6195 (N_6195,N_5810,N_5898);
xor U6196 (N_6196,N_5765,N_5970);
or U6197 (N_6197,N_5781,N_5809);
nor U6198 (N_6198,N_5775,N_5846);
or U6199 (N_6199,N_5926,N_5874);
or U6200 (N_6200,N_5881,N_5957);
and U6201 (N_6201,N_5787,N_5872);
nor U6202 (N_6202,N_5819,N_5974);
nand U6203 (N_6203,N_5825,N_5800);
or U6204 (N_6204,N_5781,N_5770);
and U6205 (N_6205,N_5959,N_5910);
nor U6206 (N_6206,N_5941,N_5777);
or U6207 (N_6207,N_5800,N_5891);
or U6208 (N_6208,N_5910,N_5763);
xor U6209 (N_6209,N_5906,N_5925);
or U6210 (N_6210,N_5985,N_5861);
and U6211 (N_6211,N_5941,N_5771);
nor U6212 (N_6212,N_5873,N_5770);
nand U6213 (N_6213,N_5788,N_5934);
or U6214 (N_6214,N_5843,N_5994);
xor U6215 (N_6215,N_5877,N_5992);
nor U6216 (N_6216,N_5934,N_5895);
or U6217 (N_6217,N_5918,N_5981);
nand U6218 (N_6218,N_5885,N_5781);
xor U6219 (N_6219,N_5949,N_5853);
or U6220 (N_6220,N_5902,N_5905);
nand U6221 (N_6221,N_5923,N_5926);
nand U6222 (N_6222,N_5827,N_5991);
xnor U6223 (N_6223,N_5948,N_5965);
nor U6224 (N_6224,N_5774,N_5768);
nand U6225 (N_6225,N_5853,N_5978);
nor U6226 (N_6226,N_5773,N_5842);
and U6227 (N_6227,N_5794,N_5770);
or U6228 (N_6228,N_5886,N_5766);
or U6229 (N_6229,N_5905,N_5783);
and U6230 (N_6230,N_5812,N_5859);
and U6231 (N_6231,N_5845,N_5800);
and U6232 (N_6232,N_5962,N_5850);
or U6233 (N_6233,N_5925,N_5792);
xnor U6234 (N_6234,N_5870,N_5777);
and U6235 (N_6235,N_5861,N_5994);
and U6236 (N_6236,N_5927,N_5851);
or U6237 (N_6237,N_5801,N_5862);
xor U6238 (N_6238,N_5809,N_5889);
or U6239 (N_6239,N_5991,N_5750);
or U6240 (N_6240,N_5855,N_5953);
or U6241 (N_6241,N_5938,N_5978);
or U6242 (N_6242,N_5888,N_5921);
nand U6243 (N_6243,N_5887,N_5944);
nor U6244 (N_6244,N_5769,N_5757);
xnor U6245 (N_6245,N_5764,N_5825);
nand U6246 (N_6246,N_5851,N_5875);
xor U6247 (N_6247,N_5945,N_5775);
nor U6248 (N_6248,N_5979,N_5801);
nand U6249 (N_6249,N_5775,N_5783);
xnor U6250 (N_6250,N_6124,N_6072);
nand U6251 (N_6251,N_6184,N_6240);
nand U6252 (N_6252,N_6014,N_6189);
or U6253 (N_6253,N_6019,N_6183);
nand U6254 (N_6254,N_6174,N_6077);
nand U6255 (N_6255,N_6016,N_6045);
nand U6256 (N_6256,N_6056,N_6148);
and U6257 (N_6257,N_6241,N_6228);
or U6258 (N_6258,N_6164,N_6041);
and U6259 (N_6259,N_6073,N_6139);
and U6260 (N_6260,N_6163,N_6201);
or U6261 (N_6261,N_6219,N_6125);
or U6262 (N_6262,N_6243,N_6051);
and U6263 (N_6263,N_6237,N_6210);
xor U6264 (N_6264,N_6142,N_6030);
or U6265 (N_6265,N_6234,N_6246);
nor U6266 (N_6266,N_6196,N_6160);
nand U6267 (N_6267,N_6191,N_6082);
or U6268 (N_6268,N_6070,N_6166);
and U6269 (N_6269,N_6224,N_6040);
nand U6270 (N_6270,N_6225,N_6043);
and U6271 (N_6271,N_6169,N_6068);
nor U6272 (N_6272,N_6107,N_6208);
or U6273 (N_6273,N_6116,N_6104);
nor U6274 (N_6274,N_6145,N_6152);
and U6275 (N_6275,N_6007,N_6170);
and U6276 (N_6276,N_6144,N_6121);
or U6277 (N_6277,N_6231,N_6071);
or U6278 (N_6278,N_6001,N_6146);
and U6279 (N_6279,N_6226,N_6161);
or U6280 (N_6280,N_6044,N_6110);
and U6281 (N_6281,N_6180,N_6186);
and U6282 (N_6282,N_6054,N_6049);
xor U6283 (N_6283,N_6017,N_6179);
nor U6284 (N_6284,N_6015,N_6046);
or U6285 (N_6285,N_6010,N_6035);
nand U6286 (N_6286,N_6178,N_6118);
nand U6287 (N_6287,N_6000,N_6157);
nand U6288 (N_6288,N_6165,N_6091);
nor U6289 (N_6289,N_6038,N_6022);
and U6290 (N_6290,N_6233,N_6206);
nand U6291 (N_6291,N_6079,N_6111);
nand U6292 (N_6292,N_6136,N_6052);
nand U6293 (N_6293,N_6032,N_6130);
or U6294 (N_6294,N_6090,N_6102);
nand U6295 (N_6295,N_6173,N_6100);
nand U6296 (N_6296,N_6115,N_6135);
or U6297 (N_6297,N_6171,N_6021);
nor U6298 (N_6298,N_6209,N_6167);
or U6299 (N_6299,N_6057,N_6013);
or U6300 (N_6300,N_6245,N_6024);
xnor U6301 (N_6301,N_6006,N_6080);
nand U6302 (N_6302,N_6204,N_6195);
nand U6303 (N_6303,N_6222,N_6012);
nor U6304 (N_6304,N_6004,N_6154);
and U6305 (N_6305,N_6093,N_6158);
nor U6306 (N_6306,N_6060,N_6203);
nand U6307 (N_6307,N_6005,N_6112);
xnor U6308 (N_6308,N_6064,N_6009);
xor U6309 (N_6309,N_6036,N_6128);
or U6310 (N_6310,N_6094,N_6211);
nand U6311 (N_6311,N_6058,N_6229);
nand U6312 (N_6312,N_6027,N_6218);
or U6313 (N_6313,N_6141,N_6114);
or U6314 (N_6314,N_6248,N_6202);
xnor U6315 (N_6315,N_6159,N_6087);
nor U6316 (N_6316,N_6227,N_6101);
nor U6317 (N_6317,N_6134,N_6236);
nand U6318 (N_6318,N_6177,N_6081);
or U6319 (N_6319,N_6023,N_6132);
and U6320 (N_6320,N_6108,N_6039);
nand U6321 (N_6321,N_6213,N_6175);
nor U6322 (N_6322,N_6042,N_6232);
and U6323 (N_6323,N_6026,N_6061);
xnor U6324 (N_6324,N_6053,N_6031);
nor U6325 (N_6325,N_6048,N_6181);
and U6326 (N_6326,N_6123,N_6050);
nand U6327 (N_6327,N_6214,N_6244);
and U6328 (N_6328,N_6190,N_6140);
xnor U6329 (N_6329,N_6119,N_6120);
xnor U6330 (N_6330,N_6182,N_6069);
xor U6331 (N_6331,N_6193,N_6063);
or U6332 (N_6332,N_6047,N_6137);
and U6333 (N_6333,N_6176,N_6150);
nor U6334 (N_6334,N_6127,N_6002);
and U6335 (N_6335,N_6088,N_6133);
xnor U6336 (N_6336,N_6083,N_6092);
or U6337 (N_6337,N_6067,N_6003);
nand U6338 (N_6338,N_6065,N_6008);
or U6339 (N_6339,N_6207,N_6113);
nor U6340 (N_6340,N_6199,N_6223);
nor U6341 (N_6341,N_6099,N_6095);
nor U6342 (N_6342,N_6200,N_6129);
and U6343 (N_6343,N_6242,N_6089);
nor U6344 (N_6344,N_6221,N_6230);
nand U6345 (N_6345,N_6033,N_6034);
or U6346 (N_6346,N_6062,N_6075);
and U6347 (N_6347,N_6153,N_6162);
and U6348 (N_6348,N_6247,N_6098);
and U6349 (N_6349,N_6122,N_6187);
or U6350 (N_6350,N_6212,N_6109);
nand U6351 (N_6351,N_6205,N_6025);
and U6352 (N_6352,N_6249,N_6198);
and U6353 (N_6353,N_6085,N_6097);
and U6354 (N_6354,N_6028,N_6106);
or U6355 (N_6355,N_6235,N_6151);
or U6356 (N_6356,N_6155,N_6117);
or U6357 (N_6357,N_6194,N_6188);
xor U6358 (N_6358,N_6238,N_6197);
nor U6359 (N_6359,N_6215,N_6018);
or U6360 (N_6360,N_6172,N_6192);
xor U6361 (N_6361,N_6239,N_6086);
nand U6362 (N_6362,N_6103,N_6066);
nor U6363 (N_6363,N_6185,N_6076);
xnor U6364 (N_6364,N_6084,N_6059);
xnor U6365 (N_6365,N_6029,N_6156);
nor U6366 (N_6366,N_6143,N_6147);
and U6367 (N_6367,N_6126,N_6168);
or U6368 (N_6368,N_6220,N_6078);
or U6369 (N_6369,N_6074,N_6149);
nand U6370 (N_6370,N_6217,N_6216);
and U6371 (N_6371,N_6011,N_6037);
xor U6372 (N_6372,N_6055,N_6020);
xnor U6373 (N_6373,N_6105,N_6138);
nand U6374 (N_6374,N_6096,N_6131);
xor U6375 (N_6375,N_6122,N_6090);
nor U6376 (N_6376,N_6003,N_6136);
nor U6377 (N_6377,N_6071,N_6153);
nor U6378 (N_6378,N_6117,N_6101);
or U6379 (N_6379,N_6203,N_6189);
nand U6380 (N_6380,N_6001,N_6096);
nor U6381 (N_6381,N_6209,N_6067);
and U6382 (N_6382,N_6091,N_6030);
and U6383 (N_6383,N_6014,N_6086);
and U6384 (N_6384,N_6235,N_6004);
nor U6385 (N_6385,N_6089,N_6162);
xor U6386 (N_6386,N_6017,N_6170);
and U6387 (N_6387,N_6232,N_6083);
or U6388 (N_6388,N_6170,N_6008);
nand U6389 (N_6389,N_6207,N_6086);
nor U6390 (N_6390,N_6164,N_6118);
nor U6391 (N_6391,N_6095,N_6231);
nor U6392 (N_6392,N_6094,N_6137);
and U6393 (N_6393,N_6099,N_6125);
xnor U6394 (N_6394,N_6119,N_6012);
and U6395 (N_6395,N_6056,N_6099);
xor U6396 (N_6396,N_6232,N_6149);
and U6397 (N_6397,N_6235,N_6084);
nor U6398 (N_6398,N_6128,N_6242);
and U6399 (N_6399,N_6202,N_6059);
or U6400 (N_6400,N_6159,N_6224);
or U6401 (N_6401,N_6177,N_6205);
or U6402 (N_6402,N_6204,N_6181);
or U6403 (N_6403,N_6126,N_6163);
and U6404 (N_6404,N_6163,N_6077);
and U6405 (N_6405,N_6206,N_6209);
nand U6406 (N_6406,N_6144,N_6181);
or U6407 (N_6407,N_6154,N_6196);
or U6408 (N_6408,N_6070,N_6132);
and U6409 (N_6409,N_6198,N_6219);
nand U6410 (N_6410,N_6101,N_6161);
and U6411 (N_6411,N_6066,N_6159);
or U6412 (N_6412,N_6130,N_6091);
and U6413 (N_6413,N_6132,N_6081);
and U6414 (N_6414,N_6215,N_6081);
nor U6415 (N_6415,N_6118,N_6130);
nor U6416 (N_6416,N_6090,N_6124);
nand U6417 (N_6417,N_6093,N_6052);
nand U6418 (N_6418,N_6058,N_6022);
nand U6419 (N_6419,N_6237,N_6219);
xor U6420 (N_6420,N_6087,N_6200);
nor U6421 (N_6421,N_6177,N_6178);
xor U6422 (N_6422,N_6129,N_6082);
xnor U6423 (N_6423,N_6074,N_6173);
nor U6424 (N_6424,N_6075,N_6206);
nor U6425 (N_6425,N_6120,N_6027);
or U6426 (N_6426,N_6161,N_6197);
nor U6427 (N_6427,N_6136,N_6038);
nand U6428 (N_6428,N_6072,N_6102);
nand U6429 (N_6429,N_6215,N_6167);
xnor U6430 (N_6430,N_6179,N_6079);
and U6431 (N_6431,N_6033,N_6106);
nand U6432 (N_6432,N_6162,N_6033);
nor U6433 (N_6433,N_6176,N_6011);
xor U6434 (N_6434,N_6061,N_6152);
or U6435 (N_6435,N_6228,N_6076);
nor U6436 (N_6436,N_6015,N_6004);
nand U6437 (N_6437,N_6058,N_6026);
nor U6438 (N_6438,N_6009,N_6207);
nand U6439 (N_6439,N_6136,N_6218);
or U6440 (N_6440,N_6058,N_6105);
or U6441 (N_6441,N_6012,N_6172);
and U6442 (N_6442,N_6086,N_6221);
and U6443 (N_6443,N_6240,N_6090);
or U6444 (N_6444,N_6005,N_6010);
and U6445 (N_6445,N_6206,N_6100);
xor U6446 (N_6446,N_6186,N_6116);
nor U6447 (N_6447,N_6049,N_6050);
or U6448 (N_6448,N_6127,N_6216);
and U6449 (N_6449,N_6186,N_6053);
nor U6450 (N_6450,N_6225,N_6014);
and U6451 (N_6451,N_6198,N_6213);
or U6452 (N_6452,N_6163,N_6032);
or U6453 (N_6453,N_6006,N_6063);
or U6454 (N_6454,N_6090,N_6116);
or U6455 (N_6455,N_6041,N_6147);
xnor U6456 (N_6456,N_6225,N_6218);
nand U6457 (N_6457,N_6137,N_6163);
nor U6458 (N_6458,N_6085,N_6059);
and U6459 (N_6459,N_6225,N_6033);
xnor U6460 (N_6460,N_6061,N_6228);
nand U6461 (N_6461,N_6135,N_6107);
nor U6462 (N_6462,N_6046,N_6097);
and U6463 (N_6463,N_6104,N_6212);
nor U6464 (N_6464,N_6092,N_6158);
or U6465 (N_6465,N_6052,N_6248);
nor U6466 (N_6466,N_6124,N_6112);
and U6467 (N_6467,N_6105,N_6119);
xor U6468 (N_6468,N_6110,N_6097);
xnor U6469 (N_6469,N_6109,N_6226);
nand U6470 (N_6470,N_6155,N_6019);
and U6471 (N_6471,N_6051,N_6146);
nand U6472 (N_6472,N_6205,N_6050);
nand U6473 (N_6473,N_6224,N_6061);
and U6474 (N_6474,N_6037,N_6133);
nor U6475 (N_6475,N_6230,N_6008);
nand U6476 (N_6476,N_6174,N_6114);
xnor U6477 (N_6477,N_6087,N_6036);
nand U6478 (N_6478,N_6137,N_6000);
nor U6479 (N_6479,N_6098,N_6084);
nand U6480 (N_6480,N_6214,N_6053);
nand U6481 (N_6481,N_6209,N_6050);
nor U6482 (N_6482,N_6075,N_6244);
xnor U6483 (N_6483,N_6035,N_6076);
nor U6484 (N_6484,N_6187,N_6229);
xor U6485 (N_6485,N_6148,N_6063);
or U6486 (N_6486,N_6064,N_6191);
nor U6487 (N_6487,N_6134,N_6075);
or U6488 (N_6488,N_6174,N_6078);
nor U6489 (N_6489,N_6063,N_6041);
nand U6490 (N_6490,N_6066,N_6208);
xor U6491 (N_6491,N_6132,N_6076);
xnor U6492 (N_6492,N_6133,N_6193);
and U6493 (N_6493,N_6202,N_6165);
and U6494 (N_6494,N_6143,N_6148);
and U6495 (N_6495,N_6208,N_6011);
nor U6496 (N_6496,N_6096,N_6133);
and U6497 (N_6497,N_6144,N_6015);
nand U6498 (N_6498,N_6007,N_6077);
and U6499 (N_6499,N_6122,N_6082);
nand U6500 (N_6500,N_6450,N_6397);
xnor U6501 (N_6501,N_6269,N_6388);
or U6502 (N_6502,N_6446,N_6255);
or U6503 (N_6503,N_6316,N_6320);
and U6504 (N_6504,N_6445,N_6370);
nor U6505 (N_6505,N_6404,N_6338);
nand U6506 (N_6506,N_6305,N_6321);
xnor U6507 (N_6507,N_6422,N_6266);
nand U6508 (N_6508,N_6265,N_6284);
xor U6509 (N_6509,N_6356,N_6420);
and U6510 (N_6510,N_6490,N_6415);
nor U6511 (N_6511,N_6461,N_6386);
xnor U6512 (N_6512,N_6367,N_6385);
xor U6513 (N_6513,N_6436,N_6278);
or U6514 (N_6514,N_6304,N_6492);
nor U6515 (N_6515,N_6317,N_6369);
or U6516 (N_6516,N_6300,N_6444);
nand U6517 (N_6517,N_6330,N_6270);
nor U6518 (N_6518,N_6279,N_6467);
nand U6519 (N_6519,N_6368,N_6275);
and U6520 (N_6520,N_6395,N_6455);
and U6521 (N_6521,N_6495,N_6361);
or U6522 (N_6522,N_6406,N_6257);
nand U6523 (N_6523,N_6328,N_6405);
or U6524 (N_6524,N_6417,N_6437);
nor U6525 (N_6525,N_6486,N_6323);
nand U6526 (N_6526,N_6345,N_6390);
xnor U6527 (N_6527,N_6448,N_6440);
xor U6528 (N_6528,N_6379,N_6303);
or U6529 (N_6529,N_6424,N_6343);
nand U6530 (N_6530,N_6340,N_6376);
nand U6531 (N_6531,N_6472,N_6315);
nor U6532 (N_6532,N_6362,N_6332);
xnor U6533 (N_6533,N_6423,N_6347);
nand U6534 (N_6534,N_6457,N_6425);
nand U6535 (N_6535,N_6310,N_6289);
nor U6536 (N_6536,N_6308,N_6413);
nand U6537 (N_6537,N_6476,N_6274);
nor U6538 (N_6538,N_6337,N_6479);
or U6539 (N_6539,N_6253,N_6291);
xor U6540 (N_6540,N_6276,N_6416);
nor U6541 (N_6541,N_6375,N_6348);
and U6542 (N_6542,N_6401,N_6427);
nor U6543 (N_6543,N_6473,N_6281);
xor U6544 (N_6544,N_6288,N_6329);
or U6545 (N_6545,N_6497,N_6311);
nor U6546 (N_6546,N_6392,N_6491);
or U6547 (N_6547,N_6421,N_6418);
nor U6548 (N_6548,N_6434,N_6474);
and U6549 (N_6549,N_6261,N_6327);
nor U6550 (N_6550,N_6494,N_6373);
xor U6551 (N_6551,N_6341,N_6384);
or U6552 (N_6552,N_6358,N_6426);
xnor U6553 (N_6553,N_6339,N_6410);
or U6554 (N_6554,N_6258,N_6462);
nand U6555 (N_6555,N_6283,N_6357);
xor U6556 (N_6556,N_6334,N_6351);
nand U6557 (N_6557,N_6331,N_6353);
xor U6558 (N_6558,N_6391,N_6471);
or U6559 (N_6559,N_6380,N_6251);
or U6560 (N_6560,N_6447,N_6412);
or U6561 (N_6561,N_6419,N_6302);
and U6562 (N_6562,N_6458,N_6371);
nor U6563 (N_6563,N_6408,N_6484);
xnor U6564 (N_6564,N_6293,N_6411);
xor U6565 (N_6565,N_6493,N_6359);
and U6566 (N_6566,N_6483,N_6468);
xor U6567 (N_6567,N_6326,N_6459);
xor U6568 (N_6568,N_6460,N_6451);
xnor U6569 (N_6569,N_6272,N_6453);
nand U6570 (N_6570,N_6350,N_6499);
nor U6571 (N_6571,N_6287,N_6466);
nand U6572 (N_6572,N_6435,N_6475);
nor U6573 (N_6573,N_6360,N_6309);
xor U6574 (N_6574,N_6498,N_6433);
nand U6575 (N_6575,N_6485,N_6478);
nor U6576 (N_6576,N_6409,N_6470);
nor U6577 (N_6577,N_6374,N_6324);
or U6578 (N_6578,N_6496,N_6430);
nand U6579 (N_6579,N_6322,N_6268);
or U6580 (N_6580,N_6403,N_6344);
or U6581 (N_6581,N_6355,N_6277);
and U6582 (N_6582,N_6271,N_6456);
nor U6583 (N_6583,N_6264,N_6299);
nand U6584 (N_6584,N_6439,N_6377);
or U6585 (N_6585,N_6346,N_6307);
xor U6586 (N_6586,N_6394,N_6432);
or U6587 (N_6587,N_6364,N_6400);
xnor U6588 (N_6588,N_6488,N_6489);
nor U6589 (N_6589,N_6336,N_6342);
nand U6590 (N_6590,N_6306,N_6431);
xnor U6591 (N_6591,N_6482,N_6452);
or U6592 (N_6592,N_6442,N_6396);
or U6593 (N_6593,N_6301,N_6366);
xor U6594 (N_6594,N_6469,N_6449);
nand U6595 (N_6595,N_6298,N_6428);
and U6596 (N_6596,N_6319,N_6335);
nor U6597 (N_6597,N_6349,N_6398);
xnor U6598 (N_6598,N_6480,N_6481);
or U6599 (N_6599,N_6267,N_6352);
or U6600 (N_6600,N_6254,N_6429);
and U6601 (N_6601,N_6312,N_6443);
and U6602 (N_6602,N_6282,N_6280);
and U6603 (N_6603,N_6313,N_6365);
nor U6604 (N_6604,N_6262,N_6399);
xor U6605 (N_6605,N_6387,N_6381);
xor U6606 (N_6606,N_6441,N_6393);
or U6607 (N_6607,N_6250,N_6260);
xor U6608 (N_6608,N_6252,N_6256);
nor U6609 (N_6609,N_6285,N_6454);
and U6610 (N_6610,N_6383,N_6389);
nand U6611 (N_6611,N_6438,N_6318);
xnor U6612 (N_6612,N_6487,N_6477);
nor U6613 (N_6613,N_6286,N_6333);
or U6614 (N_6614,N_6263,N_6402);
nor U6615 (N_6615,N_6273,N_6295);
and U6616 (N_6616,N_6382,N_6363);
nand U6617 (N_6617,N_6378,N_6354);
and U6618 (N_6618,N_6290,N_6407);
nor U6619 (N_6619,N_6414,N_6465);
or U6620 (N_6620,N_6463,N_6297);
and U6621 (N_6621,N_6296,N_6325);
nand U6622 (N_6622,N_6259,N_6372);
xor U6623 (N_6623,N_6294,N_6314);
or U6624 (N_6624,N_6292,N_6464);
or U6625 (N_6625,N_6493,N_6273);
or U6626 (N_6626,N_6489,N_6318);
nor U6627 (N_6627,N_6325,N_6363);
or U6628 (N_6628,N_6402,N_6253);
and U6629 (N_6629,N_6491,N_6444);
nor U6630 (N_6630,N_6483,N_6497);
xor U6631 (N_6631,N_6301,N_6257);
or U6632 (N_6632,N_6365,N_6327);
nand U6633 (N_6633,N_6299,N_6459);
and U6634 (N_6634,N_6258,N_6426);
or U6635 (N_6635,N_6498,N_6334);
and U6636 (N_6636,N_6495,N_6381);
nand U6637 (N_6637,N_6451,N_6353);
nand U6638 (N_6638,N_6388,N_6297);
and U6639 (N_6639,N_6411,N_6294);
xnor U6640 (N_6640,N_6442,N_6278);
nand U6641 (N_6641,N_6485,N_6326);
and U6642 (N_6642,N_6327,N_6257);
nor U6643 (N_6643,N_6461,N_6456);
nor U6644 (N_6644,N_6413,N_6493);
xor U6645 (N_6645,N_6499,N_6288);
nor U6646 (N_6646,N_6480,N_6489);
nand U6647 (N_6647,N_6469,N_6424);
nand U6648 (N_6648,N_6298,N_6250);
or U6649 (N_6649,N_6422,N_6377);
and U6650 (N_6650,N_6305,N_6363);
xnor U6651 (N_6651,N_6442,N_6404);
and U6652 (N_6652,N_6452,N_6428);
nand U6653 (N_6653,N_6452,N_6445);
nor U6654 (N_6654,N_6498,N_6430);
nand U6655 (N_6655,N_6460,N_6303);
nand U6656 (N_6656,N_6398,N_6487);
xor U6657 (N_6657,N_6464,N_6442);
nor U6658 (N_6658,N_6293,N_6401);
or U6659 (N_6659,N_6349,N_6471);
xnor U6660 (N_6660,N_6254,N_6459);
and U6661 (N_6661,N_6441,N_6299);
nor U6662 (N_6662,N_6422,N_6440);
nor U6663 (N_6663,N_6481,N_6460);
nor U6664 (N_6664,N_6448,N_6273);
or U6665 (N_6665,N_6372,N_6268);
nand U6666 (N_6666,N_6434,N_6323);
nor U6667 (N_6667,N_6262,N_6452);
nand U6668 (N_6668,N_6313,N_6463);
xor U6669 (N_6669,N_6355,N_6314);
xnor U6670 (N_6670,N_6342,N_6273);
and U6671 (N_6671,N_6336,N_6474);
or U6672 (N_6672,N_6476,N_6324);
or U6673 (N_6673,N_6345,N_6398);
or U6674 (N_6674,N_6464,N_6307);
or U6675 (N_6675,N_6272,N_6417);
and U6676 (N_6676,N_6475,N_6428);
nor U6677 (N_6677,N_6276,N_6474);
or U6678 (N_6678,N_6320,N_6491);
or U6679 (N_6679,N_6370,N_6373);
nand U6680 (N_6680,N_6370,N_6264);
nand U6681 (N_6681,N_6305,N_6425);
nand U6682 (N_6682,N_6275,N_6480);
nand U6683 (N_6683,N_6306,N_6395);
nand U6684 (N_6684,N_6361,N_6277);
and U6685 (N_6685,N_6490,N_6287);
xor U6686 (N_6686,N_6382,N_6451);
or U6687 (N_6687,N_6274,N_6494);
xnor U6688 (N_6688,N_6384,N_6450);
nand U6689 (N_6689,N_6397,N_6389);
and U6690 (N_6690,N_6479,N_6415);
nor U6691 (N_6691,N_6303,N_6474);
xnor U6692 (N_6692,N_6384,N_6442);
and U6693 (N_6693,N_6331,N_6259);
and U6694 (N_6694,N_6299,N_6399);
and U6695 (N_6695,N_6456,N_6382);
xnor U6696 (N_6696,N_6279,N_6352);
nor U6697 (N_6697,N_6329,N_6263);
nand U6698 (N_6698,N_6362,N_6303);
and U6699 (N_6699,N_6266,N_6389);
and U6700 (N_6700,N_6295,N_6259);
xor U6701 (N_6701,N_6289,N_6250);
and U6702 (N_6702,N_6470,N_6328);
nor U6703 (N_6703,N_6267,N_6394);
or U6704 (N_6704,N_6388,N_6453);
and U6705 (N_6705,N_6466,N_6444);
or U6706 (N_6706,N_6291,N_6369);
nor U6707 (N_6707,N_6335,N_6494);
nor U6708 (N_6708,N_6423,N_6388);
or U6709 (N_6709,N_6362,N_6446);
nand U6710 (N_6710,N_6481,N_6305);
or U6711 (N_6711,N_6434,N_6440);
or U6712 (N_6712,N_6445,N_6399);
and U6713 (N_6713,N_6360,N_6341);
xor U6714 (N_6714,N_6270,N_6488);
xor U6715 (N_6715,N_6443,N_6437);
nand U6716 (N_6716,N_6339,N_6463);
nor U6717 (N_6717,N_6400,N_6425);
nand U6718 (N_6718,N_6283,N_6359);
nand U6719 (N_6719,N_6365,N_6309);
or U6720 (N_6720,N_6338,N_6360);
nand U6721 (N_6721,N_6302,N_6401);
and U6722 (N_6722,N_6301,N_6452);
and U6723 (N_6723,N_6352,N_6325);
or U6724 (N_6724,N_6302,N_6417);
nor U6725 (N_6725,N_6465,N_6340);
or U6726 (N_6726,N_6369,N_6374);
or U6727 (N_6727,N_6418,N_6318);
xnor U6728 (N_6728,N_6272,N_6438);
xnor U6729 (N_6729,N_6254,N_6345);
and U6730 (N_6730,N_6329,N_6253);
nor U6731 (N_6731,N_6337,N_6372);
nor U6732 (N_6732,N_6396,N_6498);
or U6733 (N_6733,N_6336,N_6482);
xnor U6734 (N_6734,N_6268,N_6346);
or U6735 (N_6735,N_6334,N_6313);
and U6736 (N_6736,N_6397,N_6377);
or U6737 (N_6737,N_6497,N_6460);
nor U6738 (N_6738,N_6474,N_6282);
or U6739 (N_6739,N_6292,N_6408);
nor U6740 (N_6740,N_6265,N_6383);
nor U6741 (N_6741,N_6250,N_6252);
or U6742 (N_6742,N_6372,N_6409);
nand U6743 (N_6743,N_6416,N_6428);
or U6744 (N_6744,N_6329,N_6317);
nand U6745 (N_6745,N_6360,N_6315);
or U6746 (N_6746,N_6366,N_6373);
xor U6747 (N_6747,N_6495,N_6483);
xnor U6748 (N_6748,N_6439,N_6349);
xnor U6749 (N_6749,N_6306,N_6250);
nand U6750 (N_6750,N_6587,N_6676);
xnor U6751 (N_6751,N_6720,N_6674);
or U6752 (N_6752,N_6571,N_6748);
and U6753 (N_6753,N_6539,N_6522);
nor U6754 (N_6754,N_6541,N_6591);
nor U6755 (N_6755,N_6697,N_6655);
nor U6756 (N_6756,N_6555,N_6511);
or U6757 (N_6757,N_6521,N_6683);
or U6758 (N_6758,N_6735,N_6698);
xor U6759 (N_6759,N_6560,N_6611);
nand U6760 (N_6760,N_6726,N_6542);
or U6761 (N_6761,N_6667,N_6614);
or U6762 (N_6762,N_6656,N_6669);
nand U6763 (N_6763,N_6524,N_6512);
and U6764 (N_6764,N_6604,N_6568);
and U6765 (N_6765,N_6585,N_6581);
xnor U6766 (N_6766,N_6579,N_6594);
or U6767 (N_6767,N_6742,N_6505);
nor U6768 (N_6768,N_6686,N_6537);
nor U6769 (N_6769,N_6724,N_6596);
nor U6770 (N_6770,N_6658,N_6528);
or U6771 (N_6771,N_6730,N_6629);
xor U6772 (N_6772,N_6688,N_6651);
or U6773 (N_6773,N_6603,N_6507);
and U6774 (N_6774,N_6544,N_6520);
and U6775 (N_6775,N_6561,N_6642);
xor U6776 (N_6776,N_6586,N_6734);
and U6777 (N_6777,N_6733,N_6725);
nor U6778 (N_6778,N_6705,N_6648);
or U6779 (N_6779,N_6677,N_6646);
or U6780 (N_6780,N_6740,N_6540);
nand U6781 (N_6781,N_6523,N_6535);
xnor U6782 (N_6782,N_6639,N_6550);
and U6783 (N_6783,N_6504,N_6506);
nand U6784 (N_6784,N_6700,N_6517);
nor U6785 (N_6785,N_6678,N_6563);
nor U6786 (N_6786,N_6617,N_6671);
nand U6787 (N_6787,N_6577,N_6737);
nand U6788 (N_6788,N_6682,N_6628);
and U6789 (N_6789,N_6710,N_6619);
or U6790 (N_6790,N_6592,N_6572);
and U6791 (N_6791,N_6680,N_6547);
and U6792 (N_6792,N_6690,N_6719);
xor U6793 (N_6793,N_6643,N_6721);
or U6794 (N_6794,N_6749,N_6723);
xor U6795 (N_6795,N_6534,N_6549);
nand U6796 (N_6796,N_6607,N_6708);
nand U6797 (N_6797,N_6653,N_6746);
nor U6798 (N_6798,N_6613,N_6546);
xnor U6799 (N_6799,N_6608,N_6558);
xnor U6800 (N_6800,N_6625,N_6557);
or U6801 (N_6801,N_6716,N_6576);
nor U6802 (N_6802,N_6574,N_6510);
nand U6803 (N_6803,N_6623,N_6747);
xnor U6804 (N_6804,N_6508,N_6519);
xor U6805 (N_6805,N_6564,N_6500);
nand U6806 (N_6806,N_6631,N_6538);
nand U6807 (N_6807,N_6530,N_6638);
and U6808 (N_6808,N_6715,N_6627);
nand U6809 (N_6809,N_6703,N_6728);
xor U6810 (N_6810,N_6736,N_6531);
and U6811 (N_6811,N_6729,N_6569);
or U6812 (N_6812,N_6717,N_6684);
or U6813 (N_6813,N_6709,N_6652);
or U6814 (N_6814,N_6565,N_6552);
or U6815 (N_6815,N_6609,N_6695);
and U6816 (N_6816,N_6696,N_6647);
nand U6817 (N_6817,N_6559,N_6529);
nand U6818 (N_6818,N_6692,N_6584);
or U6819 (N_6819,N_6553,N_6636);
nor U6820 (N_6820,N_6722,N_6621);
nand U6821 (N_6821,N_6616,N_6713);
xor U6822 (N_6822,N_6578,N_6668);
nand U6823 (N_6823,N_6699,N_6644);
nor U6824 (N_6824,N_6583,N_6641);
nor U6825 (N_6825,N_6650,N_6707);
nand U6826 (N_6826,N_6660,N_6687);
and U6827 (N_6827,N_6675,N_6597);
and U6828 (N_6828,N_6704,N_6595);
xor U6829 (N_6829,N_6706,N_6635);
nor U6830 (N_6830,N_6731,N_6543);
xor U6831 (N_6831,N_6554,N_6526);
nand U6832 (N_6832,N_6665,N_6702);
and U6833 (N_6833,N_6527,N_6714);
and U6834 (N_6834,N_6501,N_6634);
or U6835 (N_6835,N_6610,N_6691);
or U6836 (N_6836,N_6605,N_6514);
and U6837 (N_6837,N_6502,N_6633);
and U6838 (N_6838,N_6666,N_6602);
nor U6839 (N_6839,N_6516,N_6532);
or U6840 (N_6840,N_6640,N_6590);
xnor U6841 (N_6841,N_6601,N_6738);
xor U6842 (N_6842,N_6575,N_6562);
nor U6843 (N_6843,N_6661,N_6657);
nand U6844 (N_6844,N_6600,N_6548);
nor U6845 (N_6845,N_6518,N_6712);
and U6846 (N_6846,N_6679,N_6622);
nor U6847 (N_6847,N_6567,N_6566);
or U6848 (N_6848,N_6632,N_6582);
and U6849 (N_6849,N_6689,N_6670);
or U6850 (N_6850,N_6525,N_6626);
and U6851 (N_6851,N_6615,N_6630);
nor U6852 (N_6852,N_6649,N_6588);
or U6853 (N_6853,N_6744,N_6533);
nand U6854 (N_6854,N_6741,N_6645);
nor U6855 (N_6855,N_6593,N_6745);
nor U6856 (N_6856,N_6606,N_6673);
or U6857 (N_6857,N_6551,N_6718);
nand U6858 (N_6858,N_6727,N_6599);
or U6859 (N_6859,N_6598,N_6503);
nor U6860 (N_6860,N_6681,N_6589);
or U6861 (N_6861,N_6637,N_6570);
nor U6862 (N_6862,N_6513,N_6672);
and U6863 (N_6863,N_6685,N_6663);
xor U6864 (N_6864,N_6694,N_6739);
and U6865 (N_6865,N_6620,N_6509);
and U6866 (N_6866,N_6693,N_6743);
nor U6867 (N_6867,N_6659,N_6536);
xor U6868 (N_6868,N_6612,N_6701);
xnor U6869 (N_6869,N_6732,N_6545);
xor U6870 (N_6870,N_6573,N_6664);
nand U6871 (N_6871,N_6624,N_6580);
nor U6872 (N_6872,N_6711,N_6515);
or U6873 (N_6873,N_6556,N_6662);
nand U6874 (N_6874,N_6654,N_6618);
xor U6875 (N_6875,N_6747,N_6690);
nor U6876 (N_6876,N_6603,N_6708);
nor U6877 (N_6877,N_6502,N_6509);
or U6878 (N_6878,N_6570,N_6745);
or U6879 (N_6879,N_6735,N_6749);
and U6880 (N_6880,N_6552,N_6657);
and U6881 (N_6881,N_6649,N_6517);
xor U6882 (N_6882,N_6693,N_6667);
nor U6883 (N_6883,N_6748,N_6612);
xor U6884 (N_6884,N_6656,N_6704);
nor U6885 (N_6885,N_6519,N_6559);
and U6886 (N_6886,N_6570,N_6723);
xor U6887 (N_6887,N_6583,N_6684);
nor U6888 (N_6888,N_6522,N_6628);
nand U6889 (N_6889,N_6661,N_6588);
nand U6890 (N_6890,N_6557,N_6617);
nand U6891 (N_6891,N_6596,N_6529);
nor U6892 (N_6892,N_6516,N_6708);
xnor U6893 (N_6893,N_6679,N_6550);
and U6894 (N_6894,N_6521,N_6706);
nand U6895 (N_6895,N_6511,N_6716);
and U6896 (N_6896,N_6582,N_6658);
nand U6897 (N_6897,N_6517,N_6625);
xor U6898 (N_6898,N_6651,N_6563);
or U6899 (N_6899,N_6731,N_6645);
or U6900 (N_6900,N_6731,N_6728);
or U6901 (N_6901,N_6521,N_6501);
nor U6902 (N_6902,N_6630,N_6662);
or U6903 (N_6903,N_6660,N_6595);
xnor U6904 (N_6904,N_6713,N_6742);
nand U6905 (N_6905,N_6643,N_6595);
xor U6906 (N_6906,N_6730,N_6521);
nor U6907 (N_6907,N_6726,N_6734);
xor U6908 (N_6908,N_6700,N_6719);
nor U6909 (N_6909,N_6527,N_6505);
nor U6910 (N_6910,N_6550,N_6575);
or U6911 (N_6911,N_6656,N_6702);
nand U6912 (N_6912,N_6548,N_6703);
nand U6913 (N_6913,N_6515,N_6661);
nor U6914 (N_6914,N_6679,N_6594);
or U6915 (N_6915,N_6633,N_6738);
and U6916 (N_6916,N_6581,N_6526);
or U6917 (N_6917,N_6541,N_6678);
nand U6918 (N_6918,N_6590,N_6500);
and U6919 (N_6919,N_6613,N_6521);
nor U6920 (N_6920,N_6663,N_6608);
or U6921 (N_6921,N_6709,N_6590);
nor U6922 (N_6922,N_6724,N_6538);
and U6923 (N_6923,N_6621,N_6630);
xnor U6924 (N_6924,N_6720,N_6614);
xnor U6925 (N_6925,N_6700,N_6661);
or U6926 (N_6926,N_6576,N_6591);
xor U6927 (N_6927,N_6559,N_6605);
and U6928 (N_6928,N_6648,N_6655);
xor U6929 (N_6929,N_6584,N_6696);
or U6930 (N_6930,N_6518,N_6749);
nor U6931 (N_6931,N_6701,N_6589);
xor U6932 (N_6932,N_6593,N_6742);
nand U6933 (N_6933,N_6631,N_6590);
xor U6934 (N_6934,N_6562,N_6732);
or U6935 (N_6935,N_6568,N_6556);
nor U6936 (N_6936,N_6554,N_6640);
xor U6937 (N_6937,N_6510,N_6511);
nand U6938 (N_6938,N_6722,N_6578);
xor U6939 (N_6939,N_6748,N_6594);
xnor U6940 (N_6940,N_6574,N_6590);
or U6941 (N_6941,N_6609,N_6716);
or U6942 (N_6942,N_6627,N_6631);
nor U6943 (N_6943,N_6579,N_6736);
nor U6944 (N_6944,N_6532,N_6645);
xnor U6945 (N_6945,N_6615,N_6610);
and U6946 (N_6946,N_6521,N_6698);
nand U6947 (N_6947,N_6675,N_6741);
or U6948 (N_6948,N_6607,N_6573);
and U6949 (N_6949,N_6505,N_6528);
nor U6950 (N_6950,N_6688,N_6572);
nand U6951 (N_6951,N_6655,N_6661);
xnor U6952 (N_6952,N_6678,N_6510);
xnor U6953 (N_6953,N_6533,N_6581);
xnor U6954 (N_6954,N_6743,N_6716);
or U6955 (N_6955,N_6577,N_6663);
nand U6956 (N_6956,N_6515,N_6541);
xor U6957 (N_6957,N_6546,N_6588);
nor U6958 (N_6958,N_6645,N_6570);
xnor U6959 (N_6959,N_6585,N_6711);
or U6960 (N_6960,N_6636,N_6584);
and U6961 (N_6961,N_6661,N_6508);
or U6962 (N_6962,N_6704,N_6653);
xnor U6963 (N_6963,N_6514,N_6691);
or U6964 (N_6964,N_6719,N_6671);
and U6965 (N_6965,N_6662,N_6599);
or U6966 (N_6966,N_6641,N_6726);
and U6967 (N_6967,N_6650,N_6593);
xnor U6968 (N_6968,N_6537,N_6731);
xnor U6969 (N_6969,N_6580,N_6566);
or U6970 (N_6970,N_6633,N_6504);
and U6971 (N_6971,N_6558,N_6658);
xor U6972 (N_6972,N_6601,N_6699);
nand U6973 (N_6973,N_6621,N_6700);
or U6974 (N_6974,N_6570,N_6587);
nand U6975 (N_6975,N_6616,N_6509);
nand U6976 (N_6976,N_6717,N_6665);
nand U6977 (N_6977,N_6582,N_6542);
or U6978 (N_6978,N_6746,N_6633);
nand U6979 (N_6979,N_6663,N_6740);
and U6980 (N_6980,N_6699,N_6713);
nor U6981 (N_6981,N_6722,N_6558);
xnor U6982 (N_6982,N_6549,N_6513);
xnor U6983 (N_6983,N_6554,N_6599);
or U6984 (N_6984,N_6529,N_6744);
and U6985 (N_6985,N_6673,N_6538);
xor U6986 (N_6986,N_6512,N_6502);
or U6987 (N_6987,N_6514,N_6626);
nand U6988 (N_6988,N_6734,N_6608);
nor U6989 (N_6989,N_6572,N_6699);
xnor U6990 (N_6990,N_6627,N_6701);
nor U6991 (N_6991,N_6696,N_6635);
nor U6992 (N_6992,N_6589,N_6646);
nand U6993 (N_6993,N_6687,N_6603);
xor U6994 (N_6994,N_6530,N_6713);
xor U6995 (N_6995,N_6507,N_6741);
xnor U6996 (N_6996,N_6517,N_6533);
nor U6997 (N_6997,N_6586,N_6603);
nor U6998 (N_6998,N_6738,N_6509);
and U6999 (N_6999,N_6706,N_6697);
and U7000 (N_7000,N_6910,N_6958);
and U7001 (N_7001,N_6920,N_6783);
xor U7002 (N_7002,N_6908,N_6784);
nor U7003 (N_7003,N_6935,N_6772);
xor U7004 (N_7004,N_6871,N_6954);
nand U7005 (N_7005,N_6970,N_6808);
xnor U7006 (N_7006,N_6893,N_6775);
nor U7007 (N_7007,N_6869,N_6939);
or U7008 (N_7008,N_6953,N_6926);
nand U7009 (N_7009,N_6999,N_6917);
nand U7010 (N_7010,N_6802,N_6795);
and U7011 (N_7011,N_6858,N_6866);
and U7012 (N_7012,N_6750,N_6986);
nor U7013 (N_7013,N_6764,N_6888);
and U7014 (N_7014,N_6900,N_6812);
nand U7015 (N_7015,N_6885,N_6853);
nor U7016 (N_7016,N_6843,N_6805);
xnor U7017 (N_7017,N_6849,N_6797);
nor U7018 (N_7018,N_6791,N_6967);
or U7019 (N_7019,N_6835,N_6988);
nand U7020 (N_7020,N_6921,N_6989);
xnor U7021 (N_7021,N_6878,N_6886);
xor U7022 (N_7022,N_6879,N_6841);
xnor U7023 (N_7023,N_6934,N_6994);
nor U7024 (N_7024,N_6862,N_6963);
nor U7025 (N_7025,N_6813,N_6826);
nand U7026 (N_7026,N_6766,N_6777);
nor U7027 (N_7027,N_6758,N_6966);
or U7028 (N_7028,N_6972,N_6923);
xor U7029 (N_7029,N_6851,N_6798);
and U7030 (N_7030,N_6832,N_6883);
nor U7031 (N_7031,N_6976,N_6768);
nand U7032 (N_7032,N_6864,N_6760);
xnor U7033 (N_7033,N_6933,N_6937);
or U7034 (N_7034,N_6904,N_6997);
xnor U7035 (N_7035,N_6973,N_6932);
and U7036 (N_7036,N_6964,N_6844);
xnor U7037 (N_7037,N_6957,N_6815);
xor U7038 (N_7038,N_6992,N_6831);
and U7039 (N_7039,N_6762,N_6945);
and U7040 (N_7040,N_6870,N_6996);
or U7041 (N_7041,N_6820,N_6956);
nor U7042 (N_7042,N_6856,N_6852);
nand U7043 (N_7043,N_6756,N_6889);
nand U7044 (N_7044,N_6974,N_6860);
or U7045 (N_7045,N_6824,N_6773);
nand U7046 (N_7046,N_6821,N_6898);
and U7047 (N_7047,N_6882,N_6948);
nor U7048 (N_7048,N_6874,N_6848);
or U7049 (N_7049,N_6891,N_6785);
nand U7050 (N_7050,N_6761,N_6838);
or U7051 (N_7051,N_6823,N_6825);
or U7052 (N_7052,N_6982,N_6919);
nor U7053 (N_7053,N_6828,N_6909);
or U7054 (N_7054,N_6924,N_6985);
xor U7055 (N_7055,N_6936,N_6940);
xnor U7056 (N_7056,N_6961,N_6931);
xnor U7057 (N_7057,N_6959,N_6837);
or U7058 (N_7058,N_6819,N_6987);
nor U7059 (N_7059,N_6839,N_6788);
nand U7060 (N_7060,N_6751,N_6941);
or U7061 (N_7061,N_6875,N_6930);
or U7062 (N_7062,N_6814,N_6822);
or U7063 (N_7063,N_6840,N_6955);
nand U7064 (N_7064,N_6859,N_6770);
xor U7065 (N_7065,N_6884,N_6833);
and U7066 (N_7066,N_6807,N_6857);
xor U7067 (N_7067,N_6845,N_6984);
or U7068 (N_7068,N_6971,N_6975);
nand U7069 (N_7069,N_6754,N_6960);
nand U7070 (N_7070,N_6951,N_6901);
or U7071 (N_7071,N_6755,N_6769);
or U7072 (N_7072,N_6969,N_6850);
nand U7073 (N_7073,N_6816,N_6804);
or U7074 (N_7074,N_6836,N_6776);
or U7075 (N_7075,N_6890,N_6896);
xor U7076 (N_7076,N_6803,N_6922);
xnor U7077 (N_7077,N_6993,N_6846);
nor U7078 (N_7078,N_6911,N_6944);
nor U7079 (N_7079,N_6752,N_6962);
or U7080 (N_7080,N_6765,N_6912);
nor U7081 (N_7081,N_6927,N_6790);
nand U7082 (N_7082,N_6905,N_6757);
nand U7083 (N_7083,N_6779,N_6918);
xnor U7084 (N_7084,N_6753,N_6983);
nand U7085 (N_7085,N_6865,N_6925);
or U7086 (N_7086,N_6800,N_6782);
xor U7087 (N_7087,N_6799,N_6977);
nor U7088 (N_7088,N_6834,N_6899);
nor U7089 (N_7089,N_6915,N_6965);
nor U7090 (N_7090,N_6950,N_6842);
xnor U7091 (N_7091,N_6902,N_6952);
and U7092 (N_7092,N_6979,N_6781);
or U7093 (N_7093,N_6947,N_6981);
and U7094 (N_7094,N_6867,N_6787);
and U7095 (N_7095,N_6903,N_6863);
and U7096 (N_7096,N_6907,N_6827);
xor U7097 (N_7097,N_6792,N_6786);
xnor U7098 (N_7098,N_6793,N_6771);
nand U7099 (N_7099,N_6811,N_6817);
or U7100 (N_7100,N_6990,N_6906);
nor U7101 (N_7101,N_6914,N_6929);
nand U7102 (N_7102,N_6855,N_6794);
and U7103 (N_7103,N_6818,N_6778);
nand U7104 (N_7104,N_6942,N_6991);
or U7105 (N_7105,N_6916,N_6913);
xor U7106 (N_7106,N_6767,N_6763);
nand U7107 (N_7107,N_6928,N_6774);
nor U7108 (N_7108,N_6895,N_6892);
or U7109 (N_7109,N_6995,N_6759);
nand U7110 (N_7110,N_6868,N_6980);
or U7111 (N_7111,N_6810,N_6887);
or U7112 (N_7112,N_6830,N_6806);
nor U7113 (N_7113,N_6861,N_6978);
xnor U7114 (N_7114,N_6897,N_6881);
or U7115 (N_7115,N_6872,N_6946);
and U7116 (N_7116,N_6943,N_6880);
or U7117 (N_7117,N_6998,N_6938);
xnor U7118 (N_7118,N_6796,N_6854);
and U7119 (N_7119,N_6809,N_6877);
xor U7120 (N_7120,N_6949,N_6894);
nand U7121 (N_7121,N_6789,N_6829);
nand U7122 (N_7122,N_6780,N_6876);
or U7123 (N_7123,N_6968,N_6801);
and U7124 (N_7124,N_6873,N_6847);
or U7125 (N_7125,N_6834,N_6859);
nor U7126 (N_7126,N_6765,N_6837);
or U7127 (N_7127,N_6951,N_6941);
xor U7128 (N_7128,N_6898,N_6789);
and U7129 (N_7129,N_6892,N_6925);
nand U7130 (N_7130,N_6838,N_6807);
and U7131 (N_7131,N_6834,N_6867);
and U7132 (N_7132,N_6939,N_6999);
and U7133 (N_7133,N_6855,N_6771);
or U7134 (N_7134,N_6979,N_6806);
nor U7135 (N_7135,N_6961,N_6886);
nand U7136 (N_7136,N_6846,N_6770);
xnor U7137 (N_7137,N_6896,N_6825);
xor U7138 (N_7138,N_6965,N_6945);
and U7139 (N_7139,N_6936,N_6781);
and U7140 (N_7140,N_6985,N_6799);
or U7141 (N_7141,N_6815,N_6755);
nor U7142 (N_7142,N_6793,N_6835);
nor U7143 (N_7143,N_6916,N_6852);
nand U7144 (N_7144,N_6996,N_6887);
and U7145 (N_7145,N_6955,N_6822);
or U7146 (N_7146,N_6818,N_6865);
xor U7147 (N_7147,N_6820,N_6977);
or U7148 (N_7148,N_6922,N_6785);
nand U7149 (N_7149,N_6816,N_6862);
or U7150 (N_7150,N_6838,N_6998);
xor U7151 (N_7151,N_6856,N_6910);
and U7152 (N_7152,N_6840,N_6898);
nand U7153 (N_7153,N_6836,N_6976);
or U7154 (N_7154,N_6970,N_6978);
nor U7155 (N_7155,N_6895,N_6917);
nand U7156 (N_7156,N_6907,N_6934);
nor U7157 (N_7157,N_6921,N_6911);
and U7158 (N_7158,N_6787,N_6911);
and U7159 (N_7159,N_6796,N_6787);
and U7160 (N_7160,N_6930,N_6764);
nor U7161 (N_7161,N_6968,N_6950);
xnor U7162 (N_7162,N_6759,N_6792);
nor U7163 (N_7163,N_6857,N_6785);
nor U7164 (N_7164,N_6869,N_6911);
and U7165 (N_7165,N_6810,N_6933);
xnor U7166 (N_7166,N_6866,N_6959);
nand U7167 (N_7167,N_6976,N_6911);
nor U7168 (N_7168,N_6795,N_6912);
nand U7169 (N_7169,N_6845,N_6831);
nand U7170 (N_7170,N_6881,N_6752);
nand U7171 (N_7171,N_6867,N_6971);
and U7172 (N_7172,N_6994,N_6890);
nand U7173 (N_7173,N_6905,N_6875);
or U7174 (N_7174,N_6793,N_6981);
nand U7175 (N_7175,N_6901,N_6974);
nor U7176 (N_7176,N_6917,N_6846);
xor U7177 (N_7177,N_6788,N_6929);
and U7178 (N_7178,N_6860,N_6859);
nor U7179 (N_7179,N_6758,N_6848);
xor U7180 (N_7180,N_6932,N_6981);
and U7181 (N_7181,N_6985,N_6836);
nor U7182 (N_7182,N_6924,N_6975);
nor U7183 (N_7183,N_6998,N_6786);
and U7184 (N_7184,N_6909,N_6850);
nor U7185 (N_7185,N_6916,N_6960);
or U7186 (N_7186,N_6832,N_6794);
nor U7187 (N_7187,N_6916,N_6765);
nand U7188 (N_7188,N_6829,N_6917);
or U7189 (N_7189,N_6785,N_6980);
nor U7190 (N_7190,N_6824,N_6855);
and U7191 (N_7191,N_6772,N_6912);
or U7192 (N_7192,N_6764,N_6786);
nand U7193 (N_7193,N_6794,N_6859);
nand U7194 (N_7194,N_6793,N_6916);
nand U7195 (N_7195,N_6913,N_6934);
xor U7196 (N_7196,N_6764,N_6893);
nor U7197 (N_7197,N_6825,N_6966);
or U7198 (N_7198,N_6872,N_6764);
nand U7199 (N_7199,N_6869,N_6775);
nand U7200 (N_7200,N_6853,N_6770);
nor U7201 (N_7201,N_6843,N_6926);
or U7202 (N_7202,N_6945,N_6967);
nor U7203 (N_7203,N_6758,N_6894);
or U7204 (N_7204,N_6987,N_6783);
nand U7205 (N_7205,N_6925,N_6778);
nand U7206 (N_7206,N_6969,N_6772);
nor U7207 (N_7207,N_6813,N_6912);
and U7208 (N_7208,N_6844,N_6783);
nor U7209 (N_7209,N_6842,N_6943);
or U7210 (N_7210,N_6893,N_6832);
or U7211 (N_7211,N_6888,N_6842);
and U7212 (N_7212,N_6859,N_6787);
and U7213 (N_7213,N_6868,N_6879);
nand U7214 (N_7214,N_6977,N_6942);
and U7215 (N_7215,N_6792,N_6761);
nor U7216 (N_7216,N_6882,N_6979);
nand U7217 (N_7217,N_6827,N_6931);
nor U7218 (N_7218,N_6871,N_6808);
nand U7219 (N_7219,N_6970,N_6811);
nand U7220 (N_7220,N_6890,N_6796);
xnor U7221 (N_7221,N_6865,N_6929);
and U7222 (N_7222,N_6790,N_6916);
nor U7223 (N_7223,N_6774,N_6865);
and U7224 (N_7224,N_6997,N_6760);
xor U7225 (N_7225,N_6771,N_6903);
xnor U7226 (N_7226,N_6920,N_6758);
xnor U7227 (N_7227,N_6961,N_6893);
or U7228 (N_7228,N_6955,N_6891);
and U7229 (N_7229,N_6980,N_6797);
or U7230 (N_7230,N_6817,N_6764);
or U7231 (N_7231,N_6876,N_6806);
or U7232 (N_7232,N_6953,N_6898);
and U7233 (N_7233,N_6853,N_6850);
nor U7234 (N_7234,N_6842,N_6920);
and U7235 (N_7235,N_6810,N_6787);
and U7236 (N_7236,N_6779,N_6884);
xnor U7237 (N_7237,N_6940,N_6839);
or U7238 (N_7238,N_6813,N_6875);
and U7239 (N_7239,N_6778,N_6809);
nor U7240 (N_7240,N_6939,N_6819);
and U7241 (N_7241,N_6797,N_6861);
nor U7242 (N_7242,N_6825,N_6894);
nand U7243 (N_7243,N_6906,N_6955);
nor U7244 (N_7244,N_6866,N_6800);
xnor U7245 (N_7245,N_6859,N_6987);
or U7246 (N_7246,N_6857,N_6887);
and U7247 (N_7247,N_6931,N_6954);
nand U7248 (N_7248,N_6873,N_6875);
and U7249 (N_7249,N_6859,N_6999);
xor U7250 (N_7250,N_7095,N_7196);
nor U7251 (N_7251,N_7060,N_7072);
xor U7252 (N_7252,N_7200,N_7046);
nand U7253 (N_7253,N_7164,N_7030);
and U7254 (N_7254,N_7103,N_7153);
xor U7255 (N_7255,N_7013,N_7109);
xor U7256 (N_7256,N_7117,N_7105);
nand U7257 (N_7257,N_7067,N_7217);
xor U7258 (N_7258,N_7209,N_7182);
xnor U7259 (N_7259,N_7215,N_7239);
nor U7260 (N_7260,N_7057,N_7144);
or U7261 (N_7261,N_7143,N_7224);
and U7262 (N_7262,N_7044,N_7045);
nor U7263 (N_7263,N_7027,N_7149);
and U7264 (N_7264,N_7228,N_7134);
nand U7265 (N_7265,N_7058,N_7246);
nand U7266 (N_7266,N_7194,N_7053);
or U7267 (N_7267,N_7146,N_7202);
nand U7268 (N_7268,N_7042,N_7245);
nor U7269 (N_7269,N_7137,N_7176);
nand U7270 (N_7270,N_7115,N_7133);
and U7271 (N_7271,N_7000,N_7163);
and U7272 (N_7272,N_7210,N_7028);
nand U7273 (N_7273,N_7010,N_7162);
nor U7274 (N_7274,N_7238,N_7090);
xor U7275 (N_7275,N_7247,N_7086);
nand U7276 (N_7276,N_7119,N_7054);
xnor U7277 (N_7277,N_7066,N_7130);
or U7278 (N_7278,N_7125,N_7032);
or U7279 (N_7279,N_7197,N_7244);
and U7280 (N_7280,N_7108,N_7055);
or U7281 (N_7281,N_7173,N_7212);
nor U7282 (N_7282,N_7107,N_7026);
or U7283 (N_7283,N_7225,N_7183);
or U7284 (N_7284,N_7214,N_7074);
and U7285 (N_7285,N_7004,N_7236);
and U7286 (N_7286,N_7089,N_7123);
xnor U7287 (N_7287,N_7240,N_7015);
nor U7288 (N_7288,N_7036,N_7181);
or U7289 (N_7289,N_7094,N_7129);
and U7290 (N_7290,N_7088,N_7160);
or U7291 (N_7291,N_7069,N_7185);
or U7292 (N_7292,N_7116,N_7120);
nor U7293 (N_7293,N_7077,N_7121);
nor U7294 (N_7294,N_7114,N_7083);
and U7295 (N_7295,N_7049,N_7039);
and U7296 (N_7296,N_7193,N_7171);
xor U7297 (N_7297,N_7242,N_7081);
or U7298 (N_7298,N_7172,N_7213);
xnor U7299 (N_7299,N_7093,N_7061);
and U7300 (N_7300,N_7111,N_7034);
nand U7301 (N_7301,N_7110,N_7147);
nand U7302 (N_7302,N_7249,N_7248);
xor U7303 (N_7303,N_7082,N_7007);
nand U7304 (N_7304,N_7070,N_7140);
or U7305 (N_7305,N_7131,N_7220);
and U7306 (N_7306,N_7189,N_7047);
and U7307 (N_7307,N_7018,N_7159);
and U7308 (N_7308,N_7006,N_7218);
xnor U7309 (N_7309,N_7161,N_7051);
or U7310 (N_7310,N_7241,N_7195);
xnor U7311 (N_7311,N_7087,N_7166);
nor U7312 (N_7312,N_7017,N_7151);
nand U7313 (N_7313,N_7226,N_7184);
xor U7314 (N_7314,N_7056,N_7048);
nand U7315 (N_7315,N_7100,N_7025);
and U7316 (N_7316,N_7136,N_7127);
or U7317 (N_7317,N_7216,N_7063);
xor U7318 (N_7318,N_7002,N_7158);
or U7319 (N_7319,N_7098,N_7050);
or U7320 (N_7320,N_7168,N_7229);
nor U7321 (N_7321,N_7179,N_7085);
or U7322 (N_7322,N_7118,N_7235);
xnor U7323 (N_7323,N_7169,N_7174);
nand U7324 (N_7324,N_7008,N_7033);
xor U7325 (N_7325,N_7198,N_7142);
xor U7326 (N_7326,N_7165,N_7078);
nor U7327 (N_7327,N_7029,N_7122);
nand U7328 (N_7328,N_7068,N_7112);
xor U7329 (N_7329,N_7148,N_7052);
xnor U7330 (N_7330,N_7124,N_7170);
and U7331 (N_7331,N_7227,N_7191);
nor U7332 (N_7332,N_7208,N_7156);
xnor U7333 (N_7333,N_7001,N_7099);
or U7334 (N_7334,N_7155,N_7237);
nand U7335 (N_7335,N_7073,N_7186);
and U7336 (N_7336,N_7097,N_7092);
nor U7337 (N_7337,N_7175,N_7222);
xor U7338 (N_7338,N_7150,N_7014);
and U7339 (N_7339,N_7177,N_7201);
and U7340 (N_7340,N_7205,N_7113);
and U7341 (N_7341,N_7021,N_7234);
and U7342 (N_7342,N_7012,N_7091);
nor U7343 (N_7343,N_7106,N_7101);
nand U7344 (N_7344,N_7138,N_7104);
and U7345 (N_7345,N_7003,N_7035);
xnor U7346 (N_7346,N_7080,N_7231);
nor U7347 (N_7347,N_7232,N_7145);
xor U7348 (N_7348,N_7178,N_7059);
or U7349 (N_7349,N_7141,N_7011);
xor U7350 (N_7350,N_7199,N_7024);
nor U7351 (N_7351,N_7204,N_7243);
nand U7352 (N_7352,N_7223,N_7132);
or U7353 (N_7353,N_7020,N_7190);
or U7354 (N_7354,N_7219,N_7043);
and U7355 (N_7355,N_7009,N_7016);
or U7356 (N_7356,N_7102,N_7152);
and U7357 (N_7357,N_7037,N_7192);
nor U7358 (N_7358,N_7207,N_7188);
nor U7359 (N_7359,N_7031,N_7221);
nand U7360 (N_7360,N_7211,N_7128);
nor U7361 (N_7361,N_7203,N_7038);
nand U7362 (N_7362,N_7076,N_7096);
xnor U7363 (N_7363,N_7019,N_7135);
or U7364 (N_7364,N_7233,N_7139);
nor U7365 (N_7365,N_7180,N_7167);
nand U7366 (N_7366,N_7230,N_7126);
and U7367 (N_7367,N_7084,N_7022);
and U7368 (N_7368,N_7040,N_7065);
nand U7369 (N_7369,N_7075,N_7154);
xnor U7370 (N_7370,N_7041,N_7071);
xor U7371 (N_7371,N_7062,N_7064);
and U7372 (N_7372,N_7079,N_7157);
and U7373 (N_7373,N_7206,N_7005);
and U7374 (N_7374,N_7187,N_7023);
and U7375 (N_7375,N_7117,N_7101);
nor U7376 (N_7376,N_7012,N_7048);
nand U7377 (N_7377,N_7085,N_7165);
xnor U7378 (N_7378,N_7019,N_7167);
nor U7379 (N_7379,N_7223,N_7003);
nand U7380 (N_7380,N_7160,N_7150);
or U7381 (N_7381,N_7098,N_7179);
xnor U7382 (N_7382,N_7068,N_7212);
nor U7383 (N_7383,N_7050,N_7101);
and U7384 (N_7384,N_7117,N_7090);
and U7385 (N_7385,N_7180,N_7190);
xnor U7386 (N_7386,N_7017,N_7022);
and U7387 (N_7387,N_7044,N_7154);
nor U7388 (N_7388,N_7066,N_7055);
and U7389 (N_7389,N_7091,N_7160);
and U7390 (N_7390,N_7196,N_7199);
nor U7391 (N_7391,N_7027,N_7184);
nand U7392 (N_7392,N_7207,N_7155);
and U7393 (N_7393,N_7227,N_7205);
nand U7394 (N_7394,N_7098,N_7062);
nor U7395 (N_7395,N_7195,N_7067);
and U7396 (N_7396,N_7005,N_7236);
nor U7397 (N_7397,N_7192,N_7036);
and U7398 (N_7398,N_7121,N_7078);
or U7399 (N_7399,N_7194,N_7247);
nor U7400 (N_7400,N_7068,N_7163);
xnor U7401 (N_7401,N_7010,N_7013);
and U7402 (N_7402,N_7207,N_7241);
nor U7403 (N_7403,N_7132,N_7168);
nand U7404 (N_7404,N_7141,N_7025);
nor U7405 (N_7405,N_7161,N_7038);
xor U7406 (N_7406,N_7045,N_7144);
or U7407 (N_7407,N_7001,N_7207);
nor U7408 (N_7408,N_7050,N_7124);
nand U7409 (N_7409,N_7220,N_7021);
nand U7410 (N_7410,N_7179,N_7216);
xnor U7411 (N_7411,N_7157,N_7074);
xnor U7412 (N_7412,N_7140,N_7231);
or U7413 (N_7413,N_7148,N_7085);
nor U7414 (N_7414,N_7186,N_7194);
nand U7415 (N_7415,N_7165,N_7054);
nand U7416 (N_7416,N_7225,N_7210);
xnor U7417 (N_7417,N_7152,N_7198);
xor U7418 (N_7418,N_7098,N_7065);
xor U7419 (N_7419,N_7062,N_7163);
and U7420 (N_7420,N_7098,N_7010);
xor U7421 (N_7421,N_7052,N_7161);
nor U7422 (N_7422,N_7213,N_7137);
and U7423 (N_7423,N_7088,N_7033);
or U7424 (N_7424,N_7232,N_7204);
or U7425 (N_7425,N_7173,N_7016);
xnor U7426 (N_7426,N_7217,N_7215);
or U7427 (N_7427,N_7178,N_7028);
and U7428 (N_7428,N_7190,N_7007);
or U7429 (N_7429,N_7102,N_7022);
and U7430 (N_7430,N_7147,N_7080);
and U7431 (N_7431,N_7072,N_7123);
or U7432 (N_7432,N_7237,N_7087);
nand U7433 (N_7433,N_7174,N_7172);
nor U7434 (N_7434,N_7199,N_7053);
nand U7435 (N_7435,N_7006,N_7135);
xnor U7436 (N_7436,N_7065,N_7153);
or U7437 (N_7437,N_7165,N_7231);
xnor U7438 (N_7438,N_7208,N_7062);
xor U7439 (N_7439,N_7175,N_7047);
nor U7440 (N_7440,N_7046,N_7071);
and U7441 (N_7441,N_7140,N_7216);
nand U7442 (N_7442,N_7113,N_7227);
xnor U7443 (N_7443,N_7146,N_7156);
nor U7444 (N_7444,N_7162,N_7242);
xor U7445 (N_7445,N_7168,N_7054);
xor U7446 (N_7446,N_7155,N_7124);
xor U7447 (N_7447,N_7056,N_7100);
nand U7448 (N_7448,N_7114,N_7159);
or U7449 (N_7449,N_7087,N_7089);
xnor U7450 (N_7450,N_7023,N_7134);
and U7451 (N_7451,N_7182,N_7157);
or U7452 (N_7452,N_7033,N_7245);
or U7453 (N_7453,N_7118,N_7043);
xor U7454 (N_7454,N_7013,N_7027);
and U7455 (N_7455,N_7113,N_7054);
or U7456 (N_7456,N_7138,N_7207);
xor U7457 (N_7457,N_7050,N_7241);
or U7458 (N_7458,N_7010,N_7020);
nand U7459 (N_7459,N_7014,N_7061);
nor U7460 (N_7460,N_7105,N_7224);
and U7461 (N_7461,N_7093,N_7114);
nor U7462 (N_7462,N_7139,N_7050);
nor U7463 (N_7463,N_7119,N_7088);
or U7464 (N_7464,N_7126,N_7207);
and U7465 (N_7465,N_7197,N_7126);
nor U7466 (N_7466,N_7216,N_7173);
nor U7467 (N_7467,N_7125,N_7179);
and U7468 (N_7468,N_7023,N_7205);
nand U7469 (N_7469,N_7010,N_7113);
and U7470 (N_7470,N_7108,N_7201);
nand U7471 (N_7471,N_7176,N_7206);
or U7472 (N_7472,N_7150,N_7207);
and U7473 (N_7473,N_7085,N_7163);
nor U7474 (N_7474,N_7225,N_7194);
nor U7475 (N_7475,N_7157,N_7035);
xnor U7476 (N_7476,N_7065,N_7156);
xnor U7477 (N_7477,N_7014,N_7103);
or U7478 (N_7478,N_7200,N_7085);
and U7479 (N_7479,N_7124,N_7115);
and U7480 (N_7480,N_7190,N_7121);
or U7481 (N_7481,N_7192,N_7103);
or U7482 (N_7482,N_7213,N_7080);
and U7483 (N_7483,N_7155,N_7127);
and U7484 (N_7484,N_7218,N_7184);
xnor U7485 (N_7485,N_7188,N_7171);
xnor U7486 (N_7486,N_7112,N_7168);
nand U7487 (N_7487,N_7240,N_7048);
nand U7488 (N_7488,N_7135,N_7156);
or U7489 (N_7489,N_7248,N_7055);
and U7490 (N_7490,N_7204,N_7201);
nor U7491 (N_7491,N_7149,N_7247);
nor U7492 (N_7492,N_7219,N_7098);
nand U7493 (N_7493,N_7008,N_7054);
nand U7494 (N_7494,N_7238,N_7240);
xor U7495 (N_7495,N_7160,N_7209);
and U7496 (N_7496,N_7014,N_7241);
nor U7497 (N_7497,N_7241,N_7248);
and U7498 (N_7498,N_7016,N_7248);
and U7499 (N_7499,N_7126,N_7199);
xor U7500 (N_7500,N_7458,N_7252);
xor U7501 (N_7501,N_7491,N_7441);
or U7502 (N_7502,N_7492,N_7277);
nand U7503 (N_7503,N_7432,N_7361);
xnor U7504 (N_7504,N_7427,N_7276);
nand U7505 (N_7505,N_7319,N_7425);
or U7506 (N_7506,N_7393,N_7264);
or U7507 (N_7507,N_7478,N_7274);
or U7508 (N_7508,N_7338,N_7485);
and U7509 (N_7509,N_7453,N_7394);
nand U7510 (N_7510,N_7279,N_7424);
nand U7511 (N_7511,N_7429,N_7422);
and U7512 (N_7512,N_7272,N_7299);
nand U7513 (N_7513,N_7423,N_7268);
nor U7514 (N_7514,N_7368,N_7489);
xnor U7515 (N_7515,N_7280,N_7402);
xor U7516 (N_7516,N_7460,N_7262);
nor U7517 (N_7517,N_7426,N_7371);
xnor U7518 (N_7518,N_7396,N_7303);
or U7519 (N_7519,N_7323,N_7488);
xnor U7520 (N_7520,N_7365,N_7446);
nand U7521 (N_7521,N_7398,N_7285);
nor U7522 (N_7522,N_7411,N_7315);
nand U7523 (N_7523,N_7366,N_7403);
xor U7524 (N_7524,N_7344,N_7360);
nor U7525 (N_7525,N_7340,N_7376);
xnor U7526 (N_7526,N_7459,N_7454);
nor U7527 (N_7527,N_7490,N_7378);
xnor U7528 (N_7528,N_7477,N_7325);
xor U7529 (N_7529,N_7468,N_7307);
nand U7530 (N_7530,N_7320,N_7289);
nand U7531 (N_7531,N_7281,N_7282);
or U7532 (N_7532,N_7342,N_7461);
nand U7533 (N_7533,N_7254,N_7436);
or U7534 (N_7534,N_7362,N_7256);
nand U7535 (N_7535,N_7389,N_7487);
and U7536 (N_7536,N_7367,N_7373);
and U7537 (N_7537,N_7442,N_7352);
nor U7538 (N_7538,N_7415,N_7390);
or U7539 (N_7539,N_7283,N_7295);
xnor U7540 (N_7540,N_7462,N_7261);
xnor U7541 (N_7541,N_7294,N_7348);
nor U7542 (N_7542,N_7486,N_7474);
or U7543 (N_7543,N_7407,N_7472);
nand U7544 (N_7544,N_7435,N_7316);
xnor U7545 (N_7545,N_7431,N_7329);
nand U7546 (N_7546,N_7408,N_7418);
and U7547 (N_7547,N_7273,N_7440);
or U7548 (N_7548,N_7457,N_7395);
nor U7549 (N_7549,N_7387,N_7363);
or U7550 (N_7550,N_7445,N_7349);
nor U7551 (N_7551,N_7437,N_7259);
and U7552 (N_7552,N_7484,N_7374);
xor U7553 (N_7553,N_7413,N_7317);
nand U7554 (N_7554,N_7251,N_7287);
nor U7555 (N_7555,N_7313,N_7479);
nor U7556 (N_7556,N_7356,N_7466);
nor U7557 (N_7557,N_7265,N_7300);
xnor U7558 (N_7558,N_7253,N_7383);
nand U7559 (N_7559,N_7420,N_7357);
or U7560 (N_7560,N_7339,N_7439);
nand U7561 (N_7561,N_7456,N_7305);
and U7562 (N_7562,N_7380,N_7297);
nand U7563 (N_7563,N_7464,N_7377);
nor U7564 (N_7564,N_7333,N_7433);
or U7565 (N_7565,N_7482,N_7290);
xor U7566 (N_7566,N_7270,N_7399);
or U7567 (N_7567,N_7417,N_7406);
and U7568 (N_7568,N_7263,N_7269);
and U7569 (N_7569,N_7298,N_7308);
xor U7570 (N_7570,N_7469,N_7260);
or U7571 (N_7571,N_7286,N_7449);
nand U7572 (N_7572,N_7421,N_7384);
and U7573 (N_7573,N_7291,N_7444);
nor U7574 (N_7574,N_7447,N_7443);
xor U7575 (N_7575,N_7463,N_7467);
or U7576 (N_7576,N_7330,N_7312);
xnor U7577 (N_7577,N_7400,N_7428);
or U7578 (N_7578,N_7284,N_7379);
nor U7579 (N_7579,N_7345,N_7288);
nand U7580 (N_7580,N_7306,N_7385);
and U7581 (N_7581,N_7324,N_7480);
nand U7582 (N_7582,N_7388,N_7471);
nand U7583 (N_7583,N_7434,N_7386);
and U7584 (N_7584,N_7301,N_7416);
xnor U7585 (N_7585,N_7498,N_7304);
nor U7586 (N_7586,N_7354,N_7359);
xor U7587 (N_7587,N_7318,N_7255);
and U7588 (N_7588,N_7372,N_7326);
and U7589 (N_7589,N_7404,N_7452);
nand U7590 (N_7590,N_7419,N_7293);
nand U7591 (N_7591,N_7322,N_7438);
and U7592 (N_7592,N_7369,N_7475);
and U7593 (N_7593,N_7309,N_7258);
and U7594 (N_7594,N_7481,N_7292);
or U7595 (N_7595,N_7391,N_7493);
and U7596 (N_7596,N_7430,N_7499);
xor U7597 (N_7597,N_7401,N_7314);
and U7598 (N_7598,N_7267,N_7355);
and U7599 (N_7599,N_7358,N_7311);
and U7600 (N_7600,N_7364,N_7341);
and U7601 (N_7601,N_7278,N_7450);
and U7602 (N_7602,N_7375,N_7353);
and U7603 (N_7603,N_7448,N_7343);
or U7604 (N_7604,N_7302,N_7332);
xor U7605 (N_7605,N_7405,N_7381);
or U7606 (N_7606,N_7455,N_7382);
nor U7607 (N_7607,N_7331,N_7337);
nand U7608 (N_7608,N_7271,N_7397);
nor U7609 (N_7609,N_7328,N_7346);
and U7610 (N_7610,N_7327,N_7476);
and U7611 (N_7611,N_7296,N_7496);
or U7612 (N_7612,N_7321,N_7412);
nand U7613 (N_7613,N_7470,N_7347);
or U7614 (N_7614,N_7275,N_7494);
nor U7615 (N_7615,N_7414,N_7392);
or U7616 (N_7616,N_7370,N_7310);
and U7617 (N_7617,N_7410,N_7465);
xnor U7618 (N_7618,N_7335,N_7257);
nor U7619 (N_7619,N_7334,N_7336);
xnor U7620 (N_7620,N_7451,N_7483);
or U7621 (N_7621,N_7497,N_7409);
and U7622 (N_7622,N_7250,N_7351);
or U7623 (N_7623,N_7350,N_7266);
and U7624 (N_7624,N_7473,N_7495);
nor U7625 (N_7625,N_7266,N_7330);
and U7626 (N_7626,N_7383,N_7380);
and U7627 (N_7627,N_7306,N_7476);
and U7628 (N_7628,N_7282,N_7372);
nand U7629 (N_7629,N_7462,N_7461);
and U7630 (N_7630,N_7447,N_7445);
or U7631 (N_7631,N_7486,N_7350);
or U7632 (N_7632,N_7315,N_7305);
nand U7633 (N_7633,N_7346,N_7337);
nor U7634 (N_7634,N_7377,N_7422);
and U7635 (N_7635,N_7453,N_7399);
or U7636 (N_7636,N_7451,N_7252);
xor U7637 (N_7637,N_7319,N_7273);
nor U7638 (N_7638,N_7297,N_7414);
and U7639 (N_7639,N_7446,N_7416);
xor U7640 (N_7640,N_7254,N_7313);
xor U7641 (N_7641,N_7359,N_7446);
nand U7642 (N_7642,N_7418,N_7402);
nand U7643 (N_7643,N_7433,N_7411);
nand U7644 (N_7644,N_7258,N_7352);
nand U7645 (N_7645,N_7492,N_7458);
nor U7646 (N_7646,N_7308,N_7389);
xor U7647 (N_7647,N_7461,N_7398);
or U7648 (N_7648,N_7465,N_7351);
nor U7649 (N_7649,N_7356,N_7433);
nor U7650 (N_7650,N_7275,N_7457);
or U7651 (N_7651,N_7357,N_7333);
or U7652 (N_7652,N_7312,N_7390);
or U7653 (N_7653,N_7428,N_7385);
and U7654 (N_7654,N_7388,N_7299);
xor U7655 (N_7655,N_7276,N_7441);
or U7656 (N_7656,N_7277,N_7257);
xnor U7657 (N_7657,N_7499,N_7318);
and U7658 (N_7658,N_7442,N_7326);
and U7659 (N_7659,N_7302,N_7250);
nor U7660 (N_7660,N_7408,N_7384);
xor U7661 (N_7661,N_7424,N_7357);
and U7662 (N_7662,N_7341,N_7298);
and U7663 (N_7663,N_7390,N_7428);
or U7664 (N_7664,N_7459,N_7480);
nand U7665 (N_7665,N_7349,N_7487);
nand U7666 (N_7666,N_7444,N_7438);
or U7667 (N_7667,N_7356,N_7439);
xor U7668 (N_7668,N_7429,N_7344);
nand U7669 (N_7669,N_7355,N_7307);
xor U7670 (N_7670,N_7497,N_7325);
and U7671 (N_7671,N_7393,N_7467);
nand U7672 (N_7672,N_7329,N_7408);
or U7673 (N_7673,N_7355,N_7371);
nor U7674 (N_7674,N_7296,N_7487);
or U7675 (N_7675,N_7354,N_7255);
or U7676 (N_7676,N_7377,N_7492);
nand U7677 (N_7677,N_7436,N_7455);
and U7678 (N_7678,N_7258,N_7305);
xnor U7679 (N_7679,N_7278,N_7308);
nor U7680 (N_7680,N_7472,N_7491);
nor U7681 (N_7681,N_7378,N_7368);
xor U7682 (N_7682,N_7278,N_7303);
xor U7683 (N_7683,N_7285,N_7453);
xor U7684 (N_7684,N_7468,N_7390);
nor U7685 (N_7685,N_7261,N_7485);
or U7686 (N_7686,N_7416,N_7326);
xnor U7687 (N_7687,N_7376,N_7375);
nor U7688 (N_7688,N_7371,N_7297);
nand U7689 (N_7689,N_7364,N_7318);
xnor U7690 (N_7690,N_7260,N_7302);
or U7691 (N_7691,N_7343,N_7487);
or U7692 (N_7692,N_7438,N_7406);
xnor U7693 (N_7693,N_7361,N_7397);
nor U7694 (N_7694,N_7382,N_7329);
or U7695 (N_7695,N_7290,N_7484);
nor U7696 (N_7696,N_7287,N_7376);
nor U7697 (N_7697,N_7442,N_7291);
nand U7698 (N_7698,N_7393,N_7267);
nor U7699 (N_7699,N_7370,N_7268);
or U7700 (N_7700,N_7336,N_7378);
and U7701 (N_7701,N_7341,N_7467);
and U7702 (N_7702,N_7317,N_7495);
nor U7703 (N_7703,N_7293,N_7274);
and U7704 (N_7704,N_7313,N_7368);
xor U7705 (N_7705,N_7363,N_7419);
nand U7706 (N_7706,N_7294,N_7378);
and U7707 (N_7707,N_7344,N_7271);
nor U7708 (N_7708,N_7382,N_7480);
or U7709 (N_7709,N_7266,N_7319);
xor U7710 (N_7710,N_7269,N_7313);
or U7711 (N_7711,N_7413,N_7286);
xnor U7712 (N_7712,N_7376,N_7495);
and U7713 (N_7713,N_7324,N_7359);
and U7714 (N_7714,N_7396,N_7295);
or U7715 (N_7715,N_7379,N_7352);
and U7716 (N_7716,N_7483,N_7449);
and U7717 (N_7717,N_7457,N_7309);
and U7718 (N_7718,N_7259,N_7418);
xnor U7719 (N_7719,N_7317,N_7362);
nor U7720 (N_7720,N_7468,N_7292);
and U7721 (N_7721,N_7432,N_7479);
nand U7722 (N_7722,N_7398,N_7307);
and U7723 (N_7723,N_7490,N_7261);
xnor U7724 (N_7724,N_7373,N_7399);
xor U7725 (N_7725,N_7260,N_7389);
nand U7726 (N_7726,N_7400,N_7345);
nor U7727 (N_7727,N_7446,N_7279);
or U7728 (N_7728,N_7359,N_7312);
or U7729 (N_7729,N_7346,N_7427);
nor U7730 (N_7730,N_7477,N_7314);
nor U7731 (N_7731,N_7355,N_7434);
xnor U7732 (N_7732,N_7431,N_7301);
xor U7733 (N_7733,N_7480,N_7423);
and U7734 (N_7734,N_7348,N_7457);
nand U7735 (N_7735,N_7401,N_7357);
and U7736 (N_7736,N_7402,N_7398);
or U7737 (N_7737,N_7360,N_7258);
and U7738 (N_7738,N_7312,N_7429);
or U7739 (N_7739,N_7446,N_7329);
and U7740 (N_7740,N_7391,N_7322);
nor U7741 (N_7741,N_7380,N_7270);
nor U7742 (N_7742,N_7323,N_7327);
and U7743 (N_7743,N_7396,N_7422);
xnor U7744 (N_7744,N_7272,N_7313);
nor U7745 (N_7745,N_7379,N_7340);
xor U7746 (N_7746,N_7326,N_7376);
nor U7747 (N_7747,N_7461,N_7302);
or U7748 (N_7748,N_7257,N_7329);
and U7749 (N_7749,N_7387,N_7486);
nor U7750 (N_7750,N_7581,N_7513);
nor U7751 (N_7751,N_7610,N_7516);
and U7752 (N_7752,N_7655,N_7570);
and U7753 (N_7753,N_7534,N_7543);
or U7754 (N_7754,N_7510,N_7735);
nand U7755 (N_7755,N_7631,N_7638);
or U7756 (N_7756,N_7528,N_7727);
and U7757 (N_7757,N_7734,N_7575);
or U7758 (N_7758,N_7608,N_7685);
nand U7759 (N_7759,N_7676,N_7566);
or U7760 (N_7760,N_7544,N_7607);
and U7761 (N_7761,N_7527,N_7593);
xor U7762 (N_7762,N_7582,N_7609);
and U7763 (N_7763,N_7693,N_7512);
nand U7764 (N_7764,N_7591,N_7634);
and U7765 (N_7765,N_7517,N_7697);
nand U7766 (N_7766,N_7622,N_7678);
nor U7767 (N_7767,N_7669,N_7508);
xor U7768 (N_7768,N_7690,N_7630);
xor U7769 (N_7769,N_7579,N_7551);
and U7770 (N_7770,N_7511,N_7604);
or U7771 (N_7771,N_7686,N_7715);
nor U7772 (N_7772,N_7673,N_7650);
nor U7773 (N_7773,N_7589,N_7654);
and U7774 (N_7774,N_7649,N_7747);
or U7775 (N_7775,N_7620,N_7500);
nor U7776 (N_7776,N_7530,N_7545);
or U7777 (N_7777,N_7587,N_7521);
nor U7778 (N_7778,N_7702,N_7536);
or U7779 (N_7779,N_7635,N_7615);
xnor U7780 (N_7780,N_7731,N_7675);
nand U7781 (N_7781,N_7680,N_7647);
nand U7782 (N_7782,N_7558,N_7606);
nand U7783 (N_7783,N_7605,N_7574);
nor U7784 (N_7784,N_7665,N_7656);
xor U7785 (N_7785,N_7539,N_7623);
and U7786 (N_7786,N_7648,N_7519);
xor U7787 (N_7787,N_7710,N_7625);
nor U7788 (N_7788,N_7719,N_7645);
xor U7789 (N_7789,N_7586,N_7677);
xor U7790 (N_7790,N_7522,N_7712);
and U7791 (N_7791,N_7687,N_7723);
xnor U7792 (N_7792,N_7658,N_7699);
nand U7793 (N_7793,N_7695,N_7639);
nand U7794 (N_7794,N_7692,N_7629);
nor U7795 (N_7795,N_7703,N_7742);
and U7796 (N_7796,N_7683,N_7666);
xor U7797 (N_7797,N_7599,N_7580);
nand U7798 (N_7798,N_7611,N_7661);
nand U7799 (N_7799,N_7515,N_7573);
nand U7800 (N_7800,N_7506,N_7553);
or U7801 (N_7801,N_7636,N_7529);
nand U7802 (N_7802,N_7555,N_7721);
xnor U7803 (N_7803,N_7722,N_7706);
or U7804 (N_7804,N_7682,N_7664);
or U7805 (N_7805,N_7642,N_7595);
or U7806 (N_7806,N_7532,N_7616);
xor U7807 (N_7807,N_7660,N_7741);
nand U7808 (N_7808,N_7739,N_7514);
nand U7809 (N_7809,N_7691,N_7708);
nand U7810 (N_7810,N_7569,N_7507);
and U7811 (N_7811,N_7641,N_7567);
nand U7812 (N_7812,N_7749,N_7711);
nand U7813 (N_7813,N_7704,N_7644);
and U7814 (N_7814,N_7748,N_7554);
and U7815 (N_7815,N_7643,N_7707);
and U7816 (N_7816,N_7738,N_7612);
xor U7817 (N_7817,N_7559,N_7689);
nor U7818 (N_7818,N_7657,N_7526);
nor U7819 (N_7819,N_7621,N_7557);
nand U7820 (N_7820,N_7552,N_7520);
nor U7821 (N_7821,N_7672,N_7578);
xor U7822 (N_7822,N_7617,N_7577);
or U7823 (N_7823,N_7670,N_7568);
or U7824 (N_7824,N_7726,N_7540);
and U7825 (N_7825,N_7600,N_7533);
or U7826 (N_7826,N_7740,N_7572);
xnor U7827 (N_7827,N_7681,N_7561);
or U7828 (N_7828,N_7700,N_7646);
and U7829 (N_7829,N_7556,N_7518);
nand U7830 (N_7830,N_7531,N_7729);
xnor U7831 (N_7831,N_7602,N_7730);
nor U7832 (N_7832,N_7619,N_7637);
nor U7833 (N_7833,N_7594,N_7541);
xnor U7834 (N_7834,N_7598,N_7549);
or U7835 (N_7835,N_7583,N_7732);
nand U7836 (N_7836,N_7714,N_7563);
nor U7837 (N_7837,N_7588,N_7736);
nor U7838 (N_7838,N_7705,N_7524);
or U7839 (N_7839,N_7746,N_7659);
nand U7840 (N_7840,N_7724,N_7560);
nor U7841 (N_7841,N_7501,N_7674);
nor U7842 (N_7842,N_7684,N_7671);
nor U7843 (N_7843,N_7603,N_7547);
xor U7844 (N_7844,N_7505,N_7716);
nand U7845 (N_7845,N_7624,N_7584);
xnor U7846 (N_7846,N_7627,N_7546);
xnor U7847 (N_7847,N_7662,N_7628);
and U7848 (N_7848,N_7633,N_7663);
and U7849 (N_7849,N_7701,N_7550);
xnor U7850 (N_7850,N_7696,N_7614);
and U7851 (N_7851,N_7733,N_7640);
or U7852 (N_7852,N_7651,N_7679);
nor U7853 (N_7853,N_7668,N_7717);
or U7854 (N_7854,N_7535,N_7564);
and U7855 (N_7855,N_7523,N_7652);
and U7856 (N_7856,N_7653,N_7713);
nand U7857 (N_7857,N_7525,N_7562);
nor U7858 (N_7858,N_7698,N_7728);
xor U7859 (N_7859,N_7720,N_7509);
nor U7860 (N_7860,N_7709,N_7718);
nor U7861 (N_7861,N_7502,N_7632);
or U7862 (N_7862,N_7601,N_7571);
xnor U7863 (N_7863,N_7745,N_7618);
xnor U7864 (N_7864,N_7596,N_7597);
nor U7865 (N_7865,N_7694,N_7542);
nor U7866 (N_7866,N_7667,N_7504);
nor U7867 (N_7867,N_7613,N_7725);
xnor U7868 (N_7868,N_7737,N_7537);
nor U7869 (N_7869,N_7590,N_7592);
xnor U7870 (N_7870,N_7744,N_7743);
or U7871 (N_7871,N_7585,N_7548);
or U7872 (N_7872,N_7626,N_7576);
nor U7873 (N_7873,N_7565,N_7688);
nor U7874 (N_7874,N_7503,N_7538);
or U7875 (N_7875,N_7696,N_7684);
xor U7876 (N_7876,N_7603,N_7611);
xnor U7877 (N_7877,N_7509,N_7712);
xor U7878 (N_7878,N_7687,N_7596);
xnor U7879 (N_7879,N_7606,N_7738);
nand U7880 (N_7880,N_7714,N_7640);
nor U7881 (N_7881,N_7739,N_7566);
and U7882 (N_7882,N_7561,N_7604);
nand U7883 (N_7883,N_7518,N_7721);
and U7884 (N_7884,N_7537,N_7580);
nand U7885 (N_7885,N_7501,N_7646);
and U7886 (N_7886,N_7505,N_7583);
and U7887 (N_7887,N_7708,N_7686);
or U7888 (N_7888,N_7622,N_7744);
nand U7889 (N_7889,N_7724,N_7721);
nand U7890 (N_7890,N_7602,N_7684);
and U7891 (N_7891,N_7719,N_7680);
nor U7892 (N_7892,N_7687,N_7727);
xnor U7893 (N_7893,N_7577,N_7551);
or U7894 (N_7894,N_7693,N_7664);
nor U7895 (N_7895,N_7723,N_7581);
xor U7896 (N_7896,N_7533,N_7523);
or U7897 (N_7897,N_7708,N_7695);
and U7898 (N_7898,N_7636,N_7667);
nand U7899 (N_7899,N_7642,N_7715);
xor U7900 (N_7900,N_7619,N_7647);
and U7901 (N_7901,N_7534,N_7730);
and U7902 (N_7902,N_7648,N_7553);
nor U7903 (N_7903,N_7502,N_7731);
and U7904 (N_7904,N_7542,N_7574);
or U7905 (N_7905,N_7550,N_7739);
and U7906 (N_7906,N_7512,N_7613);
nand U7907 (N_7907,N_7610,N_7739);
or U7908 (N_7908,N_7594,N_7627);
nand U7909 (N_7909,N_7728,N_7583);
xor U7910 (N_7910,N_7691,N_7553);
and U7911 (N_7911,N_7518,N_7717);
nor U7912 (N_7912,N_7739,N_7543);
and U7913 (N_7913,N_7618,N_7698);
or U7914 (N_7914,N_7683,N_7684);
and U7915 (N_7915,N_7537,N_7683);
nand U7916 (N_7916,N_7630,N_7560);
and U7917 (N_7917,N_7504,N_7732);
nand U7918 (N_7918,N_7678,N_7584);
nand U7919 (N_7919,N_7588,N_7683);
nor U7920 (N_7920,N_7586,N_7680);
or U7921 (N_7921,N_7577,N_7668);
nand U7922 (N_7922,N_7515,N_7670);
or U7923 (N_7923,N_7693,N_7662);
or U7924 (N_7924,N_7748,N_7715);
nor U7925 (N_7925,N_7530,N_7562);
nand U7926 (N_7926,N_7691,N_7551);
nor U7927 (N_7927,N_7679,N_7649);
nand U7928 (N_7928,N_7674,N_7612);
nand U7929 (N_7929,N_7702,N_7689);
or U7930 (N_7930,N_7736,N_7581);
nor U7931 (N_7931,N_7631,N_7574);
xor U7932 (N_7932,N_7710,N_7507);
xnor U7933 (N_7933,N_7748,N_7536);
xnor U7934 (N_7934,N_7535,N_7573);
xor U7935 (N_7935,N_7516,N_7662);
xnor U7936 (N_7936,N_7533,N_7560);
nor U7937 (N_7937,N_7554,N_7597);
nor U7938 (N_7938,N_7707,N_7625);
xnor U7939 (N_7939,N_7519,N_7549);
nor U7940 (N_7940,N_7597,N_7736);
or U7941 (N_7941,N_7707,N_7533);
or U7942 (N_7942,N_7699,N_7617);
or U7943 (N_7943,N_7547,N_7659);
xor U7944 (N_7944,N_7562,N_7615);
xor U7945 (N_7945,N_7638,N_7703);
or U7946 (N_7946,N_7539,N_7687);
xor U7947 (N_7947,N_7604,N_7575);
xnor U7948 (N_7948,N_7665,N_7568);
nand U7949 (N_7949,N_7630,N_7535);
nand U7950 (N_7950,N_7744,N_7735);
nand U7951 (N_7951,N_7636,N_7647);
nor U7952 (N_7952,N_7708,N_7527);
and U7953 (N_7953,N_7604,N_7622);
nor U7954 (N_7954,N_7693,N_7630);
or U7955 (N_7955,N_7636,N_7747);
nand U7956 (N_7956,N_7542,N_7518);
nand U7957 (N_7957,N_7647,N_7745);
xnor U7958 (N_7958,N_7697,N_7600);
xor U7959 (N_7959,N_7575,N_7576);
nand U7960 (N_7960,N_7574,N_7621);
xnor U7961 (N_7961,N_7605,N_7633);
or U7962 (N_7962,N_7523,N_7697);
xor U7963 (N_7963,N_7667,N_7527);
nor U7964 (N_7964,N_7669,N_7612);
or U7965 (N_7965,N_7532,N_7652);
or U7966 (N_7966,N_7502,N_7649);
or U7967 (N_7967,N_7706,N_7610);
nand U7968 (N_7968,N_7521,N_7710);
xnor U7969 (N_7969,N_7530,N_7528);
and U7970 (N_7970,N_7581,N_7643);
and U7971 (N_7971,N_7614,N_7617);
nand U7972 (N_7972,N_7601,N_7542);
nand U7973 (N_7973,N_7593,N_7674);
and U7974 (N_7974,N_7636,N_7664);
or U7975 (N_7975,N_7644,N_7594);
xnor U7976 (N_7976,N_7688,N_7693);
and U7977 (N_7977,N_7505,N_7699);
nor U7978 (N_7978,N_7582,N_7506);
or U7979 (N_7979,N_7617,N_7681);
nor U7980 (N_7980,N_7682,N_7685);
nor U7981 (N_7981,N_7538,N_7699);
or U7982 (N_7982,N_7567,N_7706);
xor U7983 (N_7983,N_7689,N_7649);
xnor U7984 (N_7984,N_7500,N_7542);
nand U7985 (N_7985,N_7677,N_7587);
nor U7986 (N_7986,N_7632,N_7689);
or U7987 (N_7987,N_7746,N_7709);
or U7988 (N_7988,N_7521,N_7658);
xnor U7989 (N_7989,N_7602,N_7503);
or U7990 (N_7990,N_7521,N_7684);
or U7991 (N_7991,N_7738,N_7659);
nor U7992 (N_7992,N_7505,N_7571);
nand U7993 (N_7993,N_7717,N_7676);
nand U7994 (N_7994,N_7532,N_7555);
or U7995 (N_7995,N_7695,N_7663);
nand U7996 (N_7996,N_7748,N_7736);
and U7997 (N_7997,N_7594,N_7602);
nand U7998 (N_7998,N_7594,N_7612);
nor U7999 (N_7999,N_7516,N_7673);
nor U8000 (N_8000,N_7882,N_7893);
xnor U8001 (N_8001,N_7873,N_7834);
or U8002 (N_8002,N_7789,N_7990);
nand U8003 (N_8003,N_7799,N_7813);
xor U8004 (N_8004,N_7877,N_7851);
or U8005 (N_8005,N_7751,N_7975);
and U8006 (N_8006,N_7819,N_7782);
nand U8007 (N_8007,N_7901,N_7937);
xor U8008 (N_8008,N_7750,N_7986);
xor U8009 (N_8009,N_7856,N_7870);
nor U8010 (N_8010,N_7818,N_7754);
xnor U8011 (N_8011,N_7933,N_7858);
and U8012 (N_8012,N_7991,N_7864);
xnor U8013 (N_8013,N_7906,N_7766);
or U8014 (N_8014,N_7950,N_7898);
xor U8015 (N_8015,N_7938,N_7796);
nand U8016 (N_8016,N_7866,N_7757);
nand U8017 (N_8017,N_7768,N_7949);
xor U8018 (N_8018,N_7935,N_7921);
xnor U8019 (N_8019,N_7947,N_7971);
nor U8020 (N_8020,N_7784,N_7867);
nand U8021 (N_8021,N_7832,N_7781);
and U8022 (N_8022,N_7923,N_7995);
xor U8023 (N_8023,N_7999,N_7835);
nand U8024 (N_8024,N_7918,N_7831);
and U8025 (N_8025,N_7814,N_7763);
or U8026 (N_8026,N_7964,N_7854);
or U8027 (N_8027,N_7869,N_7974);
nand U8028 (N_8028,N_7857,N_7800);
and U8029 (N_8029,N_7953,N_7759);
xor U8030 (N_8030,N_7826,N_7977);
and U8031 (N_8031,N_7954,N_7761);
and U8032 (N_8032,N_7758,N_7778);
xnor U8033 (N_8033,N_7776,N_7876);
xnor U8034 (N_8034,N_7978,N_7773);
nor U8035 (N_8035,N_7994,N_7943);
nand U8036 (N_8036,N_7793,N_7765);
xnor U8037 (N_8037,N_7913,N_7828);
or U8038 (N_8038,N_7902,N_7880);
nor U8039 (N_8039,N_7941,N_7993);
nor U8040 (N_8040,N_7997,N_7878);
nor U8041 (N_8041,N_7900,N_7940);
and U8042 (N_8042,N_7904,N_7968);
xnor U8043 (N_8043,N_7770,N_7909);
and U8044 (N_8044,N_7946,N_7973);
and U8045 (N_8045,N_7772,N_7911);
xor U8046 (N_8046,N_7910,N_7969);
and U8047 (N_8047,N_7847,N_7932);
or U8048 (N_8048,N_7797,N_7895);
or U8049 (N_8049,N_7959,N_7767);
nor U8050 (N_8050,N_7822,N_7861);
xnor U8051 (N_8051,N_7794,N_7920);
nand U8052 (N_8052,N_7887,N_7816);
or U8053 (N_8053,N_7976,N_7981);
xnor U8054 (N_8054,N_7802,N_7939);
and U8055 (N_8055,N_7865,N_7982);
nand U8056 (N_8056,N_7827,N_7868);
and U8057 (N_8057,N_7899,N_7948);
and U8058 (N_8058,N_7843,N_7779);
nand U8059 (N_8059,N_7956,N_7919);
and U8060 (N_8060,N_7934,N_7842);
xnor U8061 (N_8061,N_7889,N_7836);
nand U8062 (N_8062,N_7989,N_7785);
nand U8063 (N_8063,N_7891,N_7775);
and U8064 (N_8064,N_7958,N_7855);
nor U8065 (N_8065,N_7929,N_7965);
xor U8066 (N_8066,N_7885,N_7848);
nor U8067 (N_8067,N_7945,N_7801);
and U8068 (N_8068,N_7815,N_7984);
nor U8069 (N_8069,N_7853,N_7985);
nand U8070 (N_8070,N_7980,N_7809);
xnor U8071 (N_8071,N_7849,N_7908);
xnor U8072 (N_8072,N_7783,N_7774);
xor U8073 (N_8073,N_7825,N_7924);
and U8074 (N_8074,N_7795,N_7798);
and U8075 (N_8075,N_7962,N_7996);
nand U8076 (N_8076,N_7808,N_7823);
nor U8077 (N_8077,N_7931,N_7963);
or U8078 (N_8078,N_7803,N_7805);
nand U8079 (N_8079,N_7916,N_7791);
and U8080 (N_8080,N_7756,N_7896);
xor U8081 (N_8081,N_7979,N_7957);
or U8082 (N_8082,N_7915,N_7804);
or U8083 (N_8083,N_7967,N_7886);
nor U8084 (N_8084,N_7839,N_7860);
nor U8085 (N_8085,N_7951,N_7983);
or U8086 (N_8086,N_7961,N_7926);
xor U8087 (N_8087,N_7811,N_7883);
or U8088 (N_8088,N_7787,N_7907);
or U8089 (N_8089,N_7960,N_7764);
or U8090 (N_8090,N_7824,N_7755);
xor U8091 (N_8091,N_7844,N_7894);
and U8092 (N_8092,N_7928,N_7936);
or U8093 (N_8093,N_7863,N_7771);
or U8094 (N_8094,N_7897,N_7806);
nor U8095 (N_8095,N_7927,N_7917);
and U8096 (N_8096,N_7753,N_7871);
or U8097 (N_8097,N_7905,N_7884);
and U8098 (N_8098,N_7888,N_7859);
xnor U8099 (N_8099,N_7792,N_7872);
or U8100 (N_8100,N_7762,N_7972);
nand U8101 (N_8101,N_7966,N_7875);
xnor U8102 (N_8102,N_7852,N_7970);
and U8103 (N_8103,N_7944,N_7833);
nor U8104 (N_8104,N_7846,N_7838);
nor U8105 (N_8105,N_7845,N_7812);
xor U8106 (N_8106,N_7769,N_7998);
or U8107 (N_8107,N_7925,N_7837);
and U8108 (N_8108,N_7777,N_7879);
xnor U8109 (N_8109,N_7850,N_7942);
xnor U8110 (N_8110,N_7820,N_7788);
xnor U8111 (N_8111,N_7952,N_7760);
xnor U8112 (N_8112,N_7922,N_7914);
or U8113 (N_8113,N_7830,N_7874);
nand U8114 (N_8114,N_7807,N_7930);
xor U8115 (N_8115,N_7786,N_7790);
nand U8116 (N_8116,N_7841,N_7988);
nor U8117 (N_8117,N_7892,N_7829);
or U8118 (N_8118,N_7862,N_7912);
and U8119 (N_8119,N_7890,N_7840);
nand U8120 (N_8120,N_7780,N_7752);
or U8121 (N_8121,N_7821,N_7987);
xnor U8122 (N_8122,N_7881,N_7903);
nor U8123 (N_8123,N_7955,N_7810);
nor U8124 (N_8124,N_7817,N_7992);
nand U8125 (N_8125,N_7834,N_7885);
nand U8126 (N_8126,N_7852,N_7950);
xor U8127 (N_8127,N_7992,N_7828);
xnor U8128 (N_8128,N_7939,N_7919);
and U8129 (N_8129,N_7839,N_7859);
nor U8130 (N_8130,N_7814,N_7766);
and U8131 (N_8131,N_7900,N_7812);
and U8132 (N_8132,N_7970,N_7912);
and U8133 (N_8133,N_7985,N_7824);
xnor U8134 (N_8134,N_7969,N_7776);
or U8135 (N_8135,N_7937,N_7998);
nor U8136 (N_8136,N_7755,N_7893);
nor U8137 (N_8137,N_7762,N_7885);
nor U8138 (N_8138,N_7864,N_7850);
or U8139 (N_8139,N_7798,N_7937);
or U8140 (N_8140,N_7994,N_7858);
xor U8141 (N_8141,N_7753,N_7908);
xnor U8142 (N_8142,N_7915,N_7797);
or U8143 (N_8143,N_7754,N_7780);
xnor U8144 (N_8144,N_7876,N_7896);
and U8145 (N_8145,N_7945,N_7907);
nor U8146 (N_8146,N_7769,N_7945);
nand U8147 (N_8147,N_7864,N_7967);
nand U8148 (N_8148,N_7843,N_7753);
or U8149 (N_8149,N_7981,N_7869);
nand U8150 (N_8150,N_7836,N_7863);
nor U8151 (N_8151,N_7999,N_7752);
nand U8152 (N_8152,N_7910,N_7977);
and U8153 (N_8153,N_7873,N_7919);
or U8154 (N_8154,N_7888,N_7780);
nor U8155 (N_8155,N_7897,N_7847);
or U8156 (N_8156,N_7806,N_7867);
or U8157 (N_8157,N_7894,N_7847);
or U8158 (N_8158,N_7983,N_7985);
nor U8159 (N_8159,N_7992,N_7889);
or U8160 (N_8160,N_7826,N_7750);
nor U8161 (N_8161,N_7980,N_7988);
and U8162 (N_8162,N_7943,N_7786);
and U8163 (N_8163,N_7939,N_7948);
or U8164 (N_8164,N_7795,N_7805);
nor U8165 (N_8165,N_7751,N_7771);
xnor U8166 (N_8166,N_7855,N_7856);
or U8167 (N_8167,N_7783,N_7921);
nand U8168 (N_8168,N_7995,N_7948);
or U8169 (N_8169,N_7829,N_7891);
and U8170 (N_8170,N_7852,N_7751);
or U8171 (N_8171,N_7894,N_7820);
nand U8172 (N_8172,N_7987,N_7803);
nor U8173 (N_8173,N_7945,N_7783);
or U8174 (N_8174,N_7791,N_7982);
and U8175 (N_8175,N_7863,N_7933);
or U8176 (N_8176,N_7866,N_7820);
nor U8177 (N_8177,N_7817,N_7807);
nand U8178 (N_8178,N_7872,N_7846);
and U8179 (N_8179,N_7841,N_7892);
nor U8180 (N_8180,N_7757,N_7898);
nor U8181 (N_8181,N_7808,N_7802);
nor U8182 (N_8182,N_7901,N_7974);
nor U8183 (N_8183,N_7908,N_7859);
nor U8184 (N_8184,N_7990,N_7889);
xnor U8185 (N_8185,N_7902,N_7981);
nor U8186 (N_8186,N_7887,N_7933);
nand U8187 (N_8187,N_7774,N_7990);
xor U8188 (N_8188,N_7794,N_7909);
nand U8189 (N_8189,N_7770,N_7998);
or U8190 (N_8190,N_7974,N_7883);
nor U8191 (N_8191,N_7843,N_7821);
and U8192 (N_8192,N_7847,N_7951);
and U8193 (N_8193,N_7936,N_7895);
nand U8194 (N_8194,N_7986,N_7897);
nor U8195 (N_8195,N_7961,N_7925);
nor U8196 (N_8196,N_7849,N_7859);
xnor U8197 (N_8197,N_7864,N_7898);
xor U8198 (N_8198,N_7817,N_7829);
and U8199 (N_8199,N_7808,N_7789);
nor U8200 (N_8200,N_7757,N_7873);
and U8201 (N_8201,N_7768,N_7751);
xnor U8202 (N_8202,N_7919,N_7923);
and U8203 (N_8203,N_7931,N_7949);
nor U8204 (N_8204,N_7933,N_7826);
xor U8205 (N_8205,N_7913,N_7815);
nand U8206 (N_8206,N_7827,N_7997);
nand U8207 (N_8207,N_7849,N_7975);
xnor U8208 (N_8208,N_7950,N_7783);
and U8209 (N_8209,N_7835,N_7936);
nand U8210 (N_8210,N_7773,N_7951);
and U8211 (N_8211,N_7795,N_7913);
xnor U8212 (N_8212,N_7799,N_7769);
or U8213 (N_8213,N_7866,N_7998);
and U8214 (N_8214,N_7997,N_7828);
and U8215 (N_8215,N_7761,N_7825);
and U8216 (N_8216,N_7804,N_7936);
xnor U8217 (N_8217,N_7758,N_7985);
nand U8218 (N_8218,N_7857,N_7759);
nor U8219 (N_8219,N_7956,N_7766);
nand U8220 (N_8220,N_7766,N_7793);
nand U8221 (N_8221,N_7823,N_7948);
or U8222 (N_8222,N_7863,N_7907);
and U8223 (N_8223,N_7942,N_7767);
and U8224 (N_8224,N_7942,N_7967);
nor U8225 (N_8225,N_7769,N_7855);
and U8226 (N_8226,N_7911,N_7885);
or U8227 (N_8227,N_7985,N_7860);
or U8228 (N_8228,N_7795,N_7964);
and U8229 (N_8229,N_7913,N_7961);
nor U8230 (N_8230,N_7828,N_7951);
and U8231 (N_8231,N_7876,N_7765);
xnor U8232 (N_8232,N_7974,N_7965);
nand U8233 (N_8233,N_7853,N_7764);
nand U8234 (N_8234,N_7839,N_7797);
nor U8235 (N_8235,N_7968,N_7825);
and U8236 (N_8236,N_7876,N_7907);
and U8237 (N_8237,N_7835,N_7918);
or U8238 (N_8238,N_7777,N_7832);
nor U8239 (N_8239,N_7868,N_7914);
or U8240 (N_8240,N_7997,N_7837);
and U8241 (N_8241,N_7766,N_7976);
nand U8242 (N_8242,N_7882,N_7824);
nand U8243 (N_8243,N_7863,N_7879);
or U8244 (N_8244,N_7890,N_7957);
xor U8245 (N_8245,N_7848,N_7927);
xor U8246 (N_8246,N_7780,N_7920);
nor U8247 (N_8247,N_7933,N_7924);
nand U8248 (N_8248,N_7854,N_7999);
nand U8249 (N_8249,N_7920,N_7752);
or U8250 (N_8250,N_8216,N_8140);
or U8251 (N_8251,N_8009,N_8185);
and U8252 (N_8252,N_8070,N_8133);
nand U8253 (N_8253,N_8197,N_8227);
nor U8254 (N_8254,N_8134,N_8199);
xnor U8255 (N_8255,N_8006,N_8025);
or U8256 (N_8256,N_8183,N_8231);
nor U8257 (N_8257,N_8058,N_8213);
and U8258 (N_8258,N_8132,N_8000);
nor U8259 (N_8259,N_8243,N_8080);
or U8260 (N_8260,N_8190,N_8019);
or U8261 (N_8261,N_8012,N_8201);
xor U8262 (N_8262,N_8163,N_8142);
nand U8263 (N_8263,N_8114,N_8097);
or U8264 (N_8264,N_8008,N_8159);
nand U8265 (N_8265,N_8221,N_8143);
and U8266 (N_8266,N_8071,N_8095);
and U8267 (N_8267,N_8115,N_8112);
and U8268 (N_8268,N_8144,N_8057);
or U8269 (N_8269,N_8053,N_8018);
nor U8270 (N_8270,N_8076,N_8034);
xor U8271 (N_8271,N_8189,N_8020);
nor U8272 (N_8272,N_8068,N_8110);
and U8273 (N_8273,N_8127,N_8055);
nor U8274 (N_8274,N_8172,N_8167);
and U8275 (N_8275,N_8072,N_8026);
or U8276 (N_8276,N_8249,N_8177);
nand U8277 (N_8277,N_8063,N_8091);
xnor U8278 (N_8278,N_8088,N_8036);
and U8279 (N_8279,N_8217,N_8168);
xnor U8280 (N_8280,N_8105,N_8222);
nor U8281 (N_8281,N_8089,N_8078);
or U8282 (N_8282,N_8171,N_8161);
and U8283 (N_8283,N_8215,N_8062);
and U8284 (N_8284,N_8052,N_8146);
nand U8285 (N_8285,N_8073,N_8176);
or U8286 (N_8286,N_8113,N_8188);
or U8287 (N_8287,N_8067,N_8193);
nand U8288 (N_8288,N_8048,N_8103);
and U8289 (N_8289,N_8044,N_8242);
xnor U8290 (N_8290,N_8029,N_8016);
xnor U8291 (N_8291,N_8230,N_8210);
and U8292 (N_8292,N_8235,N_8107);
xnor U8293 (N_8293,N_8118,N_8245);
xor U8294 (N_8294,N_8028,N_8138);
nor U8295 (N_8295,N_8056,N_8017);
nand U8296 (N_8296,N_8220,N_8094);
xor U8297 (N_8297,N_8131,N_8060);
nor U8298 (N_8298,N_8077,N_8137);
or U8299 (N_8299,N_8125,N_8169);
or U8300 (N_8300,N_8240,N_8027);
and U8301 (N_8301,N_8074,N_8150);
and U8302 (N_8302,N_8135,N_8152);
nand U8303 (N_8303,N_8211,N_8079);
or U8304 (N_8304,N_8180,N_8236);
nor U8305 (N_8305,N_8232,N_8153);
nor U8306 (N_8306,N_8139,N_8010);
and U8307 (N_8307,N_8162,N_8156);
xnor U8308 (N_8308,N_8015,N_8084);
xor U8309 (N_8309,N_8164,N_8234);
xnor U8310 (N_8310,N_8149,N_8247);
nor U8311 (N_8311,N_8106,N_8136);
xor U8312 (N_8312,N_8109,N_8181);
and U8313 (N_8313,N_8011,N_8233);
or U8314 (N_8314,N_8130,N_8219);
and U8315 (N_8315,N_8204,N_8248);
nor U8316 (N_8316,N_8206,N_8087);
nand U8317 (N_8317,N_8148,N_8226);
nor U8318 (N_8318,N_8075,N_8117);
and U8319 (N_8319,N_8225,N_8104);
or U8320 (N_8320,N_8124,N_8207);
nor U8321 (N_8321,N_8154,N_8013);
or U8322 (N_8322,N_8166,N_8228);
or U8323 (N_8323,N_8175,N_8155);
or U8324 (N_8324,N_8083,N_8041);
nor U8325 (N_8325,N_8195,N_8239);
nand U8326 (N_8326,N_8099,N_8005);
nor U8327 (N_8327,N_8157,N_8066);
and U8328 (N_8328,N_8192,N_8173);
or U8329 (N_8329,N_8049,N_8209);
and U8330 (N_8330,N_8065,N_8021);
and U8331 (N_8331,N_8059,N_8102);
or U8332 (N_8332,N_8141,N_8208);
xor U8333 (N_8333,N_8024,N_8246);
xnor U8334 (N_8334,N_8128,N_8238);
xnor U8335 (N_8335,N_8223,N_8047);
and U8336 (N_8336,N_8182,N_8050);
or U8337 (N_8337,N_8096,N_8160);
nor U8338 (N_8338,N_8002,N_8100);
xnor U8339 (N_8339,N_8186,N_8165);
nor U8340 (N_8340,N_8198,N_8122);
nand U8341 (N_8341,N_8241,N_8203);
nand U8342 (N_8342,N_8212,N_8061);
nor U8343 (N_8343,N_8196,N_8126);
or U8344 (N_8344,N_8040,N_8145);
nand U8345 (N_8345,N_8116,N_8121);
nand U8346 (N_8346,N_8064,N_8101);
and U8347 (N_8347,N_8174,N_8093);
xnor U8348 (N_8348,N_8200,N_8123);
nand U8349 (N_8349,N_8082,N_8007);
or U8350 (N_8350,N_8111,N_8098);
nor U8351 (N_8351,N_8014,N_8214);
nor U8352 (N_8352,N_8042,N_8086);
or U8353 (N_8353,N_8187,N_8218);
xor U8354 (N_8354,N_8129,N_8037);
nand U8355 (N_8355,N_8205,N_8184);
xnor U8356 (N_8356,N_8229,N_8244);
or U8357 (N_8357,N_8081,N_8033);
nor U8358 (N_8358,N_8202,N_8085);
nor U8359 (N_8359,N_8237,N_8120);
nor U8360 (N_8360,N_8035,N_8147);
or U8361 (N_8361,N_8158,N_8046);
xor U8362 (N_8362,N_8069,N_8045);
nand U8363 (N_8363,N_8090,N_8004);
nor U8364 (N_8364,N_8032,N_8108);
or U8365 (N_8365,N_8179,N_8038);
nand U8366 (N_8366,N_8191,N_8031);
or U8367 (N_8367,N_8054,N_8030);
nor U8368 (N_8368,N_8022,N_8170);
nand U8369 (N_8369,N_8001,N_8023);
or U8370 (N_8370,N_8051,N_8178);
xor U8371 (N_8371,N_8194,N_8151);
nor U8372 (N_8372,N_8092,N_8119);
and U8373 (N_8373,N_8039,N_8003);
nand U8374 (N_8374,N_8224,N_8043);
xnor U8375 (N_8375,N_8094,N_8007);
nor U8376 (N_8376,N_8092,N_8156);
nor U8377 (N_8377,N_8039,N_8040);
and U8378 (N_8378,N_8084,N_8151);
nor U8379 (N_8379,N_8075,N_8113);
xnor U8380 (N_8380,N_8050,N_8169);
nand U8381 (N_8381,N_8074,N_8055);
and U8382 (N_8382,N_8044,N_8020);
xnor U8383 (N_8383,N_8228,N_8237);
and U8384 (N_8384,N_8189,N_8127);
xor U8385 (N_8385,N_8097,N_8071);
nand U8386 (N_8386,N_8247,N_8108);
nand U8387 (N_8387,N_8044,N_8093);
and U8388 (N_8388,N_8097,N_8175);
nand U8389 (N_8389,N_8235,N_8006);
or U8390 (N_8390,N_8166,N_8045);
or U8391 (N_8391,N_8135,N_8057);
or U8392 (N_8392,N_8047,N_8019);
and U8393 (N_8393,N_8059,N_8050);
nor U8394 (N_8394,N_8165,N_8178);
or U8395 (N_8395,N_8170,N_8245);
nand U8396 (N_8396,N_8139,N_8104);
xnor U8397 (N_8397,N_8243,N_8153);
or U8398 (N_8398,N_8099,N_8087);
or U8399 (N_8399,N_8107,N_8193);
and U8400 (N_8400,N_8213,N_8234);
or U8401 (N_8401,N_8213,N_8176);
xor U8402 (N_8402,N_8119,N_8093);
and U8403 (N_8403,N_8009,N_8059);
xor U8404 (N_8404,N_8241,N_8082);
and U8405 (N_8405,N_8099,N_8200);
or U8406 (N_8406,N_8028,N_8211);
and U8407 (N_8407,N_8015,N_8174);
nand U8408 (N_8408,N_8237,N_8019);
or U8409 (N_8409,N_8125,N_8081);
and U8410 (N_8410,N_8103,N_8112);
or U8411 (N_8411,N_8004,N_8184);
or U8412 (N_8412,N_8229,N_8248);
xor U8413 (N_8413,N_8079,N_8064);
nand U8414 (N_8414,N_8173,N_8239);
and U8415 (N_8415,N_8068,N_8237);
xnor U8416 (N_8416,N_8012,N_8236);
or U8417 (N_8417,N_8059,N_8133);
nand U8418 (N_8418,N_8090,N_8129);
and U8419 (N_8419,N_8218,N_8224);
xor U8420 (N_8420,N_8201,N_8065);
or U8421 (N_8421,N_8014,N_8104);
nand U8422 (N_8422,N_8235,N_8154);
and U8423 (N_8423,N_8035,N_8041);
nand U8424 (N_8424,N_8243,N_8059);
nor U8425 (N_8425,N_8206,N_8225);
xnor U8426 (N_8426,N_8014,N_8225);
xnor U8427 (N_8427,N_8059,N_8001);
nor U8428 (N_8428,N_8204,N_8035);
xor U8429 (N_8429,N_8225,N_8111);
or U8430 (N_8430,N_8123,N_8130);
xor U8431 (N_8431,N_8033,N_8106);
xnor U8432 (N_8432,N_8249,N_8085);
nor U8433 (N_8433,N_8135,N_8231);
or U8434 (N_8434,N_8030,N_8092);
nor U8435 (N_8435,N_8234,N_8093);
or U8436 (N_8436,N_8009,N_8060);
nand U8437 (N_8437,N_8210,N_8217);
or U8438 (N_8438,N_8128,N_8092);
or U8439 (N_8439,N_8029,N_8031);
nand U8440 (N_8440,N_8018,N_8129);
nand U8441 (N_8441,N_8213,N_8188);
nand U8442 (N_8442,N_8114,N_8027);
and U8443 (N_8443,N_8067,N_8180);
nand U8444 (N_8444,N_8126,N_8167);
and U8445 (N_8445,N_8077,N_8098);
nor U8446 (N_8446,N_8154,N_8139);
nor U8447 (N_8447,N_8129,N_8055);
or U8448 (N_8448,N_8007,N_8046);
nor U8449 (N_8449,N_8198,N_8152);
or U8450 (N_8450,N_8213,N_8091);
and U8451 (N_8451,N_8216,N_8207);
nor U8452 (N_8452,N_8085,N_8156);
nor U8453 (N_8453,N_8155,N_8180);
nand U8454 (N_8454,N_8163,N_8147);
xor U8455 (N_8455,N_8239,N_8164);
xnor U8456 (N_8456,N_8073,N_8153);
nor U8457 (N_8457,N_8150,N_8019);
nor U8458 (N_8458,N_8059,N_8207);
or U8459 (N_8459,N_8130,N_8134);
nor U8460 (N_8460,N_8114,N_8079);
and U8461 (N_8461,N_8010,N_8050);
nand U8462 (N_8462,N_8063,N_8026);
xor U8463 (N_8463,N_8070,N_8089);
xor U8464 (N_8464,N_8007,N_8042);
nor U8465 (N_8465,N_8157,N_8090);
xor U8466 (N_8466,N_8212,N_8169);
nand U8467 (N_8467,N_8046,N_8192);
or U8468 (N_8468,N_8022,N_8011);
and U8469 (N_8469,N_8111,N_8210);
and U8470 (N_8470,N_8056,N_8028);
nor U8471 (N_8471,N_8225,N_8031);
nand U8472 (N_8472,N_8180,N_8198);
nor U8473 (N_8473,N_8088,N_8178);
or U8474 (N_8474,N_8009,N_8165);
xnor U8475 (N_8475,N_8073,N_8005);
nor U8476 (N_8476,N_8203,N_8159);
xor U8477 (N_8477,N_8025,N_8038);
or U8478 (N_8478,N_8015,N_8217);
or U8479 (N_8479,N_8201,N_8195);
nor U8480 (N_8480,N_8161,N_8109);
or U8481 (N_8481,N_8236,N_8204);
nor U8482 (N_8482,N_8030,N_8102);
xnor U8483 (N_8483,N_8149,N_8171);
xnor U8484 (N_8484,N_8113,N_8073);
and U8485 (N_8485,N_8211,N_8026);
xnor U8486 (N_8486,N_8080,N_8000);
nor U8487 (N_8487,N_8082,N_8073);
xor U8488 (N_8488,N_8181,N_8137);
nor U8489 (N_8489,N_8045,N_8134);
or U8490 (N_8490,N_8202,N_8134);
nor U8491 (N_8491,N_8112,N_8223);
and U8492 (N_8492,N_8062,N_8013);
and U8493 (N_8493,N_8246,N_8163);
xor U8494 (N_8494,N_8151,N_8065);
or U8495 (N_8495,N_8086,N_8055);
and U8496 (N_8496,N_8063,N_8025);
nand U8497 (N_8497,N_8147,N_8206);
xor U8498 (N_8498,N_8241,N_8043);
nand U8499 (N_8499,N_8038,N_8136);
or U8500 (N_8500,N_8323,N_8303);
and U8501 (N_8501,N_8468,N_8403);
nor U8502 (N_8502,N_8496,N_8493);
xnor U8503 (N_8503,N_8474,N_8434);
xnor U8504 (N_8504,N_8495,N_8290);
xor U8505 (N_8505,N_8302,N_8274);
nand U8506 (N_8506,N_8492,N_8327);
and U8507 (N_8507,N_8344,N_8418);
nand U8508 (N_8508,N_8367,N_8338);
or U8509 (N_8509,N_8253,N_8266);
nor U8510 (N_8510,N_8309,N_8473);
or U8511 (N_8511,N_8422,N_8314);
or U8512 (N_8512,N_8384,N_8287);
nor U8513 (N_8513,N_8446,N_8307);
xnor U8514 (N_8514,N_8297,N_8352);
nand U8515 (N_8515,N_8386,N_8340);
nor U8516 (N_8516,N_8481,N_8391);
xnor U8517 (N_8517,N_8280,N_8353);
nor U8518 (N_8518,N_8431,N_8430);
or U8519 (N_8519,N_8469,N_8343);
or U8520 (N_8520,N_8285,N_8470);
xnor U8521 (N_8521,N_8402,N_8480);
or U8522 (N_8522,N_8254,N_8362);
or U8523 (N_8523,N_8483,N_8273);
nor U8524 (N_8524,N_8256,N_8310);
xor U8525 (N_8525,N_8326,N_8337);
or U8526 (N_8526,N_8479,N_8284);
xnor U8527 (N_8527,N_8417,N_8251);
and U8528 (N_8528,N_8459,N_8399);
nor U8529 (N_8529,N_8457,N_8361);
nor U8530 (N_8530,N_8433,N_8421);
nor U8531 (N_8531,N_8313,N_8382);
xor U8532 (N_8532,N_8317,N_8330);
xnor U8533 (N_8533,N_8356,N_8372);
xnor U8534 (N_8534,N_8415,N_8250);
nand U8535 (N_8535,N_8440,N_8265);
and U8536 (N_8536,N_8429,N_8363);
or U8537 (N_8537,N_8445,N_8279);
nor U8538 (N_8538,N_8490,N_8437);
nand U8539 (N_8539,N_8351,N_8405);
nor U8540 (N_8540,N_8296,N_8370);
nand U8541 (N_8541,N_8312,N_8349);
xor U8542 (N_8542,N_8329,N_8319);
nor U8543 (N_8543,N_8424,N_8278);
nor U8544 (N_8544,N_8339,N_8321);
nand U8545 (N_8545,N_8258,N_8320);
or U8546 (N_8546,N_8393,N_8288);
nor U8547 (N_8547,N_8374,N_8301);
nand U8548 (N_8548,N_8420,N_8345);
or U8549 (N_8549,N_8419,N_8277);
and U8550 (N_8550,N_8414,N_8252);
xor U8551 (N_8551,N_8447,N_8442);
nor U8552 (N_8552,N_8272,N_8260);
or U8553 (N_8553,N_8293,N_8304);
nor U8554 (N_8554,N_8315,N_8289);
or U8555 (N_8555,N_8400,N_8439);
and U8556 (N_8556,N_8358,N_8416);
or U8557 (N_8557,N_8404,N_8281);
nor U8558 (N_8558,N_8471,N_8385);
or U8559 (N_8559,N_8291,N_8380);
xor U8560 (N_8560,N_8411,N_8466);
nor U8561 (N_8561,N_8295,N_8394);
xor U8562 (N_8562,N_8488,N_8465);
nor U8563 (N_8563,N_8462,N_8375);
nand U8564 (N_8564,N_8268,N_8441);
nand U8565 (N_8565,N_8426,N_8498);
nor U8566 (N_8566,N_8423,N_8267);
and U8567 (N_8567,N_8453,N_8478);
nor U8568 (N_8568,N_8491,N_8325);
nor U8569 (N_8569,N_8334,N_8472);
and U8570 (N_8570,N_8322,N_8324);
or U8571 (N_8571,N_8379,N_8298);
xor U8572 (N_8572,N_8275,N_8286);
xnor U8573 (N_8573,N_8332,N_8477);
or U8574 (N_8574,N_8333,N_8276);
or U8575 (N_8575,N_8341,N_8262);
and U8576 (N_8576,N_8456,N_8318);
nor U8577 (N_8577,N_8255,N_8408);
nor U8578 (N_8578,N_8264,N_8450);
nand U8579 (N_8579,N_8406,N_8387);
xnor U8580 (N_8580,N_8371,N_8342);
xnor U8581 (N_8581,N_8388,N_8427);
or U8582 (N_8582,N_8475,N_8487);
xor U8583 (N_8583,N_8395,N_8270);
or U8584 (N_8584,N_8463,N_8455);
or U8585 (N_8585,N_8397,N_8355);
nor U8586 (N_8586,N_8452,N_8360);
and U8587 (N_8587,N_8428,N_8389);
nand U8588 (N_8588,N_8294,N_8454);
nor U8589 (N_8589,N_8282,N_8464);
and U8590 (N_8590,N_8259,N_8368);
or U8591 (N_8591,N_8438,N_8377);
nand U8592 (N_8592,N_8366,N_8482);
or U8593 (N_8593,N_8269,N_8392);
nor U8594 (N_8594,N_8410,N_8364);
nand U8595 (N_8595,N_8444,N_8308);
nor U8596 (N_8596,N_8489,N_8436);
or U8597 (N_8597,N_8497,N_8299);
nand U8598 (N_8598,N_8376,N_8486);
nor U8599 (N_8599,N_8316,N_8373);
and U8600 (N_8600,N_8409,N_8331);
nor U8601 (N_8601,N_8396,N_8398);
and U8602 (N_8602,N_8357,N_8413);
or U8603 (N_8603,N_8476,N_8369);
and U8604 (N_8604,N_8350,N_8346);
nor U8605 (N_8605,N_8263,N_8261);
xor U8606 (N_8606,N_8365,N_8407);
and U8607 (N_8607,N_8435,N_8311);
nand U8608 (N_8608,N_8432,N_8328);
or U8609 (N_8609,N_8494,N_8401);
and U8610 (N_8610,N_8467,N_8347);
nor U8611 (N_8611,N_8461,N_8378);
and U8612 (N_8612,N_8448,N_8484);
and U8613 (N_8613,N_8292,N_8499);
xnor U8614 (N_8614,N_8381,N_8348);
xor U8615 (N_8615,N_8300,N_8306);
nand U8616 (N_8616,N_8257,N_8336);
xnor U8617 (N_8617,N_8354,N_8359);
or U8618 (N_8618,N_8283,N_8383);
nor U8619 (N_8619,N_8271,N_8425);
nor U8620 (N_8620,N_8412,N_8458);
xor U8621 (N_8621,N_8390,N_8485);
and U8622 (N_8622,N_8335,N_8460);
xor U8623 (N_8623,N_8443,N_8305);
or U8624 (N_8624,N_8451,N_8449);
and U8625 (N_8625,N_8393,N_8493);
xnor U8626 (N_8626,N_8283,N_8254);
and U8627 (N_8627,N_8287,N_8293);
and U8628 (N_8628,N_8401,N_8307);
xor U8629 (N_8629,N_8389,N_8252);
or U8630 (N_8630,N_8294,N_8431);
and U8631 (N_8631,N_8345,N_8266);
or U8632 (N_8632,N_8402,N_8290);
and U8633 (N_8633,N_8329,N_8460);
or U8634 (N_8634,N_8374,N_8417);
or U8635 (N_8635,N_8346,N_8267);
or U8636 (N_8636,N_8483,N_8336);
xor U8637 (N_8637,N_8377,N_8295);
nor U8638 (N_8638,N_8308,N_8451);
xnor U8639 (N_8639,N_8385,N_8403);
or U8640 (N_8640,N_8418,N_8435);
nand U8641 (N_8641,N_8423,N_8402);
or U8642 (N_8642,N_8322,N_8450);
or U8643 (N_8643,N_8279,N_8439);
or U8644 (N_8644,N_8465,N_8463);
nand U8645 (N_8645,N_8374,N_8351);
or U8646 (N_8646,N_8419,N_8298);
and U8647 (N_8647,N_8457,N_8327);
or U8648 (N_8648,N_8379,N_8377);
or U8649 (N_8649,N_8474,N_8252);
xor U8650 (N_8650,N_8486,N_8467);
xor U8651 (N_8651,N_8484,N_8312);
and U8652 (N_8652,N_8256,N_8327);
nand U8653 (N_8653,N_8342,N_8492);
or U8654 (N_8654,N_8364,N_8442);
or U8655 (N_8655,N_8465,N_8257);
and U8656 (N_8656,N_8260,N_8448);
nand U8657 (N_8657,N_8391,N_8263);
nand U8658 (N_8658,N_8358,N_8274);
nor U8659 (N_8659,N_8422,N_8438);
or U8660 (N_8660,N_8257,N_8269);
nor U8661 (N_8661,N_8449,N_8349);
or U8662 (N_8662,N_8456,N_8434);
or U8663 (N_8663,N_8359,N_8442);
xor U8664 (N_8664,N_8405,N_8465);
and U8665 (N_8665,N_8389,N_8353);
or U8666 (N_8666,N_8455,N_8316);
or U8667 (N_8667,N_8256,N_8267);
nand U8668 (N_8668,N_8379,N_8458);
and U8669 (N_8669,N_8473,N_8288);
xnor U8670 (N_8670,N_8429,N_8478);
and U8671 (N_8671,N_8388,N_8341);
nor U8672 (N_8672,N_8278,N_8477);
or U8673 (N_8673,N_8327,N_8302);
xor U8674 (N_8674,N_8455,N_8280);
xor U8675 (N_8675,N_8351,N_8364);
nand U8676 (N_8676,N_8399,N_8439);
and U8677 (N_8677,N_8279,N_8339);
xnor U8678 (N_8678,N_8478,N_8454);
and U8679 (N_8679,N_8332,N_8474);
nand U8680 (N_8680,N_8288,N_8497);
nor U8681 (N_8681,N_8440,N_8481);
xnor U8682 (N_8682,N_8417,N_8444);
nor U8683 (N_8683,N_8365,N_8440);
and U8684 (N_8684,N_8428,N_8324);
nor U8685 (N_8685,N_8451,N_8317);
nand U8686 (N_8686,N_8313,N_8354);
and U8687 (N_8687,N_8296,N_8277);
or U8688 (N_8688,N_8499,N_8377);
or U8689 (N_8689,N_8359,N_8449);
or U8690 (N_8690,N_8481,N_8323);
nand U8691 (N_8691,N_8295,N_8416);
nor U8692 (N_8692,N_8253,N_8382);
and U8693 (N_8693,N_8403,N_8388);
or U8694 (N_8694,N_8286,N_8443);
nor U8695 (N_8695,N_8287,N_8354);
nor U8696 (N_8696,N_8439,N_8333);
nor U8697 (N_8697,N_8393,N_8386);
nand U8698 (N_8698,N_8449,N_8496);
nor U8699 (N_8699,N_8263,N_8401);
nand U8700 (N_8700,N_8469,N_8426);
or U8701 (N_8701,N_8255,N_8432);
or U8702 (N_8702,N_8356,N_8322);
xnor U8703 (N_8703,N_8403,N_8278);
xnor U8704 (N_8704,N_8487,N_8361);
and U8705 (N_8705,N_8361,N_8311);
or U8706 (N_8706,N_8427,N_8443);
xnor U8707 (N_8707,N_8325,N_8400);
or U8708 (N_8708,N_8366,N_8288);
xor U8709 (N_8709,N_8475,N_8344);
and U8710 (N_8710,N_8486,N_8431);
xor U8711 (N_8711,N_8381,N_8275);
nand U8712 (N_8712,N_8474,N_8429);
nand U8713 (N_8713,N_8291,N_8423);
nor U8714 (N_8714,N_8336,N_8293);
or U8715 (N_8715,N_8495,N_8289);
or U8716 (N_8716,N_8419,N_8265);
and U8717 (N_8717,N_8487,N_8327);
xor U8718 (N_8718,N_8396,N_8420);
nand U8719 (N_8719,N_8392,N_8464);
and U8720 (N_8720,N_8279,N_8370);
or U8721 (N_8721,N_8358,N_8360);
nand U8722 (N_8722,N_8443,N_8287);
or U8723 (N_8723,N_8261,N_8438);
and U8724 (N_8724,N_8291,N_8383);
and U8725 (N_8725,N_8426,N_8441);
or U8726 (N_8726,N_8437,N_8402);
nor U8727 (N_8727,N_8272,N_8413);
nand U8728 (N_8728,N_8425,N_8264);
or U8729 (N_8729,N_8422,N_8316);
or U8730 (N_8730,N_8491,N_8259);
and U8731 (N_8731,N_8366,N_8303);
xor U8732 (N_8732,N_8469,N_8326);
xor U8733 (N_8733,N_8428,N_8469);
nor U8734 (N_8734,N_8377,N_8478);
nand U8735 (N_8735,N_8428,N_8401);
nand U8736 (N_8736,N_8359,N_8263);
or U8737 (N_8737,N_8354,N_8266);
or U8738 (N_8738,N_8408,N_8331);
or U8739 (N_8739,N_8274,N_8413);
or U8740 (N_8740,N_8268,N_8376);
or U8741 (N_8741,N_8301,N_8404);
nand U8742 (N_8742,N_8308,N_8363);
or U8743 (N_8743,N_8392,N_8260);
and U8744 (N_8744,N_8284,N_8409);
nand U8745 (N_8745,N_8274,N_8416);
nor U8746 (N_8746,N_8434,N_8343);
and U8747 (N_8747,N_8296,N_8436);
nor U8748 (N_8748,N_8276,N_8444);
or U8749 (N_8749,N_8349,N_8414);
or U8750 (N_8750,N_8671,N_8507);
xnor U8751 (N_8751,N_8593,N_8609);
nand U8752 (N_8752,N_8521,N_8512);
or U8753 (N_8753,N_8683,N_8705);
nor U8754 (N_8754,N_8649,N_8738);
nor U8755 (N_8755,N_8673,N_8713);
xnor U8756 (N_8756,N_8504,N_8742);
xnor U8757 (N_8757,N_8689,N_8720);
or U8758 (N_8758,N_8726,N_8582);
nand U8759 (N_8759,N_8623,N_8709);
nor U8760 (N_8760,N_8680,N_8694);
nand U8761 (N_8761,N_8578,N_8606);
nor U8762 (N_8762,N_8585,N_8640);
and U8763 (N_8763,N_8515,N_8668);
nor U8764 (N_8764,N_8723,N_8731);
or U8765 (N_8765,N_8711,N_8580);
or U8766 (N_8766,N_8641,N_8547);
or U8767 (N_8767,N_8610,N_8749);
and U8768 (N_8768,N_8612,N_8535);
nor U8769 (N_8769,N_8701,N_8599);
xor U8770 (N_8770,N_8747,N_8614);
nor U8771 (N_8771,N_8702,N_8618);
nor U8772 (N_8772,N_8716,N_8644);
nor U8773 (N_8773,N_8533,N_8532);
nand U8774 (N_8774,N_8707,N_8652);
nor U8775 (N_8775,N_8691,N_8621);
and U8776 (N_8776,N_8516,N_8660);
and U8777 (N_8777,N_8733,N_8522);
or U8778 (N_8778,N_8639,N_8546);
or U8779 (N_8779,N_8571,N_8717);
nor U8780 (N_8780,N_8622,N_8737);
xor U8781 (N_8781,N_8613,N_8527);
xnor U8782 (N_8782,N_8574,N_8589);
nand U8783 (N_8783,N_8645,N_8520);
nor U8784 (N_8784,N_8678,N_8509);
and U8785 (N_8785,N_8669,N_8583);
and U8786 (N_8786,N_8525,N_8595);
nor U8787 (N_8787,N_8604,N_8581);
xnor U8788 (N_8788,N_8727,N_8714);
and U8789 (N_8789,N_8562,N_8659);
nor U8790 (N_8790,N_8626,N_8696);
or U8791 (N_8791,N_8684,N_8576);
or U8792 (N_8792,N_8634,N_8569);
and U8793 (N_8793,N_8647,N_8545);
or U8794 (N_8794,N_8706,N_8698);
xnor U8795 (N_8795,N_8615,N_8724);
and U8796 (N_8796,N_8534,N_8558);
nand U8797 (N_8797,N_8503,N_8560);
nor U8798 (N_8798,N_8686,N_8566);
or U8799 (N_8799,N_8631,N_8564);
and U8800 (N_8800,N_8554,N_8537);
nand U8801 (N_8801,N_8551,N_8518);
and U8802 (N_8802,N_8514,N_8519);
or U8803 (N_8803,N_8510,N_8642);
or U8804 (N_8804,N_8744,N_8540);
or U8805 (N_8805,N_8570,N_8638);
and U8806 (N_8806,N_8529,N_8505);
nor U8807 (N_8807,N_8708,N_8693);
nor U8808 (N_8808,N_8557,N_8667);
and U8809 (N_8809,N_8601,N_8506);
xnor U8810 (N_8810,N_8665,N_8718);
or U8811 (N_8811,N_8555,N_8625);
nor U8812 (N_8812,N_8653,N_8677);
nor U8813 (N_8813,N_8685,N_8650);
and U8814 (N_8814,N_8501,N_8704);
nor U8815 (N_8815,N_8655,N_8648);
nand U8816 (N_8816,N_8633,N_8594);
nor U8817 (N_8817,N_8538,N_8591);
and U8818 (N_8818,N_8661,N_8695);
or U8819 (N_8819,N_8587,N_8736);
nand U8820 (N_8820,N_8561,N_8740);
or U8821 (N_8821,N_8681,N_8605);
or U8822 (N_8822,N_8703,N_8636);
and U8823 (N_8823,N_8692,N_8539);
xnor U8824 (N_8824,N_8656,N_8602);
nand U8825 (N_8825,N_8741,N_8628);
and U8826 (N_8826,N_8542,N_8635);
xor U8827 (N_8827,N_8600,N_8666);
or U8828 (N_8828,N_8586,N_8573);
nor U8829 (N_8829,N_8739,N_8597);
xor U8830 (N_8830,N_8528,N_8745);
or U8831 (N_8831,N_8556,N_8688);
nand U8832 (N_8832,N_8676,N_8632);
or U8833 (N_8833,N_8712,N_8577);
nor U8834 (N_8834,N_8729,N_8511);
and U8835 (N_8835,N_8603,N_8579);
nand U8836 (N_8836,N_8746,N_8710);
or U8837 (N_8837,N_8548,N_8624);
or U8838 (N_8838,N_8619,N_8721);
nand U8839 (N_8839,N_8517,N_8734);
and U8840 (N_8840,N_8531,N_8616);
xnor U8841 (N_8841,N_8743,N_8663);
or U8842 (N_8842,N_8552,N_8735);
or U8843 (N_8843,N_8617,N_8611);
nand U8844 (N_8844,N_8502,N_8620);
nor U8845 (N_8845,N_8662,N_8651);
or U8846 (N_8846,N_8563,N_8536);
xnor U8847 (N_8847,N_8584,N_8526);
xnor U8848 (N_8848,N_8544,N_8728);
and U8849 (N_8849,N_8699,N_8670);
or U8850 (N_8850,N_8657,N_8513);
or U8851 (N_8851,N_8572,N_8658);
nand U8852 (N_8852,N_8588,N_8700);
or U8853 (N_8853,N_8508,N_8565);
nand U8854 (N_8854,N_8500,N_8559);
and U8855 (N_8855,N_8541,N_8549);
xor U8856 (N_8856,N_8654,N_8715);
nor U8857 (N_8857,N_8608,N_8719);
xor U8858 (N_8858,N_8530,N_8598);
nand U8859 (N_8859,N_8629,N_8607);
nand U8860 (N_8860,N_8567,N_8697);
xnor U8861 (N_8861,N_8687,N_8590);
nor U8862 (N_8862,N_8553,N_8722);
nor U8863 (N_8863,N_8748,N_8646);
xnor U8864 (N_8864,N_8675,N_8732);
and U8865 (N_8865,N_8524,N_8592);
nor U8866 (N_8866,N_8725,N_8690);
or U8867 (N_8867,N_8637,N_8682);
xor U8868 (N_8868,N_8630,N_8543);
and U8869 (N_8869,N_8679,N_8664);
nand U8870 (N_8870,N_8674,N_8550);
nor U8871 (N_8871,N_8643,N_8730);
or U8872 (N_8872,N_8523,N_8627);
nor U8873 (N_8873,N_8568,N_8596);
xnor U8874 (N_8874,N_8575,N_8672);
xnor U8875 (N_8875,N_8546,N_8560);
xnor U8876 (N_8876,N_8591,N_8621);
nand U8877 (N_8877,N_8739,N_8630);
nor U8878 (N_8878,N_8570,N_8515);
and U8879 (N_8879,N_8735,N_8515);
xnor U8880 (N_8880,N_8634,N_8688);
nand U8881 (N_8881,N_8642,N_8530);
and U8882 (N_8882,N_8644,N_8597);
xor U8883 (N_8883,N_8653,N_8552);
or U8884 (N_8884,N_8728,N_8702);
and U8885 (N_8885,N_8583,N_8641);
or U8886 (N_8886,N_8515,N_8631);
or U8887 (N_8887,N_8635,N_8689);
nor U8888 (N_8888,N_8659,N_8701);
xor U8889 (N_8889,N_8530,N_8523);
nand U8890 (N_8890,N_8523,N_8564);
nand U8891 (N_8891,N_8525,N_8658);
nor U8892 (N_8892,N_8726,N_8711);
xor U8893 (N_8893,N_8635,N_8529);
or U8894 (N_8894,N_8684,N_8539);
xor U8895 (N_8895,N_8670,N_8734);
xnor U8896 (N_8896,N_8526,N_8599);
nor U8897 (N_8897,N_8563,N_8540);
nor U8898 (N_8898,N_8671,N_8578);
xor U8899 (N_8899,N_8703,N_8514);
or U8900 (N_8900,N_8669,N_8540);
nand U8901 (N_8901,N_8539,N_8634);
nor U8902 (N_8902,N_8511,N_8524);
or U8903 (N_8903,N_8715,N_8690);
xnor U8904 (N_8904,N_8573,N_8538);
nand U8905 (N_8905,N_8677,N_8509);
nor U8906 (N_8906,N_8526,N_8672);
and U8907 (N_8907,N_8708,N_8566);
nor U8908 (N_8908,N_8698,N_8586);
or U8909 (N_8909,N_8566,N_8537);
and U8910 (N_8910,N_8605,N_8592);
xnor U8911 (N_8911,N_8501,N_8664);
xor U8912 (N_8912,N_8611,N_8728);
or U8913 (N_8913,N_8556,N_8594);
nor U8914 (N_8914,N_8656,N_8743);
xor U8915 (N_8915,N_8577,N_8568);
or U8916 (N_8916,N_8641,N_8573);
xor U8917 (N_8917,N_8578,N_8501);
xor U8918 (N_8918,N_8551,N_8535);
xnor U8919 (N_8919,N_8704,N_8508);
xnor U8920 (N_8920,N_8748,N_8525);
nand U8921 (N_8921,N_8732,N_8552);
nor U8922 (N_8922,N_8662,N_8507);
xor U8923 (N_8923,N_8500,N_8532);
or U8924 (N_8924,N_8737,N_8540);
and U8925 (N_8925,N_8612,N_8593);
or U8926 (N_8926,N_8734,N_8723);
xor U8927 (N_8927,N_8530,N_8718);
xor U8928 (N_8928,N_8645,N_8534);
nand U8929 (N_8929,N_8747,N_8672);
nor U8930 (N_8930,N_8670,N_8652);
xor U8931 (N_8931,N_8727,N_8512);
or U8932 (N_8932,N_8660,N_8636);
and U8933 (N_8933,N_8672,N_8610);
or U8934 (N_8934,N_8569,N_8576);
xor U8935 (N_8935,N_8635,N_8735);
xor U8936 (N_8936,N_8558,N_8717);
or U8937 (N_8937,N_8629,N_8558);
and U8938 (N_8938,N_8664,N_8720);
xor U8939 (N_8939,N_8504,N_8668);
or U8940 (N_8940,N_8620,N_8721);
nand U8941 (N_8941,N_8603,N_8738);
or U8942 (N_8942,N_8514,N_8504);
xor U8943 (N_8943,N_8701,N_8549);
or U8944 (N_8944,N_8592,N_8631);
nand U8945 (N_8945,N_8643,N_8516);
nor U8946 (N_8946,N_8551,N_8706);
nor U8947 (N_8947,N_8503,N_8618);
nor U8948 (N_8948,N_8717,N_8744);
or U8949 (N_8949,N_8534,N_8741);
or U8950 (N_8950,N_8515,N_8613);
or U8951 (N_8951,N_8512,N_8559);
nor U8952 (N_8952,N_8728,N_8739);
xnor U8953 (N_8953,N_8718,N_8504);
or U8954 (N_8954,N_8600,N_8715);
nor U8955 (N_8955,N_8692,N_8723);
and U8956 (N_8956,N_8736,N_8555);
and U8957 (N_8957,N_8646,N_8674);
xor U8958 (N_8958,N_8747,N_8642);
nor U8959 (N_8959,N_8682,N_8618);
and U8960 (N_8960,N_8611,N_8510);
nand U8961 (N_8961,N_8699,N_8609);
and U8962 (N_8962,N_8508,N_8509);
xor U8963 (N_8963,N_8718,N_8720);
nand U8964 (N_8964,N_8671,N_8595);
nand U8965 (N_8965,N_8584,N_8708);
nand U8966 (N_8966,N_8704,N_8535);
nand U8967 (N_8967,N_8645,N_8727);
nor U8968 (N_8968,N_8611,N_8603);
nor U8969 (N_8969,N_8563,N_8531);
nand U8970 (N_8970,N_8588,N_8585);
nor U8971 (N_8971,N_8508,N_8649);
xor U8972 (N_8972,N_8616,N_8610);
xnor U8973 (N_8973,N_8683,N_8563);
xor U8974 (N_8974,N_8725,N_8528);
nand U8975 (N_8975,N_8718,N_8545);
and U8976 (N_8976,N_8721,N_8635);
nand U8977 (N_8977,N_8670,N_8629);
nand U8978 (N_8978,N_8613,N_8598);
nor U8979 (N_8979,N_8546,N_8553);
nand U8980 (N_8980,N_8690,N_8682);
xor U8981 (N_8981,N_8745,N_8727);
or U8982 (N_8982,N_8720,N_8642);
nor U8983 (N_8983,N_8720,N_8731);
xnor U8984 (N_8984,N_8504,N_8575);
xnor U8985 (N_8985,N_8722,N_8687);
xor U8986 (N_8986,N_8592,N_8701);
and U8987 (N_8987,N_8687,N_8583);
xnor U8988 (N_8988,N_8680,N_8678);
or U8989 (N_8989,N_8665,N_8691);
or U8990 (N_8990,N_8616,N_8535);
nor U8991 (N_8991,N_8717,N_8693);
and U8992 (N_8992,N_8639,N_8700);
nand U8993 (N_8993,N_8657,N_8563);
or U8994 (N_8994,N_8730,N_8686);
nor U8995 (N_8995,N_8528,N_8537);
xor U8996 (N_8996,N_8712,N_8550);
nor U8997 (N_8997,N_8694,N_8633);
and U8998 (N_8998,N_8537,N_8585);
or U8999 (N_8999,N_8718,N_8683);
and U9000 (N_9000,N_8960,N_8979);
nand U9001 (N_9001,N_8840,N_8919);
nand U9002 (N_9002,N_8957,N_8874);
xor U9003 (N_9003,N_8969,N_8879);
or U9004 (N_9004,N_8811,N_8793);
xnor U9005 (N_9005,N_8931,N_8906);
or U9006 (N_9006,N_8910,N_8984);
nor U9007 (N_9007,N_8948,N_8917);
nand U9008 (N_9008,N_8780,N_8781);
nor U9009 (N_9009,N_8928,N_8756);
nand U9010 (N_9010,N_8823,N_8998);
nand U9011 (N_9011,N_8849,N_8880);
nand U9012 (N_9012,N_8930,N_8888);
or U9013 (N_9013,N_8959,N_8981);
nor U9014 (N_9014,N_8853,N_8895);
nor U9015 (N_9015,N_8947,N_8800);
nor U9016 (N_9016,N_8950,N_8873);
nand U9017 (N_9017,N_8905,N_8783);
xor U9018 (N_9018,N_8819,N_8884);
and U9019 (N_9019,N_8820,N_8878);
nor U9020 (N_9020,N_8903,N_8914);
nor U9021 (N_9021,N_8958,N_8806);
and U9022 (N_9022,N_8864,N_8992);
or U9023 (N_9023,N_8834,N_8771);
nor U9024 (N_9024,N_8752,N_8773);
nand U9025 (N_9025,N_8900,N_8818);
nor U9026 (N_9026,N_8893,N_8927);
or U9027 (N_9027,N_8935,N_8760);
xor U9028 (N_9028,N_8908,N_8824);
and U9029 (N_9029,N_8922,N_8925);
xor U9030 (N_9030,N_8942,N_8988);
nand U9031 (N_9031,N_8858,N_8938);
xnor U9032 (N_9032,N_8945,N_8837);
nand U9033 (N_9033,N_8937,N_8758);
xnor U9034 (N_9034,N_8841,N_8923);
nor U9035 (N_9035,N_8932,N_8795);
and U9036 (N_9036,N_8851,N_8902);
nand U9037 (N_9037,N_8882,N_8828);
and U9038 (N_9038,N_8845,N_8926);
xor U9039 (N_9039,N_8993,N_8863);
nor U9040 (N_9040,N_8813,N_8843);
nor U9041 (N_9041,N_8775,N_8815);
and U9042 (N_9042,N_8904,N_8989);
or U9043 (N_9043,N_8964,N_8861);
xnor U9044 (N_9044,N_8929,N_8894);
or U9045 (N_9045,N_8850,N_8751);
nor U9046 (N_9046,N_8953,N_8844);
xnor U9047 (N_9047,N_8933,N_8961);
nand U9048 (N_9048,N_8791,N_8808);
nor U9049 (N_9049,N_8867,N_8829);
nand U9050 (N_9050,N_8899,N_8831);
nand U9051 (N_9051,N_8772,N_8870);
or U9052 (N_9052,N_8762,N_8881);
or U9053 (N_9053,N_8936,N_8782);
and U9054 (N_9054,N_8860,N_8750);
xnor U9055 (N_9055,N_8779,N_8842);
or U9056 (N_9056,N_8798,N_8921);
xor U9057 (N_9057,N_8912,N_8934);
or U9058 (N_9058,N_8866,N_8803);
or U9059 (N_9059,N_8761,N_8913);
xor U9060 (N_9060,N_8941,N_8862);
nor U9061 (N_9061,N_8901,N_8907);
nor U9062 (N_9062,N_8986,N_8794);
and U9063 (N_9063,N_8802,N_8789);
and U9064 (N_9064,N_8943,N_8892);
and U9065 (N_9065,N_8816,N_8804);
or U9066 (N_9066,N_8786,N_8757);
nor U9067 (N_9067,N_8963,N_8763);
nor U9068 (N_9068,N_8974,N_8826);
or U9069 (N_9069,N_8952,N_8918);
nor U9070 (N_9070,N_8975,N_8822);
and U9071 (N_9071,N_8890,N_8753);
nor U9072 (N_9072,N_8944,N_8769);
xnor U9073 (N_9073,N_8848,N_8896);
xnor U9074 (N_9074,N_8877,N_8871);
nor U9075 (N_9075,N_8774,N_8911);
xnor U9076 (N_9076,N_8856,N_8833);
and U9077 (N_9077,N_8970,N_8966);
and U9078 (N_9078,N_8859,N_8865);
or U9079 (N_9079,N_8857,N_8836);
nand U9080 (N_9080,N_8799,N_8814);
or U9081 (N_9081,N_8968,N_8962);
or U9082 (N_9082,N_8990,N_8886);
nand U9083 (N_9083,N_8994,N_8770);
and U9084 (N_9084,N_8830,N_8764);
nor U9085 (N_9085,N_8790,N_8939);
xnor U9086 (N_9086,N_8792,N_8805);
or U9087 (N_9087,N_8885,N_8976);
nor U9088 (N_9088,N_8983,N_8765);
or U9089 (N_9089,N_8997,N_8973);
nor U9090 (N_9090,N_8995,N_8991);
nand U9091 (N_9091,N_8915,N_8787);
nor U9092 (N_9092,N_8784,N_8827);
nand U9093 (N_9093,N_8839,N_8982);
nor U9094 (N_9094,N_8891,N_8872);
xor U9095 (N_9095,N_8797,N_8889);
and U9096 (N_9096,N_8951,N_8846);
or U9097 (N_9097,N_8766,N_8817);
xor U9098 (N_9098,N_8898,N_8999);
nand U9099 (N_9099,N_8847,N_8977);
nand U9100 (N_9100,N_8909,N_8996);
nand U9101 (N_9101,N_8809,N_8949);
and U9102 (N_9102,N_8776,N_8876);
nand U9103 (N_9103,N_8924,N_8778);
and U9104 (N_9104,N_8854,N_8883);
or U9105 (N_9105,N_8887,N_8920);
or U9106 (N_9106,N_8955,N_8852);
or U9107 (N_9107,N_8777,N_8875);
xnor U9108 (N_9108,N_8972,N_8855);
or U9109 (N_9109,N_8868,N_8946);
nand U9110 (N_9110,N_8940,N_8812);
or U9111 (N_9111,N_8788,N_8987);
or U9112 (N_9112,N_8967,N_8954);
nor U9113 (N_9113,N_8807,N_8835);
or U9114 (N_9114,N_8755,N_8838);
xor U9115 (N_9115,N_8810,N_8801);
nand U9116 (N_9116,N_8825,N_8767);
and U9117 (N_9117,N_8897,N_8796);
nand U9118 (N_9118,N_8768,N_8832);
or U9119 (N_9119,N_8978,N_8785);
and U9120 (N_9120,N_8985,N_8916);
or U9121 (N_9121,N_8971,N_8980);
and U9122 (N_9122,N_8965,N_8759);
xnor U9123 (N_9123,N_8869,N_8821);
or U9124 (N_9124,N_8754,N_8956);
xor U9125 (N_9125,N_8916,N_8927);
and U9126 (N_9126,N_8885,N_8988);
xor U9127 (N_9127,N_8792,N_8879);
nand U9128 (N_9128,N_8872,N_8761);
nor U9129 (N_9129,N_8914,N_8820);
xor U9130 (N_9130,N_8905,N_8841);
nor U9131 (N_9131,N_8844,N_8987);
nand U9132 (N_9132,N_8849,N_8824);
or U9133 (N_9133,N_8975,N_8850);
xor U9134 (N_9134,N_8960,N_8902);
xnor U9135 (N_9135,N_8876,N_8868);
nor U9136 (N_9136,N_8950,N_8808);
nor U9137 (N_9137,N_8963,N_8846);
xnor U9138 (N_9138,N_8754,N_8791);
or U9139 (N_9139,N_8947,N_8955);
xnor U9140 (N_9140,N_8885,N_8894);
xnor U9141 (N_9141,N_8850,N_8923);
or U9142 (N_9142,N_8781,N_8794);
nand U9143 (N_9143,N_8983,N_8833);
or U9144 (N_9144,N_8791,N_8855);
and U9145 (N_9145,N_8864,N_8760);
nand U9146 (N_9146,N_8750,N_8977);
and U9147 (N_9147,N_8830,N_8783);
xor U9148 (N_9148,N_8954,N_8766);
xnor U9149 (N_9149,N_8965,N_8982);
xnor U9150 (N_9150,N_8846,N_8757);
xor U9151 (N_9151,N_8804,N_8810);
nor U9152 (N_9152,N_8850,N_8849);
nor U9153 (N_9153,N_8778,N_8873);
nor U9154 (N_9154,N_8822,N_8777);
nand U9155 (N_9155,N_8760,N_8776);
nand U9156 (N_9156,N_8960,N_8905);
nor U9157 (N_9157,N_8980,N_8880);
nand U9158 (N_9158,N_8757,N_8887);
or U9159 (N_9159,N_8783,N_8827);
nand U9160 (N_9160,N_8751,N_8757);
nand U9161 (N_9161,N_8899,N_8838);
or U9162 (N_9162,N_8870,N_8794);
nor U9163 (N_9163,N_8799,N_8831);
xor U9164 (N_9164,N_8846,N_8785);
or U9165 (N_9165,N_8895,N_8792);
nor U9166 (N_9166,N_8911,N_8778);
or U9167 (N_9167,N_8854,N_8798);
or U9168 (N_9168,N_8761,N_8882);
nor U9169 (N_9169,N_8857,N_8860);
and U9170 (N_9170,N_8907,N_8963);
nor U9171 (N_9171,N_8755,N_8985);
or U9172 (N_9172,N_8922,N_8799);
xor U9173 (N_9173,N_8867,N_8788);
or U9174 (N_9174,N_8993,N_8763);
and U9175 (N_9175,N_8837,N_8933);
nor U9176 (N_9176,N_8864,N_8918);
xor U9177 (N_9177,N_8988,N_8751);
xnor U9178 (N_9178,N_8813,N_8999);
and U9179 (N_9179,N_8792,N_8788);
nand U9180 (N_9180,N_8782,N_8824);
and U9181 (N_9181,N_8913,N_8932);
nand U9182 (N_9182,N_8828,N_8957);
nor U9183 (N_9183,N_8897,N_8977);
nand U9184 (N_9184,N_8992,N_8917);
or U9185 (N_9185,N_8824,N_8963);
nor U9186 (N_9186,N_8857,N_8829);
nor U9187 (N_9187,N_8845,N_8905);
and U9188 (N_9188,N_8793,N_8858);
nor U9189 (N_9189,N_8940,N_8844);
nor U9190 (N_9190,N_8856,N_8766);
nand U9191 (N_9191,N_8816,N_8959);
or U9192 (N_9192,N_8851,N_8983);
xnor U9193 (N_9193,N_8952,N_8914);
nor U9194 (N_9194,N_8899,N_8812);
xnor U9195 (N_9195,N_8908,N_8954);
or U9196 (N_9196,N_8995,N_8812);
xnor U9197 (N_9197,N_8831,N_8863);
and U9198 (N_9198,N_8794,N_8933);
xor U9199 (N_9199,N_8968,N_8839);
or U9200 (N_9200,N_8845,N_8779);
or U9201 (N_9201,N_8755,N_8990);
xor U9202 (N_9202,N_8989,N_8950);
xnor U9203 (N_9203,N_8972,N_8812);
nor U9204 (N_9204,N_8833,N_8750);
and U9205 (N_9205,N_8871,N_8787);
or U9206 (N_9206,N_8956,N_8906);
nand U9207 (N_9207,N_8898,N_8794);
xor U9208 (N_9208,N_8798,N_8783);
nor U9209 (N_9209,N_8938,N_8804);
and U9210 (N_9210,N_8824,N_8911);
nor U9211 (N_9211,N_8895,N_8774);
xor U9212 (N_9212,N_8972,N_8768);
nand U9213 (N_9213,N_8826,N_8768);
and U9214 (N_9214,N_8906,N_8839);
xor U9215 (N_9215,N_8850,N_8991);
xor U9216 (N_9216,N_8886,N_8829);
or U9217 (N_9217,N_8838,N_8920);
xnor U9218 (N_9218,N_8965,N_8894);
nand U9219 (N_9219,N_8976,N_8929);
nand U9220 (N_9220,N_8860,N_8951);
or U9221 (N_9221,N_8770,N_8817);
nand U9222 (N_9222,N_8773,N_8950);
nand U9223 (N_9223,N_8922,N_8975);
nor U9224 (N_9224,N_8795,N_8870);
and U9225 (N_9225,N_8847,N_8995);
nor U9226 (N_9226,N_8877,N_8754);
nor U9227 (N_9227,N_8923,N_8772);
and U9228 (N_9228,N_8846,N_8993);
or U9229 (N_9229,N_8787,N_8870);
nand U9230 (N_9230,N_8937,N_8993);
or U9231 (N_9231,N_8899,N_8806);
and U9232 (N_9232,N_8829,N_8865);
xor U9233 (N_9233,N_8803,N_8857);
or U9234 (N_9234,N_8773,N_8915);
xor U9235 (N_9235,N_8970,N_8793);
and U9236 (N_9236,N_8819,N_8805);
nor U9237 (N_9237,N_8893,N_8750);
and U9238 (N_9238,N_8896,N_8943);
or U9239 (N_9239,N_8943,N_8993);
nor U9240 (N_9240,N_8779,N_8839);
and U9241 (N_9241,N_8965,N_8775);
or U9242 (N_9242,N_8782,N_8842);
nor U9243 (N_9243,N_8933,N_8856);
xor U9244 (N_9244,N_8858,N_8999);
or U9245 (N_9245,N_8872,N_8847);
xnor U9246 (N_9246,N_8899,N_8822);
and U9247 (N_9247,N_8774,N_8822);
nor U9248 (N_9248,N_8793,N_8952);
xnor U9249 (N_9249,N_8808,N_8752);
or U9250 (N_9250,N_9171,N_9072);
or U9251 (N_9251,N_9211,N_9141);
nor U9252 (N_9252,N_9239,N_9125);
nor U9253 (N_9253,N_9126,N_9229);
nor U9254 (N_9254,N_9187,N_9087);
and U9255 (N_9255,N_9085,N_9051);
and U9256 (N_9256,N_9216,N_9226);
nand U9257 (N_9257,N_9227,N_9071);
and U9258 (N_9258,N_9246,N_9102);
nand U9259 (N_9259,N_9215,N_9005);
xnor U9260 (N_9260,N_9219,N_9164);
nand U9261 (N_9261,N_9017,N_9243);
and U9262 (N_9262,N_9007,N_9237);
xnor U9263 (N_9263,N_9185,N_9058);
nand U9264 (N_9264,N_9070,N_9065);
nor U9265 (N_9265,N_9184,N_9146);
nand U9266 (N_9266,N_9041,N_9175);
nor U9267 (N_9267,N_9116,N_9046);
or U9268 (N_9268,N_9090,N_9201);
xor U9269 (N_9269,N_9242,N_9173);
xor U9270 (N_9270,N_9180,N_9160);
nand U9271 (N_9271,N_9142,N_9018);
xnor U9272 (N_9272,N_9131,N_9095);
nand U9273 (N_9273,N_9044,N_9148);
nand U9274 (N_9274,N_9213,N_9040);
xor U9275 (N_9275,N_9078,N_9038);
and U9276 (N_9276,N_9117,N_9106);
or U9277 (N_9277,N_9129,N_9054);
nor U9278 (N_9278,N_9144,N_9120);
and U9279 (N_9279,N_9168,N_9154);
nand U9280 (N_9280,N_9205,N_9064);
and U9281 (N_9281,N_9199,N_9019);
and U9282 (N_9282,N_9084,N_9220);
or U9283 (N_9283,N_9133,N_9190);
nor U9284 (N_9284,N_9032,N_9218);
or U9285 (N_9285,N_9152,N_9158);
and U9286 (N_9286,N_9088,N_9143);
or U9287 (N_9287,N_9021,N_9127);
nor U9288 (N_9288,N_9022,N_9138);
xor U9289 (N_9289,N_9162,N_9189);
nand U9290 (N_9290,N_9204,N_9115);
and U9291 (N_9291,N_9196,N_9140);
nor U9292 (N_9292,N_9155,N_9092);
and U9293 (N_9293,N_9156,N_9006);
nor U9294 (N_9294,N_9232,N_9212);
or U9295 (N_9295,N_9027,N_9030);
nor U9296 (N_9296,N_9012,N_9100);
nand U9297 (N_9297,N_9009,N_9233);
or U9298 (N_9298,N_9104,N_9014);
nor U9299 (N_9299,N_9101,N_9248);
nand U9300 (N_9300,N_9025,N_9222);
nor U9301 (N_9301,N_9136,N_9034);
nand U9302 (N_9302,N_9134,N_9228);
and U9303 (N_9303,N_9119,N_9214);
and U9304 (N_9304,N_9057,N_9153);
and U9305 (N_9305,N_9235,N_9209);
and U9306 (N_9306,N_9003,N_9109);
nand U9307 (N_9307,N_9182,N_9050);
xnor U9308 (N_9308,N_9198,N_9193);
or U9309 (N_9309,N_9161,N_9128);
xnor U9310 (N_9310,N_9147,N_9091);
or U9311 (N_9311,N_9063,N_9149);
xnor U9312 (N_9312,N_9067,N_9062);
and U9313 (N_9313,N_9011,N_9016);
nand U9314 (N_9314,N_9124,N_9112);
nor U9315 (N_9315,N_9086,N_9165);
and U9316 (N_9316,N_9080,N_9004);
xor U9317 (N_9317,N_9197,N_9111);
nand U9318 (N_9318,N_9183,N_9000);
and U9319 (N_9319,N_9052,N_9172);
xnor U9320 (N_9320,N_9047,N_9028);
and U9321 (N_9321,N_9029,N_9073);
xor U9322 (N_9322,N_9236,N_9123);
nor U9323 (N_9323,N_9039,N_9079);
nand U9324 (N_9324,N_9001,N_9135);
xnor U9325 (N_9325,N_9075,N_9181);
xnor U9326 (N_9326,N_9176,N_9060);
or U9327 (N_9327,N_9178,N_9169);
nand U9328 (N_9328,N_9230,N_9093);
nor U9329 (N_9329,N_9094,N_9240);
xor U9330 (N_9330,N_9068,N_9174);
xor U9331 (N_9331,N_9121,N_9200);
and U9332 (N_9332,N_9048,N_9056);
nor U9333 (N_9333,N_9122,N_9188);
and U9334 (N_9334,N_9217,N_9043);
or U9335 (N_9335,N_9231,N_9145);
or U9336 (N_9336,N_9234,N_9108);
nor U9337 (N_9337,N_9024,N_9049);
and U9338 (N_9338,N_9035,N_9077);
and U9339 (N_9339,N_9076,N_9081);
or U9340 (N_9340,N_9033,N_9066);
nor U9341 (N_9341,N_9244,N_9074);
nor U9342 (N_9342,N_9191,N_9008);
and U9343 (N_9343,N_9241,N_9036);
nor U9344 (N_9344,N_9118,N_9026);
nand U9345 (N_9345,N_9031,N_9113);
and U9346 (N_9346,N_9042,N_9015);
nand U9347 (N_9347,N_9208,N_9249);
xor U9348 (N_9348,N_9107,N_9099);
or U9349 (N_9349,N_9096,N_9195);
nand U9350 (N_9350,N_9202,N_9045);
and U9351 (N_9351,N_9139,N_9069);
and U9352 (N_9352,N_9223,N_9137);
nand U9353 (N_9353,N_9192,N_9194);
xor U9354 (N_9354,N_9103,N_9132);
and U9355 (N_9355,N_9157,N_9166);
and U9356 (N_9356,N_9224,N_9053);
and U9357 (N_9357,N_9114,N_9177);
or U9358 (N_9358,N_9206,N_9020);
and U9359 (N_9359,N_9105,N_9013);
or U9360 (N_9360,N_9159,N_9059);
nand U9361 (N_9361,N_9179,N_9150);
and U9362 (N_9362,N_9151,N_9002);
or U9363 (N_9363,N_9167,N_9061);
nand U9364 (N_9364,N_9082,N_9083);
xnor U9365 (N_9365,N_9225,N_9089);
nor U9366 (N_9366,N_9110,N_9221);
or U9367 (N_9367,N_9238,N_9170);
xor U9368 (N_9368,N_9163,N_9247);
and U9369 (N_9369,N_9207,N_9097);
xnor U9370 (N_9370,N_9130,N_9186);
or U9371 (N_9371,N_9010,N_9023);
and U9372 (N_9372,N_9203,N_9055);
and U9373 (N_9373,N_9037,N_9245);
and U9374 (N_9374,N_9098,N_9210);
nor U9375 (N_9375,N_9138,N_9241);
xnor U9376 (N_9376,N_9082,N_9218);
xor U9377 (N_9377,N_9038,N_9109);
or U9378 (N_9378,N_9028,N_9185);
and U9379 (N_9379,N_9001,N_9115);
xor U9380 (N_9380,N_9043,N_9223);
nor U9381 (N_9381,N_9130,N_9082);
xnor U9382 (N_9382,N_9189,N_9047);
or U9383 (N_9383,N_9189,N_9027);
or U9384 (N_9384,N_9043,N_9212);
nor U9385 (N_9385,N_9146,N_9173);
and U9386 (N_9386,N_9248,N_9038);
xor U9387 (N_9387,N_9057,N_9178);
nand U9388 (N_9388,N_9152,N_9025);
xnor U9389 (N_9389,N_9100,N_9217);
nand U9390 (N_9390,N_9184,N_9073);
and U9391 (N_9391,N_9177,N_9049);
nor U9392 (N_9392,N_9038,N_9066);
nor U9393 (N_9393,N_9165,N_9170);
or U9394 (N_9394,N_9218,N_9085);
or U9395 (N_9395,N_9155,N_9117);
nand U9396 (N_9396,N_9098,N_9165);
nand U9397 (N_9397,N_9055,N_9187);
xor U9398 (N_9398,N_9100,N_9161);
xor U9399 (N_9399,N_9184,N_9148);
or U9400 (N_9400,N_9231,N_9121);
or U9401 (N_9401,N_9230,N_9073);
xnor U9402 (N_9402,N_9021,N_9057);
nor U9403 (N_9403,N_9163,N_9211);
and U9404 (N_9404,N_9160,N_9145);
or U9405 (N_9405,N_9140,N_9143);
nand U9406 (N_9406,N_9224,N_9110);
nand U9407 (N_9407,N_9180,N_9052);
nor U9408 (N_9408,N_9121,N_9232);
and U9409 (N_9409,N_9063,N_9222);
or U9410 (N_9410,N_9037,N_9177);
or U9411 (N_9411,N_9146,N_9218);
or U9412 (N_9412,N_9012,N_9082);
nand U9413 (N_9413,N_9017,N_9177);
nor U9414 (N_9414,N_9064,N_9147);
and U9415 (N_9415,N_9109,N_9010);
nor U9416 (N_9416,N_9023,N_9146);
nand U9417 (N_9417,N_9094,N_9067);
or U9418 (N_9418,N_9171,N_9168);
nor U9419 (N_9419,N_9186,N_9231);
nor U9420 (N_9420,N_9182,N_9141);
nand U9421 (N_9421,N_9141,N_9049);
or U9422 (N_9422,N_9176,N_9148);
and U9423 (N_9423,N_9167,N_9022);
or U9424 (N_9424,N_9173,N_9108);
xnor U9425 (N_9425,N_9192,N_9238);
nor U9426 (N_9426,N_9112,N_9032);
nor U9427 (N_9427,N_9101,N_9034);
or U9428 (N_9428,N_9109,N_9122);
or U9429 (N_9429,N_9097,N_9211);
xor U9430 (N_9430,N_9048,N_9094);
nor U9431 (N_9431,N_9024,N_9202);
nor U9432 (N_9432,N_9219,N_9158);
and U9433 (N_9433,N_9068,N_9026);
xnor U9434 (N_9434,N_9112,N_9013);
or U9435 (N_9435,N_9011,N_9066);
xnor U9436 (N_9436,N_9054,N_9099);
and U9437 (N_9437,N_9228,N_9096);
xnor U9438 (N_9438,N_9063,N_9111);
nor U9439 (N_9439,N_9142,N_9049);
or U9440 (N_9440,N_9226,N_9052);
nor U9441 (N_9441,N_9193,N_9015);
or U9442 (N_9442,N_9188,N_9149);
and U9443 (N_9443,N_9035,N_9056);
nor U9444 (N_9444,N_9045,N_9150);
nand U9445 (N_9445,N_9211,N_9022);
nor U9446 (N_9446,N_9211,N_9110);
and U9447 (N_9447,N_9012,N_9061);
nor U9448 (N_9448,N_9174,N_9145);
xnor U9449 (N_9449,N_9086,N_9232);
or U9450 (N_9450,N_9032,N_9015);
nor U9451 (N_9451,N_9164,N_9006);
nand U9452 (N_9452,N_9184,N_9239);
nor U9453 (N_9453,N_9064,N_9160);
nor U9454 (N_9454,N_9185,N_9206);
nor U9455 (N_9455,N_9116,N_9108);
xor U9456 (N_9456,N_9222,N_9245);
xnor U9457 (N_9457,N_9064,N_9159);
nand U9458 (N_9458,N_9182,N_9092);
and U9459 (N_9459,N_9213,N_9177);
and U9460 (N_9460,N_9222,N_9158);
or U9461 (N_9461,N_9190,N_9051);
xor U9462 (N_9462,N_9044,N_9147);
nor U9463 (N_9463,N_9223,N_9080);
or U9464 (N_9464,N_9062,N_9039);
xor U9465 (N_9465,N_9181,N_9053);
xor U9466 (N_9466,N_9187,N_9067);
or U9467 (N_9467,N_9166,N_9227);
or U9468 (N_9468,N_9145,N_9019);
xnor U9469 (N_9469,N_9087,N_9249);
and U9470 (N_9470,N_9186,N_9048);
xor U9471 (N_9471,N_9068,N_9008);
nor U9472 (N_9472,N_9155,N_9050);
nand U9473 (N_9473,N_9206,N_9029);
nand U9474 (N_9474,N_9198,N_9117);
xor U9475 (N_9475,N_9125,N_9027);
xor U9476 (N_9476,N_9238,N_9030);
xnor U9477 (N_9477,N_9205,N_9170);
and U9478 (N_9478,N_9130,N_9108);
or U9479 (N_9479,N_9172,N_9199);
nand U9480 (N_9480,N_9128,N_9164);
nor U9481 (N_9481,N_9139,N_9128);
nor U9482 (N_9482,N_9217,N_9238);
or U9483 (N_9483,N_9067,N_9124);
or U9484 (N_9484,N_9162,N_9167);
nand U9485 (N_9485,N_9062,N_9111);
xnor U9486 (N_9486,N_9103,N_9073);
nand U9487 (N_9487,N_9092,N_9226);
or U9488 (N_9488,N_9226,N_9158);
nor U9489 (N_9489,N_9109,N_9039);
xnor U9490 (N_9490,N_9115,N_9065);
nand U9491 (N_9491,N_9026,N_9206);
nor U9492 (N_9492,N_9246,N_9178);
xnor U9493 (N_9493,N_9143,N_9106);
nand U9494 (N_9494,N_9080,N_9063);
and U9495 (N_9495,N_9138,N_9183);
xnor U9496 (N_9496,N_9046,N_9043);
nand U9497 (N_9497,N_9220,N_9052);
nand U9498 (N_9498,N_9116,N_9129);
nand U9499 (N_9499,N_9071,N_9180);
and U9500 (N_9500,N_9268,N_9496);
nand U9501 (N_9501,N_9338,N_9300);
and U9502 (N_9502,N_9307,N_9330);
or U9503 (N_9503,N_9255,N_9295);
and U9504 (N_9504,N_9408,N_9264);
and U9505 (N_9505,N_9350,N_9400);
or U9506 (N_9506,N_9263,N_9390);
nor U9507 (N_9507,N_9477,N_9323);
and U9508 (N_9508,N_9495,N_9283);
nor U9509 (N_9509,N_9388,N_9416);
or U9510 (N_9510,N_9250,N_9449);
nand U9511 (N_9511,N_9378,N_9393);
or U9512 (N_9512,N_9498,N_9485);
or U9513 (N_9513,N_9431,N_9309);
or U9514 (N_9514,N_9404,N_9442);
xor U9515 (N_9515,N_9341,N_9468);
nand U9516 (N_9516,N_9418,N_9474);
nor U9517 (N_9517,N_9412,N_9486);
nor U9518 (N_9518,N_9406,N_9292);
nand U9519 (N_9519,N_9277,N_9335);
and U9520 (N_9520,N_9458,N_9274);
or U9521 (N_9521,N_9415,N_9376);
nand U9522 (N_9522,N_9320,N_9435);
and U9523 (N_9523,N_9297,N_9301);
or U9524 (N_9524,N_9384,N_9351);
xnor U9525 (N_9525,N_9342,N_9251);
xnor U9526 (N_9526,N_9348,N_9352);
nand U9527 (N_9527,N_9327,N_9271);
or U9528 (N_9528,N_9355,N_9401);
or U9529 (N_9529,N_9332,N_9482);
nor U9530 (N_9530,N_9366,N_9334);
or U9531 (N_9531,N_9325,N_9278);
and U9532 (N_9532,N_9360,N_9481);
nor U9533 (N_9533,N_9361,N_9272);
or U9534 (N_9534,N_9319,N_9454);
nand U9535 (N_9535,N_9463,N_9261);
nand U9536 (N_9536,N_9398,N_9354);
or U9537 (N_9537,N_9318,N_9465);
nand U9538 (N_9538,N_9279,N_9281);
nor U9539 (N_9539,N_9441,N_9254);
nand U9540 (N_9540,N_9467,N_9275);
or U9541 (N_9541,N_9356,N_9430);
nor U9542 (N_9542,N_9464,N_9294);
xnor U9543 (N_9543,N_9417,N_9440);
nand U9544 (N_9544,N_9284,N_9296);
nor U9545 (N_9545,N_9450,N_9478);
nand U9546 (N_9546,N_9276,N_9339);
nor U9547 (N_9547,N_9266,N_9453);
xor U9548 (N_9548,N_9490,N_9291);
and U9549 (N_9549,N_9428,N_9422);
nor U9550 (N_9550,N_9448,N_9475);
nand U9551 (N_9551,N_9363,N_9405);
or U9552 (N_9552,N_9306,N_9429);
xor U9553 (N_9553,N_9317,N_9460);
nor U9554 (N_9554,N_9310,N_9259);
xor U9555 (N_9555,N_9353,N_9253);
and U9556 (N_9556,N_9434,N_9364);
nor U9557 (N_9557,N_9423,N_9371);
nor U9558 (N_9558,N_9311,N_9432);
xnor U9559 (N_9559,N_9439,N_9346);
or U9560 (N_9560,N_9324,N_9402);
xnor U9561 (N_9561,N_9312,N_9492);
or U9562 (N_9562,N_9369,N_9394);
xnor U9563 (N_9563,N_9403,N_9359);
nand U9564 (N_9564,N_9375,N_9345);
xnor U9565 (N_9565,N_9443,N_9451);
and U9566 (N_9566,N_9285,N_9321);
nand U9567 (N_9567,N_9397,N_9273);
xnor U9568 (N_9568,N_9270,N_9480);
nand U9569 (N_9569,N_9305,N_9461);
xor U9570 (N_9570,N_9373,N_9304);
nor U9571 (N_9571,N_9298,N_9379);
nor U9572 (N_9572,N_9466,N_9267);
nand U9573 (N_9573,N_9370,N_9333);
nand U9574 (N_9574,N_9337,N_9436);
and U9575 (N_9575,N_9372,N_9316);
xnor U9576 (N_9576,N_9433,N_9489);
or U9577 (N_9577,N_9258,N_9488);
xor U9578 (N_9578,N_9265,N_9389);
or U9579 (N_9579,N_9471,N_9347);
or U9580 (N_9580,N_9315,N_9368);
nor U9581 (N_9581,N_9289,N_9459);
nand U9582 (N_9582,N_9446,N_9457);
nor U9583 (N_9583,N_9262,N_9437);
or U9584 (N_9584,N_9447,N_9326);
and U9585 (N_9585,N_9269,N_9286);
nor U9586 (N_9586,N_9425,N_9426);
nor U9587 (N_9587,N_9445,N_9421);
or U9588 (N_9588,N_9462,N_9328);
nor U9589 (N_9589,N_9280,N_9407);
and U9590 (N_9590,N_9419,N_9483);
nor U9591 (N_9591,N_9493,N_9329);
and U9592 (N_9592,N_9479,N_9331);
xor U9593 (N_9593,N_9497,N_9455);
xor U9594 (N_9594,N_9487,N_9476);
or U9595 (N_9595,N_9287,N_9340);
nor U9596 (N_9596,N_9392,N_9472);
nand U9597 (N_9597,N_9322,N_9336);
and U9598 (N_9598,N_9499,N_9395);
or U9599 (N_9599,N_9420,N_9387);
or U9600 (N_9600,N_9383,N_9452);
and U9601 (N_9601,N_9424,N_9380);
and U9602 (N_9602,N_9374,N_9293);
and U9603 (N_9603,N_9299,N_9494);
xor U9604 (N_9604,N_9357,N_9362);
and U9605 (N_9605,N_9365,N_9381);
nand U9606 (N_9606,N_9396,N_9456);
nand U9607 (N_9607,N_9413,N_9314);
nand U9608 (N_9608,N_9367,N_9469);
or U9609 (N_9609,N_9411,N_9252);
or U9610 (N_9610,N_9308,N_9399);
nand U9611 (N_9611,N_9484,N_9391);
and U9612 (N_9612,N_9386,N_9491);
xor U9613 (N_9613,N_9382,N_9260);
or U9614 (N_9614,N_9343,N_9409);
xor U9615 (N_9615,N_9444,N_9438);
nor U9616 (N_9616,N_9470,N_9257);
or U9617 (N_9617,N_9358,N_9377);
nor U9618 (N_9618,N_9410,N_9290);
xor U9619 (N_9619,N_9427,N_9288);
xnor U9620 (N_9620,N_9302,N_9303);
xor U9621 (N_9621,N_9349,N_9282);
or U9622 (N_9622,N_9385,N_9313);
nor U9623 (N_9623,N_9256,N_9473);
xor U9624 (N_9624,N_9414,N_9344);
nor U9625 (N_9625,N_9448,N_9280);
and U9626 (N_9626,N_9317,N_9396);
nand U9627 (N_9627,N_9269,N_9260);
xnor U9628 (N_9628,N_9396,N_9307);
nor U9629 (N_9629,N_9397,N_9327);
or U9630 (N_9630,N_9251,N_9363);
nand U9631 (N_9631,N_9467,N_9491);
xor U9632 (N_9632,N_9283,N_9302);
and U9633 (N_9633,N_9302,N_9440);
nand U9634 (N_9634,N_9460,N_9368);
and U9635 (N_9635,N_9394,N_9430);
xor U9636 (N_9636,N_9285,N_9267);
nor U9637 (N_9637,N_9405,N_9252);
or U9638 (N_9638,N_9423,N_9287);
or U9639 (N_9639,N_9463,N_9269);
and U9640 (N_9640,N_9357,N_9255);
nor U9641 (N_9641,N_9405,N_9468);
nand U9642 (N_9642,N_9285,N_9308);
or U9643 (N_9643,N_9433,N_9280);
nand U9644 (N_9644,N_9280,N_9493);
or U9645 (N_9645,N_9492,N_9254);
nor U9646 (N_9646,N_9489,N_9373);
nor U9647 (N_9647,N_9471,N_9456);
nand U9648 (N_9648,N_9472,N_9399);
nand U9649 (N_9649,N_9343,N_9277);
xor U9650 (N_9650,N_9457,N_9439);
or U9651 (N_9651,N_9308,N_9485);
nand U9652 (N_9652,N_9309,N_9263);
nand U9653 (N_9653,N_9487,N_9489);
nor U9654 (N_9654,N_9425,N_9348);
and U9655 (N_9655,N_9391,N_9392);
or U9656 (N_9656,N_9347,N_9254);
nor U9657 (N_9657,N_9390,N_9260);
nor U9658 (N_9658,N_9382,N_9492);
nor U9659 (N_9659,N_9409,N_9405);
and U9660 (N_9660,N_9378,N_9320);
nand U9661 (N_9661,N_9397,N_9378);
nand U9662 (N_9662,N_9327,N_9418);
nand U9663 (N_9663,N_9351,N_9413);
nand U9664 (N_9664,N_9466,N_9432);
nor U9665 (N_9665,N_9313,N_9453);
or U9666 (N_9666,N_9451,N_9477);
nand U9667 (N_9667,N_9322,N_9357);
or U9668 (N_9668,N_9404,N_9401);
xnor U9669 (N_9669,N_9266,N_9284);
or U9670 (N_9670,N_9251,N_9306);
nand U9671 (N_9671,N_9312,N_9310);
and U9672 (N_9672,N_9305,N_9390);
nor U9673 (N_9673,N_9366,N_9289);
xor U9674 (N_9674,N_9410,N_9309);
nor U9675 (N_9675,N_9394,N_9447);
xor U9676 (N_9676,N_9496,N_9439);
nand U9677 (N_9677,N_9268,N_9466);
or U9678 (N_9678,N_9282,N_9309);
nand U9679 (N_9679,N_9339,N_9408);
and U9680 (N_9680,N_9342,N_9490);
nor U9681 (N_9681,N_9368,N_9462);
nor U9682 (N_9682,N_9364,N_9394);
and U9683 (N_9683,N_9416,N_9358);
and U9684 (N_9684,N_9451,N_9345);
or U9685 (N_9685,N_9490,N_9478);
nand U9686 (N_9686,N_9395,N_9347);
and U9687 (N_9687,N_9440,N_9405);
or U9688 (N_9688,N_9315,N_9359);
or U9689 (N_9689,N_9415,N_9371);
and U9690 (N_9690,N_9265,N_9321);
or U9691 (N_9691,N_9286,N_9312);
nand U9692 (N_9692,N_9274,N_9492);
and U9693 (N_9693,N_9344,N_9374);
nor U9694 (N_9694,N_9371,N_9298);
nor U9695 (N_9695,N_9259,N_9432);
nand U9696 (N_9696,N_9368,N_9331);
or U9697 (N_9697,N_9335,N_9478);
and U9698 (N_9698,N_9475,N_9317);
nor U9699 (N_9699,N_9475,N_9349);
and U9700 (N_9700,N_9481,N_9382);
nand U9701 (N_9701,N_9498,N_9492);
and U9702 (N_9702,N_9376,N_9394);
or U9703 (N_9703,N_9358,N_9420);
nand U9704 (N_9704,N_9436,N_9416);
xnor U9705 (N_9705,N_9456,N_9295);
and U9706 (N_9706,N_9306,N_9269);
nor U9707 (N_9707,N_9483,N_9470);
and U9708 (N_9708,N_9497,N_9405);
nor U9709 (N_9709,N_9487,N_9362);
xnor U9710 (N_9710,N_9290,N_9334);
or U9711 (N_9711,N_9467,N_9359);
nand U9712 (N_9712,N_9262,N_9306);
or U9713 (N_9713,N_9488,N_9490);
nand U9714 (N_9714,N_9417,N_9478);
nor U9715 (N_9715,N_9401,N_9327);
and U9716 (N_9716,N_9449,N_9481);
xor U9717 (N_9717,N_9365,N_9369);
nand U9718 (N_9718,N_9454,N_9255);
nand U9719 (N_9719,N_9457,N_9256);
xor U9720 (N_9720,N_9362,N_9371);
nor U9721 (N_9721,N_9343,N_9454);
nand U9722 (N_9722,N_9414,N_9332);
xnor U9723 (N_9723,N_9385,N_9338);
nor U9724 (N_9724,N_9347,N_9352);
nor U9725 (N_9725,N_9416,N_9468);
xnor U9726 (N_9726,N_9263,N_9431);
nor U9727 (N_9727,N_9304,N_9486);
and U9728 (N_9728,N_9368,N_9392);
nor U9729 (N_9729,N_9275,N_9370);
xnor U9730 (N_9730,N_9464,N_9281);
nand U9731 (N_9731,N_9421,N_9364);
and U9732 (N_9732,N_9332,N_9401);
or U9733 (N_9733,N_9378,N_9419);
nor U9734 (N_9734,N_9479,N_9350);
nor U9735 (N_9735,N_9497,N_9454);
xor U9736 (N_9736,N_9265,N_9258);
nand U9737 (N_9737,N_9422,N_9486);
and U9738 (N_9738,N_9464,N_9390);
nor U9739 (N_9739,N_9284,N_9283);
and U9740 (N_9740,N_9339,N_9318);
nand U9741 (N_9741,N_9286,N_9338);
nor U9742 (N_9742,N_9473,N_9270);
nor U9743 (N_9743,N_9296,N_9467);
nor U9744 (N_9744,N_9318,N_9269);
and U9745 (N_9745,N_9353,N_9445);
xnor U9746 (N_9746,N_9312,N_9499);
nor U9747 (N_9747,N_9339,N_9434);
nand U9748 (N_9748,N_9313,N_9352);
and U9749 (N_9749,N_9497,N_9396);
xor U9750 (N_9750,N_9605,N_9522);
nand U9751 (N_9751,N_9709,N_9525);
nor U9752 (N_9752,N_9598,N_9712);
xnor U9753 (N_9753,N_9713,N_9737);
and U9754 (N_9754,N_9549,N_9682);
xnor U9755 (N_9755,N_9546,N_9530);
xnor U9756 (N_9756,N_9721,N_9670);
xnor U9757 (N_9757,N_9618,N_9631);
or U9758 (N_9758,N_9654,N_9628);
or U9759 (N_9759,N_9526,N_9511);
nand U9760 (N_9760,N_9616,N_9700);
and U9761 (N_9761,N_9567,N_9537);
and U9762 (N_9762,N_9678,N_9610);
and U9763 (N_9763,N_9746,N_9542);
nor U9764 (N_9764,N_9749,N_9699);
nor U9765 (N_9765,N_9738,N_9646);
and U9766 (N_9766,N_9614,N_9603);
or U9767 (N_9767,N_9505,N_9544);
and U9768 (N_9768,N_9674,N_9729);
xnor U9769 (N_9769,N_9748,N_9509);
or U9770 (N_9770,N_9568,N_9510);
nor U9771 (N_9771,N_9705,N_9565);
nand U9772 (N_9772,N_9643,N_9516);
xor U9773 (N_9773,N_9664,N_9677);
and U9774 (N_9774,N_9629,N_9571);
xnor U9775 (N_9775,N_9651,N_9706);
nand U9776 (N_9776,N_9653,N_9722);
nor U9777 (N_9777,N_9715,N_9588);
or U9778 (N_9778,N_9523,N_9625);
nand U9779 (N_9779,N_9644,N_9547);
and U9780 (N_9780,N_9666,N_9504);
or U9781 (N_9781,N_9650,N_9680);
nand U9782 (N_9782,N_9711,N_9639);
or U9783 (N_9783,N_9668,N_9580);
and U9784 (N_9784,N_9617,N_9661);
and U9785 (N_9785,N_9636,N_9707);
or U9786 (N_9786,N_9663,N_9601);
nor U9787 (N_9787,N_9689,N_9669);
nor U9788 (N_9788,N_9742,N_9622);
or U9789 (N_9789,N_9620,N_9691);
nor U9790 (N_9790,N_9648,N_9553);
and U9791 (N_9791,N_9692,N_9735);
xor U9792 (N_9792,N_9672,N_9671);
xnor U9793 (N_9793,N_9695,N_9703);
xnor U9794 (N_9794,N_9569,N_9665);
nor U9795 (N_9795,N_9717,N_9624);
and U9796 (N_9796,N_9658,N_9513);
xor U9797 (N_9797,N_9655,N_9556);
and U9798 (N_9798,N_9607,N_9589);
and U9799 (N_9799,N_9550,N_9633);
or U9800 (N_9800,N_9652,N_9538);
or U9801 (N_9801,N_9533,N_9576);
nand U9802 (N_9802,N_9638,N_9731);
nand U9803 (N_9803,N_9545,N_9627);
or U9804 (N_9804,N_9583,N_9529);
or U9805 (N_9805,N_9602,N_9611);
and U9806 (N_9806,N_9649,N_9608);
nor U9807 (N_9807,N_9570,N_9720);
nand U9808 (N_9808,N_9600,N_9623);
xnor U9809 (N_9809,N_9515,N_9687);
xor U9810 (N_9810,N_9562,N_9710);
or U9811 (N_9811,N_9554,N_9535);
nand U9812 (N_9812,N_9585,N_9503);
xor U9813 (N_9813,N_9718,N_9564);
nor U9814 (N_9814,N_9514,N_9642);
nor U9815 (N_9815,N_9698,N_9667);
nand U9816 (N_9816,N_9701,N_9739);
nor U9817 (N_9817,N_9688,N_9641);
or U9818 (N_9818,N_9679,N_9743);
and U9819 (N_9819,N_9512,N_9536);
and U9820 (N_9820,N_9581,N_9590);
nor U9821 (N_9821,N_9508,N_9745);
nand U9822 (N_9822,N_9675,N_9543);
xnor U9823 (N_9823,N_9632,N_9541);
and U9824 (N_9824,N_9615,N_9500);
nor U9825 (N_9825,N_9577,N_9621);
nor U9826 (N_9826,N_9724,N_9694);
or U9827 (N_9827,N_9747,N_9728);
nor U9828 (N_9828,N_9683,N_9723);
xnor U9829 (N_9829,N_9502,N_9626);
nor U9830 (N_9830,N_9593,N_9563);
xor U9831 (N_9831,N_9708,N_9609);
nor U9832 (N_9832,N_9551,N_9596);
nor U9833 (N_9833,N_9534,N_9696);
or U9834 (N_9834,N_9582,N_9591);
xor U9835 (N_9835,N_9555,N_9730);
and U9836 (N_9836,N_9528,N_9519);
xor U9837 (N_9837,N_9613,N_9634);
or U9838 (N_9838,N_9662,N_9734);
nand U9839 (N_9839,N_9531,N_9726);
and U9840 (N_9840,N_9579,N_9527);
nor U9841 (N_9841,N_9704,N_9685);
xnor U9842 (N_9842,N_9572,N_9524);
nor U9843 (N_9843,N_9659,N_9584);
xnor U9844 (N_9844,N_9635,N_9732);
xnor U9845 (N_9845,N_9714,N_9673);
nand U9846 (N_9846,N_9540,N_9690);
and U9847 (N_9847,N_9716,N_9606);
nand U9848 (N_9848,N_9693,N_9578);
xor U9849 (N_9849,N_9561,N_9560);
nand U9850 (N_9850,N_9592,N_9660);
or U9851 (N_9851,N_9647,N_9597);
xor U9852 (N_9852,N_9744,N_9566);
and U9853 (N_9853,N_9645,N_9740);
xor U9854 (N_9854,N_9575,N_9686);
and U9855 (N_9855,N_9559,N_9521);
nor U9856 (N_9856,N_9736,N_9640);
nand U9857 (N_9857,N_9595,N_9619);
nor U9858 (N_9858,N_9637,N_9676);
or U9859 (N_9859,N_9587,N_9725);
nor U9860 (N_9860,N_9719,N_9697);
and U9861 (N_9861,N_9532,N_9702);
xnor U9862 (N_9862,N_9558,N_9501);
and U9863 (N_9863,N_9539,N_9557);
nor U9864 (N_9864,N_9604,N_9741);
and U9865 (N_9865,N_9594,N_9520);
nand U9866 (N_9866,N_9630,N_9684);
nor U9867 (N_9867,N_9586,N_9657);
nor U9868 (N_9868,N_9548,N_9656);
or U9869 (N_9869,N_9681,N_9506);
and U9870 (N_9870,N_9552,N_9727);
nor U9871 (N_9871,N_9517,N_9612);
xnor U9872 (N_9872,N_9507,N_9599);
nor U9873 (N_9873,N_9733,N_9518);
and U9874 (N_9874,N_9573,N_9574);
nand U9875 (N_9875,N_9504,N_9733);
nand U9876 (N_9876,N_9672,N_9692);
nand U9877 (N_9877,N_9687,N_9711);
xnor U9878 (N_9878,N_9734,N_9686);
xor U9879 (N_9879,N_9620,N_9593);
and U9880 (N_9880,N_9641,N_9573);
nand U9881 (N_9881,N_9535,N_9627);
nand U9882 (N_9882,N_9741,N_9515);
nor U9883 (N_9883,N_9697,N_9614);
or U9884 (N_9884,N_9549,N_9528);
nand U9885 (N_9885,N_9693,N_9543);
or U9886 (N_9886,N_9590,N_9673);
or U9887 (N_9887,N_9583,N_9540);
and U9888 (N_9888,N_9507,N_9508);
nor U9889 (N_9889,N_9741,N_9665);
nand U9890 (N_9890,N_9618,N_9719);
xnor U9891 (N_9891,N_9706,N_9566);
nand U9892 (N_9892,N_9621,N_9607);
nand U9893 (N_9893,N_9570,N_9707);
xor U9894 (N_9894,N_9746,N_9713);
xor U9895 (N_9895,N_9601,N_9709);
nand U9896 (N_9896,N_9517,N_9681);
nor U9897 (N_9897,N_9625,N_9670);
xor U9898 (N_9898,N_9739,N_9643);
nand U9899 (N_9899,N_9601,N_9616);
nor U9900 (N_9900,N_9524,N_9660);
nand U9901 (N_9901,N_9557,N_9694);
nand U9902 (N_9902,N_9607,N_9574);
nand U9903 (N_9903,N_9686,N_9634);
xor U9904 (N_9904,N_9669,N_9683);
nor U9905 (N_9905,N_9536,N_9733);
xnor U9906 (N_9906,N_9695,N_9592);
or U9907 (N_9907,N_9665,N_9614);
and U9908 (N_9908,N_9581,N_9611);
nand U9909 (N_9909,N_9525,N_9573);
nor U9910 (N_9910,N_9559,N_9527);
xnor U9911 (N_9911,N_9504,N_9689);
or U9912 (N_9912,N_9536,N_9577);
nand U9913 (N_9913,N_9639,N_9745);
nand U9914 (N_9914,N_9548,N_9557);
nor U9915 (N_9915,N_9540,N_9616);
and U9916 (N_9916,N_9545,N_9534);
and U9917 (N_9917,N_9511,N_9601);
nor U9918 (N_9918,N_9578,N_9629);
nand U9919 (N_9919,N_9545,N_9609);
nor U9920 (N_9920,N_9651,N_9627);
and U9921 (N_9921,N_9625,N_9598);
xnor U9922 (N_9922,N_9560,N_9616);
or U9923 (N_9923,N_9578,N_9683);
nand U9924 (N_9924,N_9653,N_9689);
or U9925 (N_9925,N_9520,N_9719);
and U9926 (N_9926,N_9537,N_9733);
nor U9927 (N_9927,N_9594,N_9744);
or U9928 (N_9928,N_9561,N_9646);
nor U9929 (N_9929,N_9642,N_9564);
or U9930 (N_9930,N_9657,N_9575);
xnor U9931 (N_9931,N_9510,N_9713);
xnor U9932 (N_9932,N_9670,N_9615);
xnor U9933 (N_9933,N_9581,N_9733);
xnor U9934 (N_9934,N_9640,N_9742);
nor U9935 (N_9935,N_9638,N_9519);
xnor U9936 (N_9936,N_9632,N_9674);
or U9937 (N_9937,N_9629,N_9528);
nor U9938 (N_9938,N_9540,N_9658);
or U9939 (N_9939,N_9686,N_9593);
nor U9940 (N_9940,N_9570,N_9656);
xnor U9941 (N_9941,N_9678,N_9657);
nand U9942 (N_9942,N_9720,N_9557);
or U9943 (N_9943,N_9644,N_9557);
and U9944 (N_9944,N_9664,N_9719);
and U9945 (N_9945,N_9518,N_9621);
nor U9946 (N_9946,N_9629,N_9597);
and U9947 (N_9947,N_9714,N_9663);
and U9948 (N_9948,N_9590,N_9602);
or U9949 (N_9949,N_9514,N_9630);
or U9950 (N_9950,N_9620,N_9508);
nand U9951 (N_9951,N_9640,N_9601);
and U9952 (N_9952,N_9707,N_9687);
or U9953 (N_9953,N_9682,N_9562);
xnor U9954 (N_9954,N_9527,N_9624);
or U9955 (N_9955,N_9551,N_9593);
or U9956 (N_9956,N_9578,N_9700);
nor U9957 (N_9957,N_9685,N_9541);
and U9958 (N_9958,N_9588,N_9646);
or U9959 (N_9959,N_9676,N_9650);
nor U9960 (N_9960,N_9534,N_9581);
or U9961 (N_9961,N_9654,N_9514);
or U9962 (N_9962,N_9617,N_9685);
and U9963 (N_9963,N_9557,N_9670);
xor U9964 (N_9964,N_9574,N_9627);
nor U9965 (N_9965,N_9749,N_9606);
and U9966 (N_9966,N_9614,N_9655);
and U9967 (N_9967,N_9681,N_9690);
nor U9968 (N_9968,N_9601,N_9512);
or U9969 (N_9969,N_9596,N_9715);
xnor U9970 (N_9970,N_9596,N_9744);
nand U9971 (N_9971,N_9711,N_9675);
nor U9972 (N_9972,N_9741,N_9678);
nor U9973 (N_9973,N_9551,N_9685);
and U9974 (N_9974,N_9694,N_9693);
or U9975 (N_9975,N_9703,N_9712);
nand U9976 (N_9976,N_9569,N_9696);
or U9977 (N_9977,N_9603,N_9648);
xor U9978 (N_9978,N_9577,N_9721);
or U9979 (N_9979,N_9618,N_9654);
and U9980 (N_9980,N_9502,N_9598);
or U9981 (N_9981,N_9633,N_9625);
and U9982 (N_9982,N_9623,N_9655);
or U9983 (N_9983,N_9592,N_9544);
xnor U9984 (N_9984,N_9651,N_9726);
or U9985 (N_9985,N_9630,N_9534);
or U9986 (N_9986,N_9525,N_9629);
and U9987 (N_9987,N_9699,N_9715);
or U9988 (N_9988,N_9679,N_9584);
or U9989 (N_9989,N_9587,N_9576);
nand U9990 (N_9990,N_9624,N_9736);
and U9991 (N_9991,N_9664,N_9646);
xor U9992 (N_9992,N_9717,N_9524);
xnor U9993 (N_9993,N_9697,N_9705);
or U9994 (N_9994,N_9649,N_9714);
xor U9995 (N_9995,N_9560,N_9701);
xnor U9996 (N_9996,N_9606,N_9577);
xnor U9997 (N_9997,N_9749,N_9532);
or U9998 (N_9998,N_9686,N_9573);
nor U9999 (N_9999,N_9699,N_9642);
xnor U10000 (N_10000,N_9757,N_9882);
nor U10001 (N_10001,N_9895,N_9926);
nor U10002 (N_10002,N_9871,N_9950);
or U10003 (N_10003,N_9905,N_9838);
and U10004 (N_10004,N_9922,N_9992);
nand U10005 (N_10005,N_9886,N_9982);
nor U10006 (N_10006,N_9811,N_9888);
and U10007 (N_10007,N_9891,N_9807);
xor U10008 (N_10008,N_9818,N_9832);
or U10009 (N_10009,N_9932,N_9983);
xnor U10010 (N_10010,N_9842,N_9835);
and U10011 (N_10011,N_9930,N_9773);
or U10012 (N_10012,N_9981,N_9989);
or U10013 (N_10013,N_9795,N_9791);
xor U10014 (N_10014,N_9986,N_9846);
nor U10015 (N_10015,N_9924,N_9940);
nand U10016 (N_10016,N_9761,N_9917);
xnor U10017 (N_10017,N_9855,N_9767);
xnor U10018 (N_10018,N_9850,N_9921);
and U10019 (N_10019,N_9862,N_9839);
xnor U10020 (N_10020,N_9763,N_9885);
xnor U10021 (N_10021,N_9897,N_9931);
and U10022 (N_10022,N_9792,N_9994);
or U10023 (N_10023,N_9789,N_9975);
or U10024 (N_10024,N_9856,N_9787);
or U10025 (N_10025,N_9949,N_9809);
nand U10026 (N_10026,N_9851,N_9802);
and U10027 (N_10027,N_9942,N_9863);
nor U10028 (N_10028,N_9974,N_9883);
nor U10029 (N_10029,N_9904,N_9826);
nand U10030 (N_10030,N_9817,N_9947);
or U10031 (N_10031,N_9812,N_9998);
nor U10032 (N_10032,N_9770,N_9796);
xnor U10033 (N_10033,N_9887,N_9841);
xnor U10034 (N_10034,N_9870,N_9938);
nor U10035 (N_10035,N_9878,N_9972);
and U10036 (N_10036,N_9793,N_9805);
nor U10037 (N_10037,N_9900,N_9837);
nor U10038 (N_10038,N_9939,N_9753);
nand U10039 (N_10039,N_9772,N_9962);
nand U10040 (N_10040,N_9788,N_9991);
nand U10041 (N_10041,N_9967,N_9781);
xnor U10042 (N_10042,N_9903,N_9859);
nand U10043 (N_10043,N_9806,N_9799);
xor U10044 (N_10044,N_9907,N_9929);
xnor U10045 (N_10045,N_9840,N_9768);
nand U10046 (N_10046,N_9816,N_9906);
xnor U10047 (N_10047,N_9979,N_9785);
xor U10048 (N_10048,N_9877,N_9915);
or U10049 (N_10049,N_9892,N_9783);
nand U10050 (N_10050,N_9918,N_9861);
nor U10051 (N_10051,N_9923,N_9977);
nor U10052 (N_10052,N_9869,N_9825);
nand U10053 (N_10053,N_9821,N_9755);
xnor U10054 (N_10054,N_9800,N_9928);
nor U10055 (N_10055,N_9954,N_9779);
xnor U10056 (N_10056,N_9759,N_9758);
or U10057 (N_10057,N_9899,N_9893);
nand U10058 (N_10058,N_9955,N_9970);
or U10059 (N_10059,N_9958,N_9890);
or U10060 (N_10060,N_9762,N_9920);
nor U10061 (N_10061,N_9952,N_9808);
and U10062 (N_10062,N_9771,N_9898);
or U10063 (N_10063,N_9803,N_9910);
nor U10064 (N_10064,N_9911,N_9980);
xor U10065 (N_10065,N_9804,N_9822);
or U10066 (N_10066,N_9925,N_9819);
or U10067 (N_10067,N_9833,N_9765);
or U10068 (N_10068,N_9971,N_9913);
and U10069 (N_10069,N_9896,N_9784);
or U10070 (N_10070,N_9852,N_9941);
and U10071 (N_10071,N_9916,N_9756);
and U10072 (N_10072,N_9857,N_9985);
and U10073 (N_10073,N_9769,N_9797);
xnor U10074 (N_10074,N_9914,N_9960);
xor U10075 (N_10075,N_9936,N_9946);
nor U10076 (N_10076,N_9849,N_9937);
nor U10077 (N_10077,N_9865,N_9969);
or U10078 (N_10078,N_9814,N_9775);
xor U10079 (N_10079,N_9810,N_9860);
xor U10080 (N_10080,N_9894,N_9996);
or U10081 (N_10081,N_9935,N_9827);
or U10082 (N_10082,N_9909,N_9782);
nor U10083 (N_10083,N_9957,N_9964);
and U10084 (N_10084,N_9750,N_9948);
and U10085 (N_10085,N_9828,N_9927);
and U10086 (N_10086,N_9831,N_9798);
xor U10087 (N_10087,N_9966,N_9824);
nand U10088 (N_10088,N_9754,N_9976);
nor U10089 (N_10089,N_9943,N_9843);
nor U10090 (N_10090,N_9766,N_9780);
or U10091 (N_10091,N_9760,N_9813);
nand U10092 (N_10092,N_9845,N_9873);
nor U10093 (N_10093,N_9847,N_9984);
and U10094 (N_10094,N_9945,N_9751);
xor U10095 (N_10095,N_9978,N_9778);
nor U10096 (N_10096,N_9956,N_9786);
nor U10097 (N_10097,N_9874,N_9987);
xnor U10098 (N_10098,N_9790,N_9968);
nor U10099 (N_10099,N_9944,N_9752);
nor U10100 (N_10100,N_9844,N_9777);
or U10101 (N_10101,N_9988,N_9919);
xor U10102 (N_10102,N_9934,N_9953);
and U10103 (N_10103,N_9858,N_9901);
nand U10104 (N_10104,N_9866,N_9848);
xnor U10105 (N_10105,N_9872,N_9963);
xnor U10106 (N_10106,N_9961,N_9801);
nand U10107 (N_10107,N_9868,N_9997);
nand U10108 (N_10108,N_9834,N_9836);
nor U10109 (N_10109,N_9959,N_9951);
and U10110 (N_10110,N_9830,N_9879);
nand U10111 (N_10111,N_9908,N_9889);
or U10112 (N_10112,N_9820,N_9995);
nand U10113 (N_10113,N_9829,N_9999);
xor U10114 (N_10114,N_9881,N_9933);
nand U10115 (N_10115,N_9884,N_9815);
xor U10116 (N_10116,N_9864,N_9875);
nand U10117 (N_10117,N_9993,N_9823);
or U10118 (N_10118,N_9853,N_9854);
xor U10119 (N_10119,N_9902,N_9965);
and U10120 (N_10120,N_9776,N_9973);
nand U10121 (N_10121,N_9764,N_9990);
xor U10122 (N_10122,N_9912,N_9876);
nor U10123 (N_10123,N_9774,N_9880);
xnor U10124 (N_10124,N_9794,N_9867);
and U10125 (N_10125,N_9801,N_9771);
and U10126 (N_10126,N_9840,N_9892);
or U10127 (N_10127,N_9944,N_9921);
nor U10128 (N_10128,N_9982,N_9798);
and U10129 (N_10129,N_9803,N_9792);
or U10130 (N_10130,N_9845,N_9766);
or U10131 (N_10131,N_9770,N_9914);
or U10132 (N_10132,N_9802,N_9937);
nand U10133 (N_10133,N_9807,N_9976);
xnor U10134 (N_10134,N_9905,N_9982);
nand U10135 (N_10135,N_9979,N_9966);
xnor U10136 (N_10136,N_9828,N_9774);
and U10137 (N_10137,N_9895,N_9855);
or U10138 (N_10138,N_9898,N_9839);
nand U10139 (N_10139,N_9892,N_9946);
xor U10140 (N_10140,N_9839,N_9891);
xnor U10141 (N_10141,N_9849,N_9932);
nor U10142 (N_10142,N_9785,N_9827);
nand U10143 (N_10143,N_9851,N_9913);
or U10144 (N_10144,N_9790,N_9751);
nor U10145 (N_10145,N_9769,N_9793);
nand U10146 (N_10146,N_9984,N_9909);
nor U10147 (N_10147,N_9973,N_9851);
nand U10148 (N_10148,N_9968,N_9863);
nand U10149 (N_10149,N_9897,N_9798);
nor U10150 (N_10150,N_9764,N_9887);
or U10151 (N_10151,N_9840,N_9791);
xnor U10152 (N_10152,N_9759,N_9815);
nand U10153 (N_10153,N_9933,N_9778);
xnor U10154 (N_10154,N_9970,N_9861);
or U10155 (N_10155,N_9811,N_9951);
and U10156 (N_10156,N_9818,N_9795);
or U10157 (N_10157,N_9885,N_9890);
nor U10158 (N_10158,N_9919,N_9778);
xor U10159 (N_10159,N_9898,N_9881);
or U10160 (N_10160,N_9901,N_9958);
nand U10161 (N_10161,N_9799,N_9772);
xor U10162 (N_10162,N_9947,N_9872);
or U10163 (N_10163,N_9895,N_9811);
nor U10164 (N_10164,N_9892,N_9863);
nor U10165 (N_10165,N_9776,N_9886);
or U10166 (N_10166,N_9917,N_9999);
xnor U10167 (N_10167,N_9911,N_9886);
or U10168 (N_10168,N_9858,N_9806);
xnor U10169 (N_10169,N_9857,N_9900);
and U10170 (N_10170,N_9797,N_9878);
or U10171 (N_10171,N_9940,N_9783);
nor U10172 (N_10172,N_9892,N_9896);
and U10173 (N_10173,N_9879,N_9791);
and U10174 (N_10174,N_9865,N_9784);
nor U10175 (N_10175,N_9897,N_9887);
nand U10176 (N_10176,N_9819,N_9774);
nand U10177 (N_10177,N_9922,N_9870);
and U10178 (N_10178,N_9849,N_9803);
xnor U10179 (N_10179,N_9903,N_9782);
nor U10180 (N_10180,N_9886,N_9817);
nor U10181 (N_10181,N_9844,N_9947);
and U10182 (N_10182,N_9851,N_9935);
nor U10183 (N_10183,N_9855,N_9948);
or U10184 (N_10184,N_9903,N_9841);
xor U10185 (N_10185,N_9765,N_9762);
or U10186 (N_10186,N_9913,N_9973);
and U10187 (N_10187,N_9969,N_9975);
nor U10188 (N_10188,N_9854,N_9805);
and U10189 (N_10189,N_9934,N_9994);
nor U10190 (N_10190,N_9821,N_9890);
and U10191 (N_10191,N_9772,N_9774);
or U10192 (N_10192,N_9932,N_9853);
and U10193 (N_10193,N_9766,N_9943);
nand U10194 (N_10194,N_9935,N_9848);
nor U10195 (N_10195,N_9853,N_9980);
nand U10196 (N_10196,N_9921,N_9847);
nor U10197 (N_10197,N_9760,N_9809);
nor U10198 (N_10198,N_9911,N_9891);
nand U10199 (N_10199,N_9759,N_9814);
nand U10200 (N_10200,N_9913,N_9969);
nor U10201 (N_10201,N_9921,N_9753);
xnor U10202 (N_10202,N_9976,N_9773);
nand U10203 (N_10203,N_9991,N_9918);
and U10204 (N_10204,N_9755,N_9822);
and U10205 (N_10205,N_9893,N_9980);
xnor U10206 (N_10206,N_9985,N_9786);
xnor U10207 (N_10207,N_9871,N_9878);
nand U10208 (N_10208,N_9850,N_9773);
nor U10209 (N_10209,N_9838,N_9795);
xnor U10210 (N_10210,N_9958,N_9915);
nand U10211 (N_10211,N_9752,N_9870);
nand U10212 (N_10212,N_9757,N_9992);
xnor U10213 (N_10213,N_9986,N_9929);
nor U10214 (N_10214,N_9854,N_9877);
and U10215 (N_10215,N_9938,N_9946);
nand U10216 (N_10216,N_9866,N_9847);
xnor U10217 (N_10217,N_9855,N_9935);
and U10218 (N_10218,N_9817,N_9801);
and U10219 (N_10219,N_9986,N_9828);
nand U10220 (N_10220,N_9844,N_9849);
and U10221 (N_10221,N_9964,N_9840);
nor U10222 (N_10222,N_9761,N_9999);
nor U10223 (N_10223,N_9986,N_9971);
and U10224 (N_10224,N_9855,N_9853);
xnor U10225 (N_10225,N_9969,N_9873);
and U10226 (N_10226,N_9844,N_9934);
nor U10227 (N_10227,N_9925,N_9936);
and U10228 (N_10228,N_9852,N_9964);
nand U10229 (N_10229,N_9835,N_9833);
nand U10230 (N_10230,N_9969,N_9759);
nor U10231 (N_10231,N_9813,N_9990);
xor U10232 (N_10232,N_9783,N_9791);
or U10233 (N_10233,N_9875,N_9905);
xnor U10234 (N_10234,N_9970,N_9866);
nor U10235 (N_10235,N_9860,N_9986);
or U10236 (N_10236,N_9750,N_9760);
nor U10237 (N_10237,N_9860,N_9916);
nor U10238 (N_10238,N_9814,N_9852);
and U10239 (N_10239,N_9799,N_9928);
nor U10240 (N_10240,N_9972,N_9768);
nand U10241 (N_10241,N_9824,N_9921);
and U10242 (N_10242,N_9755,N_9847);
or U10243 (N_10243,N_9781,N_9793);
nand U10244 (N_10244,N_9993,N_9980);
nand U10245 (N_10245,N_9984,N_9871);
nor U10246 (N_10246,N_9958,N_9790);
nand U10247 (N_10247,N_9870,N_9901);
nand U10248 (N_10248,N_9999,N_9936);
xor U10249 (N_10249,N_9917,N_9853);
nand U10250 (N_10250,N_10099,N_10085);
nor U10251 (N_10251,N_10176,N_10249);
nor U10252 (N_10252,N_10219,N_10220);
and U10253 (N_10253,N_10229,N_10157);
and U10254 (N_10254,N_10245,N_10094);
and U10255 (N_10255,N_10064,N_10096);
xnor U10256 (N_10256,N_10208,N_10165);
nand U10257 (N_10257,N_10013,N_10228);
and U10258 (N_10258,N_10083,N_10057);
or U10259 (N_10259,N_10188,N_10135);
and U10260 (N_10260,N_10158,N_10224);
xnor U10261 (N_10261,N_10177,N_10233);
nor U10262 (N_10262,N_10078,N_10113);
and U10263 (N_10263,N_10049,N_10215);
xnor U10264 (N_10264,N_10124,N_10092);
or U10265 (N_10265,N_10054,N_10050);
or U10266 (N_10266,N_10112,N_10030);
and U10267 (N_10267,N_10015,N_10175);
xor U10268 (N_10268,N_10174,N_10155);
nor U10269 (N_10269,N_10067,N_10202);
and U10270 (N_10270,N_10042,N_10173);
and U10271 (N_10271,N_10110,N_10193);
or U10272 (N_10272,N_10171,N_10051);
nand U10273 (N_10273,N_10243,N_10031);
and U10274 (N_10274,N_10120,N_10076);
nor U10275 (N_10275,N_10068,N_10218);
xor U10276 (N_10276,N_10119,N_10232);
xnor U10277 (N_10277,N_10070,N_10037);
nand U10278 (N_10278,N_10035,N_10194);
nor U10279 (N_10279,N_10074,N_10235);
xnor U10280 (N_10280,N_10114,N_10234);
and U10281 (N_10281,N_10205,N_10145);
nand U10282 (N_10282,N_10223,N_10097);
nand U10283 (N_10283,N_10126,N_10059);
xnor U10284 (N_10284,N_10024,N_10192);
nor U10285 (N_10285,N_10216,N_10069);
or U10286 (N_10286,N_10199,N_10156);
and U10287 (N_10287,N_10217,N_10018);
nor U10288 (N_10288,N_10221,N_10009);
nand U10289 (N_10289,N_10066,N_10038);
nor U10290 (N_10290,N_10246,N_10209);
nand U10291 (N_10291,N_10008,N_10147);
nand U10292 (N_10292,N_10123,N_10003);
and U10293 (N_10293,N_10153,N_10213);
and U10294 (N_10294,N_10162,N_10247);
or U10295 (N_10295,N_10212,N_10043);
nor U10296 (N_10296,N_10071,N_10084);
and U10297 (N_10297,N_10026,N_10190);
or U10298 (N_10298,N_10065,N_10241);
nor U10299 (N_10299,N_10117,N_10130);
xor U10300 (N_10300,N_10014,N_10102);
nor U10301 (N_10301,N_10197,N_10012);
nand U10302 (N_10302,N_10116,N_10081);
and U10303 (N_10303,N_10151,N_10007);
or U10304 (N_10304,N_10144,N_10248);
and U10305 (N_10305,N_10138,N_10131);
nor U10306 (N_10306,N_10106,N_10109);
and U10307 (N_10307,N_10187,N_10060);
xor U10308 (N_10308,N_10047,N_10041);
or U10309 (N_10309,N_10207,N_10089);
nand U10310 (N_10310,N_10146,N_10046);
or U10311 (N_10311,N_10204,N_10226);
xor U10312 (N_10312,N_10062,N_10164);
nand U10313 (N_10313,N_10108,N_10056);
or U10314 (N_10314,N_10104,N_10191);
and U10315 (N_10315,N_10020,N_10163);
and U10316 (N_10316,N_10048,N_10105);
and U10317 (N_10317,N_10230,N_10134);
xor U10318 (N_10318,N_10027,N_10128);
and U10319 (N_10319,N_10023,N_10159);
or U10320 (N_10320,N_10045,N_10107);
xor U10321 (N_10321,N_10198,N_10161);
and U10322 (N_10322,N_10040,N_10001);
or U10323 (N_10323,N_10087,N_10022);
xor U10324 (N_10324,N_10139,N_10214);
or U10325 (N_10325,N_10111,N_10180);
and U10326 (N_10326,N_10010,N_10236);
nand U10327 (N_10327,N_10005,N_10167);
nor U10328 (N_10328,N_10179,N_10033);
xnor U10329 (N_10329,N_10152,N_10160);
and U10330 (N_10330,N_10017,N_10121);
xor U10331 (N_10331,N_10178,N_10227);
nand U10332 (N_10332,N_10052,N_10090);
nor U10333 (N_10333,N_10073,N_10142);
nand U10334 (N_10334,N_10240,N_10129);
or U10335 (N_10335,N_10200,N_10053);
nand U10336 (N_10336,N_10029,N_10168);
xor U10337 (N_10337,N_10028,N_10086);
nand U10338 (N_10338,N_10034,N_10036);
xnor U10339 (N_10339,N_10184,N_10203);
nor U10340 (N_10340,N_10075,N_10183);
xnor U10341 (N_10341,N_10237,N_10118);
or U10342 (N_10342,N_10201,N_10011);
and U10343 (N_10343,N_10141,N_10206);
and U10344 (N_10344,N_10149,N_10063);
or U10345 (N_10345,N_10181,N_10132);
nand U10346 (N_10346,N_10189,N_10133);
xnor U10347 (N_10347,N_10079,N_10143);
and U10348 (N_10348,N_10025,N_10055);
and U10349 (N_10349,N_10244,N_10150);
xnor U10350 (N_10350,N_10231,N_10021);
nor U10351 (N_10351,N_10032,N_10137);
xnor U10352 (N_10352,N_10115,N_10122);
nor U10353 (N_10353,N_10101,N_10077);
and U10354 (N_10354,N_10098,N_10100);
nand U10355 (N_10355,N_10211,N_10169);
and U10356 (N_10356,N_10093,N_10006);
nor U10357 (N_10357,N_10166,N_10127);
nand U10358 (N_10358,N_10154,N_10039);
and U10359 (N_10359,N_10210,N_10019);
and U10360 (N_10360,N_10002,N_10000);
xor U10361 (N_10361,N_10185,N_10016);
and U10362 (N_10362,N_10095,N_10196);
and U10363 (N_10363,N_10088,N_10172);
nand U10364 (N_10364,N_10004,N_10186);
or U10365 (N_10365,N_10238,N_10091);
or U10366 (N_10366,N_10195,N_10242);
and U10367 (N_10367,N_10082,N_10239);
nor U10368 (N_10368,N_10136,N_10148);
xnor U10369 (N_10369,N_10140,N_10072);
nor U10370 (N_10370,N_10044,N_10103);
and U10371 (N_10371,N_10170,N_10061);
and U10372 (N_10372,N_10225,N_10058);
nand U10373 (N_10373,N_10182,N_10125);
nand U10374 (N_10374,N_10080,N_10222);
nand U10375 (N_10375,N_10018,N_10004);
xor U10376 (N_10376,N_10119,N_10214);
and U10377 (N_10377,N_10200,N_10072);
nor U10378 (N_10378,N_10145,N_10184);
nand U10379 (N_10379,N_10154,N_10203);
nand U10380 (N_10380,N_10231,N_10172);
or U10381 (N_10381,N_10032,N_10144);
nor U10382 (N_10382,N_10064,N_10237);
and U10383 (N_10383,N_10237,N_10164);
nand U10384 (N_10384,N_10222,N_10237);
or U10385 (N_10385,N_10048,N_10204);
or U10386 (N_10386,N_10115,N_10195);
nor U10387 (N_10387,N_10155,N_10188);
nor U10388 (N_10388,N_10186,N_10053);
or U10389 (N_10389,N_10120,N_10177);
xor U10390 (N_10390,N_10114,N_10232);
nor U10391 (N_10391,N_10205,N_10235);
nand U10392 (N_10392,N_10083,N_10113);
or U10393 (N_10393,N_10153,N_10181);
nor U10394 (N_10394,N_10226,N_10066);
nor U10395 (N_10395,N_10101,N_10058);
nor U10396 (N_10396,N_10000,N_10011);
or U10397 (N_10397,N_10122,N_10108);
and U10398 (N_10398,N_10109,N_10203);
xor U10399 (N_10399,N_10060,N_10051);
and U10400 (N_10400,N_10224,N_10065);
nor U10401 (N_10401,N_10097,N_10220);
and U10402 (N_10402,N_10200,N_10004);
nor U10403 (N_10403,N_10001,N_10020);
xnor U10404 (N_10404,N_10242,N_10152);
nor U10405 (N_10405,N_10015,N_10192);
nor U10406 (N_10406,N_10165,N_10171);
xor U10407 (N_10407,N_10145,N_10050);
and U10408 (N_10408,N_10015,N_10133);
xnor U10409 (N_10409,N_10179,N_10232);
xor U10410 (N_10410,N_10153,N_10096);
and U10411 (N_10411,N_10137,N_10001);
and U10412 (N_10412,N_10074,N_10009);
or U10413 (N_10413,N_10099,N_10203);
and U10414 (N_10414,N_10044,N_10188);
and U10415 (N_10415,N_10208,N_10152);
xor U10416 (N_10416,N_10235,N_10165);
xnor U10417 (N_10417,N_10047,N_10074);
nand U10418 (N_10418,N_10141,N_10021);
nand U10419 (N_10419,N_10027,N_10085);
or U10420 (N_10420,N_10049,N_10045);
and U10421 (N_10421,N_10072,N_10086);
nand U10422 (N_10422,N_10199,N_10069);
or U10423 (N_10423,N_10019,N_10151);
nand U10424 (N_10424,N_10042,N_10057);
nand U10425 (N_10425,N_10008,N_10164);
and U10426 (N_10426,N_10063,N_10076);
xnor U10427 (N_10427,N_10051,N_10180);
and U10428 (N_10428,N_10001,N_10076);
xnor U10429 (N_10429,N_10003,N_10008);
xor U10430 (N_10430,N_10145,N_10123);
nand U10431 (N_10431,N_10179,N_10143);
xor U10432 (N_10432,N_10092,N_10242);
xor U10433 (N_10433,N_10075,N_10069);
nand U10434 (N_10434,N_10026,N_10128);
xnor U10435 (N_10435,N_10016,N_10234);
xor U10436 (N_10436,N_10170,N_10066);
xor U10437 (N_10437,N_10020,N_10066);
nor U10438 (N_10438,N_10067,N_10134);
nand U10439 (N_10439,N_10138,N_10108);
or U10440 (N_10440,N_10134,N_10128);
or U10441 (N_10441,N_10076,N_10248);
nor U10442 (N_10442,N_10239,N_10038);
nor U10443 (N_10443,N_10223,N_10129);
xnor U10444 (N_10444,N_10145,N_10096);
xor U10445 (N_10445,N_10192,N_10219);
or U10446 (N_10446,N_10037,N_10071);
and U10447 (N_10447,N_10154,N_10128);
or U10448 (N_10448,N_10127,N_10206);
nand U10449 (N_10449,N_10130,N_10062);
and U10450 (N_10450,N_10006,N_10097);
nand U10451 (N_10451,N_10084,N_10067);
nand U10452 (N_10452,N_10124,N_10212);
or U10453 (N_10453,N_10074,N_10147);
or U10454 (N_10454,N_10240,N_10110);
nor U10455 (N_10455,N_10105,N_10088);
or U10456 (N_10456,N_10200,N_10097);
nor U10457 (N_10457,N_10031,N_10006);
xor U10458 (N_10458,N_10101,N_10109);
nor U10459 (N_10459,N_10157,N_10143);
nor U10460 (N_10460,N_10130,N_10122);
or U10461 (N_10461,N_10078,N_10131);
or U10462 (N_10462,N_10009,N_10081);
nand U10463 (N_10463,N_10127,N_10085);
xor U10464 (N_10464,N_10081,N_10232);
or U10465 (N_10465,N_10204,N_10055);
xnor U10466 (N_10466,N_10218,N_10067);
or U10467 (N_10467,N_10047,N_10138);
nor U10468 (N_10468,N_10145,N_10028);
xnor U10469 (N_10469,N_10134,N_10177);
and U10470 (N_10470,N_10187,N_10089);
xnor U10471 (N_10471,N_10082,N_10129);
and U10472 (N_10472,N_10093,N_10224);
or U10473 (N_10473,N_10093,N_10083);
nor U10474 (N_10474,N_10180,N_10142);
nand U10475 (N_10475,N_10181,N_10142);
xor U10476 (N_10476,N_10069,N_10042);
xnor U10477 (N_10477,N_10195,N_10225);
xnor U10478 (N_10478,N_10189,N_10218);
nor U10479 (N_10479,N_10101,N_10114);
nand U10480 (N_10480,N_10096,N_10089);
nand U10481 (N_10481,N_10154,N_10249);
or U10482 (N_10482,N_10136,N_10241);
nand U10483 (N_10483,N_10097,N_10188);
or U10484 (N_10484,N_10042,N_10130);
xnor U10485 (N_10485,N_10090,N_10051);
nand U10486 (N_10486,N_10113,N_10242);
xor U10487 (N_10487,N_10061,N_10129);
nor U10488 (N_10488,N_10215,N_10247);
and U10489 (N_10489,N_10024,N_10087);
nor U10490 (N_10490,N_10052,N_10220);
and U10491 (N_10491,N_10037,N_10237);
xor U10492 (N_10492,N_10187,N_10003);
nor U10493 (N_10493,N_10170,N_10244);
xor U10494 (N_10494,N_10181,N_10135);
and U10495 (N_10495,N_10211,N_10150);
xor U10496 (N_10496,N_10167,N_10162);
or U10497 (N_10497,N_10095,N_10099);
nand U10498 (N_10498,N_10008,N_10117);
and U10499 (N_10499,N_10075,N_10100);
and U10500 (N_10500,N_10415,N_10443);
or U10501 (N_10501,N_10371,N_10261);
xor U10502 (N_10502,N_10425,N_10323);
or U10503 (N_10503,N_10354,N_10473);
and U10504 (N_10504,N_10464,N_10360);
or U10505 (N_10505,N_10277,N_10375);
and U10506 (N_10506,N_10402,N_10389);
nor U10507 (N_10507,N_10343,N_10430);
xor U10508 (N_10508,N_10357,N_10484);
nand U10509 (N_10509,N_10385,N_10413);
and U10510 (N_10510,N_10376,N_10468);
or U10511 (N_10511,N_10374,N_10365);
and U10512 (N_10512,N_10363,N_10284);
or U10513 (N_10513,N_10315,N_10431);
xor U10514 (N_10514,N_10319,N_10251);
xor U10515 (N_10515,N_10423,N_10308);
nor U10516 (N_10516,N_10309,N_10373);
or U10517 (N_10517,N_10252,N_10451);
xor U10518 (N_10518,N_10460,N_10495);
nand U10519 (N_10519,N_10299,N_10419);
or U10520 (N_10520,N_10456,N_10401);
and U10521 (N_10521,N_10280,N_10429);
and U10522 (N_10522,N_10381,N_10480);
xnor U10523 (N_10523,N_10388,N_10259);
or U10524 (N_10524,N_10421,N_10379);
and U10525 (N_10525,N_10344,N_10338);
or U10526 (N_10526,N_10481,N_10270);
or U10527 (N_10527,N_10330,N_10477);
or U10528 (N_10528,N_10262,N_10314);
and U10529 (N_10529,N_10355,N_10485);
xor U10530 (N_10530,N_10351,N_10488);
and U10531 (N_10531,N_10457,N_10318);
nor U10532 (N_10532,N_10469,N_10298);
and U10533 (N_10533,N_10336,N_10254);
xor U10534 (N_10534,N_10367,N_10274);
nand U10535 (N_10535,N_10491,N_10417);
nand U10536 (N_10536,N_10493,N_10292);
or U10537 (N_10537,N_10387,N_10452);
or U10538 (N_10538,N_10487,N_10310);
xnor U10539 (N_10539,N_10332,N_10321);
xnor U10540 (N_10540,N_10348,N_10405);
xnor U10541 (N_10541,N_10478,N_10392);
or U10542 (N_10542,N_10303,N_10359);
nor U10543 (N_10543,N_10312,N_10275);
xnor U10544 (N_10544,N_10253,N_10337);
and U10545 (N_10545,N_10424,N_10483);
nand U10546 (N_10546,N_10448,N_10276);
and U10547 (N_10547,N_10449,N_10340);
nand U10548 (N_10548,N_10459,N_10300);
xnor U10549 (N_10549,N_10438,N_10324);
or U10550 (N_10550,N_10441,N_10263);
nand U10551 (N_10551,N_10442,N_10322);
nor U10552 (N_10552,N_10260,N_10326);
nor U10553 (N_10553,N_10497,N_10406);
and U10554 (N_10554,N_10472,N_10454);
nand U10555 (N_10555,N_10462,N_10268);
nor U10556 (N_10556,N_10409,N_10283);
or U10557 (N_10557,N_10297,N_10383);
nand U10558 (N_10558,N_10432,N_10285);
nor U10559 (N_10559,N_10437,N_10341);
xor U10560 (N_10560,N_10311,N_10320);
nand U10561 (N_10561,N_10411,N_10289);
and U10562 (N_10562,N_10279,N_10498);
nor U10563 (N_10563,N_10372,N_10331);
or U10564 (N_10564,N_10258,N_10418);
nor U10565 (N_10565,N_10307,N_10410);
nor U10566 (N_10566,N_10296,N_10403);
or U10567 (N_10567,N_10433,N_10272);
nand U10568 (N_10568,N_10269,N_10470);
xor U10569 (N_10569,N_10382,N_10486);
xor U10570 (N_10570,N_10368,N_10455);
or U10571 (N_10571,N_10306,N_10316);
nor U10572 (N_10572,N_10463,N_10444);
and U10573 (N_10573,N_10345,N_10290);
or U10574 (N_10574,N_10352,N_10339);
nand U10575 (N_10575,N_10302,N_10386);
and U10576 (N_10576,N_10362,N_10428);
nor U10577 (N_10577,N_10445,N_10346);
and U10578 (N_10578,N_10476,N_10400);
or U10579 (N_10579,N_10416,N_10396);
nand U10580 (N_10580,N_10466,N_10490);
nor U10581 (N_10581,N_10447,N_10328);
nand U10582 (N_10582,N_10333,N_10439);
nor U10583 (N_10583,N_10349,N_10356);
and U10584 (N_10584,N_10286,N_10364);
nor U10585 (N_10585,N_10391,N_10287);
nand U10586 (N_10586,N_10426,N_10271);
nand U10587 (N_10587,N_10369,N_10407);
and U10588 (N_10588,N_10397,N_10325);
xor U10589 (N_10589,N_10334,N_10264);
nor U10590 (N_10590,N_10335,N_10499);
and U10591 (N_10591,N_10398,N_10265);
nand U10592 (N_10592,N_10453,N_10446);
or U10593 (N_10593,N_10390,N_10278);
nor U10594 (N_10594,N_10380,N_10420);
or U10595 (N_10595,N_10347,N_10267);
and U10596 (N_10596,N_10305,N_10288);
nor U10597 (N_10597,N_10291,N_10293);
and U10598 (N_10598,N_10378,N_10301);
and U10599 (N_10599,N_10329,N_10294);
nor U10600 (N_10600,N_10327,N_10450);
nor U10601 (N_10601,N_10479,N_10496);
xnor U10602 (N_10602,N_10361,N_10358);
nand U10603 (N_10603,N_10494,N_10250);
or U10604 (N_10604,N_10366,N_10458);
or U10605 (N_10605,N_10257,N_10474);
or U10606 (N_10606,N_10467,N_10404);
and U10607 (N_10607,N_10434,N_10377);
or U10608 (N_10608,N_10422,N_10435);
nor U10609 (N_10609,N_10482,N_10412);
and U10610 (N_10610,N_10273,N_10436);
and U10611 (N_10611,N_10394,N_10282);
xnor U10612 (N_10612,N_10489,N_10313);
or U10613 (N_10613,N_10256,N_10492);
nor U10614 (N_10614,N_10342,N_10471);
xnor U10615 (N_10615,N_10427,N_10281);
or U10616 (N_10616,N_10295,N_10393);
or U10617 (N_10617,N_10395,N_10399);
xnor U10618 (N_10618,N_10461,N_10255);
nor U10619 (N_10619,N_10370,N_10440);
xor U10620 (N_10620,N_10266,N_10350);
and U10621 (N_10621,N_10414,N_10475);
xor U10622 (N_10622,N_10408,N_10384);
or U10623 (N_10623,N_10317,N_10353);
and U10624 (N_10624,N_10304,N_10465);
and U10625 (N_10625,N_10343,N_10394);
nand U10626 (N_10626,N_10427,N_10349);
xor U10627 (N_10627,N_10266,N_10303);
and U10628 (N_10628,N_10368,N_10280);
xnor U10629 (N_10629,N_10257,N_10442);
xor U10630 (N_10630,N_10327,N_10439);
nand U10631 (N_10631,N_10488,N_10380);
nand U10632 (N_10632,N_10479,N_10378);
nand U10633 (N_10633,N_10459,N_10281);
nand U10634 (N_10634,N_10419,N_10340);
and U10635 (N_10635,N_10475,N_10498);
xor U10636 (N_10636,N_10285,N_10485);
nor U10637 (N_10637,N_10491,N_10458);
nor U10638 (N_10638,N_10438,N_10466);
xnor U10639 (N_10639,N_10478,N_10321);
nor U10640 (N_10640,N_10375,N_10286);
and U10641 (N_10641,N_10337,N_10355);
nor U10642 (N_10642,N_10451,N_10337);
xnor U10643 (N_10643,N_10352,N_10295);
nor U10644 (N_10644,N_10418,N_10311);
xnor U10645 (N_10645,N_10445,N_10391);
xnor U10646 (N_10646,N_10252,N_10400);
nor U10647 (N_10647,N_10462,N_10495);
nor U10648 (N_10648,N_10408,N_10374);
xnor U10649 (N_10649,N_10400,N_10292);
nor U10650 (N_10650,N_10284,N_10273);
nor U10651 (N_10651,N_10443,N_10319);
and U10652 (N_10652,N_10436,N_10471);
xor U10653 (N_10653,N_10292,N_10485);
and U10654 (N_10654,N_10291,N_10395);
nor U10655 (N_10655,N_10295,N_10273);
and U10656 (N_10656,N_10397,N_10369);
xnor U10657 (N_10657,N_10415,N_10420);
or U10658 (N_10658,N_10365,N_10289);
xnor U10659 (N_10659,N_10308,N_10268);
nand U10660 (N_10660,N_10490,N_10430);
nand U10661 (N_10661,N_10395,N_10282);
xor U10662 (N_10662,N_10318,N_10426);
nor U10663 (N_10663,N_10411,N_10372);
nor U10664 (N_10664,N_10459,N_10444);
and U10665 (N_10665,N_10292,N_10291);
or U10666 (N_10666,N_10435,N_10463);
nor U10667 (N_10667,N_10481,N_10395);
xnor U10668 (N_10668,N_10261,N_10400);
and U10669 (N_10669,N_10278,N_10370);
nor U10670 (N_10670,N_10269,N_10445);
and U10671 (N_10671,N_10288,N_10423);
xnor U10672 (N_10672,N_10360,N_10452);
and U10673 (N_10673,N_10452,N_10388);
nor U10674 (N_10674,N_10440,N_10358);
xnor U10675 (N_10675,N_10496,N_10332);
xor U10676 (N_10676,N_10366,N_10377);
nand U10677 (N_10677,N_10319,N_10395);
nor U10678 (N_10678,N_10364,N_10389);
and U10679 (N_10679,N_10423,N_10294);
and U10680 (N_10680,N_10267,N_10346);
nor U10681 (N_10681,N_10377,N_10354);
xor U10682 (N_10682,N_10307,N_10272);
nand U10683 (N_10683,N_10262,N_10392);
or U10684 (N_10684,N_10444,N_10380);
nor U10685 (N_10685,N_10397,N_10464);
nand U10686 (N_10686,N_10335,N_10312);
and U10687 (N_10687,N_10451,N_10319);
or U10688 (N_10688,N_10360,N_10446);
nand U10689 (N_10689,N_10464,N_10316);
or U10690 (N_10690,N_10495,N_10404);
xnor U10691 (N_10691,N_10290,N_10368);
xnor U10692 (N_10692,N_10494,N_10381);
xnor U10693 (N_10693,N_10325,N_10357);
nor U10694 (N_10694,N_10378,N_10390);
or U10695 (N_10695,N_10393,N_10461);
or U10696 (N_10696,N_10330,N_10496);
and U10697 (N_10697,N_10389,N_10499);
nand U10698 (N_10698,N_10392,N_10282);
nor U10699 (N_10699,N_10384,N_10321);
and U10700 (N_10700,N_10339,N_10273);
and U10701 (N_10701,N_10477,N_10475);
and U10702 (N_10702,N_10467,N_10425);
or U10703 (N_10703,N_10491,N_10447);
xnor U10704 (N_10704,N_10297,N_10273);
xnor U10705 (N_10705,N_10375,N_10291);
nand U10706 (N_10706,N_10375,N_10335);
xnor U10707 (N_10707,N_10281,N_10289);
nor U10708 (N_10708,N_10472,N_10387);
nand U10709 (N_10709,N_10473,N_10474);
xnor U10710 (N_10710,N_10336,N_10355);
or U10711 (N_10711,N_10397,N_10437);
xnor U10712 (N_10712,N_10387,N_10271);
nor U10713 (N_10713,N_10490,N_10378);
and U10714 (N_10714,N_10499,N_10310);
nor U10715 (N_10715,N_10348,N_10327);
and U10716 (N_10716,N_10297,N_10321);
and U10717 (N_10717,N_10494,N_10391);
nand U10718 (N_10718,N_10479,N_10324);
xor U10719 (N_10719,N_10254,N_10308);
nand U10720 (N_10720,N_10251,N_10294);
and U10721 (N_10721,N_10491,N_10440);
or U10722 (N_10722,N_10427,N_10416);
and U10723 (N_10723,N_10351,N_10370);
and U10724 (N_10724,N_10276,N_10365);
and U10725 (N_10725,N_10354,N_10375);
or U10726 (N_10726,N_10346,N_10271);
nand U10727 (N_10727,N_10373,N_10403);
nand U10728 (N_10728,N_10297,N_10452);
nor U10729 (N_10729,N_10396,N_10304);
nor U10730 (N_10730,N_10286,N_10307);
xnor U10731 (N_10731,N_10493,N_10414);
and U10732 (N_10732,N_10308,N_10432);
or U10733 (N_10733,N_10371,N_10312);
or U10734 (N_10734,N_10312,N_10420);
or U10735 (N_10735,N_10459,N_10397);
and U10736 (N_10736,N_10328,N_10298);
xnor U10737 (N_10737,N_10438,N_10388);
xor U10738 (N_10738,N_10324,N_10329);
xor U10739 (N_10739,N_10373,N_10462);
and U10740 (N_10740,N_10467,N_10279);
or U10741 (N_10741,N_10374,N_10364);
and U10742 (N_10742,N_10445,N_10354);
nor U10743 (N_10743,N_10469,N_10447);
and U10744 (N_10744,N_10441,N_10342);
nor U10745 (N_10745,N_10389,N_10379);
or U10746 (N_10746,N_10346,N_10349);
and U10747 (N_10747,N_10341,N_10295);
or U10748 (N_10748,N_10252,N_10423);
or U10749 (N_10749,N_10397,N_10284);
xor U10750 (N_10750,N_10643,N_10570);
xnor U10751 (N_10751,N_10745,N_10612);
xor U10752 (N_10752,N_10529,N_10700);
nand U10753 (N_10753,N_10602,N_10569);
and U10754 (N_10754,N_10607,N_10559);
xnor U10755 (N_10755,N_10621,N_10568);
and U10756 (N_10756,N_10699,N_10705);
nor U10757 (N_10757,N_10601,N_10566);
nand U10758 (N_10758,N_10723,N_10671);
nand U10759 (N_10759,N_10544,N_10692);
and U10760 (N_10760,N_10708,N_10632);
or U10761 (N_10761,N_10684,N_10517);
nand U10762 (N_10762,N_10717,N_10626);
and U10763 (N_10763,N_10653,N_10500);
and U10764 (N_10764,N_10552,N_10604);
xor U10765 (N_10765,N_10744,N_10651);
and U10766 (N_10766,N_10514,N_10625);
nor U10767 (N_10767,N_10659,N_10713);
nor U10768 (N_10768,N_10518,N_10715);
or U10769 (N_10769,N_10526,N_10513);
or U10770 (N_10770,N_10593,N_10637);
or U10771 (N_10771,N_10528,N_10524);
xor U10772 (N_10772,N_10596,N_10688);
xnor U10773 (N_10773,N_10535,N_10660);
nor U10774 (N_10774,N_10633,N_10698);
nand U10775 (N_10775,N_10606,N_10550);
or U10776 (N_10776,N_10507,N_10690);
nor U10777 (N_10777,N_10649,N_10622);
and U10778 (N_10778,N_10648,N_10561);
nor U10779 (N_10779,N_10576,N_10672);
and U10780 (N_10780,N_10541,N_10650);
or U10781 (N_10781,N_10691,N_10595);
xnor U10782 (N_10782,N_10610,N_10512);
nor U10783 (N_10783,N_10530,N_10666);
nand U10784 (N_10784,N_10718,N_10635);
nand U10785 (N_10785,N_10729,N_10597);
nor U10786 (N_10786,N_10532,N_10712);
and U10787 (N_10787,N_10673,N_10686);
nand U10788 (N_10788,N_10710,N_10581);
xnor U10789 (N_10789,N_10640,N_10669);
xor U10790 (N_10790,N_10516,N_10732);
nand U10791 (N_10791,N_10628,N_10676);
and U10792 (N_10792,N_10742,N_10703);
or U10793 (N_10793,N_10582,N_10682);
xor U10794 (N_10794,N_10583,N_10521);
and U10795 (N_10795,N_10501,N_10531);
or U10796 (N_10796,N_10548,N_10656);
nor U10797 (N_10797,N_10525,N_10587);
xor U10798 (N_10798,N_10667,N_10670);
nand U10799 (N_10799,N_10685,N_10733);
and U10800 (N_10800,N_10590,N_10749);
nor U10801 (N_10801,N_10617,N_10665);
nor U10802 (N_10802,N_10502,N_10679);
nand U10803 (N_10803,N_10573,N_10549);
nand U10804 (N_10804,N_10722,N_10592);
and U10805 (N_10805,N_10724,N_10735);
or U10806 (N_10806,N_10564,N_10618);
nand U10807 (N_10807,N_10695,N_10748);
nor U10808 (N_10808,N_10726,N_10509);
and U10809 (N_10809,N_10589,N_10603);
nor U10810 (N_10810,N_10580,N_10681);
and U10811 (N_10811,N_10563,N_10701);
and U10812 (N_10812,N_10615,N_10533);
or U10813 (N_10813,N_10731,N_10645);
or U10814 (N_10814,N_10508,N_10664);
nand U10815 (N_10815,N_10702,N_10554);
and U10816 (N_10816,N_10584,N_10599);
nand U10817 (N_10817,N_10738,N_10646);
nand U10818 (N_10818,N_10697,N_10553);
or U10819 (N_10819,N_10678,N_10709);
nand U10820 (N_10820,N_10539,N_10503);
and U10821 (N_10821,N_10739,N_10620);
xor U10822 (N_10822,N_10694,N_10523);
xor U10823 (N_10823,N_10630,N_10647);
xnor U10824 (N_10824,N_10641,N_10668);
xnor U10825 (N_10825,N_10661,N_10683);
nor U10826 (N_10826,N_10510,N_10736);
xor U10827 (N_10827,N_10662,N_10560);
and U10828 (N_10828,N_10588,N_10652);
nor U10829 (N_10829,N_10727,N_10556);
nand U10830 (N_10830,N_10574,N_10687);
and U10831 (N_10831,N_10614,N_10693);
and U10832 (N_10832,N_10627,N_10545);
nor U10833 (N_10833,N_10734,N_10740);
xor U10834 (N_10834,N_10600,N_10707);
xor U10835 (N_10835,N_10585,N_10543);
xor U10836 (N_10836,N_10711,N_10675);
or U10837 (N_10837,N_10706,N_10655);
nor U10838 (N_10838,N_10639,N_10663);
nor U10839 (N_10839,N_10657,N_10540);
and U10840 (N_10840,N_10537,N_10730);
and U10841 (N_10841,N_10565,N_10506);
xnor U10842 (N_10842,N_10598,N_10538);
or U10843 (N_10843,N_10624,N_10551);
nand U10844 (N_10844,N_10546,N_10746);
or U10845 (N_10845,N_10611,N_10747);
nor U10846 (N_10846,N_10642,N_10578);
nand U10847 (N_10847,N_10572,N_10674);
and U10848 (N_10848,N_10536,N_10534);
or U10849 (N_10849,N_10605,N_10623);
or U10850 (N_10850,N_10558,N_10555);
xor U10851 (N_10851,N_10577,N_10504);
and U10852 (N_10852,N_10571,N_10579);
xnor U10853 (N_10853,N_10519,N_10644);
or U10854 (N_10854,N_10562,N_10720);
nor U10855 (N_10855,N_10696,N_10638);
and U10856 (N_10856,N_10704,N_10658);
xnor U10857 (N_10857,N_10608,N_10609);
nor U10858 (N_10858,N_10616,N_10586);
xor U10859 (N_10859,N_10636,N_10542);
or U10860 (N_10860,N_10721,N_10520);
nor U10861 (N_10861,N_10631,N_10728);
nor U10862 (N_10862,N_10680,N_10591);
nor U10863 (N_10863,N_10619,N_10527);
xnor U10864 (N_10864,N_10515,N_10567);
nand U10865 (N_10865,N_10689,N_10505);
xor U10866 (N_10866,N_10575,N_10719);
or U10867 (N_10867,N_10594,N_10522);
and U10868 (N_10868,N_10511,N_10654);
xnor U10869 (N_10869,N_10725,N_10716);
and U10870 (N_10870,N_10547,N_10613);
or U10871 (N_10871,N_10714,N_10741);
nand U10872 (N_10872,N_10677,N_10743);
nand U10873 (N_10873,N_10634,N_10629);
and U10874 (N_10874,N_10557,N_10737);
nor U10875 (N_10875,N_10631,N_10644);
and U10876 (N_10876,N_10719,N_10695);
and U10877 (N_10877,N_10534,N_10587);
xor U10878 (N_10878,N_10737,N_10639);
xor U10879 (N_10879,N_10623,N_10594);
xnor U10880 (N_10880,N_10630,N_10555);
and U10881 (N_10881,N_10616,N_10647);
xnor U10882 (N_10882,N_10709,N_10629);
xnor U10883 (N_10883,N_10516,N_10523);
nor U10884 (N_10884,N_10605,N_10696);
nand U10885 (N_10885,N_10503,N_10548);
xor U10886 (N_10886,N_10606,N_10697);
nor U10887 (N_10887,N_10696,N_10503);
nor U10888 (N_10888,N_10501,N_10719);
nand U10889 (N_10889,N_10543,N_10530);
nor U10890 (N_10890,N_10500,N_10503);
or U10891 (N_10891,N_10739,N_10547);
nand U10892 (N_10892,N_10682,N_10698);
nand U10893 (N_10893,N_10743,N_10558);
xor U10894 (N_10894,N_10680,N_10551);
xor U10895 (N_10895,N_10613,N_10555);
and U10896 (N_10896,N_10551,N_10534);
or U10897 (N_10897,N_10677,N_10642);
or U10898 (N_10898,N_10724,N_10707);
xnor U10899 (N_10899,N_10515,N_10514);
nand U10900 (N_10900,N_10507,N_10684);
nor U10901 (N_10901,N_10684,N_10526);
and U10902 (N_10902,N_10596,N_10699);
xnor U10903 (N_10903,N_10509,N_10566);
nand U10904 (N_10904,N_10565,N_10514);
and U10905 (N_10905,N_10685,N_10593);
or U10906 (N_10906,N_10588,N_10747);
and U10907 (N_10907,N_10509,N_10610);
or U10908 (N_10908,N_10570,N_10608);
xor U10909 (N_10909,N_10519,N_10675);
nor U10910 (N_10910,N_10521,N_10577);
xor U10911 (N_10911,N_10644,N_10590);
nand U10912 (N_10912,N_10553,N_10621);
nor U10913 (N_10913,N_10530,N_10624);
nor U10914 (N_10914,N_10541,N_10583);
xnor U10915 (N_10915,N_10591,N_10565);
and U10916 (N_10916,N_10708,N_10506);
xor U10917 (N_10917,N_10614,N_10726);
nor U10918 (N_10918,N_10529,N_10663);
nand U10919 (N_10919,N_10587,N_10664);
and U10920 (N_10920,N_10662,N_10716);
xnor U10921 (N_10921,N_10599,N_10512);
or U10922 (N_10922,N_10618,N_10658);
and U10923 (N_10923,N_10570,N_10518);
and U10924 (N_10924,N_10510,N_10649);
or U10925 (N_10925,N_10645,N_10633);
nor U10926 (N_10926,N_10628,N_10511);
and U10927 (N_10927,N_10555,N_10697);
and U10928 (N_10928,N_10593,N_10554);
or U10929 (N_10929,N_10540,N_10665);
or U10930 (N_10930,N_10706,N_10698);
nand U10931 (N_10931,N_10550,N_10500);
nand U10932 (N_10932,N_10629,N_10664);
nand U10933 (N_10933,N_10748,N_10678);
and U10934 (N_10934,N_10525,N_10575);
and U10935 (N_10935,N_10707,N_10573);
nand U10936 (N_10936,N_10674,N_10707);
xnor U10937 (N_10937,N_10525,N_10663);
xnor U10938 (N_10938,N_10692,N_10667);
xor U10939 (N_10939,N_10658,N_10659);
and U10940 (N_10940,N_10646,N_10535);
or U10941 (N_10941,N_10724,N_10520);
nor U10942 (N_10942,N_10521,N_10626);
or U10943 (N_10943,N_10584,N_10713);
or U10944 (N_10944,N_10539,N_10743);
xnor U10945 (N_10945,N_10556,N_10690);
or U10946 (N_10946,N_10709,N_10675);
or U10947 (N_10947,N_10716,N_10704);
and U10948 (N_10948,N_10505,N_10693);
nand U10949 (N_10949,N_10689,N_10730);
and U10950 (N_10950,N_10588,N_10575);
and U10951 (N_10951,N_10748,N_10559);
nand U10952 (N_10952,N_10585,N_10672);
and U10953 (N_10953,N_10712,N_10505);
and U10954 (N_10954,N_10542,N_10674);
xor U10955 (N_10955,N_10676,N_10626);
xnor U10956 (N_10956,N_10545,N_10501);
xor U10957 (N_10957,N_10723,N_10748);
xnor U10958 (N_10958,N_10551,N_10562);
or U10959 (N_10959,N_10731,N_10723);
or U10960 (N_10960,N_10502,N_10708);
or U10961 (N_10961,N_10574,N_10655);
nand U10962 (N_10962,N_10711,N_10580);
or U10963 (N_10963,N_10688,N_10561);
or U10964 (N_10964,N_10525,N_10729);
nand U10965 (N_10965,N_10554,N_10630);
and U10966 (N_10966,N_10546,N_10610);
and U10967 (N_10967,N_10599,N_10529);
and U10968 (N_10968,N_10551,N_10661);
nor U10969 (N_10969,N_10698,N_10665);
nand U10970 (N_10970,N_10700,N_10668);
xor U10971 (N_10971,N_10504,N_10744);
and U10972 (N_10972,N_10614,N_10569);
nor U10973 (N_10973,N_10539,N_10580);
and U10974 (N_10974,N_10552,N_10661);
nor U10975 (N_10975,N_10544,N_10600);
xnor U10976 (N_10976,N_10643,N_10652);
nand U10977 (N_10977,N_10693,N_10566);
or U10978 (N_10978,N_10735,N_10677);
or U10979 (N_10979,N_10744,N_10671);
xor U10980 (N_10980,N_10573,N_10566);
xor U10981 (N_10981,N_10714,N_10545);
nor U10982 (N_10982,N_10508,N_10630);
nor U10983 (N_10983,N_10651,N_10712);
and U10984 (N_10984,N_10662,N_10562);
nor U10985 (N_10985,N_10569,N_10565);
and U10986 (N_10986,N_10745,N_10641);
and U10987 (N_10987,N_10735,N_10584);
nor U10988 (N_10988,N_10637,N_10706);
xor U10989 (N_10989,N_10640,N_10630);
nor U10990 (N_10990,N_10691,N_10725);
and U10991 (N_10991,N_10741,N_10506);
nor U10992 (N_10992,N_10556,N_10671);
xor U10993 (N_10993,N_10646,N_10607);
and U10994 (N_10994,N_10696,N_10599);
xor U10995 (N_10995,N_10507,N_10583);
nand U10996 (N_10996,N_10652,N_10514);
xnor U10997 (N_10997,N_10514,N_10731);
nand U10998 (N_10998,N_10654,N_10546);
nand U10999 (N_10999,N_10539,N_10575);
and U11000 (N_11000,N_10907,N_10930);
xor U11001 (N_11001,N_10796,N_10923);
and U11002 (N_11002,N_10925,N_10883);
and U11003 (N_11003,N_10965,N_10833);
xnor U11004 (N_11004,N_10958,N_10910);
or U11005 (N_11005,N_10757,N_10808);
or U11006 (N_11006,N_10999,N_10998);
nand U11007 (N_11007,N_10760,N_10820);
nand U11008 (N_11008,N_10886,N_10946);
nor U11009 (N_11009,N_10920,N_10981);
nor U11010 (N_11010,N_10761,N_10991);
nor U11011 (N_11011,N_10764,N_10750);
or U11012 (N_11012,N_10976,N_10982);
and U11013 (N_11013,N_10824,N_10900);
nand U11014 (N_11014,N_10873,N_10966);
nor U11015 (N_11015,N_10924,N_10852);
nor U11016 (N_11016,N_10983,N_10850);
nand U11017 (N_11017,N_10768,N_10839);
xor U11018 (N_11018,N_10967,N_10904);
nand U11019 (N_11019,N_10832,N_10866);
or U11020 (N_11020,N_10985,N_10987);
nand U11021 (N_11021,N_10960,N_10812);
nor U11022 (N_11022,N_10955,N_10937);
or U11023 (N_11023,N_10962,N_10766);
or U11024 (N_11024,N_10860,N_10804);
nor U11025 (N_11025,N_10959,N_10936);
nor U11026 (N_11026,N_10989,N_10783);
or U11027 (N_11027,N_10969,N_10977);
nor U11028 (N_11028,N_10993,N_10971);
nor U11029 (N_11029,N_10836,N_10954);
xnor U11030 (N_11030,N_10891,N_10885);
xnor U11031 (N_11031,N_10805,N_10827);
nor U11032 (N_11032,N_10895,N_10919);
xor U11033 (N_11033,N_10874,N_10818);
and U11034 (N_11034,N_10849,N_10879);
xor U11035 (N_11035,N_10821,N_10806);
or U11036 (N_11036,N_10775,N_10935);
nor U11037 (N_11037,N_10945,N_10964);
or U11038 (N_11038,N_10884,N_10961);
or U11039 (N_11039,N_10845,N_10858);
nor U11040 (N_11040,N_10974,N_10751);
nand U11041 (N_11041,N_10765,N_10933);
and U11042 (N_11042,N_10938,N_10787);
nor U11043 (N_11043,N_10917,N_10830);
xnor U11044 (N_11044,N_10892,N_10888);
or U11045 (N_11045,N_10815,N_10986);
nand U11046 (N_11046,N_10857,N_10844);
xor U11047 (N_11047,N_10791,N_10831);
nand U11048 (N_11048,N_10887,N_10995);
nor U11049 (N_11049,N_10784,N_10973);
nand U11050 (N_11050,N_10863,N_10842);
nand U11051 (N_11051,N_10763,N_10828);
xnor U11052 (N_11052,N_10841,N_10855);
nand U11053 (N_11053,N_10869,N_10931);
xnor U11054 (N_11054,N_10947,N_10780);
or U11055 (N_11055,N_10984,N_10755);
and U11056 (N_11056,N_10898,N_10968);
and U11057 (N_11057,N_10978,N_10943);
and U11058 (N_11058,N_10880,N_10810);
xor U11059 (N_11059,N_10980,N_10809);
nand U11060 (N_11060,N_10890,N_10990);
nor U11061 (N_11061,N_10752,N_10903);
and U11062 (N_11062,N_10889,N_10778);
or U11063 (N_11063,N_10940,N_10926);
and U11064 (N_11064,N_10792,N_10758);
nor U11065 (N_11065,N_10905,N_10941);
xnor U11066 (N_11066,N_10862,N_10807);
nand U11067 (N_11067,N_10826,N_10846);
nor U11068 (N_11068,N_10944,N_10753);
or U11069 (N_11069,N_10882,N_10795);
nor U11070 (N_11070,N_10773,N_10918);
nand U11071 (N_11071,N_10922,N_10875);
and U11072 (N_11072,N_10909,N_10835);
and U11073 (N_11073,N_10988,N_10861);
nand U11074 (N_11074,N_10975,N_10851);
nand U11075 (N_11075,N_10756,N_10819);
or U11076 (N_11076,N_10929,N_10994);
nor U11077 (N_11077,N_10798,N_10848);
nand U11078 (N_11078,N_10899,N_10865);
nand U11079 (N_11079,N_10951,N_10913);
xor U11080 (N_11080,N_10782,N_10801);
or U11081 (N_11081,N_10825,N_10928);
xor U11082 (N_11082,N_10970,N_10871);
and U11083 (N_11083,N_10894,N_10878);
nand U11084 (N_11084,N_10811,N_10814);
and U11085 (N_11085,N_10754,N_10859);
or U11086 (N_11086,N_10876,N_10897);
nand U11087 (N_11087,N_10896,N_10800);
nor U11088 (N_11088,N_10816,N_10797);
and U11089 (N_11089,N_10762,N_10877);
nand U11090 (N_11090,N_10881,N_10785);
nor U11091 (N_11091,N_10992,N_10777);
nor U11092 (N_11092,N_10834,N_10906);
and U11093 (N_11093,N_10934,N_10759);
or U11094 (N_11094,N_10914,N_10956);
xnor U11095 (N_11095,N_10789,N_10823);
nor U11096 (N_11096,N_10912,N_10843);
or U11097 (N_11097,N_10864,N_10911);
or U11098 (N_11098,N_10948,N_10942);
or U11099 (N_11099,N_10953,N_10997);
nand U11100 (N_11100,N_10817,N_10867);
xor U11101 (N_11101,N_10829,N_10932);
nand U11102 (N_11102,N_10915,N_10803);
nand U11103 (N_11103,N_10972,N_10957);
nor U11104 (N_11104,N_10921,N_10779);
or U11105 (N_11105,N_10793,N_10794);
xnor U11106 (N_11106,N_10908,N_10769);
and U11107 (N_11107,N_10788,N_10979);
and U11108 (N_11108,N_10774,N_10799);
or U11109 (N_11109,N_10901,N_10868);
nor U11110 (N_11110,N_10902,N_10838);
and U11111 (N_11111,N_10802,N_10813);
nor U11112 (N_11112,N_10927,N_10916);
and U11113 (N_11113,N_10837,N_10949);
xnor U11114 (N_11114,N_10772,N_10939);
or U11115 (N_11115,N_10950,N_10847);
xor U11116 (N_11116,N_10776,N_10996);
nand U11117 (N_11117,N_10770,N_10856);
and U11118 (N_11118,N_10790,N_10853);
nand U11119 (N_11119,N_10963,N_10854);
xnor U11120 (N_11120,N_10781,N_10767);
xor U11121 (N_11121,N_10893,N_10872);
nand U11122 (N_11122,N_10870,N_10952);
nand U11123 (N_11123,N_10771,N_10786);
or U11124 (N_11124,N_10840,N_10822);
or U11125 (N_11125,N_10870,N_10776);
nor U11126 (N_11126,N_10885,N_10850);
and U11127 (N_11127,N_10782,N_10779);
or U11128 (N_11128,N_10949,N_10989);
or U11129 (N_11129,N_10902,N_10904);
nor U11130 (N_11130,N_10856,N_10861);
xor U11131 (N_11131,N_10922,N_10862);
and U11132 (N_11132,N_10769,N_10915);
nor U11133 (N_11133,N_10891,N_10775);
or U11134 (N_11134,N_10988,N_10883);
xnor U11135 (N_11135,N_10967,N_10765);
or U11136 (N_11136,N_10841,N_10943);
nand U11137 (N_11137,N_10989,N_10790);
and U11138 (N_11138,N_10882,N_10915);
nor U11139 (N_11139,N_10951,N_10985);
nand U11140 (N_11140,N_10907,N_10851);
nand U11141 (N_11141,N_10822,N_10879);
nor U11142 (N_11142,N_10854,N_10790);
and U11143 (N_11143,N_10796,N_10907);
xor U11144 (N_11144,N_10916,N_10998);
nor U11145 (N_11145,N_10985,N_10765);
nor U11146 (N_11146,N_10828,N_10792);
xor U11147 (N_11147,N_10927,N_10840);
nand U11148 (N_11148,N_10912,N_10945);
and U11149 (N_11149,N_10820,N_10877);
nand U11150 (N_11150,N_10892,N_10874);
or U11151 (N_11151,N_10931,N_10883);
xor U11152 (N_11152,N_10882,N_10930);
nor U11153 (N_11153,N_10994,N_10783);
nor U11154 (N_11154,N_10840,N_10753);
and U11155 (N_11155,N_10912,N_10947);
nand U11156 (N_11156,N_10769,N_10879);
and U11157 (N_11157,N_10975,N_10942);
or U11158 (N_11158,N_10812,N_10803);
nor U11159 (N_11159,N_10954,N_10801);
and U11160 (N_11160,N_10894,N_10985);
and U11161 (N_11161,N_10963,N_10972);
nand U11162 (N_11162,N_10918,N_10809);
nor U11163 (N_11163,N_10832,N_10810);
and U11164 (N_11164,N_10861,N_10877);
nand U11165 (N_11165,N_10770,N_10860);
nor U11166 (N_11166,N_10841,N_10806);
and U11167 (N_11167,N_10901,N_10927);
nand U11168 (N_11168,N_10901,N_10832);
nor U11169 (N_11169,N_10921,N_10930);
nor U11170 (N_11170,N_10869,N_10994);
and U11171 (N_11171,N_10956,N_10752);
xor U11172 (N_11172,N_10905,N_10878);
or U11173 (N_11173,N_10915,N_10844);
nand U11174 (N_11174,N_10861,N_10790);
or U11175 (N_11175,N_10967,N_10902);
or U11176 (N_11176,N_10959,N_10756);
nand U11177 (N_11177,N_10750,N_10779);
and U11178 (N_11178,N_10914,N_10989);
xnor U11179 (N_11179,N_10818,N_10887);
and U11180 (N_11180,N_10909,N_10965);
nor U11181 (N_11181,N_10883,N_10945);
nand U11182 (N_11182,N_10798,N_10966);
or U11183 (N_11183,N_10801,N_10876);
nor U11184 (N_11184,N_10815,N_10840);
or U11185 (N_11185,N_10824,N_10835);
and U11186 (N_11186,N_10852,N_10861);
nand U11187 (N_11187,N_10924,N_10964);
nor U11188 (N_11188,N_10752,N_10976);
and U11189 (N_11189,N_10821,N_10864);
nand U11190 (N_11190,N_10796,N_10874);
and U11191 (N_11191,N_10815,N_10868);
nand U11192 (N_11192,N_10804,N_10832);
nor U11193 (N_11193,N_10994,N_10766);
xnor U11194 (N_11194,N_10777,N_10860);
or U11195 (N_11195,N_10754,N_10866);
nand U11196 (N_11196,N_10808,N_10892);
nand U11197 (N_11197,N_10845,N_10889);
and U11198 (N_11198,N_10753,N_10765);
xnor U11199 (N_11199,N_10837,N_10778);
and U11200 (N_11200,N_10760,N_10879);
nor U11201 (N_11201,N_10819,N_10799);
or U11202 (N_11202,N_10902,N_10845);
and U11203 (N_11203,N_10809,N_10860);
nor U11204 (N_11204,N_10874,N_10764);
nor U11205 (N_11205,N_10852,N_10905);
nor U11206 (N_11206,N_10972,N_10889);
xnor U11207 (N_11207,N_10763,N_10799);
nor U11208 (N_11208,N_10815,N_10847);
nand U11209 (N_11209,N_10992,N_10932);
nor U11210 (N_11210,N_10931,N_10996);
nand U11211 (N_11211,N_10999,N_10917);
nor U11212 (N_11212,N_10831,N_10966);
and U11213 (N_11213,N_10787,N_10997);
or U11214 (N_11214,N_10830,N_10789);
nor U11215 (N_11215,N_10927,N_10907);
and U11216 (N_11216,N_10817,N_10960);
xor U11217 (N_11217,N_10978,N_10811);
and U11218 (N_11218,N_10846,N_10818);
xor U11219 (N_11219,N_10825,N_10778);
and U11220 (N_11220,N_10939,N_10781);
or U11221 (N_11221,N_10763,N_10893);
xnor U11222 (N_11222,N_10919,N_10975);
or U11223 (N_11223,N_10990,N_10802);
and U11224 (N_11224,N_10987,N_10929);
and U11225 (N_11225,N_10923,N_10964);
nand U11226 (N_11226,N_10978,N_10825);
xor U11227 (N_11227,N_10751,N_10885);
nor U11228 (N_11228,N_10804,N_10960);
xor U11229 (N_11229,N_10989,N_10873);
nor U11230 (N_11230,N_10795,N_10767);
nand U11231 (N_11231,N_10753,N_10824);
nand U11232 (N_11232,N_10876,N_10943);
xor U11233 (N_11233,N_10917,N_10865);
xnor U11234 (N_11234,N_10993,N_10956);
xor U11235 (N_11235,N_10878,N_10771);
and U11236 (N_11236,N_10829,N_10788);
xor U11237 (N_11237,N_10878,N_10993);
and U11238 (N_11238,N_10777,N_10961);
nand U11239 (N_11239,N_10806,N_10944);
nor U11240 (N_11240,N_10867,N_10769);
nor U11241 (N_11241,N_10831,N_10768);
and U11242 (N_11242,N_10846,N_10992);
or U11243 (N_11243,N_10948,N_10988);
xor U11244 (N_11244,N_10837,N_10871);
nor U11245 (N_11245,N_10941,N_10813);
nor U11246 (N_11246,N_10885,N_10896);
or U11247 (N_11247,N_10960,N_10854);
nand U11248 (N_11248,N_10785,N_10802);
nand U11249 (N_11249,N_10858,N_10838);
or U11250 (N_11250,N_11096,N_11152);
nor U11251 (N_11251,N_11157,N_11153);
nor U11252 (N_11252,N_11122,N_11180);
xnor U11253 (N_11253,N_11205,N_11033);
and U11254 (N_11254,N_11161,N_11210);
nand U11255 (N_11255,N_11069,N_11187);
and U11256 (N_11256,N_11068,N_11091);
or U11257 (N_11257,N_11075,N_11226);
nor U11258 (N_11258,N_11195,N_11162);
xnor U11259 (N_11259,N_11243,N_11028);
nor U11260 (N_11260,N_11006,N_11144);
nor U11261 (N_11261,N_11116,N_11125);
nand U11262 (N_11262,N_11023,N_11179);
nand U11263 (N_11263,N_11121,N_11192);
nand U11264 (N_11264,N_11127,N_11111);
xnor U11265 (N_11265,N_11124,N_11146);
nand U11266 (N_11266,N_11175,N_11126);
nor U11267 (N_11267,N_11246,N_11206);
nand U11268 (N_11268,N_11012,N_11099);
xnor U11269 (N_11269,N_11224,N_11200);
nand U11270 (N_11270,N_11040,N_11242);
and U11271 (N_11271,N_11035,N_11108);
nor U11272 (N_11272,N_11186,N_11154);
xnor U11273 (N_11273,N_11183,N_11016);
xor U11274 (N_11274,N_11148,N_11163);
and U11275 (N_11275,N_11042,N_11107);
and U11276 (N_11276,N_11184,N_11014);
xnor U11277 (N_11277,N_11201,N_11082);
nand U11278 (N_11278,N_11051,N_11238);
or U11279 (N_11279,N_11032,N_11249);
xor U11280 (N_11280,N_11139,N_11057);
or U11281 (N_11281,N_11156,N_11070);
and U11282 (N_11282,N_11106,N_11048);
nand U11283 (N_11283,N_11169,N_11209);
xnor U11284 (N_11284,N_11113,N_11245);
nand U11285 (N_11285,N_11248,N_11022);
xnor U11286 (N_11286,N_11076,N_11176);
nand U11287 (N_11287,N_11207,N_11149);
nand U11288 (N_11288,N_11208,N_11067);
or U11289 (N_11289,N_11086,N_11083);
xnor U11290 (N_11290,N_11109,N_11034);
or U11291 (N_11291,N_11142,N_11103);
xor U11292 (N_11292,N_11056,N_11232);
nor U11293 (N_11293,N_11030,N_11219);
xnor U11294 (N_11294,N_11204,N_11087);
or U11295 (N_11295,N_11138,N_11172);
nor U11296 (N_11296,N_11236,N_11053);
nand U11297 (N_11297,N_11101,N_11058);
or U11298 (N_11298,N_11079,N_11095);
xor U11299 (N_11299,N_11078,N_11001);
nor U11300 (N_11300,N_11047,N_11151);
nand U11301 (N_11301,N_11059,N_11160);
or U11302 (N_11302,N_11131,N_11196);
and U11303 (N_11303,N_11025,N_11158);
nor U11304 (N_11304,N_11165,N_11027);
xor U11305 (N_11305,N_11188,N_11159);
nand U11306 (N_11306,N_11054,N_11197);
nand U11307 (N_11307,N_11074,N_11228);
nor U11308 (N_11308,N_11223,N_11105);
and U11309 (N_11309,N_11050,N_11155);
nand U11310 (N_11310,N_11168,N_11136);
nand U11311 (N_11311,N_11063,N_11038);
and U11312 (N_11312,N_11120,N_11072);
nand U11313 (N_11313,N_11227,N_11071);
nand U11314 (N_11314,N_11150,N_11134);
nand U11315 (N_11315,N_11088,N_11164);
or U11316 (N_11316,N_11191,N_11044);
or U11317 (N_11317,N_11235,N_11066);
nand U11318 (N_11318,N_11026,N_11178);
and U11319 (N_11319,N_11190,N_11181);
nand U11320 (N_11320,N_11185,N_11216);
or U11321 (N_11321,N_11119,N_11129);
and U11322 (N_11322,N_11143,N_11231);
or U11323 (N_11323,N_11046,N_11189);
nand U11324 (N_11324,N_11017,N_11173);
nor U11325 (N_11325,N_11049,N_11128);
and U11326 (N_11326,N_11104,N_11110);
xor U11327 (N_11327,N_11080,N_11031);
nor U11328 (N_11328,N_11174,N_11112);
nand U11329 (N_11329,N_11199,N_11005);
nor U11330 (N_11330,N_11000,N_11130);
and U11331 (N_11331,N_11222,N_11182);
and U11332 (N_11332,N_11081,N_11177);
nor U11333 (N_11333,N_11247,N_11132);
nor U11334 (N_11334,N_11013,N_11092);
and U11335 (N_11335,N_11098,N_11003);
xnor U11336 (N_11336,N_11039,N_11221);
nand U11337 (N_11337,N_11037,N_11115);
nand U11338 (N_11338,N_11141,N_11041);
and U11339 (N_11339,N_11089,N_11011);
nand U11340 (N_11340,N_11093,N_11237);
and U11341 (N_11341,N_11020,N_11045);
nor U11342 (N_11342,N_11123,N_11090);
and U11343 (N_11343,N_11244,N_11052);
or U11344 (N_11344,N_11133,N_11215);
xnor U11345 (N_11345,N_11055,N_11214);
xnor U11346 (N_11346,N_11203,N_11036);
nand U11347 (N_11347,N_11193,N_11230);
nand U11348 (N_11348,N_11211,N_11225);
xnor U11349 (N_11349,N_11029,N_11217);
or U11350 (N_11350,N_11194,N_11114);
and U11351 (N_11351,N_11220,N_11018);
nand U11352 (N_11352,N_11145,N_11137);
or U11353 (N_11353,N_11117,N_11170);
and U11354 (N_11354,N_11213,N_11010);
xnor U11355 (N_11355,N_11097,N_11118);
xnor U11356 (N_11356,N_11140,N_11240);
and U11357 (N_11357,N_11021,N_11085);
nor U11358 (N_11358,N_11094,N_11004);
nor U11359 (N_11359,N_11147,N_11212);
xor U11360 (N_11360,N_11100,N_11202);
nand U11361 (N_11361,N_11229,N_11135);
nand U11362 (N_11362,N_11008,N_11009);
xor U11363 (N_11363,N_11241,N_11198);
nor U11364 (N_11364,N_11002,N_11171);
or U11365 (N_11365,N_11233,N_11015);
nand U11366 (N_11366,N_11060,N_11064);
and U11367 (N_11367,N_11084,N_11065);
and U11368 (N_11368,N_11102,N_11019);
xnor U11369 (N_11369,N_11239,N_11061);
nand U11370 (N_11370,N_11234,N_11024);
nor U11371 (N_11371,N_11062,N_11218);
nor U11372 (N_11372,N_11166,N_11073);
xnor U11373 (N_11373,N_11077,N_11167);
or U11374 (N_11374,N_11007,N_11043);
and U11375 (N_11375,N_11013,N_11035);
nor U11376 (N_11376,N_11188,N_11001);
nor U11377 (N_11377,N_11059,N_11203);
xor U11378 (N_11378,N_11231,N_11032);
nor U11379 (N_11379,N_11049,N_11075);
or U11380 (N_11380,N_11184,N_11154);
nand U11381 (N_11381,N_11034,N_11097);
xnor U11382 (N_11382,N_11054,N_11190);
nor U11383 (N_11383,N_11199,N_11103);
nor U11384 (N_11384,N_11162,N_11048);
nand U11385 (N_11385,N_11228,N_11028);
and U11386 (N_11386,N_11206,N_11013);
nor U11387 (N_11387,N_11027,N_11053);
xor U11388 (N_11388,N_11183,N_11221);
nor U11389 (N_11389,N_11089,N_11187);
xnor U11390 (N_11390,N_11159,N_11141);
and U11391 (N_11391,N_11212,N_11056);
or U11392 (N_11392,N_11240,N_11058);
and U11393 (N_11393,N_11176,N_11066);
and U11394 (N_11394,N_11173,N_11106);
nor U11395 (N_11395,N_11200,N_11226);
nand U11396 (N_11396,N_11065,N_11081);
nor U11397 (N_11397,N_11045,N_11247);
nor U11398 (N_11398,N_11043,N_11028);
or U11399 (N_11399,N_11142,N_11106);
nor U11400 (N_11400,N_11204,N_11001);
and U11401 (N_11401,N_11149,N_11150);
and U11402 (N_11402,N_11075,N_11120);
and U11403 (N_11403,N_11179,N_11111);
or U11404 (N_11404,N_11247,N_11099);
or U11405 (N_11405,N_11094,N_11068);
xor U11406 (N_11406,N_11129,N_11094);
and U11407 (N_11407,N_11011,N_11033);
nand U11408 (N_11408,N_11234,N_11118);
xnor U11409 (N_11409,N_11012,N_11036);
or U11410 (N_11410,N_11044,N_11085);
xor U11411 (N_11411,N_11228,N_11179);
and U11412 (N_11412,N_11060,N_11240);
nand U11413 (N_11413,N_11025,N_11248);
nor U11414 (N_11414,N_11136,N_11069);
xor U11415 (N_11415,N_11076,N_11237);
and U11416 (N_11416,N_11032,N_11180);
and U11417 (N_11417,N_11001,N_11115);
or U11418 (N_11418,N_11229,N_11074);
or U11419 (N_11419,N_11002,N_11006);
nor U11420 (N_11420,N_11021,N_11126);
nor U11421 (N_11421,N_11041,N_11137);
nand U11422 (N_11422,N_11141,N_11054);
xor U11423 (N_11423,N_11013,N_11149);
or U11424 (N_11424,N_11169,N_11050);
and U11425 (N_11425,N_11092,N_11184);
nor U11426 (N_11426,N_11185,N_11155);
xnor U11427 (N_11427,N_11104,N_11010);
nor U11428 (N_11428,N_11166,N_11225);
nor U11429 (N_11429,N_11051,N_11025);
and U11430 (N_11430,N_11189,N_11095);
or U11431 (N_11431,N_11129,N_11242);
and U11432 (N_11432,N_11111,N_11064);
or U11433 (N_11433,N_11128,N_11058);
nand U11434 (N_11434,N_11041,N_11145);
nand U11435 (N_11435,N_11057,N_11090);
xor U11436 (N_11436,N_11050,N_11022);
and U11437 (N_11437,N_11004,N_11215);
or U11438 (N_11438,N_11188,N_11055);
xnor U11439 (N_11439,N_11007,N_11150);
or U11440 (N_11440,N_11009,N_11214);
xor U11441 (N_11441,N_11046,N_11058);
or U11442 (N_11442,N_11096,N_11153);
nor U11443 (N_11443,N_11215,N_11182);
and U11444 (N_11444,N_11109,N_11107);
xnor U11445 (N_11445,N_11213,N_11118);
nor U11446 (N_11446,N_11101,N_11052);
and U11447 (N_11447,N_11098,N_11027);
and U11448 (N_11448,N_11087,N_11111);
and U11449 (N_11449,N_11118,N_11226);
and U11450 (N_11450,N_11042,N_11138);
xor U11451 (N_11451,N_11112,N_11096);
xor U11452 (N_11452,N_11183,N_11110);
nand U11453 (N_11453,N_11127,N_11053);
nand U11454 (N_11454,N_11178,N_11188);
nor U11455 (N_11455,N_11130,N_11212);
nor U11456 (N_11456,N_11100,N_11025);
nand U11457 (N_11457,N_11193,N_11062);
nor U11458 (N_11458,N_11013,N_11054);
nor U11459 (N_11459,N_11097,N_11036);
nor U11460 (N_11460,N_11037,N_11025);
or U11461 (N_11461,N_11236,N_11247);
and U11462 (N_11462,N_11214,N_11004);
and U11463 (N_11463,N_11179,N_11214);
xnor U11464 (N_11464,N_11082,N_11050);
or U11465 (N_11465,N_11044,N_11039);
nand U11466 (N_11466,N_11173,N_11034);
and U11467 (N_11467,N_11020,N_11010);
nand U11468 (N_11468,N_11113,N_11101);
nand U11469 (N_11469,N_11110,N_11200);
nor U11470 (N_11470,N_11166,N_11058);
xor U11471 (N_11471,N_11237,N_11086);
or U11472 (N_11472,N_11210,N_11154);
nor U11473 (N_11473,N_11014,N_11202);
xnor U11474 (N_11474,N_11110,N_11068);
or U11475 (N_11475,N_11023,N_11191);
nor U11476 (N_11476,N_11074,N_11044);
xnor U11477 (N_11477,N_11120,N_11156);
and U11478 (N_11478,N_11068,N_11167);
nand U11479 (N_11479,N_11002,N_11181);
nor U11480 (N_11480,N_11185,N_11183);
nor U11481 (N_11481,N_11014,N_11226);
xnor U11482 (N_11482,N_11084,N_11040);
and U11483 (N_11483,N_11019,N_11009);
nor U11484 (N_11484,N_11248,N_11047);
and U11485 (N_11485,N_11216,N_11010);
and U11486 (N_11486,N_11029,N_11155);
xor U11487 (N_11487,N_11079,N_11050);
nor U11488 (N_11488,N_11053,N_11241);
nor U11489 (N_11489,N_11145,N_11148);
or U11490 (N_11490,N_11103,N_11218);
xnor U11491 (N_11491,N_11112,N_11122);
or U11492 (N_11492,N_11007,N_11130);
nor U11493 (N_11493,N_11113,N_11170);
nand U11494 (N_11494,N_11060,N_11160);
nand U11495 (N_11495,N_11146,N_11022);
nand U11496 (N_11496,N_11206,N_11208);
or U11497 (N_11497,N_11195,N_11168);
xor U11498 (N_11498,N_11230,N_11021);
xor U11499 (N_11499,N_11095,N_11185);
or U11500 (N_11500,N_11413,N_11365);
or U11501 (N_11501,N_11266,N_11425);
nor U11502 (N_11502,N_11357,N_11279);
or U11503 (N_11503,N_11389,N_11320);
and U11504 (N_11504,N_11453,N_11264);
nand U11505 (N_11505,N_11498,N_11326);
or U11506 (N_11506,N_11407,N_11390);
xnor U11507 (N_11507,N_11341,N_11434);
nor U11508 (N_11508,N_11317,N_11386);
nor U11509 (N_11509,N_11415,N_11333);
and U11510 (N_11510,N_11487,N_11294);
nand U11511 (N_11511,N_11472,N_11420);
nor U11512 (N_11512,N_11358,N_11275);
nand U11513 (N_11513,N_11366,N_11342);
and U11514 (N_11514,N_11285,N_11426);
and U11515 (N_11515,N_11397,N_11381);
or U11516 (N_11516,N_11405,N_11374);
xnor U11517 (N_11517,N_11388,N_11402);
xor U11518 (N_11518,N_11488,N_11411);
xor U11519 (N_11519,N_11376,N_11297);
xnor U11520 (N_11520,N_11310,N_11471);
and U11521 (N_11521,N_11475,N_11322);
or U11522 (N_11522,N_11296,N_11336);
or U11523 (N_11523,N_11258,N_11451);
or U11524 (N_11524,N_11339,N_11346);
and U11525 (N_11525,N_11482,N_11491);
nor U11526 (N_11526,N_11465,N_11267);
nor U11527 (N_11527,N_11316,N_11394);
nand U11528 (N_11528,N_11458,N_11305);
or U11529 (N_11529,N_11486,N_11495);
nand U11530 (N_11530,N_11292,N_11309);
nand U11531 (N_11531,N_11259,N_11382);
or U11532 (N_11532,N_11327,N_11353);
or U11533 (N_11533,N_11470,N_11417);
and U11534 (N_11534,N_11436,N_11330);
nor U11535 (N_11535,N_11334,N_11485);
xnor U11536 (N_11536,N_11331,N_11449);
nor U11537 (N_11537,N_11340,N_11403);
nor U11538 (N_11538,N_11370,N_11489);
and U11539 (N_11539,N_11301,N_11396);
or U11540 (N_11540,N_11308,N_11429);
and U11541 (N_11541,N_11430,N_11328);
xor U11542 (N_11542,N_11363,N_11354);
and U11543 (N_11543,N_11469,N_11271);
nor U11544 (N_11544,N_11424,N_11461);
nor U11545 (N_11545,N_11319,N_11385);
or U11546 (N_11546,N_11355,N_11277);
and U11547 (N_11547,N_11398,N_11421);
nand U11548 (N_11548,N_11378,N_11287);
nand U11549 (N_11549,N_11373,N_11265);
and U11550 (N_11550,N_11454,N_11474);
nand U11551 (N_11551,N_11377,N_11293);
nor U11552 (N_11552,N_11312,N_11250);
or U11553 (N_11553,N_11414,N_11372);
nor U11554 (N_11554,N_11438,N_11300);
xnor U11555 (N_11555,N_11478,N_11416);
nand U11556 (N_11556,N_11337,N_11401);
xnor U11557 (N_11557,N_11443,N_11349);
or U11558 (N_11558,N_11352,N_11291);
nand U11559 (N_11559,N_11384,N_11400);
xnor U11560 (N_11560,N_11289,N_11280);
or U11561 (N_11561,N_11364,N_11383);
nand U11562 (N_11562,N_11410,N_11418);
and U11563 (N_11563,N_11332,N_11295);
and U11564 (N_11564,N_11253,N_11281);
and U11565 (N_11565,N_11404,N_11412);
or U11566 (N_11566,N_11367,N_11483);
nand U11567 (N_11567,N_11329,N_11387);
xnor U11568 (N_11568,N_11447,N_11439);
or U11569 (N_11569,N_11276,N_11392);
nor U11570 (N_11570,N_11255,N_11282);
and U11571 (N_11571,N_11419,N_11311);
and U11572 (N_11572,N_11252,N_11269);
nand U11573 (N_11573,N_11284,N_11379);
nand U11574 (N_11574,N_11359,N_11272);
and U11575 (N_11575,N_11318,N_11494);
nor U11576 (N_11576,N_11395,N_11440);
nor U11577 (N_11577,N_11362,N_11496);
or U11578 (N_11578,N_11497,N_11446);
or U11579 (N_11579,N_11302,N_11490);
and U11580 (N_11580,N_11423,N_11298);
xnor U11581 (N_11581,N_11473,N_11463);
xnor U11582 (N_11582,N_11441,N_11278);
xnor U11583 (N_11583,N_11462,N_11481);
and U11584 (N_11584,N_11314,N_11480);
and U11585 (N_11585,N_11257,N_11315);
nor U11586 (N_11586,N_11256,N_11468);
nor U11587 (N_11587,N_11290,N_11299);
nor U11588 (N_11588,N_11306,N_11369);
nand U11589 (N_11589,N_11325,N_11262);
and U11590 (N_11590,N_11324,N_11406);
and U11591 (N_11591,N_11459,N_11457);
xor U11592 (N_11592,N_11445,N_11452);
nand U11593 (N_11593,N_11273,N_11492);
nand U11594 (N_11594,N_11428,N_11260);
nor U11595 (N_11595,N_11391,N_11350);
nand U11596 (N_11596,N_11270,N_11288);
nor U11597 (N_11597,N_11466,N_11343);
nand U11598 (N_11598,N_11435,N_11450);
nor U11599 (N_11599,N_11476,N_11347);
nor U11600 (N_11600,N_11304,N_11261);
nand U11601 (N_11601,N_11393,N_11338);
xnor U11602 (N_11602,N_11427,N_11499);
and U11603 (N_11603,N_11408,N_11456);
nand U11604 (N_11604,N_11433,N_11254);
or U11605 (N_11605,N_11448,N_11335);
and U11606 (N_11606,N_11251,N_11348);
nor U11607 (N_11607,N_11307,N_11321);
xor U11608 (N_11608,N_11477,N_11380);
xnor U11609 (N_11609,N_11399,N_11437);
xor U11610 (N_11610,N_11442,N_11432);
nand U11611 (N_11611,N_11444,N_11493);
nand U11612 (N_11612,N_11351,N_11479);
xnor U11613 (N_11613,N_11345,N_11356);
nand U11614 (N_11614,N_11431,N_11375);
and U11615 (N_11615,N_11263,N_11360);
xor U11616 (N_11616,N_11283,N_11467);
xnor U11617 (N_11617,N_11274,N_11368);
nand U11618 (N_11618,N_11323,N_11371);
or U11619 (N_11619,N_11361,N_11313);
or U11620 (N_11620,N_11286,N_11455);
nor U11621 (N_11621,N_11344,N_11409);
or U11622 (N_11622,N_11484,N_11268);
or U11623 (N_11623,N_11460,N_11464);
and U11624 (N_11624,N_11303,N_11422);
or U11625 (N_11625,N_11480,N_11351);
xnor U11626 (N_11626,N_11414,N_11499);
or U11627 (N_11627,N_11260,N_11302);
or U11628 (N_11628,N_11423,N_11383);
or U11629 (N_11629,N_11437,N_11363);
nand U11630 (N_11630,N_11285,N_11397);
xor U11631 (N_11631,N_11412,N_11393);
nor U11632 (N_11632,N_11276,N_11418);
xnor U11633 (N_11633,N_11326,N_11305);
nand U11634 (N_11634,N_11251,N_11303);
and U11635 (N_11635,N_11446,N_11486);
xor U11636 (N_11636,N_11473,N_11373);
and U11637 (N_11637,N_11275,N_11412);
or U11638 (N_11638,N_11343,N_11475);
xor U11639 (N_11639,N_11388,N_11349);
or U11640 (N_11640,N_11434,N_11381);
nor U11641 (N_11641,N_11356,N_11418);
and U11642 (N_11642,N_11412,N_11421);
nor U11643 (N_11643,N_11274,N_11373);
or U11644 (N_11644,N_11253,N_11329);
nand U11645 (N_11645,N_11266,N_11364);
nor U11646 (N_11646,N_11484,N_11252);
and U11647 (N_11647,N_11304,N_11258);
nor U11648 (N_11648,N_11388,N_11359);
nand U11649 (N_11649,N_11492,N_11279);
nand U11650 (N_11650,N_11459,N_11296);
xor U11651 (N_11651,N_11299,N_11497);
xnor U11652 (N_11652,N_11485,N_11440);
nand U11653 (N_11653,N_11339,N_11296);
and U11654 (N_11654,N_11266,N_11329);
xnor U11655 (N_11655,N_11316,N_11330);
or U11656 (N_11656,N_11319,N_11454);
and U11657 (N_11657,N_11413,N_11444);
xnor U11658 (N_11658,N_11328,N_11295);
and U11659 (N_11659,N_11282,N_11413);
nor U11660 (N_11660,N_11314,N_11499);
nor U11661 (N_11661,N_11433,N_11307);
nor U11662 (N_11662,N_11391,N_11430);
nand U11663 (N_11663,N_11439,N_11426);
and U11664 (N_11664,N_11341,N_11296);
and U11665 (N_11665,N_11253,N_11493);
and U11666 (N_11666,N_11264,N_11408);
xor U11667 (N_11667,N_11448,N_11282);
or U11668 (N_11668,N_11292,N_11458);
nor U11669 (N_11669,N_11490,N_11433);
and U11670 (N_11670,N_11379,N_11357);
nand U11671 (N_11671,N_11417,N_11309);
nor U11672 (N_11672,N_11252,N_11370);
and U11673 (N_11673,N_11467,N_11323);
and U11674 (N_11674,N_11266,N_11316);
nand U11675 (N_11675,N_11301,N_11340);
nand U11676 (N_11676,N_11320,N_11407);
nand U11677 (N_11677,N_11310,N_11380);
and U11678 (N_11678,N_11322,N_11476);
xnor U11679 (N_11679,N_11367,N_11380);
or U11680 (N_11680,N_11412,N_11389);
or U11681 (N_11681,N_11411,N_11494);
nand U11682 (N_11682,N_11441,N_11393);
and U11683 (N_11683,N_11262,N_11447);
or U11684 (N_11684,N_11295,N_11390);
nor U11685 (N_11685,N_11372,N_11370);
and U11686 (N_11686,N_11291,N_11339);
and U11687 (N_11687,N_11317,N_11385);
xnor U11688 (N_11688,N_11439,N_11486);
or U11689 (N_11689,N_11411,N_11290);
and U11690 (N_11690,N_11293,N_11301);
xnor U11691 (N_11691,N_11261,N_11342);
xnor U11692 (N_11692,N_11470,N_11296);
or U11693 (N_11693,N_11408,N_11354);
nor U11694 (N_11694,N_11436,N_11307);
and U11695 (N_11695,N_11315,N_11343);
xor U11696 (N_11696,N_11426,N_11424);
nand U11697 (N_11697,N_11466,N_11280);
or U11698 (N_11698,N_11252,N_11330);
xor U11699 (N_11699,N_11466,N_11296);
nand U11700 (N_11700,N_11288,N_11363);
or U11701 (N_11701,N_11481,N_11260);
and U11702 (N_11702,N_11328,N_11406);
or U11703 (N_11703,N_11263,N_11464);
nor U11704 (N_11704,N_11289,N_11317);
xnor U11705 (N_11705,N_11459,N_11269);
or U11706 (N_11706,N_11428,N_11493);
nor U11707 (N_11707,N_11293,N_11488);
nand U11708 (N_11708,N_11388,N_11498);
xnor U11709 (N_11709,N_11375,N_11354);
or U11710 (N_11710,N_11324,N_11355);
xor U11711 (N_11711,N_11280,N_11467);
nand U11712 (N_11712,N_11362,N_11305);
nor U11713 (N_11713,N_11298,N_11260);
or U11714 (N_11714,N_11283,N_11391);
nor U11715 (N_11715,N_11477,N_11296);
and U11716 (N_11716,N_11316,N_11362);
or U11717 (N_11717,N_11417,N_11401);
nand U11718 (N_11718,N_11487,N_11250);
and U11719 (N_11719,N_11251,N_11466);
xor U11720 (N_11720,N_11301,N_11377);
xnor U11721 (N_11721,N_11252,N_11346);
nor U11722 (N_11722,N_11476,N_11267);
and U11723 (N_11723,N_11467,N_11474);
xnor U11724 (N_11724,N_11455,N_11376);
xnor U11725 (N_11725,N_11250,N_11351);
xor U11726 (N_11726,N_11304,N_11337);
nor U11727 (N_11727,N_11411,N_11256);
and U11728 (N_11728,N_11370,N_11330);
nor U11729 (N_11729,N_11419,N_11267);
or U11730 (N_11730,N_11497,N_11290);
nor U11731 (N_11731,N_11438,N_11420);
nand U11732 (N_11732,N_11303,N_11298);
nand U11733 (N_11733,N_11272,N_11435);
nor U11734 (N_11734,N_11424,N_11352);
xnor U11735 (N_11735,N_11279,N_11351);
nand U11736 (N_11736,N_11483,N_11473);
nand U11737 (N_11737,N_11299,N_11348);
xor U11738 (N_11738,N_11484,N_11343);
and U11739 (N_11739,N_11446,N_11261);
or U11740 (N_11740,N_11367,N_11455);
nand U11741 (N_11741,N_11436,N_11454);
or U11742 (N_11742,N_11273,N_11428);
nor U11743 (N_11743,N_11467,N_11356);
nand U11744 (N_11744,N_11406,N_11289);
nand U11745 (N_11745,N_11367,N_11454);
nor U11746 (N_11746,N_11457,N_11464);
and U11747 (N_11747,N_11315,N_11298);
or U11748 (N_11748,N_11437,N_11273);
or U11749 (N_11749,N_11282,N_11488);
and U11750 (N_11750,N_11584,N_11520);
xnor U11751 (N_11751,N_11658,N_11716);
nor U11752 (N_11752,N_11577,N_11605);
xnor U11753 (N_11753,N_11656,N_11714);
or U11754 (N_11754,N_11504,N_11612);
xor U11755 (N_11755,N_11683,N_11553);
and U11756 (N_11756,N_11527,N_11704);
nor U11757 (N_11757,N_11549,N_11544);
or U11758 (N_11758,N_11503,N_11691);
xnor U11759 (N_11759,N_11705,N_11611);
and U11760 (N_11760,N_11719,N_11635);
and U11761 (N_11761,N_11746,N_11508);
xor U11762 (N_11762,N_11685,N_11689);
or U11763 (N_11763,N_11540,N_11608);
xor U11764 (N_11764,N_11668,N_11614);
and U11765 (N_11765,N_11695,N_11600);
xor U11766 (N_11766,N_11736,N_11715);
and U11767 (N_11767,N_11517,N_11519);
or U11768 (N_11768,N_11598,N_11633);
nand U11769 (N_11769,N_11707,N_11609);
and U11770 (N_11770,N_11725,N_11570);
or U11771 (N_11771,N_11562,N_11653);
or U11772 (N_11772,N_11603,N_11610);
and U11773 (N_11773,N_11500,N_11558);
xor U11774 (N_11774,N_11576,N_11632);
or U11775 (N_11775,N_11506,N_11712);
nor U11776 (N_11776,N_11700,N_11703);
and U11777 (N_11777,N_11734,N_11659);
nand U11778 (N_11778,N_11551,N_11711);
or U11779 (N_11779,N_11618,N_11702);
and U11780 (N_11780,N_11665,N_11568);
xnor U11781 (N_11781,N_11642,N_11567);
or U11782 (N_11782,N_11539,N_11621);
nand U11783 (N_11783,N_11640,N_11529);
or U11784 (N_11784,N_11522,N_11729);
and U11785 (N_11785,N_11571,N_11597);
nor U11786 (N_11786,N_11726,N_11616);
or U11787 (N_11787,N_11613,N_11696);
or U11788 (N_11788,N_11518,N_11550);
and U11789 (N_11789,N_11559,N_11583);
nand U11790 (N_11790,N_11681,N_11588);
nand U11791 (N_11791,N_11606,N_11575);
nand U11792 (N_11792,N_11666,N_11629);
or U11793 (N_11793,N_11652,N_11552);
nor U11794 (N_11794,N_11505,N_11645);
nor U11795 (N_11795,N_11515,N_11692);
or U11796 (N_11796,N_11599,N_11667);
nor U11797 (N_11797,N_11582,N_11595);
nor U11798 (N_11798,N_11533,N_11679);
nor U11799 (N_11799,N_11536,N_11651);
nand U11800 (N_11800,N_11676,N_11573);
and U11801 (N_11801,N_11628,N_11678);
and U11802 (N_11802,N_11743,N_11747);
or U11803 (N_11803,N_11622,N_11523);
nand U11804 (N_11804,N_11706,N_11675);
and U11805 (N_11805,N_11671,N_11569);
nand U11806 (N_11806,N_11578,N_11542);
xor U11807 (N_11807,N_11580,N_11641);
nor U11808 (N_11808,N_11722,N_11643);
or U11809 (N_11809,N_11620,N_11636);
xnor U11810 (N_11810,N_11661,N_11626);
nor U11811 (N_11811,N_11528,N_11555);
or U11812 (N_11812,N_11574,N_11596);
nand U11813 (N_11813,N_11548,N_11634);
and U11814 (N_11814,N_11623,N_11524);
and U11815 (N_11815,N_11727,N_11561);
and U11816 (N_11816,N_11501,N_11644);
xnor U11817 (N_11817,N_11602,N_11662);
and U11818 (N_11818,N_11708,N_11516);
xnor U11819 (N_11819,N_11650,N_11615);
nand U11820 (N_11820,N_11547,N_11686);
nand U11821 (N_11821,N_11673,N_11565);
or U11822 (N_11822,N_11740,N_11607);
nor U11823 (N_11823,N_11739,N_11731);
xor U11824 (N_11824,N_11509,N_11737);
nand U11825 (N_11825,N_11625,N_11532);
and U11826 (N_11826,N_11677,N_11717);
or U11827 (N_11827,N_11732,N_11535);
xnor U11828 (N_11828,N_11587,N_11735);
xor U11829 (N_11829,N_11638,N_11698);
xnor U11830 (N_11830,N_11639,N_11512);
and U11831 (N_11831,N_11543,N_11723);
nor U11832 (N_11832,N_11728,N_11687);
xnor U11833 (N_11833,N_11713,N_11637);
or U11834 (N_11834,N_11564,N_11647);
or U11835 (N_11835,N_11579,N_11537);
or U11836 (N_11836,N_11545,N_11557);
nor U11837 (N_11837,N_11680,N_11507);
or U11838 (N_11838,N_11738,N_11589);
nand U11839 (N_11839,N_11590,N_11742);
and U11840 (N_11840,N_11631,N_11572);
xnor U11841 (N_11841,N_11601,N_11699);
nand U11842 (N_11842,N_11660,N_11513);
xnor U11843 (N_11843,N_11664,N_11733);
nor U11844 (N_11844,N_11655,N_11525);
xor U11845 (N_11845,N_11534,N_11649);
xor U11846 (N_11846,N_11709,N_11682);
or U11847 (N_11847,N_11730,N_11749);
xnor U11848 (N_11848,N_11627,N_11657);
nor U11849 (N_11849,N_11669,N_11648);
nand U11850 (N_11850,N_11581,N_11566);
nor U11851 (N_11851,N_11748,N_11617);
or U11852 (N_11852,N_11521,N_11514);
nand U11853 (N_11853,N_11663,N_11697);
xor U11854 (N_11854,N_11619,N_11591);
or U11855 (N_11855,N_11721,N_11585);
xnor U11856 (N_11856,N_11604,N_11554);
xnor U11857 (N_11857,N_11724,N_11541);
or U11858 (N_11858,N_11510,N_11674);
or U11859 (N_11859,N_11538,N_11690);
or U11860 (N_11860,N_11593,N_11526);
nor U11861 (N_11861,N_11672,N_11688);
and U11862 (N_11862,N_11630,N_11701);
or U11863 (N_11863,N_11693,N_11531);
nand U11864 (N_11864,N_11718,N_11720);
or U11865 (N_11865,N_11560,N_11694);
or U11866 (N_11866,N_11556,N_11546);
nor U11867 (N_11867,N_11710,N_11646);
nor U11868 (N_11868,N_11670,N_11624);
and U11869 (N_11869,N_11563,N_11502);
and U11870 (N_11870,N_11744,N_11530);
nor U11871 (N_11871,N_11745,N_11592);
or U11872 (N_11872,N_11684,N_11586);
nand U11873 (N_11873,N_11511,N_11594);
nor U11874 (N_11874,N_11741,N_11654);
nand U11875 (N_11875,N_11686,N_11680);
xnor U11876 (N_11876,N_11548,N_11577);
and U11877 (N_11877,N_11578,N_11721);
and U11878 (N_11878,N_11641,N_11748);
nor U11879 (N_11879,N_11700,N_11533);
xnor U11880 (N_11880,N_11559,N_11544);
nor U11881 (N_11881,N_11677,N_11614);
and U11882 (N_11882,N_11593,N_11592);
or U11883 (N_11883,N_11649,N_11603);
xor U11884 (N_11884,N_11658,N_11736);
nand U11885 (N_11885,N_11555,N_11722);
and U11886 (N_11886,N_11542,N_11734);
or U11887 (N_11887,N_11630,N_11749);
xnor U11888 (N_11888,N_11507,N_11610);
or U11889 (N_11889,N_11700,N_11660);
nand U11890 (N_11890,N_11555,N_11519);
or U11891 (N_11891,N_11536,N_11643);
nand U11892 (N_11892,N_11580,N_11696);
and U11893 (N_11893,N_11552,N_11678);
and U11894 (N_11894,N_11641,N_11695);
nand U11895 (N_11895,N_11663,N_11737);
xor U11896 (N_11896,N_11555,N_11706);
and U11897 (N_11897,N_11523,N_11672);
xor U11898 (N_11898,N_11505,N_11583);
or U11899 (N_11899,N_11550,N_11557);
xnor U11900 (N_11900,N_11565,N_11577);
or U11901 (N_11901,N_11646,N_11749);
xor U11902 (N_11902,N_11549,N_11507);
and U11903 (N_11903,N_11630,N_11664);
xnor U11904 (N_11904,N_11589,N_11586);
or U11905 (N_11905,N_11639,N_11656);
or U11906 (N_11906,N_11680,N_11604);
nand U11907 (N_11907,N_11588,N_11557);
or U11908 (N_11908,N_11576,N_11562);
nand U11909 (N_11909,N_11639,N_11694);
xnor U11910 (N_11910,N_11548,N_11534);
or U11911 (N_11911,N_11644,N_11575);
and U11912 (N_11912,N_11730,N_11677);
nor U11913 (N_11913,N_11716,N_11583);
nand U11914 (N_11914,N_11741,N_11692);
nand U11915 (N_11915,N_11591,N_11654);
nor U11916 (N_11916,N_11660,N_11732);
and U11917 (N_11917,N_11562,N_11717);
or U11918 (N_11918,N_11583,N_11612);
nand U11919 (N_11919,N_11682,N_11668);
nand U11920 (N_11920,N_11614,N_11686);
nand U11921 (N_11921,N_11530,N_11586);
and U11922 (N_11922,N_11587,N_11714);
nor U11923 (N_11923,N_11678,N_11509);
or U11924 (N_11924,N_11630,N_11730);
or U11925 (N_11925,N_11521,N_11528);
nand U11926 (N_11926,N_11528,N_11613);
xnor U11927 (N_11927,N_11717,N_11542);
nand U11928 (N_11928,N_11546,N_11506);
xnor U11929 (N_11929,N_11660,N_11531);
and U11930 (N_11930,N_11548,N_11617);
xnor U11931 (N_11931,N_11502,N_11653);
xor U11932 (N_11932,N_11724,N_11523);
and U11933 (N_11933,N_11643,N_11552);
nand U11934 (N_11934,N_11637,N_11516);
and U11935 (N_11935,N_11747,N_11506);
and U11936 (N_11936,N_11633,N_11630);
and U11937 (N_11937,N_11534,N_11706);
nand U11938 (N_11938,N_11542,N_11648);
nand U11939 (N_11939,N_11712,N_11571);
nor U11940 (N_11940,N_11666,N_11657);
nor U11941 (N_11941,N_11548,N_11552);
nor U11942 (N_11942,N_11500,N_11657);
nand U11943 (N_11943,N_11705,N_11692);
nand U11944 (N_11944,N_11581,N_11685);
or U11945 (N_11945,N_11674,N_11683);
xnor U11946 (N_11946,N_11539,N_11590);
or U11947 (N_11947,N_11551,N_11667);
and U11948 (N_11948,N_11616,N_11600);
or U11949 (N_11949,N_11608,N_11622);
nand U11950 (N_11950,N_11680,N_11662);
and U11951 (N_11951,N_11556,N_11649);
nand U11952 (N_11952,N_11559,N_11659);
xor U11953 (N_11953,N_11596,N_11624);
nand U11954 (N_11954,N_11640,N_11685);
or U11955 (N_11955,N_11715,N_11580);
or U11956 (N_11956,N_11619,N_11724);
xnor U11957 (N_11957,N_11576,N_11699);
nand U11958 (N_11958,N_11516,N_11503);
nand U11959 (N_11959,N_11726,N_11591);
xor U11960 (N_11960,N_11699,N_11646);
nand U11961 (N_11961,N_11679,N_11507);
xor U11962 (N_11962,N_11673,N_11663);
and U11963 (N_11963,N_11661,N_11599);
nand U11964 (N_11964,N_11706,N_11617);
nor U11965 (N_11965,N_11669,N_11746);
xor U11966 (N_11966,N_11641,N_11722);
nand U11967 (N_11967,N_11584,N_11538);
and U11968 (N_11968,N_11558,N_11620);
and U11969 (N_11969,N_11594,N_11619);
nand U11970 (N_11970,N_11709,N_11566);
nand U11971 (N_11971,N_11552,N_11688);
xor U11972 (N_11972,N_11550,N_11549);
nor U11973 (N_11973,N_11684,N_11529);
nand U11974 (N_11974,N_11628,N_11644);
and U11975 (N_11975,N_11678,N_11555);
xor U11976 (N_11976,N_11502,N_11695);
or U11977 (N_11977,N_11509,N_11716);
and U11978 (N_11978,N_11640,N_11545);
and U11979 (N_11979,N_11605,N_11563);
xnor U11980 (N_11980,N_11617,N_11648);
and U11981 (N_11981,N_11623,N_11600);
and U11982 (N_11982,N_11680,N_11719);
nor U11983 (N_11983,N_11674,N_11591);
or U11984 (N_11984,N_11688,N_11630);
and U11985 (N_11985,N_11663,N_11670);
and U11986 (N_11986,N_11696,N_11748);
nor U11987 (N_11987,N_11743,N_11541);
nand U11988 (N_11988,N_11542,N_11624);
nor U11989 (N_11989,N_11675,N_11538);
xnor U11990 (N_11990,N_11700,N_11626);
nand U11991 (N_11991,N_11571,N_11619);
xor U11992 (N_11992,N_11565,N_11538);
nor U11993 (N_11993,N_11741,N_11530);
and U11994 (N_11994,N_11594,N_11697);
and U11995 (N_11995,N_11646,N_11738);
xnor U11996 (N_11996,N_11567,N_11653);
xor U11997 (N_11997,N_11711,N_11725);
and U11998 (N_11998,N_11705,N_11577);
and U11999 (N_11999,N_11735,N_11741);
nand U12000 (N_12000,N_11798,N_11751);
nor U12001 (N_12001,N_11869,N_11871);
and U12002 (N_12002,N_11912,N_11758);
xor U12003 (N_12003,N_11952,N_11995);
nor U12004 (N_12004,N_11951,N_11884);
and U12005 (N_12005,N_11803,N_11794);
or U12006 (N_12006,N_11859,N_11934);
nor U12007 (N_12007,N_11970,N_11811);
or U12008 (N_12008,N_11854,N_11950);
xnor U12009 (N_12009,N_11752,N_11855);
or U12010 (N_12010,N_11770,N_11864);
nor U12011 (N_12011,N_11755,N_11833);
and U12012 (N_12012,N_11832,N_11886);
or U12013 (N_12013,N_11947,N_11954);
or U12014 (N_12014,N_11787,N_11987);
and U12015 (N_12015,N_11763,N_11984);
nand U12016 (N_12016,N_11812,N_11856);
nand U12017 (N_12017,N_11932,N_11780);
nand U12018 (N_12018,N_11822,N_11773);
nand U12019 (N_12019,N_11893,N_11767);
nor U12020 (N_12020,N_11988,N_11777);
nor U12021 (N_12021,N_11820,N_11776);
xor U12022 (N_12022,N_11843,N_11894);
nor U12023 (N_12023,N_11924,N_11940);
and U12024 (N_12024,N_11759,N_11983);
xnor U12025 (N_12025,N_11809,N_11910);
or U12026 (N_12026,N_11975,N_11909);
nor U12027 (N_12027,N_11817,N_11901);
or U12028 (N_12028,N_11906,N_11830);
nor U12029 (N_12029,N_11921,N_11764);
xnor U12030 (N_12030,N_11927,N_11985);
or U12031 (N_12031,N_11892,N_11899);
or U12032 (N_12032,N_11997,N_11781);
and U12033 (N_12033,N_11907,N_11753);
nand U12034 (N_12034,N_11862,N_11880);
nor U12035 (N_12035,N_11806,N_11937);
nor U12036 (N_12036,N_11786,N_11800);
or U12037 (N_12037,N_11805,N_11902);
or U12038 (N_12038,N_11966,N_11925);
xor U12039 (N_12039,N_11978,N_11877);
or U12040 (N_12040,N_11979,N_11846);
nor U12041 (N_12041,N_11953,N_11908);
and U12042 (N_12042,N_11897,N_11818);
nand U12043 (N_12043,N_11814,N_11891);
nor U12044 (N_12044,N_11918,N_11771);
xnor U12045 (N_12045,N_11876,N_11959);
and U12046 (N_12046,N_11993,N_11990);
nand U12047 (N_12047,N_11841,N_11955);
nor U12048 (N_12048,N_11939,N_11831);
and U12049 (N_12049,N_11792,N_11836);
xnor U12050 (N_12050,N_11903,N_11980);
and U12051 (N_12051,N_11956,N_11797);
or U12052 (N_12052,N_11839,N_11941);
nor U12053 (N_12053,N_11900,N_11948);
or U12054 (N_12054,N_11935,N_11772);
nand U12055 (N_12055,N_11972,N_11850);
or U12056 (N_12056,N_11863,N_11957);
and U12057 (N_12057,N_11982,N_11890);
nor U12058 (N_12058,N_11881,N_11791);
and U12059 (N_12059,N_11840,N_11765);
xor U12060 (N_12060,N_11878,N_11821);
nand U12061 (N_12061,N_11824,N_11938);
xnor U12062 (N_12062,N_11834,N_11922);
xor U12063 (N_12063,N_11969,N_11904);
nand U12064 (N_12064,N_11981,N_11775);
nand U12065 (N_12065,N_11998,N_11828);
nor U12066 (N_12066,N_11783,N_11882);
xnor U12067 (N_12067,N_11913,N_11852);
and U12068 (N_12068,N_11860,N_11845);
nand U12069 (N_12069,N_11802,N_11813);
xnor U12070 (N_12070,N_11804,N_11867);
or U12071 (N_12071,N_11889,N_11919);
xor U12072 (N_12072,N_11847,N_11936);
and U12073 (N_12073,N_11848,N_11961);
nor U12074 (N_12074,N_11943,N_11819);
and U12075 (N_12075,N_11887,N_11866);
and U12076 (N_12076,N_11992,N_11960);
and U12077 (N_12077,N_11815,N_11928);
and U12078 (N_12078,N_11874,N_11778);
or U12079 (N_12079,N_11849,N_11789);
xor U12080 (N_12080,N_11949,N_11754);
or U12081 (N_12081,N_11795,N_11760);
nand U12082 (N_12082,N_11930,N_11996);
and U12083 (N_12083,N_11926,N_11766);
nand U12084 (N_12084,N_11933,N_11994);
or U12085 (N_12085,N_11929,N_11790);
nor U12086 (N_12086,N_11973,N_11838);
xnor U12087 (N_12087,N_11875,N_11762);
and U12088 (N_12088,N_11757,N_11808);
and U12089 (N_12089,N_11788,N_11816);
nor U12090 (N_12090,N_11837,N_11911);
nor U12091 (N_12091,N_11785,N_11826);
xor U12092 (N_12092,N_11879,N_11750);
xor U12093 (N_12093,N_11774,N_11905);
xor U12094 (N_12094,N_11835,N_11977);
xnor U12095 (N_12095,N_11945,N_11931);
nor U12096 (N_12096,N_11883,N_11768);
or U12097 (N_12097,N_11844,N_11923);
xnor U12098 (N_12098,N_11915,N_11976);
or U12099 (N_12099,N_11917,N_11944);
nor U12100 (N_12100,N_11963,N_11916);
xnor U12101 (N_12101,N_11756,N_11807);
nor U12102 (N_12102,N_11896,N_11971);
or U12103 (N_12103,N_11872,N_11962);
nor U12104 (N_12104,N_11853,N_11991);
nor U12105 (N_12105,N_11793,N_11868);
and U12106 (N_12106,N_11827,N_11858);
nand U12107 (N_12107,N_11810,N_11865);
nor U12108 (N_12108,N_11801,N_11974);
nand U12109 (N_12109,N_11895,N_11825);
and U12110 (N_12110,N_11769,N_11842);
xor U12111 (N_12111,N_11779,N_11999);
or U12112 (N_12112,N_11888,N_11958);
xor U12113 (N_12113,N_11942,N_11761);
or U12114 (N_12114,N_11898,N_11799);
nand U12115 (N_12115,N_11986,N_11823);
and U12116 (N_12116,N_11782,N_11920);
nor U12117 (N_12117,N_11796,N_11946);
nor U12118 (N_12118,N_11914,N_11989);
or U12119 (N_12119,N_11964,N_11857);
nand U12120 (N_12120,N_11870,N_11861);
nand U12121 (N_12121,N_11968,N_11885);
xor U12122 (N_12122,N_11967,N_11829);
xor U12123 (N_12123,N_11851,N_11873);
nor U12124 (N_12124,N_11965,N_11784);
xor U12125 (N_12125,N_11889,N_11922);
nand U12126 (N_12126,N_11877,N_11898);
xnor U12127 (N_12127,N_11917,N_11938);
xnor U12128 (N_12128,N_11924,N_11767);
xor U12129 (N_12129,N_11791,N_11807);
nand U12130 (N_12130,N_11768,N_11913);
nor U12131 (N_12131,N_11755,N_11905);
nor U12132 (N_12132,N_11977,N_11992);
nand U12133 (N_12133,N_11956,N_11839);
xnor U12134 (N_12134,N_11966,N_11855);
xnor U12135 (N_12135,N_11788,N_11944);
or U12136 (N_12136,N_11959,N_11877);
nor U12137 (N_12137,N_11943,N_11854);
nand U12138 (N_12138,N_11843,N_11945);
nor U12139 (N_12139,N_11862,N_11761);
nand U12140 (N_12140,N_11867,N_11963);
xor U12141 (N_12141,N_11943,N_11931);
nand U12142 (N_12142,N_11792,N_11851);
nor U12143 (N_12143,N_11840,N_11773);
or U12144 (N_12144,N_11793,N_11785);
or U12145 (N_12145,N_11903,N_11887);
or U12146 (N_12146,N_11983,N_11919);
nor U12147 (N_12147,N_11834,N_11806);
nor U12148 (N_12148,N_11756,N_11903);
or U12149 (N_12149,N_11869,N_11998);
or U12150 (N_12150,N_11982,N_11855);
or U12151 (N_12151,N_11812,N_11860);
xor U12152 (N_12152,N_11799,N_11763);
and U12153 (N_12153,N_11979,N_11965);
nand U12154 (N_12154,N_11790,N_11816);
or U12155 (N_12155,N_11964,N_11848);
xnor U12156 (N_12156,N_11785,N_11767);
and U12157 (N_12157,N_11829,N_11923);
and U12158 (N_12158,N_11991,N_11832);
nand U12159 (N_12159,N_11861,N_11855);
nor U12160 (N_12160,N_11985,N_11899);
and U12161 (N_12161,N_11954,N_11904);
and U12162 (N_12162,N_11818,N_11947);
xor U12163 (N_12163,N_11753,N_11853);
xor U12164 (N_12164,N_11918,N_11755);
nand U12165 (N_12165,N_11903,N_11820);
or U12166 (N_12166,N_11908,N_11883);
nor U12167 (N_12167,N_11922,N_11974);
xor U12168 (N_12168,N_11948,N_11856);
nor U12169 (N_12169,N_11914,N_11915);
or U12170 (N_12170,N_11918,N_11842);
nor U12171 (N_12171,N_11838,N_11899);
and U12172 (N_12172,N_11907,N_11771);
nor U12173 (N_12173,N_11895,N_11845);
xor U12174 (N_12174,N_11772,N_11811);
nand U12175 (N_12175,N_11756,N_11765);
and U12176 (N_12176,N_11757,N_11821);
and U12177 (N_12177,N_11838,N_11792);
xnor U12178 (N_12178,N_11790,N_11851);
nor U12179 (N_12179,N_11948,N_11848);
xor U12180 (N_12180,N_11850,N_11976);
nand U12181 (N_12181,N_11934,N_11827);
or U12182 (N_12182,N_11984,N_11978);
nor U12183 (N_12183,N_11899,N_11960);
and U12184 (N_12184,N_11839,N_11930);
nand U12185 (N_12185,N_11866,N_11973);
and U12186 (N_12186,N_11886,N_11808);
and U12187 (N_12187,N_11851,N_11993);
nand U12188 (N_12188,N_11883,N_11774);
xor U12189 (N_12189,N_11786,N_11833);
nand U12190 (N_12190,N_11810,N_11753);
nor U12191 (N_12191,N_11856,N_11750);
xnor U12192 (N_12192,N_11956,N_11891);
nor U12193 (N_12193,N_11991,N_11779);
and U12194 (N_12194,N_11867,N_11970);
and U12195 (N_12195,N_11840,N_11825);
xnor U12196 (N_12196,N_11880,N_11945);
nand U12197 (N_12197,N_11995,N_11756);
nor U12198 (N_12198,N_11970,N_11856);
nor U12199 (N_12199,N_11925,N_11913);
and U12200 (N_12200,N_11978,N_11824);
and U12201 (N_12201,N_11795,N_11891);
nand U12202 (N_12202,N_11782,N_11916);
nand U12203 (N_12203,N_11907,N_11899);
or U12204 (N_12204,N_11913,N_11797);
nand U12205 (N_12205,N_11891,N_11920);
and U12206 (N_12206,N_11902,N_11792);
xor U12207 (N_12207,N_11833,N_11821);
or U12208 (N_12208,N_11850,N_11819);
nand U12209 (N_12209,N_11889,N_11936);
or U12210 (N_12210,N_11999,N_11858);
and U12211 (N_12211,N_11772,N_11948);
xnor U12212 (N_12212,N_11926,N_11902);
and U12213 (N_12213,N_11876,N_11764);
and U12214 (N_12214,N_11797,N_11927);
and U12215 (N_12215,N_11766,N_11896);
or U12216 (N_12216,N_11795,N_11762);
nor U12217 (N_12217,N_11808,N_11811);
and U12218 (N_12218,N_11956,N_11998);
and U12219 (N_12219,N_11853,N_11875);
and U12220 (N_12220,N_11766,N_11781);
xnor U12221 (N_12221,N_11788,N_11810);
or U12222 (N_12222,N_11854,N_11926);
and U12223 (N_12223,N_11990,N_11815);
nor U12224 (N_12224,N_11886,N_11830);
and U12225 (N_12225,N_11819,N_11890);
nand U12226 (N_12226,N_11984,N_11982);
nand U12227 (N_12227,N_11808,N_11951);
xnor U12228 (N_12228,N_11975,N_11871);
and U12229 (N_12229,N_11962,N_11983);
or U12230 (N_12230,N_11849,N_11836);
xnor U12231 (N_12231,N_11819,N_11772);
and U12232 (N_12232,N_11950,N_11759);
nand U12233 (N_12233,N_11959,N_11919);
xnor U12234 (N_12234,N_11892,N_11854);
or U12235 (N_12235,N_11954,N_11977);
nand U12236 (N_12236,N_11795,N_11850);
and U12237 (N_12237,N_11954,N_11806);
and U12238 (N_12238,N_11870,N_11820);
nor U12239 (N_12239,N_11794,N_11989);
and U12240 (N_12240,N_11855,N_11961);
and U12241 (N_12241,N_11846,N_11931);
and U12242 (N_12242,N_11771,N_11868);
xor U12243 (N_12243,N_11804,N_11764);
nor U12244 (N_12244,N_11775,N_11897);
nor U12245 (N_12245,N_11762,N_11781);
xor U12246 (N_12246,N_11854,N_11993);
and U12247 (N_12247,N_11906,N_11859);
nor U12248 (N_12248,N_11892,N_11855);
nand U12249 (N_12249,N_11874,N_11889);
nor U12250 (N_12250,N_12027,N_12109);
xor U12251 (N_12251,N_12208,N_12074);
and U12252 (N_12252,N_12091,N_12225);
and U12253 (N_12253,N_12167,N_12116);
nor U12254 (N_12254,N_12089,N_12187);
and U12255 (N_12255,N_12186,N_12001);
and U12256 (N_12256,N_12192,N_12141);
or U12257 (N_12257,N_12016,N_12182);
nand U12258 (N_12258,N_12242,N_12088);
nor U12259 (N_12259,N_12097,N_12220);
and U12260 (N_12260,N_12232,N_12000);
or U12261 (N_12261,N_12139,N_12176);
or U12262 (N_12262,N_12107,N_12226);
or U12263 (N_12263,N_12179,N_12050);
and U12264 (N_12264,N_12193,N_12124);
or U12265 (N_12265,N_12244,N_12163);
nand U12266 (N_12266,N_12130,N_12235);
xor U12267 (N_12267,N_12102,N_12047);
and U12268 (N_12268,N_12128,N_12070);
or U12269 (N_12269,N_12165,N_12080);
and U12270 (N_12270,N_12065,N_12009);
nor U12271 (N_12271,N_12048,N_12157);
and U12272 (N_12272,N_12202,N_12207);
and U12273 (N_12273,N_12022,N_12061);
or U12274 (N_12274,N_12029,N_12223);
or U12275 (N_12275,N_12201,N_12227);
and U12276 (N_12276,N_12203,N_12085);
xnor U12277 (N_12277,N_12018,N_12087);
or U12278 (N_12278,N_12121,N_12114);
and U12279 (N_12279,N_12147,N_12049);
and U12280 (N_12280,N_12233,N_12161);
nand U12281 (N_12281,N_12012,N_12038);
or U12282 (N_12282,N_12180,N_12237);
and U12283 (N_12283,N_12246,N_12150);
or U12284 (N_12284,N_12210,N_12031);
and U12285 (N_12285,N_12055,N_12026);
and U12286 (N_12286,N_12195,N_12046);
nor U12287 (N_12287,N_12007,N_12052);
xor U12288 (N_12288,N_12185,N_12005);
or U12289 (N_12289,N_12083,N_12229);
nor U12290 (N_12290,N_12146,N_12216);
xor U12291 (N_12291,N_12213,N_12148);
and U12292 (N_12292,N_12138,N_12191);
nor U12293 (N_12293,N_12175,N_12212);
xor U12294 (N_12294,N_12108,N_12006);
and U12295 (N_12295,N_12096,N_12156);
or U12296 (N_12296,N_12234,N_12002);
nand U12297 (N_12297,N_12069,N_12020);
nand U12298 (N_12298,N_12200,N_12219);
or U12299 (N_12299,N_12172,N_12155);
xor U12300 (N_12300,N_12238,N_12249);
and U12301 (N_12301,N_12145,N_12053);
nand U12302 (N_12302,N_12159,N_12215);
xnor U12303 (N_12303,N_12066,N_12181);
nor U12304 (N_12304,N_12170,N_12057);
nand U12305 (N_12305,N_12032,N_12098);
and U12306 (N_12306,N_12158,N_12160);
nand U12307 (N_12307,N_12072,N_12077);
xor U12308 (N_12308,N_12034,N_12094);
xor U12309 (N_12309,N_12151,N_12221);
and U12310 (N_12310,N_12039,N_12214);
xor U12311 (N_12311,N_12103,N_12051);
xor U12312 (N_12312,N_12131,N_12117);
nand U12313 (N_12313,N_12198,N_12013);
xnor U12314 (N_12314,N_12037,N_12075);
xor U12315 (N_12315,N_12059,N_12188);
or U12316 (N_12316,N_12073,N_12078);
and U12317 (N_12317,N_12174,N_12101);
nor U12318 (N_12318,N_12149,N_12190);
and U12319 (N_12319,N_12123,N_12166);
xor U12320 (N_12320,N_12122,N_12060);
xnor U12321 (N_12321,N_12062,N_12135);
or U12322 (N_12322,N_12171,N_12177);
nor U12323 (N_12323,N_12133,N_12230);
nand U12324 (N_12324,N_12241,N_12017);
xnor U12325 (N_12325,N_12025,N_12239);
and U12326 (N_12326,N_12127,N_12144);
and U12327 (N_12327,N_12086,N_12248);
nand U12328 (N_12328,N_12132,N_12054);
nor U12329 (N_12329,N_12040,N_12152);
or U12330 (N_12330,N_12110,N_12119);
or U12331 (N_12331,N_12236,N_12134);
and U12332 (N_12332,N_12042,N_12224);
nor U12333 (N_12333,N_12045,N_12196);
nor U12334 (N_12334,N_12010,N_12036);
xnor U12335 (N_12335,N_12169,N_12071);
nor U12336 (N_12336,N_12205,N_12021);
xnor U12337 (N_12337,N_12211,N_12243);
and U12338 (N_12338,N_12093,N_12184);
xor U12339 (N_12339,N_12014,N_12104);
nand U12340 (N_12340,N_12126,N_12106);
nor U12341 (N_12341,N_12199,N_12011);
xor U12342 (N_12342,N_12063,N_12068);
nand U12343 (N_12343,N_12090,N_12217);
nor U12344 (N_12344,N_12115,N_12153);
or U12345 (N_12345,N_12081,N_12245);
nor U12346 (N_12346,N_12113,N_12173);
nand U12347 (N_12347,N_12008,N_12092);
xor U12348 (N_12348,N_12168,N_12218);
and U12349 (N_12349,N_12143,N_12003);
or U12350 (N_12350,N_12222,N_12056);
nor U12351 (N_12351,N_12118,N_12247);
xor U12352 (N_12352,N_12064,N_12120);
xnor U12353 (N_12353,N_12076,N_12240);
nand U12354 (N_12354,N_12183,N_12082);
xor U12355 (N_12355,N_12228,N_12004);
nor U12356 (N_12356,N_12154,N_12197);
nor U12357 (N_12357,N_12043,N_12084);
or U12358 (N_12358,N_12044,N_12111);
and U12359 (N_12359,N_12079,N_12125);
xnor U12360 (N_12360,N_12058,N_12015);
xnor U12361 (N_12361,N_12105,N_12129);
and U12362 (N_12362,N_12140,N_12033);
or U12363 (N_12363,N_12194,N_12178);
or U12364 (N_12364,N_12019,N_12136);
or U12365 (N_12365,N_12231,N_12095);
or U12366 (N_12366,N_12112,N_12023);
and U12367 (N_12367,N_12041,N_12162);
xnor U12368 (N_12368,N_12028,N_12164);
and U12369 (N_12369,N_12189,N_12030);
xnor U12370 (N_12370,N_12024,N_12142);
nand U12371 (N_12371,N_12206,N_12137);
nand U12372 (N_12372,N_12035,N_12209);
nand U12373 (N_12373,N_12204,N_12099);
xnor U12374 (N_12374,N_12067,N_12100);
and U12375 (N_12375,N_12176,N_12126);
and U12376 (N_12376,N_12040,N_12013);
nor U12377 (N_12377,N_12022,N_12097);
xnor U12378 (N_12378,N_12035,N_12215);
nand U12379 (N_12379,N_12069,N_12081);
nor U12380 (N_12380,N_12084,N_12041);
nand U12381 (N_12381,N_12099,N_12037);
xnor U12382 (N_12382,N_12201,N_12015);
xnor U12383 (N_12383,N_12145,N_12222);
nand U12384 (N_12384,N_12148,N_12089);
nand U12385 (N_12385,N_12087,N_12111);
nand U12386 (N_12386,N_12132,N_12236);
or U12387 (N_12387,N_12079,N_12168);
or U12388 (N_12388,N_12177,N_12016);
and U12389 (N_12389,N_12021,N_12072);
and U12390 (N_12390,N_12163,N_12065);
and U12391 (N_12391,N_12248,N_12168);
or U12392 (N_12392,N_12001,N_12081);
or U12393 (N_12393,N_12168,N_12214);
nor U12394 (N_12394,N_12125,N_12188);
nor U12395 (N_12395,N_12169,N_12127);
nand U12396 (N_12396,N_12057,N_12174);
and U12397 (N_12397,N_12156,N_12019);
or U12398 (N_12398,N_12123,N_12026);
nand U12399 (N_12399,N_12115,N_12151);
or U12400 (N_12400,N_12018,N_12131);
nand U12401 (N_12401,N_12054,N_12105);
xnor U12402 (N_12402,N_12210,N_12052);
nor U12403 (N_12403,N_12115,N_12227);
nand U12404 (N_12404,N_12165,N_12233);
xnor U12405 (N_12405,N_12229,N_12113);
nor U12406 (N_12406,N_12112,N_12204);
or U12407 (N_12407,N_12235,N_12049);
xor U12408 (N_12408,N_12242,N_12126);
nand U12409 (N_12409,N_12201,N_12217);
and U12410 (N_12410,N_12171,N_12121);
nand U12411 (N_12411,N_12082,N_12087);
nand U12412 (N_12412,N_12244,N_12215);
nand U12413 (N_12413,N_12018,N_12215);
xnor U12414 (N_12414,N_12014,N_12023);
or U12415 (N_12415,N_12241,N_12194);
or U12416 (N_12416,N_12141,N_12044);
and U12417 (N_12417,N_12126,N_12172);
or U12418 (N_12418,N_12204,N_12096);
xor U12419 (N_12419,N_12163,N_12102);
and U12420 (N_12420,N_12212,N_12039);
nand U12421 (N_12421,N_12231,N_12115);
nor U12422 (N_12422,N_12060,N_12244);
or U12423 (N_12423,N_12050,N_12248);
or U12424 (N_12424,N_12215,N_12249);
and U12425 (N_12425,N_12117,N_12080);
nand U12426 (N_12426,N_12055,N_12079);
xor U12427 (N_12427,N_12089,N_12017);
or U12428 (N_12428,N_12234,N_12166);
nand U12429 (N_12429,N_12230,N_12209);
nand U12430 (N_12430,N_12171,N_12207);
or U12431 (N_12431,N_12024,N_12242);
nand U12432 (N_12432,N_12107,N_12133);
nand U12433 (N_12433,N_12213,N_12205);
and U12434 (N_12434,N_12049,N_12106);
nor U12435 (N_12435,N_12161,N_12148);
nor U12436 (N_12436,N_12129,N_12137);
and U12437 (N_12437,N_12151,N_12043);
and U12438 (N_12438,N_12083,N_12167);
xnor U12439 (N_12439,N_12192,N_12122);
and U12440 (N_12440,N_12000,N_12231);
and U12441 (N_12441,N_12045,N_12125);
nand U12442 (N_12442,N_12040,N_12011);
xnor U12443 (N_12443,N_12101,N_12062);
nor U12444 (N_12444,N_12054,N_12079);
or U12445 (N_12445,N_12227,N_12049);
or U12446 (N_12446,N_12055,N_12193);
xor U12447 (N_12447,N_12222,N_12158);
nor U12448 (N_12448,N_12243,N_12033);
nor U12449 (N_12449,N_12216,N_12023);
nand U12450 (N_12450,N_12214,N_12128);
nand U12451 (N_12451,N_12179,N_12047);
nor U12452 (N_12452,N_12091,N_12241);
nor U12453 (N_12453,N_12249,N_12043);
and U12454 (N_12454,N_12062,N_12063);
or U12455 (N_12455,N_12025,N_12012);
or U12456 (N_12456,N_12211,N_12028);
xnor U12457 (N_12457,N_12005,N_12090);
xor U12458 (N_12458,N_12161,N_12220);
xnor U12459 (N_12459,N_12140,N_12131);
xor U12460 (N_12460,N_12205,N_12023);
nor U12461 (N_12461,N_12065,N_12120);
xor U12462 (N_12462,N_12058,N_12087);
nor U12463 (N_12463,N_12192,N_12018);
or U12464 (N_12464,N_12240,N_12245);
or U12465 (N_12465,N_12101,N_12072);
nand U12466 (N_12466,N_12060,N_12173);
xor U12467 (N_12467,N_12226,N_12191);
nand U12468 (N_12468,N_12102,N_12037);
xor U12469 (N_12469,N_12082,N_12076);
or U12470 (N_12470,N_12133,N_12220);
nand U12471 (N_12471,N_12117,N_12213);
nand U12472 (N_12472,N_12003,N_12022);
nand U12473 (N_12473,N_12188,N_12082);
nand U12474 (N_12474,N_12080,N_12194);
nand U12475 (N_12475,N_12025,N_12110);
nand U12476 (N_12476,N_12110,N_12216);
and U12477 (N_12477,N_12105,N_12133);
nand U12478 (N_12478,N_12109,N_12242);
xor U12479 (N_12479,N_12117,N_12052);
nand U12480 (N_12480,N_12064,N_12063);
and U12481 (N_12481,N_12217,N_12103);
nor U12482 (N_12482,N_12197,N_12065);
and U12483 (N_12483,N_12215,N_12126);
xor U12484 (N_12484,N_12200,N_12164);
and U12485 (N_12485,N_12067,N_12245);
and U12486 (N_12486,N_12237,N_12203);
or U12487 (N_12487,N_12212,N_12116);
xor U12488 (N_12488,N_12130,N_12124);
nor U12489 (N_12489,N_12105,N_12036);
nor U12490 (N_12490,N_12216,N_12249);
and U12491 (N_12491,N_12085,N_12069);
nor U12492 (N_12492,N_12037,N_12089);
or U12493 (N_12493,N_12192,N_12184);
and U12494 (N_12494,N_12159,N_12212);
nor U12495 (N_12495,N_12062,N_12134);
nand U12496 (N_12496,N_12112,N_12212);
xor U12497 (N_12497,N_12227,N_12008);
nor U12498 (N_12498,N_12247,N_12085);
nor U12499 (N_12499,N_12068,N_12192);
or U12500 (N_12500,N_12413,N_12332);
nand U12501 (N_12501,N_12496,N_12422);
or U12502 (N_12502,N_12337,N_12471);
xnor U12503 (N_12503,N_12437,N_12364);
nand U12504 (N_12504,N_12392,N_12490);
and U12505 (N_12505,N_12426,N_12411);
and U12506 (N_12506,N_12367,N_12481);
and U12507 (N_12507,N_12450,N_12268);
xnor U12508 (N_12508,N_12498,N_12475);
and U12509 (N_12509,N_12431,N_12476);
xnor U12510 (N_12510,N_12400,N_12321);
and U12511 (N_12511,N_12446,N_12410);
xor U12512 (N_12512,N_12483,N_12439);
nand U12513 (N_12513,N_12432,N_12380);
nand U12514 (N_12514,N_12457,N_12463);
and U12515 (N_12515,N_12438,N_12362);
and U12516 (N_12516,N_12479,N_12289);
nor U12517 (N_12517,N_12276,N_12312);
nand U12518 (N_12518,N_12478,N_12454);
nand U12519 (N_12519,N_12255,N_12453);
nand U12520 (N_12520,N_12383,N_12279);
and U12521 (N_12521,N_12421,N_12396);
and U12522 (N_12522,N_12253,N_12336);
xnor U12523 (N_12523,N_12342,N_12323);
nand U12524 (N_12524,N_12294,N_12274);
and U12525 (N_12525,N_12424,N_12464);
and U12526 (N_12526,N_12442,N_12301);
nor U12527 (N_12527,N_12252,N_12415);
nor U12528 (N_12528,N_12369,N_12462);
or U12529 (N_12529,N_12365,N_12313);
nor U12530 (N_12530,N_12254,N_12260);
xor U12531 (N_12531,N_12455,N_12472);
and U12532 (N_12532,N_12390,N_12360);
nand U12533 (N_12533,N_12314,N_12347);
xnor U12534 (N_12534,N_12309,N_12250);
or U12535 (N_12535,N_12381,N_12370);
and U12536 (N_12536,N_12290,N_12468);
nor U12537 (N_12537,N_12328,N_12441);
nand U12538 (N_12538,N_12382,N_12348);
nor U12539 (N_12539,N_12378,N_12251);
or U12540 (N_12540,N_12448,N_12277);
nand U12541 (N_12541,N_12489,N_12435);
and U12542 (N_12542,N_12401,N_12358);
xor U12543 (N_12543,N_12419,N_12458);
and U12544 (N_12544,N_12376,N_12461);
xnor U12545 (N_12545,N_12263,N_12258);
and U12546 (N_12546,N_12283,N_12331);
or U12547 (N_12547,N_12354,N_12452);
nand U12548 (N_12548,N_12257,N_12470);
nand U12549 (N_12549,N_12480,N_12357);
xor U12550 (N_12550,N_12408,N_12318);
xnor U12551 (N_12551,N_12388,N_12375);
nand U12552 (N_12552,N_12266,N_12265);
or U12553 (N_12553,N_12291,N_12394);
and U12554 (N_12554,N_12350,N_12406);
nand U12555 (N_12555,N_12412,N_12443);
and U12556 (N_12556,N_12271,N_12418);
or U12557 (N_12557,N_12273,N_12428);
and U12558 (N_12558,N_12414,N_12387);
or U12559 (N_12559,N_12272,N_12329);
or U12560 (N_12560,N_12397,N_12379);
nor U12561 (N_12561,N_12398,N_12305);
xnor U12562 (N_12562,N_12349,N_12430);
or U12563 (N_12563,N_12297,N_12356);
or U12564 (N_12564,N_12353,N_12303);
xor U12565 (N_12565,N_12493,N_12316);
nand U12566 (N_12566,N_12287,N_12307);
and U12567 (N_12567,N_12427,N_12491);
and U12568 (N_12568,N_12420,N_12447);
or U12569 (N_12569,N_12460,N_12366);
and U12570 (N_12570,N_12296,N_12386);
nor U12571 (N_12571,N_12256,N_12359);
nand U12572 (N_12572,N_12492,N_12264);
nor U12573 (N_12573,N_12324,N_12445);
nand U12574 (N_12574,N_12341,N_12485);
or U12575 (N_12575,N_12395,N_12298);
or U12576 (N_12576,N_12330,N_12488);
and U12577 (N_12577,N_12494,N_12320);
nand U12578 (N_12578,N_12327,N_12474);
nor U12579 (N_12579,N_12477,N_12299);
and U12580 (N_12580,N_12280,N_12262);
xnor U12581 (N_12581,N_12319,N_12345);
xnor U12582 (N_12582,N_12292,N_12417);
or U12583 (N_12583,N_12482,N_12304);
nand U12584 (N_12584,N_12267,N_12338);
nor U12585 (N_12585,N_12334,N_12285);
and U12586 (N_12586,N_12377,N_12434);
and U12587 (N_12587,N_12355,N_12436);
nand U12588 (N_12588,N_12429,N_12259);
or U12589 (N_12589,N_12344,N_12384);
or U12590 (N_12590,N_12315,N_12310);
and U12591 (N_12591,N_12393,N_12391);
or U12592 (N_12592,N_12282,N_12371);
xnor U12593 (N_12593,N_12293,N_12444);
and U12594 (N_12594,N_12402,N_12286);
nor U12595 (N_12595,N_12278,N_12425);
nand U12596 (N_12596,N_12407,N_12335);
or U12597 (N_12597,N_12340,N_12456);
nor U12598 (N_12598,N_12373,N_12487);
nand U12599 (N_12599,N_12311,N_12459);
xor U12600 (N_12600,N_12451,N_12449);
and U12601 (N_12601,N_12295,N_12308);
nand U12602 (N_12602,N_12306,N_12486);
and U12603 (N_12603,N_12372,N_12275);
xor U12604 (N_12604,N_12317,N_12467);
nor U12605 (N_12605,N_12404,N_12339);
xor U12606 (N_12606,N_12469,N_12440);
nand U12607 (N_12607,N_12385,N_12288);
nor U12608 (N_12608,N_12423,N_12433);
nand U12609 (N_12609,N_12261,N_12333);
nor U12610 (N_12610,N_12363,N_12405);
and U12611 (N_12611,N_12322,N_12473);
nor U12612 (N_12612,N_12300,N_12325);
xor U12613 (N_12613,N_12352,N_12343);
xnor U12614 (N_12614,N_12269,N_12399);
and U12615 (N_12615,N_12346,N_12416);
xnor U12616 (N_12616,N_12495,N_12409);
and U12617 (N_12617,N_12302,N_12361);
nand U12618 (N_12618,N_12497,N_12284);
xnor U12619 (N_12619,N_12351,N_12499);
or U12620 (N_12620,N_12403,N_12270);
or U12621 (N_12621,N_12466,N_12326);
or U12622 (N_12622,N_12374,N_12465);
xnor U12623 (N_12623,N_12389,N_12484);
xor U12624 (N_12624,N_12368,N_12281);
or U12625 (N_12625,N_12295,N_12391);
nor U12626 (N_12626,N_12259,N_12418);
nor U12627 (N_12627,N_12385,N_12343);
nor U12628 (N_12628,N_12326,N_12296);
nand U12629 (N_12629,N_12371,N_12307);
and U12630 (N_12630,N_12353,N_12478);
nor U12631 (N_12631,N_12464,N_12311);
nor U12632 (N_12632,N_12332,N_12417);
or U12633 (N_12633,N_12342,N_12347);
and U12634 (N_12634,N_12497,N_12355);
nand U12635 (N_12635,N_12260,N_12489);
xnor U12636 (N_12636,N_12451,N_12347);
and U12637 (N_12637,N_12258,N_12446);
nor U12638 (N_12638,N_12329,N_12276);
or U12639 (N_12639,N_12391,N_12433);
xnor U12640 (N_12640,N_12413,N_12439);
nand U12641 (N_12641,N_12426,N_12423);
nor U12642 (N_12642,N_12280,N_12424);
or U12643 (N_12643,N_12377,N_12278);
nor U12644 (N_12644,N_12375,N_12401);
nor U12645 (N_12645,N_12291,N_12331);
or U12646 (N_12646,N_12489,N_12418);
nor U12647 (N_12647,N_12382,N_12261);
and U12648 (N_12648,N_12453,N_12311);
and U12649 (N_12649,N_12470,N_12439);
and U12650 (N_12650,N_12482,N_12381);
nand U12651 (N_12651,N_12429,N_12466);
and U12652 (N_12652,N_12486,N_12352);
nor U12653 (N_12653,N_12258,N_12434);
nor U12654 (N_12654,N_12418,N_12373);
xnor U12655 (N_12655,N_12401,N_12302);
nand U12656 (N_12656,N_12299,N_12455);
or U12657 (N_12657,N_12342,N_12370);
or U12658 (N_12658,N_12363,N_12398);
and U12659 (N_12659,N_12319,N_12309);
xor U12660 (N_12660,N_12338,N_12381);
and U12661 (N_12661,N_12413,N_12299);
nand U12662 (N_12662,N_12464,N_12314);
xor U12663 (N_12663,N_12405,N_12341);
or U12664 (N_12664,N_12310,N_12382);
and U12665 (N_12665,N_12255,N_12495);
and U12666 (N_12666,N_12357,N_12426);
xor U12667 (N_12667,N_12390,N_12269);
and U12668 (N_12668,N_12255,N_12280);
nand U12669 (N_12669,N_12470,N_12494);
xor U12670 (N_12670,N_12389,N_12316);
nor U12671 (N_12671,N_12484,N_12302);
nor U12672 (N_12672,N_12339,N_12382);
and U12673 (N_12673,N_12273,N_12435);
or U12674 (N_12674,N_12342,N_12356);
xnor U12675 (N_12675,N_12499,N_12343);
and U12676 (N_12676,N_12365,N_12488);
and U12677 (N_12677,N_12365,N_12499);
and U12678 (N_12678,N_12488,N_12326);
nand U12679 (N_12679,N_12397,N_12414);
or U12680 (N_12680,N_12381,N_12384);
nor U12681 (N_12681,N_12470,N_12436);
nand U12682 (N_12682,N_12365,N_12420);
or U12683 (N_12683,N_12413,N_12459);
and U12684 (N_12684,N_12426,N_12274);
nor U12685 (N_12685,N_12343,N_12257);
or U12686 (N_12686,N_12467,N_12487);
or U12687 (N_12687,N_12418,N_12459);
xnor U12688 (N_12688,N_12382,N_12437);
or U12689 (N_12689,N_12317,N_12482);
nand U12690 (N_12690,N_12345,N_12430);
or U12691 (N_12691,N_12341,N_12270);
nand U12692 (N_12692,N_12498,N_12362);
nand U12693 (N_12693,N_12334,N_12311);
or U12694 (N_12694,N_12481,N_12422);
or U12695 (N_12695,N_12400,N_12260);
and U12696 (N_12696,N_12461,N_12499);
xnor U12697 (N_12697,N_12343,N_12429);
and U12698 (N_12698,N_12425,N_12444);
nor U12699 (N_12699,N_12486,N_12401);
nand U12700 (N_12700,N_12381,N_12366);
and U12701 (N_12701,N_12320,N_12300);
nand U12702 (N_12702,N_12376,N_12453);
and U12703 (N_12703,N_12486,N_12494);
xnor U12704 (N_12704,N_12349,N_12456);
or U12705 (N_12705,N_12286,N_12294);
or U12706 (N_12706,N_12288,N_12330);
and U12707 (N_12707,N_12411,N_12387);
nor U12708 (N_12708,N_12376,N_12472);
nand U12709 (N_12709,N_12448,N_12428);
and U12710 (N_12710,N_12390,N_12314);
xor U12711 (N_12711,N_12339,N_12361);
xor U12712 (N_12712,N_12327,N_12265);
or U12713 (N_12713,N_12328,N_12325);
nand U12714 (N_12714,N_12365,N_12469);
nor U12715 (N_12715,N_12490,N_12323);
and U12716 (N_12716,N_12481,N_12350);
nand U12717 (N_12717,N_12439,N_12419);
nor U12718 (N_12718,N_12484,N_12288);
xor U12719 (N_12719,N_12472,N_12415);
or U12720 (N_12720,N_12377,N_12470);
nor U12721 (N_12721,N_12477,N_12403);
and U12722 (N_12722,N_12295,N_12470);
xor U12723 (N_12723,N_12355,N_12393);
and U12724 (N_12724,N_12433,N_12469);
nor U12725 (N_12725,N_12405,N_12435);
nand U12726 (N_12726,N_12474,N_12336);
or U12727 (N_12727,N_12488,N_12293);
and U12728 (N_12728,N_12303,N_12260);
xor U12729 (N_12729,N_12298,N_12434);
and U12730 (N_12730,N_12310,N_12336);
and U12731 (N_12731,N_12438,N_12284);
nor U12732 (N_12732,N_12279,N_12411);
nand U12733 (N_12733,N_12313,N_12380);
nor U12734 (N_12734,N_12337,N_12379);
nand U12735 (N_12735,N_12366,N_12453);
or U12736 (N_12736,N_12269,N_12326);
and U12737 (N_12737,N_12387,N_12403);
or U12738 (N_12738,N_12270,N_12371);
xnor U12739 (N_12739,N_12338,N_12445);
or U12740 (N_12740,N_12300,N_12303);
xnor U12741 (N_12741,N_12346,N_12378);
nand U12742 (N_12742,N_12494,N_12304);
nand U12743 (N_12743,N_12297,N_12388);
nand U12744 (N_12744,N_12391,N_12252);
nor U12745 (N_12745,N_12320,N_12422);
nor U12746 (N_12746,N_12467,N_12337);
and U12747 (N_12747,N_12290,N_12378);
nor U12748 (N_12748,N_12444,N_12364);
or U12749 (N_12749,N_12281,N_12341);
nand U12750 (N_12750,N_12619,N_12656);
nor U12751 (N_12751,N_12731,N_12543);
nand U12752 (N_12752,N_12686,N_12623);
and U12753 (N_12753,N_12676,N_12661);
nand U12754 (N_12754,N_12624,N_12561);
nor U12755 (N_12755,N_12635,N_12627);
nand U12756 (N_12756,N_12654,N_12707);
nor U12757 (N_12757,N_12533,N_12601);
xor U12758 (N_12758,N_12515,N_12532);
nor U12759 (N_12759,N_12675,N_12735);
nor U12760 (N_12760,N_12650,N_12743);
or U12761 (N_12761,N_12663,N_12726);
nand U12762 (N_12762,N_12699,N_12598);
nor U12763 (N_12763,N_12683,N_12667);
or U12764 (N_12764,N_12727,N_12700);
xnor U12765 (N_12765,N_12556,N_12634);
and U12766 (N_12766,N_12510,N_12748);
xor U12767 (N_12767,N_12528,N_12722);
and U12768 (N_12768,N_12523,N_12689);
xnor U12769 (N_12769,N_12670,N_12617);
xor U12770 (N_12770,N_12549,N_12544);
or U12771 (N_12771,N_12606,N_12738);
nand U12772 (N_12772,N_12503,N_12733);
nand U12773 (N_12773,N_12567,N_12541);
nand U12774 (N_12774,N_12691,N_12604);
and U12775 (N_12775,N_12747,N_12698);
nand U12776 (N_12776,N_12580,N_12694);
or U12777 (N_12777,N_12653,N_12592);
or U12778 (N_12778,N_12512,N_12704);
or U12779 (N_12779,N_12578,N_12616);
or U12780 (N_12780,N_12520,N_12640);
nand U12781 (N_12781,N_12588,N_12516);
nand U12782 (N_12782,N_12701,N_12690);
and U12783 (N_12783,N_12552,N_12570);
or U12784 (N_12784,N_12711,N_12702);
or U12785 (N_12785,N_12706,N_12665);
xor U12786 (N_12786,N_12524,N_12594);
nand U12787 (N_12787,N_12553,N_12527);
nand U12788 (N_12788,N_12664,N_12557);
xnor U12789 (N_12789,N_12540,N_12697);
or U12790 (N_12790,N_12547,N_12657);
nor U12791 (N_12791,N_12692,N_12724);
and U12792 (N_12792,N_12521,N_12501);
and U12793 (N_12793,N_12680,N_12509);
nand U12794 (N_12794,N_12517,N_12639);
and U12795 (N_12795,N_12646,N_12749);
or U12796 (N_12796,N_12741,N_12551);
xor U12797 (N_12797,N_12530,N_12609);
or U12798 (N_12798,N_12630,N_12579);
xnor U12799 (N_12799,N_12576,N_12581);
nand U12800 (N_12800,N_12710,N_12622);
or U12801 (N_12801,N_12574,N_12648);
and U12802 (N_12802,N_12525,N_12560);
or U12803 (N_12803,N_12500,N_12573);
nor U12804 (N_12804,N_12720,N_12607);
or U12805 (N_12805,N_12638,N_12502);
nor U12806 (N_12806,N_12587,N_12746);
nor U12807 (N_12807,N_12569,N_12677);
nand U12808 (N_12808,N_12681,N_12734);
or U12809 (N_12809,N_12662,N_12531);
xor U12810 (N_12810,N_12596,N_12508);
nor U12811 (N_12811,N_12542,N_12687);
or U12812 (N_12812,N_12562,N_12513);
xor U12813 (N_12813,N_12545,N_12721);
nor U12814 (N_12814,N_12709,N_12673);
and U12815 (N_12815,N_12659,N_12614);
nor U12816 (N_12816,N_12636,N_12712);
xnor U12817 (N_12817,N_12685,N_12708);
and U12818 (N_12818,N_12565,N_12647);
xor U12819 (N_12819,N_12625,N_12688);
and U12820 (N_12820,N_12511,N_12572);
and U12821 (N_12821,N_12593,N_12526);
xor U12822 (N_12822,N_12589,N_12671);
or U12823 (N_12823,N_12714,N_12571);
nor U12824 (N_12824,N_12591,N_12739);
xnor U12825 (N_12825,N_12737,N_12705);
nand U12826 (N_12826,N_12534,N_12518);
nor U12827 (N_12827,N_12610,N_12716);
or U12828 (N_12828,N_12672,N_12555);
nand U12829 (N_12829,N_12548,N_12669);
xor U12830 (N_12830,N_12725,N_12558);
nand U12831 (N_12831,N_12641,N_12618);
nor U12832 (N_12832,N_12584,N_12608);
nor U12833 (N_12833,N_12583,N_12730);
nand U12834 (N_12834,N_12660,N_12719);
or U12835 (N_12835,N_12693,N_12695);
or U12836 (N_12836,N_12744,N_12713);
or U12837 (N_12837,N_12577,N_12504);
xor U12838 (N_12838,N_12679,N_12535);
nor U12839 (N_12839,N_12642,N_12736);
and U12840 (N_12840,N_12651,N_12684);
or U12841 (N_12841,N_12613,N_12633);
xor U12842 (N_12842,N_12703,N_12729);
nand U12843 (N_12843,N_12696,N_12546);
or U12844 (N_12844,N_12582,N_12529);
nor U12845 (N_12845,N_12507,N_12644);
nor U12846 (N_12846,N_12637,N_12728);
nor U12847 (N_12847,N_12599,N_12615);
nor U12848 (N_12848,N_12732,N_12514);
or U12849 (N_12849,N_12666,N_12575);
xnor U12850 (N_12850,N_12522,N_12559);
xor U12851 (N_12851,N_12519,N_12742);
nor U12852 (N_12852,N_12745,N_12643);
or U12853 (N_12853,N_12539,N_12629);
and U12854 (N_12854,N_12658,N_12717);
nor U12855 (N_12855,N_12612,N_12674);
xor U12856 (N_12856,N_12621,N_12632);
and U12857 (N_12857,N_12740,N_12537);
nor U12858 (N_12858,N_12586,N_12723);
xor U12859 (N_12859,N_12595,N_12611);
xnor U12860 (N_12860,N_12602,N_12585);
and U12861 (N_12861,N_12626,N_12649);
and U12862 (N_12862,N_12550,N_12563);
or U12863 (N_12863,N_12597,N_12568);
and U12864 (N_12864,N_12590,N_12628);
and U12865 (N_12865,N_12600,N_12718);
or U12866 (N_12866,N_12655,N_12554);
nand U12867 (N_12867,N_12620,N_12564);
and U12868 (N_12868,N_12603,N_12506);
or U12869 (N_12869,N_12715,N_12566);
or U12870 (N_12870,N_12538,N_12631);
and U12871 (N_12871,N_12678,N_12536);
and U12872 (N_12872,N_12668,N_12645);
nor U12873 (N_12873,N_12605,N_12652);
and U12874 (N_12874,N_12505,N_12682);
nor U12875 (N_12875,N_12504,N_12571);
nor U12876 (N_12876,N_12720,N_12609);
nor U12877 (N_12877,N_12721,N_12673);
nand U12878 (N_12878,N_12675,N_12515);
nor U12879 (N_12879,N_12733,N_12713);
and U12880 (N_12880,N_12743,N_12533);
and U12881 (N_12881,N_12722,N_12657);
or U12882 (N_12882,N_12697,N_12736);
and U12883 (N_12883,N_12525,N_12696);
nand U12884 (N_12884,N_12602,N_12714);
xor U12885 (N_12885,N_12550,N_12639);
xnor U12886 (N_12886,N_12721,N_12665);
nor U12887 (N_12887,N_12721,N_12533);
nand U12888 (N_12888,N_12645,N_12708);
xnor U12889 (N_12889,N_12604,N_12574);
xor U12890 (N_12890,N_12604,N_12597);
nand U12891 (N_12891,N_12589,N_12655);
nor U12892 (N_12892,N_12557,N_12668);
or U12893 (N_12893,N_12629,N_12698);
and U12894 (N_12894,N_12723,N_12503);
and U12895 (N_12895,N_12569,N_12609);
nand U12896 (N_12896,N_12725,N_12731);
nand U12897 (N_12897,N_12514,N_12572);
or U12898 (N_12898,N_12737,N_12671);
or U12899 (N_12899,N_12630,N_12674);
and U12900 (N_12900,N_12704,N_12642);
nand U12901 (N_12901,N_12637,N_12591);
and U12902 (N_12902,N_12716,N_12556);
nand U12903 (N_12903,N_12645,N_12502);
nand U12904 (N_12904,N_12611,N_12522);
or U12905 (N_12905,N_12689,N_12526);
nor U12906 (N_12906,N_12672,N_12625);
or U12907 (N_12907,N_12505,N_12560);
and U12908 (N_12908,N_12563,N_12672);
or U12909 (N_12909,N_12672,N_12690);
xnor U12910 (N_12910,N_12519,N_12579);
nor U12911 (N_12911,N_12724,N_12677);
nor U12912 (N_12912,N_12641,N_12696);
or U12913 (N_12913,N_12641,N_12713);
xor U12914 (N_12914,N_12651,N_12749);
xnor U12915 (N_12915,N_12661,N_12509);
xor U12916 (N_12916,N_12673,N_12637);
or U12917 (N_12917,N_12607,N_12590);
and U12918 (N_12918,N_12706,N_12596);
nand U12919 (N_12919,N_12543,N_12654);
nand U12920 (N_12920,N_12650,N_12684);
or U12921 (N_12921,N_12726,N_12644);
and U12922 (N_12922,N_12582,N_12560);
nand U12923 (N_12923,N_12511,N_12677);
and U12924 (N_12924,N_12584,N_12649);
nor U12925 (N_12925,N_12742,N_12713);
xor U12926 (N_12926,N_12540,N_12520);
and U12927 (N_12927,N_12708,N_12533);
nor U12928 (N_12928,N_12659,N_12742);
and U12929 (N_12929,N_12705,N_12603);
or U12930 (N_12930,N_12733,N_12596);
nor U12931 (N_12931,N_12653,N_12654);
nand U12932 (N_12932,N_12573,N_12560);
and U12933 (N_12933,N_12631,N_12615);
or U12934 (N_12934,N_12563,N_12592);
or U12935 (N_12935,N_12695,N_12657);
nand U12936 (N_12936,N_12663,N_12526);
xnor U12937 (N_12937,N_12631,N_12562);
or U12938 (N_12938,N_12580,N_12687);
or U12939 (N_12939,N_12626,N_12671);
nand U12940 (N_12940,N_12572,N_12685);
xor U12941 (N_12941,N_12617,N_12610);
xor U12942 (N_12942,N_12745,N_12673);
nand U12943 (N_12943,N_12522,N_12518);
nand U12944 (N_12944,N_12551,N_12738);
xnor U12945 (N_12945,N_12714,N_12541);
xor U12946 (N_12946,N_12667,N_12582);
nor U12947 (N_12947,N_12513,N_12661);
nand U12948 (N_12948,N_12605,N_12597);
xnor U12949 (N_12949,N_12705,N_12556);
nor U12950 (N_12950,N_12590,N_12585);
nor U12951 (N_12951,N_12589,N_12713);
or U12952 (N_12952,N_12666,N_12722);
and U12953 (N_12953,N_12596,N_12691);
nand U12954 (N_12954,N_12676,N_12745);
xnor U12955 (N_12955,N_12677,N_12726);
nor U12956 (N_12956,N_12651,N_12656);
and U12957 (N_12957,N_12746,N_12657);
nand U12958 (N_12958,N_12553,N_12614);
or U12959 (N_12959,N_12645,N_12523);
nand U12960 (N_12960,N_12527,N_12614);
or U12961 (N_12961,N_12567,N_12540);
nor U12962 (N_12962,N_12679,N_12670);
nor U12963 (N_12963,N_12695,N_12505);
xor U12964 (N_12964,N_12743,N_12562);
xor U12965 (N_12965,N_12682,N_12707);
or U12966 (N_12966,N_12553,N_12560);
xor U12967 (N_12967,N_12740,N_12651);
xor U12968 (N_12968,N_12711,N_12623);
nor U12969 (N_12969,N_12683,N_12642);
or U12970 (N_12970,N_12605,N_12737);
nand U12971 (N_12971,N_12672,N_12521);
and U12972 (N_12972,N_12575,N_12715);
nor U12973 (N_12973,N_12646,N_12676);
and U12974 (N_12974,N_12507,N_12603);
nand U12975 (N_12975,N_12572,N_12636);
or U12976 (N_12976,N_12592,N_12604);
nand U12977 (N_12977,N_12545,N_12661);
nor U12978 (N_12978,N_12514,N_12712);
xnor U12979 (N_12979,N_12700,N_12721);
nor U12980 (N_12980,N_12606,N_12731);
and U12981 (N_12981,N_12548,N_12578);
and U12982 (N_12982,N_12720,N_12598);
xnor U12983 (N_12983,N_12610,N_12718);
xor U12984 (N_12984,N_12697,N_12704);
xor U12985 (N_12985,N_12621,N_12595);
xor U12986 (N_12986,N_12508,N_12531);
nor U12987 (N_12987,N_12632,N_12545);
xor U12988 (N_12988,N_12622,N_12577);
xor U12989 (N_12989,N_12557,N_12631);
nand U12990 (N_12990,N_12684,N_12506);
nand U12991 (N_12991,N_12523,N_12694);
xor U12992 (N_12992,N_12663,N_12510);
xnor U12993 (N_12993,N_12710,N_12704);
or U12994 (N_12994,N_12675,N_12666);
nand U12995 (N_12995,N_12639,N_12630);
xor U12996 (N_12996,N_12625,N_12566);
xnor U12997 (N_12997,N_12643,N_12683);
xnor U12998 (N_12998,N_12729,N_12668);
or U12999 (N_12999,N_12664,N_12700);
nand U13000 (N_13000,N_12871,N_12811);
or U13001 (N_13001,N_12884,N_12752);
and U13002 (N_13002,N_12993,N_12788);
or U13003 (N_13003,N_12976,N_12923);
nor U13004 (N_13004,N_12964,N_12830);
nor U13005 (N_13005,N_12892,N_12781);
nand U13006 (N_13006,N_12889,N_12912);
or U13007 (N_13007,N_12835,N_12833);
or U13008 (N_13008,N_12821,N_12768);
xnor U13009 (N_13009,N_12972,N_12860);
nor U13010 (N_13010,N_12966,N_12981);
xor U13011 (N_13011,N_12828,N_12757);
or U13012 (N_13012,N_12777,N_12843);
nor U13013 (N_13013,N_12837,N_12775);
xor U13014 (N_13014,N_12822,N_12868);
or U13015 (N_13015,N_12787,N_12965);
and U13016 (N_13016,N_12987,N_12997);
nand U13017 (N_13017,N_12790,N_12797);
xor U13018 (N_13018,N_12883,N_12862);
nor U13019 (N_13019,N_12808,N_12975);
and U13020 (N_13020,N_12970,N_12967);
or U13021 (N_13021,N_12979,N_12971);
and U13022 (N_13022,N_12906,N_12824);
or U13023 (N_13023,N_12859,N_12818);
nor U13024 (N_13024,N_12815,N_12942);
xor U13025 (N_13025,N_12990,N_12956);
nor U13026 (N_13026,N_12928,N_12802);
nand U13027 (N_13027,N_12764,N_12769);
or U13028 (N_13028,N_12834,N_12766);
or U13029 (N_13029,N_12772,N_12849);
or U13030 (N_13030,N_12907,N_12973);
and U13031 (N_13031,N_12948,N_12844);
nor U13032 (N_13032,N_12897,N_12886);
nor U13033 (N_13033,N_12969,N_12831);
xor U13034 (N_13034,N_12845,N_12911);
and U13035 (N_13035,N_12957,N_12870);
and U13036 (N_13036,N_12899,N_12910);
nor U13037 (N_13037,N_12915,N_12995);
nand U13038 (N_13038,N_12991,N_12782);
or U13039 (N_13039,N_12994,N_12934);
and U13040 (N_13040,N_12959,N_12778);
xor U13041 (N_13041,N_12807,N_12930);
or U13042 (N_13042,N_12920,N_12945);
nand U13043 (N_13043,N_12767,N_12881);
or U13044 (N_13044,N_12874,N_12761);
and U13045 (N_13045,N_12864,N_12953);
nor U13046 (N_13046,N_12820,N_12756);
nor U13047 (N_13047,N_12776,N_12992);
nor U13048 (N_13048,N_12943,N_12983);
or U13049 (N_13049,N_12935,N_12898);
nor U13050 (N_13050,N_12861,N_12851);
nand U13051 (N_13051,N_12890,N_12875);
nand U13052 (N_13052,N_12853,N_12936);
nor U13053 (N_13053,N_12783,N_12784);
nor U13054 (N_13054,N_12937,N_12801);
or U13055 (N_13055,N_12917,N_12896);
nand U13056 (N_13056,N_12751,N_12809);
nand U13057 (N_13057,N_12939,N_12765);
xnor U13058 (N_13058,N_12872,N_12839);
xor U13059 (N_13059,N_12805,N_12867);
nand U13060 (N_13060,N_12893,N_12940);
nor U13061 (N_13061,N_12929,N_12825);
nand U13062 (N_13062,N_12977,N_12826);
and U13063 (N_13063,N_12963,N_12792);
nor U13064 (N_13064,N_12786,N_12858);
nand U13065 (N_13065,N_12998,N_12914);
nor U13066 (N_13066,N_12755,N_12789);
xnor U13067 (N_13067,N_12806,N_12799);
xnor U13068 (N_13068,N_12955,N_12773);
xor U13069 (N_13069,N_12954,N_12947);
nand U13070 (N_13070,N_12838,N_12978);
nand U13071 (N_13071,N_12932,N_12841);
and U13072 (N_13072,N_12840,N_12796);
or U13073 (N_13073,N_12924,N_12901);
or U13074 (N_13074,N_12869,N_12762);
nor U13075 (N_13075,N_12836,N_12895);
nor U13076 (N_13076,N_12800,N_12759);
xor U13077 (N_13077,N_12961,N_12779);
and U13078 (N_13078,N_12951,N_12996);
nand U13079 (N_13079,N_12829,N_12926);
nand U13080 (N_13080,N_12812,N_12949);
xor U13081 (N_13081,N_12985,N_12793);
nand U13082 (N_13082,N_12946,N_12863);
nand U13083 (N_13083,N_12832,N_12780);
nor U13084 (N_13084,N_12988,N_12952);
nand U13085 (N_13085,N_12882,N_12823);
and U13086 (N_13086,N_12760,N_12877);
and U13087 (N_13087,N_12904,N_12891);
and U13088 (N_13088,N_12927,N_12753);
nor U13089 (N_13089,N_12921,N_12804);
or U13090 (N_13090,N_12931,N_12887);
and U13091 (N_13091,N_12894,N_12850);
or U13092 (N_13092,N_12770,N_12922);
nor U13093 (N_13093,N_12908,N_12791);
nor U13094 (N_13094,N_12750,N_12879);
xnor U13095 (N_13095,N_12763,N_12857);
nor U13096 (N_13096,N_12758,N_12974);
xnor U13097 (N_13097,N_12810,N_12980);
nor U13098 (N_13098,N_12916,N_12986);
or U13099 (N_13099,N_12817,N_12885);
nand U13100 (N_13100,N_12933,N_12827);
nor U13101 (N_13101,N_12968,N_12880);
and U13102 (N_13102,N_12842,N_12794);
xor U13103 (N_13103,N_12847,N_12754);
nand U13104 (N_13104,N_12785,N_12846);
nand U13105 (N_13105,N_12771,N_12876);
and U13106 (N_13106,N_12960,N_12774);
nor U13107 (N_13107,N_12903,N_12803);
nand U13108 (N_13108,N_12962,N_12798);
and U13109 (N_13109,N_12856,N_12795);
or U13110 (N_13110,N_12813,N_12919);
or U13111 (N_13111,N_12944,N_12938);
or U13112 (N_13112,N_12866,N_12913);
nand U13113 (N_13113,N_12819,N_12984);
or U13114 (N_13114,N_12873,N_12918);
xor U13115 (N_13115,N_12902,N_12854);
xnor U13116 (N_13116,N_12888,N_12814);
nand U13117 (N_13117,N_12989,N_12950);
nor U13118 (N_13118,N_12982,N_12958);
nand U13119 (N_13119,N_12909,N_12852);
and U13120 (N_13120,N_12878,N_12855);
nand U13121 (N_13121,N_12900,N_12816);
and U13122 (N_13122,N_12941,N_12865);
or U13123 (N_13123,N_12999,N_12925);
xor U13124 (N_13124,N_12848,N_12905);
or U13125 (N_13125,N_12970,N_12908);
xor U13126 (N_13126,N_12825,N_12790);
nor U13127 (N_13127,N_12792,N_12927);
nor U13128 (N_13128,N_12840,N_12870);
nand U13129 (N_13129,N_12846,N_12893);
nor U13130 (N_13130,N_12811,N_12756);
nand U13131 (N_13131,N_12985,N_12788);
nor U13132 (N_13132,N_12907,N_12827);
or U13133 (N_13133,N_12895,N_12807);
xor U13134 (N_13134,N_12871,N_12810);
nand U13135 (N_13135,N_12897,N_12789);
xor U13136 (N_13136,N_12992,N_12850);
xor U13137 (N_13137,N_12883,N_12755);
or U13138 (N_13138,N_12989,N_12910);
nand U13139 (N_13139,N_12942,N_12906);
nor U13140 (N_13140,N_12980,N_12901);
nand U13141 (N_13141,N_12759,N_12905);
or U13142 (N_13142,N_12865,N_12786);
nand U13143 (N_13143,N_12880,N_12866);
xor U13144 (N_13144,N_12865,N_12953);
nor U13145 (N_13145,N_12833,N_12752);
xnor U13146 (N_13146,N_12987,N_12975);
nand U13147 (N_13147,N_12848,N_12846);
and U13148 (N_13148,N_12907,N_12842);
and U13149 (N_13149,N_12973,N_12825);
xor U13150 (N_13150,N_12981,N_12812);
or U13151 (N_13151,N_12890,N_12755);
and U13152 (N_13152,N_12946,N_12828);
or U13153 (N_13153,N_12834,N_12840);
nand U13154 (N_13154,N_12968,N_12930);
and U13155 (N_13155,N_12974,N_12839);
and U13156 (N_13156,N_12920,N_12772);
nand U13157 (N_13157,N_12939,N_12845);
nor U13158 (N_13158,N_12992,N_12761);
and U13159 (N_13159,N_12778,N_12886);
xor U13160 (N_13160,N_12874,N_12929);
nand U13161 (N_13161,N_12971,N_12773);
or U13162 (N_13162,N_12960,N_12945);
or U13163 (N_13163,N_12902,N_12805);
xor U13164 (N_13164,N_12985,N_12910);
and U13165 (N_13165,N_12929,N_12993);
nand U13166 (N_13166,N_12919,N_12842);
nor U13167 (N_13167,N_12820,N_12973);
xor U13168 (N_13168,N_12808,N_12840);
xor U13169 (N_13169,N_12995,N_12894);
nor U13170 (N_13170,N_12910,N_12851);
nor U13171 (N_13171,N_12838,N_12751);
xnor U13172 (N_13172,N_12805,N_12933);
nand U13173 (N_13173,N_12965,N_12792);
and U13174 (N_13174,N_12950,N_12909);
nand U13175 (N_13175,N_12970,N_12895);
or U13176 (N_13176,N_12945,N_12820);
and U13177 (N_13177,N_12954,N_12924);
xor U13178 (N_13178,N_12813,N_12784);
and U13179 (N_13179,N_12918,N_12962);
or U13180 (N_13180,N_12860,N_12794);
nand U13181 (N_13181,N_12761,N_12930);
or U13182 (N_13182,N_12835,N_12793);
nand U13183 (N_13183,N_12834,N_12831);
and U13184 (N_13184,N_12891,N_12812);
nand U13185 (N_13185,N_12897,N_12930);
nand U13186 (N_13186,N_12783,N_12816);
nand U13187 (N_13187,N_12861,N_12795);
or U13188 (N_13188,N_12893,N_12800);
or U13189 (N_13189,N_12946,N_12900);
and U13190 (N_13190,N_12979,N_12959);
nor U13191 (N_13191,N_12758,N_12787);
and U13192 (N_13192,N_12959,N_12787);
or U13193 (N_13193,N_12881,N_12995);
nand U13194 (N_13194,N_12785,N_12829);
or U13195 (N_13195,N_12760,N_12836);
nor U13196 (N_13196,N_12753,N_12828);
or U13197 (N_13197,N_12804,N_12780);
nand U13198 (N_13198,N_12864,N_12803);
nand U13199 (N_13199,N_12836,N_12851);
and U13200 (N_13200,N_12891,N_12752);
and U13201 (N_13201,N_12984,N_12912);
nor U13202 (N_13202,N_12767,N_12942);
nor U13203 (N_13203,N_12854,N_12977);
nor U13204 (N_13204,N_12865,N_12806);
or U13205 (N_13205,N_12882,N_12768);
or U13206 (N_13206,N_12929,N_12889);
nor U13207 (N_13207,N_12998,N_12839);
nand U13208 (N_13208,N_12806,N_12856);
nand U13209 (N_13209,N_12831,N_12948);
nor U13210 (N_13210,N_12858,N_12877);
and U13211 (N_13211,N_12894,N_12779);
or U13212 (N_13212,N_12930,N_12791);
or U13213 (N_13213,N_12831,N_12892);
xnor U13214 (N_13214,N_12989,N_12865);
xnor U13215 (N_13215,N_12992,N_12798);
nor U13216 (N_13216,N_12840,N_12992);
xor U13217 (N_13217,N_12941,N_12988);
nand U13218 (N_13218,N_12965,N_12838);
nand U13219 (N_13219,N_12934,N_12799);
nor U13220 (N_13220,N_12786,N_12981);
xor U13221 (N_13221,N_12989,N_12862);
xor U13222 (N_13222,N_12986,N_12903);
and U13223 (N_13223,N_12754,N_12980);
nor U13224 (N_13224,N_12784,N_12899);
xor U13225 (N_13225,N_12949,N_12781);
nor U13226 (N_13226,N_12908,N_12895);
xnor U13227 (N_13227,N_12795,N_12962);
and U13228 (N_13228,N_12932,N_12902);
nor U13229 (N_13229,N_12825,N_12814);
nor U13230 (N_13230,N_12797,N_12817);
nand U13231 (N_13231,N_12848,N_12917);
and U13232 (N_13232,N_12790,N_12774);
nand U13233 (N_13233,N_12923,N_12907);
xnor U13234 (N_13234,N_12842,N_12882);
and U13235 (N_13235,N_12875,N_12772);
xnor U13236 (N_13236,N_12913,N_12816);
xnor U13237 (N_13237,N_12870,N_12875);
nand U13238 (N_13238,N_12805,N_12854);
xnor U13239 (N_13239,N_12971,N_12906);
nand U13240 (N_13240,N_12825,N_12960);
or U13241 (N_13241,N_12931,N_12814);
and U13242 (N_13242,N_12925,N_12761);
nand U13243 (N_13243,N_12818,N_12948);
xor U13244 (N_13244,N_12811,N_12974);
xor U13245 (N_13245,N_12750,N_12842);
nor U13246 (N_13246,N_12968,N_12911);
xnor U13247 (N_13247,N_12832,N_12769);
xor U13248 (N_13248,N_12961,N_12892);
xnor U13249 (N_13249,N_12940,N_12971);
xor U13250 (N_13250,N_13151,N_13086);
nand U13251 (N_13251,N_13230,N_13225);
xnor U13252 (N_13252,N_13173,N_13073);
nand U13253 (N_13253,N_13050,N_13215);
and U13254 (N_13254,N_13197,N_13051);
xor U13255 (N_13255,N_13060,N_13011);
and U13256 (N_13256,N_13111,N_13201);
xnor U13257 (N_13257,N_13037,N_13226);
nor U13258 (N_13258,N_13216,N_13188);
and U13259 (N_13259,N_13057,N_13033);
nand U13260 (N_13260,N_13117,N_13077);
nand U13261 (N_13261,N_13032,N_13042);
nand U13262 (N_13262,N_13114,N_13192);
nor U13263 (N_13263,N_13135,N_13047);
xnor U13264 (N_13264,N_13180,N_13206);
nor U13265 (N_13265,N_13098,N_13001);
and U13266 (N_13266,N_13070,N_13132);
or U13267 (N_13267,N_13140,N_13222);
xor U13268 (N_13268,N_13103,N_13155);
and U13269 (N_13269,N_13150,N_13221);
nand U13270 (N_13270,N_13228,N_13016);
xnor U13271 (N_13271,N_13071,N_13119);
xnor U13272 (N_13272,N_13019,N_13021);
nor U13273 (N_13273,N_13058,N_13045);
nand U13274 (N_13274,N_13131,N_13249);
nor U13275 (N_13275,N_13167,N_13052);
or U13276 (N_13276,N_13189,N_13109);
nand U13277 (N_13277,N_13066,N_13059);
nand U13278 (N_13278,N_13072,N_13218);
nand U13279 (N_13279,N_13046,N_13208);
or U13280 (N_13280,N_13024,N_13194);
nand U13281 (N_13281,N_13010,N_13017);
xor U13282 (N_13282,N_13012,N_13003);
and U13283 (N_13283,N_13005,N_13023);
nand U13284 (N_13284,N_13061,N_13008);
nor U13285 (N_13285,N_13107,N_13013);
or U13286 (N_13286,N_13153,N_13095);
or U13287 (N_13287,N_13120,N_13231);
nand U13288 (N_13288,N_13078,N_13090);
or U13289 (N_13289,N_13105,N_13154);
or U13290 (N_13290,N_13092,N_13220);
or U13291 (N_13291,N_13136,N_13196);
xor U13292 (N_13292,N_13234,N_13067);
or U13293 (N_13293,N_13184,N_13123);
or U13294 (N_13294,N_13191,N_13161);
or U13295 (N_13295,N_13204,N_13079);
or U13296 (N_13296,N_13169,N_13193);
or U13297 (N_13297,N_13171,N_13101);
or U13298 (N_13298,N_13063,N_13202);
and U13299 (N_13299,N_13020,N_13049);
nand U13300 (N_13300,N_13183,N_13022);
and U13301 (N_13301,N_13246,N_13076);
xnor U13302 (N_13302,N_13243,N_13223);
xor U13303 (N_13303,N_13018,N_13178);
nand U13304 (N_13304,N_13043,N_13240);
xor U13305 (N_13305,N_13190,N_13121);
xnor U13306 (N_13306,N_13038,N_13144);
xnor U13307 (N_13307,N_13143,N_13235);
and U13308 (N_13308,N_13142,N_13091);
and U13309 (N_13309,N_13237,N_13083);
nor U13310 (N_13310,N_13162,N_13082);
nand U13311 (N_13311,N_13089,N_13242);
nand U13312 (N_13312,N_13233,N_13069);
and U13313 (N_13313,N_13214,N_13200);
and U13314 (N_13314,N_13207,N_13232);
nor U13315 (N_13315,N_13075,N_13165);
and U13316 (N_13316,N_13236,N_13080);
and U13317 (N_13317,N_13199,N_13148);
or U13318 (N_13318,N_13040,N_13124);
or U13319 (N_13319,N_13170,N_13035);
nand U13320 (N_13320,N_13068,N_13122);
xnor U13321 (N_13321,N_13127,N_13056);
xor U13322 (N_13322,N_13039,N_13177);
or U13323 (N_13323,N_13074,N_13026);
nor U13324 (N_13324,N_13000,N_13158);
nand U13325 (N_13325,N_13041,N_13108);
or U13326 (N_13326,N_13025,N_13146);
or U13327 (N_13327,N_13245,N_13128);
nand U13328 (N_13328,N_13044,N_13093);
nand U13329 (N_13329,N_13130,N_13096);
and U13330 (N_13330,N_13164,N_13247);
and U13331 (N_13331,N_13027,N_13084);
nand U13332 (N_13332,N_13203,N_13125);
nand U13333 (N_13333,N_13209,N_13172);
or U13334 (N_13334,N_13181,N_13007);
and U13335 (N_13335,N_13004,N_13137);
nor U13336 (N_13336,N_13248,N_13244);
nand U13337 (N_13337,N_13212,N_13157);
xor U13338 (N_13338,N_13210,N_13227);
or U13339 (N_13339,N_13166,N_13036);
and U13340 (N_13340,N_13168,N_13065);
and U13341 (N_13341,N_13085,N_13138);
nand U13342 (N_13342,N_13126,N_13100);
nand U13343 (N_13343,N_13029,N_13159);
nor U13344 (N_13344,N_13113,N_13015);
nor U13345 (N_13345,N_13149,N_13179);
xnor U13346 (N_13346,N_13106,N_13034);
or U13347 (N_13347,N_13134,N_13028);
xor U13348 (N_13348,N_13147,N_13115);
xor U13349 (N_13349,N_13133,N_13185);
nand U13350 (N_13350,N_13112,N_13099);
nand U13351 (N_13351,N_13053,N_13116);
or U13352 (N_13352,N_13102,N_13213);
or U13353 (N_13353,N_13219,N_13186);
or U13354 (N_13354,N_13176,N_13006);
xor U13355 (N_13355,N_13229,N_13163);
and U13356 (N_13356,N_13081,N_13064);
xor U13357 (N_13357,N_13088,N_13239);
and U13358 (N_13358,N_13104,N_13110);
nand U13359 (N_13359,N_13224,N_13174);
and U13360 (N_13360,N_13002,N_13139);
xor U13361 (N_13361,N_13009,N_13195);
xor U13362 (N_13362,N_13097,N_13030);
or U13363 (N_13363,N_13087,N_13156);
nor U13364 (N_13364,N_13241,N_13141);
and U13365 (N_13365,N_13205,N_13014);
nor U13366 (N_13366,N_13129,N_13175);
nor U13367 (N_13367,N_13054,N_13238);
nor U13368 (N_13368,N_13152,N_13031);
and U13369 (N_13369,N_13145,N_13211);
nor U13370 (N_13370,N_13187,N_13048);
and U13371 (N_13371,N_13055,N_13118);
xnor U13372 (N_13372,N_13094,N_13160);
nor U13373 (N_13373,N_13182,N_13198);
xnor U13374 (N_13374,N_13062,N_13217);
nor U13375 (N_13375,N_13129,N_13242);
xnor U13376 (N_13376,N_13132,N_13080);
nor U13377 (N_13377,N_13191,N_13202);
xnor U13378 (N_13378,N_13058,N_13066);
xnor U13379 (N_13379,N_13210,N_13063);
nor U13380 (N_13380,N_13164,N_13185);
or U13381 (N_13381,N_13004,N_13133);
nor U13382 (N_13382,N_13191,N_13037);
and U13383 (N_13383,N_13167,N_13012);
nor U13384 (N_13384,N_13103,N_13207);
or U13385 (N_13385,N_13247,N_13213);
nor U13386 (N_13386,N_13042,N_13055);
nor U13387 (N_13387,N_13048,N_13244);
xor U13388 (N_13388,N_13083,N_13071);
nand U13389 (N_13389,N_13121,N_13196);
nor U13390 (N_13390,N_13013,N_13064);
nor U13391 (N_13391,N_13079,N_13243);
nor U13392 (N_13392,N_13001,N_13169);
xnor U13393 (N_13393,N_13230,N_13111);
or U13394 (N_13394,N_13170,N_13140);
nor U13395 (N_13395,N_13173,N_13145);
nor U13396 (N_13396,N_13069,N_13190);
or U13397 (N_13397,N_13099,N_13177);
xor U13398 (N_13398,N_13164,N_13187);
and U13399 (N_13399,N_13013,N_13158);
nand U13400 (N_13400,N_13129,N_13123);
and U13401 (N_13401,N_13175,N_13066);
nor U13402 (N_13402,N_13161,N_13217);
and U13403 (N_13403,N_13075,N_13194);
nand U13404 (N_13404,N_13086,N_13177);
nor U13405 (N_13405,N_13094,N_13155);
nand U13406 (N_13406,N_13144,N_13054);
xor U13407 (N_13407,N_13113,N_13234);
xor U13408 (N_13408,N_13212,N_13040);
nand U13409 (N_13409,N_13178,N_13004);
and U13410 (N_13410,N_13023,N_13194);
nand U13411 (N_13411,N_13114,N_13093);
or U13412 (N_13412,N_13197,N_13102);
or U13413 (N_13413,N_13239,N_13134);
nor U13414 (N_13414,N_13109,N_13176);
or U13415 (N_13415,N_13104,N_13230);
and U13416 (N_13416,N_13246,N_13139);
nor U13417 (N_13417,N_13048,N_13085);
nor U13418 (N_13418,N_13117,N_13015);
nand U13419 (N_13419,N_13149,N_13163);
nand U13420 (N_13420,N_13189,N_13024);
nand U13421 (N_13421,N_13229,N_13131);
nand U13422 (N_13422,N_13205,N_13036);
xnor U13423 (N_13423,N_13058,N_13216);
or U13424 (N_13424,N_13019,N_13020);
nand U13425 (N_13425,N_13186,N_13175);
xor U13426 (N_13426,N_13023,N_13147);
xor U13427 (N_13427,N_13230,N_13020);
xnor U13428 (N_13428,N_13051,N_13119);
and U13429 (N_13429,N_13070,N_13034);
and U13430 (N_13430,N_13173,N_13165);
and U13431 (N_13431,N_13061,N_13241);
nor U13432 (N_13432,N_13162,N_13036);
or U13433 (N_13433,N_13082,N_13183);
xor U13434 (N_13434,N_13007,N_13077);
or U13435 (N_13435,N_13088,N_13042);
or U13436 (N_13436,N_13047,N_13004);
nor U13437 (N_13437,N_13112,N_13150);
and U13438 (N_13438,N_13206,N_13117);
or U13439 (N_13439,N_13130,N_13050);
and U13440 (N_13440,N_13186,N_13134);
nor U13441 (N_13441,N_13151,N_13045);
nand U13442 (N_13442,N_13091,N_13195);
or U13443 (N_13443,N_13160,N_13195);
nor U13444 (N_13444,N_13015,N_13201);
xnor U13445 (N_13445,N_13068,N_13104);
nand U13446 (N_13446,N_13166,N_13182);
nand U13447 (N_13447,N_13124,N_13085);
or U13448 (N_13448,N_13196,N_13246);
and U13449 (N_13449,N_13066,N_13028);
or U13450 (N_13450,N_13006,N_13013);
and U13451 (N_13451,N_13132,N_13091);
nand U13452 (N_13452,N_13170,N_13190);
nand U13453 (N_13453,N_13222,N_13211);
and U13454 (N_13454,N_13059,N_13231);
nand U13455 (N_13455,N_13175,N_13106);
and U13456 (N_13456,N_13197,N_13133);
nand U13457 (N_13457,N_13026,N_13018);
xor U13458 (N_13458,N_13047,N_13093);
nor U13459 (N_13459,N_13209,N_13040);
nor U13460 (N_13460,N_13156,N_13174);
and U13461 (N_13461,N_13063,N_13120);
xnor U13462 (N_13462,N_13092,N_13038);
xor U13463 (N_13463,N_13234,N_13191);
nor U13464 (N_13464,N_13063,N_13232);
nand U13465 (N_13465,N_13058,N_13195);
xor U13466 (N_13466,N_13034,N_13025);
or U13467 (N_13467,N_13117,N_13222);
nand U13468 (N_13468,N_13166,N_13097);
nor U13469 (N_13469,N_13023,N_13160);
xor U13470 (N_13470,N_13002,N_13183);
xor U13471 (N_13471,N_13087,N_13089);
xor U13472 (N_13472,N_13145,N_13075);
nor U13473 (N_13473,N_13093,N_13080);
nor U13474 (N_13474,N_13208,N_13246);
and U13475 (N_13475,N_13207,N_13048);
nand U13476 (N_13476,N_13240,N_13093);
and U13477 (N_13477,N_13019,N_13169);
nor U13478 (N_13478,N_13008,N_13085);
and U13479 (N_13479,N_13134,N_13163);
nor U13480 (N_13480,N_13175,N_13231);
nand U13481 (N_13481,N_13121,N_13238);
xor U13482 (N_13482,N_13210,N_13141);
xor U13483 (N_13483,N_13220,N_13024);
nor U13484 (N_13484,N_13054,N_13176);
and U13485 (N_13485,N_13226,N_13247);
xor U13486 (N_13486,N_13024,N_13076);
nor U13487 (N_13487,N_13220,N_13238);
or U13488 (N_13488,N_13111,N_13147);
or U13489 (N_13489,N_13058,N_13246);
and U13490 (N_13490,N_13135,N_13160);
and U13491 (N_13491,N_13119,N_13009);
or U13492 (N_13492,N_13241,N_13225);
nand U13493 (N_13493,N_13221,N_13045);
nor U13494 (N_13494,N_13101,N_13216);
nand U13495 (N_13495,N_13109,N_13142);
nor U13496 (N_13496,N_13107,N_13245);
nand U13497 (N_13497,N_13022,N_13161);
xor U13498 (N_13498,N_13105,N_13095);
nand U13499 (N_13499,N_13215,N_13078);
xor U13500 (N_13500,N_13449,N_13459);
and U13501 (N_13501,N_13446,N_13375);
nor U13502 (N_13502,N_13488,N_13489);
and U13503 (N_13503,N_13405,N_13484);
xnor U13504 (N_13504,N_13250,N_13477);
xnor U13505 (N_13505,N_13291,N_13454);
and U13506 (N_13506,N_13279,N_13347);
and U13507 (N_13507,N_13326,N_13403);
and U13508 (N_13508,N_13378,N_13401);
and U13509 (N_13509,N_13428,N_13303);
nand U13510 (N_13510,N_13338,N_13260);
nand U13511 (N_13511,N_13388,N_13340);
or U13512 (N_13512,N_13299,N_13476);
xor U13513 (N_13513,N_13381,N_13386);
or U13514 (N_13514,N_13302,N_13322);
xor U13515 (N_13515,N_13370,N_13290);
or U13516 (N_13516,N_13461,N_13305);
and U13517 (N_13517,N_13486,N_13392);
and U13518 (N_13518,N_13493,N_13409);
or U13519 (N_13519,N_13438,N_13481);
nand U13520 (N_13520,N_13376,N_13464);
xor U13521 (N_13521,N_13437,N_13344);
and U13522 (N_13522,N_13342,N_13424);
xnor U13523 (N_13523,N_13465,N_13274);
or U13524 (N_13524,N_13447,N_13293);
nor U13525 (N_13525,N_13468,N_13318);
nand U13526 (N_13526,N_13374,N_13479);
and U13527 (N_13527,N_13373,N_13275);
xnor U13528 (N_13528,N_13263,N_13445);
or U13529 (N_13529,N_13289,N_13482);
nand U13530 (N_13530,N_13496,N_13491);
nand U13531 (N_13531,N_13255,N_13295);
or U13532 (N_13532,N_13404,N_13483);
xnor U13533 (N_13533,N_13257,N_13492);
xnor U13534 (N_13534,N_13329,N_13287);
nor U13535 (N_13535,N_13470,N_13414);
xnor U13536 (N_13536,N_13252,N_13394);
and U13537 (N_13537,N_13306,N_13314);
and U13538 (N_13538,N_13367,N_13389);
xor U13539 (N_13539,N_13364,N_13431);
and U13540 (N_13540,N_13460,N_13412);
nand U13541 (N_13541,N_13312,N_13282);
xor U13542 (N_13542,N_13360,N_13321);
nand U13543 (N_13543,N_13408,N_13485);
xnor U13544 (N_13544,N_13363,N_13472);
or U13545 (N_13545,N_13361,N_13425);
and U13546 (N_13546,N_13390,N_13422);
and U13547 (N_13547,N_13264,N_13372);
or U13548 (N_13548,N_13297,N_13358);
xnor U13549 (N_13549,N_13308,N_13272);
nor U13550 (N_13550,N_13396,N_13448);
nor U13551 (N_13551,N_13262,N_13383);
and U13552 (N_13552,N_13490,N_13324);
xor U13553 (N_13553,N_13443,N_13456);
and U13554 (N_13554,N_13377,N_13391);
nor U13555 (N_13555,N_13284,N_13379);
or U13556 (N_13556,N_13467,N_13296);
and U13557 (N_13557,N_13265,N_13382);
and U13558 (N_13558,N_13330,N_13256);
nor U13559 (N_13559,N_13385,N_13328);
or U13560 (N_13560,N_13339,N_13353);
nor U13561 (N_13561,N_13271,N_13371);
xnor U13562 (N_13562,N_13395,N_13301);
or U13563 (N_13563,N_13410,N_13427);
nand U13564 (N_13564,N_13354,N_13327);
xor U13565 (N_13565,N_13345,N_13475);
or U13566 (N_13566,N_13288,N_13268);
nand U13567 (N_13567,N_13309,N_13463);
nand U13568 (N_13568,N_13341,N_13399);
xnor U13569 (N_13569,N_13286,N_13458);
and U13570 (N_13570,N_13254,N_13436);
xor U13571 (N_13571,N_13429,N_13320);
or U13572 (N_13572,N_13259,N_13304);
or U13573 (N_13573,N_13285,N_13368);
or U13574 (N_13574,N_13397,N_13407);
xnor U13575 (N_13575,N_13450,N_13380);
or U13576 (N_13576,N_13315,N_13319);
nand U13577 (N_13577,N_13426,N_13300);
xor U13578 (N_13578,N_13499,N_13495);
xnor U13579 (N_13579,N_13417,N_13267);
and U13580 (N_13580,N_13270,N_13433);
nor U13581 (N_13581,N_13423,N_13421);
xor U13582 (N_13582,N_13440,N_13384);
and U13583 (N_13583,N_13452,N_13335);
xnor U13584 (N_13584,N_13451,N_13469);
xor U13585 (N_13585,N_13273,N_13439);
nor U13586 (N_13586,N_13416,N_13498);
and U13587 (N_13587,N_13334,N_13455);
or U13588 (N_13588,N_13462,N_13292);
nand U13589 (N_13589,N_13473,N_13434);
nand U13590 (N_13590,N_13415,N_13356);
nand U13591 (N_13591,N_13253,N_13346);
and U13592 (N_13592,N_13336,N_13413);
nor U13593 (N_13593,N_13294,N_13317);
nand U13594 (N_13594,N_13350,N_13352);
nor U13595 (N_13595,N_13359,N_13369);
nor U13596 (N_13596,N_13280,N_13420);
nor U13597 (N_13597,N_13400,N_13349);
nor U13598 (N_13598,N_13365,N_13251);
and U13599 (N_13599,N_13487,N_13269);
nor U13600 (N_13600,N_13419,N_13266);
xnor U13601 (N_13601,N_13362,N_13457);
or U13602 (N_13602,N_13310,N_13337);
or U13603 (N_13603,N_13283,N_13466);
nor U13604 (N_13604,N_13333,N_13343);
and U13605 (N_13605,N_13281,N_13357);
nor U13606 (N_13606,N_13398,N_13307);
and U13607 (N_13607,N_13430,N_13471);
nor U13608 (N_13608,N_13480,N_13402);
nor U13609 (N_13609,N_13278,N_13316);
or U13610 (N_13610,N_13442,N_13348);
xor U13611 (N_13611,N_13298,N_13387);
xor U13612 (N_13612,N_13435,N_13311);
and U13613 (N_13613,N_13323,N_13277);
xor U13614 (N_13614,N_13497,N_13411);
xor U13615 (N_13615,N_13261,N_13406);
xnor U13616 (N_13616,N_13351,N_13366);
nor U13617 (N_13617,N_13332,N_13453);
or U13618 (N_13618,N_13355,N_13441);
and U13619 (N_13619,N_13474,N_13313);
nor U13620 (N_13620,N_13432,N_13393);
nand U13621 (N_13621,N_13494,N_13418);
and U13622 (N_13622,N_13331,N_13258);
nand U13623 (N_13623,N_13444,N_13276);
and U13624 (N_13624,N_13325,N_13478);
nand U13625 (N_13625,N_13434,N_13367);
and U13626 (N_13626,N_13366,N_13392);
nor U13627 (N_13627,N_13376,N_13449);
nor U13628 (N_13628,N_13304,N_13491);
nand U13629 (N_13629,N_13266,N_13432);
and U13630 (N_13630,N_13364,N_13323);
nor U13631 (N_13631,N_13367,N_13302);
xnor U13632 (N_13632,N_13470,N_13424);
or U13633 (N_13633,N_13346,N_13437);
or U13634 (N_13634,N_13308,N_13426);
nand U13635 (N_13635,N_13428,N_13493);
nor U13636 (N_13636,N_13493,N_13364);
xor U13637 (N_13637,N_13312,N_13359);
nand U13638 (N_13638,N_13410,N_13481);
nor U13639 (N_13639,N_13309,N_13302);
xor U13640 (N_13640,N_13339,N_13322);
nor U13641 (N_13641,N_13435,N_13343);
nor U13642 (N_13642,N_13275,N_13401);
nand U13643 (N_13643,N_13393,N_13486);
and U13644 (N_13644,N_13334,N_13333);
or U13645 (N_13645,N_13347,N_13485);
xor U13646 (N_13646,N_13454,N_13345);
nor U13647 (N_13647,N_13432,N_13250);
xor U13648 (N_13648,N_13308,N_13393);
nor U13649 (N_13649,N_13426,N_13302);
nor U13650 (N_13650,N_13269,N_13348);
and U13651 (N_13651,N_13417,N_13415);
xor U13652 (N_13652,N_13422,N_13465);
xor U13653 (N_13653,N_13262,N_13284);
nand U13654 (N_13654,N_13480,N_13370);
or U13655 (N_13655,N_13372,N_13311);
nor U13656 (N_13656,N_13318,N_13494);
xor U13657 (N_13657,N_13269,N_13367);
nor U13658 (N_13658,N_13374,N_13427);
xor U13659 (N_13659,N_13438,N_13490);
nor U13660 (N_13660,N_13417,N_13356);
nand U13661 (N_13661,N_13298,N_13366);
nand U13662 (N_13662,N_13400,N_13389);
and U13663 (N_13663,N_13255,N_13473);
or U13664 (N_13664,N_13359,N_13381);
nand U13665 (N_13665,N_13284,N_13407);
xor U13666 (N_13666,N_13491,N_13418);
nand U13667 (N_13667,N_13483,N_13452);
and U13668 (N_13668,N_13271,N_13347);
and U13669 (N_13669,N_13380,N_13375);
or U13670 (N_13670,N_13257,N_13380);
and U13671 (N_13671,N_13420,N_13458);
nor U13672 (N_13672,N_13491,N_13317);
nor U13673 (N_13673,N_13258,N_13292);
nand U13674 (N_13674,N_13306,N_13405);
or U13675 (N_13675,N_13450,N_13428);
xnor U13676 (N_13676,N_13484,N_13416);
or U13677 (N_13677,N_13255,N_13380);
xor U13678 (N_13678,N_13330,N_13446);
and U13679 (N_13679,N_13260,N_13302);
or U13680 (N_13680,N_13365,N_13373);
or U13681 (N_13681,N_13250,N_13404);
and U13682 (N_13682,N_13412,N_13484);
and U13683 (N_13683,N_13282,N_13485);
nand U13684 (N_13684,N_13300,N_13313);
nor U13685 (N_13685,N_13363,N_13299);
and U13686 (N_13686,N_13410,N_13464);
nand U13687 (N_13687,N_13425,N_13410);
nor U13688 (N_13688,N_13251,N_13384);
and U13689 (N_13689,N_13499,N_13437);
xor U13690 (N_13690,N_13300,N_13483);
nand U13691 (N_13691,N_13395,N_13397);
or U13692 (N_13692,N_13484,N_13382);
and U13693 (N_13693,N_13459,N_13439);
and U13694 (N_13694,N_13491,N_13364);
nor U13695 (N_13695,N_13433,N_13277);
xnor U13696 (N_13696,N_13377,N_13317);
nand U13697 (N_13697,N_13355,N_13474);
nor U13698 (N_13698,N_13277,N_13437);
and U13699 (N_13699,N_13305,N_13407);
or U13700 (N_13700,N_13480,N_13422);
and U13701 (N_13701,N_13492,N_13455);
xnor U13702 (N_13702,N_13346,N_13495);
nor U13703 (N_13703,N_13320,N_13439);
nor U13704 (N_13704,N_13368,N_13459);
nor U13705 (N_13705,N_13279,N_13482);
xnor U13706 (N_13706,N_13304,N_13382);
nor U13707 (N_13707,N_13326,N_13270);
and U13708 (N_13708,N_13425,N_13253);
or U13709 (N_13709,N_13250,N_13396);
nor U13710 (N_13710,N_13281,N_13278);
nand U13711 (N_13711,N_13322,N_13334);
xnor U13712 (N_13712,N_13424,N_13273);
xor U13713 (N_13713,N_13318,N_13297);
nor U13714 (N_13714,N_13441,N_13367);
xnor U13715 (N_13715,N_13285,N_13340);
nand U13716 (N_13716,N_13381,N_13273);
or U13717 (N_13717,N_13284,N_13258);
nand U13718 (N_13718,N_13263,N_13319);
nand U13719 (N_13719,N_13342,N_13259);
nand U13720 (N_13720,N_13451,N_13396);
nand U13721 (N_13721,N_13346,N_13466);
nand U13722 (N_13722,N_13442,N_13325);
nand U13723 (N_13723,N_13373,N_13388);
nor U13724 (N_13724,N_13339,N_13401);
nor U13725 (N_13725,N_13294,N_13444);
nor U13726 (N_13726,N_13283,N_13297);
nor U13727 (N_13727,N_13330,N_13486);
xor U13728 (N_13728,N_13449,N_13273);
xnor U13729 (N_13729,N_13481,N_13311);
or U13730 (N_13730,N_13499,N_13339);
or U13731 (N_13731,N_13311,N_13335);
nand U13732 (N_13732,N_13367,N_13432);
nor U13733 (N_13733,N_13472,N_13282);
nor U13734 (N_13734,N_13325,N_13446);
and U13735 (N_13735,N_13418,N_13329);
and U13736 (N_13736,N_13275,N_13446);
nor U13737 (N_13737,N_13473,N_13491);
xnor U13738 (N_13738,N_13308,N_13381);
xor U13739 (N_13739,N_13383,N_13278);
or U13740 (N_13740,N_13402,N_13498);
and U13741 (N_13741,N_13256,N_13329);
or U13742 (N_13742,N_13491,N_13253);
and U13743 (N_13743,N_13270,N_13383);
and U13744 (N_13744,N_13487,N_13303);
and U13745 (N_13745,N_13347,N_13302);
and U13746 (N_13746,N_13353,N_13449);
and U13747 (N_13747,N_13410,N_13339);
nand U13748 (N_13748,N_13422,N_13284);
and U13749 (N_13749,N_13374,N_13491);
and U13750 (N_13750,N_13644,N_13574);
nand U13751 (N_13751,N_13746,N_13711);
xor U13752 (N_13752,N_13560,N_13501);
xnor U13753 (N_13753,N_13611,N_13518);
and U13754 (N_13754,N_13582,N_13689);
nand U13755 (N_13755,N_13536,N_13655);
or U13756 (N_13756,N_13683,N_13537);
nand U13757 (N_13757,N_13595,N_13699);
nor U13758 (N_13758,N_13717,N_13728);
and U13759 (N_13759,N_13712,N_13718);
xnor U13760 (N_13760,N_13734,N_13620);
xnor U13761 (N_13761,N_13538,N_13657);
or U13762 (N_13762,N_13552,N_13740);
and U13763 (N_13763,N_13569,N_13545);
nor U13764 (N_13764,N_13523,N_13573);
and U13765 (N_13765,N_13708,N_13615);
nor U13766 (N_13766,N_13621,N_13547);
nor U13767 (N_13767,N_13736,N_13589);
xor U13768 (N_13768,N_13727,N_13730);
and U13769 (N_13769,N_13558,N_13515);
nor U13770 (N_13770,N_13576,N_13745);
or U13771 (N_13771,N_13667,N_13610);
xnor U13772 (N_13772,N_13668,N_13660);
or U13773 (N_13773,N_13663,N_13577);
xnor U13774 (N_13774,N_13700,N_13679);
nand U13775 (N_13775,N_13642,N_13529);
and U13776 (N_13776,N_13629,N_13672);
or U13777 (N_13777,N_13594,N_13648);
or U13778 (N_13778,N_13540,N_13692);
nor U13779 (N_13779,N_13721,N_13739);
and U13780 (N_13780,N_13680,N_13639);
nand U13781 (N_13781,N_13720,N_13659);
xor U13782 (N_13782,N_13505,N_13618);
nor U13783 (N_13783,N_13617,N_13517);
or U13784 (N_13784,N_13521,N_13693);
or U13785 (N_13785,N_13698,N_13656);
xnor U13786 (N_13786,N_13563,N_13530);
nor U13787 (N_13787,N_13670,N_13592);
nand U13788 (N_13788,N_13666,N_13599);
or U13789 (N_13789,N_13645,N_13612);
and U13790 (N_13790,N_13604,N_13622);
and U13791 (N_13791,N_13519,N_13535);
or U13792 (N_13792,N_13635,N_13516);
and U13793 (N_13793,N_13676,N_13714);
or U13794 (N_13794,N_13743,N_13562);
or U13795 (N_13795,N_13633,N_13735);
and U13796 (N_13796,N_13571,N_13559);
and U13797 (N_13797,N_13598,N_13682);
and U13798 (N_13798,N_13502,N_13684);
nor U13799 (N_13799,N_13691,N_13688);
nand U13800 (N_13800,N_13681,N_13677);
xor U13801 (N_13801,N_13747,N_13634);
or U13802 (N_13802,N_13719,N_13555);
or U13803 (N_13803,N_13614,N_13565);
xor U13804 (N_13804,N_13546,N_13627);
nor U13805 (N_13805,N_13525,N_13626);
nand U13806 (N_13806,N_13613,N_13588);
nor U13807 (N_13807,N_13715,N_13570);
xor U13808 (N_13808,N_13543,N_13685);
nor U13809 (N_13809,N_13605,N_13556);
and U13810 (N_13810,N_13528,N_13616);
nand U13811 (N_13811,N_13632,N_13504);
nand U13812 (N_13812,N_13726,N_13513);
nand U13813 (N_13813,N_13653,N_13514);
xnor U13814 (N_13814,N_13609,N_13686);
nor U13815 (N_13815,N_13650,N_13703);
or U13816 (N_13816,N_13586,N_13646);
and U13817 (N_13817,N_13671,N_13548);
nand U13818 (N_13818,N_13500,N_13637);
or U13819 (N_13819,N_13640,N_13597);
nand U13820 (N_13820,N_13673,N_13600);
nor U13821 (N_13821,N_13511,N_13596);
and U13822 (N_13822,N_13579,N_13506);
xor U13823 (N_13823,N_13695,N_13580);
xor U13824 (N_13824,N_13707,N_13606);
and U13825 (N_13825,N_13702,N_13625);
nand U13826 (N_13826,N_13531,N_13510);
nor U13827 (N_13827,N_13549,N_13520);
xor U13828 (N_13828,N_13508,N_13624);
or U13829 (N_13829,N_13704,N_13738);
nor U13830 (N_13830,N_13553,N_13722);
nand U13831 (N_13831,N_13705,N_13664);
or U13832 (N_13832,N_13534,N_13723);
and U13833 (N_13833,N_13697,N_13716);
nand U13834 (N_13834,N_13643,N_13593);
or U13835 (N_13835,N_13527,N_13578);
or U13836 (N_13836,N_13742,N_13602);
or U13837 (N_13837,N_13607,N_13503);
and U13838 (N_13838,N_13690,N_13591);
nand U13839 (N_13839,N_13628,N_13674);
nand U13840 (N_13840,N_13512,N_13636);
and U13841 (N_13841,N_13631,N_13678);
or U13842 (N_13842,N_13741,N_13572);
nor U13843 (N_13843,N_13647,N_13585);
and U13844 (N_13844,N_13732,N_13564);
and U13845 (N_13845,N_13524,N_13551);
nor U13846 (N_13846,N_13661,N_13675);
or U13847 (N_13847,N_13541,N_13603);
xor U13848 (N_13848,N_13638,N_13557);
and U13849 (N_13849,N_13561,N_13729);
and U13850 (N_13850,N_13507,N_13567);
and U13851 (N_13851,N_13584,N_13566);
nor U13852 (N_13852,N_13608,N_13619);
nand U13853 (N_13853,N_13737,N_13694);
or U13854 (N_13854,N_13554,N_13601);
nor U13855 (N_13855,N_13696,N_13590);
xnor U13856 (N_13856,N_13669,N_13533);
and U13857 (N_13857,N_13744,N_13724);
nand U13858 (N_13858,N_13649,N_13522);
and U13859 (N_13859,N_13542,N_13550);
and U13860 (N_13860,N_13733,N_13748);
nor U13861 (N_13861,N_13568,N_13709);
xor U13862 (N_13862,N_13731,N_13641);
nand U13863 (N_13863,N_13575,N_13652);
nand U13864 (N_13864,N_13687,N_13539);
and U13865 (N_13865,N_13532,N_13710);
nand U13866 (N_13866,N_13701,N_13658);
xnor U13867 (N_13867,N_13706,N_13654);
nor U13868 (N_13868,N_13749,N_13665);
nor U13869 (N_13869,N_13630,N_13526);
and U13870 (N_13870,N_13623,N_13713);
xor U13871 (N_13871,N_13509,N_13587);
nand U13872 (N_13872,N_13583,N_13581);
and U13873 (N_13873,N_13662,N_13725);
nand U13874 (N_13874,N_13544,N_13651);
nand U13875 (N_13875,N_13734,N_13682);
and U13876 (N_13876,N_13591,N_13746);
xnor U13877 (N_13877,N_13528,N_13728);
xor U13878 (N_13878,N_13636,N_13685);
nand U13879 (N_13879,N_13660,N_13616);
xnor U13880 (N_13880,N_13710,N_13736);
nor U13881 (N_13881,N_13593,N_13601);
and U13882 (N_13882,N_13570,N_13548);
xor U13883 (N_13883,N_13531,N_13591);
and U13884 (N_13884,N_13576,N_13692);
or U13885 (N_13885,N_13670,N_13504);
nand U13886 (N_13886,N_13569,N_13518);
nand U13887 (N_13887,N_13560,N_13676);
and U13888 (N_13888,N_13713,N_13687);
xnor U13889 (N_13889,N_13680,N_13656);
nor U13890 (N_13890,N_13588,N_13586);
and U13891 (N_13891,N_13597,N_13528);
and U13892 (N_13892,N_13534,N_13517);
or U13893 (N_13893,N_13546,N_13611);
or U13894 (N_13894,N_13654,N_13574);
nor U13895 (N_13895,N_13697,N_13668);
and U13896 (N_13896,N_13527,N_13638);
nand U13897 (N_13897,N_13540,N_13711);
and U13898 (N_13898,N_13647,N_13631);
or U13899 (N_13899,N_13571,N_13658);
xor U13900 (N_13900,N_13612,N_13513);
or U13901 (N_13901,N_13673,N_13517);
xor U13902 (N_13902,N_13712,N_13687);
or U13903 (N_13903,N_13661,N_13745);
or U13904 (N_13904,N_13648,N_13552);
and U13905 (N_13905,N_13579,N_13607);
xor U13906 (N_13906,N_13616,N_13535);
and U13907 (N_13907,N_13659,N_13722);
nor U13908 (N_13908,N_13593,N_13603);
and U13909 (N_13909,N_13569,N_13508);
or U13910 (N_13910,N_13642,N_13620);
nor U13911 (N_13911,N_13697,N_13560);
nand U13912 (N_13912,N_13732,N_13539);
or U13913 (N_13913,N_13668,N_13649);
or U13914 (N_13914,N_13538,N_13695);
or U13915 (N_13915,N_13504,N_13592);
or U13916 (N_13916,N_13705,N_13594);
xor U13917 (N_13917,N_13569,N_13541);
or U13918 (N_13918,N_13532,N_13543);
nor U13919 (N_13919,N_13593,N_13533);
nand U13920 (N_13920,N_13710,N_13722);
and U13921 (N_13921,N_13551,N_13725);
xnor U13922 (N_13922,N_13656,N_13551);
nor U13923 (N_13923,N_13593,N_13705);
xnor U13924 (N_13924,N_13736,N_13564);
xor U13925 (N_13925,N_13565,N_13610);
nand U13926 (N_13926,N_13745,N_13548);
xor U13927 (N_13927,N_13746,N_13563);
xnor U13928 (N_13928,N_13573,N_13716);
nand U13929 (N_13929,N_13566,N_13630);
xor U13930 (N_13930,N_13694,N_13675);
and U13931 (N_13931,N_13508,N_13690);
and U13932 (N_13932,N_13551,N_13617);
nor U13933 (N_13933,N_13570,N_13708);
nor U13934 (N_13934,N_13658,N_13603);
and U13935 (N_13935,N_13611,N_13644);
xnor U13936 (N_13936,N_13672,N_13684);
nand U13937 (N_13937,N_13593,N_13576);
xnor U13938 (N_13938,N_13676,N_13517);
and U13939 (N_13939,N_13718,N_13597);
nand U13940 (N_13940,N_13692,N_13647);
xnor U13941 (N_13941,N_13688,N_13509);
nor U13942 (N_13942,N_13637,N_13563);
or U13943 (N_13943,N_13560,N_13656);
and U13944 (N_13944,N_13685,N_13637);
nand U13945 (N_13945,N_13507,N_13706);
nor U13946 (N_13946,N_13558,N_13516);
or U13947 (N_13947,N_13691,N_13507);
nor U13948 (N_13948,N_13656,N_13696);
nor U13949 (N_13949,N_13695,N_13537);
and U13950 (N_13950,N_13703,N_13583);
nor U13951 (N_13951,N_13619,N_13618);
xor U13952 (N_13952,N_13656,N_13564);
nand U13953 (N_13953,N_13653,N_13584);
and U13954 (N_13954,N_13560,N_13633);
nor U13955 (N_13955,N_13624,N_13639);
or U13956 (N_13956,N_13568,N_13646);
nand U13957 (N_13957,N_13692,N_13650);
nor U13958 (N_13958,N_13690,N_13552);
and U13959 (N_13959,N_13581,N_13675);
xor U13960 (N_13960,N_13645,N_13580);
nand U13961 (N_13961,N_13624,N_13586);
or U13962 (N_13962,N_13519,N_13544);
xnor U13963 (N_13963,N_13618,N_13532);
xor U13964 (N_13964,N_13639,N_13521);
or U13965 (N_13965,N_13592,N_13704);
nand U13966 (N_13966,N_13696,N_13531);
nor U13967 (N_13967,N_13706,N_13517);
xor U13968 (N_13968,N_13541,N_13653);
nand U13969 (N_13969,N_13548,N_13615);
xor U13970 (N_13970,N_13725,N_13647);
nor U13971 (N_13971,N_13571,N_13652);
or U13972 (N_13972,N_13702,N_13543);
or U13973 (N_13973,N_13734,N_13716);
and U13974 (N_13974,N_13529,N_13567);
xnor U13975 (N_13975,N_13650,N_13514);
and U13976 (N_13976,N_13703,N_13592);
nor U13977 (N_13977,N_13595,N_13553);
and U13978 (N_13978,N_13682,N_13736);
or U13979 (N_13979,N_13584,N_13583);
nor U13980 (N_13980,N_13540,N_13550);
nor U13981 (N_13981,N_13689,N_13516);
nand U13982 (N_13982,N_13503,N_13504);
xor U13983 (N_13983,N_13689,N_13586);
and U13984 (N_13984,N_13727,N_13686);
or U13985 (N_13985,N_13742,N_13685);
nand U13986 (N_13986,N_13664,N_13505);
or U13987 (N_13987,N_13698,N_13745);
and U13988 (N_13988,N_13553,N_13528);
xnor U13989 (N_13989,N_13679,N_13518);
nor U13990 (N_13990,N_13529,N_13657);
nor U13991 (N_13991,N_13746,N_13683);
or U13992 (N_13992,N_13715,N_13615);
nand U13993 (N_13993,N_13515,N_13589);
nor U13994 (N_13994,N_13536,N_13692);
nor U13995 (N_13995,N_13566,N_13662);
or U13996 (N_13996,N_13531,N_13588);
or U13997 (N_13997,N_13528,N_13737);
xor U13998 (N_13998,N_13623,N_13701);
or U13999 (N_13999,N_13705,N_13696);
nor U14000 (N_14000,N_13820,N_13761);
and U14001 (N_14001,N_13816,N_13953);
and U14002 (N_14002,N_13838,N_13832);
xnor U14003 (N_14003,N_13946,N_13769);
xnor U14004 (N_14004,N_13985,N_13972);
xor U14005 (N_14005,N_13883,N_13920);
nor U14006 (N_14006,N_13803,N_13767);
nand U14007 (N_14007,N_13963,N_13940);
nand U14008 (N_14008,N_13868,N_13853);
xnor U14009 (N_14009,N_13912,N_13882);
nand U14010 (N_14010,N_13856,N_13751);
and U14011 (N_14011,N_13768,N_13980);
nor U14012 (N_14012,N_13781,N_13861);
or U14013 (N_14013,N_13798,N_13894);
or U14014 (N_14014,N_13927,N_13814);
or U14015 (N_14015,N_13904,N_13784);
nor U14016 (N_14016,N_13961,N_13810);
and U14017 (N_14017,N_13930,N_13959);
nor U14018 (N_14018,N_13867,N_13783);
and U14019 (N_14019,N_13939,N_13759);
nand U14020 (N_14020,N_13976,N_13905);
nand U14021 (N_14021,N_13764,N_13924);
xnor U14022 (N_14022,N_13776,N_13873);
xnor U14023 (N_14023,N_13969,N_13921);
xor U14024 (N_14024,N_13862,N_13922);
or U14025 (N_14025,N_13994,N_13943);
or U14026 (N_14026,N_13808,N_13762);
and U14027 (N_14027,N_13971,N_13931);
xor U14028 (N_14028,N_13944,N_13806);
xor U14029 (N_14029,N_13797,N_13955);
or U14030 (N_14030,N_13859,N_13965);
nand U14031 (N_14031,N_13978,N_13849);
nand U14032 (N_14032,N_13765,N_13854);
nor U14033 (N_14033,N_13909,N_13893);
nand U14034 (N_14034,N_13879,N_13991);
or U14035 (N_14035,N_13997,N_13903);
nor U14036 (N_14036,N_13778,N_13787);
and U14037 (N_14037,N_13844,N_13998);
xor U14038 (N_14038,N_13852,N_13827);
nor U14039 (N_14039,N_13990,N_13851);
nor U14040 (N_14040,N_13910,N_13865);
nand U14041 (N_14041,N_13823,N_13896);
nand U14042 (N_14042,N_13902,N_13796);
nor U14043 (N_14043,N_13753,N_13917);
and U14044 (N_14044,N_13766,N_13949);
or U14045 (N_14045,N_13967,N_13870);
nor U14046 (N_14046,N_13821,N_13822);
nor U14047 (N_14047,N_13885,N_13929);
xor U14048 (N_14048,N_13895,N_13842);
and U14049 (N_14049,N_13906,N_13891);
nor U14050 (N_14050,N_13809,N_13775);
xor U14051 (N_14051,N_13860,N_13750);
and U14052 (N_14052,N_13941,N_13829);
nand U14053 (N_14053,N_13817,N_13892);
nand U14054 (N_14054,N_13938,N_13918);
xor U14055 (N_14055,N_13973,N_13807);
and U14056 (N_14056,N_13913,N_13935);
or U14057 (N_14057,N_13874,N_13984);
nand U14058 (N_14058,N_13995,N_13794);
xnor U14059 (N_14059,N_13779,N_13916);
or U14060 (N_14060,N_13933,N_13900);
xnor U14061 (N_14061,N_13830,N_13754);
nand U14062 (N_14062,N_13804,N_13825);
and U14063 (N_14063,N_13872,N_13780);
or U14064 (N_14064,N_13826,N_13947);
nor U14065 (N_14065,N_13926,N_13818);
and U14066 (N_14066,N_13907,N_13790);
or U14067 (N_14067,N_13974,N_13898);
or U14068 (N_14068,N_13958,N_13878);
or U14069 (N_14069,N_13999,N_13792);
nor U14070 (N_14070,N_13982,N_13773);
and U14071 (N_14071,N_13875,N_13763);
nand U14072 (N_14072,N_13964,N_13815);
and U14073 (N_14073,N_13819,N_13956);
xnor U14074 (N_14074,N_13869,N_13977);
and U14075 (N_14075,N_13756,N_13881);
nand U14076 (N_14076,N_13925,N_13937);
or U14077 (N_14077,N_13805,N_13975);
and U14078 (N_14078,N_13758,N_13855);
nand U14079 (N_14079,N_13850,N_13752);
nor U14080 (N_14080,N_13957,N_13845);
or U14081 (N_14081,N_13770,N_13760);
and U14082 (N_14082,N_13960,N_13880);
xnor U14083 (N_14083,N_13840,N_13934);
xnor U14084 (N_14084,N_13901,N_13877);
or U14085 (N_14085,N_13962,N_13890);
or U14086 (N_14086,N_13908,N_13788);
and U14087 (N_14087,N_13811,N_13847);
or U14088 (N_14088,N_13889,N_13858);
xnor U14089 (N_14089,N_13757,N_13755);
or U14090 (N_14090,N_13897,N_13813);
nor U14091 (N_14091,N_13951,N_13800);
or U14092 (N_14092,N_13911,N_13771);
nand U14093 (N_14093,N_13942,N_13979);
nor U14094 (N_14094,N_13950,N_13836);
or U14095 (N_14095,N_13993,N_13786);
and U14096 (N_14096,N_13782,N_13841);
nand U14097 (N_14097,N_13795,N_13884);
xor U14098 (N_14098,N_13986,N_13923);
nor U14099 (N_14099,N_13802,N_13831);
xnor U14100 (N_14100,N_13772,N_13987);
nand U14101 (N_14101,N_13936,N_13899);
and U14102 (N_14102,N_13888,N_13774);
nand U14103 (N_14103,N_13848,N_13812);
nand U14104 (N_14104,N_13989,N_13945);
xnor U14105 (N_14105,N_13835,N_13843);
nor U14106 (N_14106,N_13833,N_13793);
xnor U14107 (N_14107,N_13863,N_13970);
xor U14108 (N_14108,N_13914,N_13866);
xor U14109 (N_14109,N_13968,N_13992);
nor U14110 (N_14110,N_13948,N_13864);
and U14111 (N_14111,N_13857,N_13983);
and U14112 (N_14112,N_13824,N_13915);
nand U14113 (N_14113,N_13828,N_13846);
nor U14114 (N_14114,N_13919,N_13966);
nor U14115 (N_14115,N_13954,N_13871);
xnor U14116 (N_14116,N_13876,N_13799);
nand U14117 (N_14117,N_13932,N_13887);
and U14118 (N_14118,N_13928,N_13886);
xnor U14119 (N_14119,N_13791,N_13801);
nand U14120 (N_14120,N_13785,N_13981);
nor U14121 (N_14121,N_13834,N_13777);
or U14122 (N_14122,N_13837,N_13839);
and U14123 (N_14123,N_13789,N_13988);
and U14124 (N_14124,N_13996,N_13952);
nor U14125 (N_14125,N_13810,N_13762);
xnor U14126 (N_14126,N_13885,N_13817);
nor U14127 (N_14127,N_13906,N_13956);
nand U14128 (N_14128,N_13791,N_13769);
and U14129 (N_14129,N_13889,N_13815);
xor U14130 (N_14130,N_13854,N_13928);
and U14131 (N_14131,N_13771,N_13789);
nor U14132 (N_14132,N_13814,N_13951);
nor U14133 (N_14133,N_13846,N_13804);
nor U14134 (N_14134,N_13937,N_13753);
or U14135 (N_14135,N_13869,N_13966);
xor U14136 (N_14136,N_13945,N_13914);
nand U14137 (N_14137,N_13951,N_13804);
nand U14138 (N_14138,N_13891,N_13858);
nand U14139 (N_14139,N_13892,N_13779);
and U14140 (N_14140,N_13958,N_13857);
or U14141 (N_14141,N_13765,N_13826);
nor U14142 (N_14142,N_13881,N_13848);
nand U14143 (N_14143,N_13928,N_13750);
nor U14144 (N_14144,N_13839,N_13761);
nand U14145 (N_14145,N_13982,N_13894);
and U14146 (N_14146,N_13996,N_13805);
nand U14147 (N_14147,N_13887,N_13960);
and U14148 (N_14148,N_13972,N_13945);
xor U14149 (N_14149,N_13844,N_13785);
or U14150 (N_14150,N_13816,N_13957);
or U14151 (N_14151,N_13841,N_13931);
and U14152 (N_14152,N_13828,N_13942);
and U14153 (N_14153,N_13780,N_13834);
nor U14154 (N_14154,N_13857,N_13901);
or U14155 (N_14155,N_13764,N_13762);
nand U14156 (N_14156,N_13963,N_13783);
and U14157 (N_14157,N_13875,N_13780);
or U14158 (N_14158,N_13942,N_13998);
or U14159 (N_14159,N_13791,N_13929);
and U14160 (N_14160,N_13807,N_13884);
nor U14161 (N_14161,N_13809,N_13918);
nor U14162 (N_14162,N_13799,N_13878);
xnor U14163 (N_14163,N_13850,N_13861);
nor U14164 (N_14164,N_13925,N_13786);
nor U14165 (N_14165,N_13841,N_13828);
nand U14166 (N_14166,N_13789,N_13857);
xor U14167 (N_14167,N_13916,N_13841);
nand U14168 (N_14168,N_13856,N_13970);
nor U14169 (N_14169,N_13960,N_13943);
xnor U14170 (N_14170,N_13767,N_13906);
nand U14171 (N_14171,N_13841,N_13781);
and U14172 (N_14172,N_13809,N_13911);
nand U14173 (N_14173,N_13979,N_13971);
and U14174 (N_14174,N_13843,N_13836);
nand U14175 (N_14175,N_13984,N_13885);
and U14176 (N_14176,N_13963,N_13816);
nor U14177 (N_14177,N_13912,N_13781);
and U14178 (N_14178,N_13974,N_13931);
or U14179 (N_14179,N_13930,N_13866);
nor U14180 (N_14180,N_13938,N_13845);
nor U14181 (N_14181,N_13773,N_13955);
xnor U14182 (N_14182,N_13863,N_13866);
xnor U14183 (N_14183,N_13772,N_13770);
nor U14184 (N_14184,N_13783,N_13978);
nor U14185 (N_14185,N_13755,N_13854);
nand U14186 (N_14186,N_13819,N_13894);
or U14187 (N_14187,N_13980,N_13877);
nor U14188 (N_14188,N_13963,N_13791);
xnor U14189 (N_14189,N_13768,N_13952);
nand U14190 (N_14190,N_13931,N_13938);
nand U14191 (N_14191,N_13825,N_13882);
nand U14192 (N_14192,N_13826,N_13975);
and U14193 (N_14193,N_13999,N_13773);
and U14194 (N_14194,N_13787,N_13869);
nand U14195 (N_14195,N_13764,N_13974);
and U14196 (N_14196,N_13757,N_13880);
nor U14197 (N_14197,N_13750,N_13953);
or U14198 (N_14198,N_13775,N_13850);
nand U14199 (N_14199,N_13997,N_13967);
nor U14200 (N_14200,N_13936,N_13930);
xor U14201 (N_14201,N_13837,N_13811);
and U14202 (N_14202,N_13841,N_13844);
and U14203 (N_14203,N_13992,N_13771);
and U14204 (N_14204,N_13900,N_13915);
nor U14205 (N_14205,N_13791,N_13771);
nor U14206 (N_14206,N_13993,N_13961);
nor U14207 (N_14207,N_13774,N_13799);
nand U14208 (N_14208,N_13886,N_13768);
and U14209 (N_14209,N_13985,N_13952);
or U14210 (N_14210,N_13794,N_13886);
xor U14211 (N_14211,N_13904,N_13763);
nor U14212 (N_14212,N_13786,N_13959);
xor U14213 (N_14213,N_13867,N_13897);
nor U14214 (N_14214,N_13943,N_13853);
xnor U14215 (N_14215,N_13934,N_13831);
nor U14216 (N_14216,N_13874,N_13928);
xnor U14217 (N_14217,N_13983,N_13929);
and U14218 (N_14218,N_13794,N_13927);
xor U14219 (N_14219,N_13824,N_13846);
and U14220 (N_14220,N_13843,N_13834);
xnor U14221 (N_14221,N_13779,N_13799);
nand U14222 (N_14222,N_13821,N_13948);
nand U14223 (N_14223,N_13990,N_13906);
nor U14224 (N_14224,N_13874,N_13978);
xnor U14225 (N_14225,N_13964,N_13945);
xnor U14226 (N_14226,N_13852,N_13953);
nand U14227 (N_14227,N_13960,N_13781);
or U14228 (N_14228,N_13839,N_13961);
nor U14229 (N_14229,N_13976,N_13806);
and U14230 (N_14230,N_13756,N_13951);
and U14231 (N_14231,N_13848,N_13865);
or U14232 (N_14232,N_13807,N_13882);
or U14233 (N_14233,N_13934,N_13855);
nand U14234 (N_14234,N_13840,N_13962);
and U14235 (N_14235,N_13779,N_13951);
xor U14236 (N_14236,N_13802,N_13852);
nor U14237 (N_14237,N_13846,N_13922);
and U14238 (N_14238,N_13983,N_13806);
xnor U14239 (N_14239,N_13941,N_13981);
or U14240 (N_14240,N_13809,N_13858);
or U14241 (N_14241,N_13854,N_13919);
or U14242 (N_14242,N_13787,N_13777);
xnor U14243 (N_14243,N_13931,N_13864);
xnor U14244 (N_14244,N_13956,N_13750);
nor U14245 (N_14245,N_13938,N_13960);
xnor U14246 (N_14246,N_13900,N_13957);
xor U14247 (N_14247,N_13888,N_13968);
and U14248 (N_14248,N_13826,N_13875);
xor U14249 (N_14249,N_13805,N_13894);
xnor U14250 (N_14250,N_14049,N_14048);
nor U14251 (N_14251,N_14232,N_14115);
xor U14252 (N_14252,N_14228,N_14112);
and U14253 (N_14253,N_14052,N_14069);
nand U14254 (N_14254,N_14153,N_14167);
nand U14255 (N_14255,N_14160,N_14072);
or U14256 (N_14256,N_14059,N_14119);
nor U14257 (N_14257,N_14187,N_14008);
and U14258 (N_14258,N_14233,N_14066);
or U14259 (N_14259,N_14138,N_14158);
nor U14260 (N_14260,N_14230,N_14067);
xor U14261 (N_14261,N_14116,N_14007);
nor U14262 (N_14262,N_14142,N_14204);
nor U14263 (N_14263,N_14225,N_14223);
xnor U14264 (N_14264,N_14071,N_14041);
or U14265 (N_14265,N_14010,N_14015);
and U14266 (N_14266,N_14194,N_14175);
nor U14267 (N_14267,N_14002,N_14079);
nand U14268 (N_14268,N_14099,N_14201);
or U14269 (N_14269,N_14030,N_14000);
nand U14270 (N_14270,N_14149,N_14062);
nand U14271 (N_14271,N_14024,N_14168);
xnor U14272 (N_14272,N_14109,N_14156);
nand U14273 (N_14273,N_14060,N_14183);
or U14274 (N_14274,N_14128,N_14065);
nor U14275 (N_14275,N_14198,N_14213);
and U14276 (N_14276,N_14018,N_14245);
nand U14277 (N_14277,N_14005,N_14141);
or U14278 (N_14278,N_14101,N_14053);
or U14279 (N_14279,N_14044,N_14098);
xnor U14280 (N_14280,N_14016,N_14170);
and U14281 (N_14281,N_14061,N_14218);
and U14282 (N_14282,N_14100,N_14102);
nor U14283 (N_14283,N_14165,N_14083);
nand U14284 (N_14284,N_14082,N_14241);
nand U14285 (N_14285,N_14246,N_14191);
and U14286 (N_14286,N_14238,N_14051);
and U14287 (N_14287,N_14169,N_14211);
or U14288 (N_14288,N_14186,N_14039);
or U14289 (N_14289,N_14074,N_14023);
nor U14290 (N_14290,N_14017,N_14031);
xor U14291 (N_14291,N_14013,N_14038);
nor U14292 (N_14292,N_14094,N_14093);
and U14293 (N_14293,N_14081,N_14162);
and U14294 (N_14294,N_14210,N_14003);
nand U14295 (N_14295,N_14085,N_14215);
nand U14296 (N_14296,N_14147,N_14047);
or U14297 (N_14297,N_14011,N_14027);
or U14298 (N_14298,N_14064,N_14086);
nand U14299 (N_14299,N_14208,N_14090);
or U14300 (N_14300,N_14217,N_14173);
or U14301 (N_14301,N_14224,N_14164);
and U14302 (N_14302,N_14172,N_14136);
nand U14303 (N_14303,N_14155,N_14125);
xor U14304 (N_14304,N_14229,N_14212);
or U14305 (N_14305,N_14133,N_14236);
and U14306 (N_14306,N_14121,N_14103);
nand U14307 (N_14307,N_14248,N_14058);
xor U14308 (N_14308,N_14050,N_14097);
and U14309 (N_14309,N_14028,N_14239);
or U14310 (N_14310,N_14089,N_14104);
xnor U14311 (N_14311,N_14012,N_14056);
nand U14312 (N_14312,N_14130,N_14219);
nand U14313 (N_14313,N_14077,N_14095);
and U14314 (N_14314,N_14159,N_14148);
nand U14315 (N_14315,N_14004,N_14196);
xnor U14316 (N_14316,N_14057,N_14195);
and U14317 (N_14317,N_14131,N_14105);
and U14318 (N_14318,N_14087,N_14190);
nand U14319 (N_14319,N_14139,N_14197);
and U14320 (N_14320,N_14111,N_14075);
nor U14321 (N_14321,N_14040,N_14009);
xor U14322 (N_14322,N_14084,N_14227);
nand U14323 (N_14323,N_14129,N_14078);
nor U14324 (N_14324,N_14035,N_14042);
nand U14325 (N_14325,N_14171,N_14014);
nor U14326 (N_14326,N_14037,N_14118);
and U14327 (N_14327,N_14214,N_14157);
nor U14328 (N_14328,N_14123,N_14140);
xor U14329 (N_14329,N_14221,N_14120);
xor U14330 (N_14330,N_14126,N_14179);
nand U14331 (N_14331,N_14143,N_14006);
and U14332 (N_14332,N_14240,N_14184);
nand U14333 (N_14333,N_14154,N_14046);
nor U14334 (N_14334,N_14045,N_14091);
and U14335 (N_14335,N_14193,N_14205);
xor U14336 (N_14336,N_14033,N_14114);
nand U14337 (N_14337,N_14163,N_14203);
nor U14338 (N_14338,N_14063,N_14055);
and U14339 (N_14339,N_14178,N_14202);
nand U14340 (N_14340,N_14073,N_14092);
nand U14341 (N_14341,N_14088,N_14200);
nand U14342 (N_14342,N_14242,N_14247);
and U14343 (N_14343,N_14001,N_14220);
nand U14344 (N_14344,N_14110,N_14080);
and U14345 (N_14345,N_14036,N_14113);
xnor U14346 (N_14346,N_14032,N_14132);
and U14347 (N_14347,N_14150,N_14207);
xnor U14348 (N_14348,N_14068,N_14026);
or U14349 (N_14349,N_14152,N_14209);
nor U14350 (N_14350,N_14182,N_14234);
nor U14351 (N_14351,N_14025,N_14226);
nor U14352 (N_14352,N_14166,N_14107);
xnor U14353 (N_14353,N_14244,N_14022);
nand U14354 (N_14354,N_14176,N_14124);
and U14355 (N_14355,N_14043,N_14145);
or U14356 (N_14356,N_14134,N_14237);
nor U14357 (N_14357,N_14181,N_14146);
nand U14358 (N_14358,N_14021,N_14188);
nand U14359 (N_14359,N_14020,N_14216);
nand U14360 (N_14360,N_14127,N_14135);
or U14361 (N_14361,N_14144,N_14019);
nand U14362 (N_14362,N_14137,N_14249);
nand U14363 (N_14363,N_14222,N_14070);
or U14364 (N_14364,N_14029,N_14185);
nor U14365 (N_14365,N_14122,N_14106);
nor U14366 (N_14366,N_14161,N_14174);
xnor U14367 (N_14367,N_14054,N_14192);
xor U14368 (N_14368,N_14206,N_14034);
or U14369 (N_14369,N_14177,N_14108);
or U14370 (N_14370,N_14096,N_14199);
or U14371 (N_14371,N_14235,N_14243);
nand U14372 (N_14372,N_14076,N_14180);
or U14373 (N_14373,N_14117,N_14231);
or U14374 (N_14374,N_14189,N_14151);
nor U14375 (N_14375,N_14109,N_14052);
nor U14376 (N_14376,N_14188,N_14057);
or U14377 (N_14377,N_14015,N_14086);
and U14378 (N_14378,N_14018,N_14011);
xnor U14379 (N_14379,N_14067,N_14228);
nor U14380 (N_14380,N_14059,N_14204);
and U14381 (N_14381,N_14199,N_14217);
nand U14382 (N_14382,N_14089,N_14065);
and U14383 (N_14383,N_14055,N_14180);
and U14384 (N_14384,N_14040,N_14010);
or U14385 (N_14385,N_14070,N_14145);
and U14386 (N_14386,N_14158,N_14190);
nand U14387 (N_14387,N_14151,N_14002);
and U14388 (N_14388,N_14054,N_14188);
and U14389 (N_14389,N_14241,N_14004);
or U14390 (N_14390,N_14029,N_14226);
nor U14391 (N_14391,N_14196,N_14132);
nor U14392 (N_14392,N_14060,N_14017);
nor U14393 (N_14393,N_14213,N_14114);
xor U14394 (N_14394,N_14049,N_14238);
or U14395 (N_14395,N_14017,N_14226);
or U14396 (N_14396,N_14243,N_14057);
nor U14397 (N_14397,N_14018,N_14067);
and U14398 (N_14398,N_14166,N_14148);
and U14399 (N_14399,N_14172,N_14237);
nor U14400 (N_14400,N_14170,N_14118);
nor U14401 (N_14401,N_14011,N_14110);
xor U14402 (N_14402,N_14193,N_14011);
and U14403 (N_14403,N_14041,N_14166);
and U14404 (N_14404,N_14225,N_14246);
and U14405 (N_14405,N_14238,N_14151);
or U14406 (N_14406,N_14247,N_14034);
or U14407 (N_14407,N_14245,N_14184);
or U14408 (N_14408,N_14133,N_14235);
nor U14409 (N_14409,N_14152,N_14178);
xnor U14410 (N_14410,N_14213,N_14130);
and U14411 (N_14411,N_14058,N_14243);
or U14412 (N_14412,N_14135,N_14164);
xor U14413 (N_14413,N_14052,N_14018);
nor U14414 (N_14414,N_14093,N_14012);
or U14415 (N_14415,N_14249,N_14165);
xor U14416 (N_14416,N_14162,N_14221);
and U14417 (N_14417,N_14064,N_14114);
xnor U14418 (N_14418,N_14202,N_14128);
nor U14419 (N_14419,N_14071,N_14122);
nand U14420 (N_14420,N_14038,N_14223);
xor U14421 (N_14421,N_14203,N_14028);
and U14422 (N_14422,N_14233,N_14188);
xor U14423 (N_14423,N_14237,N_14217);
nand U14424 (N_14424,N_14071,N_14234);
and U14425 (N_14425,N_14010,N_14082);
and U14426 (N_14426,N_14134,N_14087);
nor U14427 (N_14427,N_14179,N_14017);
nand U14428 (N_14428,N_14163,N_14226);
xor U14429 (N_14429,N_14156,N_14060);
and U14430 (N_14430,N_14097,N_14141);
or U14431 (N_14431,N_14084,N_14056);
xor U14432 (N_14432,N_14004,N_14003);
xnor U14433 (N_14433,N_14037,N_14140);
or U14434 (N_14434,N_14246,N_14243);
and U14435 (N_14435,N_14144,N_14186);
nand U14436 (N_14436,N_14227,N_14130);
or U14437 (N_14437,N_14215,N_14200);
nand U14438 (N_14438,N_14178,N_14095);
nor U14439 (N_14439,N_14014,N_14080);
and U14440 (N_14440,N_14124,N_14214);
xor U14441 (N_14441,N_14105,N_14021);
xnor U14442 (N_14442,N_14126,N_14237);
xor U14443 (N_14443,N_14158,N_14111);
and U14444 (N_14444,N_14197,N_14244);
or U14445 (N_14445,N_14145,N_14231);
or U14446 (N_14446,N_14019,N_14210);
nand U14447 (N_14447,N_14058,N_14108);
or U14448 (N_14448,N_14048,N_14056);
and U14449 (N_14449,N_14133,N_14076);
and U14450 (N_14450,N_14226,N_14164);
or U14451 (N_14451,N_14113,N_14166);
and U14452 (N_14452,N_14047,N_14092);
nand U14453 (N_14453,N_14230,N_14018);
and U14454 (N_14454,N_14215,N_14197);
or U14455 (N_14455,N_14242,N_14097);
nor U14456 (N_14456,N_14046,N_14008);
and U14457 (N_14457,N_14194,N_14230);
nor U14458 (N_14458,N_14171,N_14237);
nor U14459 (N_14459,N_14082,N_14027);
nand U14460 (N_14460,N_14091,N_14207);
and U14461 (N_14461,N_14242,N_14156);
and U14462 (N_14462,N_14054,N_14088);
xnor U14463 (N_14463,N_14056,N_14176);
nand U14464 (N_14464,N_14221,N_14151);
or U14465 (N_14465,N_14162,N_14145);
and U14466 (N_14466,N_14117,N_14130);
or U14467 (N_14467,N_14036,N_14233);
nor U14468 (N_14468,N_14145,N_14236);
nand U14469 (N_14469,N_14160,N_14091);
or U14470 (N_14470,N_14065,N_14071);
xnor U14471 (N_14471,N_14169,N_14244);
or U14472 (N_14472,N_14239,N_14175);
xnor U14473 (N_14473,N_14237,N_14210);
xor U14474 (N_14474,N_14030,N_14119);
and U14475 (N_14475,N_14041,N_14057);
or U14476 (N_14476,N_14236,N_14142);
xor U14477 (N_14477,N_14073,N_14135);
nand U14478 (N_14478,N_14119,N_14140);
and U14479 (N_14479,N_14109,N_14161);
nand U14480 (N_14480,N_14057,N_14232);
nand U14481 (N_14481,N_14140,N_14224);
or U14482 (N_14482,N_14193,N_14243);
xor U14483 (N_14483,N_14166,N_14228);
nor U14484 (N_14484,N_14065,N_14139);
nor U14485 (N_14485,N_14013,N_14083);
or U14486 (N_14486,N_14065,N_14181);
nand U14487 (N_14487,N_14047,N_14145);
nor U14488 (N_14488,N_14065,N_14067);
nand U14489 (N_14489,N_14078,N_14116);
nand U14490 (N_14490,N_14176,N_14242);
or U14491 (N_14491,N_14014,N_14087);
and U14492 (N_14492,N_14105,N_14210);
nor U14493 (N_14493,N_14004,N_14087);
nand U14494 (N_14494,N_14229,N_14132);
and U14495 (N_14495,N_14035,N_14189);
nand U14496 (N_14496,N_14226,N_14050);
xor U14497 (N_14497,N_14049,N_14009);
nor U14498 (N_14498,N_14218,N_14161);
nor U14499 (N_14499,N_14172,N_14226);
nand U14500 (N_14500,N_14458,N_14395);
and U14501 (N_14501,N_14485,N_14368);
and U14502 (N_14502,N_14382,N_14445);
nor U14503 (N_14503,N_14479,N_14302);
and U14504 (N_14504,N_14491,N_14356);
nand U14505 (N_14505,N_14380,N_14406);
and U14506 (N_14506,N_14296,N_14473);
nand U14507 (N_14507,N_14437,N_14285);
nand U14508 (N_14508,N_14439,N_14456);
and U14509 (N_14509,N_14346,N_14374);
or U14510 (N_14510,N_14323,N_14405);
nor U14511 (N_14511,N_14492,N_14418);
and U14512 (N_14512,N_14328,N_14274);
xor U14513 (N_14513,N_14273,N_14284);
xnor U14514 (N_14514,N_14367,N_14304);
xor U14515 (N_14515,N_14394,N_14385);
nand U14516 (N_14516,N_14480,N_14411);
nor U14517 (N_14517,N_14435,N_14313);
nor U14518 (N_14518,N_14287,N_14468);
and U14519 (N_14519,N_14431,N_14444);
nor U14520 (N_14520,N_14258,N_14353);
nor U14521 (N_14521,N_14282,N_14376);
or U14522 (N_14522,N_14389,N_14465);
nor U14523 (N_14523,N_14331,N_14317);
or U14524 (N_14524,N_14446,N_14404);
and U14525 (N_14525,N_14267,N_14416);
or U14526 (N_14526,N_14292,N_14270);
xnor U14527 (N_14527,N_14255,N_14291);
xnor U14528 (N_14528,N_14316,N_14470);
nor U14529 (N_14529,N_14257,N_14459);
nand U14530 (N_14530,N_14432,N_14361);
xnor U14531 (N_14531,N_14345,N_14472);
or U14532 (N_14532,N_14303,N_14461);
and U14533 (N_14533,N_14397,N_14334);
xor U14534 (N_14534,N_14253,N_14484);
or U14535 (N_14535,N_14378,N_14436);
or U14536 (N_14536,N_14275,N_14424);
xor U14537 (N_14537,N_14454,N_14381);
or U14538 (N_14538,N_14386,N_14280);
nor U14539 (N_14539,N_14347,N_14490);
nor U14540 (N_14540,N_14268,N_14339);
nand U14541 (N_14541,N_14442,N_14261);
nand U14542 (N_14542,N_14494,N_14354);
nand U14543 (N_14543,N_14363,N_14489);
nor U14544 (N_14544,N_14350,N_14362);
xnor U14545 (N_14545,N_14466,N_14384);
and U14546 (N_14546,N_14355,N_14340);
nor U14547 (N_14547,N_14252,N_14392);
nor U14548 (N_14548,N_14370,N_14495);
and U14549 (N_14549,N_14441,N_14281);
xnor U14550 (N_14550,N_14409,N_14271);
and U14551 (N_14551,N_14452,N_14430);
nor U14552 (N_14552,N_14419,N_14414);
or U14553 (N_14553,N_14289,N_14415);
or U14554 (N_14554,N_14369,N_14398);
xor U14555 (N_14555,N_14401,N_14259);
xnor U14556 (N_14556,N_14309,N_14410);
xor U14557 (N_14557,N_14457,N_14278);
nand U14558 (N_14558,N_14402,N_14462);
xnor U14559 (N_14559,N_14360,N_14262);
or U14560 (N_14560,N_14320,N_14417);
or U14561 (N_14561,N_14447,N_14412);
nor U14562 (N_14562,N_14375,N_14455);
or U14563 (N_14563,N_14383,N_14254);
nor U14564 (N_14564,N_14326,N_14312);
xor U14565 (N_14565,N_14464,N_14348);
nor U14566 (N_14566,N_14475,N_14276);
xor U14567 (N_14567,N_14372,N_14335);
nand U14568 (N_14568,N_14493,N_14482);
and U14569 (N_14569,N_14336,N_14449);
nand U14570 (N_14570,N_14467,N_14498);
nor U14571 (N_14571,N_14358,N_14342);
nor U14572 (N_14572,N_14440,N_14427);
and U14573 (N_14573,N_14433,N_14425);
or U14574 (N_14574,N_14264,N_14423);
nand U14575 (N_14575,N_14443,N_14306);
xnor U14576 (N_14576,N_14251,N_14408);
xor U14577 (N_14577,N_14448,N_14298);
and U14578 (N_14578,N_14365,N_14438);
nor U14579 (N_14579,N_14341,N_14390);
nand U14580 (N_14580,N_14277,N_14332);
and U14581 (N_14581,N_14400,N_14453);
xnor U14582 (N_14582,N_14393,N_14329);
nand U14583 (N_14583,N_14325,N_14283);
and U14584 (N_14584,N_14359,N_14481);
or U14585 (N_14585,N_14295,N_14499);
xnor U14586 (N_14586,N_14256,N_14308);
nor U14587 (N_14587,N_14450,N_14290);
and U14588 (N_14588,N_14310,N_14429);
xor U14589 (N_14589,N_14265,N_14352);
nor U14590 (N_14590,N_14266,N_14351);
nand U14591 (N_14591,N_14421,N_14388);
xnor U14592 (N_14592,N_14324,N_14319);
nand U14593 (N_14593,N_14269,N_14338);
nor U14594 (N_14594,N_14428,N_14333);
nor U14595 (N_14595,N_14377,N_14311);
nand U14596 (N_14596,N_14396,N_14272);
xor U14597 (N_14597,N_14318,N_14260);
or U14598 (N_14598,N_14297,N_14460);
nand U14599 (N_14599,N_14330,N_14477);
nand U14600 (N_14600,N_14294,N_14315);
xor U14601 (N_14601,N_14496,N_14349);
nor U14602 (N_14602,N_14486,N_14366);
xnor U14603 (N_14603,N_14391,N_14305);
xor U14604 (N_14604,N_14407,N_14288);
nand U14605 (N_14605,N_14344,N_14343);
xnor U14606 (N_14606,N_14426,N_14488);
nand U14607 (N_14607,N_14371,N_14293);
nand U14608 (N_14608,N_14422,N_14286);
xor U14609 (N_14609,N_14497,N_14463);
nor U14610 (N_14610,N_14483,N_14471);
nor U14611 (N_14611,N_14476,N_14403);
and U14612 (N_14612,N_14300,N_14322);
nor U14613 (N_14613,N_14469,N_14413);
nor U14614 (N_14614,N_14420,N_14379);
and U14615 (N_14615,N_14399,N_14487);
or U14616 (N_14616,N_14357,N_14279);
nor U14617 (N_14617,N_14263,N_14478);
or U14618 (N_14618,N_14364,N_14337);
nor U14619 (N_14619,N_14307,N_14321);
nor U14620 (N_14620,N_14314,N_14387);
and U14621 (N_14621,N_14327,N_14373);
xnor U14622 (N_14622,N_14474,N_14434);
nor U14623 (N_14623,N_14299,N_14301);
or U14624 (N_14624,N_14250,N_14451);
and U14625 (N_14625,N_14465,N_14293);
xnor U14626 (N_14626,N_14428,N_14455);
xnor U14627 (N_14627,N_14405,N_14410);
xnor U14628 (N_14628,N_14417,N_14267);
xor U14629 (N_14629,N_14396,N_14320);
nor U14630 (N_14630,N_14485,N_14370);
nor U14631 (N_14631,N_14318,N_14390);
nor U14632 (N_14632,N_14387,N_14363);
nor U14633 (N_14633,N_14358,N_14498);
nor U14634 (N_14634,N_14321,N_14328);
and U14635 (N_14635,N_14388,N_14466);
xor U14636 (N_14636,N_14449,N_14418);
or U14637 (N_14637,N_14310,N_14341);
nand U14638 (N_14638,N_14333,N_14438);
xnor U14639 (N_14639,N_14436,N_14498);
or U14640 (N_14640,N_14441,N_14373);
nand U14641 (N_14641,N_14335,N_14259);
nand U14642 (N_14642,N_14382,N_14263);
nand U14643 (N_14643,N_14437,N_14387);
and U14644 (N_14644,N_14463,N_14382);
nor U14645 (N_14645,N_14489,N_14264);
xor U14646 (N_14646,N_14478,N_14494);
nand U14647 (N_14647,N_14253,N_14427);
nor U14648 (N_14648,N_14441,N_14493);
xor U14649 (N_14649,N_14430,N_14392);
nor U14650 (N_14650,N_14272,N_14325);
nand U14651 (N_14651,N_14480,N_14305);
or U14652 (N_14652,N_14330,N_14344);
or U14653 (N_14653,N_14366,N_14278);
and U14654 (N_14654,N_14434,N_14263);
and U14655 (N_14655,N_14490,N_14265);
and U14656 (N_14656,N_14493,N_14409);
nand U14657 (N_14657,N_14455,N_14454);
and U14658 (N_14658,N_14340,N_14330);
and U14659 (N_14659,N_14420,N_14402);
xnor U14660 (N_14660,N_14363,N_14428);
nand U14661 (N_14661,N_14304,N_14347);
xnor U14662 (N_14662,N_14282,N_14498);
nor U14663 (N_14663,N_14381,N_14425);
and U14664 (N_14664,N_14267,N_14292);
xnor U14665 (N_14665,N_14404,N_14314);
or U14666 (N_14666,N_14254,N_14293);
nand U14667 (N_14667,N_14324,N_14337);
nand U14668 (N_14668,N_14445,N_14316);
and U14669 (N_14669,N_14463,N_14271);
and U14670 (N_14670,N_14301,N_14474);
nor U14671 (N_14671,N_14269,N_14374);
nor U14672 (N_14672,N_14398,N_14496);
or U14673 (N_14673,N_14455,N_14350);
xor U14674 (N_14674,N_14487,N_14304);
nand U14675 (N_14675,N_14385,N_14281);
and U14676 (N_14676,N_14460,N_14395);
xnor U14677 (N_14677,N_14367,N_14427);
and U14678 (N_14678,N_14366,N_14356);
or U14679 (N_14679,N_14392,N_14298);
or U14680 (N_14680,N_14490,N_14337);
nand U14681 (N_14681,N_14423,N_14480);
nand U14682 (N_14682,N_14346,N_14415);
nor U14683 (N_14683,N_14312,N_14447);
or U14684 (N_14684,N_14355,N_14433);
nand U14685 (N_14685,N_14368,N_14401);
and U14686 (N_14686,N_14394,N_14424);
and U14687 (N_14687,N_14444,N_14478);
nor U14688 (N_14688,N_14253,N_14379);
or U14689 (N_14689,N_14340,N_14314);
nor U14690 (N_14690,N_14470,N_14459);
nand U14691 (N_14691,N_14396,N_14476);
nor U14692 (N_14692,N_14337,N_14400);
and U14693 (N_14693,N_14398,N_14393);
nor U14694 (N_14694,N_14433,N_14478);
nand U14695 (N_14695,N_14274,N_14259);
and U14696 (N_14696,N_14395,N_14427);
xor U14697 (N_14697,N_14468,N_14483);
or U14698 (N_14698,N_14401,N_14406);
and U14699 (N_14699,N_14394,N_14255);
and U14700 (N_14700,N_14251,N_14327);
or U14701 (N_14701,N_14431,N_14477);
xnor U14702 (N_14702,N_14275,N_14347);
or U14703 (N_14703,N_14285,N_14456);
nor U14704 (N_14704,N_14489,N_14384);
xnor U14705 (N_14705,N_14361,N_14469);
or U14706 (N_14706,N_14264,N_14263);
nand U14707 (N_14707,N_14417,N_14336);
nor U14708 (N_14708,N_14322,N_14269);
nor U14709 (N_14709,N_14477,N_14460);
or U14710 (N_14710,N_14412,N_14367);
or U14711 (N_14711,N_14487,N_14403);
and U14712 (N_14712,N_14257,N_14340);
and U14713 (N_14713,N_14436,N_14298);
xnor U14714 (N_14714,N_14295,N_14340);
nand U14715 (N_14715,N_14431,N_14322);
xor U14716 (N_14716,N_14484,N_14352);
xnor U14717 (N_14717,N_14378,N_14291);
xor U14718 (N_14718,N_14323,N_14425);
nand U14719 (N_14719,N_14431,N_14493);
and U14720 (N_14720,N_14333,N_14271);
nand U14721 (N_14721,N_14483,N_14462);
nand U14722 (N_14722,N_14329,N_14340);
and U14723 (N_14723,N_14250,N_14459);
or U14724 (N_14724,N_14466,N_14360);
and U14725 (N_14725,N_14495,N_14288);
or U14726 (N_14726,N_14498,N_14313);
and U14727 (N_14727,N_14323,N_14404);
xor U14728 (N_14728,N_14328,N_14466);
and U14729 (N_14729,N_14441,N_14443);
nand U14730 (N_14730,N_14264,N_14480);
nor U14731 (N_14731,N_14317,N_14375);
or U14732 (N_14732,N_14439,N_14263);
and U14733 (N_14733,N_14358,N_14316);
or U14734 (N_14734,N_14399,N_14465);
xnor U14735 (N_14735,N_14302,N_14462);
nand U14736 (N_14736,N_14297,N_14495);
xnor U14737 (N_14737,N_14351,N_14462);
nor U14738 (N_14738,N_14414,N_14287);
nand U14739 (N_14739,N_14294,N_14443);
xor U14740 (N_14740,N_14389,N_14410);
nand U14741 (N_14741,N_14440,N_14410);
or U14742 (N_14742,N_14355,N_14414);
nand U14743 (N_14743,N_14266,N_14278);
nor U14744 (N_14744,N_14455,N_14422);
or U14745 (N_14745,N_14327,N_14467);
nand U14746 (N_14746,N_14420,N_14475);
and U14747 (N_14747,N_14266,N_14489);
nand U14748 (N_14748,N_14475,N_14295);
xnor U14749 (N_14749,N_14332,N_14250);
and U14750 (N_14750,N_14569,N_14556);
nand U14751 (N_14751,N_14606,N_14715);
nor U14752 (N_14752,N_14589,N_14561);
and U14753 (N_14753,N_14597,N_14554);
nand U14754 (N_14754,N_14619,N_14633);
nand U14755 (N_14755,N_14696,N_14737);
nand U14756 (N_14756,N_14601,N_14711);
or U14757 (N_14757,N_14681,N_14721);
nand U14758 (N_14758,N_14677,N_14583);
nand U14759 (N_14759,N_14519,N_14625);
nor U14760 (N_14760,N_14725,N_14507);
nor U14761 (N_14761,N_14615,N_14623);
and U14762 (N_14762,N_14684,N_14523);
nand U14763 (N_14763,N_14539,N_14707);
nand U14764 (N_14764,N_14632,N_14511);
xnor U14765 (N_14765,N_14645,N_14697);
or U14766 (N_14766,N_14610,N_14567);
and U14767 (N_14767,N_14718,N_14660);
or U14768 (N_14768,N_14653,N_14662);
and U14769 (N_14769,N_14515,N_14525);
nand U14770 (N_14770,N_14592,N_14622);
xor U14771 (N_14771,N_14573,N_14527);
nand U14772 (N_14772,N_14686,N_14731);
xnor U14773 (N_14773,N_14643,N_14650);
nor U14774 (N_14774,N_14698,N_14616);
nand U14775 (N_14775,N_14548,N_14655);
nor U14776 (N_14776,N_14690,N_14739);
or U14777 (N_14777,N_14602,N_14713);
nand U14778 (N_14778,N_14672,N_14605);
nor U14779 (N_14779,N_14661,N_14505);
nand U14780 (N_14780,N_14745,N_14692);
xor U14781 (N_14781,N_14678,N_14641);
xor U14782 (N_14782,N_14566,N_14716);
xnor U14783 (N_14783,N_14666,N_14652);
nand U14784 (N_14784,N_14517,N_14720);
or U14785 (N_14785,N_14549,N_14559);
xor U14786 (N_14786,N_14552,N_14571);
nor U14787 (N_14787,N_14538,N_14603);
nor U14788 (N_14788,N_14504,N_14740);
or U14789 (N_14789,N_14636,N_14607);
and U14790 (N_14790,N_14732,N_14639);
nor U14791 (N_14791,N_14679,N_14565);
and U14792 (N_14792,N_14594,N_14516);
or U14793 (N_14793,N_14506,N_14503);
nor U14794 (N_14794,N_14695,N_14669);
or U14795 (N_14795,N_14500,N_14544);
and U14796 (N_14796,N_14744,N_14621);
and U14797 (N_14797,N_14665,N_14614);
and U14798 (N_14798,N_14532,N_14522);
or U14799 (N_14799,N_14746,N_14629);
nor U14800 (N_14800,N_14627,N_14749);
nor U14801 (N_14801,N_14723,N_14689);
xnor U14802 (N_14802,N_14591,N_14572);
and U14803 (N_14803,N_14575,N_14588);
or U14804 (N_14804,N_14590,N_14545);
or U14805 (N_14805,N_14617,N_14620);
or U14806 (N_14806,N_14685,N_14694);
or U14807 (N_14807,N_14743,N_14709);
nor U14808 (N_14808,N_14509,N_14563);
nor U14809 (N_14809,N_14675,N_14520);
or U14810 (N_14810,N_14624,N_14700);
xnor U14811 (N_14811,N_14705,N_14608);
xnor U14812 (N_14812,N_14541,N_14670);
and U14813 (N_14813,N_14646,N_14609);
xor U14814 (N_14814,N_14564,N_14706);
xnor U14815 (N_14815,N_14726,N_14659);
xnor U14816 (N_14816,N_14668,N_14654);
nand U14817 (N_14817,N_14699,N_14693);
or U14818 (N_14818,N_14687,N_14562);
and U14819 (N_14819,N_14635,N_14585);
and U14820 (N_14820,N_14704,N_14547);
or U14821 (N_14821,N_14719,N_14702);
or U14822 (N_14822,N_14531,N_14703);
nand U14823 (N_14823,N_14557,N_14664);
and U14824 (N_14824,N_14528,N_14742);
xor U14825 (N_14825,N_14510,N_14667);
nor U14826 (N_14826,N_14513,N_14570);
nand U14827 (N_14827,N_14551,N_14651);
nand U14828 (N_14828,N_14582,N_14644);
nor U14829 (N_14829,N_14530,N_14501);
and U14830 (N_14830,N_14735,N_14658);
or U14831 (N_14831,N_14701,N_14648);
nor U14832 (N_14832,N_14529,N_14730);
xor U14833 (N_14833,N_14598,N_14508);
and U14834 (N_14834,N_14656,N_14680);
xnor U14835 (N_14835,N_14595,N_14568);
nor U14836 (N_14836,N_14533,N_14657);
or U14837 (N_14837,N_14581,N_14683);
or U14838 (N_14838,N_14674,N_14748);
xnor U14839 (N_14839,N_14543,N_14577);
nor U14840 (N_14840,N_14593,N_14682);
or U14841 (N_14841,N_14712,N_14612);
nand U14842 (N_14842,N_14663,N_14546);
or U14843 (N_14843,N_14618,N_14555);
xnor U14844 (N_14844,N_14710,N_14521);
xnor U14845 (N_14845,N_14741,N_14637);
xor U14846 (N_14846,N_14550,N_14553);
nor U14847 (N_14847,N_14526,N_14537);
xor U14848 (N_14848,N_14728,N_14604);
nand U14849 (N_14849,N_14611,N_14596);
and U14850 (N_14850,N_14724,N_14586);
or U14851 (N_14851,N_14542,N_14640);
and U14852 (N_14852,N_14536,N_14722);
xnor U14853 (N_14853,N_14673,N_14736);
and U14854 (N_14854,N_14691,N_14524);
and U14855 (N_14855,N_14512,N_14579);
and U14856 (N_14856,N_14688,N_14626);
and U14857 (N_14857,N_14738,N_14642);
nor U14858 (N_14858,N_14714,N_14647);
xnor U14859 (N_14859,N_14708,N_14560);
and U14860 (N_14860,N_14613,N_14638);
xor U14861 (N_14861,N_14584,N_14733);
and U14862 (N_14862,N_14534,N_14558);
nand U14863 (N_14863,N_14540,N_14599);
nand U14864 (N_14864,N_14747,N_14514);
or U14865 (N_14865,N_14502,N_14631);
nor U14866 (N_14866,N_14676,N_14535);
and U14867 (N_14867,N_14649,N_14671);
nand U14868 (N_14868,N_14518,N_14576);
or U14869 (N_14869,N_14600,N_14717);
and U14870 (N_14870,N_14587,N_14630);
nand U14871 (N_14871,N_14574,N_14580);
or U14872 (N_14872,N_14729,N_14634);
or U14873 (N_14873,N_14628,N_14578);
xor U14874 (N_14874,N_14734,N_14727);
and U14875 (N_14875,N_14572,N_14590);
xnor U14876 (N_14876,N_14686,N_14597);
xnor U14877 (N_14877,N_14607,N_14585);
xor U14878 (N_14878,N_14637,N_14601);
nor U14879 (N_14879,N_14561,N_14685);
nor U14880 (N_14880,N_14566,N_14701);
or U14881 (N_14881,N_14738,N_14637);
xor U14882 (N_14882,N_14728,N_14729);
xor U14883 (N_14883,N_14502,N_14585);
or U14884 (N_14884,N_14562,N_14642);
xnor U14885 (N_14885,N_14538,N_14533);
xnor U14886 (N_14886,N_14614,N_14657);
nand U14887 (N_14887,N_14570,N_14675);
nand U14888 (N_14888,N_14596,N_14711);
or U14889 (N_14889,N_14524,N_14657);
and U14890 (N_14890,N_14590,N_14662);
nor U14891 (N_14891,N_14741,N_14537);
xnor U14892 (N_14892,N_14517,N_14719);
nor U14893 (N_14893,N_14663,N_14729);
nand U14894 (N_14894,N_14615,N_14720);
or U14895 (N_14895,N_14535,N_14598);
nor U14896 (N_14896,N_14707,N_14741);
nor U14897 (N_14897,N_14660,N_14692);
nand U14898 (N_14898,N_14541,N_14636);
xor U14899 (N_14899,N_14599,N_14737);
nor U14900 (N_14900,N_14635,N_14637);
or U14901 (N_14901,N_14739,N_14687);
nor U14902 (N_14902,N_14563,N_14626);
nor U14903 (N_14903,N_14598,N_14696);
nor U14904 (N_14904,N_14543,N_14600);
and U14905 (N_14905,N_14704,N_14740);
xor U14906 (N_14906,N_14543,N_14558);
or U14907 (N_14907,N_14615,N_14590);
nand U14908 (N_14908,N_14642,N_14535);
and U14909 (N_14909,N_14507,N_14560);
nand U14910 (N_14910,N_14668,N_14737);
nor U14911 (N_14911,N_14615,N_14649);
or U14912 (N_14912,N_14561,N_14704);
or U14913 (N_14913,N_14508,N_14678);
and U14914 (N_14914,N_14522,N_14717);
nand U14915 (N_14915,N_14738,N_14673);
nor U14916 (N_14916,N_14722,N_14525);
and U14917 (N_14917,N_14617,N_14734);
or U14918 (N_14918,N_14702,N_14600);
and U14919 (N_14919,N_14581,N_14675);
nand U14920 (N_14920,N_14731,N_14706);
nor U14921 (N_14921,N_14683,N_14631);
and U14922 (N_14922,N_14716,N_14500);
xnor U14923 (N_14923,N_14504,N_14672);
nand U14924 (N_14924,N_14578,N_14637);
xnor U14925 (N_14925,N_14515,N_14618);
nor U14926 (N_14926,N_14588,N_14717);
nand U14927 (N_14927,N_14706,N_14631);
nor U14928 (N_14928,N_14640,N_14669);
and U14929 (N_14929,N_14667,N_14715);
and U14930 (N_14930,N_14683,N_14586);
nor U14931 (N_14931,N_14653,N_14566);
xor U14932 (N_14932,N_14658,N_14612);
or U14933 (N_14933,N_14747,N_14726);
nor U14934 (N_14934,N_14661,N_14671);
nand U14935 (N_14935,N_14526,N_14626);
and U14936 (N_14936,N_14696,N_14686);
xor U14937 (N_14937,N_14703,N_14535);
nand U14938 (N_14938,N_14593,N_14690);
and U14939 (N_14939,N_14705,N_14708);
or U14940 (N_14940,N_14641,N_14546);
or U14941 (N_14941,N_14538,N_14568);
or U14942 (N_14942,N_14531,N_14541);
nor U14943 (N_14943,N_14594,N_14734);
or U14944 (N_14944,N_14676,N_14561);
or U14945 (N_14945,N_14688,N_14591);
nand U14946 (N_14946,N_14546,N_14544);
nor U14947 (N_14947,N_14717,N_14617);
or U14948 (N_14948,N_14621,N_14721);
xnor U14949 (N_14949,N_14704,N_14708);
nand U14950 (N_14950,N_14697,N_14614);
xnor U14951 (N_14951,N_14639,N_14728);
xor U14952 (N_14952,N_14677,N_14736);
and U14953 (N_14953,N_14693,N_14605);
or U14954 (N_14954,N_14710,N_14511);
nand U14955 (N_14955,N_14606,N_14575);
nand U14956 (N_14956,N_14594,N_14682);
or U14957 (N_14957,N_14685,N_14668);
nor U14958 (N_14958,N_14687,N_14578);
or U14959 (N_14959,N_14517,N_14635);
nor U14960 (N_14960,N_14655,N_14563);
xor U14961 (N_14961,N_14732,N_14599);
or U14962 (N_14962,N_14512,N_14740);
nor U14963 (N_14963,N_14513,N_14671);
or U14964 (N_14964,N_14656,N_14725);
nand U14965 (N_14965,N_14591,N_14675);
nand U14966 (N_14966,N_14510,N_14719);
nor U14967 (N_14967,N_14690,N_14671);
nand U14968 (N_14968,N_14724,N_14692);
nor U14969 (N_14969,N_14530,N_14670);
and U14970 (N_14970,N_14589,N_14587);
and U14971 (N_14971,N_14729,N_14549);
or U14972 (N_14972,N_14748,N_14747);
xnor U14973 (N_14973,N_14501,N_14643);
nor U14974 (N_14974,N_14601,N_14713);
nand U14975 (N_14975,N_14654,N_14547);
and U14976 (N_14976,N_14721,N_14608);
or U14977 (N_14977,N_14513,N_14721);
nor U14978 (N_14978,N_14573,N_14612);
nand U14979 (N_14979,N_14561,N_14584);
or U14980 (N_14980,N_14741,N_14566);
and U14981 (N_14981,N_14685,N_14705);
and U14982 (N_14982,N_14733,N_14534);
xor U14983 (N_14983,N_14655,N_14576);
and U14984 (N_14984,N_14622,N_14586);
or U14985 (N_14985,N_14613,N_14629);
nor U14986 (N_14986,N_14742,N_14677);
nor U14987 (N_14987,N_14568,N_14596);
and U14988 (N_14988,N_14622,N_14519);
or U14989 (N_14989,N_14740,N_14531);
and U14990 (N_14990,N_14566,N_14557);
xor U14991 (N_14991,N_14664,N_14653);
or U14992 (N_14992,N_14592,N_14733);
nand U14993 (N_14993,N_14593,N_14669);
nand U14994 (N_14994,N_14579,N_14710);
and U14995 (N_14995,N_14734,N_14660);
nor U14996 (N_14996,N_14740,N_14570);
nor U14997 (N_14997,N_14720,N_14548);
nand U14998 (N_14998,N_14674,N_14745);
or U14999 (N_14999,N_14525,N_14629);
nand U15000 (N_15000,N_14930,N_14856);
or U15001 (N_15001,N_14802,N_14808);
and U15002 (N_15002,N_14803,N_14754);
nand U15003 (N_15003,N_14801,N_14948);
nor U15004 (N_15004,N_14775,N_14950);
xnor U15005 (N_15005,N_14986,N_14816);
xor U15006 (N_15006,N_14954,N_14752);
xnor U15007 (N_15007,N_14955,N_14866);
xnor U15008 (N_15008,N_14818,N_14860);
or U15009 (N_15009,N_14916,N_14852);
nor U15010 (N_15010,N_14871,N_14770);
nand U15011 (N_15011,N_14791,N_14780);
xnor U15012 (N_15012,N_14769,N_14756);
or U15013 (N_15013,N_14751,N_14865);
and U15014 (N_15014,N_14807,N_14913);
xor U15015 (N_15015,N_14755,N_14843);
or U15016 (N_15016,N_14973,N_14840);
nand U15017 (N_15017,N_14814,N_14790);
or U15018 (N_15018,N_14925,N_14792);
nand U15019 (N_15019,N_14810,N_14868);
nand U15020 (N_15020,N_14823,N_14895);
xor U15021 (N_15021,N_14881,N_14809);
nor U15022 (N_15022,N_14857,N_14966);
xnor U15023 (N_15023,N_14781,N_14822);
and U15024 (N_15024,N_14936,N_14864);
nor U15025 (N_15025,N_14982,N_14761);
nand U15026 (N_15026,N_14838,N_14952);
or U15027 (N_15027,N_14820,N_14889);
or U15028 (N_15028,N_14960,N_14855);
or U15029 (N_15029,N_14945,N_14934);
and U15030 (N_15030,N_14845,N_14773);
or U15031 (N_15031,N_14812,N_14772);
xor U15032 (N_15032,N_14819,N_14869);
or U15033 (N_15033,N_14905,N_14969);
and U15034 (N_15034,N_14922,N_14964);
or U15035 (N_15035,N_14811,N_14861);
and U15036 (N_15036,N_14963,N_14996);
xnor U15037 (N_15037,N_14981,N_14940);
and U15038 (N_15038,N_14989,N_14898);
and U15039 (N_15039,N_14927,N_14893);
or U15040 (N_15040,N_14891,N_14980);
nand U15041 (N_15041,N_14892,N_14879);
and U15042 (N_15042,N_14763,N_14789);
or U15043 (N_15043,N_14910,N_14970);
xor U15044 (N_15044,N_14759,N_14830);
nor U15045 (N_15045,N_14967,N_14815);
nand U15046 (N_15046,N_14962,N_14887);
xnor U15047 (N_15047,N_14782,N_14771);
nand U15048 (N_15048,N_14831,N_14833);
nand U15049 (N_15049,N_14850,N_14941);
or U15050 (N_15050,N_14854,N_14827);
nand U15051 (N_15051,N_14999,N_14939);
nor U15052 (N_15052,N_14894,N_14768);
nor U15053 (N_15053,N_14975,N_14813);
xor U15054 (N_15054,N_14929,N_14979);
nand U15055 (N_15055,N_14900,N_14906);
xnor U15056 (N_15056,N_14907,N_14937);
xnor U15057 (N_15057,N_14961,N_14841);
or U15058 (N_15058,N_14793,N_14901);
xor U15059 (N_15059,N_14786,N_14990);
xnor U15060 (N_15060,N_14824,N_14978);
nand U15061 (N_15061,N_14836,N_14942);
and U15062 (N_15062,N_14796,N_14779);
nand U15063 (N_15063,N_14911,N_14873);
xnor U15064 (N_15064,N_14806,N_14784);
nor U15065 (N_15065,N_14971,N_14988);
or U15066 (N_15066,N_14985,N_14870);
xnor U15067 (N_15067,N_14821,N_14798);
xnor U15068 (N_15068,N_14992,N_14957);
nand U15069 (N_15069,N_14919,N_14914);
nand U15070 (N_15070,N_14849,N_14917);
and U15071 (N_15071,N_14903,N_14926);
xnor U15072 (N_15072,N_14765,N_14826);
xor U15073 (N_15073,N_14890,N_14876);
xor U15074 (N_15074,N_14783,N_14977);
xor U15075 (N_15075,N_14994,N_14909);
nor U15076 (N_15076,N_14760,N_14983);
or U15077 (N_15077,N_14825,N_14885);
or U15078 (N_15078,N_14976,N_14928);
xnor U15079 (N_15079,N_14923,N_14920);
xnor U15080 (N_15080,N_14764,N_14993);
xor U15081 (N_15081,N_14959,N_14884);
or U15082 (N_15082,N_14848,N_14767);
nor U15083 (N_15083,N_14862,N_14987);
nand U15084 (N_15084,N_14997,N_14880);
xor U15085 (N_15085,N_14766,N_14839);
xor U15086 (N_15086,N_14785,N_14932);
and U15087 (N_15087,N_14776,N_14956);
nor U15088 (N_15088,N_14858,N_14757);
nand U15089 (N_15089,N_14953,N_14853);
and U15090 (N_15090,N_14998,N_14800);
and U15091 (N_15091,N_14777,N_14859);
nand U15092 (N_15092,N_14947,N_14797);
xor U15093 (N_15093,N_14875,N_14794);
and U15094 (N_15094,N_14995,N_14762);
xnor U15095 (N_15095,N_14984,N_14787);
nor U15096 (N_15096,N_14874,N_14842);
xnor U15097 (N_15097,N_14750,N_14896);
or U15098 (N_15098,N_14958,N_14944);
and U15099 (N_15099,N_14908,N_14883);
or U15100 (N_15100,N_14795,N_14935);
and U15101 (N_15101,N_14804,N_14835);
nor U15102 (N_15102,N_14888,N_14991);
nand U15103 (N_15103,N_14946,N_14968);
or U15104 (N_15104,N_14758,N_14844);
nand U15105 (N_15105,N_14886,N_14828);
or U15106 (N_15106,N_14933,N_14882);
xor U15107 (N_15107,N_14912,N_14846);
or U15108 (N_15108,N_14943,N_14878);
nand U15109 (N_15109,N_14863,N_14938);
and U15110 (N_15110,N_14931,N_14872);
xnor U15111 (N_15111,N_14974,N_14949);
xnor U15112 (N_15112,N_14832,N_14837);
nand U15113 (N_15113,N_14902,N_14753);
and U15114 (N_15114,N_14774,N_14897);
xor U15115 (N_15115,N_14817,N_14921);
or U15116 (N_15116,N_14778,N_14847);
or U15117 (N_15117,N_14904,N_14877);
nand U15118 (N_15118,N_14965,N_14915);
nand U15119 (N_15119,N_14972,N_14951);
or U15120 (N_15120,N_14834,N_14829);
or U15121 (N_15121,N_14899,N_14918);
xnor U15122 (N_15122,N_14924,N_14867);
or U15123 (N_15123,N_14851,N_14805);
or U15124 (N_15124,N_14788,N_14799);
nor U15125 (N_15125,N_14916,N_14813);
or U15126 (N_15126,N_14908,N_14833);
nand U15127 (N_15127,N_14771,N_14992);
nand U15128 (N_15128,N_14796,N_14863);
xnor U15129 (N_15129,N_14950,N_14827);
xnor U15130 (N_15130,N_14809,N_14765);
and U15131 (N_15131,N_14817,N_14770);
and U15132 (N_15132,N_14955,N_14990);
or U15133 (N_15133,N_14927,N_14998);
xor U15134 (N_15134,N_14929,N_14971);
and U15135 (N_15135,N_14967,N_14901);
and U15136 (N_15136,N_14807,N_14923);
xnor U15137 (N_15137,N_14839,N_14927);
or U15138 (N_15138,N_14863,N_14967);
or U15139 (N_15139,N_14913,N_14803);
or U15140 (N_15140,N_14996,N_14940);
nand U15141 (N_15141,N_14913,N_14909);
and U15142 (N_15142,N_14836,N_14935);
xor U15143 (N_15143,N_14966,N_14894);
or U15144 (N_15144,N_14820,N_14874);
xor U15145 (N_15145,N_14838,N_14900);
or U15146 (N_15146,N_14763,N_14924);
and U15147 (N_15147,N_14910,N_14824);
or U15148 (N_15148,N_14981,N_14782);
or U15149 (N_15149,N_14818,N_14940);
xnor U15150 (N_15150,N_14822,N_14948);
nand U15151 (N_15151,N_14963,N_14990);
nand U15152 (N_15152,N_14803,N_14760);
nor U15153 (N_15153,N_14804,N_14993);
nand U15154 (N_15154,N_14777,N_14766);
or U15155 (N_15155,N_14805,N_14885);
or U15156 (N_15156,N_14883,N_14865);
nor U15157 (N_15157,N_14812,N_14767);
or U15158 (N_15158,N_14900,N_14845);
xnor U15159 (N_15159,N_14932,N_14975);
or U15160 (N_15160,N_14988,N_14764);
and U15161 (N_15161,N_14923,N_14795);
xor U15162 (N_15162,N_14947,N_14953);
nor U15163 (N_15163,N_14754,N_14982);
nor U15164 (N_15164,N_14877,N_14799);
or U15165 (N_15165,N_14833,N_14822);
nand U15166 (N_15166,N_14864,N_14900);
xor U15167 (N_15167,N_14868,N_14897);
nand U15168 (N_15168,N_14833,N_14952);
nor U15169 (N_15169,N_14844,N_14896);
nand U15170 (N_15170,N_14996,N_14842);
nor U15171 (N_15171,N_14764,N_14966);
nor U15172 (N_15172,N_14782,N_14899);
nor U15173 (N_15173,N_14856,N_14877);
nor U15174 (N_15174,N_14955,N_14879);
xnor U15175 (N_15175,N_14933,N_14874);
nor U15176 (N_15176,N_14750,N_14907);
nand U15177 (N_15177,N_14830,N_14851);
and U15178 (N_15178,N_14820,N_14764);
nor U15179 (N_15179,N_14900,N_14954);
nor U15180 (N_15180,N_14792,N_14835);
nor U15181 (N_15181,N_14946,N_14878);
nand U15182 (N_15182,N_14875,N_14956);
nand U15183 (N_15183,N_14775,N_14987);
or U15184 (N_15184,N_14872,N_14863);
and U15185 (N_15185,N_14870,N_14855);
nor U15186 (N_15186,N_14788,N_14871);
nand U15187 (N_15187,N_14773,N_14825);
nor U15188 (N_15188,N_14949,N_14986);
nand U15189 (N_15189,N_14758,N_14757);
nand U15190 (N_15190,N_14970,N_14939);
and U15191 (N_15191,N_14942,N_14797);
and U15192 (N_15192,N_14792,N_14794);
and U15193 (N_15193,N_14758,N_14763);
nor U15194 (N_15194,N_14878,N_14797);
nor U15195 (N_15195,N_14883,N_14752);
and U15196 (N_15196,N_14802,N_14769);
xnor U15197 (N_15197,N_14753,N_14952);
nand U15198 (N_15198,N_14883,N_14761);
and U15199 (N_15199,N_14750,N_14922);
nand U15200 (N_15200,N_14941,N_14860);
nor U15201 (N_15201,N_14847,N_14914);
nor U15202 (N_15202,N_14867,N_14831);
nor U15203 (N_15203,N_14862,N_14793);
xor U15204 (N_15204,N_14807,N_14915);
and U15205 (N_15205,N_14879,N_14841);
or U15206 (N_15206,N_14971,N_14765);
nor U15207 (N_15207,N_14796,N_14981);
nor U15208 (N_15208,N_14911,N_14967);
and U15209 (N_15209,N_14980,N_14959);
xor U15210 (N_15210,N_14863,N_14870);
xnor U15211 (N_15211,N_14810,N_14865);
xor U15212 (N_15212,N_14819,N_14814);
and U15213 (N_15213,N_14901,N_14783);
and U15214 (N_15214,N_14900,N_14976);
nor U15215 (N_15215,N_14872,N_14907);
nand U15216 (N_15216,N_14971,N_14870);
or U15217 (N_15217,N_14859,N_14815);
or U15218 (N_15218,N_14851,N_14827);
and U15219 (N_15219,N_14875,N_14872);
and U15220 (N_15220,N_14826,N_14910);
and U15221 (N_15221,N_14771,N_14971);
or U15222 (N_15222,N_14774,N_14830);
nor U15223 (N_15223,N_14964,N_14767);
or U15224 (N_15224,N_14914,N_14897);
or U15225 (N_15225,N_14814,N_14874);
and U15226 (N_15226,N_14915,N_14958);
nor U15227 (N_15227,N_14825,N_14811);
nand U15228 (N_15228,N_14788,N_14760);
nand U15229 (N_15229,N_14962,N_14797);
nor U15230 (N_15230,N_14750,N_14790);
xnor U15231 (N_15231,N_14906,N_14910);
nand U15232 (N_15232,N_14851,N_14997);
nand U15233 (N_15233,N_14768,N_14938);
xnor U15234 (N_15234,N_14916,N_14822);
nand U15235 (N_15235,N_14965,N_14814);
nand U15236 (N_15236,N_14969,N_14853);
or U15237 (N_15237,N_14750,N_14805);
and U15238 (N_15238,N_14867,N_14925);
nor U15239 (N_15239,N_14809,N_14894);
xnor U15240 (N_15240,N_14772,N_14952);
nor U15241 (N_15241,N_14960,N_14998);
or U15242 (N_15242,N_14784,N_14768);
nor U15243 (N_15243,N_14888,N_14942);
and U15244 (N_15244,N_14935,N_14793);
and U15245 (N_15245,N_14890,N_14874);
and U15246 (N_15246,N_14865,N_14945);
xor U15247 (N_15247,N_14940,N_14777);
nor U15248 (N_15248,N_14854,N_14808);
nand U15249 (N_15249,N_14972,N_14804);
or U15250 (N_15250,N_15032,N_15217);
nor U15251 (N_15251,N_15016,N_15006);
nor U15252 (N_15252,N_15180,N_15161);
xor U15253 (N_15253,N_15202,N_15068);
xnor U15254 (N_15254,N_15082,N_15079);
and U15255 (N_15255,N_15237,N_15156);
nand U15256 (N_15256,N_15048,N_15046);
nor U15257 (N_15257,N_15229,N_15085);
xor U15258 (N_15258,N_15001,N_15223);
and U15259 (N_15259,N_15000,N_15135);
xnor U15260 (N_15260,N_15240,N_15113);
or U15261 (N_15261,N_15060,N_15219);
nor U15262 (N_15262,N_15211,N_15033);
nand U15263 (N_15263,N_15142,N_15152);
nor U15264 (N_15264,N_15066,N_15083);
and U15265 (N_15265,N_15153,N_15174);
nor U15266 (N_15266,N_15058,N_15191);
nor U15267 (N_15267,N_15200,N_15099);
xnor U15268 (N_15268,N_15248,N_15098);
nor U15269 (N_15269,N_15246,N_15055);
xor U15270 (N_15270,N_15100,N_15057);
and U15271 (N_15271,N_15070,N_15104);
or U15272 (N_15272,N_15195,N_15030);
or U15273 (N_15273,N_15044,N_15197);
nand U15274 (N_15274,N_15102,N_15158);
nand U15275 (N_15275,N_15242,N_15128);
or U15276 (N_15276,N_15029,N_15167);
nor U15277 (N_15277,N_15010,N_15247);
and U15278 (N_15278,N_15218,N_15215);
nor U15279 (N_15279,N_15072,N_15097);
nor U15280 (N_15280,N_15022,N_15148);
nand U15281 (N_15281,N_15230,N_15224);
xnor U15282 (N_15282,N_15101,N_15053);
xor U15283 (N_15283,N_15170,N_15189);
xor U15284 (N_15284,N_15020,N_15141);
and U15285 (N_15285,N_15171,N_15005);
and U15286 (N_15286,N_15225,N_15136);
or U15287 (N_15287,N_15162,N_15067);
and U15288 (N_15288,N_15077,N_15241);
or U15289 (N_15289,N_15210,N_15112);
or U15290 (N_15290,N_15155,N_15041);
and U15291 (N_15291,N_15184,N_15092);
nand U15292 (N_15292,N_15090,N_15179);
xnor U15293 (N_15293,N_15123,N_15081);
nor U15294 (N_15294,N_15235,N_15116);
and U15295 (N_15295,N_15183,N_15047);
xor U15296 (N_15296,N_15182,N_15118);
xor U15297 (N_15297,N_15011,N_15159);
nor U15298 (N_15298,N_15025,N_15103);
nand U15299 (N_15299,N_15244,N_15089);
nand U15300 (N_15300,N_15194,N_15017);
nand U15301 (N_15301,N_15173,N_15201);
or U15302 (N_15302,N_15045,N_15243);
xnor U15303 (N_15303,N_15132,N_15086);
and U15304 (N_15304,N_15004,N_15088);
nand U15305 (N_15305,N_15129,N_15054);
and U15306 (N_15306,N_15015,N_15056);
or U15307 (N_15307,N_15114,N_15140);
xor U15308 (N_15308,N_15075,N_15169);
nor U15309 (N_15309,N_15065,N_15121);
nor U15310 (N_15310,N_15013,N_15122);
nand U15311 (N_15311,N_15134,N_15031);
nor U15312 (N_15312,N_15049,N_15186);
or U15313 (N_15313,N_15238,N_15157);
xnor U15314 (N_15314,N_15145,N_15038);
nand U15315 (N_15315,N_15115,N_15062);
and U15316 (N_15316,N_15052,N_15014);
and U15317 (N_15317,N_15151,N_15027);
nor U15318 (N_15318,N_15138,N_15106);
nand U15319 (N_15319,N_15076,N_15193);
xor U15320 (N_15320,N_15133,N_15207);
xnor U15321 (N_15321,N_15190,N_15074);
nor U15322 (N_15322,N_15231,N_15012);
and U15323 (N_15323,N_15177,N_15119);
nand U15324 (N_15324,N_15236,N_15093);
or U15325 (N_15325,N_15149,N_15042);
nand U15326 (N_15326,N_15192,N_15245);
nor U15327 (N_15327,N_15080,N_15203);
and U15328 (N_15328,N_15221,N_15206);
and U15329 (N_15329,N_15214,N_15143);
and U15330 (N_15330,N_15063,N_15127);
nor U15331 (N_15331,N_15036,N_15213);
and U15332 (N_15332,N_15175,N_15007);
or U15333 (N_15333,N_15043,N_15146);
nand U15334 (N_15334,N_15154,N_15094);
nand U15335 (N_15335,N_15227,N_15050);
nor U15336 (N_15336,N_15196,N_15105);
xor U15337 (N_15337,N_15232,N_15234);
nor U15338 (N_15338,N_15096,N_15208);
or U15339 (N_15339,N_15233,N_15126);
and U15340 (N_15340,N_15051,N_15163);
nand U15341 (N_15341,N_15064,N_15160);
nand U15342 (N_15342,N_15034,N_15239);
or U15343 (N_15343,N_15108,N_15249);
or U15344 (N_15344,N_15125,N_15059);
nor U15345 (N_15345,N_15139,N_15131);
or U15346 (N_15346,N_15166,N_15087);
xnor U15347 (N_15347,N_15039,N_15117);
xnor U15348 (N_15348,N_15084,N_15176);
or U15349 (N_15349,N_15222,N_15040);
xnor U15350 (N_15350,N_15003,N_15061);
and U15351 (N_15351,N_15037,N_15181);
and U15352 (N_15352,N_15008,N_15091);
or U15353 (N_15353,N_15172,N_15187);
nand U15354 (N_15354,N_15147,N_15120);
and U15355 (N_15355,N_15071,N_15204);
and U15356 (N_15356,N_15110,N_15107);
xor U15357 (N_15357,N_15002,N_15073);
and U15358 (N_15358,N_15009,N_15111);
xnor U15359 (N_15359,N_15124,N_15216);
nor U15360 (N_15360,N_15028,N_15026);
nor U15361 (N_15361,N_15220,N_15212);
xor U15362 (N_15362,N_15095,N_15198);
xor U15363 (N_15363,N_15165,N_15069);
nor U15364 (N_15364,N_15178,N_15078);
nand U15365 (N_15365,N_15185,N_15188);
nand U15366 (N_15366,N_15137,N_15023);
or U15367 (N_15367,N_15035,N_15019);
nand U15368 (N_15368,N_15130,N_15018);
or U15369 (N_15369,N_15021,N_15205);
nor U15370 (N_15370,N_15168,N_15226);
xnor U15371 (N_15371,N_15164,N_15228);
and U15372 (N_15372,N_15024,N_15209);
nor U15373 (N_15373,N_15150,N_15199);
nand U15374 (N_15374,N_15144,N_15109);
nand U15375 (N_15375,N_15020,N_15021);
nand U15376 (N_15376,N_15096,N_15151);
nor U15377 (N_15377,N_15207,N_15120);
and U15378 (N_15378,N_15188,N_15028);
and U15379 (N_15379,N_15072,N_15011);
and U15380 (N_15380,N_15234,N_15139);
nor U15381 (N_15381,N_15128,N_15023);
or U15382 (N_15382,N_15067,N_15148);
nor U15383 (N_15383,N_15015,N_15171);
and U15384 (N_15384,N_15183,N_15153);
or U15385 (N_15385,N_15162,N_15108);
xor U15386 (N_15386,N_15129,N_15004);
and U15387 (N_15387,N_15139,N_15089);
xor U15388 (N_15388,N_15247,N_15043);
nand U15389 (N_15389,N_15180,N_15244);
xnor U15390 (N_15390,N_15017,N_15166);
or U15391 (N_15391,N_15007,N_15099);
nor U15392 (N_15392,N_15212,N_15173);
nor U15393 (N_15393,N_15045,N_15189);
nand U15394 (N_15394,N_15002,N_15190);
nor U15395 (N_15395,N_15119,N_15081);
xnor U15396 (N_15396,N_15135,N_15043);
or U15397 (N_15397,N_15093,N_15005);
and U15398 (N_15398,N_15175,N_15078);
and U15399 (N_15399,N_15158,N_15209);
or U15400 (N_15400,N_15226,N_15044);
or U15401 (N_15401,N_15049,N_15217);
nand U15402 (N_15402,N_15236,N_15042);
and U15403 (N_15403,N_15014,N_15060);
xor U15404 (N_15404,N_15222,N_15042);
and U15405 (N_15405,N_15187,N_15173);
nand U15406 (N_15406,N_15204,N_15181);
xor U15407 (N_15407,N_15043,N_15061);
and U15408 (N_15408,N_15240,N_15044);
and U15409 (N_15409,N_15052,N_15194);
or U15410 (N_15410,N_15107,N_15198);
nor U15411 (N_15411,N_15148,N_15045);
nor U15412 (N_15412,N_15021,N_15067);
and U15413 (N_15413,N_15201,N_15096);
and U15414 (N_15414,N_15012,N_15019);
nand U15415 (N_15415,N_15166,N_15245);
nor U15416 (N_15416,N_15049,N_15132);
nor U15417 (N_15417,N_15054,N_15034);
nor U15418 (N_15418,N_15014,N_15219);
or U15419 (N_15419,N_15144,N_15220);
or U15420 (N_15420,N_15013,N_15031);
nor U15421 (N_15421,N_15173,N_15189);
nand U15422 (N_15422,N_15124,N_15119);
and U15423 (N_15423,N_15234,N_15146);
or U15424 (N_15424,N_15213,N_15193);
xor U15425 (N_15425,N_15181,N_15216);
nor U15426 (N_15426,N_15151,N_15099);
xnor U15427 (N_15427,N_15249,N_15211);
xor U15428 (N_15428,N_15200,N_15091);
nor U15429 (N_15429,N_15032,N_15245);
xor U15430 (N_15430,N_15143,N_15035);
nand U15431 (N_15431,N_15121,N_15150);
nor U15432 (N_15432,N_15102,N_15020);
or U15433 (N_15433,N_15098,N_15008);
nor U15434 (N_15434,N_15248,N_15175);
or U15435 (N_15435,N_15131,N_15192);
or U15436 (N_15436,N_15185,N_15036);
nand U15437 (N_15437,N_15161,N_15162);
nor U15438 (N_15438,N_15040,N_15198);
nand U15439 (N_15439,N_15010,N_15081);
xnor U15440 (N_15440,N_15050,N_15156);
nand U15441 (N_15441,N_15009,N_15043);
xnor U15442 (N_15442,N_15083,N_15014);
and U15443 (N_15443,N_15236,N_15147);
nor U15444 (N_15444,N_15008,N_15248);
xnor U15445 (N_15445,N_15058,N_15196);
nand U15446 (N_15446,N_15234,N_15168);
xor U15447 (N_15447,N_15061,N_15089);
and U15448 (N_15448,N_15018,N_15121);
and U15449 (N_15449,N_15010,N_15056);
nor U15450 (N_15450,N_15016,N_15022);
and U15451 (N_15451,N_15079,N_15126);
nor U15452 (N_15452,N_15126,N_15000);
xor U15453 (N_15453,N_15039,N_15005);
nor U15454 (N_15454,N_15027,N_15100);
or U15455 (N_15455,N_15234,N_15020);
or U15456 (N_15456,N_15192,N_15098);
nor U15457 (N_15457,N_15184,N_15015);
or U15458 (N_15458,N_15208,N_15113);
and U15459 (N_15459,N_15120,N_15102);
or U15460 (N_15460,N_15210,N_15220);
nor U15461 (N_15461,N_15121,N_15100);
or U15462 (N_15462,N_15237,N_15197);
or U15463 (N_15463,N_15059,N_15204);
nand U15464 (N_15464,N_15103,N_15055);
and U15465 (N_15465,N_15006,N_15125);
xor U15466 (N_15466,N_15074,N_15033);
and U15467 (N_15467,N_15171,N_15097);
xor U15468 (N_15468,N_15177,N_15208);
or U15469 (N_15469,N_15133,N_15007);
nand U15470 (N_15470,N_15203,N_15156);
and U15471 (N_15471,N_15046,N_15040);
or U15472 (N_15472,N_15068,N_15214);
nor U15473 (N_15473,N_15206,N_15187);
nand U15474 (N_15474,N_15070,N_15185);
nor U15475 (N_15475,N_15141,N_15072);
nand U15476 (N_15476,N_15103,N_15083);
nor U15477 (N_15477,N_15036,N_15123);
nor U15478 (N_15478,N_15104,N_15248);
and U15479 (N_15479,N_15209,N_15100);
and U15480 (N_15480,N_15053,N_15149);
nand U15481 (N_15481,N_15172,N_15157);
xor U15482 (N_15482,N_15023,N_15174);
nand U15483 (N_15483,N_15077,N_15006);
xnor U15484 (N_15484,N_15216,N_15076);
nor U15485 (N_15485,N_15010,N_15174);
nor U15486 (N_15486,N_15211,N_15225);
nor U15487 (N_15487,N_15013,N_15152);
nand U15488 (N_15488,N_15010,N_15121);
and U15489 (N_15489,N_15232,N_15070);
or U15490 (N_15490,N_15196,N_15166);
nand U15491 (N_15491,N_15122,N_15022);
nand U15492 (N_15492,N_15069,N_15091);
nor U15493 (N_15493,N_15003,N_15247);
nand U15494 (N_15494,N_15230,N_15212);
xnor U15495 (N_15495,N_15191,N_15168);
and U15496 (N_15496,N_15152,N_15079);
nor U15497 (N_15497,N_15225,N_15046);
nand U15498 (N_15498,N_15004,N_15243);
nand U15499 (N_15499,N_15183,N_15185);
nor U15500 (N_15500,N_15457,N_15400);
xor U15501 (N_15501,N_15268,N_15372);
xnor U15502 (N_15502,N_15353,N_15467);
nand U15503 (N_15503,N_15395,N_15284);
nand U15504 (N_15504,N_15498,N_15490);
or U15505 (N_15505,N_15319,N_15443);
and U15506 (N_15506,N_15332,N_15465);
nand U15507 (N_15507,N_15253,N_15391);
nor U15508 (N_15508,N_15338,N_15299);
nand U15509 (N_15509,N_15325,N_15286);
xor U15510 (N_15510,N_15252,N_15274);
nor U15511 (N_15511,N_15261,N_15331);
and U15512 (N_15512,N_15458,N_15424);
nand U15513 (N_15513,N_15446,N_15451);
and U15514 (N_15514,N_15399,N_15484);
and U15515 (N_15515,N_15383,N_15321);
xnor U15516 (N_15516,N_15406,N_15276);
xor U15517 (N_15517,N_15340,N_15402);
nor U15518 (N_15518,N_15384,N_15262);
or U15519 (N_15519,N_15493,N_15295);
or U15520 (N_15520,N_15355,N_15474);
nor U15521 (N_15521,N_15327,N_15390);
and U15522 (N_15522,N_15448,N_15287);
nor U15523 (N_15523,N_15480,N_15344);
nand U15524 (N_15524,N_15449,N_15296);
nor U15525 (N_15525,N_15258,N_15320);
nand U15526 (N_15526,N_15360,N_15381);
and U15527 (N_15527,N_15460,N_15461);
nand U15528 (N_15528,N_15368,N_15456);
xnor U15529 (N_15529,N_15481,N_15339);
nor U15530 (N_15530,N_15293,N_15445);
nor U15531 (N_15531,N_15373,N_15291);
nand U15532 (N_15532,N_15462,N_15315);
nand U15533 (N_15533,N_15447,N_15453);
or U15534 (N_15534,N_15463,N_15392);
xnor U15535 (N_15535,N_15289,N_15483);
or U15536 (N_15536,N_15455,N_15397);
nor U15537 (N_15537,N_15354,N_15270);
xor U15538 (N_15538,N_15301,N_15468);
nor U15539 (N_15539,N_15413,N_15426);
nand U15540 (N_15540,N_15494,N_15288);
nor U15541 (N_15541,N_15491,N_15441);
nor U15542 (N_15542,N_15290,N_15294);
nand U15543 (N_15543,N_15361,N_15489);
or U15544 (N_15544,N_15285,N_15358);
or U15545 (N_15545,N_15302,N_15431);
and U15546 (N_15546,N_15422,N_15326);
xor U15547 (N_15547,N_15470,N_15305);
nor U15548 (N_15548,N_15350,N_15322);
nand U15549 (N_15549,N_15442,N_15382);
and U15550 (N_15550,N_15309,N_15370);
or U15551 (N_15551,N_15497,N_15419);
and U15552 (N_15552,N_15313,N_15495);
xnor U15553 (N_15553,N_15312,N_15482);
or U15554 (N_15554,N_15439,N_15298);
or U15555 (N_15555,N_15264,N_15410);
nor U15556 (N_15556,N_15415,N_15496);
nand U15557 (N_15557,N_15477,N_15267);
nor U15558 (N_15558,N_15405,N_15271);
nand U15559 (N_15559,N_15421,N_15367);
nand U15560 (N_15560,N_15371,N_15475);
nor U15561 (N_15561,N_15254,N_15394);
or U15562 (N_15562,N_15452,N_15377);
xnor U15563 (N_15563,N_15388,N_15478);
xnor U15564 (N_15564,N_15323,N_15356);
and U15565 (N_15565,N_15306,N_15255);
nor U15566 (N_15566,N_15308,N_15420);
nand U15567 (N_15567,N_15486,N_15333);
nand U15568 (N_15568,N_15300,N_15435);
nand U15569 (N_15569,N_15438,N_15335);
and U15570 (N_15570,N_15260,N_15444);
xnor U15571 (N_15571,N_15411,N_15436);
nor U15572 (N_15572,N_15385,N_15269);
xor U15573 (N_15573,N_15409,N_15487);
xor U15574 (N_15574,N_15430,N_15351);
nor U15575 (N_15575,N_15259,N_15330);
and U15576 (N_15576,N_15279,N_15433);
or U15577 (N_15577,N_15250,N_15380);
and U15578 (N_15578,N_15423,N_15329);
or U15579 (N_15579,N_15292,N_15317);
xor U15580 (N_15580,N_15282,N_15256);
xor U15581 (N_15581,N_15459,N_15398);
and U15582 (N_15582,N_15464,N_15473);
nand U15583 (N_15583,N_15472,N_15469);
nand U15584 (N_15584,N_15364,N_15277);
or U15585 (N_15585,N_15348,N_15281);
and U15586 (N_15586,N_15311,N_15432);
and U15587 (N_15587,N_15283,N_15429);
xor U15588 (N_15588,N_15393,N_15273);
nor U15589 (N_15589,N_15466,N_15280);
nor U15590 (N_15590,N_15412,N_15278);
xnor U15591 (N_15591,N_15341,N_15297);
and U15592 (N_15592,N_15345,N_15265);
and U15593 (N_15593,N_15407,N_15352);
nand U15594 (N_15594,N_15314,N_15499);
xnor U15595 (N_15595,N_15266,N_15272);
or U15596 (N_15596,N_15303,N_15428);
nand U15597 (N_15597,N_15257,N_15401);
xnor U15598 (N_15598,N_15434,N_15378);
or U15599 (N_15599,N_15427,N_15359);
nand U15600 (N_15600,N_15369,N_15307);
xor U15601 (N_15601,N_15471,N_15337);
xnor U15602 (N_15602,N_15347,N_15416);
nand U15603 (N_15603,N_15349,N_15488);
nand U15604 (N_15604,N_15414,N_15404);
nor U15605 (N_15605,N_15476,N_15437);
nor U15606 (N_15606,N_15479,N_15366);
nor U15607 (N_15607,N_15316,N_15417);
xor U15608 (N_15608,N_15365,N_15275);
xnor U15609 (N_15609,N_15454,N_15357);
and U15610 (N_15610,N_15304,N_15374);
and U15611 (N_15611,N_15362,N_15425);
or U15612 (N_15612,N_15328,N_15387);
and U15613 (N_15613,N_15440,N_15396);
and U15614 (N_15614,N_15334,N_15251);
xor U15615 (N_15615,N_15324,N_15263);
or U15616 (N_15616,N_15450,N_15492);
and U15617 (N_15617,N_15485,N_15318);
nor U15618 (N_15618,N_15386,N_15408);
and U15619 (N_15619,N_15418,N_15336);
nand U15620 (N_15620,N_15375,N_15346);
or U15621 (N_15621,N_15376,N_15389);
nand U15622 (N_15622,N_15403,N_15363);
nand U15623 (N_15623,N_15342,N_15343);
nand U15624 (N_15624,N_15310,N_15379);
and U15625 (N_15625,N_15299,N_15405);
nand U15626 (N_15626,N_15499,N_15406);
nand U15627 (N_15627,N_15329,N_15309);
nand U15628 (N_15628,N_15346,N_15393);
or U15629 (N_15629,N_15495,N_15399);
or U15630 (N_15630,N_15308,N_15400);
xnor U15631 (N_15631,N_15320,N_15408);
nand U15632 (N_15632,N_15424,N_15426);
or U15633 (N_15633,N_15382,N_15386);
nor U15634 (N_15634,N_15328,N_15316);
nand U15635 (N_15635,N_15283,N_15461);
or U15636 (N_15636,N_15447,N_15467);
xor U15637 (N_15637,N_15433,N_15417);
or U15638 (N_15638,N_15405,N_15252);
and U15639 (N_15639,N_15453,N_15279);
and U15640 (N_15640,N_15418,N_15470);
or U15641 (N_15641,N_15311,N_15454);
xnor U15642 (N_15642,N_15420,N_15406);
xor U15643 (N_15643,N_15360,N_15253);
nor U15644 (N_15644,N_15399,N_15429);
nand U15645 (N_15645,N_15314,N_15372);
xor U15646 (N_15646,N_15403,N_15316);
or U15647 (N_15647,N_15307,N_15370);
and U15648 (N_15648,N_15256,N_15421);
xnor U15649 (N_15649,N_15379,N_15448);
nor U15650 (N_15650,N_15302,N_15434);
nor U15651 (N_15651,N_15253,N_15445);
or U15652 (N_15652,N_15467,N_15383);
xnor U15653 (N_15653,N_15415,N_15318);
xor U15654 (N_15654,N_15379,N_15461);
nor U15655 (N_15655,N_15497,N_15400);
or U15656 (N_15656,N_15283,N_15412);
and U15657 (N_15657,N_15467,N_15269);
nand U15658 (N_15658,N_15368,N_15462);
or U15659 (N_15659,N_15471,N_15330);
or U15660 (N_15660,N_15477,N_15427);
and U15661 (N_15661,N_15292,N_15365);
nand U15662 (N_15662,N_15473,N_15439);
or U15663 (N_15663,N_15391,N_15459);
nand U15664 (N_15664,N_15366,N_15262);
nand U15665 (N_15665,N_15473,N_15481);
nor U15666 (N_15666,N_15295,N_15416);
or U15667 (N_15667,N_15372,N_15371);
or U15668 (N_15668,N_15295,N_15411);
or U15669 (N_15669,N_15449,N_15405);
nand U15670 (N_15670,N_15499,N_15380);
or U15671 (N_15671,N_15305,N_15386);
or U15672 (N_15672,N_15272,N_15277);
nand U15673 (N_15673,N_15289,N_15294);
nand U15674 (N_15674,N_15371,N_15333);
and U15675 (N_15675,N_15257,N_15383);
or U15676 (N_15676,N_15396,N_15304);
and U15677 (N_15677,N_15390,N_15379);
or U15678 (N_15678,N_15468,N_15317);
nand U15679 (N_15679,N_15402,N_15443);
xnor U15680 (N_15680,N_15263,N_15461);
nor U15681 (N_15681,N_15294,N_15326);
and U15682 (N_15682,N_15432,N_15320);
and U15683 (N_15683,N_15429,N_15328);
nor U15684 (N_15684,N_15430,N_15476);
nor U15685 (N_15685,N_15292,N_15285);
nor U15686 (N_15686,N_15345,N_15445);
xnor U15687 (N_15687,N_15487,N_15351);
or U15688 (N_15688,N_15428,N_15449);
nand U15689 (N_15689,N_15493,N_15480);
xnor U15690 (N_15690,N_15338,N_15270);
or U15691 (N_15691,N_15465,N_15497);
nand U15692 (N_15692,N_15332,N_15492);
and U15693 (N_15693,N_15422,N_15459);
nand U15694 (N_15694,N_15466,N_15266);
xor U15695 (N_15695,N_15284,N_15354);
nand U15696 (N_15696,N_15388,N_15477);
or U15697 (N_15697,N_15276,N_15369);
nor U15698 (N_15698,N_15349,N_15433);
xnor U15699 (N_15699,N_15493,N_15462);
nand U15700 (N_15700,N_15422,N_15353);
nand U15701 (N_15701,N_15319,N_15275);
and U15702 (N_15702,N_15484,N_15350);
nand U15703 (N_15703,N_15262,N_15383);
and U15704 (N_15704,N_15391,N_15337);
nor U15705 (N_15705,N_15436,N_15422);
or U15706 (N_15706,N_15301,N_15419);
nor U15707 (N_15707,N_15430,N_15493);
xor U15708 (N_15708,N_15286,N_15295);
nand U15709 (N_15709,N_15430,N_15325);
or U15710 (N_15710,N_15353,N_15299);
and U15711 (N_15711,N_15425,N_15383);
nand U15712 (N_15712,N_15278,N_15366);
nand U15713 (N_15713,N_15495,N_15321);
and U15714 (N_15714,N_15409,N_15278);
and U15715 (N_15715,N_15431,N_15257);
or U15716 (N_15716,N_15351,N_15358);
nand U15717 (N_15717,N_15468,N_15322);
nand U15718 (N_15718,N_15421,N_15391);
or U15719 (N_15719,N_15475,N_15349);
nand U15720 (N_15720,N_15274,N_15412);
or U15721 (N_15721,N_15392,N_15408);
nor U15722 (N_15722,N_15447,N_15470);
nand U15723 (N_15723,N_15390,N_15436);
nor U15724 (N_15724,N_15422,N_15287);
nand U15725 (N_15725,N_15474,N_15349);
nor U15726 (N_15726,N_15331,N_15475);
and U15727 (N_15727,N_15474,N_15314);
and U15728 (N_15728,N_15472,N_15307);
nor U15729 (N_15729,N_15454,N_15414);
and U15730 (N_15730,N_15478,N_15433);
or U15731 (N_15731,N_15475,N_15469);
nand U15732 (N_15732,N_15278,N_15399);
xnor U15733 (N_15733,N_15423,N_15480);
or U15734 (N_15734,N_15344,N_15388);
or U15735 (N_15735,N_15284,N_15494);
and U15736 (N_15736,N_15492,N_15281);
and U15737 (N_15737,N_15345,N_15368);
nand U15738 (N_15738,N_15471,N_15459);
xor U15739 (N_15739,N_15306,N_15339);
nand U15740 (N_15740,N_15495,N_15400);
nor U15741 (N_15741,N_15419,N_15478);
xor U15742 (N_15742,N_15347,N_15269);
and U15743 (N_15743,N_15273,N_15424);
nand U15744 (N_15744,N_15445,N_15275);
nor U15745 (N_15745,N_15482,N_15439);
nor U15746 (N_15746,N_15412,N_15267);
nor U15747 (N_15747,N_15283,N_15420);
and U15748 (N_15748,N_15461,N_15454);
or U15749 (N_15749,N_15369,N_15345);
and U15750 (N_15750,N_15662,N_15622);
nand U15751 (N_15751,N_15613,N_15587);
and U15752 (N_15752,N_15734,N_15569);
and U15753 (N_15753,N_15501,N_15733);
nand U15754 (N_15754,N_15723,N_15642);
xnor U15755 (N_15755,N_15655,N_15696);
nand U15756 (N_15756,N_15740,N_15619);
nor U15757 (N_15757,N_15534,N_15540);
nor U15758 (N_15758,N_15611,N_15718);
nand U15759 (N_15759,N_15679,N_15665);
nor U15760 (N_15760,N_15566,N_15584);
and U15761 (N_15761,N_15511,N_15513);
nor U15762 (N_15762,N_15575,N_15564);
and U15763 (N_15763,N_15746,N_15601);
and U15764 (N_15764,N_15657,N_15681);
nand U15765 (N_15765,N_15710,N_15557);
xnor U15766 (N_15766,N_15570,N_15689);
xor U15767 (N_15767,N_15546,N_15519);
and U15768 (N_15768,N_15634,N_15735);
nand U15769 (N_15769,N_15686,N_15701);
nor U15770 (N_15770,N_15552,N_15661);
nand U15771 (N_15771,N_15722,N_15521);
nor U15772 (N_15772,N_15737,N_15747);
nand U15773 (N_15773,N_15709,N_15640);
xnor U15774 (N_15774,N_15639,N_15563);
nand U15775 (N_15775,N_15620,N_15700);
xnor U15776 (N_15776,N_15533,N_15726);
and U15777 (N_15777,N_15731,N_15715);
xnor U15778 (N_15778,N_15678,N_15724);
and U15779 (N_15779,N_15676,N_15561);
nor U15780 (N_15780,N_15633,N_15605);
nor U15781 (N_15781,N_15682,N_15548);
and U15782 (N_15782,N_15515,N_15608);
xnor U15783 (N_15783,N_15594,N_15738);
or U15784 (N_15784,N_15606,N_15537);
xnor U15785 (N_15785,N_15695,N_15616);
nor U15786 (N_15786,N_15705,N_15547);
and U15787 (N_15787,N_15562,N_15531);
xor U15788 (N_15788,N_15697,N_15589);
and U15789 (N_15789,N_15579,N_15692);
and U15790 (N_15790,N_15627,N_15524);
or U15791 (N_15791,N_15615,N_15716);
nor U15792 (N_15792,N_15599,N_15727);
xnor U15793 (N_15793,N_15623,N_15712);
nand U15794 (N_15794,N_15556,N_15590);
nor U15795 (N_15795,N_15516,N_15517);
nand U15796 (N_15796,N_15539,N_15603);
or U15797 (N_15797,N_15593,N_15532);
nand U15798 (N_15798,N_15672,N_15577);
nand U15799 (N_15799,N_15667,N_15576);
or U15800 (N_15800,N_15635,N_15550);
nand U15801 (N_15801,N_15506,N_15578);
or U15802 (N_15802,N_15643,N_15670);
xor U15803 (N_15803,N_15703,N_15560);
and U15804 (N_15804,N_15505,N_15596);
nand U15805 (N_15805,N_15637,N_15600);
xor U15806 (N_15806,N_15720,N_15618);
nand U15807 (N_15807,N_15729,N_15598);
nand U15808 (N_15808,N_15545,N_15510);
nand U15809 (N_15809,N_15650,N_15630);
nor U15810 (N_15810,N_15684,N_15725);
nor U15811 (N_15811,N_15535,N_15629);
nor U15812 (N_15812,N_15527,N_15607);
and U15813 (N_15813,N_15581,N_15612);
or U15814 (N_15814,N_15644,N_15651);
nor U15815 (N_15815,N_15688,N_15741);
xor U15816 (N_15816,N_15707,N_15687);
and U15817 (N_15817,N_15685,N_15553);
nand U15818 (N_15818,N_15500,N_15572);
nand U15819 (N_15819,N_15609,N_15558);
nand U15820 (N_15820,N_15628,N_15698);
nand U15821 (N_15821,N_15702,N_15694);
nor U15822 (N_15822,N_15666,N_15509);
nor U15823 (N_15823,N_15660,N_15713);
or U15824 (N_15824,N_15652,N_15543);
xnor U15825 (N_15825,N_15518,N_15631);
nand U15826 (N_15826,N_15659,N_15503);
xnor U15827 (N_15827,N_15743,N_15699);
nor U15828 (N_15828,N_15522,N_15582);
or U15829 (N_15829,N_15573,N_15654);
nand U15830 (N_15830,N_15744,N_15568);
nor U15831 (N_15831,N_15604,N_15626);
nand U15832 (N_15832,N_15526,N_15529);
nor U15833 (N_15833,N_15621,N_15711);
nand U15834 (N_15834,N_15671,N_15632);
or U15835 (N_15835,N_15656,N_15648);
or U15836 (N_15836,N_15664,N_15583);
nand U15837 (N_15837,N_15719,N_15544);
xor U15838 (N_15838,N_15668,N_15580);
or U15839 (N_15839,N_15617,N_15536);
xnor U15840 (N_15840,N_15514,N_15591);
or U15841 (N_15841,N_15653,N_15571);
nand U15842 (N_15842,N_15624,N_15704);
and U15843 (N_15843,N_15675,N_15592);
and U15844 (N_15844,N_15673,N_15646);
nor U15845 (N_15845,N_15555,N_15677);
xor U15846 (N_15846,N_15717,N_15645);
or U15847 (N_15847,N_15721,N_15597);
and U15848 (N_15848,N_15706,N_15625);
xor U15849 (N_15849,N_15610,N_15502);
and U15850 (N_15850,N_15736,N_15647);
nand U15851 (N_15851,N_15554,N_15745);
nand U15852 (N_15852,N_15525,N_15551);
and U15853 (N_15853,N_15638,N_15728);
or U15854 (N_15854,N_15574,N_15549);
xnor U15855 (N_15855,N_15586,N_15614);
xor U15856 (N_15856,N_15504,N_15641);
or U15857 (N_15857,N_15742,N_15542);
nand U15858 (N_15858,N_15663,N_15749);
nand U15859 (N_15859,N_15538,N_15658);
and U15860 (N_15860,N_15680,N_15541);
nor U15861 (N_15861,N_15565,N_15520);
xor U15862 (N_15862,N_15714,N_15748);
nand U15863 (N_15863,N_15674,N_15530);
nor U15864 (N_15864,N_15512,N_15690);
xnor U15865 (N_15865,N_15567,N_15507);
xnor U15866 (N_15866,N_15730,N_15691);
or U15867 (N_15867,N_15528,N_15602);
nor U15868 (N_15868,N_15636,N_15588);
nor U15869 (N_15869,N_15708,N_15669);
nand U15870 (N_15870,N_15523,N_15508);
nor U15871 (N_15871,N_15739,N_15595);
and U15872 (N_15872,N_15732,N_15649);
and U15873 (N_15873,N_15559,N_15693);
xor U15874 (N_15874,N_15585,N_15683);
nor U15875 (N_15875,N_15712,N_15708);
xnor U15876 (N_15876,N_15747,N_15529);
and U15877 (N_15877,N_15554,N_15721);
or U15878 (N_15878,N_15653,N_15735);
nand U15879 (N_15879,N_15575,N_15583);
nand U15880 (N_15880,N_15604,N_15593);
or U15881 (N_15881,N_15734,N_15662);
xnor U15882 (N_15882,N_15616,N_15636);
and U15883 (N_15883,N_15704,N_15650);
or U15884 (N_15884,N_15730,N_15574);
xor U15885 (N_15885,N_15502,N_15651);
nand U15886 (N_15886,N_15698,N_15718);
xnor U15887 (N_15887,N_15704,N_15642);
nand U15888 (N_15888,N_15544,N_15640);
nor U15889 (N_15889,N_15721,N_15596);
xnor U15890 (N_15890,N_15663,N_15701);
and U15891 (N_15891,N_15504,N_15682);
nor U15892 (N_15892,N_15521,N_15602);
and U15893 (N_15893,N_15543,N_15553);
nor U15894 (N_15894,N_15728,N_15747);
nor U15895 (N_15895,N_15658,N_15596);
or U15896 (N_15896,N_15592,N_15711);
and U15897 (N_15897,N_15503,N_15695);
xor U15898 (N_15898,N_15630,N_15695);
xnor U15899 (N_15899,N_15653,N_15576);
xor U15900 (N_15900,N_15696,N_15683);
xor U15901 (N_15901,N_15635,N_15655);
xor U15902 (N_15902,N_15538,N_15501);
and U15903 (N_15903,N_15520,N_15716);
xor U15904 (N_15904,N_15691,N_15520);
or U15905 (N_15905,N_15535,N_15659);
nand U15906 (N_15906,N_15748,N_15720);
or U15907 (N_15907,N_15629,N_15560);
xor U15908 (N_15908,N_15562,N_15585);
xor U15909 (N_15909,N_15678,N_15680);
xor U15910 (N_15910,N_15560,N_15577);
nor U15911 (N_15911,N_15609,N_15567);
nor U15912 (N_15912,N_15712,N_15558);
xnor U15913 (N_15913,N_15590,N_15579);
xnor U15914 (N_15914,N_15615,N_15522);
xor U15915 (N_15915,N_15540,N_15554);
nand U15916 (N_15916,N_15586,N_15546);
xor U15917 (N_15917,N_15640,N_15743);
xor U15918 (N_15918,N_15652,N_15712);
nand U15919 (N_15919,N_15629,N_15640);
xor U15920 (N_15920,N_15546,N_15514);
nor U15921 (N_15921,N_15719,N_15725);
and U15922 (N_15922,N_15672,N_15538);
xnor U15923 (N_15923,N_15582,N_15672);
nor U15924 (N_15924,N_15617,N_15506);
or U15925 (N_15925,N_15678,N_15523);
nand U15926 (N_15926,N_15515,N_15634);
xnor U15927 (N_15927,N_15653,N_15515);
nand U15928 (N_15928,N_15629,N_15607);
nand U15929 (N_15929,N_15578,N_15548);
nand U15930 (N_15930,N_15577,N_15711);
nor U15931 (N_15931,N_15503,N_15712);
nand U15932 (N_15932,N_15665,N_15502);
and U15933 (N_15933,N_15597,N_15538);
nor U15934 (N_15934,N_15656,N_15562);
nand U15935 (N_15935,N_15717,N_15588);
nor U15936 (N_15936,N_15689,N_15739);
nor U15937 (N_15937,N_15647,N_15738);
and U15938 (N_15938,N_15626,N_15749);
and U15939 (N_15939,N_15716,N_15601);
nand U15940 (N_15940,N_15514,N_15624);
nand U15941 (N_15941,N_15556,N_15670);
or U15942 (N_15942,N_15680,N_15518);
xor U15943 (N_15943,N_15712,N_15703);
nand U15944 (N_15944,N_15659,N_15611);
xor U15945 (N_15945,N_15669,N_15608);
and U15946 (N_15946,N_15716,N_15645);
nor U15947 (N_15947,N_15654,N_15508);
nor U15948 (N_15948,N_15632,N_15609);
nand U15949 (N_15949,N_15722,N_15708);
and U15950 (N_15950,N_15509,N_15522);
and U15951 (N_15951,N_15669,N_15582);
nor U15952 (N_15952,N_15658,N_15668);
xor U15953 (N_15953,N_15582,N_15648);
or U15954 (N_15954,N_15572,N_15577);
nand U15955 (N_15955,N_15577,N_15549);
nor U15956 (N_15956,N_15543,N_15714);
xnor U15957 (N_15957,N_15601,N_15654);
xnor U15958 (N_15958,N_15596,N_15555);
and U15959 (N_15959,N_15633,N_15585);
or U15960 (N_15960,N_15711,N_15748);
or U15961 (N_15961,N_15637,N_15575);
and U15962 (N_15962,N_15585,N_15528);
or U15963 (N_15963,N_15648,N_15686);
or U15964 (N_15964,N_15506,N_15679);
and U15965 (N_15965,N_15621,N_15598);
xor U15966 (N_15966,N_15630,N_15611);
and U15967 (N_15967,N_15519,N_15647);
or U15968 (N_15968,N_15690,N_15532);
and U15969 (N_15969,N_15725,N_15697);
nor U15970 (N_15970,N_15655,N_15710);
xnor U15971 (N_15971,N_15572,N_15510);
nand U15972 (N_15972,N_15591,N_15557);
and U15973 (N_15973,N_15666,N_15695);
xor U15974 (N_15974,N_15626,N_15651);
nand U15975 (N_15975,N_15633,N_15511);
xor U15976 (N_15976,N_15540,N_15706);
and U15977 (N_15977,N_15728,N_15749);
nand U15978 (N_15978,N_15648,N_15748);
or U15979 (N_15979,N_15500,N_15726);
nand U15980 (N_15980,N_15580,N_15521);
and U15981 (N_15981,N_15680,N_15659);
or U15982 (N_15982,N_15517,N_15510);
nand U15983 (N_15983,N_15534,N_15668);
xor U15984 (N_15984,N_15630,N_15701);
nand U15985 (N_15985,N_15508,N_15525);
nor U15986 (N_15986,N_15706,N_15504);
or U15987 (N_15987,N_15641,N_15747);
nand U15988 (N_15988,N_15732,N_15553);
or U15989 (N_15989,N_15721,N_15575);
xnor U15990 (N_15990,N_15567,N_15740);
nand U15991 (N_15991,N_15724,N_15574);
nor U15992 (N_15992,N_15632,N_15672);
nor U15993 (N_15993,N_15706,N_15545);
xor U15994 (N_15994,N_15542,N_15670);
nor U15995 (N_15995,N_15736,N_15667);
or U15996 (N_15996,N_15593,N_15524);
xnor U15997 (N_15997,N_15590,N_15624);
xnor U15998 (N_15998,N_15558,N_15604);
xnor U15999 (N_15999,N_15670,N_15728);
xnor U16000 (N_16000,N_15870,N_15964);
nor U16001 (N_16001,N_15782,N_15807);
xnor U16002 (N_16002,N_15878,N_15804);
xnor U16003 (N_16003,N_15792,N_15967);
or U16004 (N_16004,N_15852,N_15850);
and U16005 (N_16005,N_15948,N_15906);
xnor U16006 (N_16006,N_15924,N_15921);
and U16007 (N_16007,N_15923,N_15874);
nor U16008 (N_16008,N_15800,N_15755);
or U16009 (N_16009,N_15882,N_15866);
or U16010 (N_16010,N_15846,N_15803);
nor U16011 (N_16011,N_15822,N_15865);
nand U16012 (N_16012,N_15828,N_15756);
xor U16013 (N_16013,N_15830,N_15780);
and U16014 (N_16014,N_15986,N_15890);
xor U16015 (N_16015,N_15784,N_15899);
nor U16016 (N_16016,N_15911,N_15930);
or U16017 (N_16017,N_15751,N_15753);
nand U16018 (N_16018,N_15788,N_15801);
or U16019 (N_16019,N_15974,N_15959);
nor U16020 (N_16020,N_15954,N_15876);
xor U16021 (N_16021,N_15936,N_15851);
nand U16022 (N_16022,N_15848,N_15881);
and U16023 (N_16023,N_15928,N_15957);
xnor U16024 (N_16024,N_15977,N_15945);
nor U16025 (N_16025,N_15769,N_15833);
and U16026 (N_16026,N_15777,N_15982);
and U16027 (N_16027,N_15836,N_15860);
nand U16028 (N_16028,N_15942,N_15900);
nand U16029 (N_16029,N_15898,N_15922);
or U16030 (N_16030,N_15888,N_15950);
and U16031 (N_16031,N_15919,N_15775);
nand U16032 (N_16032,N_15884,N_15811);
or U16033 (N_16033,N_15829,N_15990);
nand U16034 (N_16034,N_15845,N_15816);
and U16035 (N_16035,N_15952,N_15812);
xor U16036 (N_16036,N_15937,N_15971);
nor U16037 (N_16037,N_15931,N_15806);
and U16038 (N_16038,N_15904,N_15757);
nor U16039 (N_16039,N_15824,N_15781);
nor U16040 (N_16040,N_15809,N_15759);
nor U16041 (N_16041,N_15991,N_15794);
nand U16042 (N_16042,N_15879,N_15933);
and U16043 (N_16043,N_15880,N_15802);
and U16044 (N_16044,N_15849,N_15868);
or U16045 (N_16045,N_15791,N_15892);
nor U16046 (N_16046,N_15883,N_15955);
and U16047 (N_16047,N_15915,N_15787);
xnor U16048 (N_16048,N_15839,N_15820);
xor U16049 (N_16049,N_15987,N_15926);
xnor U16050 (N_16050,N_15980,N_15981);
nor U16051 (N_16051,N_15979,N_15855);
or U16052 (N_16052,N_15963,N_15815);
and U16053 (N_16053,N_15873,N_15946);
or U16054 (N_16054,N_15993,N_15837);
nand U16055 (N_16055,N_15841,N_15790);
xor U16056 (N_16056,N_15944,N_15972);
or U16057 (N_16057,N_15795,N_15893);
or U16058 (N_16058,N_15998,N_15798);
xor U16059 (N_16059,N_15786,N_15854);
xor U16060 (N_16060,N_15975,N_15932);
or U16061 (N_16061,N_15805,N_15894);
and U16062 (N_16062,N_15821,N_15970);
and U16063 (N_16063,N_15825,N_15988);
nand U16064 (N_16064,N_15917,N_15760);
xor U16065 (N_16065,N_15861,N_15961);
and U16066 (N_16066,N_15886,N_15871);
xor U16067 (N_16067,N_15918,N_15857);
or U16068 (N_16068,N_15983,N_15935);
and U16069 (N_16069,N_15907,N_15842);
and U16070 (N_16070,N_15997,N_15843);
and U16071 (N_16071,N_15808,N_15896);
or U16072 (N_16072,N_15902,N_15762);
nor U16073 (N_16073,N_15996,N_15771);
nand U16074 (N_16074,N_15814,N_15768);
and U16075 (N_16075,N_15909,N_15877);
nand U16076 (N_16076,N_15976,N_15774);
and U16077 (N_16077,N_15826,N_15905);
nor U16078 (N_16078,N_15785,N_15847);
xor U16079 (N_16079,N_15838,N_15966);
nor U16080 (N_16080,N_15872,N_15913);
and U16081 (N_16081,N_15891,N_15853);
nor U16082 (N_16082,N_15773,N_15914);
nand U16083 (N_16083,N_15764,N_15863);
nand U16084 (N_16084,N_15925,N_15940);
nor U16085 (N_16085,N_15969,N_15889);
nor U16086 (N_16086,N_15758,N_15844);
nand U16087 (N_16087,N_15953,N_15817);
nor U16088 (N_16088,N_15763,N_15875);
nor U16089 (N_16089,N_15897,N_15778);
nand U16090 (N_16090,N_15761,N_15765);
nand U16091 (N_16091,N_15831,N_15810);
and U16092 (N_16092,N_15832,N_15989);
nor U16093 (N_16093,N_15951,N_15862);
nand U16094 (N_16094,N_15772,N_15797);
nor U16095 (N_16095,N_15965,N_15984);
nor U16096 (N_16096,N_15799,N_15869);
or U16097 (N_16097,N_15985,N_15962);
nor U16098 (N_16098,N_15903,N_15767);
nor U16099 (N_16099,N_15920,N_15819);
nor U16100 (N_16100,N_15859,N_15941);
and U16101 (N_16101,N_15929,N_15856);
or U16102 (N_16102,N_15835,N_15895);
and U16103 (N_16103,N_15999,N_15938);
nand U16104 (N_16104,N_15834,N_15864);
or U16105 (N_16105,N_15947,N_15916);
xnor U16106 (N_16106,N_15956,N_15910);
nor U16107 (N_16107,N_15960,N_15992);
nand U16108 (N_16108,N_15912,N_15949);
nand U16109 (N_16109,N_15973,N_15968);
or U16110 (N_16110,N_15823,N_15934);
or U16111 (N_16111,N_15943,N_15939);
nor U16112 (N_16112,N_15858,N_15818);
xnor U16113 (N_16113,N_15754,N_15783);
nand U16114 (N_16114,N_15994,N_15908);
and U16115 (N_16115,N_15789,N_15813);
xor U16116 (N_16116,N_15901,N_15796);
nor U16117 (N_16117,N_15776,N_15793);
xnor U16118 (N_16118,N_15779,N_15958);
xnor U16119 (N_16119,N_15927,N_15766);
or U16120 (N_16120,N_15840,N_15885);
or U16121 (N_16121,N_15770,N_15752);
xor U16122 (N_16122,N_15867,N_15978);
xnor U16123 (N_16123,N_15887,N_15995);
and U16124 (N_16124,N_15750,N_15827);
nor U16125 (N_16125,N_15840,N_15818);
or U16126 (N_16126,N_15919,N_15790);
xnor U16127 (N_16127,N_15999,N_15876);
xor U16128 (N_16128,N_15960,N_15774);
or U16129 (N_16129,N_15918,N_15786);
and U16130 (N_16130,N_15838,N_15820);
nor U16131 (N_16131,N_15870,N_15790);
xor U16132 (N_16132,N_15822,N_15981);
nor U16133 (N_16133,N_15998,N_15768);
xor U16134 (N_16134,N_15812,N_15822);
and U16135 (N_16135,N_15906,N_15946);
or U16136 (N_16136,N_15806,N_15852);
nor U16137 (N_16137,N_15990,N_15764);
and U16138 (N_16138,N_15983,N_15840);
or U16139 (N_16139,N_15908,N_15990);
nand U16140 (N_16140,N_15853,N_15984);
and U16141 (N_16141,N_15810,N_15938);
nor U16142 (N_16142,N_15804,N_15906);
and U16143 (N_16143,N_15888,N_15796);
xor U16144 (N_16144,N_15868,N_15925);
xnor U16145 (N_16145,N_15937,N_15980);
xor U16146 (N_16146,N_15762,N_15929);
nand U16147 (N_16147,N_15792,N_15909);
xor U16148 (N_16148,N_15983,N_15815);
xnor U16149 (N_16149,N_15965,N_15993);
nor U16150 (N_16150,N_15854,N_15971);
or U16151 (N_16151,N_15877,N_15899);
nand U16152 (N_16152,N_15855,N_15848);
xor U16153 (N_16153,N_15774,N_15884);
or U16154 (N_16154,N_15835,N_15803);
and U16155 (N_16155,N_15785,N_15859);
nor U16156 (N_16156,N_15949,N_15907);
xnor U16157 (N_16157,N_15971,N_15870);
or U16158 (N_16158,N_15821,N_15856);
nor U16159 (N_16159,N_15775,N_15768);
nor U16160 (N_16160,N_15774,N_15876);
nand U16161 (N_16161,N_15810,N_15829);
or U16162 (N_16162,N_15946,N_15806);
or U16163 (N_16163,N_15821,N_15812);
nor U16164 (N_16164,N_15922,N_15943);
nor U16165 (N_16165,N_15915,N_15849);
nor U16166 (N_16166,N_15787,N_15840);
nor U16167 (N_16167,N_15934,N_15793);
nor U16168 (N_16168,N_15924,N_15946);
and U16169 (N_16169,N_15932,N_15971);
or U16170 (N_16170,N_15782,N_15973);
xor U16171 (N_16171,N_15997,N_15974);
xnor U16172 (N_16172,N_15870,N_15878);
and U16173 (N_16173,N_15799,N_15853);
and U16174 (N_16174,N_15794,N_15903);
xor U16175 (N_16175,N_15917,N_15813);
xnor U16176 (N_16176,N_15791,N_15943);
nand U16177 (N_16177,N_15836,N_15761);
nor U16178 (N_16178,N_15906,N_15914);
and U16179 (N_16179,N_15974,N_15763);
and U16180 (N_16180,N_15895,N_15964);
xor U16181 (N_16181,N_15896,N_15841);
xor U16182 (N_16182,N_15825,N_15945);
nand U16183 (N_16183,N_15821,N_15807);
and U16184 (N_16184,N_15765,N_15766);
and U16185 (N_16185,N_15808,N_15948);
xor U16186 (N_16186,N_15899,N_15790);
or U16187 (N_16187,N_15839,N_15750);
nand U16188 (N_16188,N_15779,N_15876);
or U16189 (N_16189,N_15814,N_15901);
and U16190 (N_16190,N_15963,N_15988);
and U16191 (N_16191,N_15833,N_15945);
nor U16192 (N_16192,N_15788,N_15919);
and U16193 (N_16193,N_15878,N_15774);
and U16194 (N_16194,N_15923,N_15876);
and U16195 (N_16195,N_15904,N_15921);
and U16196 (N_16196,N_15910,N_15976);
nor U16197 (N_16197,N_15765,N_15801);
nor U16198 (N_16198,N_15761,N_15858);
nor U16199 (N_16199,N_15883,N_15983);
or U16200 (N_16200,N_15945,N_15920);
nor U16201 (N_16201,N_15966,N_15958);
nor U16202 (N_16202,N_15896,N_15964);
xnor U16203 (N_16203,N_15872,N_15961);
xnor U16204 (N_16204,N_15771,N_15784);
or U16205 (N_16205,N_15830,N_15905);
nand U16206 (N_16206,N_15820,N_15997);
or U16207 (N_16207,N_15882,N_15821);
or U16208 (N_16208,N_15950,N_15940);
and U16209 (N_16209,N_15914,N_15887);
nand U16210 (N_16210,N_15845,N_15762);
and U16211 (N_16211,N_15976,N_15802);
or U16212 (N_16212,N_15755,N_15815);
and U16213 (N_16213,N_15909,N_15842);
nand U16214 (N_16214,N_15998,N_15999);
nor U16215 (N_16215,N_15978,N_15989);
nand U16216 (N_16216,N_15777,N_15923);
nor U16217 (N_16217,N_15766,N_15975);
nor U16218 (N_16218,N_15919,N_15768);
nor U16219 (N_16219,N_15811,N_15845);
nor U16220 (N_16220,N_15951,N_15905);
xnor U16221 (N_16221,N_15807,N_15769);
nand U16222 (N_16222,N_15875,N_15805);
nand U16223 (N_16223,N_15900,N_15948);
xnor U16224 (N_16224,N_15863,N_15958);
xnor U16225 (N_16225,N_15772,N_15851);
or U16226 (N_16226,N_15901,N_15893);
nand U16227 (N_16227,N_15816,N_15831);
or U16228 (N_16228,N_15978,N_15841);
nor U16229 (N_16229,N_15915,N_15964);
xor U16230 (N_16230,N_15815,N_15882);
nand U16231 (N_16231,N_15789,N_15751);
xor U16232 (N_16232,N_15981,N_15879);
xor U16233 (N_16233,N_15896,N_15908);
xnor U16234 (N_16234,N_15928,N_15980);
or U16235 (N_16235,N_15999,N_15996);
and U16236 (N_16236,N_15893,N_15887);
nand U16237 (N_16237,N_15832,N_15818);
xnor U16238 (N_16238,N_15757,N_15779);
or U16239 (N_16239,N_15957,N_15986);
nand U16240 (N_16240,N_15912,N_15832);
and U16241 (N_16241,N_15772,N_15890);
nand U16242 (N_16242,N_15912,N_15825);
nor U16243 (N_16243,N_15958,N_15794);
nor U16244 (N_16244,N_15952,N_15979);
nor U16245 (N_16245,N_15762,N_15754);
and U16246 (N_16246,N_15804,N_15940);
nand U16247 (N_16247,N_15808,N_15858);
nand U16248 (N_16248,N_15981,N_15751);
nor U16249 (N_16249,N_15990,N_15773);
or U16250 (N_16250,N_16105,N_16026);
or U16251 (N_16251,N_16154,N_16085);
and U16252 (N_16252,N_16129,N_16127);
or U16253 (N_16253,N_16191,N_16039);
nand U16254 (N_16254,N_16153,N_16041);
or U16255 (N_16255,N_16000,N_16066);
nor U16256 (N_16256,N_16131,N_16175);
and U16257 (N_16257,N_16144,N_16187);
nand U16258 (N_16258,N_16225,N_16184);
xor U16259 (N_16259,N_16083,N_16014);
or U16260 (N_16260,N_16001,N_16005);
nor U16261 (N_16261,N_16013,N_16167);
xnor U16262 (N_16262,N_16218,N_16242);
and U16263 (N_16263,N_16065,N_16090);
nand U16264 (N_16264,N_16019,N_16150);
or U16265 (N_16265,N_16202,N_16155);
and U16266 (N_16266,N_16199,N_16089);
xnor U16267 (N_16267,N_16226,N_16067);
xnor U16268 (N_16268,N_16018,N_16055);
xnor U16269 (N_16269,N_16248,N_16042);
or U16270 (N_16270,N_16078,N_16186);
or U16271 (N_16271,N_16074,N_16180);
nor U16272 (N_16272,N_16240,N_16033);
xnor U16273 (N_16273,N_16221,N_16237);
or U16274 (N_16274,N_16052,N_16235);
nor U16275 (N_16275,N_16209,N_16061);
xor U16276 (N_16276,N_16149,N_16081);
nand U16277 (N_16277,N_16071,N_16073);
nand U16278 (N_16278,N_16134,N_16053);
or U16279 (N_16279,N_16166,N_16130);
or U16280 (N_16280,N_16012,N_16158);
or U16281 (N_16281,N_16137,N_16157);
xor U16282 (N_16282,N_16206,N_16190);
xor U16283 (N_16283,N_16011,N_16006);
or U16284 (N_16284,N_16016,N_16020);
or U16285 (N_16285,N_16007,N_16223);
or U16286 (N_16286,N_16063,N_16173);
nor U16287 (N_16287,N_16247,N_16239);
nand U16288 (N_16288,N_16102,N_16048);
nand U16289 (N_16289,N_16062,N_16230);
nor U16290 (N_16290,N_16058,N_16093);
nor U16291 (N_16291,N_16091,N_16022);
and U16292 (N_16292,N_16215,N_16231);
xnor U16293 (N_16293,N_16243,N_16148);
and U16294 (N_16294,N_16076,N_16030);
xnor U16295 (N_16295,N_16249,N_16228);
xor U16296 (N_16296,N_16161,N_16100);
and U16297 (N_16297,N_16170,N_16171);
and U16298 (N_16298,N_16200,N_16109);
nand U16299 (N_16299,N_16165,N_16128);
nor U16300 (N_16300,N_16234,N_16211);
nor U16301 (N_16301,N_16116,N_16207);
nand U16302 (N_16302,N_16194,N_16138);
and U16303 (N_16303,N_16101,N_16140);
and U16304 (N_16304,N_16189,N_16133);
nor U16305 (N_16305,N_16050,N_16132);
nor U16306 (N_16306,N_16110,N_16070);
nand U16307 (N_16307,N_16009,N_16195);
nor U16308 (N_16308,N_16147,N_16217);
and U16309 (N_16309,N_16172,N_16010);
nand U16310 (N_16310,N_16185,N_16029);
nor U16311 (N_16311,N_16142,N_16017);
nor U16312 (N_16312,N_16168,N_16193);
nand U16313 (N_16313,N_16238,N_16222);
nor U16314 (N_16314,N_16205,N_16088);
or U16315 (N_16315,N_16097,N_16210);
and U16316 (N_16316,N_16213,N_16106);
and U16317 (N_16317,N_16117,N_16037);
nand U16318 (N_16318,N_16060,N_16245);
nor U16319 (N_16319,N_16141,N_16214);
nand U16320 (N_16320,N_16179,N_16224);
or U16321 (N_16321,N_16069,N_16040);
nand U16322 (N_16322,N_16241,N_16125);
and U16323 (N_16323,N_16178,N_16034);
or U16324 (N_16324,N_16181,N_16182);
and U16325 (N_16325,N_16056,N_16162);
nor U16326 (N_16326,N_16087,N_16216);
and U16327 (N_16327,N_16196,N_16021);
xor U16328 (N_16328,N_16108,N_16064);
nor U16329 (N_16329,N_16152,N_16111);
and U16330 (N_16330,N_16057,N_16054);
nor U16331 (N_16331,N_16188,N_16049);
or U16332 (N_16332,N_16115,N_16123);
or U16333 (N_16333,N_16232,N_16164);
nand U16334 (N_16334,N_16004,N_16135);
or U16335 (N_16335,N_16159,N_16174);
xor U16336 (N_16336,N_16051,N_16032);
nor U16337 (N_16337,N_16015,N_16119);
xnor U16338 (N_16338,N_16104,N_16028);
nand U16339 (N_16339,N_16059,N_16204);
and U16340 (N_16340,N_16151,N_16080);
or U16341 (N_16341,N_16244,N_16079);
or U16342 (N_16342,N_16126,N_16068);
xnor U16343 (N_16343,N_16208,N_16008);
xnor U16344 (N_16344,N_16031,N_16113);
nand U16345 (N_16345,N_16219,N_16198);
nand U16346 (N_16346,N_16092,N_16220);
or U16347 (N_16347,N_16146,N_16003);
or U16348 (N_16348,N_16024,N_16169);
and U16349 (N_16349,N_16046,N_16229);
nor U16350 (N_16350,N_16183,N_16145);
or U16351 (N_16351,N_16095,N_16246);
nor U16352 (N_16352,N_16047,N_16099);
and U16353 (N_16353,N_16120,N_16023);
and U16354 (N_16354,N_16035,N_16025);
nor U16355 (N_16355,N_16045,N_16163);
nand U16356 (N_16356,N_16124,N_16094);
or U16357 (N_16357,N_16156,N_16143);
nand U16358 (N_16358,N_16121,N_16197);
or U16359 (N_16359,N_16139,N_16122);
nand U16360 (N_16360,N_16043,N_16114);
and U16361 (N_16361,N_16036,N_16084);
xnor U16362 (N_16362,N_16002,N_16227);
and U16363 (N_16363,N_16201,N_16096);
nor U16364 (N_16364,N_16027,N_16107);
nand U16365 (N_16365,N_16086,N_16176);
or U16366 (N_16366,N_16103,N_16192);
xor U16367 (N_16367,N_16072,N_16075);
nor U16368 (N_16368,N_16038,N_16136);
or U16369 (N_16369,N_16177,N_16077);
and U16370 (N_16370,N_16112,N_16098);
and U16371 (N_16371,N_16236,N_16082);
xnor U16372 (N_16372,N_16044,N_16118);
xnor U16373 (N_16373,N_16203,N_16212);
or U16374 (N_16374,N_16160,N_16233);
nand U16375 (N_16375,N_16230,N_16249);
and U16376 (N_16376,N_16032,N_16002);
nor U16377 (N_16377,N_16200,N_16194);
or U16378 (N_16378,N_16247,N_16055);
and U16379 (N_16379,N_16229,N_16066);
xnor U16380 (N_16380,N_16116,N_16233);
xnor U16381 (N_16381,N_16053,N_16184);
nand U16382 (N_16382,N_16019,N_16242);
xor U16383 (N_16383,N_16249,N_16010);
nand U16384 (N_16384,N_16044,N_16045);
or U16385 (N_16385,N_16004,N_16195);
nor U16386 (N_16386,N_16011,N_16152);
nand U16387 (N_16387,N_16100,N_16067);
and U16388 (N_16388,N_16236,N_16248);
and U16389 (N_16389,N_16119,N_16091);
and U16390 (N_16390,N_16019,N_16186);
nand U16391 (N_16391,N_16104,N_16237);
nand U16392 (N_16392,N_16017,N_16238);
xor U16393 (N_16393,N_16242,N_16037);
nand U16394 (N_16394,N_16013,N_16172);
xor U16395 (N_16395,N_16051,N_16110);
xor U16396 (N_16396,N_16071,N_16082);
or U16397 (N_16397,N_16172,N_16137);
or U16398 (N_16398,N_16202,N_16151);
nor U16399 (N_16399,N_16217,N_16019);
xor U16400 (N_16400,N_16238,N_16107);
xor U16401 (N_16401,N_16096,N_16184);
xor U16402 (N_16402,N_16014,N_16149);
nor U16403 (N_16403,N_16179,N_16119);
nand U16404 (N_16404,N_16189,N_16145);
nand U16405 (N_16405,N_16134,N_16048);
nor U16406 (N_16406,N_16208,N_16150);
nand U16407 (N_16407,N_16040,N_16172);
nor U16408 (N_16408,N_16167,N_16117);
nor U16409 (N_16409,N_16246,N_16152);
or U16410 (N_16410,N_16222,N_16156);
nor U16411 (N_16411,N_16159,N_16071);
xor U16412 (N_16412,N_16231,N_16096);
or U16413 (N_16413,N_16021,N_16229);
xnor U16414 (N_16414,N_16151,N_16085);
nand U16415 (N_16415,N_16183,N_16098);
xnor U16416 (N_16416,N_16244,N_16196);
xor U16417 (N_16417,N_16039,N_16115);
and U16418 (N_16418,N_16242,N_16171);
or U16419 (N_16419,N_16120,N_16125);
nor U16420 (N_16420,N_16008,N_16071);
nand U16421 (N_16421,N_16037,N_16170);
xnor U16422 (N_16422,N_16010,N_16182);
or U16423 (N_16423,N_16189,N_16220);
nor U16424 (N_16424,N_16209,N_16185);
and U16425 (N_16425,N_16111,N_16019);
xnor U16426 (N_16426,N_16238,N_16006);
nor U16427 (N_16427,N_16113,N_16049);
nor U16428 (N_16428,N_16096,N_16049);
or U16429 (N_16429,N_16116,N_16155);
xor U16430 (N_16430,N_16235,N_16227);
nand U16431 (N_16431,N_16063,N_16150);
xnor U16432 (N_16432,N_16208,N_16081);
xnor U16433 (N_16433,N_16220,N_16119);
or U16434 (N_16434,N_16214,N_16163);
xnor U16435 (N_16435,N_16116,N_16128);
nand U16436 (N_16436,N_16101,N_16157);
nor U16437 (N_16437,N_16093,N_16072);
or U16438 (N_16438,N_16237,N_16082);
xor U16439 (N_16439,N_16102,N_16186);
nor U16440 (N_16440,N_16042,N_16032);
nor U16441 (N_16441,N_16004,N_16048);
and U16442 (N_16442,N_16133,N_16209);
or U16443 (N_16443,N_16243,N_16101);
and U16444 (N_16444,N_16210,N_16167);
or U16445 (N_16445,N_16093,N_16118);
and U16446 (N_16446,N_16029,N_16065);
or U16447 (N_16447,N_16006,N_16098);
nor U16448 (N_16448,N_16010,N_16212);
nand U16449 (N_16449,N_16154,N_16064);
or U16450 (N_16450,N_16150,N_16185);
xor U16451 (N_16451,N_16085,N_16153);
nor U16452 (N_16452,N_16216,N_16122);
xnor U16453 (N_16453,N_16189,N_16087);
xnor U16454 (N_16454,N_16103,N_16021);
nand U16455 (N_16455,N_16118,N_16099);
and U16456 (N_16456,N_16099,N_16025);
or U16457 (N_16457,N_16001,N_16052);
xor U16458 (N_16458,N_16111,N_16224);
nor U16459 (N_16459,N_16028,N_16107);
nor U16460 (N_16460,N_16154,N_16197);
nor U16461 (N_16461,N_16049,N_16009);
or U16462 (N_16462,N_16116,N_16051);
nand U16463 (N_16463,N_16175,N_16021);
nor U16464 (N_16464,N_16106,N_16090);
nor U16465 (N_16465,N_16114,N_16232);
and U16466 (N_16466,N_16070,N_16086);
xor U16467 (N_16467,N_16104,N_16147);
nor U16468 (N_16468,N_16147,N_16213);
and U16469 (N_16469,N_16179,N_16107);
nor U16470 (N_16470,N_16147,N_16019);
nor U16471 (N_16471,N_16211,N_16213);
and U16472 (N_16472,N_16068,N_16090);
or U16473 (N_16473,N_16093,N_16161);
and U16474 (N_16474,N_16248,N_16233);
or U16475 (N_16475,N_16039,N_16094);
nand U16476 (N_16476,N_16135,N_16186);
nor U16477 (N_16477,N_16010,N_16066);
or U16478 (N_16478,N_16202,N_16049);
and U16479 (N_16479,N_16156,N_16165);
xor U16480 (N_16480,N_16185,N_16128);
nor U16481 (N_16481,N_16193,N_16190);
xnor U16482 (N_16482,N_16184,N_16155);
or U16483 (N_16483,N_16080,N_16014);
nor U16484 (N_16484,N_16161,N_16118);
nor U16485 (N_16485,N_16109,N_16061);
xnor U16486 (N_16486,N_16179,N_16213);
nand U16487 (N_16487,N_16066,N_16097);
or U16488 (N_16488,N_16126,N_16148);
nand U16489 (N_16489,N_16005,N_16183);
and U16490 (N_16490,N_16132,N_16163);
nand U16491 (N_16491,N_16060,N_16139);
and U16492 (N_16492,N_16194,N_16049);
nand U16493 (N_16493,N_16235,N_16003);
xor U16494 (N_16494,N_16203,N_16199);
nand U16495 (N_16495,N_16032,N_16062);
nand U16496 (N_16496,N_16062,N_16069);
and U16497 (N_16497,N_16033,N_16216);
nor U16498 (N_16498,N_16110,N_16198);
nor U16499 (N_16499,N_16049,N_16077);
nand U16500 (N_16500,N_16347,N_16314);
nor U16501 (N_16501,N_16327,N_16313);
or U16502 (N_16502,N_16364,N_16382);
or U16503 (N_16503,N_16270,N_16442);
nand U16504 (N_16504,N_16480,N_16253);
or U16505 (N_16505,N_16398,N_16300);
xnor U16506 (N_16506,N_16370,N_16404);
or U16507 (N_16507,N_16407,N_16330);
or U16508 (N_16508,N_16291,N_16338);
nor U16509 (N_16509,N_16384,N_16440);
nand U16510 (N_16510,N_16349,N_16340);
nand U16511 (N_16511,N_16392,N_16358);
nand U16512 (N_16512,N_16264,N_16299);
and U16513 (N_16513,N_16287,N_16351);
and U16514 (N_16514,N_16277,N_16254);
xor U16515 (N_16515,N_16388,N_16343);
or U16516 (N_16516,N_16454,N_16260);
and U16517 (N_16517,N_16305,N_16318);
or U16518 (N_16518,N_16280,N_16474);
xnor U16519 (N_16519,N_16290,N_16416);
and U16520 (N_16520,N_16447,N_16256);
nor U16521 (N_16521,N_16333,N_16375);
and U16522 (N_16522,N_16499,N_16345);
nor U16523 (N_16523,N_16437,N_16279);
and U16524 (N_16524,N_16337,N_16460);
xor U16525 (N_16525,N_16451,N_16430);
and U16526 (N_16526,N_16276,N_16387);
nand U16527 (N_16527,N_16262,N_16488);
nor U16528 (N_16528,N_16423,N_16329);
nand U16529 (N_16529,N_16413,N_16301);
xor U16530 (N_16530,N_16355,N_16439);
xnor U16531 (N_16531,N_16402,N_16482);
xnor U16532 (N_16532,N_16306,N_16394);
and U16533 (N_16533,N_16449,N_16255);
or U16534 (N_16534,N_16316,N_16463);
xor U16535 (N_16535,N_16289,N_16292);
xnor U16536 (N_16536,N_16293,N_16479);
and U16537 (N_16537,N_16396,N_16325);
nor U16538 (N_16538,N_16450,N_16335);
nor U16539 (N_16539,N_16434,N_16483);
nor U16540 (N_16540,N_16436,N_16432);
nand U16541 (N_16541,N_16371,N_16295);
or U16542 (N_16542,N_16465,N_16378);
nand U16543 (N_16543,N_16310,N_16428);
xor U16544 (N_16544,N_16429,N_16275);
nand U16545 (N_16545,N_16419,N_16263);
nor U16546 (N_16546,N_16328,N_16359);
nand U16547 (N_16547,N_16362,N_16354);
and U16548 (N_16548,N_16494,N_16455);
xnor U16549 (N_16549,N_16357,N_16323);
nand U16550 (N_16550,N_16433,N_16380);
nand U16551 (N_16551,N_16298,N_16485);
nand U16552 (N_16552,N_16350,N_16406);
xnor U16553 (N_16553,N_16268,N_16274);
xor U16554 (N_16554,N_16311,N_16348);
nand U16555 (N_16555,N_16484,N_16441);
and U16556 (N_16556,N_16409,N_16251);
or U16557 (N_16557,N_16444,N_16438);
and U16558 (N_16558,N_16472,N_16464);
nor U16559 (N_16559,N_16397,N_16372);
nor U16560 (N_16560,N_16495,N_16385);
and U16561 (N_16561,N_16252,N_16352);
or U16562 (N_16562,N_16284,N_16381);
nand U16563 (N_16563,N_16288,N_16400);
nor U16564 (N_16564,N_16422,N_16258);
and U16565 (N_16565,N_16377,N_16336);
xor U16566 (N_16566,N_16265,N_16391);
nor U16567 (N_16567,N_16490,N_16331);
and U16568 (N_16568,N_16273,N_16383);
xor U16569 (N_16569,N_16294,N_16346);
or U16570 (N_16570,N_16344,N_16315);
xnor U16571 (N_16571,N_16424,N_16477);
nand U16572 (N_16572,N_16443,N_16312);
xor U16573 (N_16573,N_16309,N_16373);
nand U16574 (N_16574,N_16326,N_16486);
nor U16575 (N_16575,N_16487,N_16390);
xor U16576 (N_16576,N_16417,N_16399);
or U16577 (N_16577,N_16386,N_16341);
or U16578 (N_16578,N_16420,N_16478);
nor U16579 (N_16579,N_16324,N_16456);
nor U16580 (N_16580,N_16389,N_16481);
or U16581 (N_16581,N_16403,N_16452);
and U16582 (N_16582,N_16446,N_16410);
nor U16583 (N_16583,N_16414,N_16411);
nand U16584 (N_16584,N_16368,N_16269);
nand U16585 (N_16585,N_16493,N_16489);
and U16586 (N_16586,N_16457,N_16365);
nand U16587 (N_16587,N_16283,N_16304);
nand U16588 (N_16588,N_16496,N_16469);
nor U16589 (N_16589,N_16307,N_16401);
and U16590 (N_16590,N_16425,N_16408);
and U16591 (N_16591,N_16353,N_16302);
and U16592 (N_16592,N_16459,N_16278);
nor U16593 (N_16593,N_16281,N_16285);
nand U16594 (N_16594,N_16257,N_16492);
and U16595 (N_16595,N_16320,N_16250);
or U16596 (N_16596,N_16393,N_16427);
nand U16597 (N_16597,N_16376,N_16259);
and U16598 (N_16598,N_16308,N_16470);
or U16599 (N_16599,N_16272,N_16367);
nor U16600 (N_16600,N_16426,N_16303);
xor U16601 (N_16601,N_16418,N_16475);
and U16602 (N_16602,N_16435,N_16491);
and U16603 (N_16603,N_16468,N_16461);
and U16604 (N_16604,N_16296,N_16322);
or U16605 (N_16605,N_16476,N_16356);
nand U16606 (N_16606,N_16379,N_16261);
xnor U16607 (N_16607,N_16267,N_16374);
and U16608 (N_16608,N_16366,N_16412);
and U16609 (N_16609,N_16369,N_16453);
nand U16610 (N_16610,N_16421,N_16458);
xnor U16611 (N_16611,N_16405,N_16415);
or U16612 (N_16612,N_16462,N_16473);
or U16613 (N_16613,N_16334,N_16317);
nor U16614 (N_16614,N_16497,N_16360);
xnor U16615 (N_16615,N_16395,N_16286);
or U16616 (N_16616,N_16342,N_16271);
or U16617 (N_16617,N_16321,N_16498);
nor U16618 (N_16618,N_16445,N_16319);
xnor U16619 (N_16619,N_16467,N_16363);
nand U16620 (N_16620,N_16361,N_16466);
or U16621 (N_16621,N_16431,N_16282);
or U16622 (N_16622,N_16448,N_16339);
nand U16623 (N_16623,N_16332,N_16471);
and U16624 (N_16624,N_16266,N_16297);
nor U16625 (N_16625,N_16260,N_16272);
nand U16626 (N_16626,N_16458,N_16443);
and U16627 (N_16627,N_16486,N_16494);
or U16628 (N_16628,N_16353,N_16342);
nand U16629 (N_16629,N_16307,N_16475);
nor U16630 (N_16630,N_16493,N_16408);
nor U16631 (N_16631,N_16391,N_16435);
and U16632 (N_16632,N_16346,N_16462);
xnor U16633 (N_16633,N_16471,N_16257);
and U16634 (N_16634,N_16457,N_16449);
nand U16635 (N_16635,N_16252,N_16300);
and U16636 (N_16636,N_16439,N_16446);
nor U16637 (N_16637,N_16445,N_16359);
nand U16638 (N_16638,N_16366,N_16393);
nor U16639 (N_16639,N_16406,N_16261);
and U16640 (N_16640,N_16417,N_16486);
or U16641 (N_16641,N_16397,N_16434);
or U16642 (N_16642,N_16421,N_16434);
xor U16643 (N_16643,N_16441,N_16372);
or U16644 (N_16644,N_16437,N_16413);
or U16645 (N_16645,N_16397,N_16409);
xor U16646 (N_16646,N_16446,N_16416);
nor U16647 (N_16647,N_16299,N_16347);
nand U16648 (N_16648,N_16306,N_16472);
xnor U16649 (N_16649,N_16432,N_16372);
nor U16650 (N_16650,N_16320,N_16469);
or U16651 (N_16651,N_16378,N_16380);
nand U16652 (N_16652,N_16355,N_16476);
nor U16653 (N_16653,N_16298,N_16488);
xor U16654 (N_16654,N_16279,N_16366);
nand U16655 (N_16655,N_16290,N_16352);
or U16656 (N_16656,N_16407,N_16428);
xnor U16657 (N_16657,N_16481,N_16293);
xor U16658 (N_16658,N_16410,N_16256);
nor U16659 (N_16659,N_16346,N_16468);
xor U16660 (N_16660,N_16325,N_16326);
xnor U16661 (N_16661,N_16296,N_16301);
and U16662 (N_16662,N_16338,N_16462);
or U16663 (N_16663,N_16365,N_16398);
xor U16664 (N_16664,N_16435,N_16342);
and U16665 (N_16665,N_16332,N_16349);
nand U16666 (N_16666,N_16327,N_16353);
or U16667 (N_16667,N_16303,N_16307);
nand U16668 (N_16668,N_16398,N_16263);
nand U16669 (N_16669,N_16397,N_16332);
or U16670 (N_16670,N_16333,N_16393);
nand U16671 (N_16671,N_16355,N_16374);
nor U16672 (N_16672,N_16320,N_16304);
xor U16673 (N_16673,N_16406,N_16415);
and U16674 (N_16674,N_16482,N_16322);
nand U16675 (N_16675,N_16293,N_16417);
nand U16676 (N_16676,N_16368,N_16413);
nor U16677 (N_16677,N_16364,N_16345);
nand U16678 (N_16678,N_16401,N_16389);
nand U16679 (N_16679,N_16494,N_16496);
nand U16680 (N_16680,N_16489,N_16495);
nand U16681 (N_16681,N_16484,N_16496);
nand U16682 (N_16682,N_16435,N_16394);
nor U16683 (N_16683,N_16289,N_16358);
or U16684 (N_16684,N_16467,N_16489);
or U16685 (N_16685,N_16491,N_16396);
or U16686 (N_16686,N_16425,N_16490);
nor U16687 (N_16687,N_16360,N_16383);
xor U16688 (N_16688,N_16291,N_16499);
nor U16689 (N_16689,N_16499,N_16453);
and U16690 (N_16690,N_16369,N_16281);
xor U16691 (N_16691,N_16473,N_16297);
or U16692 (N_16692,N_16452,N_16341);
nor U16693 (N_16693,N_16394,N_16368);
xor U16694 (N_16694,N_16414,N_16266);
nor U16695 (N_16695,N_16439,N_16378);
xnor U16696 (N_16696,N_16307,N_16325);
and U16697 (N_16697,N_16286,N_16341);
xnor U16698 (N_16698,N_16309,N_16393);
or U16699 (N_16699,N_16383,N_16298);
nand U16700 (N_16700,N_16497,N_16325);
and U16701 (N_16701,N_16467,N_16451);
xor U16702 (N_16702,N_16262,N_16383);
nand U16703 (N_16703,N_16430,N_16406);
nor U16704 (N_16704,N_16257,N_16258);
or U16705 (N_16705,N_16365,N_16364);
nor U16706 (N_16706,N_16280,N_16352);
xor U16707 (N_16707,N_16271,N_16337);
nor U16708 (N_16708,N_16493,N_16450);
or U16709 (N_16709,N_16278,N_16322);
nor U16710 (N_16710,N_16349,N_16393);
or U16711 (N_16711,N_16285,N_16299);
or U16712 (N_16712,N_16275,N_16469);
xnor U16713 (N_16713,N_16292,N_16265);
and U16714 (N_16714,N_16404,N_16455);
xnor U16715 (N_16715,N_16418,N_16370);
nand U16716 (N_16716,N_16327,N_16282);
nor U16717 (N_16717,N_16427,N_16277);
or U16718 (N_16718,N_16431,N_16292);
xor U16719 (N_16719,N_16493,N_16284);
and U16720 (N_16720,N_16386,N_16367);
or U16721 (N_16721,N_16402,N_16306);
nand U16722 (N_16722,N_16418,N_16314);
or U16723 (N_16723,N_16391,N_16277);
or U16724 (N_16724,N_16441,N_16429);
or U16725 (N_16725,N_16483,N_16428);
or U16726 (N_16726,N_16282,N_16382);
nor U16727 (N_16727,N_16410,N_16440);
nand U16728 (N_16728,N_16352,N_16438);
xnor U16729 (N_16729,N_16331,N_16262);
or U16730 (N_16730,N_16450,N_16466);
or U16731 (N_16731,N_16301,N_16460);
or U16732 (N_16732,N_16485,N_16450);
xnor U16733 (N_16733,N_16387,N_16460);
or U16734 (N_16734,N_16383,N_16475);
nor U16735 (N_16735,N_16256,N_16292);
nor U16736 (N_16736,N_16336,N_16347);
nand U16737 (N_16737,N_16311,N_16482);
or U16738 (N_16738,N_16319,N_16407);
nand U16739 (N_16739,N_16297,N_16491);
xor U16740 (N_16740,N_16318,N_16417);
xor U16741 (N_16741,N_16277,N_16327);
and U16742 (N_16742,N_16302,N_16327);
or U16743 (N_16743,N_16256,N_16411);
xor U16744 (N_16744,N_16281,N_16305);
xnor U16745 (N_16745,N_16400,N_16375);
nand U16746 (N_16746,N_16369,N_16318);
nand U16747 (N_16747,N_16459,N_16314);
nand U16748 (N_16748,N_16357,N_16268);
or U16749 (N_16749,N_16263,N_16301);
or U16750 (N_16750,N_16714,N_16546);
xnor U16751 (N_16751,N_16678,N_16599);
nand U16752 (N_16752,N_16561,N_16555);
xor U16753 (N_16753,N_16593,N_16648);
nor U16754 (N_16754,N_16549,N_16713);
nand U16755 (N_16755,N_16532,N_16706);
or U16756 (N_16756,N_16630,N_16540);
xnor U16757 (N_16757,N_16600,N_16594);
xnor U16758 (N_16758,N_16533,N_16591);
and U16759 (N_16759,N_16615,N_16718);
nand U16760 (N_16760,N_16659,N_16573);
or U16761 (N_16761,N_16661,N_16535);
nand U16762 (N_16762,N_16683,N_16585);
nor U16763 (N_16763,N_16622,N_16520);
or U16764 (N_16764,N_16657,N_16514);
or U16765 (N_16765,N_16551,N_16562);
or U16766 (N_16766,N_16627,N_16671);
nand U16767 (N_16767,N_16628,N_16577);
nor U16768 (N_16768,N_16595,N_16696);
nand U16769 (N_16769,N_16674,N_16726);
nand U16770 (N_16770,N_16544,N_16582);
and U16771 (N_16771,N_16724,N_16526);
or U16772 (N_16772,N_16608,N_16579);
nand U16773 (N_16773,N_16655,N_16513);
xnor U16774 (N_16774,N_16524,N_16587);
or U16775 (N_16775,N_16702,N_16580);
nand U16776 (N_16776,N_16605,N_16601);
nor U16777 (N_16777,N_16704,N_16745);
xnor U16778 (N_16778,N_16505,N_16639);
nand U16779 (N_16779,N_16735,N_16649);
xnor U16780 (N_16780,N_16565,N_16665);
or U16781 (N_16781,N_16528,N_16695);
nor U16782 (N_16782,N_16529,N_16643);
nor U16783 (N_16783,N_16684,N_16614);
xor U16784 (N_16784,N_16590,N_16530);
xor U16785 (N_16785,N_16557,N_16602);
nand U16786 (N_16786,N_16584,N_16581);
nor U16787 (N_16787,N_16663,N_16570);
xnor U16788 (N_16788,N_16617,N_16653);
nor U16789 (N_16789,N_16621,N_16693);
nor U16790 (N_16790,N_16749,N_16723);
and U16791 (N_16791,N_16554,N_16597);
xor U16792 (N_16792,N_16603,N_16728);
or U16793 (N_16793,N_16652,N_16700);
xor U16794 (N_16794,N_16576,N_16681);
xnor U16795 (N_16795,N_16673,N_16699);
or U16796 (N_16796,N_16720,N_16536);
nor U16797 (N_16797,N_16701,N_16645);
nor U16798 (N_16798,N_16690,N_16734);
and U16799 (N_16799,N_16741,N_16672);
nand U16800 (N_16800,N_16626,N_16620);
and U16801 (N_16801,N_16742,N_16527);
or U16802 (N_16802,N_16548,N_16613);
and U16803 (N_16803,N_16619,N_16710);
nor U16804 (N_16804,N_16509,N_16564);
nor U16805 (N_16805,N_16629,N_16503);
and U16806 (N_16806,N_16539,N_16574);
nor U16807 (N_16807,N_16654,N_16623);
or U16808 (N_16808,N_16521,N_16725);
nand U16809 (N_16809,N_16685,N_16666);
or U16810 (N_16810,N_16646,N_16716);
or U16811 (N_16811,N_16715,N_16598);
xnor U16812 (N_16812,N_16522,N_16586);
and U16813 (N_16813,N_16727,N_16578);
or U16814 (N_16814,N_16680,N_16531);
nand U16815 (N_16815,N_16604,N_16670);
xnor U16816 (N_16816,N_16634,N_16592);
xnor U16817 (N_16817,N_16631,N_16687);
and U16818 (N_16818,N_16553,N_16688);
nand U16819 (N_16819,N_16560,N_16607);
nand U16820 (N_16820,N_16534,N_16717);
or U16821 (N_16821,N_16606,N_16571);
nor U16822 (N_16822,N_16552,N_16675);
and U16823 (N_16823,N_16517,N_16538);
xor U16824 (N_16824,N_16677,N_16508);
and U16825 (N_16825,N_16709,N_16500);
xor U16826 (N_16826,N_16523,N_16712);
nand U16827 (N_16827,N_16545,N_16641);
xor U16828 (N_16828,N_16697,N_16501);
or U16829 (N_16829,N_16705,N_16633);
and U16830 (N_16830,N_16612,N_16518);
nor U16831 (N_16831,N_16737,N_16588);
nand U16832 (N_16832,N_16694,N_16721);
nand U16833 (N_16833,N_16610,N_16686);
nand U16834 (N_16834,N_16525,N_16719);
xnor U16835 (N_16835,N_16519,N_16502);
nor U16836 (N_16836,N_16676,N_16730);
xnor U16837 (N_16837,N_16618,N_16667);
xor U16838 (N_16838,N_16510,N_16583);
nand U16839 (N_16839,N_16572,N_16722);
or U16840 (N_16840,N_16711,N_16746);
xnor U16841 (N_16841,N_16708,N_16550);
xor U16842 (N_16842,N_16506,N_16689);
nand U16843 (N_16843,N_16732,N_16658);
xnor U16844 (N_16844,N_16691,N_16596);
or U16845 (N_16845,N_16575,N_16543);
xor U16846 (N_16846,N_16662,N_16556);
nor U16847 (N_16847,N_16512,N_16638);
or U16848 (N_16848,N_16731,N_16611);
nand U16849 (N_16849,N_16563,N_16625);
nand U16850 (N_16850,N_16747,N_16740);
nor U16851 (N_16851,N_16566,N_16568);
or U16852 (N_16852,N_16569,N_16733);
and U16853 (N_16853,N_16692,N_16542);
xnor U16854 (N_16854,N_16743,N_16609);
xnor U16855 (N_16855,N_16644,N_16748);
xnor U16856 (N_16856,N_16736,N_16729);
nor U16857 (N_16857,N_16547,N_16651);
or U16858 (N_16858,N_16637,N_16589);
or U16859 (N_16859,N_16635,N_16616);
nand U16860 (N_16860,N_16567,N_16624);
or U16861 (N_16861,N_16703,N_16647);
xnor U16862 (N_16862,N_16558,N_16507);
nand U16863 (N_16863,N_16632,N_16664);
nand U16864 (N_16864,N_16698,N_16640);
xor U16865 (N_16865,N_16636,N_16668);
nand U16866 (N_16866,N_16739,N_16679);
nor U16867 (N_16867,N_16707,N_16541);
nor U16868 (N_16868,N_16738,N_16669);
or U16869 (N_16869,N_16650,N_16642);
xor U16870 (N_16870,N_16682,N_16537);
and U16871 (N_16871,N_16515,N_16511);
nor U16872 (N_16872,N_16656,N_16516);
xor U16873 (N_16873,N_16504,N_16559);
nand U16874 (N_16874,N_16660,N_16744);
nor U16875 (N_16875,N_16515,N_16702);
nor U16876 (N_16876,N_16613,N_16516);
nand U16877 (N_16877,N_16709,N_16527);
nand U16878 (N_16878,N_16539,N_16748);
xnor U16879 (N_16879,N_16550,N_16512);
and U16880 (N_16880,N_16517,N_16523);
nor U16881 (N_16881,N_16654,N_16581);
xor U16882 (N_16882,N_16574,N_16563);
nor U16883 (N_16883,N_16545,N_16604);
or U16884 (N_16884,N_16632,N_16724);
and U16885 (N_16885,N_16656,N_16588);
nor U16886 (N_16886,N_16715,N_16521);
xnor U16887 (N_16887,N_16713,N_16584);
nand U16888 (N_16888,N_16711,N_16632);
and U16889 (N_16889,N_16700,N_16714);
or U16890 (N_16890,N_16548,N_16515);
nand U16891 (N_16891,N_16639,N_16657);
and U16892 (N_16892,N_16670,N_16737);
and U16893 (N_16893,N_16543,N_16566);
or U16894 (N_16894,N_16735,N_16584);
xnor U16895 (N_16895,N_16583,N_16667);
and U16896 (N_16896,N_16745,N_16565);
or U16897 (N_16897,N_16570,N_16727);
and U16898 (N_16898,N_16509,N_16622);
nor U16899 (N_16899,N_16660,N_16561);
or U16900 (N_16900,N_16595,N_16544);
xor U16901 (N_16901,N_16620,N_16581);
xnor U16902 (N_16902,N_16654,N_16651);
xor U16903 (N_16903,N_16605,N_16655);
or U16904 (N_16904,N_16610,N_16524);
and U16905 (N_16905,N_16509,N_16668);
and U16906 (N_16906,N_16503,N_16592);
and U16907 (N_16907,N_16689,N_16546);
xnor U16908 (N_16908,N_16561,N_16503);
nand U16909 (N_16909,N_16516,N_16587);
xnor U16910 (N_16910,N_16528,N_16582);
xnor U16911 (N_16911,N_16502,N_16594);
or U16912 (N_16912,N_16633,N_16640);
nor U16913 (N_16913,N_16584,N_16508);
xnor U16914 (N_16914,N_16600,N_16549);
xor U16915 (N_16915,N_16582,N_16713);
nor U16916 (N_16916,N_16647,N_16513);
nand U16917 (N_16917,N_16548,N_16645);
or U16918 (N_16918,N_16552,N_16713);
or U16919 (N_16919,N_16713,N_16686);
nor U16920 (N_16920,N_16579,N_16568);
and U16921 (N_16921,N_16595,N_16632);
xnor U16922 (N_16922,N_16738,N_16728);
or U16923 (N_16923,N_16619,N_16565);
nand U16924 (N_16924,N_16640,N_16693);
xnor U16925 (N_16925,N_16508,N_16749);
or U16926 (N_16926,N_16574,N_16740);
nand U16927 (N_16927,N_16590,N_16528);
nor U16928 (N_16928,N_16685,N_16633);
and U16929 (N_16929,N_16556,N_16716);
nor U16930 (N_16930,N_16697,N_16673);
xor U16931 (N_16931,N_16745,N_16663);
nor U16932 (N_16932,N_16746,N_16717);
xnor U16933 (N_16933,N_16560,N_16734);
or U16934 (N_16934,N_16609,N_16710);
and U16935 (N_16935,N_16620,N_16723);
xnor U16936 (N_16936,N_16720,N_16541);
nor U16937 (N_16937,N_16536,N_16726);
and U16938 (N_16938,N_16594,N_16696);
nor U16939 (N_16939,N_16606,N_16560);
nor U16940 (N_16940,N_16540,N_16642);
and U16941 (N_16941,N_16625,N_16714);
xnor U16942 (N_16942,N_16599,N_16639);
nand U16943 (N_16943,N_16715,N_16514);
and U16944 (N_16944,N_16580,N_16666);
and U16945 (N_16945,N_16716,N_16577);
nand U16946 (N_16946,N_16653,N_16583);
and U16947 (N_16947,N_16744,N_16624);
nand U16948 (N_16948,N_16698,N_16571);
xor U16949 (N_16949,N_16596,N_16630);
xor U16950 (N_16950,N_16557,N_16535);
and U16951 (N_16951,N_16739,N_16684);
nand U16952 (N_16952,N_16652,N_16579);
nand U16953 (N_16953,N_16719,N_16741);
nor U16954 (N_16954,N_16713,N_16519);
nor U16955 (N_16955,N_16633,N_16511);
nor U16956 (N_16956,N_16671,N_16674);
xor U16957 (N_16957,N_16745,N_16730);
or U16958 (N_16958,N_16631,N_16573);
or U16959 (N_16959,N_16603,N_16666);
and U16960 (N_16960,N_16727,N_16663);
or U16961 (N_16961,N_16648,N_16651);
or U16962 (N_16962,N_16706,N_16551);
nor U16963 (N_16963,N_16717,N_16552);
xnor U16964 (N_16964,N_16544,N_16562);
xor U16965 (N_16965,N_16618,N_16586);
xnor U16966 (N_16966,N_16575,N_16506);
xor U16967 (N_16967,N_16719,N_16593);
nand U16968 (N_16968,N_16629,N_16626);
xor U16969 (N_16969,N_16568,N_16672);
or U16970 (N_16970,N_16523,N_16708);
nor U16971 (N_16971,N_16529,N_16627);
nand U16972 (N_16972,N_16686,N_16655);
nand U16973 (N_16973,N_16542,N_16661);
and U16974 (N_16974,N_16706,N_16664);
nor U16975 (N_16975,N_16514,N_16582);
nand U16976 (N_16976,N_16507,N_16586);
or U16977 (N_16977,N_16740,N_16533);
nor U16978 (N_16978,N_16581,N_16747);
xor U16979 (N_16979,N_16606,N_16708);
or U16980 (N_16980,N_16625,N_16558);
nand U16981 (N_16981,N_16575,N_16701);
nor U16982 (N_16982,N_16666,N_16610);
or U16983 (N_16983,N_16597,N_16641);
nand U16984 (N_16984,N_16544,N_16745);
nor U16985 (N_16985,N_16707,N_16733);
and U16986 (N_16986,N_16720,N_16746);
nand U16987 (N_16987,N_16589,N_16718);
or U16988 (N_16988,N_16536,N_16719);
nand U16989 (N_16989,N_16609,N_16689);
and U16990 (N_16990,N_16508,N_16628);
or U16991 (N_16991,N_16663,N_16717);
nand U16992 (N_16992,N_16733,N_16685);
nor U16993 (N_16993,N_16728,N_16716);
or U16994 (N_16994,N_16707,N_16577);
nor U16995 (N_16995,N_16606,N_16536);
or U16996 (N_16996,N_16697,N_16561);
or U16997 (N_16997,N_16607,N_16722);
nor U16998 (N_16998,N_16563,N_16540);
nand U16999 (N_16999,N_16531,N_16677);
nor U17000 (N_17000,N_16869,N_16821);
or U17001 (N_17001,N_16839,N_16940);
and U17002 (N_17002,N_16982,N_16899);
nor U17003 (N_17003,N_16956,N_16957);
and U17004 (N_17004,N_16919,N_16845);
and U17005 (N_17005,N_16758,N_16789);
nor U17006 (N_17006,N_16999,N_16939);
xor U17007 (N_17007,N_16829,N_16917);
nor U17008 (N_17008,N_16981,N_16912);
or U17009 (N_17009,N_16870,N_16882);
and U17010 (N_17010,N_16816,N_16763);
or U17011 (N_17011,N_16905,N_16926);
nor U17012 (N_17012,N_16799,N_16815);
nand U17013 (N_17013,N_16781,N_16925);
nand U17014 (N_17014,N_16798,N_16834);
or U17015 (N_17015,N_16947,N_16787);
xor U17016 (N_17016,N_16796,N_16934);
and U17017 (N_17017,N_16991,N_16773);
xnor U17018 (N_17018,N_16804,N_16970);
nand U17019 (N_17019,N_16813,N_16814);
and U17020 (N_17020,N_16861,N_16989);
xor U17021 (N_17021,N_16797,N_16988);
and U17022 (N_17022,N_16844,N_16846);
nor U17023 (N_17023,N_16780,N_16900);
nor U17024 (N_17024,N_16998,N_16768);
or U17025 (N_17025,N_16785,N_16774);
or U17026 (N_17026,N_16874,N_16995);
nand U17027 (N_17027,N_16800,N_16848);
or U17028 (N_17028,N_16907,N_16761);
xnor U17029 (N_17029,N_16860,N_16898);
nand U17030 (N_17030,N_16836,N_16765);
and U17031 (N_17031,N_16891,N_16941);
nand U17032 (N_17032,N_16817,N_16875);
or U17033 (N_17033,N_16772,N_16760);
nor U17034 (N_17034,N_16857,N_16904);
nand U17035 (N_17035,N_16918,N_16825);
nor U17036 (N_17036,N_16767,N_16868);
nand U17037 (N_17037,N_16858,N_16952);
xor U17038 (N_17038,N_16977,N_16983);
or U17039 (N_17039,N_16835,N_16928);
or U17040 (N_17040,N_16762,N_16873);
xnor U17041 (N_17041,N_16853,N_16888);
or U17042 (N_17042,N_16943,N_16872);
nor U17043 (N_17043,N_16842,N_16938);
nand U17044 (N_17044,N_16750,N_16927);
or U17045 (N_17045,N_16903,N_16808);
nor U17046 (N_17046,N_16771,N_16911);
xor U17047 (N_17047,N_16769,N_16795);
xor U17048 (N_17048,N_16838,N_16876);
nor U17049 (N_17049,N_16935,N_16830);
and U17050 (N_17050,N_16929,N_16997);
nand U17051 (N_17051,N_16883,N_16932);
nand U17052 (N_17052,N_16752,N_16862);
or U17053 (N_17053,N_16906,N_16824);
or U17054 (N_17054,N_16877,N_16881);
nand U17055 (N_17055,N_16859,N_16777);
nand U17056 (N_17056,N_16823,N_16992);
or U17057 (N_17057,N_16990,N_16851);
xor U17058 (N_17058,N_16948,N_16993);
nand U17059 (N_17059,N_16955,N_16812);
xor U17060 (N_17060,N_16822,N_16864);
nor U17061 (N_17061,N_16967,N_16942);
nand U17062 (N_17062,N_16978,N_16811);
nor U17063 (N_17063,N_16803,N_16893);
xor U17064 (N_17064,N_16764,N_16755);
and U17065 (N_17065,N_16962,N_16958);
nand U17066 (N_17066,N_16770,N_16890);
nand U17067 (N_17067,N_16827,N_16885);
or U17068 (N_17068,N_16775,N_16985);
nand U17069 (N_17069,N_16960,N_16969);
xnor U17070 (N_17070,N_16854,N_16757);
or U17071 (N_17071,N_16951,N_16984);
or U17072 (N_17072,N_16896,N_16884);
and U17073 (N_17073,N_16843,N_16784);
xor U17074 (N_17074,N_16828,N_16949);
nor U17075 (N_17075,N_16950,N_16913);
and U17076 (N_17076,N_16779,N_16986);
and U17077 (N_17077,N_16908,N_16878);
nor U17078 (N_17078,N_16887,N_16879);
xor U17079 (N_17079,N_16966,N_16886);
and U17080 (N_17080,N_16790,N_16863);
and U17081 (N_17081,N_16806,N_16915);
and U17082 (N_17082,N_16754,N_16959);
and U17083 (N_17083,N_16867,N_16902);
or U17084 (N_17084,N_16953,N_16792);
and U17085 (N_17085,N_16963,N_16756);
and U17086 (N_17086,N_16945,N_16837);
nor U17087 (N_17087,N_16818,N_16973);
or U17088 (N_17088,N_16996,N_16944);
xnor U17089 (N_17089,N_16849,N_16931);
or U17090 (N_17090,N_16880,N_16782);
or U17091 (N_17091,N_16791,N_16909);
nand U17092 (N_17092,N_16922,N_16847);
xnor U17093 (N_17093,N_16831,N_16961);
xor U17094 (N_17094,N_16980,N_16923);
and U17095 (N_17095,N_16820,N_16901);
nor U17096 (N_17096,N_16892,N_16766);
nor U17097 (N_17097,N_16924,N_16788);
and U17098 (N_17098,N_16783,N_16810);
xor U17099 (N_17099,N_16897,N_16759);
nand U17100 (N_17100,N_16976,N_16889);
xor U17101 (N_17101,N_16916,N_16937);
or U17102 (N_17102,N_16794,N_16965);
and U17103 (N_17103,N_16833,N_16850);
or U17104 (N_17104,N_16801,N_16974);
and U17105 (N_17105,N_16778,N_16793);
xnor U17106 (N_17106,N_16936,N_16921);
nand U17107 (N_17107,N_16753,N_16910);
nand U17108 (N_17108,N_16994,N_16914);
and U17109 (N_17109,N_16865,N_16871);
or U17110 (N_17110,N_16852,N_16751);
nor U17111 (N_17111,N_16840,N_16826);
nor U17112 (N_17112,N_16895,N_16979);
xor U17113 (N_17113,N_16954,N_16975);
nand U17114 (N_17114,N_16819,N_16946);
nand U17115 (N_17115,N_16933,N_16987);
and U17116 (N_17116,N_16930,N_16832);
nand U17117 (N_17117,N_16809,N_16972);
nand U17118 (N_17118,N_16807,N_16866);
and U17119 (N_17119,N_16968,N_16894);
xnor U17120 (N_17120,N_16920,N_16855);
and U17121 (N_17121,N_16964,N_16971);
nand U17122 (N_17122,N_16856,N_16805);
and U17123 (N_17123,N_16786,N_16802);
nor U17124 (N_17124,N_16776,N_16841);
or U17125 (N_17125,N_16957,N_16793);
and U17126 (N_17126,N_16924,N_16922);
nor U17127 (N_17127,N_16812,N_16935);
nand U17128 (N_17128,N_16846,N_16901);
nand U17129 (N_17129,N_16920,N_16754);
xnor U17130 (N_17130,N_16966,N_16868);
and U17131 (N_17131,N_16940,N_16753);
or U17132 (N_17132,N_16923,N_16751);
and U17133 (N_17133,N_16849,N_16979);
and U17134 (N_17134,N_16864,N_16969);
or U17135 (N_17135,N_16827,N_16750);
nor U17136 (N_17136,N_16900,N_16987);
or U17137 (N_17137,N_16844,N_16988);
and U17138 (N_17138,N_16990,N_16960);
xnor U17139 (N_17139,N_16757,N_16754);
or U17140 (N_17140,N_16868,N_16766);
or U17141 (N_17141,N_16766,N_16929);
or U17142 (N_17142,N_16853,N_16896);
xor U17143 (N_17143,N_16926,N_16917);
or U17144 (N_17144,N_16864,N_16983);
nand U17145 (N_17145,N_16764,N_16851);
and U17146 (N_17146,N_16972,N_16793);
nand U17147 (N_17147,N_16795,N_16911);
xor U17148 (N_17148,N_16898,N_16828);
nor U17149 (N_17149,N_16882,N_16840);
nand U17150 (N_17150,N_16894,N_16840);
nor U17151 (N_17151,N_16833,N_16870);
and U17152 (N_17152,N_16793,N_16880);
nand U17153 (N_17153,N_16909,N_16763);
nand U17154 (N_17154,N_16952,N_16822);
and U17155 (N_17155,N_16993,N_16959);
nand U17156 (N_17156,N_16994,N_16985);
nand U17157 (N_17157,N_16965,N_16834);
nor U17158 (N_17158,N_16835,N_16771);
xor U17159 (N_17159,N_16775,N_16800);
nor U17160 (N_17160,N_16787,N_16791);
or U17161 (N_17161,N_16997,N_16806);
xnor U17162 (N_17162,N_16852,N_16834);
or U17163 (N_17163,N_16927,N_16841);
nand U17164 (N_17164,N_16798,N_16962);
xor U17165 (N_17165,N_16942,N_16763);
and U17166 (N_17166,N_16848,N_16894);
nand U17167 (N_17167,N_16919,N_16891);
nor U17168 (N_17168,N_16925,N_16764);
or U17169 (N_17169,N_16901,N_16795);
and U17170 (N_17170,N_16904,N_16964);
xor U17171 (N_17171,N_16769,N_16755);
and U17172 (N_17172,N_16894,N_16867);
nand U17173 (N_17173,N_16918,N_16764);
nand U17174 (N_17174,N_16897,N_16771);
or U17175 (N_17175,N_16873,N_16968);
nand U17176 (N_17176,N_16905,N_16892);
and U17177 (N_17177,N_16976,N_16877);
or U17178 (N_17178,N_16804,N_16837);
xnor U17179 (N_17179,N_16915,N_16766);
nor U17180 (N_17180,N_16901,N_16859);
xnor U17181 (N_17181,N_16800,N_16774);
xor U17182 (N_17182,N_16867,N_16832);
or U17183 (N_17183,N_16796,N_16809);
nor U17184 (N_17184,N_16920,N_16861);
and U17185 (N_17185,N_16863,N_16761);
nor U17186 (N_17186,N_16753,N_16756);
or U17187 (N_17187,N_16821,N_16888);
nand U17188 (N_17188,N_16760,N_16838);
xnor U17189 (N_17189,N_16780,N_16889);
xnor U17190 (N_17190,N_16951,N_16820);
or U17191 (N_17191,N_16898,N_16853);
xor U17192 (N_17192,N_16966,N_16863);
nor U17193 (N_17193,N_16987,N_16935);
nor U17194 (N_17194,N_16967,N_16948);
nor U17195 (N_17195,N_16861,N_16808);
xor U17196 (N_17196,N_16798,N_16794);
nand U17197 (N_17197,N_16892,N_16961);
xnor U17198 (N_17198,N_16988,N_16800);
nor U17199 (N_17199,N_16883,N_16934);
nand U17200 (N_17200,N_16753,N_16848);
and U17201 (N_17201,N_16754,N_16880);
xor U17202 (N_17202,N_16932,N_16766);
or U17203 (N_17203,N_16998,N_16965);
nand U17204 (N_17204,N_16827,N_16803);
or U17205 (N_17205,N_16807,N_16754);
nor U17206 (N_17206,N_16838,N_16991);
and U17207 (N_17207,N_16853,N_16801);
xor U17208 (N_17208,N_16916,N_16771);
nor U17209 (N_17209,N_16794,N_16806);
xor U17210 (N_17210,N_16778,N_16764);
and U17211 (N_17211,N_16903,N_16847);
nor U17212 (N_17212,N_16964,N_16922);
and U17213 (N_17213,N_16812,N_16758);
and U17214 (N_17214,N_16863,N_16948);
nor U17215 (N_17215,N_16908,N_16851);
or U17216 (N_17216,N_16833,N_16810);
or U17217 (N_17217,N_16874,N_16755);
nor U17218 (N_17218,N_16754,N_16786);
and U17219 (N_17219,N_16883,N_16998);
and U17220 (N_17220,N_16788,N_16902);
xnor U17221 (N_17221,N_16883,N_16829);
or U17222 (N_17222,N_16971,N_16863);
and U17223 (N_17223,N_16941,N_16776);
nor U17224 (N_17224,N_16912,N_16766);
xor U17225 (N_17225,N_16887,N_16852);
and U17226 (N_17226,N_16806,N_16858);
or U17227 (N_17227,N_16927,N_16870);
or U17228 (N_17228,N_16858,N_16855);
xor U17229 (N_17229,N_16817,N_16764);
and U17230 (N_17230,N_16963,N_16871);
nand U17231 (N_17231,N_16983,N_16753);
xnor U17232 (N_17232,N_16885,N_16872);
nand U17233 (N_17233,N_16834,N_16992);
or U17234 (N_17234,N_16788,N_16918);
or U17235 (N_17235,N_16987,N_16861);
or U17236 (N_17236,N_16829,N_16775);
nand U17237 (N_17237,N_16789,N_16878);
nand U17238 (N_17238,N_16919,N_16944);
nand U17239 (N_17239,N_16960,N_16925);
or U17240 (N_17240,N_16802,N_16773);
nand U17241 (N_17241,N_16802,N_16967);
nor U17242 (N_17242,N_16917,N_16918);
nor U17243 (N_17243,N_16996,N_16993);
nand U17244 (N_17244,N_16873,N_16949);
nor U17245 (N_17245,N_16912,N_16915);
nor U17246 (N_17246,N_16861,N_16925);
nor U17247 (N_17247,N_16839,N_16750);
nand U17248 (N_17248,N_16772,N_16811);
nor U17249 (N_17249,N_16773,N_16949);
xnor U17250 (N_17250,N_17001,N_17012);
xor U17251 (N_17251,N_17241,N_17133);
nand U17252 (N_17252,N_17153,N_17206);
nand U17253 (N_17253,N_17178,N_17003);
nor U17254 (N_17254,N_17075,N_17142);
nor U17255 (N_17255,N_17188,N_17038);
or U17256 (N_17256,N_17169,N_17179);
nor U17257 (N_17257,N_17187,N_17223);
nor U17258 (N_17258,N_17067,N_17129);
or U17259 (N_17259,N_17202,N_17072);
nand U17260 (N_17260,N_17174,N_17068);
nor U17261 (N_17261,N_17196,N_17126);
nor U17262 (N_17262,N_17086,N_17105);
nand U17263 (N_17263,N_17077,N_17199);
nand U17264 (N_17264,N_17132,N_17236);
and U17265 (N_17265,N_17161,N_17229);
xor U17266 (N_17266,N_17249,N_17246);
nand U17267 (N_17267,N_17085,N_17143);
xor U17268 (N_17268,N_17002,N_17225);
and U17269 (N_17269,N_17213,N_17048);
and U17270 (N_17270,N_17017,N_17130);
or U17271 (N_17271,N_17124,N_17162);
xnor U17272 (N_17272,N_17192,N_17056);
nor U17273 (N_17273,N_17014,N_17207);
nand U17274 (N_17274,N_17109,N_17146);
or U17275 (N_17275,N_17237,N_17144);
nor U17276 (N_17276,N_17200,N_17028);
xor U17277 (N_17277,N_17217,N_17155);
nor U17278 (N_17278,N_17018,N_17000);
and U17279 (N_17279,N_17070,N_17083);
and U17280 (N_17280,N_17211,N_17089);
xnor U17281 (N_17281,N_17243,N_17231);
and U17282 (N_17282,N_17063,N_17159);
or U17283 (N_17283,N_17189,N_17244);
xor U17284 (N_17284,N_17203,N_17222);
xnor U17285 (N_17285,N_17088,N_17190);
nor U17286 (N_17286,N_17157,N_17005);
or U17287 (N_17287,N_17071,N_17108);
and U17288 (N_17288,N_17042,N_17052);
or U17289 (N_17289,N_17090,N_17212);
or U17290 (N_17290,N_17182,N_17170);
nand U17291 (N_17291,N_17198,N_17111);
nand U17292 (N_17292,N_17041,N_17066);
xnor U17293 (N_17293,N_17046,N_17093);
nor U17294 (N_17294,N_17228,N_17150);
nand U17295 (N_17295,N_17175,N_17009);
nand U17296 (N_17296,N_17127,N_17107);
nand U17297 (N_17297,N_17023,N_17034);
nor U17298 (N_17298,N_17011,N_17152);
and U17299 (N_17299,N_17224,N_17247);
nand U17300 (N_17300,N_17015,N_17233);
or U17301 (N_17301,N_17087,N_17043);
and U17302 (N_17302,N_17166,N_17047);
nand U17303 (N_17303,N_17186,N_17205);
or U17304 (N_17304,N_17025,N_17053);
nor U17305 (N_17305,N_17151,N_17135);
nand U17306 (N_17306,N_17221,N_17035);
xor U17307 (N_17307,N_17158,N_17030);
xor U17308 (N_17308,N_17026,N_17165);
xor U17309 (N_17309,N_17113,N_17197);
or U17310 (N_17310,N_17171,N_17149);
or U17311 (N_17311,N_17065,N_17214);
or U17312 (N_17312,N_17074,N_17095);
xnor U17313 (N_17313,N_17008,N_17238);
nor U17314 (N_17314,N_17115,N_17116);
xor U17315 (N_17315,N_17173,N_17110);
nand U17316 (N_17316,N_17004,N_17091);
or U17317 (N_17317,N_17010,N_17201);
or U17318 (N_17318,N_17084,N_17194);
xor U17319 (N_17319,N_17069,N_17117);
and U17320 (N_17320,N_17248,N_17104);
nor U17321 (N_17321,N_17123,N_17078);
or U17322 (N_17322,N_17181,N_17195);
or U17323 (N_17323,N_17131,N_17007);
xor U17324 (N_17324,N_17059,N_17044);
xnor U17325 (N_17325,N_17096,N_17050);
or U17326 (N_17326,N_17029,N_17031);
or U17327 (N_17327,N_17128,N_17125);
and U17328 (N_17328,N_17230,N_17138);
and U17329 (N_17329,N_17098,N_17032);
xor U17330 (N_17330,N_17148,N_17055);
and U17331 (N_17331,N_17185,N_17081);
nor U17332 (N_17332,N_17016,N_17076);
xnor U17333 (N_17333,N_17177,N_17218);
nand U17334 (N_17334,N_17082,N_17168);
xor U17335 (N_17335,N_17037,N_17092);
xnor U17336 (N_17336,N_17019,N_17136);
nor U17337 (N_17337,N_17013,N_17054);
xor U17338 (N_17338,N_17160,N_17242);
or U17339 (N_17339,N_17097,N_17167);
and U17340 (N_17340,N_17040,N_17172);
nand U17341 (N_17341,N_17114,N_17139);
xor U17342 (N_17342,N_17220,N_17102);
and U17343 (N_17343,N_17079,N_17141);
nand U17344 (N_17344,N_17184,N_17122);
or U17345 (N_17345,N_17232,N_17180);
xor U17346 (N_17346,N_17210,N_17051);
nor U17347 (N_17347,N_17036,N_17020);
xor U17348 (N_17348,N_17235,N_17103);
and U17349 (N_17349,N_17120,N_17024);
or U17350 (N_17350,N_17080,N_17064);
and U17351 (N_17351,N_17073,N_17154);
nand U17352 (N_17352,N_17156,N_17006);
or U17353 (N_17353,N_17191,N_17240);
or U17354 (N_17354,N_17022,N_17208);
xor U17355 (N_17355,N_17215,N_17245);
xnor U17356 (N_17356,N_17062,N_17039);
and U17357 (N_17357,N_17140,N_17060);
xnor U17358 (N_17358,N_17147,N_17121);
nand U17359 (N_17359,N_17163,N_17227);
nor U17360 (N_17360,N_17099,N_17134);
nand U17361 (N_17361,N_17204,N_17119);
nor U17362 (N_17362,N_17137,N_17061);
nor U17363 (N_17363,N_17164,N_17112);
and U17364 (N_17364,N_17058,N_17216);
nor U17365 (N_17365,N_17118,N_17057);
nand U17366 (N_17366,N_17226,N_17027);
and U17367 (N_17367,N_17045,N_17209);
and U17368 (N_17368,N_17234,N_17106);
and U17369 (N_17369,N_17101,N_17145);
or U17370 (N_17370,N_17176,N_17033);
or U17371 (N_17371,N_17239,N_17094);
nand U17372 (N_17372,N_17219,N_17049);
and U17373 (N_17373,N_17100,N_17193);
xor U17374 (N_17374,N_17183,N_17021);
and U17375 (N_17375,N_17154,N_17223);
or U17376 (N_17376,N_17187,N_17174);
and U17377 (N_17377,N_17159,N_17068);
nor U17378 (N_17378,N_17158,N_17064);
and U17379 (N_17379,N_17151,N_17233);
nand U17380 (N_17380,N_17196,N_17247);
xor U17381 (N_17381,N_17119,N_17228);
nor U17382 (N_17382,N_17119,N_17194);
and U17383 (N_17383,N_17101,N_17144);
or U17384 (N_17384,N_17152,N_17138);
and U17385 (N_17385,N_17065,N_17223);
or U17386 (N_17386,N_17161,N_17048);
nand U17387 (N_17387,N_17170,N_17044);
and U17388 (N_17388,N_17170,N_17029);
or U17389 (N_17389,N_17223,N_17129);
and U17390 (N_17390,N_17201,N_17169);
xor U17391 (N_17391,N_17210,N_17010);
or U17392 (N_17392,N_17100,N_17102);
nor U17393 (N_17393,N_17183,N_17075);
xnor U17394 (N_17394,N_17016,N_17246);
nor U17395 (N_17395,N_17012,N_17101);
nor U17396 (N_17396,N_17230,N_17180);
and U17397 (N_17397,N_17023,N_17067);
nor U17398 (N_17398,N_17078,N_17202);
or U17399 (N_17399,N_17242,N_17108);
or U17400 (N_17400,N_17178,N_17014);
xnor U17401 (N_17401,N_17127,N_17234);
nor U17402 (N_17402,N_17207,N_17208);
xor U17403 (N_17403,N_17065,N_17173);
nand U17404 (N_17404,N_17139,N_17047);
nor U17405 (N_17405,N_17100,N_17060);
xnor U17406 (N_17406,N_17229,N_17085);
nor U17407 (N_17407,N_17002,N_17148);
xnor U17408 (N_17408,N_17189,N_17171);
and U17409 (N_17409,N_17173,N_17084);
or U17410 (N_17410,N_17102,N_17161);
or U17411 (N_17411,N_17121,N_17129);
nor U17412 (N_17412,N_17186,N_17059);
and U17413 (N_17413,N_17190,N_17199);
or U17414 (N_17414,N_17128,N_17170);
nand U17415 (N_17415,N_17033,N_17222);
nand U17416 (N_17416,N_17087,N_17100);
and U17417 (N_17417,N_17228,N_17177);
nand U17418 (N_17418,N_17072,N_17064);
and U17419 (N_17419,N_17065,N_17247);
nand U17420 (N_17420,N_17118,N_17248);
xor U17421 (N_17421,N_17047,N_17188);
and U17422 (N_17422,N_17099,N_17132);
and U17423 (N_17423,N_17123,N_17243);
xnor U17424 (N_17424,N_17173,N_17217);
nand U17425 (N_17425,N_17100,N_17225);
and U17426 (N_17426,N_17201,N_17138);
and U17427 (N_17427,N_17028,N_17017);
and U17428 (N_17428,N_17114,N_17243);
nand U17429 (N_17429,N_17011,N_17067);
or U17430 (N_17430,N_17034,N_17175);
or U17431 (N_17431,N_17054,N_17019);
nor U17432 (N_17432,N_17175,N_17201);
and U17433 (N_17433,N_17082,N_17115);
nand U17434 (N_17434,N_17072,N_17029);
nand U17435 (N_17435,N_17153,N_17223);
nand U17436 (N_17436,N_17124,N_17061);
and U17437 (N_17437,N_17145,N_17200);
and U17438 (N_17438,N_17092,N_17221);
or U17439 (N_17439,N_17093,N_17057);
nor U17440 (N_17440,N_17030,N_17155);
and U17441 (N_17441,N_17032,N_17095);
or U17442 (N_17442,N_17091,N_17031);
xor U17443 (N_17443,N_17084,N_17246);
and U17444 (N_17444,N_17199,N_17124);
and U17445 (N_17445,N_17033,N_17096);
nand U17446 (N_17446,N_17167,N_17241);
nor U17447 (N_17447,N_17071,N_17115);
nand U17448 (N_17448,N_17056,N_17220);
or U17449 (N_17449,N_17192,N_17049);
or U17450 (N_17450,N_17039,N_17158);
or U17451 (N_17451,N_17176,N_17121);
or U17452 (N_17452,N_17199,N_17101);
xor U17453 (N_17453,N_17154,N_17115);
nor U17454 (N_17454,N_17005,N_17143);
or U17455 (N_17455,N_17000,N_17089);
or U17456 (N_17456,N_17092,N_17125);
and U17457 (N_17457,N_17008,N_17168);
nand U17458 (N_17458,N_17220,N_17223);
or U17459 (N_17459,N_17068,N_17152);
nand U17460 (N_17460,N_17133,N_17066);
xnor U17461 (N_17461,N_17054,N_17026);
or U17462 (N_17462,N_17224,N_17219);
nand U17463 (N_17463,N_17098,N_17215);
xor U17464 (N_17464,N_17225,N_17094);
nor U17465 (N_17465,N_17068,N_17035);
nand U17466 (N_17466,N_17211,N_17013);
nor U17467 (N_17467,N_17013,N_17241);
nand U17468 (N_17468,N_17136,N_17137);
nand U17469 (N_17469,N_17052,N_17017);
or U17470 (N_17470,N_17145,N_17056);
and U17471 (N_17471,N_17069,N_17044);
xor U17472 (N_17472,N_17092,N_17072);
or U17473 (N_17473,N_17240,N_17178);
nand U17474 (N_17474,N_17078,N_17238);
and U17475 (N_17475,N_17003,N_17206);
and U17476 (N_17476,N_17067,N_17121);
nor U17477 (N_17477,N_17128,N_17092);
or U17478 (N_17478,N_17121,N_17010);
and U17479 (N_17479,N_17081,N_17059);
xor U17480 (N_17480,N_17089,N_17178);
or U17481 (N_17481,N_17140,N_17055);
xnor U17482 (N_17482,N_17033,N_17193);
xor U17483 (N_17483,N_17059,N_17231);
nand U17484 (N_17484,N_17023,N_17043);
nor U17485 (N_17485,N_17014,N_17118);
and U17486 (N_17486,N_17186,N_17069);
nor U17487 (N_17487,N_17242,N_17244);
and U17488 (N_17488,N_17216,N_17068);
xnor U17489 (N_17489,N_17202,N_17004);
and U17490 (N_17490,N_17216,N_17161);
nor U17491 (N_17491,N_17140,N_17205);
and U17492 (N_17492,N_17225,N_17197);
or U17493 (N_17493,N_17189,N_17174);
nand U17494 (N_17494,N_17034,N_17086);
xor U17495 (N_17495,N_17128,N_17093);
and U17496 (N_17496,N_17095,N_17110);
nor U17497 (N_17497,N_17186,N_17176);
nor U17498 (N_17498,N_17219,N_17191);
nor U17499 (N_17499,N_17042,N_17173);
xor U17500 (N_17500,N_17412,N_17294);
nor U17501 (N_17501,N_17442,N_17473);
nand U17502 (N_17502,N_17403,N_17401);
and U17503 (N_17503,N_17377,N_17288);
nand U17504 (N_17504,N_17475,N_17446);
nand U17505 (N_17505,N_17367,N_17451);
and U17506 (N_17506,N_17350,N_17281);
nand U17507 (N_17507,N_17386,N_17323);
xnor U17508 (N_17508,N_17440,N_17466);
xnor U17509 (N_17509,N_17380,N_17424);
or U17510 (N_17510,N_17351,N_17317);
and U17511 (N_17511,N_17303,N_17375);
xnor U17512 (N_17512,N_17461,N_17333);
or U17513 (N_17513,N_17346,N_17459);
nor U17514 (N_17514,N_17467,N_17425);
xnor U17515 (N_17515,N_17404,N_17414);
nor U17516 (N_17516,N_17339,N_17429);
xor U17517 (N_17517,N_17447,N_17393);
or U17518 (N_17518,N_17273,N_17343);
nor U17519 (N_17519,N_17392,N_17252);
or U17520 (N_17520,N_17301,N_17376);
xor U17521 (N_17521,N_17251,N_17371);
xor U17522 (N_17522,N_17432,N_17335);
xor U17523 (N_17523,N_17308,N_17278);
nand U17524 (N_17524,N_17313,N_17444);
xnor U17525 (N_17525,N_17280,N_17452);
nand U17526 (N_17526,N_17457,N_17314);
nor U17527 (N_17527,N_17357,N_17291);
nor U17528 (N_17528,N_17274,N_17302);
or U17529 (N_17529,N_17262,N_17470);
nor U17530 (N_17530,N_17259,N_17332);
xor U17531 (N_17531,N_17276,N_17327);
nor U17532 (N_17532,N_17315,N_17279);
and U17533 (N_17533,N_17415,N_17304);
or U17534 (N_17534,N_17493,N_17477);
nor U17535 (N_17535,N_17434,N_17471);
and U17536 (N_17536,N_17311,N_17468);
and U17537 (N_17537,N_17390,N_17497);
nand U17538 (N_17538,N_17257,N_17363);
nor U17539 (N_17539,N_17491,N_17287);
nand U17540 (N_17540,N_17438,N_17494);
or U17541 (N_17541,N_17366,N_17484);
nand U17542 (N_17542,N_17398,N_17423);
nor U17543 (N_17543,N_17261,N_17275);
or U17544 (N_17544,N_17486,N_17364);
nor U17545 (N_17545,N_17430,N_17448);
or U17546 (N_17546,N_17487,N_17331);
nor U17547 (N_17547,N_17495,N_17410);
or U17548 (N_17548,N_17458,N_17334);
and U17549 (N_17549,N_17450,N_17496);
xor U17550 (N_17550,N_17454,N_17396);
or U17551 (N_17551,N_17312,N_17298);
xnor U17552 (N_17552,N_17316,N_17268);
nor U17553 (N_17553,N_17289,N_17255);
xor U17554 (N_17554,N_17329,N_17359);
and U17555 (N_17555,N_17365,N_17420);
and U17556 (N_17556,N_17480,N_17347);
nor U17557 (N_17557,N_17264,N_17277);
nand U17558 (N_17558,N_17336,N_17483);
and U17559 (N_17559,N_17307,N_17453);
or U17560 (N_17560,N_17270,N_17456);
xnor U17561 (N_17561,N_17338,N_17319);
nand U17562 (N_17562,N_17265,N_17370);
and U17563 (N_17563,N_17260,N_17330);
nor U17564 (N_17564,N_17476,N_17326);
xor U17565 (N_17565,N_17437,N_17465);
xnor U17566 (N_17566,N_17431,N_17387);
nand U17567 (N_17567,N_17389,N_17292);
nand U17568 (N_17568,N_17356,N_17407);
nor U17569 (N_17569,N_17299,N_17488);
and U17570 (N_17570,N_17253,N_17306);
or U17571 (N_17571,N_17428,N_17406);
nor U17572 (N_17572,N_17340,N_17374);
nor U17573 (N_17573,N_17472,N_17481);
and U17574 (N_17574,N_17282,N_17441);
nor U17575 (N_17575,N_17310,N_17272);
nand U17576 (N_17576,N_17328,N_17382);
nand U17577 (N_17577,N_17271,N_17394);
or U17578 (N_17578,N_17402,N_17489);
nand U17579 (N_17579,N_17449,N_17296);
or U17580 (N_17580,N_17325,N_17416);
or U17581 (N_17581,N_17293,N_17354);
or U17582 (N_17582,N_17464,N_17254);
or U17583 (N_17583,N_17388,N_17352);
and U17584 (N_17584,N_17479,N_17405);
xor U17585 (N_17585,N_17384,N_17353);
nand U17586 (N_17586,N_17421,N_17417);
nand U17587 (N_17587,N_17320,N_17284);
xor U17588 (N_17588,N_17283,N_17318);
and U17589 (N_17589,N_17385,N_17348);
nand U17590 (N_17590,N_17263,N_17395);
nand U17591 (N_17591,N_17460,N_17290);
and U17592 (N_17592,N_17397,N_17372);
xnor U17593 (N_17593,N_17455,N_17368);
or U17594 (N_17594,N_17433,N_17345);
or U17595 (N_17595,N_17443,N_17400);
or U17596 (N_17596,N_17342,N_17435);
xnor U17597 (N_17597,N_17408,N_17482);
nor U17598 (N_17598,N_17381,N_17391);
or U17599 (N_17599,N_17485,N_17469);
nor U17600 (N_17600,N_17349,N_17399);
and U17601 (N_17601,N_17498,N_17286);
and U17602 (N_17602,N_17358,N_17355);
nand U17603 (N_17603,N_17250,N_17285);
nand U17604 (N_17604,N_17341,N_17427);
or U17605 (N_17605,N_17383,N_17360);
nor U17606 (N_17606,N_17300,N_17422);
or U17607 (N_17607,N_17321,N_17409);
xnor U17608 (N_17608,N_17379,N_17256);
and U17609 (N_17609,N_17413,N_17474);
and U17610 (N_17610,N_17478,N_17362);
nor U17611 (N_17611,N_17462,N_17269);
nor U17612 (N_17612,N_17499,N_17337);
xnor U17613 (N_17613,N_17411,N_17426);
and U17614 (N_17614,N_17418,N_17463);
xor U17615 (N_17615,N_17295,N_17258);
and U17616 (N_17616,N_17436,N_17267);
nor U17617 (N_17617,N_17305,N_17361);
or U17618 (N_17618,N_17492,N_17369);
and U17619 (N_17619,N_17373,N_17378);
or U17620 (N_17620,N_17322,N_17324);
xnor U17621 (N_17621,N_17490,N_17445);
xor U17622 (N_17622,N_17419,N_17266);
nand U17623 (N_17623,N_17309,N_17439);
xor U17624 (N_17624,N_17297,N_17344);
nand U17625 (N_17625,N_17299,N_17441);
nor U17626 (N_17626,N_17340,N_17479);
xor U17627 (N_17627,N_17470,N_17409);
xor U17628 (N_17628,N_17376,N_17331);
xnor U17629 (N_17629,N_17368,N_17352);
xor U17630 (N_17630,N_17414,N_17292);
nor U17631 (N_17631,N_17271,N_17344);
xnor U17632 (N_17632,N_17370,N_17383);
and U17633 (N_17633,N_17281,N_17309);
nand U17634 (N_17634,N_17288,N_17427);
nor U17635 (N_17635,N_17436,N_17438);
nand U17636 (N_17636,N_17402,N_17430);
nor U17637 (N_17637,N_17381,N_17368);
xnor U17638 (N_17638,N_17252,N_17286);
or U17639 (N_17639,N_17402,N_17470);
nor U17640 (N_17640,N_17427,N_17271);
or U17641 (N_17641,N_17255,N_17333);
or U17642 (N_17642,N_17255,N_17331);
nand U17643 (N_17643,N_17255,N_17459);
or U17644 (N_17644,N_17360,N_17468);
xor U17645 (N_17645,N_17301,N_17488);
or U17646 (N_17646,N_17375,N_17284);
and U17647 (N_17647,N_17348,N_17354);
or U17648 (N_17648,N_17289,N_17421);
or U17649 (N_17649,N_17355,N_17420);
nor U17650 (N_17650,N_17330,N_17345);
nor U17651 (N_17651,N_17414,N_17470);
nor U17652 (N_17652,N_17358,N_17396);
xnor U17653 (N_17653,N_17456,N_17407);
xor U17654 (N_17654,N_17251,N_17260);
or U17655 (N_17655,N_17388,N_17494);
or U17656 (N_17656,N_17270,N_17268);
or U17657 (N_17657,N_17267,N_17292);
or U17658 (N_17658,N_17387,N_17458);
nand U17659 (N_17659,N_17317,N_17324);
xnor U17660 (N_17660,N_17320,N_17453);
and U17661 (N_17661,N_17318,N_17364);
nand U17662 (N_17662,N_17377,N_17273);
nor U17663 (N_17663,N_17433,N_17385);
and U17664 (N_17664,N_17252,N_17411);
or U17665 (N_17665,N_17254,N_17392);
nor U17666 (N_17666,N_17271,N_17415);
nand U17667 (N_17667,N_17383,N_17457);
and U17668 (N_17668,N_17475,N_17277);
or U17669 (N_17669,N_17374,N_17345);
nand U17670 (N_17670,N_17375,N_17443);
and U17671 (N_17671,N_17298,N_17396);
or U17672 (N_17672,N_17423,N_17459);
nand U17673 (N_17673,N_17302,N_17404);
nor U17674 (N_17674,N_17433,N_17326);
and U17675 (N_17675,N_17254,N_17288);
nor U17676 (N_17676,N_17416,N_17306);
nand U17677 (N_17677,N_17470,N_17475);
nand U17678 (N_17678,N_17418,N_17483);
nor U17679 (N_17679,N_17301,N_17474);
and U17680 (N_17680,N_17371,N_17293);
nand U17681 (N_17681,N_17267,N_17486);
or U17682 (N_17682,N_17353,N_17498);
or U17683 (N_17683,N_17465,N_17447);
nor U17684 (N_17684,N_17395,N_17309);
and U17685 (N_17685,N_17431,N_17487);
nand U17686 (N_17686,N_17486,N_17444);
nor U17687 (N_17687,N_17284,N_17426);
and U17688 (N_17688,N_17434,N_17393);
and U17689 (N_17689,N_17326,N_17447);
nor U17690 (N_17690,N_17474,N_17257);
nand U17691 (N_17691,N_17358,N_17345);
and U17692 (N_17692,N_17482,N_17285);
and U17693 (N_17693,N_17257,N_17250);
xnor U17694 (N_17694,N_17269,N_17254);
nor U17695 (N_17695,N_17260,N_17480);
or U17696 (N_17696,N_17495,N_17254);
and U17697 (N_17697,N_17259,N_17357);
or U17698 (N_17698,N_17438,N_17264);
nand U17699 (N_17699,N_17274,N_17451);
xnor U17700 (N_17700,N_17487,N_17334);
xor U17701 (N_17701,N_17439,N_17311);
nand U17702 (N_17702,N_17290,N_17351);
nand U17703 (N_17703,N_17346,N_17393);
and U17704 (N_17704,N_17410,N_17494);
or U17705 (N_17705,N_17334,N_17299);
or U17706 (N_17706,N_17426,N_17492);
or U17707 (N_17707,N_17420,N_17367);
xor U17708 (N_17708,N_17464,N_17369);
or U17709 (N_17709,N_17404,N_17427);
or U17710 (N_17710,N_17330,N_17255);
and U17711 (N_17711,N_17298,N_17402);
or U17712 (N_17712,N_17293,N_17415);
nor U17713 (N_17713,N_17274,N_17403);
and U17714 (N_17714,N_17469,N_17391);
nor U17715 (N_17715,N_17351,N_17321);
xor U17716 (N_17716,N_17453,N_17448);
xor U17717 (N_17717,N_17336,N_17489);
nor U17718 (N_17718,N_17367,N_17421);
nand U17719 (N_17719,N_17318,N_17407);
xor U17720 (N_17720,N_17435,N_17388);
nand U17721 (N_17721,N_17342,N_17494);
xor U17722 (N_17722,N_17448,N_17319);
or U17723 (N_17723,N_17274,N_17433);
or U17724 (N_17724,N_17372,N_17365);
or U17725 (N_17725,N_17332,N_17367);
or U17726 (N_17726,N_17381,N_17453);
and U17727 (N_17727,N_17254,N_17253);
nor U17728 (N_17728,N_17468,N_17374);
xnor U17729 (N_17729,N_17473,N_17386);
nor U17730 (N_17730,N_17281,N_17361);
or U17731 (N_17731,N_17298,N_17410);
nand U17732 (N_17732,N_17464,N_17445);
or U17733 (N_17733,N_17457,N_17466);
or U17734 (N_17734,N_17274,N_17468);
nand U17735 (N_17735,N_17286,N_17465);
nor U17736 (N_17736,N_17265,N_17325);
and U17737 (N_17737,N_17276,N_17384);
xnor U17738 (N_17738,N_17353,N_17431);
nand U17739 (N_17739,N_17428,N_17351);
xor U17740 (N_17740,N_17370,N_17487);
nor U17741 (N_17741,N_17405,N_17491);
nor U17742 (N_17742,N_17499,N_17368);
nand U17743 (N_17743,N_17450,N_17398);
nor U17744 (N_17744,N_17338,N_17425);
nand U17745 (N_17745,N_17470,N_17352);
and U17746 (N_17746,N_17375,N_17278);
or U17747 (N_17747,N_17440,N_17281);
xor U17748 (N_17748,N_17254,N_17266);
or U17749 (N_17749,N_17282,N_17308);
or U17750 (N_17750,N_17537,N_17520);
and U17751 (N_17751,N_17739,N_17550);
and U17752 (N_17752,N_17710,N_17688);
nand U17753 (N_17753,N_17561,N_17672);
or U17754 (N_17754,N_17586,N_17556);
xnor U17755 (N_17755,N_17518,N_17746);
nand U17756 (N_17756,N_17660,N_17535);
and U17757 (N_17757,N_17713,N_17639);
and U17758 (N_17758,N_17645,N_17720);
xnor U17759 (N_17759,N_17597,N_17719);
nor U17760 (N_17760,N_17698,N_17749);
nor U17761 (N_17761,N_17664,N_17678);
nor U17762 (N_17762,N_17542,N_17722);
xnor U17763 (N_17763,N_17618,N_17654);
nor U17764 (N_17764,N_17551,N_17658);
nand U17765 (N_17765,N_17743,N_17516);
or U17766 (N_17766,N_17718,N_17549);
nand U17767 (N_17767,N_17711,N_17669);
or U17768 (N_17768,N_17604,N_17500);
or U17769 (N_17769,N_17595,N_17620);
xor U17770 (N_17770,N_17708,N_17745);
nor U17771 (N_17771,N_17584,N_17534);
or U17772 (N_17772,N_17650,N_17522);
nor U17773 (N_17773,N_17632,N_17587);
nor U17774 (N_17774,N_17704,N_17616);
and U17775 (N_17775,N_17526,N_17544);
xor U17776 (N_17776,N_17619,N_17610);
and U17777 (N_17777,N_17572,N_17701);
nor U17778 (N_17778,N_17726,N_17621);
nor U17779 (N_17779,N_17571,N_17733);
nor U17780 (N_17780,N_17643,N_17747);
or U17781 (N_17781,N_17657,N_17625);
nand U17782 (N_17782,N_17569,N_17504);
or U17783 (N_17783,N_17581,N_17730);
nor U17784 (N_17784,N_17729,N_17666);
nor U17785 (N_17785,N_17690,N_17721);
or U17786 (N_17786,N_17646,N_17540);
or U17787 (N_17787,N_17692,N_17714);
nand U17788 (N_17788,N_17612,N_17681);
and U17789 (N_17789,N_17555,N_17695);
or U17790 (N_17790,N_17661,N_17628);
nand U17791 (N_17791,N_17510,N_17683);
and U17792 (N_17792,N_17501,N_17741);
or U17793 (N_17793,N_17562,N_17694);
or U17794 (N_17794,N_17583,N_17573);
xor U17795 (N_17795,N_17656,N_17738);
xnor U17796 (N_17796,N_17608,N_17557);
nand U17797 (N_17797,N_17630,N_17699);
or U17798 (N_17798,N_17575,N_17631);
or U17799 (N_17799,N_17568,N_17731);
and U17800 (N_17800,N_17603,N_17601);
and U17801 (N_17801,N_17653,N_17700);
nand U17802 (N_17802,N_17696,N_17665);
xor U17803 (N_17803,N_17528,N_17543);
or U17804 (N_17804,N_17706,N_17592);
xnor U17805 (N_17805,N_17709,N_17578);
xnor U17806 (N_17806,N_17502,N_17512);
nor U17807 (N_17807,N_17716,N_17671);
xor U17808 (N_17808,N_17565,N_17647);
nand U17809 (N_17809,N_17717,N_17547);
xnor U17810 (N_17810,N_17634,N_17558);
nor U17811 (N_17811,N_17633,N_17651);
and U17812 (N_17812,N_17574,N_17677);
and U17813 (N_17813,N_17570,N_17675);
nor U17814 (N_17814,N_17517,N_17611);
and U17815 (N_17815,N_17590,N_17723);
xnor U17816 (N_17816,N_17742,N_17703);
and U17817 (N_17817,N_17652,N_17613);
xnor U17818 (N_17818,N_17624,N_17734);
nor U17819 (N_17819,N_17546,N_17670);
and U17820 (N_17820,N_17629,N_17640);
xnor U17821 (N_17821,N_17589,N_17566);
nor U17822 (N_17822,N_17591,N_17508);
or U17823 (N_17823,N_17614,N_17593);
nor U17824 (N_17824,N_17617,N_17638);
or U17825 (N_17825,N_17530,N_17539);
nand U17826 (N_17826,N_17644,N_17637);
nand U17827 (N_17827,N_17523,N_17615);
xnor U17828 (N_17828,N_17564,N_17737);
and U17829 (N_17829,N_17588,N_17548);
or U17830 (N_17830,N_17511,N_17724);
nor U17831 (N_17831,N_17662,N_17748);
nand U17832 (N_17832,N_17626,N_17663);
xnor U17833 (N_17833,N_17538,N_17689);
nand U17834 (N_17834,N_17527,N_17648);
or U17835 (N_17835,N_17679,N_17513);
and U17836 (N_17836,N_17505,N_17684);
xnor U17837 (N_17837,N_17641,N_17707);
xnor U17838 (N_17838,N_17580,N_17607);
and U17839 (N_17839,N_17507,N_17554);
or U17840 (N_17840,N_17667,N_17712);
or U17841 (N_17841,N_17577,N_17668);
or U17842 (N_17842,N_17552,N_17725);
nor U17843 (N_17843,N_17691,N_17585);
nand U17844 (N_17844,N_17627,N_17596);
xor U17845 (N_17845,N_17736,N_17576);
nand U17846 (N_17846,N_17553,N_17519);
and U17847 (N_17847,N_17702,N_17693);
nand U17848 (N_17848,N_17655,N_17529);
and U17849 (N_17849,N_17659,N_17735);
nor U17850 (N_17850,N_17649,N_17525);
xnor U17851 (N_17851,N_17536,N_17533);
nor U17852 (N_17852,N_17744,N_17635);
xor U17853 (N_17853,N_17642,N_17541);
xnor U17854 (N_17854,N_17532,N_17686);
or U17855 (N_17855,N_17685,N_17622);
or U17856 (N_17856,N_17524,N_17506);
nand U17857 (N_17857,N_17740,N_17599);
nand U17858 (N_17858,N_17567,N_17594);
xnor U17859 (N_17859,N_17727,N_17676);
or U17860 (N_17860,N_17598,N_17715);
nor U17861 (N_17861,N_17531,N_17606);
xnor U17862 (N_17862,N_17560,N_17563);
xor U17863 (N_17863,N_17521,N_17687);
nand U17864 (N_17864,N_17732,N_17602);
xor U17865 (N_17865,N_17545,N_17514);
or U17866 (N_17866,N_17559,N_17579);
xnor U17867 (N_17867,N_17705,N_17609);
nand U17868 (N_17868,N_17680,N_17503);
xor U17869 (N_17869,N_17605,N_17623);
nand U17870 (N_17870,N_17582,N_17509);
nor U17871 (N_17871,N_17682,N_17728);
xor U17872 (N_17872,N_17600,N_17674);
nor U17873 (N_17873,N_17697,N_17515);
nand U17874 (N_17874,N_17673,N_17636);
and U17875 (N_17875,N_17534,N_17518);
xor U17876 (N_17876,N_17736,N_17719);
or U17877 (N_17877,N_17636,N_17607);
and U17878 (N_17878,N_17692,N_17628);
xor U17879 (N_17879,N_17606,N_17609);
and U17880 (N_17880,N_17562,N_17591);
and U17881 (N_17881,N_17740,N_17678);
nand U17882 (N_17882,N_17686,N_17691);
nor U17883 (N_17883,N_17523,N_17732);
nand U17884 (N_17884,N_17501,N_17614);
or U17885 (N_17885,N_17676,N_17573);
and U17886 (N_17886,N_17511,N_17594);
and U17887 (N_17887,N_17691,N_17726);
or U17888 (N_17888,N_17654,N_17581);
or U17889 (N_17889,N_17645,N_17662);
or U17890 (N_17890,N_17585,N_17746);
or U17891 (N_17891,N_17749,N_17571);
and U17892 (N_17892,N_17590,N_17567);
nand U17893 (N_17893,N_17681,N_17629);
or U17894 (N_17894,N_17598,N_17522);
and U17895 (N_17895,N_17684,N_17662);
nor U17896 (N_17896,N_17738,N_17727);
nor U17897 (N_17897,N_17736,N_17555);
nor U17898 (N_17898,N_17709,N_17658);
nand U17899 (N_17899,N_17511,N_17645);
xor U17900 (N_17900,N_17591,N_17627);
or U17901 (N_17901,N_17584,N_17657);
and U17902 (N_17902,N_17746,N_17517);
xor U17903 (N_17903,N_17599,N_17631);
or U17904 (N_17904,N_17531,N_17553);
xor U17905 (N_17905,N_17519,N_17676);
nand U17906 (N_17906,N_17547,N_17556);
and U17907 (N_17907,N_17704,N_17599);
or U17908 (N_17908,N_17500,N_17650);
and U17909 (N_17909,N_17647,N_17586);
xor U17910 (N_17910,N_17719,N_17610);
xnor U17911 (N_17911,N_17597,N_17537);
or U17912 (N_17912,N_17671,N_17557);
and U17913 (N_17913,N_17511,N_17703);
xor U17914 (N_17914,N_17690,N_17717);
xnor U17915 (N_17915,N_17525,N_17695);
xnor U17916 (N_17916,N_17732,N_17595);
xnor U17917 (N_17917,N_17571,N_17535);
nand U17918 (N_17918,N_17625,N_17638);
or U17919 (N_17919,N_17649,N_17719);
nand U17920 (N_17920,N_17726,N_17714);
xnor U17921 (N_17921,N_17577,N_17506);
or U17922 (N_17922,N_17564,N_17746);
nand U17923 (N_17923,N_17741,N_17652);
or U17924 (N_17924,N_17669,N_17697);
nor U17925 (N_17925,N_17614,N_17514);
or U17926 (N_17926,N_17729,N_17698);
or U17927 (N_17927,N_17629,N_17673);
and U17928 (N_17928,N_17740,N_17590);
nor U17929 (N_17929,N_17580,N_17678);
nand U17930 (N_17930,N_17707,N_17655);
or U17931 (N_17931,N_17556,N_17673);
nand U17932 (N_17932,N_17647,N_17706);
xor U17933 (N_17933,N_17624,N_17517);
nor U17934 (N_17934,N_17625,N_17644);
xnor U17935 (N_17935,N_17565,N_17673);
nor U17936 (N_17936,N_17657,N_17546);
xor U17937 (N_17937,N_17586,N_17729);
xor U17938 (N_17938,N_17561,N_17633);
xor U17939 (N_17939,N_17506,N_17522);
xnor U17940 (N_17940,N_17748,N_17583);
and U17941 (N_17941,N_17651,N_17695);
or U17942 (N_17942,N_17594,N_17548);
xor U17943 (N_17943,N_17612,N_17592);
nor U17944 (N_17944,N_17603,N_17628);
xnor U17945 (N_17945,N_17581,N_17713);
xor U17946 (N_17946,N_17732,N_17537);
and U17947 (N_17947,N_17745,N_17722);
or U17948 (N_17948,N_17617,N_17554);
or U17949 (N_17949,N_17637,N_17724);
nor U17950 (N_17950,N_17527,N_17503);
nor U17951 (N_17951,N_17653,N_17667);
nand U17952 (N_17952,N_17692,N_17653);
nor U17953 (N_17953,N_17504,N_17623);
nor U17954 (N_17954,N_17501,N_17586);
and U17955 (N_17955,N_17630,N_17627);
nor U17956 (N_17956,N_17593,N_17653);
or U17957 (N_17957,N_17596,N_17745);
nand U17958 (N_17958,N_17699,N_17603);
or U17959 (N_17959,N_17616,N_17596);
nand U17960 (N_17960,N_17714,N_17746);
nand U17961 (N_17961,N_17553,N_17532);
xor U17962 (N_17962,N_17639,N_17637);
or U17963 (N_17963,N_17531,N_17539);
or U17964 (N_17964,N_17558,N_17690);
and U17965 (N_17965,N_17528,N_17717);
nor U17966 (N_17966,N_17593,N_17576);
and U17967 (N_17967,N_17546,N_17524);
xnor U17968 (N_17968,N_17677,N_17636);
nand U17969 (N_17969,N_17538,N_17680);
or U17970 (N_17970,N_17656,N_17525);
and U17971 (N_17971,N_17737,N_17730);
nor U17972 (N_17972,N_17600,N_17552);
nor U17973 (N_17973,N_17621,N_17695);
or U17974 (N_17974,N_17520,N_17597);
xnor U17975 (N_17975,N_17521,N_17665);
and U17976 (N_17976,N_17626,N_17537);
or U17977 (N_17977,N_17525,N_17532);
and U17978 (N_17978,N_17747,N_17708);
nor U17979 (N_17979,N_17736,N_17622);
nand U17980 (N_17980,N_17672,N_17556);
or U17981 (N_17981,N_17531,N_17668);
xor U17982 (N_17982,N_17515,N_17528);
and U17983 (N_17983,N_17690,N_17707);
nor U17984 (N_17984,N_17687,N_17646);
nand U17985 (N_17985,N_17726,N_17592);
nand U17986 (N_17986,N_17673,N_17607);
nor U17987 (N_17987,N_17589,N_17668);
nor U17988 (N_17988,N_17636,N_17675);
or U17989 (N_17989,N_17724,N_17582);
or U17990 (N_17990,N_17501,N_17672);
xor U17991 (N_17991,N_17508,N_17581);
xnor U17992 (N_17992,N_17719,N_17707);
xnor U17993 (N_17993,N_17709,N_17686);
and U17994 (N_17994,N_17519,N_17502);
nand U17995 (N_17995,N_17541,N_17734);
nand U17996 (N_17996,N_17736,N_17545);
or U17997 (N_17997,N_17709,N_17625);
nand U17998 (N_17998,N_17581,N_17698);
nor U17999 (N_17999,N_17609,N_17610);
or U18000 (N_18000,N_17985,N_17841);
xor U18001 (N_18001,N_17842,N_17852);
nor U18002 (N_18002,N_17814,N_17895);
nor U18003 (N_18003,N_17830,N_17755);
and U18004 (N_18004,N_17752,N_17946);
nor U18005 (N_18005,N_17956,N_17983);
xor U18006 (N_18006,N_17828,N_17858);
xnor U18007 (N_18007,N_17861,N_17989);
and U18008 (N_18008,N_17905,N_17951);
nand U18009 (N_18009,N_17885,N_17898);
xnor U18010 (N_18010,N_17929,N_17821);
or U18011 (N_18011,N_17772,N_17869);
xor U18012 (N_18012,N_17923,N_17974);
xnor U18013 (N_18013,N_17884,N_17896);
nand U18014 (N_18014,N_17826,N_17777);
nor U18015 (N_18015,N_17959,N_17824);
nand U18016 (N_18016,N_17787,N_17784);
or U18017 (N_18017,N_17786,N_17998);
or U18018 (N_18018,N_17897,N_17937);
and U18019 (N_18019,N_17924,N_17789);
and U18020 (N_18020,N_17878,N_17843);
nand U18021 (N_18021,N_17811,N_17846);
xnor U18022 (N_18022,N_17805,N_17753);
xnor U18023 (N_18023,N_17860,N_17851);
nor U18024 (N_18024,N_17840,N_17958);
nand U18025 (N_18025,N_17818,N_17980);
and U18026 (N_18026,N_17867,N_17750);
nand U18027 (N_18027,N_17900,N_17973);
or U18028 (N_18028,N_17854,N_17944);
nand U18029 (N_18029,N_17812,N_17835);
or U18030 (N_18030,N_17763,N_17850);
or U18031 (N_18031,N_17922,N_17836);
nand U18032 (N_18032,N_17968,N_17965);
nor U18033 (N_18033,N_17979,N_17950);
nor U18034 (N_18034,N_17890,N_17925);
nand U18035 (N_18035,N_17798,N_17916);
xor U18036 (N_18036,N_17810,N_17780);
xor U18037 (N_18037,N_17970,N_17893);
nor U18038 (N_18038,N_17794,N_17954);
xnor U18039 (N_18039,N_17957,N_17876);
or U18040 (N_18040,N_17995,N_17764);
and U18041 (N_18041,N_17797,N_17768);
nor U18042 (N_18042,N_17941,N_17803);
nand U18043 (N_18043,N_17807,N_17855);
xnor U18044 (N_18044,N_17899,N_17817);
nand U18045 (N_18045,N_17976,N_17820);
and U18046 (N_18046,N_17991,N_17868);
or U18047 (N_18047,N_17760,N_17781);
nor U18048 (N_18048,N_17879,N_17804);
nand U18049 (N_18049,N_17791,N_17907);
xnor U18050 (N_18050,N_17931,N_17782);
and U18051 (N_18051,N_17971,N_17774);
nand U18052 (N_18052,N_17845,N_17783);
and U18053 (N_18053,N_17779,N_17847);
and U18054 (N_18054,N_17833,N_17999);
or U18055 (N_18055,N_17966,N_17908);
or U18056 (N_18056,N_17862,N_17911);
nand U18057 (N_18057,N_17939,N_17880);
nand U18058 (N_18058,N_17904,N_17825);
nand U18059 (N_18059,N_17751,N_17758);
and U18060 (N_18060,N_17819,N_17775);
xor U18061 (N_18061,N_17888,N_17886);
or U18062 (N_18062,N_17994,N_17961);
or U18063 (N_18063,N_17874,N_17953);
nor U18064 (N_18064,N_17917,N_17802);
nor U18065 (N_18065,N_17938,N_17914);
nor U18066 (N_18066,N_17838,N_17770);
nor U18067 (N_18067,N_17792,N_17933);
xor U18068 (N_18068,N_17873,N_17837);
nand U18069 (N_18069,N_17864,N_17912);
xor U18070 (N_18070,N_17815,N_17800);
or U18071 (N_18071,N_17806,N_17993);
nand U18072 (N_18072,N_17975,N_17793);
or U18073 (N_18073,N_17865,N_17857);
or U18074 (N_18074,N_17813,N_17808);
xnor U18075 (N_18075,N_17769,N_17871);
xor U18076 (N_18076,N_17892,N_17952);
and U18077 (N_18077,N_17955,N_17928);
and U18078 (N_18078,N_17992,N_17771);
nor U18079 (N_18079,N_17809,N_17778);
nand U18080 (N_18080,N_17920,N_17997);
nand U18081 (N_18081,N_17894,N_17915);
nand U18082 (N_18082,N_17788,N_17767);
nor U18083 (N_18083,N_17913,N_17766);
xnor U18084 (N_18084,N_17906,N_17949);
nand U18085 (N_18085,N_17964,N_17801);
or U18086 (N_18086,N_17849,N_17754);
and U18087 (N_18087,N_17934,N_17839);
and U18088 (N_18088,N_17972,N_17773);
and U18089 (N_18089,N_17823,N_17921);
nand U18090 (N_18090,N_17856,N_17872);
nor U18091 (N_18091,N_17960,N_17910);
xor U18092 (N_18092,N_17883,N_17963);
nand U18093 (N_18093,N_17881,N_17863);
nand U18094 (N_18094,N_17932,N_17936);
nand U18095 (N_18095,N_17940,N_17848);
nand U18096 (N_18096,N_17948,N_17967);
and U18097 (N_18097,N_17984,N_17942);
xnor U18098 (N_18098,N_17796,N_17947);
nor U18099 (N_18099,N_17829,N_17762);
nor U18100 (N_18100,N_17962,N_17853);
nor U18101 (N_18101,N_17945,N_17903);
nor U18102 (N_18102,N_17919,N_17827);
xor U18103 (N_18103,N_17943,N_17875);
nand U18104 (N_18104,N_17887,N_17982);
xor U18105 (N_18105,N_17859,N_17832);
and U18106 (N_18106,N_17822,N_17834);
and U18107 (N_18107,N_17756,N_17870);
xor U18108 (N_18108,N_17877,N_17969);
nor U18109 (N_18109,N_17831,N_17990);
xor U18110 (N_18110,N_17986,N_17761);
nand U18111 (N_18111,N_17926,N_17977);
or U18112 (N_18112,N_17757,N_17987);
nand U18113 (N_18113,N_17981,N_17988);
and U18114 (N_18114,N_17978,N_17909);
and U18115 (N_18115,N_17927,N_17930);
xor U18116 (N_18116,N_17918,N_17765);
and U18117 (N_18117,N_17776,N_17901);
xnor U18118 (N_18118,N_17891,N_17795);
xnor U18119 (N_18119,N_17882,N_17816);
xnor U18120 (N_18120,N_17889,N_17785);
and U18121 (N_18121,N_17866,N_17759);
or U18122 (N_18122,N_17799,N_17844);
xnor U18123 (N_18123,N_17902,N_17996);
or U18124 (N_18124,N_17790,N_17935);
nor U18125 (N_18125,N_17814,N_17984);
nand U18126 (N_18126,N_17811,N_17752);
or U18127 (N_18127,N_17944,N_17758);
nand U18128 (N_18128,N_17971,N_17893);
nor U18129 (N_18129,N_17885,N_17975);
or U18130 (N_18130,N_17846,N_17822);
and U18131 (N_18131,N_17928,N_17988);
and U18132 (N_18132,N_17751,N_17833);
or U18133 (N_18133,N_17981,N_17813);
and U18134 (N_18134,N_17942,N_17977);
or U18135 (N_18135,N_17828,N_17938);
or U18136 (N_18136,N_17938,N_17780);
nor U18137 (N_18137,N_17912,N_17806);
nor U18138 (N_18138,N_17892,N_17991);
and U18139 (N_18139,N_17815,N_17774);
or U18140 (N_18140,N_17996,N_17949);
nand U18141 (N_18141,N_17962,N_17830);
or U18142 (N_18142,N_17941,N_17894);
xnor U18143 (N_18143,N_17974,N_17947);
xor U18144 (N_18144,N_17935,N_17783);
nand U18145 (N_18145,N_17786,N_17953);
or U18146 (N_18146,N_17987,N_17919);
xor U18147 (N_18147,N_17974,N_17833);
xnor U18148 (N_18148,N_17892,N_17776);
or U18149 (N_18149,N_17754,N_17751);
nand U18150 (N_18150,N_17881,N_17888);
nand U18151 (N_18151,N_17821,N_17858);
and U18152 (N_18152,N_17906,N_17857);
or U18153 (N_18153,N_17995,N_17942);
xnor U18154 (N_18154,N_17873,N_17994);
and U18155 (N_18155,N_17940,N_17998);
or U18156 (N_18156,N_17805,N_17948);
and U18157 (N_18157,N_17816,N_17999);
and U18158 (N_18158,N_17914,N_17843);
nor U18159 (N_18159,N_17789,N_17975);
and U18160 (N_18160,N_17964,N_17870);
nand U18161 (N_18161,N_17952,N_17942);
or U18162 (N_18162,N_17758,N_17915);
nand U18163 (N_18163,N_17878,N_17763);
nand U18164 (N_18164,N_17985,N_17792);
nor U18165 (N_18165,N_17916,N_17847);
and U18166 (N_18166,N_17988,N_17862);
nand U18167 (N_18167,N_17931,N_17839);
or U18168 (N_18168,N_17837,N_17926);
and U18169 (N_18169,N_17997,N_17996);
and U18170 (N_18170,N_17943,N_17825);
xor U18171 (N_18171,N_17782,N_17769);
nor U18172 (N_18172,N_17995,N_17868);
nor U18173 (N_18173,N_17991,N_17862);
nand U18174 (N_18174,N_17944,N_17765);
or U18175 (N_18175,N_17985,N_17750);
nor U18176 (N_18176,N_17998,N_17871);
or U18177 (N_18177,N_17796,N_17884);
nand U18178 (N_18178,N_17884,N_17844);
or U18179 (N_18179,N_17783,N_17797);
and U18180 (N_18180,N_17807,N_17885);
or U18181 (N_18181,N_17940,N_17973);
or U18182 (N_18182,N_17899,N_17804);
nor U18183 (N_18183,N_17924,N_17891);
nor U18184 (N_18184,N_17765,N_17789);
and U18185 (N_18185,N_17976,N_17863);
or U18186 (N_18186,N_17968,N_17909);
or U18187 (N_18187,N_17979,N_17988);
nor U18188 (N_18188,N_17909,N_17991);
nand U18189 (N_18189,N_17826,N_17972);
nor U18190 (N_18190,N_17773,N_17764);
and U18191 (N_18191,N_17785,N_17772);
nor U18192 (N_18192,N_17861,N_17881);
nor U18193 (N_18193,N_17831,N_17823);
nor U18194 (N_18194,N_17955,N_17790);
nor U18195 (N_18195,N_17834,N_17875);
nor U18196 (N_18196,N_17764,N_17777);
and U18197 (N_18197,N_17948,N_17778);
and U18198 (N_18198,N_17927,N_17837);
and U18199 (N_18199,N_17990,N_17801);
nand U18200 (N_18200,N_17858,N_17960);
or U18201 (N_18201,N_17821,N_17907);
and U18202 (N_18202,N_17953,N_17779);
xnor U18203 (N_18203,N_17965,N_17930);
and U18204 (N_18204,N_17898,N_17818);
nand U18205 (N_18205,N_17891,N_17959);
and U18206 (N_18206,N_17886,N_17878);
nand U18207 (N_18207,N_17788,N_17880);
nand U18208 (N_18208,N_17802,N_17801);
xor U18209 (N_18209,N_17975,N_17996);
xnor U18210 (N_18210,N_17829,N_17823);
or U18211 (N_18211,N_17926,N_17913);
and U18212 (N_18212,N_17910,N_17928);
xor U18213 (N_18213,N_17775,N_17944);
and U18214 (N_18214,N_17950,N_17813);
and U18215 (N_18215,N_17885,N_17895);
nand U18216 (N_18216,N_17845,N_17915);
nor U18217 (N_18217,N_17755,N_17765);
nand U18218 (N_18218,N_17900,N_17979);
nand U18219 (N_18219,N_17980,N_17952);
xor U18220 (N_18220,N_17785,N_17812);
and U18221 (N_18221,N_17876,N_17882);
nor U18222 (N_18222,N_17946,N_17763);
nor U18223 (N_18223,N_17975,N_17992);
and U18224 (N_18224,N_17832,N_17778);
and U18225 (N_18225,N_17930,N_17866);
and U18226 (N_18226,N_17962,N_17891);
xnor U18227 (N_18227,N_17942,N_17993);
nor U18228 (N_18228,N_17817,N_17971);
nor U18229 (N_18229,N_17843,N_17890);
or U18230 (N_18230,N_17925,N_17769);
and U18231 (N_18231,N_17962,N_17778);
and U18232 (N_18232,N_17820,N_17936);
and U18233 (N_18233,N_17872,N_17767);
or U18234 (N_18234,N_17788,N_17918);
and U18235 (N_18235,N_17917,N_17954);
xnor U18236 (N_18236,N_17822,N_17990);
nand U18237 (N_18237,N_17967,N_17848);
nand U18238 (N_18238,N_17870,N_17758);
nor U18239 (N_18239,N_17837,N_17841);
or U18240 (N_18240,N_17863,N_17902);
and U18241 (N_18241,N_17977,N_17886);
or U18242 (N_18242,N_17858,N_17971);
xnor U18243 (N_18243,N_17784,N_17973);
or U18244 (N_18244,N_17877,N_17997);
and U18245 (N_18245,N_17813,N_17988);
and U18246 (N_18246,N_17865,N_17905);
and U18247 (N_18247,N_17786,N_17896);
or U18248 (N_18248,N_17770,N_17999);
xnor U18249 (N_18249,N_17965,N_17795);
and U18250 (N_18250,N_18064,N_18244);
and U18251 (N_18251,N_18056,N_18213);
xor U18252 (N_18252,N_18216,N_18077);
xor U18253 (N_18253,N_18199,N_18089);
and U18254 (N_18254,N_18150,N_18104);
nand U18255 (N_18255,N_18074,N_18133);
xnor U18256 (N_18256,N_18190,N_18013);
nor U18257 (N_18257,N_18103,N_18241);
and U18258 (N_18258,N_18026,N_18172);
nor U18259 (N_18259,N_18095,N_18215);
nor U18260 (N_18260,N_18145,N_18003);
or U18261 (N_18261,N_18247,N_18075);
and U18262 (N_18262,N_18081,N_18094);
xor U18263 (N_18263,N_18017,N_18163);
and U18264 (N_18264,N_18186,N_18248);
xnor U18265 (N_18265,N_18041,N_18178);
and U18266 (N_18266,N_18243,N_18065);
xnor U18267 (N_18267,N_18173,N_18112);
xnor U18268 (N_18268,N_18008,N_18098);
or U18269 (N_18269,N_18036,N_18191);
nand U18270 (N_18270,N_18181,N_18130);
or U18271 (N_18271,N_18200,N_18083);
or U18272 (N_18272,N_18237,N_18023);
nand U18273 (N_18273,N_18070,N_18205);
or U18274 (N_18274,N_18234,N_18156);
nor U18275 (N_18275,N_18125,N_18019);
and U18276 (N_18276,N_18055,N_18211);
nor U18277 (N_18277,N_18227,N_18196);
nand U18278 (N_18278,N_18062,N_18082);
xor U18279 (N_18279,N_18087,N_18158);
nor U18280 (N_18280,N_18031,N_18143);
xnor U18281 (N_18281,N_18141,N_18010);
nand U18282 (N_18282,N_18048,N_18167);
xnor U18283 (N_18283,N_18151,N_18030);
or U18284 (N_18284,N_18146,N_18137);
and U18285 (N_18285,N_18240,N_18076);
or U18286 (N_18286,N_18127,N_18028);
nor U18287 (N_18287,N_18230,N_18111);
nand U18288 (N_18288,N_18035,N_18084);
xnor U18289 (N_18289,N_18113,N_18174);
xor U18290 (N_18290,N_18136,N_18233);
nand U18291 (N_18291,N_18142,N_18086);
nor U18292 (N_18292,N_18228,N_18051);
xor U18293 (N_18293,N_18022,N_18197);
or U18294 (N_18294,N_18085,N_18015);
nor U18295 (N_18295,N_18219,N_18222);
or U18296 (N_18296,N_18018,N_18162);
nor U18297 (N_18297,N_18000,N_18209);
nor U18298 (N_18298,N_18132,N_18079);
or U18299 (N_18299,N_18155,N_18067);
nor U18300 (N_18300,N_18032,N_18118);
xnor U18301 (N_18301,N_18135,N_18129);
nor U18302 (N_18302,N_18044,N_18179);
nor U18303 (N_18303,N_18193,N_18096);
or U18304 (N_18304,N_18110,N_18061);
xnor U18305 (N_18305,N_18057,N_18042);
nand U18306 (N_18306,N_18206,N_18047);
nor U18307 (N_18307,N_18012,N_18126);
or U18308 (N_18308,N_18101,N_18192);
nand U18309 (N_18309,N_18007,N_18235);
xnor U18310 (N_18310,N_18177,N_18097);
or U18311 (N_18311,N_18105,N_18168);
xor U18312 (N_18312,N_18050,N_18242);
or U18313 (N_18313,N_18232,N_18164);
or U18314 (N_18314,N_18184,N_18180);
xor U18315 (N_18315,N_18045,N_18069);
and U18316 (N_18316,N_18034,N_18198);
nand U18317 (N_18317,N_18063,N_18231);
nand U18318 (N_18318,N_18147,N_18033);
nor U18319 (N_18319,N_18040,N_18091);
and U18320 (N_18320,N_18005,N_18049);
xnor U18321 (N_18321,N_18202,N_18002);
xnor U18322 (N_18322,N_18175,N_18149);
nor U18323 (N_18323,N_18122,N_18139);
xor U18324 (N_18324,N_18249,N_18090);
nor U18325 (N_18325,N_18229,N_18188);
and U18326 (N_18326,N_18225,N_18221);
and U18327 (N_18327,N_18024,N_18208);
and U18328 (N_18328,N_18121,N_18166);
or U18329 (N_18329,N_18194,N_18115);
nand U18330 (N_18330,N_18109,N_18088);
xnor U18331 (N_18331,N_18068,N_18239);
xnor U18332 (N_18332,N_18020,N_18182);
nor U18333 (N_18333,N_18176,N_18066);
and U18334 (N_18334,N_18140,N_18171);
nor U18335 (N_18335,N_18078,N_18187);
or U18336 (N_18336,N_18059,N_18117);
and U18337 (N_18337,N_18072,N_18152);
or U18338 (N_18338,N_18224,N_18120);
nor U18339 (N_18339,N_18052,N_18071);
and U18340 (N_18340,N_18092,N_18246);
or U18341 (N_18341,N_18016,N_18226);
or U18342 (N_18342,N_18009,N_18037);
nand U18343 (N_18343,N_18159,N_18148);
nor U18344 (N_18344,N_18006,N_18093);
nand U18345 (N_18345,N_18058,N_18183);
or U18346 (N_18346,N_18038,N_18138);
or U18347 (N_18347,N_18106,N_18039);
and U18348 (N_18348,N_18201,N_18154);
and U18349 (N_18349,N_18046,N_18217);
or U18350 (N_18350,N_18124,N_18220);
and U18351 (N_18351,N_18203,N_18027);
nor U18352 (N_18352,N_18236,N_18100);
nor U18353 (N_18353,N_18128,N_18238);
and U18354 (N_18354,N_18218,N_18014);
or U18355 (N_18355,N_18204,N_18189);
or U18356 (N_18356,N_18157,N_18107);
nand U18357 (N_18357,N_18123,N_18153);
nor U18358 (N_18358,N_18195,N_18004);
and U18359 (N_18359,N_18116,N_18185);
or U18360 (N_18360,N_18073,N_18210);
nor U18361 (N_18361,N_18245,N_18161);
nor U18362 (N_18362,N_18054,N_18134);
nand U18363 (N_18363,N_18207,N_18099);
nand U18364 (N_18364,N_18025,N_18114);
or U18365 (N_18365,N_18102,N_18001);
nor U18366 (N_18366,N_18214,N_18170);
xor U18367 (N_18367,N_18108,N_18119);
and U18368 (N_18368,N_18060,N_18080);
and U18369 (N_18369,N_18011,N_18021);
nor U18370 (N_18370,N_18169,N_18212);
and U18371 (N_18371,N_18043,N_18144);
nand U18372 (N_18372,N_18053,N_18165);
or U18373 (N_18373,N_18223,N_18029);
xor U18374 (N_18374,N_18160,N_18131);
nand U18375 (N_18375,N_18007,N_18123);
xnor U18376 (N_18376,N_18219,N_18016);
nand U18377 (N_18377,N_18198,N_18197);
nand U18378 (N_18378,N_18034,N_18166);
or U18379 (N_18379,N_18007,N_18144);
nand U18380 (N_18380,N_18181,N_18167);
and U18381 (N_18381,N_18056,N_18219);
and U18382 (N_18382,N_18125,N_18029);
xnor U18383 (N_18383,N_18169,N_18050);
xor U18384 (N_18384,N_18142,N_18161);
nor U18385 (N_18385,N_18241,N_18004);
or U18386 (N_18386,N_18220,N_18149);
xnor U18387 (N_18387,N_18197,N_18244);
nand U18388 (N_18388,N_18070,N_18056);
or U18389 (N_18389,N_18175,N_18134);
nand U18390 (N_18390,N_18196,N_18190);
or U18391 (N_18391,N_18209,N_18171);
xor U18392 (N_18392,N_18002,N_18115);
or U18393 (N_18393,N_18037,N_18078);
nor U18394 (N_18394,N_18050,N_18157);
or U18395 (N_18395,N_18153,N_18049);
or U18396 (N_18396,N_18067,N_18061);
or U18397 (N_18397,N_18195,N_18012);
nand U18398 (N_18398,N_18085,N_18101);
or U18399 (N_18399,N_18201,N_18129);
or U18400 (N_18400,N_18041,N_18174);
and U18401 (N_18401,N_18032,N_18181);
or U18402 (N_18402,N_18181,N_18017);
or U18403 (N_18403,N_18087,N_18131);
nor U18404 (N_18404,N_18177,N_18122);
nor U18405 (N_18405,N_18069,N_18070);
or U18406 (N_18406,N_18035,N_18224);
nand U18407 (N_18407,N_18174,N_18020);
and U18408 (N_18408,N_18157,N_18230);
and U18409 (N_18409,N_18178,N_18015);
xor U18410 (N_18410,N_18158,N_18118);
and U18411 (N_18411,N_18239,N_18030);
xor U18412 (N_18412,N_18161,N_18188);
or U18413 (N_18413,N_18175,N_18133);
nand U18414 (N_18414,N_18144,N_18239);
xor U18415 (N_18415,N_18207,N_18138);
nor U18416 (N_18416,N_18044,N_18203);
or U18417 (N_18417,N_18119,N_18230);
nand U18418 (N_18418,N_18075,N_18158);
nor U18419 (N_18419,N_18104,N_18115);
xor U18420 (N_18420,N_18164,N_18237);
nor U18421 (N_18421,N_18085,N_18021);
or U18422 (N_18422,N_18124,N_18209);
or U18423 (N_18423,N_18166,N_18011);
or U18424 (N_18424,N_18090,N_18021);
nor U18425 (N_18425,N_18021,N_18236);
and U18426 (N_18426,N_18202,N_18159);
and U18427 (N_18427,N_18233,N_18074);
xor U18428 (N_18428,N_18198,N_18230);
or U18429 (N_18429,N_18149,N_18052);
nor U18430 (N_18430,N_18005,N_18108);
or U18431 (N_18431,N_18031,N_18014);
nor U18432 (N_18432,N_18112,N_18192);
nor U18433 (N_18433,N_18079,N_18043);
and U18434 (N_18434,N_18234,N_18208);
xnor U18435 (N_18435,N_18133,N_18237);
and U18436 (N_18436,N_18247,N_18000);
or U18437 (N_18437,N_18193,N_18145);
xor U18438 (N_18438,N_18107,N_18169);
and U18439 (N_18439,N_18077,N_18042);
and U18440 (N_18440,N_18243,N_18103);
and U18441 (N_18441,N_18006,N_18106);
xor U18442 (N_18442,N_18007,N_18164);
nand U18443 (N_18443,N_18144,N_18190);
nand U18444 (N_18444,N_18193,N_18086);
or U18445 (N_18445,N_18127,N_18195);
and U18446 (N_18446,N_18077,N_18054);
or U18447 (N_18447,N_18089,N_18017);
or U18448 (N_18448,N_18102,N_18140);
nor U18449 (N_18449,N_18008,N_18223);
and U18450 (N_18450,N_18053,N_18076);
or U18451 (N_18451,N_18030,N_18240);
nand U18452 (N_18452,N_18006,N_18127);
nand U18453 (N_18453,N_18054,N_18181);
nand U18454 (N_18454,N_18183,N_18127);
nor U18455 (N_18455,N_18131,N_18127);
xnor U18456 (N_18456,N_18222,N_18025);
nand U18457 (N_18457,N_18097,N_18213);
nor U18458 (N_18458,N_18183,N_18028);
nand U18459 (N_18459,N_18005,N_18219);
or U18460 (N_18460,N_18038,N_18059);
xor U18461 (N_18461,N_18190,N_18073);
nor U18462 (N_18462,N_18029,N_18136);
or U18463 (N_18463,N_18142,N_18087);
nor U18464 (N_18464,N_18090,N_18152);
or U18465 (N_18465,N_18171,N_18108);
nor U18466 (N_18466,N_18082,N_18234);
or U18467 (N_18467,N_18086,N_18216);
and U18468 (N_18468,N_18050,N_18118);
and U18469 (N_18469,N_18058,N_18159);
xor U18470 (N_18470,N_18059,N_18161);
or U18471 (N_18471,N_18164,N_18008);
and U18472 (N_18472,N_18056,N_18228);
and U18473 (N_18473,N_18235,N_18222);
nor U18474 (N_18474,N_18069,N_18111);
nand U18475 (N_18475,N_18215,N_18023);
nor U18476 (N_18476,N_18098,N_18168);
nand U18477 (N_18477,N_18177,N_18013);
xor U18478 (N_18478,N_18141,N_18184);
nand U18479 (N_18479,N_18131,N_18027);
xnor U18480 (N_18480,N_18233,N_18028);
nor U18481 (N_18481,N_18048,N_18125);
nand U18482 (N_18482,N_18190,N_18029);
or U18483 (N_18483,N_18037,N_18120);
nand U18484 (N_18484,N_18032,N_18085);
or U18485 (N_18485,N_18096,N_18029);
and U18486 (N_18486,N_18160,N_18209);
xnor U18487 (N_18487,N_18156,N_18218);
and U18488 (N_18488,N_18114,N_18073);
and U18489 (N_18489,N_18242,N_18176);
xor U18490 (N_18490,N_18155,N_18218);
or U18491 (N_18491,N_18071,N_18144);
nor U18492 (N_18492,N_18206,N_18111);
nor U18493 (N_18493,N_18228,N_18019);
or U18494 (N_18494,N_18241,N_18248);
nand U18495 (N_18495,N_18211,N_18127);
and U18496 (N_18496,N_18001,N_18044);
nand U18497 (N_18497,N_18076,N_18184);
xor U18498 (N_18498,N_18020,N_18071);
and U18499 (N_18499,N_18015,N_18093);
nand U18500 (N_18500,N_18446,N_18356);
nand U18501 (N_18501,N_18477,N_18443);
nand U18502 (N_18502,N_18496,N_18343);
nor U18503 (N_18503,N_18307,N_18381);
and U18504 (N_18504,N_18283,N_18452);
and U18505 (N_18505,N_18396,N_18324);
or U18506 (N_18506,N_18404,N_18401);
or U18507 (N_18507,N_18376,N_18363);
and U18508 (N_18508,N_18412,N_18304);
nand U18509 (N_18509,N_18284,N_18441);
nor U18510 (N_18510,N_18310,N_18313);
nor U18511 (N_18511,N_18489,N_18348);
xor U18512 (N_18512,N_18293,N_18382);
and U18513 (N_18513,N_18261,N_18469);
and U18514 (N_18514,N_18466,N_18357);
xnor U18515 (N_18515,N_18292,N_18306);
or U18516 (N_18516,N_18353,N_18424);
and U18517 (N_18517,N_18332,N_18388);
or U18518 (N_18518,N_18468,N_18456);
xor U18519 (N_18519,N_18354,N_18337);
and U18520 (N_18520,N_18492,N_18392);
or U18521 (N_18521,N_18482,N_18393);
nand U18522 (N_18522,N_18276,N_18488);
xor U18523 (N_18523,N_18269,N_18472);
nor U18524 (N_18524,N_18336,N_18254);
nand U18525 (N_18525,N_18440,N_18263);
xor U18526 (N_18526,N_18397,N_18335);
nand U18527 (N_18527,N_18330,N_18478);
or U18528 (N_18528,N_18314,N_18437);
nand U18529 (N_18529,N_18408,N_18334);
and U18530 (N_18530,N_18394,N_18426);
or U18531 (N_18531,N_18409,N_18458);
or U18532 (N_18532,N_18379,N_18368);
nor U18533 (N_18533,N_18296,N_18258);
nor U18534 (N_18534,N_18251,N_18250);
nor U18535 (N_18535,N_18407,N_18290);
or U18536 (N_18536,N_18374,N_18346);
and U18537 (N_18537,N_18311,N_18367);
nor U18538 (N_18538,N_18411,N_18427);
and U18539 (N_18539,N_18257,N_18453);
nand U18540 (N_18540,N_18420,N_18295);
nand U18541 (N_18541,N_18390,N_18398);
xnor U18542 (N_18542,N_18480,N_18460);
and U18543 (N_18543,N_18272,N_18385);
nand U18544 (N_18544,N_18422,N_18485);
nand U18545 (N_18545,N_18358,N_18445);
nand U18546 (N_18546,N_18282,N_18338);
nand U18547 (N_18547,N_18349,N_18359);
nand U18548 (N_18548,N_18298,N_18326);
and U18549 (N_18549,N_18444,N_18487);
xor U18550 (N_18550,N_18253,N_18289);
nand U18551 (N_18551,N_18291,N_18499);
and U18552 (N_18552,N_18389,N_18369);
nor U18553 (N_18553,N_18459,N_18302);
xnor U18554 (N_18554,N_18266,N_18341);
or U18555 (N_18555,N_18299,N_18451);
and U18556 (N_18556,N_18395,N_18345);
nor U18557 (N_18557,N_18457,N_18418);
xor U18558 (N_18558,N_18461,N_18486);
nand U18559 (N_18559,N_18277,N_18316);
and U18560 (N_18560,N_18462,N_18474);
nand U18561 (N_18561,N_18325,N_18386);
nor U18562 (N_18562,N_18429,N_18475);
and U18563 (N_18563,N_18301,N_18383);
or U18564 (N_18564,N_18320,N_18484);
xnor U18565 (N_18565,N_18373,N_18454);
or U18566 (N_18566,N_18450,N_18464);
nor U18567 (N_18567,N_18323,N_18252);
nand U18568 (N_18568,N_18271,N_18428);
nand U18569 (N_18569,N_18305,N_18435);
nand U18570 (N_18570,N_18423,N_18260);
nand U18571 (N_18571,N_18463,N_18279);
and U18572 (N_18572,N_18372,N_18285);
xnor U18573 (N_18573,N_18439,N_18491);
nand U18574 (N_18574,N_18476,N_18391);
xnor U18575 (N_18575,N_18360,N_18483);
nor U18576 (N_18576,N_18433,N_18490);
or U18577 (N_18577,N_18312,N_18402);
nor U18578 (N_18578,N_18327,N_18414);
and U18579 (N_18579,N_18415,N_18399);
nand U18580 (N_18580,N_18256,N_18430);
xor U18581 (N_18581,N_18378,N_18339);
xor U18582 (N_18582,N_18344,N_18438);
and U18583 (N_18583,N_18436,N_18361);
xnor U18584 (N_18584,N_18286,N_18403);
and U18585 (N_18585,N_18405,N_18494);
or U18586 (N_18586,N_18421,N_18364);
nand U18587 (N_18587,N_18321,N_18273);
xnor U18588 (N_18588,N_18309,N_18497);
and U18589 (N_18589,N_18384,N_18300);
xnor U18590 (N_18590,N_18465,N_18417);
nand U18591 (N_18591,N_18351,N_18375);
and U18592 (N_18592,N_18287,N_18431);
nand U18593 (N_18593,N_18493,N_18255);
nor U18594 (N_18594,N_18280,N_18328);
or U18595 (N_18595,N_18303,N_18413);
nand U18596 (N_18596,N_18371,N_18432);
and U18597 (N_18597,N_18265,N_18455);
nor U18598 (N_18598,N_18410,N_18317);
nor U18599 (N_18599,N_18340,N_18425);
nand U18600 (N_18600,N_18406,N_18275);
nand U18601 (N_18601,N_18288,N_18470);
and U18602 (N_18602,N_18362,N_18387);
or U18603 (N_18603,N_18448,N_18350);
nor U18604 (N_18604,N_18416,N_18400);
nor U18605 (N_18605,N_18467,N_18473);
nand U18606 (N_18606,N_18481,N_18281);
or U18607 (N_18607,N_18347,N_18268);
nor U18608 (N_18608,N_18449,N_18447);
and U18609 (N_18609,N_18366,N_18419);
nor U18610 (N_18610,N_18315,N_18297);
nand U18611 (N_18611,N_18495,N_18294);
nand U18612 (N_18612,N_18329,N_18274);
and U18613 (N_18613,N_18442,N_18318);
and U18614 (N_18614,N_18377,N_18319);
nand U18615 (N_18615,N_18264,N_18308);
nand U18616 (N_18616,N_18365,N_18270);
nor U18617 (N_18617,N_18262,N_18342);
and U18618 (N_18618,N_18370,N_18471);
nand U18619 (N_18619,N_18479,N_18267);
and U18620 (N_18620,N_18434,N_18331);
xnor U18621 (N_18621,N_18380,N_18259);
nand U18622 (N_18622,N_18278,N_18355);
nand U18623 (N_18623,N_18322,N_18352);
nand U18624 (N_18624,N_18333,N_18498);
nor U18625 (N_18625,N_18255,N_18289);
nor U18626 (N_18626,N_18336,N_18317);
and U18627 (N_18627,N_18456,N_18362);
and U18628 (N_18628,N_18262,N_18451);
or U18629 (N_18629,N_18455,N_18446);
nor U18630 (N_18630,N_18277,N_18418);
or U18631 (N_18631,N_18386,N_18298);
xnor U18632 (N_18632,N_18376,N_18428);
or U18633 (N_18633,N_18379,N_18287);
nand U18634 (N_18634,N_18369,N_18446);
and U18635 (N_18635,N_18332,N_18331);
nor U18636 (N_18636,N_18281,N_18330);
nor U18637 (N_18637,N_18493,N_18258);
xnor U18638 (N_18638,N_18382,N_18365);
and U18639 (N_18639,N_18447,N_18340);
and U18640 (N_18640,N_18286,N_18464);
nand U18641 (N_18641,N_18321,N_18413);
nand U18642 (N_18642,N_18290,N_18367);
and U18643 (N_18643,N_18345,N_18482);
nand U18644 (N_18644,N_18365,N_18374);
and U18645 (N_18645,N_18365,N_18427);
or U18646 (N_18646,N_18250,N_18394);
nor U18647 (N_18647,N_18401,N_18332);
nand U18648 (N_18648,N_18338,N_18398);
and U18649 (N_18649,N_18499,N_18362);
and U18650 (N_18650,N_18452,N_18295);
or U18651 (N_18651,N_18304,N_18498);
and U18652 (N_18652,N_18367,N_18280);
nor U18653 (N_18653,N_18348,N_18313);
nor U18654 (N_18654,N_18284,N_18304);
nor U18655 (N_18655,N_18324,N_18453);
nor U18656 (N_18656,N_18287,N_18279);
xor U18657 (N_18657,N_18335,N_18353);
xor U18658 (N_18658,N_18471,N_18456);
nor U18659 (N_18659,N_18434,N_18429);
nand U18660 (N_18660,N_18374,N_18370);
and U18661 (N_18661,N_18347,N_18360);
xnor U18662 (N_18662,N_18346,N_18370);
or U18663 (N_18663,N_18319,N_18347);
nand U18664 (N_18664,N_18446,N_18324);
xor U18665 (N_18665,N_18333,N_18276);
xor U18666 (N_18666,N_18462,N_18402);
nor U18667 (N_18667,N_18490,N_18379);
nand U18668 (N_18668,N_18456,N_18321);
and U18669 (N_18669,N_18496,N_18494);
nand U18670 (N_18670,N_18295,N_18474);
nand U18671 (N_18671,N_18354,N_18353);
nand U18672 (N_18672,N_18301,N_18279);
or U18673 (N_18673,N_18338,N_18431);
nor U18674 (N_18674,N_18396,N_18420);
xnor U18675 (N_18675,N_18335,N_18492);
and U18676 (N_18676,N_18314,N_18292);
or U18677 (N_18677,N_18390,N_18426);
or U18678 (N_18678,N_18359,N_18254);
nor U18679 (N_18679,N_18323,N_18464);
nor U18680 (N_18680,N_18499,N_18432);
nor U18681 (N_18681,N_18372,N_18351);
nand U18682 (N_18682,N_18432,N_18463);
xor U18683 (N_18683,N_18322,N_18308);
and U18684 (N_18684,N_18284,N_18312);
xnor U18685 (N_18685,N_18478,N_18415);
xor U18686 (N_18686,N_18304,N_18263);
nor U18687 (N_18687,N_18397,N_18481);
and U18688 (N_18688,N_18449,N_18309);
nor U18689 (N_18689,N_18314,N_18458);
nor U18690 (N_18690,N_18396,N_18426);
xnor U18691 (N_18691,N_18492,N_18266);
nor U18692 (N_18692,N_18424,N_18458);
and U18693 (N_18693,N_18431,N_18430);
xnor U18694 (N_18694,N_18312,N_18316);
and U18695 (N_18695,N_18458,N_18342);
nand U18696 (N_18696,N_18324,N_18357);
nor U18697 (N_18697,N_18439,N_18496);
nor U18698 (N_18698,N_18390,N_18337);
xor U18699 (N_18699,N_18499,N_18385);
xor U18700 (N_18700,N_18353,N_18298);
or U18701 (N_18701,N_18473,N_18251);
or U18702 (N_18702,N_18333,N_18427);
or U18703 (N_18703,N_18329,N_18312);
xor U18704 (N_18704,N_18486,N_18250);
and U18705 (N_18705,N_18327,N_18317);
and U18706 (N_18706,N_18415,N_18304);
xnor U18707 (N_18707,N_18434,N_18492);
xor U18708 (N_18708,N_18348,N_18476);
or U18709 (N_18709,N_18329,N_18490);
and U18710 (N_18710,N_18472,N_18434);
xnor U18711 (N_18711,N_18427,N_18305);
or U18712 (N_18712,N_18473,N_18401);
nor U18713 (N_18713,N_18489,N_18453);
or U18714 (N_18714,N_18391,N_18483);
nor U18715 (N_18715,N_18436,N_18326);
xnor U18716 (N_18716,N_18250,N_18485);
and U18717 (N_18717,N_18474,N_18397);
xor U18718 (N_18718,N_18492,N_18289);
or U18719 (N_18719,N_18251,N_18417);
xnor U18720 (N_18720,N_18485,N_18453);
nor U18721 (N_18721,N_18312,N_18377);
nor U18722 (N_18722,N_18311,N_18447);
xnor U18723 (N_18723,N_18462,N_18338);
nand U18724 (N_18724,N_18313,N_18264);
xnor U18725 (N_18725,N_18351,N_18456);
nand U18726 (N_18726,N_18402,N_18494);
xor U18727 (N_18727,N_18385,N_18265);
or U18728 (N_18728,N_18360,N_18468);
and U18729 (N_18729,N_18349,N_18319);
and U18730 (N_18730,N_18391,N_18475);
xnor U18731 (N_18731,N_18496,N_18412);
xor U18732 (N_18732,N_18423,N_18321);
nor U18733 (N_18733,N_18273,N_18323);
xnor U18734 (N_18734,N_18299,N_18462);
xnor U18735 (N_18735,N_18258,N_18440);
nor U18736 (N_18736,N_18379,N_18299);
and U18737 (N_18737,N_18295,N_18442);
or U18738 (N_18738,N_18456,N_18447);
xnor U18739 (N_18739,N_18482,N_18447);
nor U18740 (N_18740,N_18415,N_18434);
nor U18741 (N_18741,N_18331,N_18450);
xnor U18742 (N_18742,N_18300,N_18416);
xnor U18743 (N_18743,N_18271,N_18375);
nor U18744 (N_18744,N_18347,N_18323);
and U18745 (N_18745,N_18305,N_18409);
or U18746 (N_18746,N_18435,N_18270);
and U18747 (N_18747,N_18434,N_18441);
or U18748 (N_18748,N_18298,N_18409);
and U18749 (N_18749,N_18399,N_18497);
nor U18750 (N_18750,N_18647,N_18505);
xnor U18751 (N_18751,N_18642,N_18539);
and U18752 (N_18752,N_18560,N_18596);
nor U18753 (N_18753,N_18748,N_18711);
nor U18754 (N_18754,N_18506,N_18638);
xnor U18755 (N_18755,N_18626,N_18535);
and U18756 (N_18756,N_18671,N_18507);
and U18757 (N_18757,N_18720,N_18685);
xnor U18758 (N_18758,N_18687,N_18602);
and U18759 (N_18759,N_18588,N_18503);
or U18760 (N_18760,N_18690,N_18741);
nand U18761 (N_18761,N_18686,N_18734);
nor U18762 (N_18762,N_18661,N_18715);
and U18763 (N_18763,N_18649,N_18727);
or U18764 (N_18764,N_18616,N_18608);
or U18765 (N_18765,N_18673,N_18597);
or U18766 (N_18766,N_18603,N_18553);
or U18767 (N_18767,N_18565,N_18587);
nand U18768 (N_18768,N_18634,N_18513);
nand U18769 (N_18769,N_18563,N_18611);
xor U18770 (N_18770,N_18624,N_18509);
nand U18771 (N_18771,N_18681,N_18742);
xnor U18772 (N_18772,N_18656,N_18645);
and U18773 (N_18773,N_18538,N_18708);
or U18774 (N_18774,N_18749,N_18567);
nor U18775 (N_18775,N_18704,N_18702);
nand U18776 (N_18776,N_18590,N_18728);
xnor U18777 (N_18777,N_18536,N_18533);
nor U18778 (N_18778,N_18559,N_18598);
xor U18779 (N_18779,N_18738,N_18639);
nor U18780 (N_18780,N_18546,N_18652);
nor U18781 (N_18781,N_18610,N_18580);
nor U18782 (N_18782,N_18568,N_18705);
or U18783 (N_18783,N_18730,N_18707);
and U18784 (N_18784,N_18532,N_18571);
xor U18785 (N_18785,N_18651,N_18672);
and U18786 (N_18786,N_18576,N_18696);
and U18787 (N_18787,N_18519,N_18591);
nand U18788 (N_18788,N_18745,N_18581);
xor U18789 (N_18789,N_18692,N_18574);
and U18790 (N_18790,N_18510,N_18542);
or U18791 (N_18791,N_18721,N_18606);
nor U18792 (N_18792,N_18713,N_18660);
and U18793 (N_18793,N_18575,N_18543);
nor U18794 (N_18794,N_18619,N_18743);
and U18795 (N_18795,N_18622,N_18670);
or U18796 (N_18796,N_18736,N_18694);
or U18797 (N_18797,N_18664,N_18650);
or U18798 (N_18798,N_18526,N_18569);
nor U18799 (N_18799,N_18657,N_18528);
xnor U18800 (N_18800,N_18551,N_18502);
nor U18801 (N_18801,N_18665,N_18592);
or U18802 (N_18802,N_18655,N_18555);
nor U18803 (N_18803,N_18607,N_18527);
xnor U18804 (N_18804,N_18654,N_18724);
xor U18805 (N_18805,N_18631,N_18501);
or U18806 (N_18806,N_18677,N_18531);
nor U18807 (N_18807,N_18675,N_18632);
and U18808 (N_18808,N_18522,N_18572);
or U18809 (N_18809,N_18698,N_18732);
nor U18810 (N_18810,N_18617,N_18541);
or U18811 (N_18811,N_18700,N_18570);
and U18812 (N_18812,N_18718,N_18737);
and U18813 (N_18813,N_18682,N_18593);
and U18814 (N_18814,N_18666,N_18620);
and U18815 (N_18815,N_18552,N_18693);
or U18816 (N_18816,N_18558,N_18662);
and U18817 (N_18817,N_18544,N_18697);
nand U18818 (N_18818,N_18641,N_18517);
or U18819 (N_18819,N_18684,N_18618);
nand U18820 (N_18820,N_18594,N_18625);
xnor U18821 (N_18821,N_18706,N_18735);
or U18822 (N_18822,N_18600,N_18549);
nor U18823 (N_18823,N_18548,N_18547);
xor U18824 (N_18824,N_18747,N_18710);
nor U18825 (N_18825,N_18586,N_18613);
nand U18826 (N_18826,N_18726,N_18578);
nand U18827 (N_18827,N_18577,N_18701);
nand U18828 (N_18828,N_18729,N_18722);
or U18829 (N_18829,N_18667,N_18640);
and U18830 (N_18830,N_18523,N_18669);
or U18831 (N_18831,N_18723,N_18534);
nor U18832 (N_18832,N_18689,N_18508);
nor U18833 (N_18833,N_18561,N_18582);
and U18834 (N_18834,N_18699,N_18668);
nand U18835 (N_18835,N_18595,N_18643);
nand U18836 (N_18836,N_18601,N_18676);
or U18837 (N_18837,N_18554,N_18630);
nand U18838 (N_18838,N_18589,N_18525);
xor U18839 (N_18839,N_18733,N_18614);
nor U18840 (N_18840,N_18500,N_18512);
xnor U18841 (N_18841,N_18562,N_18717);
or U18842 (N_18842,N_18688,N_18744);
nand U18843 (N_18843,N_18663,N_18678);
nor U18844 (N_18844,N_18605,N_18530);
nor U18845 (N_18845,N_18740,N_18629);
xnor U18846 (N_18846,N_18712,N_18719);
or U18847 (N_18847,N_18623,N_18564);
and U18848 (N_18848,N_18518,N_18604);
xor U18849 (N_18849,N_18573,N_18615);
and U18850 (N_18850,N_18709,N_18556);
nor U18851 (N_18851,N_18521,N_18583);
nand U18852 (N_18852,N_18648,N_18714);
xor U18853 (N_18853,N_18646,N_18537);
nor U18854 (N_18854,N_18679,N_18550);
nand U18855 (N_18855,N_18627,N_18691);
nor U18856 (N_18856,N_18545,N_18520);
nor U18857 (N_18857,N_18584,N_18674);
nand U18858 (N_18858,N_18524,N_18612);
xnor U18859 (N_18859,N_18540,N_18621);
or U18860 (N_18860,N_18633,N_18566);
xor U18861 (N_18861,N_18680,N_18659);
nand U18862 (N_18862,N_18739,N_18636);
nor U18863 (N_18863,N_18628,N_18683);
xnor U18864 (N_18864,N_18635,N_18557);
xor U18865 (N_18865,N_18658,N_18637);
xor U18866 (N_18866,N_18609,N_18703);
nor U18867 (N_18867,N_18653,N_18514);
or U18868 (N_18868,N_18695,N_18515);
and U18869 (N_18869,N_18644,N_18725);
xnor U18870 (N_18870,N_18579,N_18504);
and U18871 (N_18871,N_18746,N_18511);
xnor U18872 (N_18872,N_18516,N_18731);
xnor U18873 (N_18873,N_18716,N_18529);
nand U18874 (N_18874,N_18585,N_18599);
xnor U18875 (N_18875,N_18583,N_18741);
and U18876 (N_18876,N_18625,N_18693);
and U18877 (N_18877,N_18626,N_18632);
nor U18878 (N_18878,N_18703,N_18651);
or U18879 (N_18879,N_18722,N_18621);
or U18880 (N_18880,N_18643,N_18652);
nand U18881 (N_18881,N_18668,N_18656);
nand U18882 (N_18882,N_18583,N_18688);
nor U18883 (N_18883,N_18689,N_18640);
and U18884 (N_18884,N_18517,N_18519);
and U18885 (N_18885,N_18594,N_18513);
or U18886 (N_18886,N_18536,N_18629);
nand U18887 (N_18887,N_18536,N_18732);
or U18888 (N_18888,N_18662,N_18525);
nor U18889 (N_18889,N_18564,N_18745);
xor U18890 (N_18890,N_18652,N_18724);
nor U18891 (N_18891,N_18622,N_18537);
xor U18892 (N_18892,N_18538,N_18717);
xnor U18893 (N_18893,N_18569,N_18574);
xnor U18894 (N_18894,N_18580,N_18650);
and U18895 (N_18895,N_18551,N_18653);
nand U18896 (N_18896,N_18696,N_18600);
and U18897 (N_18897,N_18523,N_18719);
nor U18898 (N_18898,N_18672,N_18589);
and U18899 (N_18899,N_18583,N_18731);
nand U18900 (N_18900,N_18710,N_18612);
nand U18901 (N_18901,N_18515,N_18627);
nand U18902 (N_18902,N_18707,N_18628);
and U18903 (N_18903,N_18612,N_18625);
and U18904 (N_18904,N_18608,N_18718);
or U18905 (N_18905,N_18565,N_18640);
xnor U18906 (N_18906,N_18567,N_18561);
or U18907 (N_18907,N_18532,N_18551);
and U18908 (N_18908,N_18547,N_18665);
xnor U18909 (N_18909,N_18723,N_18576);
xor U18910 (N_18910,N_18572,N_18513);
nor U18911 (N_18911,N_18506,N_18621);
nand U18912 (N_18912,N_18645,N_18584);
xor U18913 (N_18913,N_18701,N_18514);
nand U18914 (N_18914,N_18621,N_18700);
nor U18915 (N_18915,N_18613,N_18608);
xnor U18916 (N_18916,N_18541,N_18654);
and U18917 (N_18917,N_18669,N_18608);
nand U18918 (N_18918,N_18566,N_18561);
nor U18919 (N_18919,N_18698,N_18574);
nand U18920 (N_18920,N_18730,N_18702);
and U18921 (N_18921,N_18503,N_18616);
and U18922 (N_18922,N_18692,N_18635);
and U18923 (N_18923,N_18508,N_18522);
or U18924 (N_18924,N_18522,N_18538);
or U18925 (N_18925,N_18634,N_18614);
nor U18926 (N_18926,N_18727,N_18646);
and U18927 (N_18927,N_18701,N_18663);
or U18928 (N_18928,N_18695,N_18647);
or U18929 (N_18929,N_18599,N_18575);
nor U18930 (N_18930,N_18610,N_18692);
nor U18931 (N_18931,N_18562,N_18656);
xor U18932 (N_18932,N_18731,N_18602);
and U18933 (N_18933,N_18576,N_18609);
nand U18934 (N_18934,N_18682,N_18663);
nor U18935 (N_18935,N_18693,N_18688);
nand U18936 (N_18936,N_18512,N_18541);
xor U18937 (N_18937,N_18591,N_18665);
nor U18938 (N_18938,N_18505,N_18716);
and U18939 (N_18939,N_18733,N_18633);
xnor U18940 (N_18940,N_18577,N_18557);
and U18941 (N_18941,N_18600,N_18559);
xor U18942 (N_18942,N_18552,N_18704);
xnor U18943 (N_18943,N_18591,N_18695);
xnor U18944 (N_18944,N_18530,N_18688);
nand U18945 (N_18945,N_18728,N_18678);
xor U18946 (N_18946,N_18580,N_18525);
xnor U18947 (N_18947,N_18711,N_18650);
nand U18948 (N_18948,N_18728,N_18550);
and U18949 (N_18949,N_18571,N_18720);
nor U18950 (N_18950,N_18697,N_18537);
or U18951 (N_18951,N_18545,N_18616);
xnor U18952 (N_18952,N_18600,N_18601);
xor U18953 (N_18953,N_18524,N_18547);
or U18954 (N_18954,N_18707,N_18528);
nand U18955 (N_18955,N_18545,N_18585);
xnor U18956 (N_18956,N_18732,N_18679);
xnor U18957 (N_18957,N_18543,N_18690);
nand U18958 (N_18958,N_18669,N_18687);
xnor U18959 (N_18959,N_18674,N_18544);
xor U18960 (N_18960,N_18533,N_18526);
nor U18961 (N_18961,N_18500,N_18557);
nand U18962 (N_18962,N_18731,N_18628);
or U18963 (N_18963,N_18532,N_18738);
or U18964 (N_18964,N_18505,N_18727);
nand U18965 (N_18965,N_18636,N_18591);
nor U18966 (N_18966,N_18575,N_18557);
nor U18967 (N_18967,N_18707,N_18595);
nand U18968 (N_18968,N_18600,N_18553);
nand U18969 (N_18969,N_18564,N_18612);
nor U18970 (N_18970,N_18564,N_18565);
or U18971 (N_18971,N_18553,N_18670);
or U18972 (N_18972,N_18607,N_18653);
xnor U18973 (N_18973,N_18603,N_18665);
nor U18974 (N_18974,N_18543,N_18694);
xnor U18975 (N_18975,N_18626,N_18609);
and U18976 (N_18976,N_18607,N_18647);
and U18977 (N_18977,N_18593,N_18678);
or U18978 (N_18978,N_18586,N_18562);
and U18979 (N_18979,N_18549,N_18571);
nand U18980 (N_18980,N_18512,N_18719);
nand U18981 (N_18981,N_18517,N_18716);
nor U18982 (N_18982,N_18599,N_18722);
xor U18983 (N_18983,N_18676,N_18618);
xnor U18984 (N_18984,N_18544,N_18749);
nor U18985 (N_18985,N_18582,N_18738);
nor U18986 (N_18986,N_18564,N_18644);
xor U18987 (N_18987,N_18539,N_18577);
xor U18988 (N_18988,N_18639,N_18591);
or U18989 (N_18989,N_18628,N_18620);
nand U18990 (N_18990,N_18732,N_18650);
xnor U18991 (N_18991,N_18709,N_18699);
nor U18992 (N_18992,N_18659,N_18547);
or U18993 (N_18993,N_18593,N_18590);
xor U18994 (N_18994,N_18568,N_18682);
xor U18995 (N_18995,N_18611,N_18707);
and U18996 (N_18996,N_18605,N_18623);
and U18997 (N_18997,N_18729,N_18683);
nand U18998 (N_18998,N_18608,N_18586);
or U18999 (N_18999,N_18555,N_18720);
nor U19000 (N_19000,N_18855,N_18909);
nand U19001 (N_19001,N_18854,N_18872);
nor U19002 (N_19002,N_18834,N_18775);
nand U19003 (N_19003,N_18760,N_18924);
nand U19004 (N_19004,N_18891,N_18758);
or U19005 (N_19005,N_18897,N_18797);
nand U19006 (N_19006,N_18824,N_18914);
or U19007 (N_19007,N_18938,N_18860);
nand U19008 (N_19008,N_18935,N_18815);
nor U19009 (N_19009,N_18969,N_18968);
nor U19010 (N_19010,N_18772,N_18754);
nand U19011 (N_19011,N_18894,N_18796);
nor U19012 (N_19012,N_18831,N_18910);
nand U19013 (N_19013,N_18768,N_18987);
nor U19014 (N_19014,N_18845,N_18849);
and U19015 (N_19015,N_18783,N_18823);
and U19016 (N_19016,N_18808,N_18956);
and U19017 (N_19017,N_18840,N_18844);
nor U19018 (N_19018,N_18786,N_18949);
nand U19019 (N_19019,N_18853,N_18753);
xor U19020 (N_19020,N_18936,N_18958);
or U19021 (N_19021,N_18895,N_18792);
xnor U19022 (N_19022,N_18919,N_18920);
nand U19023 (N_19023,N_18795,N_18850);
nand U19024 (N_19024,N_18991,N_18807);
and U19025 (N_19025,N_18877,N_18888);
nor U19026 (N_19026,N_18826,N_18951);
or U19027 (N_19027,N_18986,N_18843);
nand U19028 (N_19028,N_18966,N_18806);
nor U19029 (N_19029,N_18839,N_18751);
or U19030 (N_19030,N_18800,N_18947);
nor U19031 (N_19031,N_18979,N_18982);
nand U19032 (N_19032,N_18945,N_18915);
xor U19033 (N_19033,N_18899,N_18943);
or U19034 (N_19034,N_18798,N_18977);
or U19035 (N_19035,N_18762,N_18925);
and U19036 (N_19036,N_18866,N_18851);
xnor U19037 (N_19037,N_18848,N_18992);
xnor U19038 (N_19038,N_18889,N_18952);
or U19039 (N_19039,N_18903,N_18811);
and U19040 (N_19040,N_18944,N_18862);
and U19041 (N_19041,N_18835,N_18939);
nand U19042 (N_19042,N_18812,N_18856);
nor U19043 (N_19043,N_18882,N_18934);
xor U19044 (N_19044,N_18879,N_18921);
xor U19045 (N_19045,N_18873,N_18801);
nand U19046 (N_19046,N_18993,N_18907);
xnor U19047 (N_19047,N_18918,N_18885);
xor U19048 (N_19048,N_18817,N_18972);
and U19049 (N_19049,N_18861,N_18828);
and U19050 (N_19050,N_18874,N_18809);
xor U19051 (N_19051,N_18859,N_18750);
or U19052 (N_19052,N_18963,N_18931);
and U19053 (N_19053,N_18830,N_18756);
xor U19054 (N_19054,N_18988,N_18832);
nor U19055 (N_19055,N_18959,N_18912);
or U19056 (N_19056,N_18770,N_18876);
xor U19057 (N_19057,N_18766,N_18976);
nor U19058 (N_19058,N_18997,N_18868);
and U19059 (N_19059,N_18759,N_18871);
or U19060 (N_19060,N_18884,N_18774);
or U19061 (N_19061,N_18927,N_18799);
nor U19062 (N_19062,N_18941,N_18793);
and U19063 (N_19063,N_18822,N_18922);
nor U19064 (N_19064,N_18781,N_18755);
nor U19065 (N_19065,N_18869,N_18838);
and U19066 (N_19066,N_18814,N_18932);
or U19067 (N_19067,N_18827,N_18883);
nand U19068 (N_19068,N_18858,N_18820);
nor U19069 (N_19069,N_18779,N_18875);
nor U19070 (N_19070,N_18771,N_18954);
or U19071 (N_19071,N_18886,N_18957);
and U19072 (N_19072,N_18788,N_18930);
nor U19073 (N_19073,N_18752,N_18893);
or U19074 (N_19074,N_18916,N_18990);
nand U19075 (N_19075,N_18777,N_18970);
and U19076 (N_19076,N_18794,N_18892);
nand U19077 (N_19077,N_18898,N_18784);
xor U19078 (N_19078,N_18950,N_18778);
nand U19079 (N_19079,N_18967,N_18785);
and U19080 (N_19080,N_18955,N_18962);
nor U19081 (N_19081,N_18940,N_18802);
nor U19082 (N_19082,N_18761,N_18965);
nand U19083 (N_19083,N_18836,N_18948);
nand U19084 (N_19084,N_18867,N_18863);
or U19085 (N_19085,N_18971,N_18902);
xor U19086 (N_19086,N_18842,N_18870);
nor U19087 (N_19087,N_18782,N_18767);
or U19088 (N_19088,N_18975,N_18923);
and U19089 (N_19089,N_18789,N_18805);
nand U19090 (N_19090,N_18906,N_18887);
nor U19091 (N_19091,N_18881,N_18757);
nor U19092 (N_19092,N_18978,N_18913);
and U19093 (N_19093,N_18937,N_18841);
nor U19094 (N_19094,N_18865,N_18900);
or U19095 (N_19095,N_18787,N_18953);
nor U19096 (N_19096,N_18780,N_18821);
xor U19097 (N_19097,N_18908,N_18880);
nand U19098 (N_19098,N_18996,N_18764);
or U19099 (N_19099,N_18928,N_18960);
or U19100 (N_19100,N_18926,N_18946);
nand U19101 (N_19101,N_18791,N_18929);
and U19102 (N_19102,N_18901,N_18973);
or U19103 (N_19103,N_18857,N_18998);
and U19104 (N_19104,N_18983,N_18829);
xnor U19105 (N_19105,N_18933,N_18911);
nand U19106 (N_19106,N_18810,N_18790);
nand U19107 (N_19107,N_18989,N_18999);
nor U19108 (N_19108,N_18890,N_18763);
nor U19109 (N_19109,N_18904,N_18819);
nor U19110 (N_19110,N_18974,N_18825);
and U19111 (N_19111,N_18776,N_18847);
xor U19112 (N_19112,N_18878,N_18942);
xor U19113 (N_19113,N_18852,N_18813);
or U19114 (N_19114,N_18837,N_18816);
xor U19115 (N_19115,N_18803,N_18964);
and U19116 (N_19116,N_18833,N_18984);
xnor U19117 (N_19117,N_18773,N_18985);
nor U19118 (N_19118,N_18846,N_18917);
nand U19119 (N_19119,N_18994,N_18981);
or U19120 (N_19120,N_18864,N_18995);
xor U19121 (N_19121,N_18961,N_18980);
or U19122 (N_19122,N_18905,N_18765);
nand U19123 (N_19123,N_18818,N_18804);
or U19124 (N_19124,N_18769,N_18896);
nand U19125 (N_19125,N_18821,N_18842);
nor U19126 (N_19126,N_18774,N_18783);
or U19127 (N_19127,N_18832,N_18762);
nor U19128 (N_19128,N_18957,N_18881);
nand U19129 (N_19129,N_18813,N_18806);
and U19130 (N_19130,N_18800,N_18935);
xor U19131 (N_19131,N_18939,N_18825);
nand U19132 (N_19132,N_18914,N_18902);
nor U19133 (N_19133,N_18794,N_18821);
or U19134 (N_19134,N_18800,N_18864);
nand U19135 (N_19135,N_18793,N_18945);
nand U19136 (N_19136,N_18923,N_18841);
and U19137 (N_19137,N_18851,N_18779);
or U19138 (N_19138,N_18865,N_18813);
and U19139 (N_19139,N_18750,N_18970);
nand U19140 (N_19140,N_18857,N_18938);
xor U19141 (N_19141,N_18999,N_18797);
xor U19142 (N_19142,N_18881,N_18909);
xor U19143 (N_19143,N_18763,N_18822);
and U19144 (N_19144,N_18861,N_18887);
nor U19145 (N_19145,N_18786,N_18852);
xor U19146 (N_19146,N_18823,N_18983);
xor U19147 (N_19147,N_18856,N_18750);
xnor U19148 (N_19148,N_18812,N_18991);
and U19149 (N_19149,N_18834,N_18975);
xnor U19150 (N_19150,N_18900,N_18987);
nor U19151 (N_19151,N_18836,N_18870);
or U19152 (N_19152,N_18784,N_18888);
and U19153 (N_19153,N_18971,N_18868);
xor U19154 (N_19154,N_18797,N_18813);
nand U19155 (N_19155,N_18973,N_18892);
xnor U19156 (N_19156,N_18865,N_18987);
and U19157 (N_19157,N_18987,N_18830);
nand U19158 (N_19158,N_18881,N_18933);
nand U19159 (N_19159,N_18771,N_18921);
and U19160 (N_19160,N_18977,N_18860);
nor U19161 (N_19161,N_18889,N_18842);
nand U19162 (N_19162,N_18929,N_18818);
xnor U19163 (N_19163,N_18757,N_18931);
and U19164 (N_19164,N_18786,N_18805);
nor U19165 (N_19165,N_18996,N_18977);
xor U19166 (N_19166,N_18792,N_18852);
or U19167 (N_19167,N_18862,N_18867);
or U19168 (N_19168,N_18771,N_18764);
xnor U19169 (N_19169,N_18835,N_18887);
nand U19170 (N_19170,N_18938,N_18933);
or U19171 (N_19171,N_18759,N_18822);
nand U19172 (N_19172,N_18982,N_18993);
xnor U19173 (N_19173,N_18907,N_18910);
xor U19174 (N_19174,N_18986,N_18844);
and U19175 (N_19175,N_18787,N_18892);
xnor U19176 (N_19176,N_18927,N_18846);
xnor U19177 (N_19177,N_18886,N_18900);
and U19178 (N_19178,N_18989,N_18835);
xor U19179 (N_19179,N_18978,N_18862);
nor U19180 (N_19180,N_18939,N_18966);
xor U19181 (N_19181,N_18887,N_18907);
nand U19182 (N_19182,N_18884,N_18983);
nand U19183 (N_19183,N_18979,N_18866);
xor U19184 (N_19184,N_18860,N_18865);
or U19185 (N_19185,N_18885,N_18805);
or U19186 (N_19186,N_18757,N_18895);
or U19187 (N_19187,N_18832,N_18837);
nor U19188 (N_19188,N_18845,N_18789);
nand U19189 (N_19189,N_18825,N_18868);
and U19190 (N_19190,N_18907,N_18946);
xor U19191 (N_19191,N_18785,N_18855);
and U19192 (N_19192,N_18905,N_18850);
or U19193 (N_19193,N_18864,N_18841);
and U19194 (N_19194,N_18985,N_18762);
nand U19195 (N_19195,N_18922,N_18751);
nor U19196 (N_19196,N_18975,N_18883);
nand U19197 (N_19197,N_18867,N_18947);
nor U19198 (N_19198,N_18944,N_18869);
xor U19199 (N_19199,N_18950,N_18862);
nand U19200 (N_19200,N_18983,N_18820);
and U19201 (N_19201,N_18850,N_18787);
xnor U19202 (N_19202,N_18815,N_18754);
and U19203 (N_19203,N_18863,N_18814);
or U19204 (N_19204,N_18760,N_18895);
or U19205 (N_19205,N_18906,N_18852);
xnor U19206 (N_19206,N_18896,N_18955);
nor U19207 (N_19207,N_18885,N_18838);
xnor U19208 (N_19208,N_18811,N_18787);
and U19209 (N_19209,N_18915,N_18846);
xor U19210 (N_19210,N_18946,N_18866);
nor U19211 (N_19211,N_18840,N_18830);
xnor U19212 (N_19212,N_18872,N_18960);
or U19213 (N_19213,N_18933,N_18854);
nand U19214 (N_19214,N_18759,N_18888);
and U19215 (N_19215,N_18914,N_18968);
nand U19216 (N_19216,N_18942,N_18911);
and U19217 (N_19217,N_18757,N_18996);
or U19218 (N_19218,N_18957,N_18955);
nor U19219 (N_19219,N_18926,N_18848);
xnor U19220 (N_19220,N_18988,N_18975);
nor U19221 (N_19221,N_18841,N_18758);
nand U19222 (N_19222,N_18922,N_18948);
or U19223 (N_19223,N_18894,N_18871);
xnor U19224 (N_19224,N_18830,N_18755);
and U19225 (N_19225,N_18912,N_18815);
nand U19226 (N_19226,N_18802,N_18911);
and U19227 (N_19227,N_18777,N_18933);
nand U19228 (N_19228,N_18826,N_18814);
nor U19229 (N_19229,N_18954,N_18780);
xor U19230 (N_19230,N_18759,N_18795);
xor U19231 (N_19231,N_18774,N_18952);
nor U19232 (N_19232,N_18935,N_18900);
nand U19233 (N_19233,N_18879,N_18763);
xnor U19234 (N_19234,N_18843,N_18944);
xnor U19235 (N_19235,N_18834,N_18957);
xor U19236 (N_19236,N_18767,N_18885);
and U19237 (N_19237,N_18840,N_18771);
and U19238 (N_19238,N_18769,N_18839);
nand U19239 (N_19239,N_18888,N_18902);
nor U19240 (N_19240,N_18829,N_18897);
nand U19241 (N_19241,N_18821,N_18888);
nor U19242 (N_19242,N_18908,N_18940);
and U19243 (N_19243,N_18845,N_18910);
nand U19244 (N_19244,N_18919,N_18953);
and U19245 (N_19245,N_18982,N_18779);
nand U19246 (N_19246,N_18833,N_18977);
and U19247 (N_19247,N_18764,N_18933);
nor U19248 (N_19248,N_18809,N_18966);
nand U19249 (N_19249,N_18875,N_18984);
nor U19250 (N_19250,N_19230,N_19212);
nand U19251 (N_19251,N_19214,N_19139);
xnor U19252 (N_19252,N_19217,N_19131);
and U19253 (N_19253,N_19065,N_19102);
and U19254 (N_19254,N_19016,N_19245);
xnor U19255 (N_19255,N_19152,N_19010);
or U19256 (N_19256,N_19101,N_19035);
or U19257 (N_19257,N_19080,N_19196);
nand U19258 (N_19258,N_19082,N_19054);
nand U19259 (N_19259,N_19206,N_19066);
nand U19260 (N_19260,N_19222,N_19036);
and U19261 (N_19261,N_19165,N_19138);
xnor U19262 (N_19262,N_19110,N_19058);
and U19263 (N_19263,N_19187,N_19098);
and U19264 (N_19264,N_19200,N_19169);
nand U19265 (N_19265,N_19103,N_19225);
and U19266 (N_19266,N_19015,N_19076);
xnor U19267 (N_19267,N_19105,N_19115);
nor U19268 (N_19268,N_19204,N_19155);
nor U19269 (N_19269,N_19123,N_19143);
xor U19270 (N_19270,N_19062,N_19229);
nor U19271 (N_19271,N_19023,N_19224);
or U19272 (N_19272,N_19022,N_19133);
nor U19273 (N_19273,N_19125,N_19072);
and U19274 (N_19274,N_19021,N_19201);
nor U19275 (N_19275,N_19051,N_19060);
nand U19276 (N_19276,N_19176,N_19179);
nor U19277 (N_19277,N_19223,N_19071);
xor U19278 (N_19278,N_19025,N_19033);
or U19279 (N_19279,N_19218,N_19151);
xnor U19280 (N_19280,N_19234,N_19128);
or U19281 (N_19281,N_19113,N_19129);
nand U19282 (N_19282,N_19183,N_19120);
or U19283 (N_19283,N_19091,N_19001);
nand U19284 (N_19284,N_19085,N_19086);
xnor U19285 (N_19285,N_19114,N_19150);
or U19286 (N_19286,N_19092,N_19089);
or U19287 (N_19287,N_19090,N_19029);
nand U19288 (N_19288,N_19147,N_19081);
and U19289 (N_19289,N_19140,N_19167);
or U19290 (N_19290,N_19097,N_19079);
xor U19291 (N_19291,N_19007,N_19148);
and U19292 (N_19292,N_19002,N_19168);
or U19293 (N_19293,N_19043,N_19017);
xnor U19294 (N_19294,N_19039,N_19184);
xnor U19295 (N_19295,N_19059,N_19178);
or U19296 (N_19296,N_19161,N_19160);
or U19297 (N_19297,N_19052,N_19207);
or U19298 (N_19298,N_19240,N_19135);
and U19299 (N_19299,N_19018,N_19117);
or U19300 (N_19300,N_19142,N_19199);
nand U19301 (N_19301,N_19056,N_19162);
and U19302 (N_19302,N_19073,N_19112);
and U19303 (N_19303,N_19188,N_19000);
nand U19304 (N_19304,N_19094,N_19186);
or U19305 (N_19305,N_19070,N_19109);
and U19306 (N_19306,N_19074,N_19239);
or U19307 (N_19307,N_19069,N_19177);
nor U19308 (N_19308,N_19087,N_19045);
nand U19309 (N_19309,N_19173,N_19132);
nand U19310 (N_19310,N_19044,N_19208);
or U19311 (N_19311,N_19158,N_19134);
or U19312 (N_19312,N_19137,N_19159);
or U19313 (N_19313,N_19193,N_19190);
xnor U19314 (N_19314,N_19191,N_19047);
nor U19315 (N_19315,N_19202,N_19198);
nand U19316 (N_19316,N_19020,N_19174);
and U19317 (N_19317,N_19083,N_19028);
or U19318 (N_19318,N_19163,N_19048);
nor U19319 (N_19319,N_19210,N_19149);
or U19320 (N_19320,N_19093,N_19146);
nand U19321 (N_19321,N_19119,N_19096);
xnor U19322 (N_19322,N_19049,N_19050);
and U19323 (N_19323,N_19130,N_19211);
and U19324 (N_19324,N_19205,N_19099);
and U19325 (N_19325,N_19121,N_19171);
nor U19326 (N_19326,N_19100,N_19249);
nor U19327 (N_19327,N_19084,N_19189);
xnor U19328 (N_19328,N_19197,N_19122);
nand U19329 (N_19329,N_19145,N_19013);
xnor U19330 (N_19330,N_19153,N_19216);
nor U19331 (N_19331,N_19172,N_19180);
nor U19332 (N_19332,N_19248,N_19246);
or U19333 (N_19333,N_19116,N_19012);
nor U19334 (N_19334,N_19034,N_19232);
or U19335 (N_19335,N_19008,N_19038);
nand U19336 (N_19336,N_19141,N_19003);
nand U19337 (N_19337,N_19019,N_19136);
nand U19338 (N_19338,N_19068,N_19215);
xor U19339 (N_19339,N_19220,N_19221);
nor U19340 (N_19340,N_19061,N_19118);
nand U19341 (N_19341,N_19027,N_19124);
and U19342 (N_19342,N_19032,N_19213);
nor U19343 (N_19343,N_19107,N_19243);
xor U19344 (N_19344,N_19088,N_19238);
nand U19345 (N_19345,N_19126,N_19209);
xnor U19346 (N_19346,N_19144,N_19233);
xnor U19347 (N_19347,N_19014,N_19077);
or U19348 (N_19348,N_19095,N_19046);
and U19349 (N_19349,N_19235,N_19011);
or U19350 (N_19350,N_19031,N_19236);
or U19351 (N_19351,N_19041,N_19004);
or U19352 (N_19352,N_19005,N_19195);
nor U19353 (N_19353,N_19231,N_19227);
and U19354 (N_19354,N_19064,N_19185);
or U19355 (N_19355,N_19164,N_19181);
nand U19356 (N_19356,N_19111,N_19040);
nor U19357 (N_19357,N_19182,N_19067);
and U19358 (N_19358,N_19237,N_19053);
and U19359 (N_19359,N_19228,N_19106);
nand U19360 (N_19360,N_19127,N_19192);
nor U19361 (N_19361,N_19055,N_19244);
or U19362 (N_19362,N_19203,N_19241);
xor U19363 (N_19363,N_19156,N_19226);
and U19364 (N_19364,N_19042,N_19037);
or U19365 (N_19365,N_19175,N_19078);
nor U19366 (N_19366,N_19075,N_19170);
nor U19367 (N_19367,N_19247,N_19242);
or U19368 (N_19368,N_19063,N_19030);
and U19369 (N_19369,N_19006,N_19157);
and U19370 (N_19370,N_19057,N_19219);
nor U19371 (N_19371,N_19104,N_19024);
nand U19372 (N_19372,N_19154,N_19009);
and U19373 (N_19373,N_19026,N_19108);
or U19374 (N_19374,N_19166,N_19194);
nand U19375 (N_19375,N_19014,N_19041);
or U19376 (N_19376,N_19021,N_19185);
or U19377 (N_19377,N_19180,N_19024);
or U19378 (N_19378,N_19070,N_19098);
nor U19379 (N_19379,N_19046,N_19120);
and U19380 (N_19380,N_19234,N_19088);
xnor U19381 (N_19381,N_19084,N_19055);
xor U19382 (N_19382,N_19110,N_19217);
and U19383 (N_19383,N_19025,N_19188);
xnor U19384 (N_19384,N_19212,N_19046);
nor U19385 (N_19385,N_19163,N_19085);
nand U19386 (N_19386,N_19184,N_19081);
and U19387 (N_19387,N_19159,N_19090);
or U19388 (N_19388,N_19095,N_19085);
nor U19389 (N_19389,N_19125,N_19033);
and U19390 (N_19390,N_19070,N_19023);
nor U19391 (N_19391,N_19166,N_19159);
nand U19392 (N_19392,N_19084,N_19143);
xor U19393 (N_19393,N_19015,N_19196);
nor U19394 (N_19394,N_19212,N_19055);
or U19395 (N_19395,N_19210,N_19136);
nor U19396 (N_19396,N_19109,N_19105);
nand U19397 (N_19397,N_19183,N_19100);
nor U19398 (N_19398,N_19145,N_19064);
nor U19399 (N_19399,N_19225,N_19074);
xor U19400 (N_19400,N_19164,N_19204);
and U19401 (N_19401,N_19233,N_19171);
xor U19402 (N_19402,N_19101,N_19190);
xnor U19403 (N_19403,N_19108,N_19064);
nand U19404 (N_19404,N_19116,N_19022);
and U19405 (N_19405,N_19007,N_19221);
nor U19406 (N_19406,N_19016,N_19083);
or U19407 (N_19407,N_19180,N_19205);
or U19408 (N_19408,N_19231,N_19169);
nor U19409 (N_19409,N_19207,N_19054);
nand U19410 (N_19410,N_19152,N_19187);
nand U19411 (N_19411,N_19033,N_19225);
nor U19412 (N_19412,N_19003,N_19060);
or U19413 (N_19413,N_19055,N_19165);
xnor U19414 (N_19414,N_19158,N_19051);
nor U19415 (N_19415,N_19161,N_19142);
xnor U19416 (N_19416,N_19044,N_19242);
nor U19417 (N_19417,N_19211,N_19215);
nor U19418 (N_19418,N_19117,N_19179);
nor U19419 (N_19419,N_19073,N_19024);
xnor U19420 (N_19420,N_19202,N_19145);
or U19421 (N_19421,N_19104,N_19050);
nor U19422 (N_19422,N_19110,N_19026);
nor U19423 (N_19423,N_19236,N_19044);
nor U19424 (N_19424,N_19053,N_19213);
or U19425 (N_19425,N_19030,N_19248);
nand U19426 (N_19426,N_19118,N_19181);
or U19427 (N_19427,N_19142,N_19042);
xnor U19428 (N_19428,N_19159,N_19174);
nor U19429 (N_19429,N_19107,N_19037);
nor U19430 (N_19430,N_19125,N_19216);
xor U19431 (N_19431,N_19149,N_19213);
and U19432 (N_19432,N_19041,N_19032);
and U19433 (N_19433,N_19001,N_19074);
xor U19434 (N_19434,N_19192,N_19156);
nor U19435 (N_19435,N_19070,N_19041);
and U19436 (N_19436,N_19089,N_19117);
and U19437 (N_19437,N_19018,N_19060);
nand U19438 (N_19438,N_19207,N_19186);
or U19439 (N_19439,N_19002,N_19131);
and U19440 (N_19440,N_19079,N_19036);
and U19441 (N_19441,N_19239,N_19090);
or U19442 (N_19442,N_19016,N_19142);
or U19443 (N_19443,N_19129,N_19059);
xnor U19444 (N_19444,N_19104,N_19120);
and U19445 (N_19445,N_19191,N_19001);
or U19446 (N_19446,N_19118,N_19157);
xnor U19447 (N_19447,N_19024,N_19172);
or U19448 (N_19448,N_19049,N_19115);
nor U19449 (N_19449,N_19200,N_19217);
nand U19450 (N_19450,N_19219,N_19146);
and U19451 (N_19451,N_19222,N_19220);
nand U19452 (N_19452,N_19147,N_19244);
and U19453 (N_19453,N_19070,N_19137);
nand U19454 (N_19454,N_19230,N_19056);
nand U19455 (N_19455,N_19115,N_19119);
and U19456 (N_19456,N_19214,N_19044);
and U19457 (N_19457,N_19029,N_19097);
or U19458 (N_19458,N_19212,N_19106);
nand U19459 (N_19459,N_19035,N_19107);
nor U19460 (N_19460,N_19218,N_19027);
nor U19461 (N_19461,N_19183,N_19037);
nand U19462 (N_19462,N_19038,N_19210);
xnor U19463 (N_19463,N_19238,N_19222);
nor U19464 (N_19464,N_19133,N_19128);
or U19465 (N_19465,N_19153,N_19026);
nand U19466 (N_19466,N_19037,N_19127);
and U19467 (N_19467,N_19029,N_19214);
or U19468 (N_19468,N_19189,N_19208);
and U19469 (N_19469,N_19223,N_19015);
nand U19470 (N_19470,N_19249,N_19085);
nor U19471 (N_19471,N_19206,N_19245);
nor U19472 (N_19472,N_19008,N_19080);
nor U19473 (N_19473,N_19172,N_19198);
xnor U19474 (N_19474,N_19140,N_19031);
and U19475 (N_19475,N_19192,N_19218);
nor U19476 (N_19476,N_19046,N_19118);
nor U19477 (N_19477,N_19149,N_19066);
or U19478 (N_19478,N_19093,N_19054);
nand U19479 (N_19479,N_19102,N_19094);
nand U19480 (N_19480,N_19181,N_19238);
nor U19481 (N_19481,N_19054,N_19100);
nor U19482 (N_19482,N_19089,N_19017);
or U19483 (N_19483,N_19066,N_19071);
nand U19484 (N_19484,N_19211,N_19056);
and U19485 (N_19485,N_19046,N_19021);
nand U19486 (N_19486,N_19053,N_19192);
nand U19487 (N_19487,N_19130,N_19036);
xnor U19488 (N_19488,N_19128,N_19227);
xnor U19489 (N_19489,N_19152,N_19035);
nand U19490 (N_19490,N_19088,N_19231);
or U19491 (N_19491,N_19060,N_19150);
xor U19492 (N_19492,N_19027,N_19214);
nand U19493 (N_19493,N_19105,N_19018);
or U19494 (N_19494,N_19184,N_19137);
nor U19495 (N_19495,N_19168,N_19133);
xnor U19496 (N_19496,N_19234,N_19025);
nor U19497 (N_19497,N_19013,N_19236);
or U19498 (N_19498,N_19103,N_19122);
or U19499 (N_19499,N_19166,N_19054);
and U19500 (N_19500,N_19313,N_19285);
nand U19501 (N_19501,N_19414,N_19418);
nor U19502 (N_19502,N_19318,N_19413);
xor U19503 (N_19503,N_19251,N_19254);
nand U19504 (N_19504,N_19462,N_19306);
xor U19505 (N_19505,N_19334,N_19496);
and U19506 (N_19506,N_19278,N_19329);
nand U19507 (N_19507,N_19384,N_19335);
and U19508 (N_19508,N_19386,N_19304);
xnor U19509 (N_19509,N_19288,N_19398);
nand U19510 (N_19510,N_19373,N_19488);
or U19511 (N_19511,N_19379,N_19308);
nor U19512 (N_19512,N_19456,N_19368);
nand U19513 (N_19513,N_19467,N_19475);
nand U19514 (N_19514,N_19487,N_19339);
nand U19515 (N_19515,N_19393,N_19265);
nor U19516 (N_19516,N_19319,N_19438);
or U19517 (N_19517,N_19415,N_19473);
nor U19518 (N_19518,N_19471,N_19321);
nand U19519 (N_19519,N_19419,N_19345);
xnor U19520 (N_19520,N_19253,N_19469);
and U19521 (N_19521,N_19344,N_19294);
or U19522 (N_19522,N_19341,N_19410);
or U19523 (N_19523,N_19360,N_19390);
xnor U19524 (N_19524,N_19424,N_19315);
and U19525 (N_19525,N_19264,N_19355);
and U19526 (N_19526,N_19406,N_19397);
or U19527 (N_19527,N_19352,N_19351);
nor U19528 (N_19528,N_19396,N_19317);
nand U19529 (N_19529,N_19322,N_19311);
or U19530 (N_19530,N_19391,N_19457);
xnor U19531 (N_19531,N_19331,N_19439);
or U19532 (N_19532,N_19299,N_19286);
nand U19533 (N_19533,N_19484,N_19409);
or U19534 (N_19534,N_19483,N_19284);
xnor U19535 (N_19535,N_19270,N_19283);
nor U19536 (N_19536,N_19408,N_19272);
nor U19537 (N_19537,N_19463,N_19369);
or U19538 (N_19538,N_19403,N_19287);
xnor U19539 (N_19539,N_19383,N_19482);
xnor U19540 (N_19540,N_19411,N_19432);
nor U19541 (N_19541,N_19450,N_19486);
and U19542 (N_19542,N_19443,N_19275);
nor U19543 (N_19543,N_19374,N_19455);
nand U19544 (N_19544,N_19367,N_19250);
nor U19545 (N_19545,N_19333,N_19256);
nand U19546 (N_19546,N_19326,N_19387);
and U19547 (N_19547,N_19301,N_19466);
nand U19548 (N_19548,N_19421,N_19268);
xnor U19549 (N_19549,N_19320,N_19499);
xnor U19550 (N_19550,N_19485,N_19402);
and U19551 (N_19551,N_19293,N_19312);
nand U19552 (N_19552,N_19337,N_19479);
xnor U19553 (N_19553,N_19343,N_19423);
xnor U19554 (N_19554,N_19420,N_19495);
nand U19555 (N_19555,N_19266,N_19362);
and U19556 (N_19556,N_19290,N_19428);
nand U19557 (N_19557,N_19459,N_19426);
xnor U19558 (N_19558,N_19282,N_19489);
nand U19559 (N_19559,N_19273,N_19399);
and U19560 (N_19560,N_19356,N_19444);
and U19561 (N_19561,N_19472,N_19279);
nand U19562 (N_19562,N_19468,N_19447);
nor U19563 (N_19563,N_19461,N_19381);
and U19564 (N_19564,N_19255,N_19493);
nor U19565 (N_19565,N_19477,N_19258);
or U19566 (N_19566,N_19276,N_19429);
xnor U19567 (N_19567,N_19371,N_19470);
and U19568 (N_19568,N_19372,N_19323);
and U19569 (N_19569,N_19385,N_19417);
xor U19570 (N_19570,N_19303,N_19349);
and U19571 (N_19571,N_19347,N_19454);
nand U19572 (N_19572,N_19401,N_19353);
nand U19573 (N_19573,N_19382,N_19434);
and U19574 (N_19574,N_19328,N_19442);
nor U19575 (N_19575,N_19464,N_19404);
xnor U19576 (N_19576,N_19370,N_19252);
nand U19577 (N_19577,N_19325,N_19448);
and U19578 (N_19578,N_19378,N_19274);
nand U19579 (N_19579,N_19269,N_19476);
nor U19580 (N_19580,N_19412,N_19297);
nor U19581 (N_19581,N_19376,N_19332);
or U19582 (N_19582,N_19395,N_19458);
xnor U19583 (N_19583,N_19261,N_19480);
nor U19584 (N_19584,N_19375,N_19316);
nand U19585 (N_19585,N_19310,N_19305);
or U19586 (N_19586,N_19291,N_19405);
or U19587 (N_19587,N_19346,N_19289);
nor U19588 (N_19588,N_19400,N_19357);
xor U19589 (N_19589,N_19430,N_19281);
or U19590 (N_19590,N_19338,N_19474);
and U19591 (N_19591,N_19452,N_19365);
xor U19592 (N_19592,N_19300,N_19497);
nor U19593 (N_19593,N_19262,N_19358);
and U19594 (N_19594,N_19465,N_19340);
and U19595 (N_19595,N_19478,N_19435);
nand U19596 (N_19596,N_19361,N_19263);
nor U19597 (N_19597,N_19498,N_19431);
xnor U19598 (N_19598,N_19441,N_19388);
and U19599 (N_19599,N_19446,N_19491);
or U19600 (N_19600,N_19425,N_19307);
nor U19601 (N_19601,N_19348,N_19257);
and U19602 (N_19602,N_19259,N_19336);
nor U19603 (N_19603,N_19377,N_19492);
xnor U19604 (N_19604,N_19359,N_19392);
and U19605 (N_19605,N_19314,N_19451);
nor U19606 (N_19606,N_19394,N_19277);
and U19607 (N_19607,N_19280,N_19422);
nor U19608 (N_19608,N_19302,N_19296);
nand U19609 (N_19609,N_19437,N_19298);
nor U19610 (N_19610,N_19324,N_19453);
xnor U19611 (N_19611,N_19267,N_19260);
nor U19612 (N_19612,N_19342,N_19309);
xnor U19613 (N_19613,N_19327,N_19427);
or U19614 (N_19614,N_19407,N_19364);
or U19615 (N_19615,N_19460,N_19481);
xor U19616 (N_19616,N_19436,N_19445);
or U19617 (N_19617,N_19350,N_19295);
nand U19618 (N_19618,N_19389,N_19292);
xor U19619 (N_19619,N_19440,N_19271);
and U19620 (N_19620,N_19366,N_19354);
nor U19621 (N_19621,N_19380,N_19449);
xnor U19622 (N_19622,N_19330,N_19363);
and U19623 (N_19623,N_19490,N_19416);
xor U19624 (N_19624,N_19494,N_19433);
or U19625 (N_19625,N_19295,N_19482);
nand U19626 (N_19626,N_19324,N_19316);
nor U19627 (N_19627,N_19336,N_19452);
nor U19628 (N_19628,N_19357,N_19264);
or U19629 (N_19629,N_19426,N_19316);
xnor U19630 (N_19630,N_19486,N_19421);
nor U19631 (N_19631,N_19359,N_19496);
xnor U19632 (N_19632,N_19411,N_19297);
nor U19633 (N_19633,N_19458,N_19304);
or U19634 (N_19634,N_19477,N_19337);
nand U19635 (N_19635,N_19270,N_19452);
and U19636 (N_19636,N_19470,N_19468);
and U19637 (N_19637,N_19322,N_19286);
nor U19638 (N_19638,N_19477,N_19362);
nand U19639 (N_19639,N_19416,N_19415);
xor U19640 (N_19640,N_19472,N_19459);
and U19641 (N_19641,N_19399,N_19254);
and U19642 (N_19642,N_19396,N_19463);
xor U19643 (N_19643,N_19485,N_19253);
xnor U19644 (N_19644,N_19400,N_19470);
and U19645 (N_19645,N_19403,N_19405);
nor U19646 (N_19646,N_19400,N_19431);
nand U19647 (N_19647,N_19487,N_19419);
or U19648 (N_19648,N_19496,N_19336);
nand U19649 (N_19649,N_19464,N_19421);
nand U19650 (N_19650,N_19399,N_19428);
xnor U19651 (N_19651,N_19433,N_19480);
or U19652 (N_19652,N_19363,N_19433);
nor U19653 (N_19653,N_19432,N_19426);
xor U19654 (N_19654,N_19278,N_19286);
or U19655 (N_19655,N_19415,N_19254);
or U19656 (N_19656,N_19413,N_19322);
or U19657 (N_19657,N_19332,N_19284);
or U19658 (N_19658,N_19285,N_19260);
nor U19659 (N_19659,N_19421,N_19319);
xnor U19660 (N_19660,N_19282,N_19264);
nand U19661 (N_19661,N_19382,N_19412);
nor U19662 (N_19662,N_19292,N_19483);
nand U19663 (N_19663,N_19342,N_19473);
and U19664 (N_19664,N_19256,N_19486);
xnor U19665 (N_19665,N_19314,N_19287);
and U19666 (N_19666,N_19478,N_19461);
xor U19667 (N_19667,N_19391,N_19399);
xor U19668 (N_19668,N_19444,N_19285);
nor U19669 (N_19669,N_19496,N_19403);
and U19670 (N_19670,N_19390,N_19352);
and U19671 (N_19671,N_19318,N_19358);
nand U19672 (N_19672,N_19255,N_19366);
xor U19673 (N_19673,N_19325,N_19405);
nand U19674 (N_19674,N_19346,N_19302);
xor U19675 (N_19675,N_19298,N_19276);
xor U19676 (N_19676,N_19266,N_19460);
nor U19677 (N_19677,N_19415,N_19448);
or U19678 (N_19678,N_19307,N_19433);
and U19679 (N_19679,N_19294,N_19487);
xor U19680 (N_19680,N_19429,N_19285);
xor U19681 (N_19681,N_19437,N_19436);
and U19682 (N_19682,N_19405,N_19374);
nand U19683 (N_19683,N_19252,N_19366);
xor U19684 (N_19684,N_19385,N_19444);
nor U19685 (N_19685,N_19396,N_19433);
nand U19686 (N_19686,N_19371,N_19448);
or U19687 (N_19687,N_19376,N_19350);
nand U19688 (N_19688,N_19475,N_19385);
and U19689 (N_19689,N_19440,N_19486);
and U19690 (N_19690,N_19469,N_19311);
or U19691 (N_19691,N_19297,N_19359);
and U19692 (N_19692,N_19343,N_19307);
nand U19693 (N_19693,N_19269,N_19344);
or U19694 (N_19694,N_19326,N_19372);
nor U19695 (N_19695,N_19461,N_19314);
and U19696 (N_19696,N_19324,N_19252);
nor U19697 (N_19697,N_19397,N_19272);
xnor U19698 (N_19698,N_19319,N_19423);
or U19699 (N_19699,N_19284,N_19360);
nand U19700 (N_19700,N_19260,N_19488);
nand U19701 (N_19701,N_19324,N_19422);
nor U19702 (N_19702,N_19402,N_19419);
xnor U19703 (N_19703,N_19334,N_19384);
or U19704 (N_19704,N_19309,N_19351);
nand U19705 (N_19705,N_19431,N_19284);
or U19706 (N_19706,N_19256,N_19493);
nand U19707 (N_19707,N_19322,N_19354);
or U19708 (N_19708,N_19384,N_19273);
nor U19709 (N_19709,N_19491,N_19356);
nor U19710 (N_19710,N_19383,N_19382);
nand U19711 (N_19711,N_19345,N_19375);
nor U19712 (N_19712,N_19324,N_19499);
nor U19713 (N_19713,N_19318,N_19268);
or U19714 (N_19714,N_19481,N_19418);
nor U19715 (N_19715,N_19466,N_19290);
or U19716 (N_19716,N_19292,N_19405);
and U19717 (N_19717,N_19328,N_19404);
xor U19718 (N_19718,N_19402,N_19478);
nand U19719 (N_19719,N_19322,N_19406);
and U19720 (N_19720,N_19264,N_19371);
or U19721 (N_19721,N_19262,N_19449);
nand U19722 (N_19722,N_19393,N_19434);
nand U19723 (N_19723,N_19252,N_19346);
and U19724 (N_19724,N_19388,N_19351);
or U19725 (N_19725,N_19484,N_19404);
xnor U19726 (N_19726,N_19496,N_19444);
and U19727 (N_19727,N_19499,N_19359);
nand U19728 (N_19728,N_19476,N_19291);
or U19729 (N_19729,N_19360,N_19374);
or U19730 (N_19730,N_19478,N_19357);
and U19731 (N_19731,N_19288,N_19381);
xor U19732 (N_19732,N_19252,N_19389);
or U19733 (N_19733,N_19405,N_19486);
nor U19734 (N_19734,N_19283,N_19346);
or U19735 (N_19735,N_19342,N_19460);
and U19736 (N_19736,N_19278,N_19267);
and U19737 (N_19737,N_19466,N_19277);
or U19738 (N_19738,N_19447,N_19388);
or U19739 (N_19739,N_19360,N_19419);
nor U19740 (N_19740,N_19468,N_19386);
nand U19741 (N_19741,N_19401,N_19495);
nand U19742 (N_19742,N_19395,N_19353);
nand U19743 (N_19743,N_19303,N_19483);
nand U19744 (N_19744,N_19319,N_19275);
xor U19745 (N_19745,N_19394,N_19462);
or U19746 (N_19746,N_19478,N_19254);
and U19747 (N_19747,N_19250,N_19483);
nand U19748 (N_19748,N_19337,N_19315);
nor U19749 (N_19749,N_19263,N_19465);
xor U19750 (N_19750,N_19633,N_19589);
nand U19751 (N_19751,N_19733,N_19556);
xnor U19752 (N_19752,N_19585,N_19545);
or U19753 (N_19753,N_19628,N_19703);
and U19754 (N_19754,N_19564,N_19739);
nor U19755 (N_19755,N_19503,N_19664);
nor U19756 (N_19756,N_19587,N_19504);
or U19757 (N_19757,N_19672,N_19525);
or U19758 (N_19758,N_19653,N_19594);
and U19759 (N_19759,N_19658,N_19674);
xnor U19760 (N_19760,N_19668,N_19605);
xor U19761 (N_19761,N_19573,N_19670);
nand U19762 (N_19762,N_19530,N_19574);
or U19763 (N_19763,N_19527,N_19519);
nor U19764 (N_19764,N_19738,N_19735);
nor U19765 (N_19765,N_19533,N_19600);
nor U19766 (N_19766,N_19637,N_19655);
nor U19767 (N_19767,N_19540,N_19693);
nor U19768 (N_19768,N_19714,N_19511);
nand U19769 (N_19769,N_19725,N_19713);
or U19770 (N_19770,N_19706,N_19737);
xor U19771 (N_19771,N_19727,N_19705);
and U19772 (N_19772,N_19623,N_19528);
or U19773 (N_19773,N_19669,N_19534);
and U19774 (N_19774,N_19657,N_19609);
nand U19775 (N_19775,N_19690,N_19515);
xnor U19776 (N_19776,N_19665,N_19698);
nor U19777 (N_19777,N_19570,N_19671);
nor U19778 (N_19778,N_19513,N_19648);
or U19779 (N_19779,N_19567,N_19640);
xnor U19780 (N_19780,N_19514,N_19641);
nor U19781 (N_19781,N_19501,N_19744);
nand U19782 (N_19782,N_19638,N_19678);
xor U19783 (N_19783,N_19632,N_19734);
or U19784 (N_19784,N_19679,N_19569);
xor U19785 (N_19785,N_19539,N_19711);
and U19786 (N_19786,N_19673,N_19741);
xnor U19787 (N_19787,N_19720,N_19607);
nand U19788 (N_19788,N_19526,N_19661);
nor U19789 (N_19789,N_19715,N_19645);
nor U19790 (N_19790,N_19561,N_19659);
xnor U19791 (N_19791,N_19642,N_19537);
or U19792 (N_19792,N_19746,N_19520);
and U19793 (N_19793,N_19508,N_19676);
xnor U19794 (N_19794,N_19553,N_19522);
xnor U19795 (N_19795,N_19736,N_19516);
and U19796 (N_19796,N_19684,N_19704);
nor U19797 (N_19797,N_19718,N_19524);
and U19798 (N_19798,N_19549,N_19689);
nand U19799 (N_19799,N_19575,N_19546);
xor U19800 (N_19800,N_19617,N_19536);
nor U19801 (N_19801,N_19558,N_19675);
nand U19802 (N_19802,N_19651,N_19506);
or U19803 (N_19803,N_19708,N_19700);
nor U19804 (N_19804,N_19505,N_19635);
and U19805 (N_19805,N_19745,N_19723);
or U19806 (N_19806,N_19572,N_19680);
nor U19807 (N_19807,N_19709,N_19716);
nor U19808 (N_19808,N_19721,N_19611);
nor U19809 (N_19809,N_19604,N_19691);
nand U19810 (N_19810,N_19666,N_19612);
and U19811 (N_19811,N_19624,N_19729);
or U19812 (N_19812,N_19634,N_19603);
or U19813 (N_19813,N_19697,N_19608);
and U19814 (N_19814,N_19582,N_19548);
nand U19815 (N_19815,N_19688,N_19584);
and U19816 (N_19816,N_19593,N_19749);
and U19817 (N_19817,N_19580,N_19523);
or U19818 (N_19818,N_19500,N_19701);
and U19819 (N_19819,N_19719,N_19748);
or U19820 (N_19820,N_19654,N_19686);
nor U19821 (N_19821,N_19578,N_19592);
or U19822 (N_19822,N_19629,N_19728);
or U19823 (N_19823,N_19535,N_19557);
xnor U19824 (N_19824,N_19597,N_19591);
nor U19825 (N_19825,N_19620,N_19588);
and U19826 (N_19826,N_19712,N_19656);
xor U19827 (N_19827,N_19724,N_19542);
nor U19828 (N_19828,N_19732,N_19627);
or U19829 (N_19829,N_19644,N_19507);
xnor U19830 (N_19830,N_19742,N_19643);
nor U19831 (N_19831,N_19681,N_19560);
xor U19832 (N_19832,N_19650,N_19631);
nor U19833 (N_19833,N_19565,N_19613);
or U19834 (N_19834,N_19717,N_19529);
nor U19835 (N_19835,N_19707,N_19722);
and U19836 (N_19836,N_19531,N_19646);
xnor U19837 (N_19837,N_19677,N_19596);
nor U19838 (N_19838,N_19509,N_19625);
nor U19839 (N_19839,N_19660,N_19598);
nand U19840 (N_19840,N_19639,N_19581);
or U19841 (N_19841,N_19630,N_19614);
nand U19842 (N_19842,N_19626,N_19583);
or U19843 (N_19843,N_19610,N_19521);
nor U19844 (N_19844,N_19579,N_19682);
or U19845 (N_19845,N_19696,N_19554);
nor U19846 (N_19846,N_19667,N_19518);
nor U19847 (N_19847,N_19694,N_19571);
or U19848 (N_19848,N_19622,N_19619);
nand U19849 (N_19849,N_19606,N_19544);
or U19850 (N_19850,N_19702,N_19685);
nand U19851 (N_19851,N_19595,N_19618);
or U19852 (N_19852,N_19543,N_19555);
nor U19853 (N_19853,N_19683,N_19502);
nor U19854 (N_19854,N_19662,N_19586);
nor U19855 (N_19855,N_19647,N_19747);
xnor U19856 (N_19856,N_19551,N_19621);
or U19857 (N_19857,N_19636,N_19652);
xnor U19858 (N_19858,N_19550,N_19552);
xnor U19859 (N_19859,N_19730,N_19740);
nand U19860 (N_19860,N_19692,N_19726);
or U19861 (N_19861,N_19731,N_19562);
nor U19862 (N_19862,N_19616,N_19576);
and U19863 (N_19863,N_19601,N_19699);
nor U19864 (N_19864,N_19559,N_19695);
or U19865 (N_19865,N_19615,N_19710);
nand U19866 (N_19866,N_19602,N_19649);
xnor U19867 (N_19867,N_19590,N_19743);
xor U19868 (N_19868,N_19538,N_19547);
xor U19869 (N_19869,N_19563,N_19577);
nor U19870 (N_19870,N_19517,N_19687);
xnor U19871 (N_19871,N_19663,N_19510);
or U19872 (N_19872,N_19512,N_19532);
xor U19873 (N_19873,N_19541,N_19566);
xor U19874 (N_19874,N_19599,N_19568);
nor U19875 (N_19875,N_19569,N_19579);
and U19876 (N_19876,N_19659,N_19558);
nand U19877 (N_19877,N_19708,N_19693);
nor U19878 (N_19878,N_19508,N_19705);
nand U19879 (N_19879,N_19619,N_19748);
nand U19880 (N_19880,N_19659,N_19532);
or U19881 (N_19881,N_19713,N_19667);
xnor U19882 (N_19882,N_19620,N_19677);
and U19883 (N_19883,N_19684,N_19601);
nand U19884 (N_19884,N_19570,N_19687);
xor U19885 (N_19885,N_19676,N_19683);
nand U19886 (N_19886,N_19591,N_19677);
nor U19887 (N_19887,N_19647,N_19557);
and U19888 (N_19888,N_19706,N_19542);
and U19889 (N_19889,N_19695,N_19548);
xnor U19890 (N_19890,N_19746,N_19528);
nand U19891 (N_19891,N_19719,N_19739);
xor U19892 (N_19892,N_19542,N_19738);
or U19893 (N_19893,N_19644,N_19621);
or U19894 (N_19894,N_19622,N_19516);
nor U19895 (N_19895,N_19531,N_19734);
nor U19896 (N_19896,N_19584,N_19617);
nand U19897 (N_19897,N_19542,N_19565);
nor U19898 (N_19898,N_19657,N_19692);
or U19899 (N_19899,N_19619,N_19580);
xor U19900 (N_19900,N_19559,N_19701);
and U19901 (N_19901,N_19531,N_19610);
nand U19902 (N_19902,N_19518,N_19574);
nor U19903 (N_19903,N_19703,N_19664);
xor U19904 (N_19904,N_19682,N_19598);
nor U19905 (N_19905,N_19661,N_19549);
nor U19906 (N_19906,N_19678,N_19550);
nor U19907 (N_19907,N_19726,N_19639);
xor U19908 (N_19908,N_19625,N_19504);
nor U19909 (N_19909,N_19738,N_19558);
nor U19910 (N_19910,N_19534,N_19704);
xnor U19911 (N_19911,N_19540,N_19591);
nand U19912 (N_19912,N_19543,N_19662);
or U19913 (N_19913,N_19639,N_19728);
xor U19914 (N_19914,N_19588,N_19650);
nand U19915 (N_19915,N_19668,N_19696);
nand U19916 (N_19916,N_19593,N_19502);
or U19917 (N_19917,N_19602,N_19670);
xor U19918 (N_19918,N_19646,N_19553);
nor U19919 (N_19919,N_19584,N_19579);
and U19920 (N_19920,N_19742,N_19560);
and U19921 (N_19921,N_19704,N_19526);
nor U19922 (N_19922,N_19635,N_19699);
nor U19923 (N_19923,N_19747,N_19544);
or U19924 (N_19924,N_19548,N_19664);
xor U19925 (N_19925,N_19542,N_19536);
nor U19926 (N_19926,N_19548,N_19530);
and U19927 (N_19927,N_19513,N_19642);
xor U19928 (N_19928,N_19618,N_19704);
nand U19929 (N_19929,N_19614,N_19723);
nor U19930 (N_19930,N_19534,N_19700);
or U19931 (N_19931,N_19630,N_19532);
or U19932 (N_19932,N_19745,N_19634);
xnor U19933 (N_19933,N_19724,N_19602);
and U19934 (N_19934,N_19572,N_19708);
and U19935 (N_19935,N_19516,N_19526);
nand U19936 (N_19936,N_19738,N_19684);
xor U19937 (N_19937,N_19527,N_19699);
nand U19938 (N_19938,N_19649,N_19509);
nand U19939 (N_19939,N_19634,N_19612);
and U19940 (N_19940,N_19500,N_19629);
and U19941 (N_19941,N_19706,N_19748);
xnor U19942 (N_19942,N_19507,N_19535);
xor U19943 (N_19943,N_19744,N_19542);
or U19944 (N_19944,N_19635,N_19581);
xor U19945 (N_19945,N_19681,N_19620);
and U19946 (N_19946,N_19645,N_19553);
nor U19947 (N_19947,N_19655,N_19713);
nor U19948 (N_19948,N_19554,N_19709);
xnor U19949 (N_19949,N_19550,N_19595);
and U19950 (N_19950,N_19557,N_19586);
or U19951 (N_19951,N_19642,N_19637);
nor U19952 (N_19952,N_19531,N_19723);
nor U19953 (N_19953,N_19531,N_19577);
and U19954 (N_19954,N_19502,N_19656);
nand U19955 (N_19955,N_19690,N_19680);
or U19956 (N_19956,N_19668,N_19708);
and U19957 (N_19957,N_19684,N_19554);
nand U19958 (N_19958,N_19519,N_19720);
nand U19959 (N_19959,N_19512,N_19553);
and U19960 (N_19960,N_19663,N_19512);
or U19961 (N_19961,N_19595,N_19699);
and U19962 (N_19962,N_19514,N_19693);
or U19963 (N_19963,N_19685,N_19697);
or U19964 (N_19964,N_19681,N_19532);
or U19965 (N_19965,N_19620,N_19727);
and U19966 (N_19966,N_19701,N_19518);
and U19967 (N_19967,N_19728,N_19542);
nand U19968 (N_19968,N_19619,N_19663);
nand U19969 (N_19969,N_19527,N_19649);
or U19970 (N_19970,N_19596,N_19594);
or U19971 (N_19971,N_19731,N_19529);
and U19972 (N_19972,N_19650,N_19576);
and U19973 (N_19973,N_19509,N_19603);
xor U19974 (N_19974,N_19702,N_19512);
xnor U19975 (N_19975,N_19604,N_19605);
and U19976 (N_19976,N_19560,N_19614);
or U19977 (N_19977,N_19721,N_19679);
or U19978 (N_19978,N_19529,N_19635);
or U19979 (N_19979,N_19691,N_19583);
xnor U19980 (N_19980,N_19598,N_19608);
and U19981 (N_19981,N_19650,N_19626);
or U19982 (N_19982,N_19706,N_19699);
or U19983 (N_19983,N_19600,N_19530);
or U19984 (N_19984,N_19660,N_19595);
and U19985 (N_19985,N_19522,N_19742);
nor U19986 (N_19986,N_19559,N_19703);
xnor U19987 (N_19987,N_19566,N_19657);
nor U19988 (N_19988,N_19703,N_19690);
or U19989 (N_19989,N_19619,N_19698);
nand U19990 (N_19990,N_19554,N_19513);
nor U19991 (N_19991,N_19610,N_19745);
and U19992 (N_19992,N_19618,N_19672);
nor U19993 (N_19993,N_19618,N_19655);
or U19994 (N_19994,N_19644,N_19537);
or U19995 (N_19995,N_19696,N_19719);
xnor U19996 (N_19996,N_19571,N_19556);
and U19997 (N_19997,N_19736,N_19636);
or U19998 (N_19998,N_19508,N_19572);
nand U19999 (N_19999,N_19709,N_19654);
nor U20000 (N_20000,N_19960,N_19806);
xnor U20001 (N_20001,N_19908,N_19757);
nand U20002 (N_20002,N_19918,N_19925);
xor U20003 (N_20003,N_19834,N_19914);
xnor U20004 (N_20004,N_19966,N_19752);
or U20005 (N_20005,N_19978,N_19758);
nand U20006 (N_20006,N_19921,N_19802);
or U20007 (N_20007,N_19778,N_19750);
nor U20008 (N_20008,N_19945,N_19933);
nor U20009 (N_20009,N_19905,N_19832);
or U20010 (N_20010,N_19965,N_19825);
nand U20011 (N_20011,N_19767,N_19899);
xnor U20012 (N_20012,N_19761,N_19873);
or U20013 (N_20013,N_19819,N_19789);
or U20014 (N_20014,N_19992,N_19958);
or U20015 (N_20015,N_19936,N_19829);
nand U20016 (N_20016,N_19956,N_19848);
nor U20017 (N_20017,N_19851,N_19976);
nand U20018 (N_20018,N_19830,N_19783);
xnor U20019 (N_20019,N_19787,N_19822);
nand U20020 (N_20020,N_19841,N_19967);
or U20021 (N_20021,N_19817,N_19809);
xnor U20022 (N_20022,N_19842,N_19970);
nand U20023 (N_20023,N_19891,N_19869);
or U20024 (N_20024,N_19799,N_19803);
or U20025 (N_20025,N_19926,N_19993);
xor U20026 (N_20026,N_19991,N_19881);
nor U20027 (N_20027,N_19919,N_19777);
and U20028 (N_20028,N_19975,N_19765);
or U20029 (N_20029,N_19900,N_19988);
xor U20030 (N_20030,N_19927,N_19795);
nor U20031 (N_20031,N_19963,N_19866);
xor U20032 (N_20032,N_19782,N_19964);
nor U20033 (N_20033,N_19801,N_19868);
nand U20034 (N_20034,N_19797,N_19931);
xnor U20035 (N_20035,N_19940,N_19860);
or U20036 (N_20036,N_19909,N_19784);
nor U20037 (N_20037,N_19995,N_19779);
or U20038 (N_20038,N_19864,N_19946);
or U20039 (N_20039,N_19838,N_19898);
nor U20040 (N_20040,N_19775,N_19769);
nand U20041 (N_20041,N_19754,N_19759);
or U20042 (N_20042,N_19911,N_19915);
xnor U20043 (N_20043,N_19969,N_19839);
nand U20044 (N_20044,N_19974,N_19895);
nor U20045 (N_20045,N_19878,N_19792);
nor U20046 (N_20046,N_19941,N_19780);
nand U20047 (N_20047,N_19984,N_19904);
xor U20048 (N_20048,N_19790,N_19875);
nor U20049 (N_20049,N_19948,N_19824);
or U20050 (N_20050,N_19858,N_19786);
and U20051 (N_20051,N_19916,N_19827);
or U20052 (N_20052,N_19844,N_19990);
xor U20053 (N_20053,N_19939,N_19770);
and U20054 (N_20054,N_19816,N_19937);
nand U20055 (N_20055,N_19962,N_19768);
nor U20056 (N_20056,N_19836,N_19961);
or U20057 (N_20057,N_19776,N_19846);
and U20058 (N_20058,N_19852,N_19883);
nand U20059 (N_20059,N_19996,N_19763);
and U20060 (N_20060,N_19913,N_19944);
or U20061 (N_20061,N_19879,N_19815);
nand U20062 (N_20062,N_19957,N_19863);
nand U20063 (N_20063,N_19753,N_19751);
xor U20064 (N_20064,N_19972,N_19896);
nor U20065 (N_20065,N_19855,N_19997);
and U20066 (N_20066,N_19843,N_19980);
and U20067 (N_20067,N_19821,N_19924);
nand U20068 (N_20068,N_19798,N_19986);
and U20069 (N_20069,N_19985,N_19870);
nor U20070 (N_20070,N_19894,N_19764);
xnor U20071 (N_20071,N_19889,N_19910);
nand U20072 (N_20072,N_19880,N_19794);
nand U20073 (N_20073,N_19892,N_19850);
xnor U20074 (N_20074,N_19952,N_19840);
nor U20075 (N_20075,N_19887,N_19968);
or U20076 (N_20076,N_19999,N_19877);
nor U20077 (N_20077,N_19781,N_19987);
or U20078 (N_20078,N_19932,N_19808);
nor U20079 (N_20079,N_19934,N_19772);
and U20080 (N_20080,N_19837,N_19849);
xnor U20081 (N_20081,N_19833,N_19818);
nand U20082 (N_20082,N_19862,N_19865);
xor U20083 (N_20083,N_19977,N_19943);
xnor U20084 (N_20084,N_19897,N_19828);
nor U20085 (N_20085,N_19859,N_19755);
nor U20086 (N_20086,N_19951,N_19930);
and U20087 (N_20087,N_19785,N_19981);
or U20088 (N_20088,N_19928,N_19774);
and U20089 (N_20089,N_19773,N_19857);
xnor U20090 (N_20090,N_19856,N_19831);
or U20091 (N_20091,N_19800,N_19923);
nand U20092 (N_20092,N_19810,N_19872);
xnor U20093 (N_20093,N_19853,N_19922);
or U20094 (N_20094,N_19998,N_19938);
nor U20095 (N_20095,N_19847,N_19813);
and U20096 (N_20096,N_19867,N_19906);
nor U20097 (N_20097,N_19955,N_19949);
and U20098 (N_20098,N_19812,N_19766);
or U20099 (N_20099,N_19912,N_19820);
nand U20100 (N_20100,N_19950,N_19788);
and U20101 (N_20101,N_19902,N_19762);
nor U20102 (N_20102,N_19882,N_19823);
nor U20103 (N_20103,N_19907,N_19884);
and U20104 (N_20104,N_19935,N_19982);
nor U20105 (N_20105,N_19953,N_19885);
nor U20106 (N_20106,N_19756,N_19903);
and U20107 (N_20107,N_19901,N_19888);
or U20108 (N_20108,N_19805,N_19973);
nor U20109 (N_20109,N_19959,N_19793);
nor U20110 (N_20110,N_19886,N_19791);
and U20111 (N_20111,N_19871,N_19971);
or U20112 (N_20112,N_19917,N_19942);
nor U20113 (N_20113,N_19771,N_19804);
xnor U20114 (N_20114,N_19994,N_19861);
nand U20115 (N_20115,N_19835,N_19826);
nor U20116 (N_20116,N_19920,N_19845);
nor U20117 (N_20117,N_19796,N_19814);
and U20118 (N_20118,N_19890,N_19979);
xor U20119 (N_20119,N_19876,N_19989);
xnor U20120 (N_20120,N_19929,N_19893);
or U20121 (N_20121,N_19760,N_19874);
and U20122 (N_20122,N_19954,N_19807);
xnor U20123 (N_20123,N_19854,N_19811);
nand U20124 (N_20124,N_19983,N_19947);
nor U20125 (N_20125,N_19992,N_19809);
nand U20126 (N_20126,N_19831,N_19982);
or U20127 (N_20127,N_19782,N_19812);
and U20128 (N_20128,N_19831,N_19848);
and U20129 (N_20129,N_19867,N_19769);
and U20130 (N_20130,N_19796,N_19977);
and U20131 (N_20131,N_19877,N_19783);
nor U20132 (N_20132,N_19933,N_19752);
nand U20133 (N_20133,N_19838,N_19773);
or U20134 (N_20134,N_19805,N_19965);
nand U20135 (N_20135,N_19971,N_19949);
xor U20136 (N_20136,N_19805,N_19855);
nor U20137 (N_20137,N_19769,N_19961);
xnor U20138 (N_20138,N_19943,N_19944);
and U20139 (N_20139,N_19873,N_19818);
and U20140 (N_20140,N_19814,N_19797);
xor U20141 (N_20141,N_19793,N_19788);
or U20142 (N_20142,N_19898,N_19867);
nand U20143 (N_20143,N_19756,N_19776);
and U20144 (N_20144,N_19751,N_19776);
and U20145 (N_20145,N_19859,N_19787);
nand U20146 (N_20146,N_19844,N_19940);
nor U20147 (N_20147,N_19961,N_19962);
and U20148 (N_20148,N_19964,N_19852);
xor U20149 (N_20149,N_19831,N_19834);
nand U20150 (N_20150,N_19923,N_19789);
or U20151 (N_20151,N_19863,N_19832);
xor U20152 (N_20152,N_19757,N_19827);
or U20153 (N_20153,N_19988,N_19875);
and U20154 (N_20154,N_19804,N_19958);
and U20155 (N_20155,N_19840,N_19856);
and U20156 (N_20156,N_19862,N_19897);
xor U20157 (N_20157,N_19820,N_19919);
or U20158 (N_20158,N_19828,N_19990);
and U20159 (N_20159,N_19917,N_19796);
nand U20160 (N_20160,N_19968,N_19776);
nand U20161 (N_20161,N_19898,N_19841);
nor U20162 (N_20162,N_19823,N_19890);
nor U20163 (N_20163,N_19941,N_19985);
or U20164 (N_20164,N_19763,N_19952);
nand U20165 (N_20165,N_19977,N_19923);
or U20166 (N_20166,N_19953,N_19987);
or U20167 (N_20167,N_19966,N_19758);
nand U20168 (N_20168,N_19942,N_19757);
and U20169 (N_20169,N_19973,N_19992);
and U20170 (N_20170,N_19845,N_19835);
nor U20171 (N_20171,N_19990,N_19854);
or U20172 (N_20172,N_19784,N_19832);
nor U20173 (N_20173,N_19944,N_19761);
or U20174 (N_20174,N_19792,N_19805);
xnor U20175 (N_20175,N_19763,N_19979);
nor U20176 (N_20176,N_19790,N_19908);
and U20177 (N_20177,N_19807,N_19960);
xor U20178 (N_20178,N_19862,N_19845);
or U20179 (N_20179,N_19835,N_19919);
or U20180 (N_20180,N_19940,N_19998);
and U20181 (N_20181,N_19834,N_19954);
nand U20182 (N_20182,N_19979,N_19986);
nand U20183 (N_20183,N_19988,N_19937);
or U20184 (N_20184,N_19861,N_19757);
and U20185 (N_20185,N_19810,N_19835);
or U20186 (N_20186,N_19817,N_19890);
nor U20187 (N_20187,N_19982,N_19854);
or U20188 (N_20188,N_19787,N_19926);
or U20189 (N_20189,N_19775,N_19759);
and U20190 (N_20190,N_19769,N_19796);
nor U20191 (N_20191,N_19992,N_19825);
nor U20192 (N_20192,N_19845,N_19876);
and U20193 (N_20193,N_19949,N_19850);
or U20194 (N_20194,N_19770,N_19809);
nand U20195 (N_20195,N_19884,N_19920);
xor U20196 (N_20196,N_19875,N_19912);
or U20197 (N_20197,N_19847,N_19868);
nand U20198 (N_20198,N_19891,N_19877);
nor U20199 (N_20199,N_19764,N_19879);
or U20200 (N_20200,N_19803,N_19764);
and U20201 (N_20201,N_19849,N_19803);
xor U20202 (N_20202,N_19952,N_19793);
xor U20203 (N_20203,N_19770,N_19814);
xnor U20204 (N_20204,N_19895,N_19852);
and U20205 (N_20205,N_19832,N_19785);
xor U20206 (N_20206,N_19799,N_19762);
and U20207 (N_20207,N_19848,N_19910);
xor U20208 (N_20208,N_19916,N_19754);
nand U20209 (N_20209,N_19854,N_19885);
xor U20210 (N_20210,N_19782,N_19923);
nor U20211 (N_20211,N_19938,N_19780);
or U20212 (N_20212,N_19776,N_19870);
or U20213 (N_20213,N_19800,N_19827);
nand U20214 (N_20214,N_19911,N_19851);
nor U20215 (N_20215,N_19922,N_19844);
xnor U20216 (N_20216,N_19771,N_19883);
xor U20217 (N_20217,N_19818,N_19920);
nor U20218 (N_20218,N_19894,N_19874);
nand U20219 (N_20219,N_19839,N_19876);
nand U20220 (N_20220,N_19814,N_19847);
xnor U20221 (N_20221,N_19907,N_19777);
and U20222 (N_20222,N_19768,N_19796);
xor U20223 (N_20223,N_19839,N_19836);
nor U20224 (N_20224,N_19988,N_19884);
or U20225 (N_20225,N_19982,N_19971);
nor U20226 (N_20226,N_19937,N_19817);
or U20227 (N_20227,N_19952,N_19767);
nand U20228 (N_20228,N_19958,N_19846);
nand U20229 (N_20229,N_19886,N_19865);
xnor U20230 (N_20230,N_19816,N_19857);
xor U20231 (N_20231,N_19947,N_19999);
and U20232 (N_20232,N_19878,N_19795);
or U20233 (N_20233,N_19945,N_19867);
xor U20234 (N_20234,N_19999,N_19940);
xnor U20235 (N_20235,N_19959,N_19772);
and U20236 (N_20236,N_19876,N_19963);
or U20237 (N_20237,N_19852,N_19761);
or U20238 (N_20238,N_19922,N_19936);
and U20239 (N_20239,N_19962,N_19906);
xor U20240 (N_20240,N_19867,N_19927);
xnor U20241 (N_20241,N_19876,N_19762);
xnor U20242 (N_20242,N_19760,N_19753);
or U20243 (N_20243,N_19840,N_19805);
nand U20244 (N_20244,N_19969,N_19850);
nor U20245 (N_20245,N_19948,N_19908);
and U20246 (N_20246,N_19753,N_19818);
nor U20247 (N_20247,N_19952,N_19969);
nor U20248 (N_20248,N_19855,N_19841);
and U20249 (N_20249,N_19867,N_19932);
nand U20250 (N_20250,N_20136,N_20085);
or U20251 (N_20251,N_20197,N_20209);
or U20252 (N_20252,N_20236,N_20006);
or U20253 (N_20253,N_20180,N_20070);
and U20254 (N_20254,N_20018,N_20160);
nor U20255 (N_20255,N_20123,N_20010);
nor U20256 (N_20256,N_20244,N_20154);
nor U20257 (N_20257,N_20113,N_20235);
xor U20258 (N_20258,N_20106,N_20164);
xnor U20259 (N_20259,N_20028,N_20091);
xnor U20260 (N_20260,N_20174,N_20147);
xor U20261 (N_20261,N_20133,N_20097);
nor U20262 (N_20262,N_20151,N_20105);
and U20263 (N_20263,N_20152,N_20109);
nand U20264 (N_20264,N_20040,N_20053);
nor U20265 (N_20265,N_20043,N_20014);
or U20266 (N_20266,N_20212,N_20068);
and U20267 (N_20267,N_20139,N_20168);
or U20268 (N_20268,N_20107,N_20046);
and U20269 (N_20269,N_20193,N_20083);
xnor U20270 (N_20270,N_20054,N_20167);
and U20271 (N_20271,N_20146,N_20149);
nand U20272 (N_20272,N_20076,N_20022);
nor U20273 (N_20273,N_20215,N_20041);
and U20274 (N_20274,N_20242,N_20108);
nand U20275 (N_20275,N_20089,N_20143);
or U20276 (N_20276,N_20065,N_20048);
or U20277 (N_20277,N_20189,N_20037);
xor U20278 (N_20278,N_20208,N_20185);
nor U20279 (N_20279,N_20052,N_20213);
or U20280 (N_20280,N_20203,N_20030);
nor U20281 (N_20281,N_20207,N_20119);
nand U20282 (N_20282,N_20093,N_20163);
nor U20283 (N_20283,N_20016,N_20138);
nand U20284 (N_20284,N_20231,N_20178);
xor U20285 (N_20285,N_20225,N_20239);
nor U20286 (N_20286,N_20223,N_20015);
xnor U20287 (N_20287,N_20087,N_20232);
and U20288 (N_20288,N_20102,N_20222);
and U20289 (N_20289,N_20063,N_20004);
nor U20290 (N_20290,N_20027,N_20058);
xnor U20291 (N_20291,N_20241,N_20033);
nand U20292 (N_20292,N_20003,N_20009);
and U20293 (N_20293,N_20243,N_20135);
xnor U20294 (N_20294,N_20158,N_20162);
nor U20295 (N_20295,N_20122,N_20165);
nand U20296 (N_20296,N_20013,N_20072);
nor U20297 (N_20297,N_20100,N_20038);
and U20298 (N_20298,N_20196,N_20140);
xor U20299 (N_20299,N_20219,N_20086);
nand U20300 (N_20300,N_20184,N_20098);
xnor U20301 (N_20301,N_20214,N_20061);
nand U20302 (N_20302,N_20036,N_20005);
or U20303 (N_20303,N_20127,N_20169);
nand U20304 (N_20304,N_20118,N_20011);
nor U20305 (N_20305,N_20090,N_20077);
nand U20306 (N_20306,N_20177,N_20148);
nor U20307 (N_20307,N_20240,N_20246);
nand U20308 (N_20308,N_20078,N_20092);
and U20309 (N_20309,N_20039,N_20190);
nand U20310 (N_20310,N_20029,N_20195);
nand U20311 (N_20311,N_20103,N_20071);
xnor U20312 (N_20312,N_20198,N_20044);
nor U20313 (N_20313,N_20073,N_20220);
nand U20314 (N_20314,N_20024,N_20238);
xor U20315 (N_20315,N_20096,N_20159);
or U20316 (N_20316,N_20045,N_20128);
or U20317 (N_20317,N_20157,N_20179);
or U20318 (N_20318,N_20171,N_20114);
nor U20319 (N_20319,N_20248,N_20069);
xor U20320 (N_20320,N_20021,N_20226);
nor U20321 (N_20321,N_20124,N_20218);
or U20322 (N_20322,N_20192,N_20064);
nand U20323 (N_20323,N_20001,N_20175);
nor U20324 (N_20324,N_20141,N_20111);
nor U20325 (N_20325,N_20026,N_20012);
and U20326 (N_20326,N_20230,N_20047);
xor U20327 (N_20327,N_20104,N_20211);
nand U20328 (N_20328,N_20199,N_20080);
and U20329 (N_20329,N_20183,N_20188);
xnor U20330 (N_20330,N_20237,N_20145);
and U20331 (N_20331,N_20150,N_20182);
and U20332 (N_20332,N_20131,N_20137);
nor U20333 (N_20333,N_20216,N_20217);
or U20334 (N_20334,N_20019,N_20191);
nand U20335 (N_20335,N_20249,N_20049);
nand U20336 (N_20336,N_20181,N_20229);
xnor U20337 (N_20337,N_20125,N_20062);
and U20338 (N_20338,N_20117,N_20099);
or U20339 (N_20339,N_20210,N_20057);
and U20340 (N_20340,N_20134,N_20166);
and U20341 (N_20341,N_20074,N_20234);
nor U20342 (N_20342,N_20101,N_20088);
and U20343 (N_20343,N_20035,N_20082);
xor U20344 (N_20344,N_20227,N_20032);
nand U20345 (N_20345,N_20200,N_20233);
and U20346 (N_20346,N_20247,N_20156);
nand U20347 (N_20347,N_20034,N_20017);
nor U20348 (N_20348,N_20060,N_20031);
nand U20349 (N_20349,N_20161,N_20186);
nand U20350 (N_20350,N_20067,N_20120);
xor U20351 (N_20351,N_20204,N_20050);
nor U20352 (N_20352,N_20023,N_20202);
or U20353 (N_20353,N_20205,N_20025);
and U20354 (N_20354,N_20116,N_20075);
or U20355 (N_20355,N_20042,N_20126);
xor U20356 (N_20356,N_20176,N_20084);
nor U20357 (N_20357,N_20142,N_20129);
or U20358 (N_20358,N_20115,N_20094);
nand U20359 (N_20359,N_20055,N_20173);
and U20360 (N_20360,N_20020,N_20007);
and U20361 (N_20361,N_20221,N_20206);
nand U20362 (N_20362,N_20081,N_20112);
nor U20363 (N_20363,N_20000,N_20132);
and U20364 (N_20364,N_20008,N_20245);
or U20365 (N_20365,N_20172,N_20153);
or U20366 (N_20366,N_20170,N_20201);
xor U20367 (N_20367,N_20110,N_20144);
or U20368 (N_20368,N_20194,N_20121);
nand U20369 (N_20369,N_20079,N_20155);
nor U20370 (N_20370,N_20066,N_20002);
and U20371 (N_20371,N_20130,N_20059);
and U20372 (N_20372,N_20095,N_20056);
nor U20373 (N_20373,N_20051,N_20224);
or U20374 (N_20374,N_20187,N_20228);
or U20375 (N_20375,N_20030,N_20193);
nor U20376 (N_20376,N_20179,N_20051);
or U20377 (N_20377,N_20197,N_20091);
nand U20378 (N_20378,N_20149,N_20016);
nand U20379 (N_20379,N_20168,N_20146);
nor U20380 (N_20380,N_20025,N_20133);
and U20381 (N_20381,N_20067,N_20156);
xnor U20382 (N_20382,N_20189,N_20041);
nand U20383 (N_20383,N_20045,N_20025);
xnor U20384 (N_20384,N_20203,N_20080);
nand U20385 (N_20385,N_20165,N_20098);
and U20386 (N_20386,N_20182,N_20001);
and U20387 (N_20387,N_20207,N_20020);
nor U20388 (N_20388,N_20069,N_20223);
and U20389 (N_20389,N_20021,N_20078);
and U20390 (N_20390,N_20168,N_20138);
nor U20391 (N_20391,N_20001,N_20223);
and U20392 (N_20392,N_20110,N_20145);
and U20393 (N_20393,N_20194,N_20159);
and U20394 (N_20394,N_20031,N_20175);
nor U20395 (N_20395,N_20238,N_20005);
xor U20396 (N_20396,N_20117,N_20229);
nand U20397 (N_20397,N_20080,N_20161);
or U20398 (N_20398,N_20242,N_20072);
nor U20399 (N_20399,N_20032,N_20246);
nor U20400 (N_20400,N_20181,N_20129);
nor U20401 (N_20401,N_20204,N_20201);
nor U20402 (N_20402,N_20106,N_20073);
or U20403 (N_20403,N_20133,N_20155);
and U20404 (N_20404,N_20130,N_20191);
nand U20405 (N_20405,N_20175,N_20199);
and U20406 (N_20406,N_20060,N_20175);
nand U20407 (N_20407,N_20004,N_20118);
or U20408 (N_20408,N_20016,N_20094);
or U20409 (N_20409,N_20086,N_20141);
xnor U20410 (N_20410,N_20139,N_20245);
and U20411 (N_20411,N_20207,N_20018);
nor U20412 (N_20412,N_20059,N_20172);
nor U20413 (N_20413,N_20245,N_20073);
or U20414 (N_20414,N_20199,N_20097);
nand U20415 (N_20415,N_20084,N_20019);
or U20416 (N_20416,N_20171,N_20238);
or U20417 (N_20417,N_20136,N_20235);
nor U20418 (N_20418,N_20189,N_20187);
nand U20419 (N_20419,N_20040,N_20042);
nand U20420 (N_20420,N_20077,N_20006);
and U20421 (N_20421,N_20099,N_20007);
xnor U20422 (N_20422,N_20132,N_20100);
nand U20423 (N_20423,N_20128,N_20050);
xor U20424 (N_20424,N_20063,N_20244);
and U20425 (N_20425,N_20147,N_20142);
xnor U20426 (N_20426,N_20103,N_20217);
or U20427 (N_20427,N_20097,N_20094);
or U20428 (N_20428,N_20014,N_20217);
or U20429 (N_20429,N_20008,N_20213);
xor U20430 (N_20430,N_20199,N_20044);
or U20431 (N_20431,N_20101,N_20164);
and U20432 (N_20432,N_20029,N_20142);
xor U20433 (N_20433,N_20217,N_20051);
nor U20434 (N_20434,N_20041,N_20031);
nand U20435 (N_20435,N_20225,N_20124);
nor U20436 (N_20436,N_20019,N_20034);
xor U20437 (N_20437,N_20128,N_20241);
xor U20438 (N_20438,N_20036,N_20172);
and U20439 (N_20439,N_20114,N_20055);
or U20440 (N_20440,N_20173,N_20062);
and U20441 (N_20441,N_20193,N_20012);
nand U20442 (N_20442,N_20066,N_20020);
or U20443 (N_20443,N_20167,N_20056);
or U20444 (N_20444,N_20025,N_20208);
nand U20445 (N_20445,N_20196,N_20127);
nand U20446 (N_20446,N_20216,N_20018);
and U20447 (N_20447,N_20152,N_20132);
nor U20448 (N_20448,N_20204,N_20011);
and U20449 (N_20449,N_20026,N_20179);
or U20450 (N_20450,N_20030,N_20047);
and U20451 (N_20451,N_20133,N_20040);
nand U20452 (N_20452,N_20205,N_20155);
nand U20453 (N_20453,N_20099,N_20146);
xnor U20454 (N_20454,N_20121,N_20075);
nor U20455 (N_20455,N_20179,N_20223);
nand U20456 (N_20456,N_20225,N_20090);
and U20457 (N_20457,N_20077,N_20062);
nand U20458 (N_20458,N_20023,N_20118);
or U20459 (N_20459,N_20222,N_20130);
and U20460 (N_20460,N_20231,N_20053);
nor U20461 (N_20461,N_20126,N_20131);
nand U20462 (N_20462,N_20108,N_20243);
or U20463 (N_20463,N_20094,N_20177);
nand U20464 (N_20464,N_20076,N_20189);
nor U20465 (N_20465,N_20109,N_20083);
nor U20466 (N_20466,N_20078,N_20107);
or U20467 (N_20467,N_20006,N_20137);
xnor U20468 (N_20468,N_20054,N_20140);
or U20469 (N_20469,N_20012,N_20137);
xnor U20470 (N_20470,N_20058,N_20137);
or U20471 (N_20471,N_20244,N_20043);
nand U20472 (N_20472,N_20046,N_20161);
or U20473 (N_20473,N_20186,N_20120);
xor U20474 (N_20474,N_20219,N_20105);
nand U20475 (N_20475,N_20166,N_20236);
or U20476 (N_20476,N_20084,N_20104);
xnor U20477 (N_20477,N_20219,N_20123);
nor U20478 (N_20478,N_20161,N_20072);
and U20479 (N_20479,N_20016,N_20106);
nand U20480 (N_20480,N_20155,N_20224);
and U20481 (N_20481,N_20047,N_20036);
xor U20482 (N_20482,N_20090,N_20118);
nor U20483 (N_20483,N_20051,N_20091);
and U20484 (N_20484,N_20096,N_20129);
xnor U20485 (N_20485,N_20185,N_20075);
and U20486 (N_20486,N_20158,N_20085);
nand U20487 (N_20487,N_20211,N_20169);
or U20488 (N_20488,N_20189,N_20043);
nor U20489 (N_20489,N_20083,N_20020);
and U20490 (N_20490,N_20175,N_20160);
nand U20491 (N_20491,N_20091,N_20110);
nor U20492 (N_20492,N_20205,N_20204);
xnor U20493 (N_20493,N_20017,N_20197);
nand U20494 (N_20494,N_20224,N_20181);
and U20495 (N_20495,N_20196,N_20054);
and U20496 (N_20496,N_20049,N_20089);
nand U20497 (N_20497,N_20001,N_20004);
and U20498 (N_20498,N_20021,N_20120);
xor U20499 (N_20499,N_20051,N_20146);
nand U20500 (N_20500,N_20381,N_20386);
or U20501 (N_20501,N_20430,N_20498);
nand U20502 (N_20502,N_20264,N_20288);
nor U20503 (N_20503,N_20298,N_20431);
nand U20504 (N_20504,N_20377,N_20297);
xor U20505 (N_20505,N_20362,N_20432);
or U20506 (N_20506,N_20373,N_20353);
or U20507 (N_20507,N_20342,N_20406);
xor U20508 (N_20508,N_20496,N_20396);
or U20509 (N_20509,N_20411,N_20367);
nor U20510 (N_20510,N_20408,N_20299);
nor U20511 (N_20511,N_20444,N_20291);
or U20512 (N_20512,N_20348,N_20319);
xnor U20513 (N_20513,N_20472,N_20439);
nor U20514 (N_20514,N_20344,N_20347);
and U20515 (N_20515,N_20417,N_20470);
or U20516 (N_20516,N_20437,N_20427);
nor U20517 (N_20517,N_20383,N_20301);
nor U20518 (N_20518,N_20407,N_20255);
and U20519 (N_20519,N_20363,N_20358);
and U20520 (N_20520,N_20372,N_20335);
xor U20521 (N_20521,N_20464,N_20390);
xor U20522 (N_20522,N_20399,N_20425);
xor U20523 (N_20523,N_20487,N_20334);
or U20524 (N_20524,N_20316,N_20389);
or U20525 (N_20525,N_20279,N_20269);
and U20526 (N_20526,N_20493,N_20458);
nand U20527 (N_20527,N_20262,N_20424);
or U20528 (N_20528,N_20480,N_20414);
or U20529 (N_20529,N_20375,N_20440);
nand U20530 (N_20530,N_20361,N_20481);
nand U20531 (N_20531,N_20345,N_20258);
nor U20532 (N_20532,N_20459,N_20446);
xor U20533 (N_20533,N_20488,N_20415);
xnor U20534 (N_20534,N_20388,N_20395);
or U20535 (N_20535,N_20420,N_20397);
nand U20536 (N_20536,N_20465,N_20378);
or U20537 (N_20537,N_20486,N_20426);
and U20538 (N_20538,N_20272,N_20312);
xnor U20539 (N_20539,N_20280,N_20351);
xnor U20540 (N_20540,N_20306,N_20254);
and U20541 (N_20541,N_20268,N_20302);
nor U20542 (N_20542,N_20359,N_20366);
and U20543 (N_20543,N_20490,N_20273);
nor U20544 (N_20544,N_20275,N_20284);
or U20545 (N_20545,N_20250,N_20277);
nand U20546 (N_20546,N_20402,N_20318);
or U20547 (N_20547,N_20341,N_20438);
or U20548 (N_20548,N_20423,N_20382);
nand U20549 (N_20549,N_20323,N_20283);
xnor U20550 (N_20550,N_20349,N_20332);
nand U20551 (N_20551,N_20292,N_20466);
nor U20552 (N_20552,N_20336,N_20267);
nor U20553 (N_20553,N_20266,N_20448);
xor U20554 (N_20554,N_20281,N_20436);
nand U20555 (N_20555,N_20494,N_20460);
or U20556 (N_20556,N_20355,N_20482);
xnor U20557 (N_20557,N_20419,N_20270);
and U20558 (N_20558,N_20308,N_20320);
nor U20559 (N_20559,N_20314,N_20433);
nand U20560 (N_20560,N_20252,N_20285);
and U20561 (N_20561,N_20309,N_20315);
or U20562 (N_20562,N_20326,N_20416);
xor U20563 (N_20563,N_20369,N_20385);
nand U20564 (N_20564,N_20303,N_20339);
and U20565 (N_20565,N_20449,N_20313);
and U20566 (N_20566,N_20421,N_20329);
or U20567 (N_20567,N_20499,N_20327);
nor U20568 (N_20568,N_20379,N_20462);
and U20569 (N_20569,N_20317,N_20461);
or U20570 (N_20570,N_20380,N_20253);
nor U20571 (N_20571,N_20333,N_20370);
or U20572 (N_20572,N_20305,N_20338);
xnor U20573 (N_20573,N_20453,N_20259);
xnor U20574 (N_20574,N_20322,N_20392);
nand U20575 (N_20575,N_20463,N_20265);
nor U20576 (N_20576,N_20489,N_20276);
or U20577 (N_20577,N_20256,N_20394);
and U20578 (N_20578,N_20450,N_20357);
and U20579 (N_20579,N_20293,N_20492);
nand U20580 (N_20580,N_20340,N_20483);
or U20581 (N_20581,N_20374,N_20434);
and U20582 (N_20582,N_20451,N_20321);
or U20583 (N_20583,N_20473,N_20296);
or U20584 (N_20584,N_20413,N_20401);
and U20585 (N_20585,N_20405,N_20376);
nor U20586 (N_20586,N_20457,N_20330);
xnor U20587 (N_20587,N_20477,N_20310);
xnor U20588 (N_20588,N_20365,N_20410);
nand U20589 (N_20589,N_20422,N_20469);
nand U20590 (N_20590,N_20282,N_20455);
and U20591 (N_20591,N_20307,N_20398);
xor U20592 (N_20592,N_20350,N_20356);
nor U20593 (N_20593,N_20328,N_20287);
xnor U20594 (N_20594,N_20471,N_20474);
xor U20595 (N_20595,N_20409,N_20484);
xor U20596 (N_20596,N_20403,N_20478);
xnor U20597 (N_20597,N_20294,N_20441);
or U20598 (N_20598,N_20452,N_20304);
and U20599 (N_20599,N_20443,N_20368);
xnor U20600 (N_20600,N_20447,N_20346);
and U20601 (N_20601,N_20271,N_20337);
or U20602 (N_20602,N_20311,N_20442);
nor U20603 (N_20603,N_20454,N_20393);
xor U20604 (N_20604,N_20468,N_20290);
nor U20605 (N_20605,N_20467,N_20387);
xor U20606 (N_20606,N_20435,N_20400);
nand U20607 (N_20607,N_20445,N_20497);
or U20608 (N_20608,N_20260,N_20371);
xnor U20609 (N_20609,N_20456,N_20325);
and U20610 (N_20610,N_20391,N_20261);
nand U20611 (N_20611,N_20412,N_20485);
or U20612 (N_20612,N_20263,N_20352);
nor U20613 (N_20613,N_20479,N_20495);
or U20614 (N_20614,N_20295,N_20429);
nand U20615 (N_20615,N_20331,N_20343);
xnor U20616 (N_20616,N_20476,N_20324);
xnor U20617 (N_20617,N_20428,N_20289);
nor U20618 (N_20618,N_20354,N_20491);
nand U20619 (N_20619,N_20300,N_20278);
xor U20620 (N_20620,N_20404,N_20418);
nand U20621 (N_20621,N_20475,N_20364);
and U20622 (N_20622,N_20257,N_20360);
xor U20623 (N_20623,N_20274,N_20384);
nand U20624 (N_20624,N_20286,N_20251);
nor U20625 (N_20625,N_20309,N_20447);
xnor U20626 (N_20626,N_20339,N_20325);
nand U20627 (N_20627,N_20294,N_20448);
xor U20628 (N_20628,N_20423,N_20486);
or U20629 (N_20629,N_20259,N_20335);
xnor U20630 (N_20630,N_20484,N_20378);
xnor U20631 (N_20631,N_20490,N_20396);
nor U20632 (N_20632,N_20416,N_20271);
or U20633 (N_20633,N_20479,N_20417);
nor U20634 (N_20634,N_20256,N_20337);
xnor U20635 (N_20635,N_20435,N_20449);
nand U20636 (N_20636,N_20384,N_20385);
and U20637 (N_20637,N_20384,N_20285);
and U20638 (N_20638,N_20365,N_20361);
or U20639 (N_20639,N_20322,N_20365);
xnor U20640 (N_20640,N_20484,N_20316);
and U20641 (N_20641,N_20337,N_20354);
nor U20642 (N_20642,N_20322,N_20440);
and U20643 (N_20643,N_20478,N_20282);
and U20644 (N_20644,N_20251,N_20331);
or U20645 (N_20645,N_20399,N_20364);
and U20646 (N_20646,N_20495,N_20323);
xor U20647 (N_20647,N_20345,N_20294);
and U20648 (N_20648,N_20422,N_20307);
or U20649 (N_20649,N_20255,N_20431);
and U20650 (N_20650,N_20464,N_20457);
nor U20651 (N_20651,N_20414,N_20289);
and U20652 (N_20652,N_20369,N_20459);
nand U20653 (N_20653,N_20465,N_20358);
nand U20654 (N_20654,N_20424,N_20329);
nor U20655 (N_20655,N_20298,N_20392);
nand U20656 (N_20656,N_20314,N_20251);
nor U20657 (N_20657,N_20418,N_20449);
or U20658 (N_20658,N_20491,N_20308);
nor U20659 (N_20659,N_20256,N_20347);
nand U20660 (N_20660,N_20430,N_20463);
or U20661 (N_20661,N_20449,N_20476);
nand U20662 (N_20662,N_20309,N_20401);
and U20663 (N_20663,N_20483,N_20409);
and U20664 (N_20664,N_20298,N_20440);
xor U20665 (N_20665,N_20369,N_20357);
nor U20666 (N_20666,N_20258,N_20375);
or U20667 (N_20667,N_20353,N_20319);
nand U20668 (N_20668,N_20304,N_20346);
nor U20669 (N_20669,N_20454,N_20308);
and U20670 (N_20670,N_20276,N_20373);
nor U20671 (N_20671,N_20497,N_20488);
or U20672 (N_20672,N_20411,N_20451);
and U20673 (N_20673,N_20394,N_20488);
or U20674 (N_20674,N_20410,N_20266);
xnor U20675 (N_20675,N_20392,N_20393);
or U20676 (N_20676,N_20467,N_20493);
nand U20677 (N_20677,N_20455,N_20444);
or U20678 (N_20678,N_20330,N_20498);
or U20679 (N_20679,N_20296,N_20448);
or U20680 (N_20680,N_20469,N_20257);
nand U20681 (N_20681,N_20261,N_20468);
and U20682 (N_20682,N_20360,N_20262);
or U20683 (N_20683,N_20421,N_20294);
nor U20684 (N_20684,N_20469,N_20309);
nor U20685 (N_20685,N_20468,N_20399);
nand U20686 (N_20686,N_20382,N_20436);
nor U20687 (N_20687,N_20446,N_20444);
and U20688 (N_20688,N_20331,N_20313);
or U20689 (N_20689,N_20281,N_20465);
or U20690 (N_20690,N_20427,N_20291);
and U20691 (N_20691,N_20477,N_20442);
nor U20692 (N_20692,N_20469,N_20275);
and U20693 (N_20693,N_20327,N_20395);
or U20694 (N_20694,N_20397,N_20490);
nand U20695 (N_20695,N_20352,N_20441);
and U20696 (N_20696,N_20475,N_20380);
or U20697 (N_20697,N_20429,N_20494);
xor U20698 (N_20698,N_20315,N_20489);
and U20699 (N_20699,N_20329,N_20406);
nand U20700 (N_20700,N_20412,N_20328);
nand U20701 (N_20701,N_20283,N_20465);
and U20702 (N_20702,N_20327,N_20468);
xnor U20703 (N_20703,N_20359,N_20302);
or U20704 (N_20704,N_20290,N_20465);
xor U20705 (N_20705,N_20493,N_20459);
or U20706 (N_20706,N_20370,N_20319);
and U20707 (N_20707,N_20472,N_20416);
or U20708 (N_20708,N_20293,N_20353);
and U20709 (N_20709,N_20441,N_20433);
nand U20710 (N_20710,N_20256,N_20290);
and U20711 (N_20711,N_20485,N_20382);
xnor U20712 (N_20712,N_20335,N_20471);
or U20713 (N_20713,N_20341,N_20453);
nor U20714 (N_20714,N_20399,N_20469);
and U20715 (N_20715,N_20464,N_20331);
or U20716 (N_20716,N_20257,N_20340);
or U20717 (N_20717,N_20337,N_20378);
xor U20718 (N_20718,N_20295,N_20445);
xor U20719 (N_20719,N_20307,N_20288);
and U20720 (N_20720,N_20254,N_20485);
nand U20721 (N_20721,N_20424,N_20451);
nand U20722 (N_20722,N_20346,N_20422);
nor U20723 (N_20723,N_20318,N_20321);
and U20724 (N_20724,N_20412,N_20421);
nand U20725 (N_20725,N_20284,N_20460);
and U20726 (N_20726,N_20335,N_20377);
or U20727 (N_20727,N_20374,N_20305);
nand U20728 (N_20728,N_20413,N_20480);
xor U20729 (N_20729,N_20317,N_20260);
and U20730 (N_20730,N_20309,N_20350);
xnor U20731 (N_20731,N_20442,N_20267);
and U20732 (N_20732,N_20402,N_20436);
or U20733 (N_20733,N_20343,N_20385);
or U20734 (N_20734,N_20408,N_20478);
and U20735 (N_20735,N_20310,N_20464);
nand U20736 (N_20736,N_20448,N_20356);
nor U20737 (N_20737,N_20420,N_20419);
nand U20738 (N_20738,N_20321,N_20442);
or U20739 (N_20739,N_20252,N_20310);
or U20740 (N_20740,N_20434,N_20410);
nand U20741 (N_20741,N_20323,N_20315);
or U20742 (N_20742,N_20384,N_20391);
and U20743 (N_20743,N_20452,N_20444);
xor U20744 (N_20744,N_20349,N_20467);
nand U20745 (N_20745,N_20361,N_20492);
or U20746 (N_20746,N_20386,N_20435);
and U20747 (N_20747,N_20319,N_20265);
or U20748 (N_20748,N_20260,N_20424);
or U20749 (N_20749,N_20398,N_20335);
and U20750 (N_20750,N_20519,N_20682);
nor U20751 (N_20751,N_20705,N_20692);
nand U20752 (N_20752,N_20616,N_20595);
and U20753 (N_20753,N_20685,N_20748);
xnor U20754 (N_20754,N_20668,N_20719);
or U20755 (N_20755,N_20712,N_20627);
or U20756 (N_20756,N_20565,N_20707);
nor U20757 (N_20757,N_20612,N_20671);
nand U20758 (N_20758,N_20728,N_20659);
xor U20759 (N_20759,N_20663,N_20655);
or U20760 (N_20760,N_20572,N_20722);
xor U20761 (N_20761,N_20573,N_20622);
and U20762 (N_20762,N_20589,N_20564);
or U20763 (N_20763,N_20513,N_20724);
xor U20764 (N_20764,N_20533,N_20648);
or U20765 (N_20765,N_20696,N_20702);
xor U20766 (N_20766,N_20545,N_20703);
or U20767 (N_20767,N_20599,N_20646);
nand U20768 (N_20768,N_20694,N_20738);
nor U20769 (N_20769,N_20571,N_20615);
and U20770 (N_20770,N_20523,N_20597);
nor U20771 (N_20771,N_20548,N_20536);
nand U20772 (N_20772,N_20594,N_20733);
xor U20773 (N_20773,N_20527,N_20674);
or U20774 (N_20774,N_20617,N_20735);
nand U20775 (N_20775,N_20718,N_20747);
nand U20776 (N_20776,N_20690,N_20505);
nor U20777 (N_20777,N_20587,N_20596);
and U20778 (N_20778,N_20567,N_20683);
or U20779 (N_20779,N_20525,N_20512);
xor U20780 (N_20780,N_20639,N_20563);
and U20781 (N_20781,N_20670,N_20501);
nand U20782 (N_20782,N_20637,N_20516);
or U20783 (N_20783,N_20720,N_20591);
xnor U20784 (N_20784,N_20559,N_20518);
and U20785 (N_20785,N_20592,N_20636);
and U20786 (N_20786,N_20699,N_20607);
nand U20787 (N_20787,N_20675,N_20613);
xor U20788 (N_20788,N_20678,N_20649);
nand U20789 (N_20789,N_20598,N_20638);
and U20790 (N_20790,N_20582,N_20725);
or U20791 (N_20791,N_20601,N_20538);
or U20792 (N_20792,N_20658,N_20584);
xnor U20793 (N_20793,N_20715,N_20546);
nor U20794 (N_20794,N_20691,N_20697);
nand U20795 (N_20795,N_20727,N_20709);
nor U20796 (N_20796,N_20628,N_20681);
or U20797 (N_20797,N_20515,N_20631);
nand U20798 (N_20798,N_20633,N_20575);
xor U20799 (N_20799,N_20570,N_20689);
or U20800 (N_20800,N_20614,N_20608);
xor U20801 (N_20801,N_20520,N_20641);
or U20802 (N_20802,N_20600,N_20632);
nand U20803 (N_20803,N_20581,N_20540);
nor U20804 (N_20804,N_20530,N_20602);
and U20805 (N_20805,N_20517,N_20693);
nand U20806 (N_20806,N_20643,N_20716);
xor U20807 (N_20807,N_20506,N_20619);
and U20808 (N_20808,N_20524,N_20574);
and U20809 (N_20809,N_20521,N_20746);
or U20810 (N_20810,N_20710,N_20629);
and U20811 (N_20811,N_20635,N_20680);
nor U20812 (N_20812,N_20620,N_20731);
nor U20813 (N_20813,N_20665,N_20726);
nand U20814 (N_20814,N_20560,N_20729);
or U20815 (N_20815,N_20645,N_20593);
and U20816 (N_20816,N_20528,N_20660);
nor U20817 (N_20817,N_20568,N_20514);
or U20818 (N_20818,N_20507,N_20654);
nand U20819 (N_20819,N_20737,N_20531);
and U20820 (N_20820,N_20606,N_20745);
or U20821 (N_20821,N_20618,N_20555);
or U20822 (N_20822,N_20554,N_20586);
nand U20823 (N_20823,N_20704,N_20624);
xor U20824 (N_20824,N_20698,N_20566);
nand U20825 (N_20825,N_20740,N_20686);
and U20826 (N_20826,N_20701,N_20662);
or U20827 (N_20827,N_20642,N_20541);
nand U20828 (N_20828,N_20644,N_20544);
xnor U20829 (N_20829,N_20552,N_20534);
nor U20830 (N_20830,N_20569,N_20713);
nor U20831 (N_20831,N_20736,N_20529);
and U20832 (N_20832,N_20577,N_20688);
or U20833 (N_20833,N_20551,N_20500);
or U20834 (N_20834,N_20610,N_20717);
or U20835 (N_20835,N_20621,N_20630);
or U20836 (N_20836,N_20650,N_20547);
and U20837 (N_20837,N_20611,N_20749);
and U20838 (N_20838,N_20604,N_20549);
and U20839 (N_20839,N_20667,N_20640);
xor U20840 (N_20840,N_20556,N_20539);
nor U20841 (N_20841,N_20625,N_20730);
or U20842 (N_20842,N_20684,N_20510);
xor U20843 (N_20843,N_20664,N_20504);
nor U20844 (N_20844,N_20669,N_20732);
xnor U20845 (N_20845,N_20700,N_20741);
and U20846 (N_20846,N_20522,N_20734);
and U20847 (N_20847,N_20511,N_20605);
or U20848 (N_20848,N_20742,N_20532);
nand U20849 (N_20849,N_20652,N_20553);
and U20850 (N_20850,N_20708,N_20537);
xor U20851 (N_20851,N_20576,N_20502);
nor U20852 (N_20852,N_20695,N_20653);
xor U20853 (N_20853,N_20590,N_20580);
or U20854 (N_20854,N_20672,N_20651);
or U20855 (N_20855,N_20744,N_20679);
or U20856 (N_20856,N_20503,N_20508);
and U20857 (N_20857,N_20550,N_20739);
xnor U20858 (N_20858,N_20673,N_20666);
and U20859 (N_20859,N_20562,N_20609);
nand U20860 (N_20860,N_20583,N_20603);
xnor U20861 (N_20861,N_20623,N_20526);
and U20862 (N_20862,N_20543,N_20626);
or U20863 (N_20863,N_20711,N_20721);
or U20864 (N_20864,N_20535,N_20743);
or U20865 (N_20865,N_20706,N_20657);
or U20866 (N_20866,N_20677,N_20634);
and U20867 (N_20867,N_20557,N_20509);
and U20868 (N_20868,N_20714,N_20561);
nand U20869 (N_20869,N_20542,N_20687);
or U20870 (N_20870,N_20588,N_20579);
xor U20871 (N_20871,N_20676,N_20647);
and U20872 (N_20872,N_20661,N_20656);
nand U20873 (N_20873,N_20578,N_20585);
xnor U20874 (N_20874,N_20723,N_20558);
or U20875 (N_20875,N_20534,N_20595);
xnor U20876 (N_20876,N_20728,N_20676);
and U20877 (N_20877,N_20549,N_20661);
xnor U20878 (N_20878,N_20733,N_20703);
xnor U20879 (N_20879,N_20680,N_20579);
nand U20880 (N_20880,N_20564,N_20707);
and U20881 (N_20881,N_20541,N_20681);
nand U20882 (N_20882,N_20718,N_20501);
xor U20883 (N_20883,N_20734,N_20661);
and U20884 (N_20884,N_20725,N_20610);
nand U20885 (N_20885,N_20563,N_20508);
or U20886 (N_20886,N_20524,N_20726);
nor U20887 (N_20887,N_20657,N_20609);
or U20888 (N_20888,N_20739,N_20622);
nand U20889 (N_20889,N_20709,N_20617);
xnor U20890 (N_20890,N_20545,N_20669);
or U20891 (N_20891,N_20733,N_20614);
nand U20892 (N_20892,N_20507,N_20730);
nand U20893 (N_20893,N_20733,N_20500);
xor U20894 (N_20894,N_20566,N_20547);
and U20895 (N_20895,N_20531,N_20559);
and U20896 (N_20896,N_20540,N_20616);
and U20897 (N_20897,N_20518,N_20536);
nand U20898 (N_20898,N_20598,N_20565);
nand U20899 (N_20899,N_20661,N_20610);
nand U20900 (N_20900,N_20639,N_20605);
nand U20901 (N_20901,N_20705,N_20699);
nand U20902 (N_20902,N_20646,N_20576);
or U20903 (N_20903,N_20715,N_20632);
or U20904 (N_20904,N_20584,N_20562);
nor U20905 (N_20905,N_20574,N_20508);
xnor U20906 (N_20906,N_20678,N_20662);
nand U20907 (N_20907,N_20685,N_20623);
or U20908 (N_20908,N_20725,N_20637);
nand U20909 (N_20909,N_20558,N_20601);
nand U20910 (N_20910,N_20632,N_20609);
nor U20911 (N_20911,N_20589,N_20646);
xnor U20912 (N_20912,N_20613,N_20506);
xnor U20913 (N_20913,N_20688,N_20646);
or U20914 (N_20914,N_20749,N_20676);
xor U20915 (N_20915,N_20599,N_20576);
nand U20916 (N_20916,N_20609,N_20615);
nor U20917 (N_20917,N_20722,N_20559);
and U20918 (N_20918,N_20632,N_20573);
or U20919 (N_20919,N_20588,N_20502);
nand U20920 (N_20920,N_20671,N_20530);
nand U20921 (N_20921,N_20557,N_20708);
and U20922 (N_20922,N_20662,N_20531);
or U20923 (N_20923,N_20584,N_20719);
nand U20924 (N_20924,N_20614,N_20729);
xor U20925 (N_20925,N_20670,N_20721);
nand U20926 (N_20926,N_20653,N_20578);
nand U20927 (N_20927,N_20730,N_20716);
nand U20928 (N_20928,N_20560,N_20565);
or U20929 (N_20929,N_20545,N_20630);
nor U20930 (N_20930,N_20633,N_20566);
or U20931 (N_20931,N_20635,N_20542);
nor U20932 (N_20932,N_20596,N_20597);
nor U20933 (N_20933,N_20717,N_20703);
and U20934 (N_20934,N_20545,N_20551);
or U20935 (N_20935,N_20748,N_20746);
nor U20936 (N_20936,N_20500,N_20716);
and U20937 (N_20937,N_20524,N_20513);
or U20938 (N_20938,N_20525,N_20600);
xnor U20939 (N_20939,N_20714,N_20503);
nand U20940 (N_20940,N_20542,N_20508);
or U20941 (N_20941,N_20631,N_20569);
nor U20942 (N_20942,N_20510,N_20518);
or U20943 (N_20943,N_20627,N_20549);
and U20944 (N_20944,N_20560,N_20685);
nor U20945 (N_20945,N_20684,N_20560);
or U20946 (N_20946,N_20703,N_20721);
nand U20947 (N_20947,N_20720,N_20555);
nor U20948 (N_20948,N_20699,N_20612);
xor U20949 (N_20949,N_20648,N_20585);
xnor U20950 (N_20950,N_20610,N_20573);
nor U20951 (N_20951,N_20547,N_20539);
or U20952 (N_20952,N_20583,N_20701);
and U20953 (N_20953,N_20531,N_20717);
xor U20954 (N_20954,N_20668,N_20591);
xor U20955 (N_20955,N_20748,N_20730);
or U20956 (N_20956,N_20505,N_20552);
or U20957 (N_20957,N_20581,N_20636);
nand U20958 (N_20958,N_20502,N_20687);
xnor U20959 (N_20959,N_20697,N_20560);
xnor U20960 (N_20960,N_20563,N_20626);
xor U20961 (N_20961,N_20600,N_20687);
xor U20962 (N_20962,N_20509,N_20622);
nor U20963 (N_20963,N_20586,N_20575);
and U20964 (N_20964,N_20557,N_20532);
nor U20965 (N_20965,N_20579,N_20547);
xnor U20966 (N_20966,N_20550,N_20659);
and U20967 (N_20967,N_20684,N_20703);
xor U20968 (N_20968,N_20631,N_20540);
and U20969 (N_20969,N_20620,N_20657);
and U20970 (N_20970,N_20589,N_20526);
or U20971 (N_20971,N_20649,N_20566);
or U20972 (N_20972,N_20567,N_20719);
and U20973 (N_20973,N_20526,N_20576);
xnor U20974 (N_20974,N_20616,N_20664);
nand U20975 (N_20975,N_20523,N_20542);
nand U20976 (N_20976,N_20671,N_20522);
or U20977 (N_20977,N_20606,N_20723);
or U20978 (N_20978,N_20732,N_20602);
and U20979 (N_20979,N_20529,N_20665);
nand U20980 (N_20980,N_20659,N_20641);
nand U20981 (N_20981,N_20596,N_20520);
nor U20982 (N_20982,N_20708,N_20680);
xnor U20983 (N_20983,N_20627,N_20546);
nand U20984 (N_20984,N_20549,N_20515);
xor U20985 (N_20985,N_20740,N_20553);
nor U20986 (N_20986,N_20604,N_20554);
nand U20987 (N_20987,N_20722,N_20734);
and U20988 (N_20988,N_20522,N_20557);
nor U20989 (N_20989,N_20577,N_20527);
or U20990 (N_20990,N_20725,N_20518);
or U20991 (N_20991,N_20519,N_20677);
or U20992 (N_20992,N_20622,N_20514);
and U20993 (N_20993,N_20703,N_20744);
nor U20994 (N_20994,N_20509,N_20684);
xor U20995 (N_20995,N_20621,N_20593);
nand U20996 (N_20996,N_20710,N_20510);
xor U20997 (N_20997,N_20577,N_20641);
or U20998 (N_20998,N_20692,N_20638);
or U20999 (N_20999,N_20696,N_20700);
or U21000 (N_21000,N_20908,N_20819);
and U21001 (N_21001,N_20751,N_20889);
and U21002 (N_21002,N_20887,N_20944);
and U21003 (N_21003,N_20897,N_20938);
or U21004 (N_21004,N_20785,N_20939);
and U21005 (N_21005,N_20970,N_20972);
or U21006 (N_21006,N_20998,N_20806);
nand U21007 (N_21007,N_20913,N_20846);
nor U21008 (N_21008,N_20865,N_20779);
nor U21009 (N_21009,N_20898,N_20880);
nor U21010 (N_21010,N_20832,N_20901);
nor U21011 (N_21011,N_20885,N_20965);
or U21012 (N_21012,N_20888,N_20878);
and U21013 (N_21013,N_20823,N_20780);
or U21014 (N_21014,N_20951,N_20886);
and U21015 (N_21015,N_20936,N_20852);
or U21016 (N_21016,N_20877,N_20802);
nor U21017 (N_21017,N_20816,N_20962);
xnor U21018 (N_21018,N_20811,N_20989);
xor U21019 (N_21019,N_20827,N_20862);
and U21020 (N_21020,N_20871,N_20756);
nor U21021 (N_21021,N_20836,N_20818);
or U21022 (N_21022,N_20991,N_20789);
nor U21023 (N_21023,N_20905,N_20792);
or U21024 (N_21024,N_20800,N_20853);
and U21025 (N_21025,N_20782,N_20775);
xnor U21026 (N_21026,N_20845,N_20955);
xnor U21027 (N_21027,N_20803,N_20759);
nor U21028 (N_21028,N_20860,N_20809);
nor U21029 (N_21029,N_20801,N_20883);
nor U21030 (N_21030,N_20837,N_20796);
nand U21031 (N_21031,N_20863,N_20753);
nor U21032 (N_21032,N_20956,N_20899);
or U21033 (N_21033,N_20927,N_20879);
and U21034 (N_21034,N_20769,N_20873);
and U21035 (N_21035,N_20976,N_20842);
or U21036 (N_21036,N_20934,N_20866);
and U21037 (N_21037,N_20850,N_20907);
or U21038 (N_21038,N_20984,N_20834);
nand U21039 (N_21039,N_20930,N_20847);
nand U21040 (N_21040,N_20815,N_20754);
or U21041 (N_21041,N_20781,N_20813);
nor U21042 (N_21042,N_20969,N_20774);
nand U21043 (N_21043,N_20841,N_20963);
or U21044 (N_21044,N_20896,N_20903);
or U21045 (N_21045,N_20977,N_20791);
and U21046 (N_21046,N_20824,N_20917);
nor U21047 (N_21047,N_20990,N_20752);
nor U21048 (N_21048,N_20855,N_20904);
nand U21049 (N_21049,N_20857,N_20831);
xor U21050 (N_21050,N_20919,N_20912);
or U21051 (N_21051,N_20999,N_20966);
nor U21052 (N_21052,N_20922,N_20772);
nand U21053 (N_21053,N_20778,N_20861);
nand U21054 (N_21054,N_20942,N_20961);
nor U21055 (N_21055,N_20994,N_20967);
nor U21056 (N_21056,N_20915,N_20825);
xnor U21057 (N_21057,N_20985,N_20810);
or U21058 (N_21058,N_20884,N_20892);
or U21059 (N_21059,N_20833,N_20790);
and U21060 (N_21060,N_20854,N_20949);
xor U21061 (N_21061,N_20788,N_20768);
xor U21062 (N_21062,N_20840,N_20895);
and U21063 (N_21063,N_20996,N_20914);
xor U21064 (N_21064,N_20925,N_20902);
xnor U21065 (N_21065,N_20900,N_20805);
nor U21066 (N_21066,N_20876,N_20979);
or U21067 (N_21067,N_20858,N_20867);
xnor U21068 (N_21068,N_20968,N_20997);
nand U21069 (N_21069,N_20807,N_20766);
xnor U21070 (N_21070,N_20828,N_20973);
nor U21071 (N_21071,N_20909,N_20921);
or U21072 (N_21072,N_20926,N_20808);
and U21073 (N_21073,N_20839,N_20987);
xnor U21074 (N_21074,N_20763,N_20954);
and U21075 (N_21075,N_20767,N_20964);
or U21076 (N_21076,N_20993,N_20894);
nor U21077 (N_21077,N_20812,N_20870);
or U21078 (N_21078,N_20829,N_20765);
and U21079 (N_21079,N_20771,N_20817);
nand U21080 (N_21080,N_20992,N_20799);
nand U21081 (N_21081,N_20868,N_20856);
nand U21082 (N_21082,N_20760,N_20947);
xnor U21083 (N_21083,N_20764,N_20821);
nor U21084 (N_21084,N_20783,N_20822);
nand U21085 (N_21085,N_20761,N_20770);
nand U21086 (N_21086,N_20784,N_20950);
or U21087 (N_21087,N_20794,N_20875);
nand U21088 (N_21088,N_20755,N_20835);
xor U21089 (N_21089,N_20971,N_20940);
or U21090 (N_21090,N_20932,N_20981);
nand U21091 (N_21091,N_20838,N_20787);
xor U21092 (N_21092,N_20804,N_20959);
nand U21093 (N_21093,N_20978,N_20937);
or U21094 (N_21094,N_20982,N_20757);
and U21095 (N_21095,N_20891,N_20980);
or U21096 (N_21096,N_20859,N_20975);
or U21097 (N_21097,N_20906,N_20928);
and U21098 (N_21098,N_20952,N_20820);
nor U21099 (N_21099,N_20974,N_20797);
and U21100 (N_21100,N_20988,N_20957);
and U21101 (N_21101,N_20777,N_20893);
nor U21102 (N_21102,N_20986,N_20793);
nor U21103 (N_21103,N_20776,N_20941);
nand U21104 (N_21104,N_20848,N_20948);
nand U21105 (N_21105,N_20851,N_20798);
and U21106 (N_21106,N_20874,N_20983);
and U21107 (N_21107,N_20864,N_20814);
and U21108 (N_21108,N_20960,N_20931);
or U21109 (N_21109,N_20943,N_20935);
or U21110 (N_21110,N_20830,N_20924);
xor U21111 (N_21111,N_20918,N_20995);
nor U21112 (N_21112,N_20881,N_20758);
nand U21113 (N_21113,N_20958,N_20849);
or U21114 (N_21114,N_20795,N_20872);
nor U21115 (N_21115,N_20773,N_20916);
xor U21116 (N_21116,N_20910,N_20920);
nor U21117 (N_21117,N_20826,N_20869);
or U21118 (N_21118,N_20923,N_20786);
or U21119 (N_21119,N_20844,N_20762);
nand U21120 (N_21120,N_20953,N_20911);
nand U21121 (N_21121,N_20750,N_20890);
nor U21122 (N_21122,N_20929,N_20882);
or U21123 (N_21123,N_20933,N_20946);
and U21124 (N_21124,N_20945,N_20843);
nand U21125 (N_21125,N_20851,N_20781);
nand U21126 (N_21126,N_20896,N_20993);
or U21127 (N_21127,N_20818,N_20928);
or U21128 (N_21128,N_20918,N_20789);
and U21129 (N_21129,N_20944,N_20991);
xnor U21130 (N_21130,N_20967,N_20901);
nor U21131 (N_21131,N_20889,N_20888);
xnor U21132 (N_21132,N_20963,N_20762);
nor U21133 (N_21133,N_20969,N_20847);
xnor U21134 (N_21134,N_20750,N_20830);
and U21135 (N_21135,N_20969,N_20951);
or U21136 (N_21136,N_20938,N_20844);
xnor U21137 (N_21137,N_20856,N_20981);
nand U21138 (N_21138,N_20954,N_20995);
nor U21139 (N_21139,N_20865,N_20917);
and U21140 (N_21140,N_20852,N_20890);
or U21141 (N_21141,N_20995,N_20962);
nor U21142 (N_21142,N_20992,N_20964);
nor U21143 (N_21143,N_20988,N_20765);
nand U21144 (N_21144,N_20780,N_20875);
and U21145 (N_21145,N_20916,N_20962);
nand U21146 (N_21146,N_20899,N_20823);
xnor U21147 (N_21147,N_20949,N_20765);
nand U21148 (N_21148,N_20869,N_20816);
nand U21149 (N_21149,N_20944,N_20819);
or U21150 (N_21150,N_20863,N_20999);
nand U21151 (N_21151,N_20955,N_20840);
nor U21152 (N_21152,N_20993,N_20998);
nor U21153 (N_21153,N_20885,N_20811);
nor U21154 (N_21154,N_20895,N_20893);
nor U21155 (N_21155,N_20786,N_20936);
nand U21156 (N_21156,N_20875,N_20873);
nor U21157 (N_21157,N_20980,N_20880);
and U21158 (N_21158,N_20762,N_20759);
nor U21159 (N_21159,N_20854,N_20978);
nor U21160 (N_21160,N_20955,N_20778);
xor U21161 (N_21161,N_20896,N_20872);
nand U21162 (N_21162,N_20915,N_20842);
and U21163 (N_21163,N_20984,N_20770);
xor U21164 (N_21164,N_20876,N_20975);
or U21165 (N_21165,N_20778,N_20967);
and U21166 (N_21166,N_20759,N_20994);
xor U21167 (N_21167,N_20765,N_20976);
xnor U21168 (N_21168,N_20838,N_20998);
and U21169 (N_21169,N_20932,N_20895);
and U21170 (N_21170,N_20838,N_20869);
xor U21171 (N_21171,N_20983,N_20927);
or U21172 (N_21172,N_20756,N_20790);
nand U21173 (N_21173,N_20816,N_20950);
or U21174 (N_21174,N_20879,N_20888);
xor U21175 (N_21175,N_20916,N_20897);
nand U21176 (N_21176,N_20906,N_20868);
nand U21177 (N_21177,N_20855,N_20947);
nand U21178 (N_21178,N_20904,N_20924);
and U21179 (N_21179,N_20932,N_20859);
nor U21180 (N_21180,N_20803,N_20877);
and U21181 (N_21181,N_20890,N_20889);
xnor U21182 (N_21182,N_20845,N_20775);
nand U21183 (N_21183,N_20806,N_20934);
nand U21184 (N_21184,N_20792,N_20868);
nand U21185 (N_21185,N_20942,N_20762);
nand U21186 (N_21186,N_20903,N_20880);
xnor U21187 (N_21187,N_20870,N_20816);
nor U21188 (N_21188,N_20805,N_20772);
and U21189 (N_21189,N_20789,N_20949);
nand U21190 (N_21190,N_20942,N_20841);
xor U21191 (N_21191,N_20845,N_20900);
nand U21192 (N_21192,N_20818,N_20760);
xnor U21193 (N_21193,N_20758,N_20977);
nand U21194 (N_21194,N_20852,N_20791);
xnor U21195 (N_21195,N_20833,N_20945);
xnor U21196 (N_21196,N_20885,N_20797);
or U21197 (N_21197,N_20910,N_20856);
or U21198 (N_21198,N_20992,N_20989);
nor U21199 (N_21199,N_20891,N_20777);
xnor U21200 (N_21200,N_20873,N_20891);
or U21201 (N_21201,N_20964,N_20987);
xnor U21202 (N_21202,N_20783,N_20789);
nor U21203 (N_21203,N_20759,N_20909);
or U21204 (N_21204,N_20881,N_20925);
and U21205 (N_21205,N_20955,N_20931);
and U21206 (N_21206,N_20891,N_20947);
nand U21207 (N_21207,N_20894,N_20790);
nand U21208 (N_21208,N_20797,N_20949);
nor U21209 (N_21209,N_20991,N_20895);
nand U21210 (N_21210,N_20799,N_20873);
nand U21211 (N_21211,N_20964,N_20799);
nor U21212 (N_21212,N_20943,N_20985);
nand U21213 (N_21213,N_20964,N_20916);
nand U21214 (N_21214,N_20871,N_20824);
xnor U21215 (N_21215,N_20856,N_20798);
nand U21216 (N_21216,N_20816,N_20804);
xor U21217 (N_21217,N_20941,N_20821);
and U21218 (N_21218,N_20837,N_20794);
xor U21219 (N_21219,N_20968,N_20893);
nor U21220 (N_21220,N_20764,N_20986);
xnor U21221 (N_21221,N_20942,N_20901);
or U21222 (N_21222,N_20984,N_20871);
or U21223 (N_21223,N_20764,N_20853);
nand U21224 (N_21224,N_20874,N_20847);
and U21225 (N_21225,N_20781,N_20935);
and U21226 (N_21226,N_20998,N_20758);
xnor U21227 (N_21227,N_20799,N_20936);
nand U21228 (N_21228,N_20901,N_20795);
and U21229 (N_21229,N_20917,N_20953);
nand U21230 (N_21230,N_20923,N_20776);
nor U21231 (N_21231,N_20858,N_20906);
and U21232 (N_21232,N_20873,N_20976);
and U21233 (N_21233,N_20936,N_20815);
nor U21234 (N_21234,N_20923,N_20937);
nor U21235 (N_21235,N_20974,N_20942);
and U21236 (N_21236,N_20835,N_20805);
nand U21237 (N_21237,N_20858,N_20802);
nand U21238 (N_21238,N_20949,N_20900);
or U21239 (N_21239,N_20768,N_20948);
xnor U21240 (N_21240,N_20758,N_20798);
xnor U21241 (N_21241,N_20975,N_20820);
nand U21242 (N_21242,N_20792,N_20766);
or U21243 (N_21243,N_20871,N_20961);
nor U21244 (N_21244,N_20919,N_20954);
nand U21245 (N_21245,N_20915,N_20763);
or U21246 (N_21246,N_20945,N_20975);
or U21247 (N_21247,N_20808,N_20894);
or U21248 (N_21248,N_20853,N_20768);
or U21249 (N_21249,N_20913,N_20990);
nor U21250 (N_21250,N_21018,N_21225);
nor U21251 (N_21251,N_21131,N_21129);
and U21252 (N_21252,N_21040,N_21221);
nor U21253 (N_21253,N_21033,N_21244);
and U21254 (N_21254,N_21156,N_21092);
or U21255 (N_21255,N_21005,N_21003);
nor U21256 (N_21256,N_21114,N_21211);
or U21257 (N_21257,N_21057,N_21187);
nand U21258 (N_21258,N_21107,N_21193);
or U21259 (N_21259,N_21242,N_21084);
nand U21260 (N_21260,N_21170,N_21215);
xor U21261 (N_21261,N_21121,N_21100);
and U21262 (N_21262,N_21074,N_21024);
nor U21263 (N_21263,N_21214,N_21019);
nor U21264 (N_21264,N_21041,N_21171);
and U21265 (N_21265,N_21063,N_21046);
or U21266 (N_21266,N_21134,N_21197);
nand U21267 (N_21267,N_21076,N_21035);
nand U21268 (N_21268,N_21128,N_21054);
nand U21269 (N_21269,N_21227,N_21009);
or U21270 (N_21270,N_21031,N_21233);
xnor U21271 (N_21271,N_21199,N_21159);
or U21272 (N_21272,N_21115,N_21013);
or U21273 (N_21273,N_21038,N_21079);
nor U21274 (N_21274,N_21144,N_21202);
xor U21275 (N_21275,N_21090,N_21234);
nand U21276 (N_21276,N_21167,N_21010);
and U21277 (N_21277,N_21047,N_21027);
or U21278 (N_21278,N_21042,N_21068);
and U21279 (N_21279,N_21058,N_21248);
xnor U21280 (N_21280,N_21191,N_21142);
xnor U21281 (N_21281,N_21071,N_21062);
or U21282 (N_21282,N_21070,N_21103);
nand U21283 (N_21283,N_21116,N_21162);
nor U21284 (N_21284,N_21059,N_21026);
and U21285 (N_21285,N_21056,N_21188);
nand U21286 (N_21286,N_21238,N_21241);
or U21287 (N_21287,N_21016,N_21132);
or U21288 (N_21288,N_21133,N_21184);
nand U21289 (N_21289,N_21179,N_21011);
or U21290 (N_21290,N_21138,N_21164);
nand U21291 (N_21291,N_21039,N_21205);
and U21292 (N_21292,N_21152,N_21073);
or U21293 (N_21293,N_21219,N_21212);
or U21294 (N_21294,N_21029,N_21185);
nand U21295 (N_21295,N_21022,N_21078);
nor U21296 (N_21296,N_21143,N_21086);
and U21297 (N_21297,N_21136,N_21232);
or U21298 (N_21298,N_21077,N_21083);
xor U21299 (N_21299,N_21175,N_21108);
nand U21300 (N_21300,N_21190,N_21235);
or U21301 (N_21301,N_21135,N_21036);
nor U21302 (N_21302,N_21157,N_21120);
nor U21303 (N_21303,N_21081,N_21025);
xnor U21304 (N_21304,N_21240,N_21151);
xnor U21305 (N_21305,N_21109,N_21066);
nor U21306 (N_21306,N_21126,N_21186);
xor U21307 (N_21307,N_21180,N_21168);
or U21308 (N_21308,N_21158,N_21097);
xor U21309 (N_21309,N_21204,N_21220);
nor U21310 (N_21310,N_21080,N_21200);
nand U21311 (N_21311,N_21223,N_21122);
nor U21312 (N_21312,N_21236,N_21119);
nor U21313 (N_21313,N_21196,N_21239);
xor U21314 (N_21314,N_21094,N_21111);
nor U21315 (N_21315,N_21104,N_21194);
and U21316 (N_21316,N_21049,N_21161);
xor U21317 (N_21317,N_21243,N_21087);
nand U21318 (N_21318,N_21028,N_21048);
and U21319 (N_21319,N_21072,N_21014);
xnor U21320 (N_21320,N_21127,N_21209);
nor U21321 (N_21321,N_21069,N_21213);
xnor U21322 (N_21322,N_21166,N_21043);
nand U21323 (N_21323,N_21089,N_21002);
and U21324 (N_21324,N_21224,N_21163);
nand U21325 (N_21325,N_21230,N_21125);
nor U21326 (N_21326,N_21155,N_21008);
and U21327 (N_21327,N_21141,N_21117);
nand U21328 (N_21328,N_21137,N_21247);
xnor U21329 (N_21329,N_21249,N_21237);
nor U21330 (N_21330,N_21000,N_21096);
xnor U21331 (N_21331,N_21004,N_21021);
nand U21332 (N_21332,N_21091,N_21061);
nor U21333 (N_21333,N_21140,N_21044);
or U21334 (N_21334,N_21208,N_21206);
nand U21335 (N_21335,N_21055,N_21112);
nor U21336 (N_21336,N_21075,N_21006);
and U21337 (N_21337,N_21139,N_21160);
and U21338 (N_21338,N_21053,N_21015);
nand U21339 (N_21339,N_21174,N_21101);
nand U21340 (N_21340,N_21182,N_21098);
or U21341 (N_21341,N_21037,N_21201);
nand U21342 (N_21342,N_21123,N_21001);
nor U21343 (N_21343,N_21034,N_21085);
xor U21344 (N_21344,N_21050,N_21118);
xor U21345 (N_21345,N_21088,N_21229);
nand U21346 (N_21346,N_21246,N_21183);
and U21347 (N_21347,N_21231,N_21023);
nor U21348 (N_21348,N_21195,N_21217);
nor U21349 (N_21349,N_21222,N_21192);
nor U21350 (N_21350,N_21177,N_21130);
nor U21351 (N_21351,N_21150,N_21095);
and U21352 (N_21352,N_21113,N_21060);
nand U21353 (N_21353,N_21189,N_21124);
nor U21354 (N_21354,N_21169,N_21012);
nor U21355 (N_21355,N_21203,N_21228);
or U21356 (N_21356,N_21145,N_21045);
nand U21357 (N_21357,N_21153,N_21065);
nor U21358 (N_21358,N_21218,N_21030);
xnor U21359 (N_21359,N_21020,N_21165);
and U21360 (N_21360,N_21176,N_21052);
nand U21361 (N_21361,N_21093,N_21181);
or U21362 (N_21362,N_21017,N_21064);
xnor U21363 (N_21363,N_21051,N_21106);
and U21364 (N_21364,N_21226,N_21198);
or U21365 (N_21365,N_21148,N_21032);
nor U21366 (N_21366,N_21207,N_21210);
or U21367 (N_21367,N_21099,N_21067);
xor U21368 (N_21368,N_21147,N_21149);
nor U21369 (N_21369,N_21110,N_21172);
xnor U21370 (N_21370,N_21007,N_21173);
nand U21371 (N_21371,N_21245,N_21146);
nand U21372 (N_21372,N_21154,N_21105);
xor U21373 (N_21373,N_21082,N_21216);
or U21374 (N_21374,N_21178,N_21102);
xnor U21375 (N_21375,N_21015,N_21104);
nor U21376 (N_21376,N_21210,N_21102);
or U21377 (N_21377,N_21072,N_21036);
nand U21378 (N_21378,N_21122,N_21004);
or U21379 (N_21379,N_21248,N_21121);
nand U21380 (N_21380,N_21135,N_21200);
xnor U21381 (N_21381,N_21139,N_21085);
nor U21382 (N_21382,N_21107,N_21087);
nor U21383 (N_21383,N_21203,N_21073);
and U21384 (N_21384,N_21202,N_21204);
nand U21385 (N_21385,N_21183,N_21033);
xor U21386 (N_21386,N_21236,N_21148);
nand U21387 (N_21387,N_21201,N_21203);
and U21388 (N_21388,N_21085,N_21146);
nand U21389 (N_21389,N_21091,N_21194);
nand U21390 (N_21390,N_21100,N_21067);
nand U21391 (N_21391,N_21164,N_21049);
xor U21392 (N_21392,N_21117,N_21047);
nand U21393 (N_21393,N_21170,N_21133);
nor U21394 (N_21394,N_21005,N_21083);
nand U21395 (N_21395,N_21117,N_21155);
or U21396 (N_21396,N_21063,N_21043);
xnor U21397 (N_21397,N_21196,N_21248);
and U21398 (N_21398,N_21225,N_21056);
nor U21399 (N_21399,N_21137,N_21001);
nand U21400 (N_21400,N_21141,N_21089);
and U21401 (N_21401,N_21212,N_21214);
xnor U21402 (N_21402,N_21118,N_21088);
or U21403 (N_21403,N_21015,N_21055);
nand U21404 (N_21404,N_21108,N_21240);
or U21405 (N_21405,N_21187,N_21007);
nand U21406 (N_21406,N_21247,N_21124);
nor U21407 (N_21407,N_21090,N_21102);
xor U21408 (N_21408,N_21147,N_21173);
nor U21409 (N_21409,N_21146,N_21166);
and U21410 (N_21410,N_21058,N_21215);
or U21411 (N_21411,N_21097,N_21225);
nand U21412 (N_21412,N_21048,N_21153);
nand U21413 (N_21413,N_21224,N_21105);
nor U21414 (N_21414,N_21016,N_21024);
or U21415 (N_21415,N_21095,N_21059);
and U21416 (N_21416,N_21201,N_21225);
nor U21417 (N_21417,N_21143,N_21055);
or U21418 (N_21418,N_21077,N_21110);
nor U21419 (N_21419,N_21111,N_21243);
nand U21420 (N_21420,N_21202,N_21066);
nand U21421 (N_21421,N_21142,N_21199);
xor U21422 (N_21422,N_21221,N_21023);
xor U21423 (N_21423,N_21234,N_21142);
or U21424 (N_21424,N_21169,N_21015);
and U21425 (N_21425,N_21161,N_21247);
nand U21426 (N_21426,N_21140,N_21109);
or U21427 (N_21427,N_21197,N_21186);
nor U21428 (N_21428,N_21011,N_21116);
nor U21429 (N_21429,N_21078,N_21197);
and U21430 (N_21430,N_21126,N_21178);
nand U21431 (N_21431,N_21146,N_21185);
or U21432 (N_21432,N_21073,N_21122);
and U21433 (N_21433,N_21113,N_21212);
nor U21434 (N_21434,N_21089,N_21150);
xnor U21435 (N_21435,N_21064,N_21232);
nor U21436 (N_21436,N_21141,N_21132);
nand U21437 (N_21437,N_21000,N_21220);
nand U21438 (N_21438,N_21113,N_21201);
nand U21439 (N_21439,N_21244,N_21134);
or U21440 (N_21440,N_21026,N_21054);
xor U21441 (N_21441,N_21153,N_21192);
nand U21442 (N_21442,N_21141,N_21100);
nand U21443 (N_21443,N_21054,N_21002);
and U21444 (N_21444,N_21229,N_21075);
or U21445 (N_21445,N_21232,N_21045);
or U21446 (N_21446,N_21097,N_21220);
and U21447 (N_21447,N_21087,N_21233);
nand U21448 (N_21448,N_21075,N_21053);
nand U21449 (N_21449,N_21022,N_21216);
and U21450 (N_21450,N_21186,N_21062);
nor U21451 (N_21451,N_21088,N_21052);
xnor U21452 (N_21452,N_21199,N_21029);
nand U21453 (N_21453,N_21000,N_21141);
xnor U21454 (N_21454,N_21054,N_21038);
or U21455 (N_21455,N_21150,N_21179);
or U21456 (N_21456,N_21028,N_21145);
xnor U21457 (N_21457,N_21084,N_21007);
or U21458 (N_21458,N_21146,N_21010);
nand U21459 (N_21459,N_21162,N_21083);
xor U21460 (N_21460,N_21059,N_21199);
or U21461 (N_21461,N_21145,N_21219);
nor U21462 (N_21462,N_21035,N_21015);
xor U21463 (N_21463,N_21065,N_21056);
or U21464 (N_21464,N_21153,N_21143);
xor U21465 (N_21465,N_21035,N_21100);
or U21466 (N_21466,N_21213,N_21216);
xnor U21467 (N_21467,N_21055,N_21178);
nor U21468 (N_21468,N_21146,N_21156);
nand U21469 (N_21469,N_21138,N_21099);
and U21470 (N_21470,N_21220,N_21159);
nand U21471 (N_21471,N_21151,N_21128);
nand U21472 (N_21472,N_21168,N_21116);
xnor U21473 (N_21473,N_21018,N_21211);
or U21474 (N_21474,N_21168,N_21204);
or U21475 (N_21475,N_21233,N_21004);
nand U21476 (N_21476,N_21127,N_21030);
and U21477 (N_21477,N_21009,N_21120);
xnor U21478 (N_21478,N_21219,N_21074);
and U21479 (N_21479,N_21131,N_21162);
nand U21480 (N_21480,N_21089,N_21238);
xnor U21481 (N_21481,N_21084,N_21113);
or U21482 (N_21482,N_21118,N_21072);
nor U21483 (N_21483,N_21155,N_21245);
and U21484 (N_21484,N_21080,N_21203);
nand U21485 (N_21485,N_21018,N_21030);
and U21486 (N_21486,N_21046,N_21061);
or U21487 (N_21487,N_21192,N_21204);
or U21488 (N_21488,N_21008,N_21178);
nand U21489 (N_21489,N_21110,N_21013);
and U21490 (N_21490,N_21047,N_21223);
nor U21491 (N_21491,N_21089,N_21134);
nand U21492 (N_21492,N_21241,N_21040);
and U21493 (N_21493,N_21233,N_21030);
nand U21494 (N_21494,N_21221,N_21164);
xnor U21495 (N_21495,N_21002,N_21141);
xor U21496 (N_21496,N_21031,N_21206);
or U21497 (N_21497,N_21192,N_21034);
and U21498 (N_21498,N_21047,N_21137);
or U21499 (N_21499,N_21095,N_21222);
and U21500 (N_21500,N_21375,N_21289);
nand U21501 (N_21501,N_21314,N_21354);
or U21502 (N_21502,N_21499,N_21473);
nor U21503 (N_21503,N_21295,N_21258);
and U21504 (N_21504,N_21411,N_21262);
xor U21505 (N_21505,N_21429,N_21460);
nand U21506 (N_21506,N_21303,N_21488);
nor U21507 (N_21507,N_21260,N_21335);
and U21508 (N_21508,N_21498,N_21450);
nand U21509 (N_21509,N_21485,N_21370);
xor U21510 (N_21510,N_21472,N_21377);
xnor U21511 (N_21511,N_21478,N_21300);
and U21512 (N_21512,N_21394,N_21287);
or U21513 (N_21513,N_21313,N_21468);
and U21514 (N_21514,N_21463,N_21364);
nand U21515 (N_21515,N_21469,N_21481);
and U21516 (N_21516,N_21366,N_21284);
or U21517 (N_21517,N_21269,N_21448);
and U21518 (N_21518,N_21343,N_21348);
nand U21519 (N_21519,N_21355,N_21255);
and U21520 (N_21520,N_21334,N_21261);
and U21521 (N_21521,N_21387,N_21357);
and U21522 (N_21522,N_21495,N_21346);
nor U21523 (N_21523,N_21254,N_21321);
nor U21524 (N_21524,N_21333,N_21363);
nand U21525 (N_21525,N_21476,N_21471);
xor U21526 (N_21526,N_21421,N_21270);
or U21527 (N_21527,N_21286,N_21408);
and U21528 (N_21528,N_21386,N_21332);
xnor U21529 (N_21529,N_21256,N_21441);
nand U21530 (N_21530,N_21446,N_21442);
or U21531 (N_21531,N_21497,N_21492);
nor U21532 (N_21532,N_21279,N_21268);
nand U21533 (N_21533,N_21414,N_21470);
nand U21534 (N_21534,N_21385,N_21451);
and U21535 (N_21535,N_21445,N_21416);
and U21536 (N_21536,N_21291,N_21253);
xnor U21537 (N_21537,N_21358,N_21402);
xnor U21538 (N_21538,N_21338,N_21317);
xor U21539 (N_21539,N_21439,N_21412);
and U21540 (N_21540,N_21459,N_21323);
and U21541 (N_21541,N_21331,N_21360);
nor U21542 (N_21542,N_21444,N_21349);
nor U21543 (N_21543,N_21251,N_21480);
and U21544 (N_21544,N_21409,N_21252);
nor U21545 (N_21545,N_21455,N_21318);
nor U21546 (N_21546,N_21427,N_21456);
xnor U21547 (N_21547,N_21423,N_21352);
and U21548 (N_21548,N_21462,N_21329);
nand U21549 (N_21549,N_21401,N_21307);
nor U21550 (N_21550,N_21336,N_21272);
or U21551 (N_21551,N_21482,N_21322);
nand U21552 (N_21552,N_21280,N_21337);
nor U21553 (N_21553,N_21396,N_21304);
nand U21554 (N_21554,N_21452,N_21486);
nand U21555 (N_21555,N_21381,N_21432);
or U21556 (N_21556,N_21392,N_21418);
xnor U21557 (N_21557,N_21404,N_21426);
xnor U21558 (N_21558,N_21433,N_21373);
and U21559 (N_21559,N_21431,N_21413);
and U21560 (N_21560,N_21395,N_21312);
nand U21561 (N_21561,N_21285,N_21308);
nand U21562 (N_21562,N_21440,N_21388);
or U21563 (N_21563,N_21449,N_21368);
and U21564 (N_21564,N_21400,N_21467);
xor U21565 (N_21565,N_21290,N_21250);
nor U21566 (N_21566,N_21484,N_21430);
xnor U21567 (N_21567,N_21325,N_21361);
or U21568 (N_21568,N_21393,N_21496);
xor U21569 (N_21569,N_21405,N_21309);
nand U21570 (N_21570,N_21347,N_21424);
xnor U21571 (N_21571,N_21390,N_21382);
xor U21572 (N_21572,N_21457,N_21282);
nand U21573 (N_21573,N_21376,N_21417);
or U21574 (N_21574,N_21380,N_21410);
nor U21575 (N_21575,N_21437,N_21297);
and U21576 (N_21576,N_21397,N_21320);
or U21577 (N_21577,N_21491,N_21306);
xor U21578 (N_21578,N_21453,N_21454);
xor U21579 (N_21579,N_21327,N_21428);
or U21580 (N_21580,N_21461,N_21316);
and U21581 (N_21581,N_21464,N_21435);
xnor U21582 (N_21582,N_21425,N_21275);
nor U21583 (N_21583,N_21447,N_21281);
nand U21584 (N_21584,N_21378,N_21293);
nor U21585 (N_21585,N_21379,N_21294);
or U21586 (N_21586,N_21266,N_21351);
nor U21587 (N_21587,N_21436,N_21443);
or U21588 (N_21588,N_21399,N_21257);
nor U21589 (N_21589,N_21438,N_21479);
nand U21590 (N_21590,N_21362,N_21263);
nor U21591 (N_21591,N_21276,N_21367);
or U21592 (N_21592,N_21489,N_21383);
or U21593 (N_21593,N_21434,N_21345);
xnor U21594 (N_21594,N_21391,N_21301);
xnor U21595 (N_21595,N_21296,N_21465);
nor U21596 (N_21596,N_21371,N_21356);
or U21597 (N_21597,N_21330,N_21283);
and U21598 (N_21598,N_21340,N_21483);
nand U21599 (N_21599,N_21415,N_21277);
nand U21600 (N_21600,N_21372,N_21288);
xnor U21601 (N_21601,N_21477,N_21389);
and U21602 (N_21602,N_21458,N_21422);
xnor U21603 (N_21603,N_21302,N_21474);
nor U21604 (N_21604,N_21299,N_21292);
nor U21605 (N_21605,N_21305,N_21264);
or U21606 (N_21606,N_21315,N_21273);
and U21607 (N_21607,N_21328,N_21466);
and U21608 (N_21608,N_21311,N_21310);
xor U21609 (N_21609,N_21344,N_21494);
and U21610 (N_21610,N_21267,N_21319);
nand U21611 (N_21611,N_21324,N_21265);
nand U21612 (N_21612,N_21420,N_21398);
or U21613 (N_21613,N_21278,N_21419);
xnor U21614 (N_21614,N_21353,N_21274);
nand U21615 (N_21615,N_21342,N_21407);
and U21616 (N_21616,N_21341,N_21326);
nor U21617 (N_21617,N_21490,N_21259);
xnor U21618 (N_21618,N_21369,N_21487);
nand U21619 (N_21619,N_21350,N_21271);
nand U21620 (N_21620,N_21493,N_21359);
and U21621 (N_21621,N_21374,N_21475);
nand U21622 (N_21622,N_21365,N_21406);
nor U21623 (N_21623,N_21384,N_21403);
nand U21624 (N_21624,N_21298,N_21339);
or U21625 (N_21625,N_21362,N_21414);
nand U21626 (N_21626,N_21354,N_21489);
or U21627 (N_21627,N_21310,N_21429);
and U21628 (N_21628,N_21371,N_21421);
nor U21629 (N_21629,N_21259,N_21265);
or U21630 (N_21630,N_21296,N_21409);
nand U21631 (N_21631,N_21352,N_21348);
or U21632 (N_21632,N_21384,N_21382);
and U21633 (N_21633,N_21309,N_21315);
xor U21634 (N_21634,N_21469,N_21301);
and U21635 (N_21635,N_21447,N_21297);
xor U21636 (N_21636,N_21387,N_21334);
xnor U21637 (N_21637,N_21375,N_21350);
nand U21638 (N_21638,N_21424,N_21406);
and U21639 (N_21639,N_21290,N_21316);
nor U21640 (N_21640,N_21499,N_21469);
nor U21641 (N_21641,N_21330,N_21352);
or U21642 (N_21642,N_21454,N_21494);
xnor U21643 (N_21643,N_21416,N_21337);
and U21644 (N_21644,N_21341,N_21449);
or U21645 (N_21645,N_21398,N_21430);
and U21646 (N_21646,N_21455,N_21383);
xnor U21647 (N_21647,N_21399,N_21387);
nor U21648 (N_21648,N_21314,N_21327);
xor U21649 (N_21649,N_21474,N_21313);
and U21650 (N_21650,N_21298,N_21452);
and U21651 (N_21651,N_21443,N_21402);
xor U21652 (N_21652,N_21363,N_21358);
and U21653 (N_21653,N_21387,N_21276);
nand U21654 (N_21654,N_21266,N_21251);
nand U21655 (N_21655,N_21316,N_21297);
xor U21656 (N_21656,N_21327,N_21497);
nor U21657 (N_21657,N_21451,N_21438);
nor U21658 (N_21658,N_21302,N_21453);
or U21659 (N_21659,N_21363,N_21405);
xnor U21660 (N_21660,N_21391,N_21267);
and U21661 (N_21661,N_21470,N_21416);
xnor U21662 (N_21662,N_21372,N_21419);
xor U21663 (N_21663,N_21447,N_21250);
nor U21664 (N_21664,N_21298,N_21436);
xnor U21665 (N_21665,N_21432,N_21318);
nor U21666 (N_21666,N_21463,N_21399);
xnor U21667 (N_21667,N_21470,N_21267);
xnor U21668 (N_21668,N_21356,N_21435);
xnor U21669 (N_21669,N_21399,N_21441);
xor U21670 (N_21670,N_21381,N_21309);
nand U21671 (N_21671,N_21389,N_21424);
nor U21672 (N_21672,N_21430,N_21444);
nor U21673 (N_21673,N_21364,N_21443);
nor U21674 (N_21674,N_21313,N_21348);
xnor U21675 (N_21675,N_21287,N_21264);
and U21676 (N_21676,N_21276,N_21302);
nand U21677 (N_21677,N_21342,N_21301);
xor U21678 (N_21678,N_21470,N_21361);
and U21679 (N_21679,N_21399,N_21352);
xnor U21680 (N_21680,N_21373,N_21357);
xor U21681 (N_21681,N_21442,N_21375);
or U21682 (N_21682,N_21484,N_21337);
and U21683 (N_21683,N_21322,N_21465);
and U21684 (N_21684,N_21493,N_21326);
nand U21685 (N_21685,N_21490,N_21398);
nand U21686 (N_21686,N_21318,N_21352);
nand U21687 (N_21687,N_21318,N_21332);
or U21688 (N_21688,N_21403,N_21461);
xnor U21689 (N_21689,N_21320,N_21475);
or U21690 (N_21690,N_21465,N_21376);
and U21691 (N_21691,N_21452,N_21291);
and U21692 (N_21692,N_21359,N_21428);
nor U21693 (N_21693,N_21476,N_21403);
or U21694 (N_21694,N_21452,N_21333);
or U21695 (N_21695,N_21459,N_21448);
and U21696 (N_21696,N_21493,N_21356);
nand U21697 (N_21697,N_21304,N_21256);
xor U21698 (N_21698,N_21484,N_21365);
xor U21699 (N_21699,N_21432,N_21388);
xor U21700 (N_21700,N_21279,N_21416);
nor U21701 (N_21701,N_21348,N_21435);
or U21702 (N_21702,N_21278,N_21286);
nand U21703 (N_21703,N_21395,N_21440);
xor U21704 (N_21704,N_21424,N_21272);
and U21705 (N_21705,N_21332,N_21299);
nor U21706 (N_21706,N_21285,N_21493);
xnor U21707 (N_21707,N_21391,N_21362);
or U21708 (N_21708,N_21291,N_21297);
xor U21709 (N_21709,N_21311,N_21452);
nor U21710 (N_21710,N_21483,N_21405);
and U21711 (N_21711,N_21351,N_21449);
nor U21712 (N_21712,N_21465,N_21289);
and U21713 (N_21713,N_21347,N_21452);
and U21714 (N_21714,N_21458,N_21382);
nor U21715 (N_21715,N_21437,N_21350);
nand U21716 (N_21716,N_21387,N_21397);
nand U21717 (N_21717,N_21283,N_21300);
or U21718 (N_21718,N_21380,N_21313);
nor U21719 (N_21719,N_21398,N_21282);
nor U21720 (N_21720,N_21302,N_21361);
xnor U21721 (N_21721,N_21451,N_21289);
xnor U21722 (N_21722,N_21350,N_21301);
and U21723 (N_21723,N_21493,N_21374);
and U21724 (N_21724,N_21437,N_21338);
xor U21725 (N_21725,N_21434,N_21255);
or U21726 (N_21726,N_21416,N_21383);
xor U21727 (N_21727,N_21486,N_21257);
nand U21728 (N_21728,N_21358,N_21455);
nor U21729 (N_21729,N_21290,N_21382);
nor U21730 (N_21730,N_21429,N_21281);
nand U21731 (N_21731,N_21390,N_21463);
and U21732 (N_21732,N_21435,N_21460);
nor U21733 (N_21733,N_21321,N_21366);
and U21734 (N_21734,N_21348,N_21300);
nor U21735 (N_21735,N_21473,N_21251);
nor U21736 (N_21736,N_21459,N_21449);
nand U21737 (N_21737,N_21331,N_21477);
nand U21738 (N_21738,N_21427,N_21431);
xnor U21739 (N_21739,N_21310,N_21339);
nand U21740 (N_21740,N_21457,N_21425);
and U21741 (N_21741,N_21400,N_21302);
nor U21742 (N_21742,N_21286,N_21411);
xnor U21743 (N_21743,N_21352,N_21495);
nand U21744 (N_21744,N_21477,N_21413);
nand U21745 (N_21745,N_21272,N_21328);
and U21746 (N_21746,N_21485,N_21494);
or U21747 (N_21747,N_21389,N_21414);
xor U21748 (N_21748,N_21254,N_21427);
xnor U21749 (N_21749,N_21372,N_21268);
nand U21750 (N_21750,N_21688,N_21665);
and U21751 (N_21751,N_21593,N_21604);
xnor U21752 (N_21752,N_21612,N_21658);
nor U21753 (N_21753,N_21541,N_21502);
or U21754 (N_21754,N_21741,N_21747);
and U21755 (N_21755,N_21616,N_21729);
nand U21756 (N_21756,N_21673,N_21719);
xor U21757 (N_21757,N_21714,N_21618);
nor U21758 (N_21758,N_21503,N_21632);
or U21759 (N_21759,N_21651,N_21600);
nand U21760 (N_21760,N_21553,N_21574);
xor U21761 (N_21761,N_21685,N_21532);
xnor U21762 (N_21762,N_21596,N_21622);
xnor U21763 (N_21763,N_21543,N_21520);
and U21764 (N_21764,N_21583,N_21689);
or U21765 (N_21765,N_21672,N_21572);
nand U21766 (N_21766,N_21645,N_21744);
and U21767 (N_21767,N_21667,N_21670);
nor U21768 (N_21768,N_21569,N_21663);
nor U21769 (N_21769,N_21727,N_21587);
nand U21770 (N_21770,N_21546,N_21551);
nand U21771 (N_21771,N_21626,N_21695);
nor U21772 (N_21772,N_21599,N_21507);
or U21773 (N_21773,N_21606,N_21588);
nor U21774 (N_21774,N_21620,N_21723);
and U21775 (N_21775,N_21565,N_21701);
nand U21776 (N_21776,N_21563,N_21638);
or U21777 (N_21777,N_21571,N_21531);
nor U21778 (N_21778,N_21677,N_21713);
nand U21779 (N_21779,N_21630,N_21578);
nand U21780 (N_21780,N_21748,N_21740);
nand U21781 (N_21781,N_21611,N_21518);
nand U21782 (N_21782,N_21662,N_21666);
nand U21783 (N_21783,N_21627,N_21691);
xnor U21784 (N_21784,N_21609,N_21601);
nor U21785 (N_21785,N_21562,N_21697);
and U21786 (N_21786,N_21679,N_21653);
nand U21787 (N_21787,N_21680,N_21742);
and U21788 (N_21788,N_21500,N_21537);
nor U21789 (N_21789,N_21542,N_21581);
and U21790 (N_21790,N_21589,N_21560);
and U21791 (N_21791,N_21639,N_21700);
nor U21792 (N_21792,N_21633,N_21746);
nor U21793 (N_21793,N_21696,N_21635);
and U21794 (N_21794,N_21745,N_21538);
nand U21795 (N_21795,N_21624,N_21737);
nand U21796 (N_21796,N_21720,N_21504);
nand U21797 (N_21797,N_21711,N_21557);
nand U21798 (N_21798,N_21617,N_21660);
nor U21799 (N_21799,N_21684,N_21510);
nand U21800 (N_21800,N_21656,N_21530);
and U21801 (N_21801,N_21734,N_21704);
or U21802 (N_21802,N_21615,N_21647);
or U21803 (N_21803,N_21605,N_21725);
xnor U21804 (N_21804,N_21515,N_21570);
xor U21805 (N_21805,N_21568,N_21610);
and U21806 (N_21806,N_21548,N_21703);
xor U21807 (N_21807,N_21523,N_21642);
nand U21808 (N_21808,N_21580,N_21712);
nand U21809 (N_21809,N_21586,N_21527);
and U21810 (N_21810,N_21733,N_21702);
and U21811 (N_21811,N_21707,N_21694);
nor U21812 (N_21812,N_21501,N_21661);
or U21813 (N_21813,N_21674,N_21705);
nor U21814 (N_21814,N_21655,N_21514);
nand U21815 (N_21815,N_21577,N_21668);
xnor U21816 (N_21816,N_21631,N_21652);
nor U21817 (N_21817,N_21513,N_21607);
xor U21818 (N_21818,N_21634,N_21730);
and U21819 (N_21819,N_21613,N_21539);
nand U21820 (N_21820,N_21686,N_21693);
and U21821 (N_21821,N_21678,N_21636);
nor U21822 (N_21822,N_21575,N_21698);
nand U21823 (N_21823,N_21544,N_21650);
or U21824 (N_21824,N_21743,N_21640);
xor U21825 (N_21825,N_21594,N_21721);
and U21826 (N_21826,N_21726,N_21584);
nand U21827 (N_21827,N_21567,N_21681);
or U21828 (N_21828,N_21576,N_21718);
nor U21829 (N_21829,N_21554,N_21710);
nand U21830 (N_21830,N_21525,N_21536);
nor U21831 (N_21831,N_21722,N_21516);
nand U21832 (N_21832,N_21706,N_21508);
and U21833 (N_21833,N_21545,N_21534);
or U21834 (N_21834,N_21522,N_21724);
and U21835 (N_21835,N_21590,N_21728);
nor U21836 (N_21836,N_21597,N_21558);
or U21837 (N_21837,N_21731,N_21664);
xor U21838 (N_21838,N_21659,N_21708);
or U21839 (N_21839,N_21529,N_21669);
xor U21840 (N_21840,N_21509,N_21732);
nand U21841 (N_21841,N_21716,N_21547);
nor U21842 (N_21842,N_21511,N_21552);
xor U21843 (N_21843,N_21619,N_21559);
nor U21844 (N_21844,N_21749,N_21550);
nand U21845 (N_21845,N_21564,N_21592);
nor U21846 (N_21846,N_21598,N_21629);
or U21847 (N_21847,N_21526,N_21528);
or U21848 (N_21848,N_21505,N_21585);
or U21849 (N_21849,N_21643,N_21683);
nand U21850 (N_21850,N_21649,N_21517);
and U21851 (N_21851,N_21582,N_21566);
or U21852 (N_21852,N_21533,N_21709);
or U21853 (N_21853,N_21573,N_21519);
nand U21854 (N_21854,N_21540,N_21603);
or U21855 (N_21855,N_21628,N_21692);
xnor U21856 (N_21856,N_21699,N_21625);
xnor U21857 (N_21857,N_21675,N_21648);
nand U21858 (N_21858,N_21591,N_21738);
and U21859 (N_21859,N_21595,N_21623);
xor U21860 (N_21860,N_21657,N_21621);
nand U21861 (N_21861,N_21676,N_21561);
and U21862 (N_21862,N_21549,N_21614);
nor U21863 (N_21863,N_21654,N_21735);
or U21864 (N_21864,N_21739,N_21687);
or U21865 (N_21865,N_21512,N_21524);
nand U21866 (N_21866,N_21644,N_21555);
nand U21867 (N_21867,N_21641,N_21535);
nand U21868 (N_21868,N_21602,N_21556);
or U21869 (N_21869,N_21506,N_21646);
nor U21870 (N_21870,N_21521,N_21579);
nor U21871 (N_21871,N_21637,N_21690);
xnor U21872 (N_21872,N_21608,N_21736);
nand U21873 (N_21873,N_21682,N_21671);
nand U21874 (N_21874,N_21715,N_21717);
xnor U21875 (N_21875,N_21587,N_21516);
xor U21876 (N_21876,N_21501,N_21595);
nand U21877 (N_21877,N_21627,N_21526);
nor U21878 (N_21878,N_21739,N_21649);
or U21879 (N_21879,N_21729,N_21585);
nor U21880 (N_21880,N_21616,N_21683);
nor U21881 (N_21881,N_21569,N_21699);
nor U21882 (N_21882,N_21553,N_21572);
nor U21883 (N_21883,N_21502,N_21742);
and U21884 (N_21884,N_21700,N_21630);
nand U21885 (N_21885,N_21643,N_21722);
xnor U21886 (N_21886,N_21696,N_21703);
nand U21887 (N_21887,N_21710,N_21566);
or U21888 (N_21888,N_21631,N_21687);
nand U21889 (N_21889,N_21628,N_21614);
nor U21890 (N_21890,N_21508,N_21611);
nand U21891 (N_21891,N_21612,N_21595);
and U21892 (N_21892,N_21733,N_21631);
nor U21893 (N_21893,N_21654,N_21596);
or U21894 (N_21894,N_21553,N_21576);
nand U21895 (N_21895,N_21638,N_21540);
nor U21896 (N_21896,N_21511,N_21646);
and U21897 (N_21897,N_21616,N_21703);
xnor U21898 (N_21898,N_21717,N_21536);
and U21899 (N_21899,N_21566,N_21507);
and U21900 (N_21900,N_21543,N_21534);
xor U21901 (N_21901,N_21551,N_21635);
nor U21902 (N_21902,N_21721,N_21500);
xnor U21903 (N_21903,N_21504,N_21717);
or U21904 (N_21904,N_21730,N_21646);
nand U21905 (N_21905,N_21636,N_21684);
nand U21906 (N_21906,N_21568,N_21501);
or U21907 (N_21907,N_21625,N_21714);
nor U21908 (N_21908,N_21650,N_21724);
or U21909 (N_21909,N_21685,N_21629);
nor U21910 (N_21910,N_21500,N_21723);
nor U21911 (N_21911,N_21691,N_21621);
nor U21912 (N_21912,N_21738,N_21544);
or U21913 (N_21913,N_21679,N_21535);
and U21914 (N_21914,N_21723,N_21720);
nand U21915 (N_21915,N_21699,N_21690);
nand U21916 (N_21916,N_21562,N_21516);
or U21917 (N_21917,N_21661,N_21601);
and U21918 (N_21918,N_21582,N_21737);
nand U21919 (N_21919,N_21601,N_21511);
and U21920 (N_21920,N_21659,N_21745);
nor U21921 (N_21921,N_21684,N_21580);
and U21922 (N_21922,N_21678,N_21662);
xor U21923 (N_21923,N_21626,N_21602);
and U21924 (N_21924,N_21682,N_21729);
and U21925 (N_21925,N_21622,N_21588);
nor U21926 (N_21926,N_21556,N_21591);
nor U21927 (N_21927,N_21632,N_21680);
nor U21928 (N_21928,N_21561,N_21572);
and U21929 (N_21929,N_21557,N_21573);
and U21930 (N_21930,N_21663,N_21529);
and U21931 (N_21931,N_21732,N_21744);
xnor U21932 (N_21932,N_21556,N_21555);
or U21933 (N_21933,N_21589,N_21549);
nor U21934 (N_21934,N_21743,N_21589);
nor U21935 (N_21935,N_21737,N_21675);
or U21936 (N_21936,N_21542,N_21698);
nor U21937 (N_21937,N_21619,N_21556);
and U21938 (N_21938,N_21575,N_21507);
nand U21939 (N_21939,N_21634,N_21529);
nor U21940 (N_21940,N_21537,N_21530);
nand U21941 (N_21941,N_21645,N_21703);
xor U21942 (N_21942,N_21605,N_21629);
and U21943 (N_21943,N_21510,N_21613);
xnor U21944 (N_21944,N_21536,N_21700);
xnor U21945 (N_21945,N_21606,N_21536);
or U21946 (N_21946,N_21749,N_21746);
or U21947 (N_21947,N_21543,N_21633);
or U21948 (N_21948,N_21530,N_21546);
nor U21949 (N_21949,N_21579,N_21690);
and U21950 (N_21950,N_21667,N_21736);
nor U21951 (N_21951,N_21738,N_21519);
and U21952 (N_21952,N_21597,N_21720);
and U21953 (N_21953,N_21664,N_21541);
or U21954 (N_21954,N_21700,N_21666);
or U21955 (N_21955,N_21715,N_21640);
and U21956 (N_21956,N_21690,N_21642);
xor U21957 (N_21957,N_21515,N_21678);
nand U21958 (N_21958,N_21508,N_21579);
and U21959 (N_21959,N_21545,N_21725);
xnor U21960 (N_21960,N_21583,N_21635);
nand U21961 (N_21961,N_21705,N_21653);
nand U21962 (N_21962,N_21546,N_21643);
and U21963 (N_21963,N_21560,N_21733);
nor U21964 (N_21964,N_21674,N_21553);
xor U21965 (N_21965,N_21586,N_21567);
xor U21966 (N_21966,N_21638,N_21506);
xnor U21967 (N_21967,N_21552,N_21621);
xnor U21968 (N_21968,N_21633,N_21749);
nor U21969 (N_21969,N_21642,N_21596);
nand U21970 (N_21970,N_21744,N_21549);
and U21971 (N_21971,N_21731,N_21543);
and U21972 (N_21972,N_21525,N_21743);
nor U21973 (N_21973,N_21587,N_21503);
or U21974 (N_21974,N_21691,N_21587);
nand U21975 (N_21975,N_21596,N_21603);
or U21976 (N_21976,N_21528,N_21581);
nand U21977 (N_21977,N_21740,N_21645);
nand U21978 (N_21978,N_21512,N_21581);
xnor U21979 (N_21979,N_21746,N_21639);
nand U21980 (N_21980,N_21710,N_21627);
and U21981 (N_21981,N_21564,N_21570);
or U21982 (N_21982,N_21652,N_21507);
xor U21983 (N_21983,N_21601,N_21703);
nand U21984 (N_21984,N_21663,N_21729);
nand U21985 (N_21985,N_21523,N_21612);
nor U21986 (N_21986,N_21574,N_21525);
xnor U21987 (N_21987,N_21505,N_21578);
or U21988 (N_21988,N_21666,N_21641);
or U21989 (N_21989,N_21593,N_21609);
nand U21990 (N_21990,N_21655,N_21665);
nand U21991 (N_21991,N_21713,N_21583);
or U21992 (N_21992,N_21554,N_21593);
nor U21993 (N_21993,N_21529,N_21657);
nand U21994 (N_21994,N_21709,N_21598);
xnor U21995 (N_21995,N_21625,N_21747);
nand U21996 (N_21996,N_21721,N_21534);
nor U21997 (N_21997,N_21726,N_21535);
nor U21998 (N_21998,N_21688,N_21633);
nand U21999 (N_21999,N_21582,N_21630);
nand U22000 (N_22000,N_21911,N_21890);
nand U22001 (N_22001,N_21830,N_21752);
xnor U22002 (N_22002,N_21802,N_21902);
and U22003 (N_22003,N_21788,N_21797);
xor U22004 (N_22004,N_21773,N_21759);
and U22005 (N_22005,N_21762,N_21825);
nand U22006 (N_22006,N_21796,N_21843);
and U22007 (N_22007,N_21756,N_21882);
or U22008 (N_22008,N_21828,N_21850);
and U22009 (N_22009,N_21760,N_21963);
xnor U22010 (N_22010,N_21897,N_21959);
and U22011 (N_22011,N_21981,N_21844);
nand U22012 (N_22012,N_21889,N_21763);
and U22013 (N_22013,N_21879,N_21861);
xor U22014 (N_22014,N_21811,N_21854);
and U22015 (N_22015,N_21877,N_21753);
or U22016 (N_22016,N_21833,N_21823);
nand U22017 (N_22017,N_21853,N_21804);
and U22018 (N_22018,N_21961,N_21829);
or U22019 (N_22019,N_21956,N_21966);
nor U22020 (N_22020,N_21867,N_21940);
or U22021 (N_22021,N_21881,N_21952);
and U22022 (N_22022,N_21781,N_21815);
and U22023 (N_22023,N_21962,N_21942);
xnor U22024 (N_22024,N_21974,N_21915);
or U22025 (N_22025,N_21986,N_21921);
nor U22026 (N_22026,N_21934,N_21895);
and U22027 (N_22027,N_21842,N_21775);
and U22028 (N_22028,N_21872,N_21798);
or U22029 (N_22029,N_21978,N_21973);
and U22030 (N_22030,N_21967,N_21770);
xnor U22031 (N_22031,N_21880,N_21808);
nand U22032 (N_22032,N_21780,N_21987);
nand U22033 (N_22033,N_21793,N_21864);
xnor U22034 (N_22034,N_21943,N_21886);
and U22035 (N_22035,N_21923,N_21900);
xor U22036 (N_22036,N_21779,N_21898);
nand U22037 (N_22037,N_21824,N_21896);
xnor U22038 (N_22038,N_21863,N_21977);
and U22039 (N_22039,N_21751,N_21789);
nand U22040 (N_22040,N_21904,N_21771);
nand U22041 (N_22041,N_21992,N_21972);
and U22042 (N_22042,N_21946,N_21822);
nand U22043 (N_22043,N_21918,N_21805);
xnor U22044 (N_22044,N_21891,N_21883);
or U22045 (N_22045,N_21807,N_21758);
xnor U22046 (N_22046,N_21985,N_21976);
nand U22047 (N_22047,N_21795,N_21984);
xor U22048 (N_22048,N_21869,N_21785);
xnor U22049 (N_22049,N_21866,N_21903);
and U22050 (N_22050,N_21953,N_21970);
and U22051 (N_22051,N_21839,N_21764);
nor U22052 (N_22052,N_21859,N_21841);
or U22053 (N_22053,N_21884,N_21988);
and U22054 (N_22054,N_21768,N_21913);
or U22055 (N_22055,N_21906,N_21993);
and U22056 (N_22056,N_21831,N_21887);
and U22057 (N_22057,N_21784,N_21874);
nor U22058 (N_22058,N_21865,N_21893);
nor U22059 (N_22059,N_21772,N_21858);
or U22060 (N_22060,N_21997,N_21980);
and U22061 (N_22061,N_21821,N_21856);
nor U22062 (N_22062,N_21927,N_21885);
or U22063 (N_22063,N_21778,N_21838);
and U22064 (N_22064,N_21782,N_21806);
or U22065 (N_22065,N_21814,N_21929);
or U22066 (N_22066,N_21991,N_21870);
and U22067 (N_22067,N_21937,N_21965);
or U22068 (N_22068,N_21916,N_21932);
or U22069 (N_22069,N_21791,N_21907);
nand U22070 (N_22070,N_21928,N_21765);
or U22071 (N_22071,N_21871,N_21809);
nand U22072 (N_22072,N_21888,N_21941);
nand U22073 (N_22073,N_21855,N_21910);
or U22074 (N_22074,N_21998,N_21920);
or U22075 (N_22075,N_21801,N_21938);
nand U22076 (N_22076,N_21786,N_21755);
nor U22077 (N_22077,N_21933,N_21852);
xor U22078 (N_22078,N_21919,N_21945);
xor U22079 (N_22079,N_21996,N_21944);
nor U22080 (N_22080,N_21847,N_21792);
nand U22081 (N_22081,N_21969,N_21794);
nor U22082 (N_22082,N_21769,N_21878);
nand U22083 (N_22083,N_21766,N_21924);
nor U22084 (N_22084,N_21813,N_21826);
nor U22085 (N_22085,N_21957,N_21818);
nor U22086 (N_22086,N_21892,N_21857);
xor U22087 (N_22087,N_21812,N_21774);
nand U22088 (N_22088,N_21840,N_21964);
or U22089 (N_22089,N_21832,N_21955);
or U22090 (N_22090,N_21909,N_21799);
xor U22091 (N_22091,N_21800,N_21926);
and U22092 (N_22092,N_21950,N_21876);
or U22093 (N_22093,N_21757,N_21954);
or U22094 (N_22094,N_21936,N_21922);
nor U22095 (N_22095,N_21894,N_21776);
xor U22096 (N_22096,N_21949,N_21851);
and U22097 (N_22097,N_21914,N_21837);
nand U22098 (N_22098,N_21960,N_21817);
and U22099 (N_22099,N_21925,N_21931);
or U22100 (N_22100,N_21860,N_21948);
nand U22101 (N_22101,N_21819,N_21787);
xnor U22102 (N_22102,N_21994,N_21803);
nand U22103 (N_22103,N_21836,N_21846);
and U22104 (N_22104,N_21777,N_21834);
nand U22105 (N_22105,N_21990,N_21971);
xor U22106 (N_22106,N_21947,N_21754);
xnor U22107 (N_22107,N_21875,N_21982);
nand U22108 (N_22108,N_21899,N_21979);
nor U22109 (N_22109,N_21939,N_21848);
and U22110 (N_22110,N_21958,N_21827);
nand U22111 (N_22111,N_21790,N_21983);
nor U22112 (N_22112,N_21868,N_21750);
nand U22113 (N_22113,N_21761,N_21862);
nor U22114 (N_22114,N_21917,N_21901);
and U22115 (N_22115,N_21935,N_21912);
and U22116 (N_22116,N_21905,N_21767);
xor U22117 (N_22117,N_21816,N_21995);
or U22118 (N_22118,N_21908,N_21989);
nor U22119 (N_22119,N_21873,N_21783);
xnor U22120 (N_22120,N_21975,N_21951);
xnor U22121 (N_22121,N_21930,N_21968);
or U22122 (N_22122,N_21999,N_21849);
xor U22123 (N_22123,N_21845,N_21835);
xor U22124 (N_22124,N_21820,N_21810);
xnor U22125 (N_22125,N_21752,N_21777);
nor U22126 (N_22126,N_21751,N_21790);
and U22127 (N_22127,N_21794,N_21980);
nand U22128 (N_22128,N_21793,N_21874);
nor U22129 (N_22129,N_21839,N_21825);
xnor U22130 (N_22130,N_21964,N_21923);
nor U22131 (N_22131,N_21962,N_21895);
and U22132 (N_22132,N_21978,N_21805);
xor U22133 (N_22133,N_21826,N_21831);
nor U22134 (N_22134,N_21966,N_21929);
nand U22135 (N_22135,N_21823,N_21871);
xnor U22136 (N_22136,N_21918,N_21833);
nand U22137 (N_22137,N_21883,N_21827);
xor U22138 (N_22138,N_21895,N_21754);
nor U22139 (N_22139,N_21844,N_21993);
nor U22140 (N_22140,N_21933,N_21758);
nor U22141 (N_22141,N_21948,N_21859);
or U22142 (N_22142,N_21887,N_21983);
and U22143 (N_22143,N_21779,N_21996);
and U22144 (N_22144,N_21890,N_21882);
nand U22145 (N_22145,N_21825,N_21903);
xor U22146 (N_22146,N_21908,N_21837);
xnor U22147 (N_22147,N_21779,N_21884);
nor U22148 (N_22148,N_21934,N_21873);
xor U22149 (N_22149,N_21947,N_21931);
nor U22150 (N_22150,N_21854,N_21796);
nand U22151 (N_22151,N_21763,N_21992);
or U22152 (N_22152,N_21887,N_21871);
nor U22153 (N_22153,N_21817,N_21836);
nand U22154 (N_22154,N_21822,N_21905);
and U22155 (N_22155,N_21954,N_21940);
or U22156 (N_22156,N_21986,N_21984);
xor U22157 (N_22157,N_21754,N_21878);
or U22158 (N_22158,N_21814,N_21816);
xor U22159 (N_22159,N_21865,N_21963);
nor U22160 (N_22160,N_21953,N_21817);
xor U22161 (N_22161,N_21757,N_21955);
xor U22162 (N_22162,N_21900,N_21973);
and U22163 (N_22163,N_21877,N_21882);
nor U22164 (N_22164,N_21979,N_21957);
and U22165 (N_22165,N_21954,N_21758);
nor U22166 (N_22166,N_21979,N_21976);
nor U22167 (N_22167,N_21796,N_21911);
xor U22168 (N_22168,N_21815,N_21863);
nand U22169 (N_22169,N_21769,N_21941);
and U22170 (N_22170,N_21817,N_21840);
and U22171 (N_22171,N_21993,N_21953);
xnor U22172 (N_22172,N_21891,N_21983);
nor U22173 (N_22173,N_21858,N_21782);
or U22174 (N_22174,N_21867,N_21948);
or U22175 (N_22175,N_21834,N_21892);
nor U22176 (N_22176,N_21843,N_21853);
xnor U22177 (N_22177,N_21796,N_21984);
or U22178 (N_22178,N_21751,N_21763);
and U22179 (N_22179,N_21772,N_21887);
and U22180 (N_22180,N_21869,N_21994);
nor U22181 (N_22181,N_21958,N_21964);
xnor U22182 (N_22182,N_21767,N_21962);
nor U22183 (N_22183,N_21805,N_21881);
and U22184 (N_22184,N_21767,N_21781);
and U22185 (N_22185,N_21753,N_21820);
nand U22186 (N_22186,N_21969,N_21859);
nor U22187 (N_22187,N_21876,N_21999);
and U22188 (N_22188,N_21900,N_21848);
xor U22189 (N_22189,N_21760,N_21857);
nor U22190 (N_22190,N_21753,N_21857);
nand U22191 (N_22191,N_21851,N_21883);
and U22192 (N_22192,N_21946,N_21981);
nor U22193 (N_22193,N_21782,N_21908);
nand U22194 (N_22194,N_21772,N_21951);
nand U22195 (N_22195,N_21955,N_21787);
or U22196 (N_22196,N_21893,N_21986);
nand U22197 (N_22197,N_21908,N_21890);
nand U22198 (N_22198,N_21994,N_21907);
or U22199 (N_22199,N_21848,N_21905);
and U22200 (N_22200,N_21787,N_21786);
xor U22201 (N_22201,N_21970,N_21880);
nor U22202 (N_22202,N_21954,N_21926);
nand U22203 (N_22203,N_21965,N_21813);
and U22204 (N_22204,N_21768,N_21785);
and U22205 (N_22205,N_21921,N_21856);
nor U22206 (N_22206,N_21959,N_21965);
nor U22207 (N_22207,N_21876,N_21966);
nand U22208 (N_22208,N_21824,N_21966);
nand U22209 (N_22209,N_21907,N_21996);
nor U22210 (N_22210,N_21760,N_21821);
or U22211 (N_22211,N_21766,N_21976);
or U22212 (N_22212,N_21767,N_21780);
and U22213 (N_22213,N_21778,N_21913);
xor U22214 (N_22214,N_21967,N_21847);
nor U22215 (N_22215,N_21838,N_21984);
or U22216 (N_22216,N_21974,N_21928);
nand U22217 (N_22217,N_21781,N_21777);
and U22218 (N_22218,N_21840,N_21801);
xnor U22219 (N_22219,N_21959,N_21860);
or U22220 (N_22220,N_21873,N_21807);
xnor U22221 (N_22221,N_21923,N_21788);
or U22222 (N_22222,N_21751,N_21797);
nand U22223 (N_22223,N_21779,N_21797);
or U22224 (N_22224,N_21822,N_21976);
nor U22225 (N_22225,N_21993,N_21760);
nor U22226 (N_22226,N_21873,N_21819);
and U22227 (N_22227,N_21876,N_21942);
or U22228 (N_22228,N_21938,N_21955);
nor U22229 (N_22229,N_21815,N_21867);
xnor U22230 (N_22230,N_21815,N_21940);
or U22231 (N_22231,N_21768,N_21841);
xor U22232 (N_22232,N_21851,N_21857);
or U22233 (N_22233,N_21898,N_21949);
nand U22234 (N_22234,N_21760,N_21813);
nand U22235 (N_22235,N_21971,N_21781);
nand U22236 (N_22236,N_21752,N_21935);
nor U22237 (N_22237,N_21856,N_21756);
nor U22238 (N_22238,N_21773,N_21993);
and U22239 (N_22239,N_21898,N_21927);
or U22240 (N_22240,N_21900,N_21857);
nor U22241 (N_22241,N_21786,N_21993);
xnor U22242 (N_22242,N_21770,N_21942);
xor U22243 (N_22243,N_21818,N_21941);
nor U22244 (N_22244,N_21922,N_21955);
or U22245 (N_22245,N_21775,N_21828);
nor U22246 (N_22246,N_21963,N_21855);
and U22247 (N_22247,N_21827,N_21840);
or U22248 (N_22248,N_21803,N_21909);
nor U22249 (N_22249,N_21789,N_21951);
and U22250 (N_22250,N_22032,N_22197);
and U22251 (N_22251,N_22077,N_22171);
nand U22252 (N_22252,N_22190,N_22206);
or U22253 (N_22253,N_22041,N_22039);
or U22254 (N_22254,N_22006,N_22212);
nand U22255 (N_22255,N_22135,N_22043);
or U22256 (N_22256,N_22137,N_22122);
nand U22257 (N_22257,N_22031,N_22113);
or U22258 (N_22258,N_22040,N_22184);
nand U22259 (N_22259,N_22233,N_22241);
or U22260 (N_22260,N_22011,N_22195);
or U22261 (N_22261,N_22243,N_22239);
or U22262 (N_22262,N_22221,N_22214);
or U22263 (N_22263,N_22194,N_22024);
nand U22264 (N_22264,N_22164,N_22125);
or U22265 (N_22265,N_22019,N_22035);
or U22266 (N_22266,N_22045,N_22231);
and U22267 (N_22267,N_22152,N_22102);
nor U22268 (N_22268,N_22225,N_22021);
and U22269 (N_22269,N_22193,N_22051);
xor U22270 (N_22270,N_22063,N_22103);
nand U22271 (N_22271,N_22201,N_22093);
xnor U22272 (N_22272,N_22244,N_22100);
or U22273 (N_22273,N_22128,N_22007);
nor U22274 (N_22274,N_22081,N_22215);
or U22275 (N_22275,N_22245,N_22058);
xor U22276 (N_22276,N_22151,N_22166);
nor U22277 (N_22277,N_22027,N_22157);
xnor U22278 (N_22278,N_22115,N_22065);
and U22279 (N_22279,N_22029,N_22238);
and U22280 (N_22280,N_22232,N_22119);
nand U22281 (N_22281,N_22175,N_22216);
and U22282 (N_22282,N_22139,N_22108);
or U22283 (N_22283,N_22237,N_22052);
nor U22284 (N_22284,N_22138,N_22106);
nand U22285 (N_22285,N_22089,N_22114);
or U22286 (N_22286,N_22149,N_22023);
nor U22287 (N_22287,N_22014,N_22046);
xor U22288 (N_22288,N_22004,N_22121);
and U22289 (N_22289,N_22200,N_22158);
and U22290 (N_22290,N_22042,N_22161);
or U22291 (N_22291,N_22159,N_22144);
and U22292 (N_22292,N_22112,N_22069);
xnor U22293 (N_22293,N_22094,N_22169);
xnor U22294 (N_22294,N_22246,N_22016);
nor U22295 (N_22295,N_22129,N_22111);
and U22296 (N_22296,N_22165,N_22049);
nand U22297 (N_22297,N_22204,N_22179);
and U22298 (N_22298,N_22229,N_22018);
xor U22299 (N_22299,N_22222,N_22067);
or U22300 (N_22300,N_22101,N_22181);
xor U22301 (N_22301,N_22022,N_22209);
and U22302 (N_22302,N_22168,N_22236);
xor U22303 (N_22303,N_22226,N_22198);
xnor U22304 (N_22304,N_22078,N_22061);
nand U22305 (N_22305,N_22010,N_22187);
or U22306 (N_22306,N_22249,N_22053);
xnor U22307 (N_22307,N_22047,N_22116);
nor U22308 (N_22308,N_22180,N_22132);
or U22309 (N_22309,N_22118,N_22167);
or U22310 (N_22310,N_22154,N_22025);
or U22311 (N_22311,N_22177,N_22015);
xor U22312 (N_22312,N_22070,N_22117);
or U22313 (N_22313,N_22218,N_22079);
xor U22314 (N_22314,N_22202,N_22134);
xnor U22315 (N_22315,N_22033,N_22148);
xnor U22316 (N_22316,N_22009,N_22105);
nand U22317 (N_22317,N_22013,N_22219);
nand U22318 (N_22318,N_22203,N_22127);
xnor U22319 (N_22319,N_22182,N_22211);
nor U22320 (N_22320,N_22110,N_22005);
and U22321 (N_22321,N_22228,N_22248);
nand U22322 (N_22322,N_22068,N_22247);
and U22323 (N_22323,N_22082,N_22059);
nand U22324 (N_22324,N_22207,N_22172);
and U22325 (N_22325,N_22131,N_22140);
or U22326 (N_22326,N_22191,N_22235);
nand U22327 (N_22327,N_22062,N_22044);
xnor U22328 (N_22328,N_22099,N_22150);
and U22329 (N_22329,N_22186,N_22143);
and U22330 (N_22330,N_22220,N_22230);
xnor U22331 (N_22331,N_22086,N_22003);
or U22332 (N_22332,N_22037,N_22170);
nand U22333 (N_22333,N_22012,N_22060);
nand U22334 (N_22334,N_22088,N_22073);
or U22335 (N_22335,N_22087,N_22071);
and U22336 (N_22336,N_22185,N_22133);
nand U22337 (N_22337,N_22155,N_22036);
xor U22338 (N_22338,N_22174,N_22120);
nand U22339 (N_22339,N_22050,N_22028);
nand U22340 (N_22340,N_22160,N_22098);
or U22341 (N_22341,N_22092,N_22156);
and U22342 (N_22342,N_22130,N_22224);
nor U22343 (N_22343,N_22026,N_22142);
nand U22344 (N_22344,N_22146,N_22208);
nor U22345 (N_22345,N_22038,N_22242);
xor U22346 (N_22346,N_22083,N_22104);
xor U22347 (N_22347,N_22107,N_22123);
nand U22348 (N_22348,N_22176,N_22136);
or U22349 (N_22349,N_22085,N_22192);
and U22350 (N_22350,N_22126,N_22227);
xor U22351 (N_22351,N_22001,N_22223);
xnor U22352 (N_22352,N_22057,N_22189);
xnor U22353 (N_22353,N_22124,N_22183);
nor U22354 (N_22354,N_22199,N_22210);
nor U22355 (N_22355,N_22234,N_22020);
xnor U22356 (N_22356,N_22091,N_22141);
nand U22357 (N_22357,N_22178,N_22188);
and U22358 (N_22358,N_22056,N_22066);
and U22359 (N_22359,N_22196,N_22084);
nor U22360 (N_22360,N_22034,N_22002);
or U22361 (N_22361,N_22008,N_22055);
or U22362 (N_22362,N_22090,N_22072);
xor U22363 (N_22363,N_22109,N_22163);
or U22364 (N_22364,N_22017,N_22000);
and U22365 (N_22365,N_22095,N_22076);
nand U22366 (N_22366,N_22173,N_22075);
nand U22367 (N_22367,N_22097,N_22080);
nor U22368 (N_22368,N_22217,N_22162);
nand U22369 (N_22369,N_22213,N_22153);
xnor U22370 (N_22370,N_22240,N_22064);
and U22371 (N_22371,N_22074,N_22030);
nor U22372 (N_22372,N_22145,N_22205);
or U22373 (N_22373,N_22048,N_22096);
nor U22374 (N_22374,N_22147,N_22054);
or U22375 (N_22375,N_22243,N_22035);
and U22376 (N_22376,N_22069,N_22036);
and U22377 (N_22377,N_22230,N_22126);
and U22378 (N_22378,N_22174,N_22071);
xor U22379 (N_22379,N_22130,N_22017);
or U22380 (N_22380,N_22157,N_22052);
xnor U22381 (N_22381,N_22062,N_22039);
nor U22382 (N_22382,N_22061,N_22130);
and U22383 (N_22383,N_22006,N_22196);
or U22384 (N_22384,N_22166,N_22038);
nor U22385 (N_22385,N_22108,N_22047);
nand U22386 (N_22386,N_22071,N_22090);
and U22387 (N_22387,N_22208,N_22042);
or U22388 (N_22388,N_22105,N_22029);
and U22389 (N_22389,N_22048,N_22202);
nand U22390 (N_22390,N_22194,N_22191);
and U22391 (N_22391,N_22036,N_22095);
nand U22392 (N_22392,N_22233,N_22042);
nor U22393 (N_22393,N_22156,N_22010);
or U22394 (N_22394,N_22012,N_22057);
nor U22395 (N_22395,N_22171,N_22076);
and U22396 (N_22396,N_22162,N_22019);
and U22397 (N_22397,N_22144,N_22184);
nand U22398 (N_22398,N_22055,N_22024);
or U22399 (N_22399,N_22203,N_22117);
and U22400 (N_22400,N_22168,N_22004);
xor U22401 (N_22401,N_22230,N_22171);
xor U22402 (N_22402,N_22231,N_22092);
nand U22403 (N_22403,N_22220,N_22158);
or U22404 (N_22404,N_22238,N_22103);
xnor U22405 (N_22405,N_22014,N_22128);
or U22406 (N_22406,N_22135,N_22085);
nor U22407 (N_22407,N_22055,N_22081);
or U22408 (N_22408,N_22122,N_22078);
xnor U22409 (N_22409,N_22182,N_22147);
nor U22410 (N_22410,N_22151,N_22080);
nand U22411 (N_22411,N_22096,N_22210);
nor U22412 (N_22412,N_22021,N_22237);
nand U22413 (N_22413,N_22217,N_22082);
and U22414 (N_22414,N_22157,N_22215);
nor U22415 (N_22415,N_22112,N_22149);
nor U22416 (N_22416,N_22161,N_22008);
xor U22417 (N_22417,N_22114,N_22123);
or U22418 (N_22418,N_22135,N_22230);
or U22419 (N_22419,N_22031,N_22003);
xnor U22420 (N_22420,N_22203,N_22144);
or U22421 (N_22421,N_22103,N_22015);
nand U22422 (N_22422,N_22140,N_22077);
xnor U22423 (N_22423,N_22243,N_22111);
nor U22424 (N_22424,N_22191,N_22068);
xnor U22425 (N_22425,N_22064,N_22202);
and U22426 (N_22426,N_22195,N_22074);
nor U22427 (N_22427,N_22001,N_22170);
xnor U22428 (N_22428,N_22055,N_22089);
nand U22429 (N_22429,N_22148,N_22125);
nor U22430 (N_22430,N_22203,N_22189);
nor U22431 (N_22431,N_22062,N_22242);
nor U22432 (N_22432,N_22111,N_22092);
nand U22433 (N_22433,N_22229,N_22063);
or U22434 (N_22434,N_22034,N_22056);
xor U22435 (N_22435,N_22083,N_22036);
nor U22436 (N_22436,N_22050,N_22042);
nand U22437 (N_22437,N_22072,N_22133);
or U22438 (N_22438,N_22185,N_22211);
xor U22439 (N_22439,N_22114,N_22040);
or U22440 (N_22440,N_22175,N_22078);
and U22441 (N_22441,N_22122,N_22038);
xnor U22442 (N_22442,N_22016,N_22221);
or U22443 (N_22443,N_22100,N_22205);
or U22444 (N_22444,N_22076,N_22098);
nor U22445 (N_22445,N_22071,N_22155);
nand U22446 (N_22446,N_22044,N_22028);
nand U22447 (N_22447,N_22191,N_22121);
nand U22448 (N_22448,N_22006,N_22157);
xor U22449 (N_22449,N_22244,N_22246);
xnor U22450 (N_22450,N_22216,N_22032);
or U22451 (N_22451,N_22019,N_22219);
xnor U22452 (N_22452,N_22014,N_22067);
nor U22453 (N_22453,N_22111,N_22203);
or U22454 (N_22454,N_22195,N_22003);
and U22455 (N_22455,N_22208,N_22099);
or U22456 (N_22456,N_22167,N_22179);
nor U22457 (N_22457,N_22049,N_22106);
nand U22458 (N_22458,N_22222,N_22247);
or U22459 (N_22459,N_22011,N_22129);
or U22460 (N_22460,N_22036,N_22013);
or U22461 (N_22461,N_22013,N_22103);
and U22462 (N_22462,N_22006,N_22056);
nor U22463 (N_22463,N_22134,N_22157);
or U22464 (N_22464,N_22054,N_22215);
or U22465 (N_22465,N_22109,N_22158);
nor U22466 (N_22466,N_22036,N_22133);
or U22467 (N_22467,N_22062,N_22149);
and U22468 (N_22468,N_22057,N_22004);
nand U22469 (N_22469,N_22177,N_22006);
or U22470 (N_22470,N_22197,N_22104);
nor U22471 (N_22471,N_22045,N_22112);
xnor U22472 (N_22472,N_22234,N_22157);
or U22473 (N_22473,N_22020,N_22162);
nand U22474 (N_22474,N_22201,N_22038);
and U22475 (N_22475,N_22009,N_22046);
nor U22476 (N_22476,N_22237,N_22228);
nor U22477 (N_22477,N_22065,N_22205);
nand U22478 (N_22478,N_22080,N_22202);
and U22479 (N_22479,N_22197,N_22145);
xor U22480 (N_22480,N_22092,N_22165);
xnor U22481 (N_22481,N_22104,N_22169);
xnor U22482 (N_22482,N_22217,N_22008);
xor U22483 (N_22483,N_22129,N_22197);
or U22484 (N_22484,N_22008,N_22223);
xor U22485 (N_22485,N_22170,N_22028);
or U22486 (N_22486,N_22105,N_22034);
nor U22487 (N_22487,N_22105,N_22088);
nand U22488 (N_22488,N_22142,N_22089);
xnor U22489 (N_22489,N_22074,N_22044);
or U22490 (N_22490,N_22196,N_22177);
or U22491 (N_22491,N_22087,N_22025);
nand U22492 (N_22492,N_22182,N_22197);
or U22493 (N_22493,N_22141,N_22209);
nor U22494 (N_22494,N_22102,N_22040);
or U22495 (N_22495,N_22207,N_22063);
and U22496 (N_22496,N_22200,N_22103);
xnor U22497 (N_22497,N_22171,N_22084);
and U22498 (N_22498,N_22014,N_22114);
or U22499 (N_22499,N_22117,N_22174);
and U22500 (N_22500,N_22392,N_22303);
xnor U22501 (N_22501,N_22262,N_22456);
nand U22502 (N_22502,N_22374,N_22423);
nand U22503 (N_22503,N_22292,N_22445);
xnor U22504 (N_22504,N_22294,N_22282);
or U22505 (N_22505,N_22307,N_22454);
xor U22506 (N_22506,N_22330,N_22408);
or U22507 (N_22507,N_22404,N_22452);
nor U22508 (N_22508,N_22337,N_22470);
xnor U22509 (N_22509,N_22293,N_22482);
or U22510 (N_22510,N_22467,N_22288);
nand U22511 (N_22511,N_22377,N_22365);
xor U22512 (N_22512,N_22356,N_22491);
nand U22513 (N_22513,N_22462,N_22298);
or U22514 (N_22514,N_22443,N_22492);
nand U22515 (N_22515,N_22353,N_22384);
and U22516 (N_22516,N_22264,N_22306);
or U22517 (N_22517,N_22344,N_22426);
nor U22518 (N_22518,N_22484,N_22327);
nand U22519 (N_22519,N_22350,N_22386);
and U22520 (N_22520,N_22419,N_22322);
xnor U22521 (N_22521,N_22255,N_22253);
nor U22522 (N_22522,N_22376,N_22336);
nor U22523 (N_22523,N_22433,N_22441);
xnor U22524 (N_22524,N_22463,N_22265);
nor U22525 (N_22525,N_22279,N_22358);
xnor U22526 (N_22526,N_22457,N_22477);
xnor U22527 (N_22527,N_22289,N_22304);
xor U22528 (N_22528,N_22494,N_22390);
xor U22529 (N_22529,N_22449,N_22340);
xor U22530 (N_22530,N_22461,N_22260);
or U22531 (N_22531,N_22319,N_22295);
xnor U22532 (N_22532,N_22422,N_22311);
and U22533 (N_22533,N_22285,N_22431);
nand U22534 (N_22534,N_22308,N_22355);
or U22535 (N_22535,N_22272,N_22380);
and U22536 (N_22536,N_22345,N_22455);
or U22537 (N_22537,N_22401,N_22284);
and U22538 (N_22538,N_22414,N_22420);
or U22539 (N_22539,N_22476,N_22465);
xnor U22540 (N_22540,N_22393,N_22447);
or U22541 (N_22541,N_22438,N_22363);
and U22542 (N_22542,N_22347,N_22409);
nor U22543 (N_22543,N_22479,N_22261);
nand U22544 (N_22544,N_22378,N_22486);
nand U22545 (N_22545,N_22362,N_22370);
and U22546 (N_22546,N_22357,N_22267);
or U22547 (N_22547,N_22475,N_22399);
and U22548 (N_22548,N_22341,N_22446);
or U22549 (N_22549,N_22373,N_22417);
nand U22550 (N_22550,N_22435,N_22381);
xor U22551 (N_22551,N_22371,N_22348);
nor U22552 (N_22552,N_22418,N_22442);
or U22553 (N_22553,N_22466,N_22331);
nor U22554 (N_22554,N_22312,N_22360);
xnor U22555 (N_22555,N_22405,N_22413);
or U22556 (N_22556,N_22459,N_22281);
or U22557 (N_22557,N_22391,N_22329);
nand U22558 (N_22558,N_22316,N_22259);
or U22559 (N_22559,N_22334,N_22415);
and U22560 (N_22560,N_22480,N_22489);
nand U22561 (N_22561,N_22254,N_22437);
nand U22562 (N_22562,N_22300,N_22483);
and U22563 (N_22563,N_22495,N_22323);
xor U22564 (N_22564,N_22448,N_22487);
xor U22565 (N_22565,N_22273,N_22296);
nand U22566 (N_22566,N_22352,N_22263);
xor U22567 (N_22567,N_22369,N_22382);
xor U22568 (N_22568,N_22326,N_22324);
nand U22569 (N_22569,N_22388,N_22299);
and U22570 (N_22570,N_22297,N_22460);
or U22571 (N_22571,N_22314,N_22497);
nor U22572 (N_22572,N_22379,N_22302);
and U22573 (N_22573,N_22343,N_22412);
nor U22574 (N_22574,N_22440,N_22389);
nor U22575 (N_22575,N_22338,N_22256);
nand U22576 (N_22576,N_22471,N_22498);
nor U22577 (N_22577,N_22428,N_22411);
xnor U22578 (N_22578,N_22367,N_22481);
or U22579 (N_22579,N_22478,N_22383);
nor U22580 (N_22580,N_22269,N_22398);
or U22581 (N_22581,N_22372,N_22385);
nand U22582 (N_22582,N_22328,N_22429);
and U22583 (N_22583,N_22280,N_22351);
nand U22584 (N_22584,N_22375,N_22349);
and U22585 (N_22585,N_22325,N_22290);
and U22586 (N_22586,N_22335,N_22275);
nor U22587 (N_22587,N_22286,N_22439);
nor U22588 (N_22588,N_22317,N_22276);
or U22589 (N_22589,N_22301,N_22485);
nor U22590 (N_22590,N_22277,N_22251);
xnor U22591 (N_22591,N_22468,N_22472);
xor U22592 (N_22592,N_22287,N_22313);
or U22593 (N_22593,N_22458,N_22396);
or U22594 (N_22594,N_22430,N_22421);
nand U22595 (N_22595,N_22271,N_22250);
xnor U22596 (N_22596,N_22333,N_22283);
nor U22597 (N_22597,N_22451,N_22403);
nand U22598 (N_22598,N_22270,N_22278);
nor U22599 (N_22599,N_22305,N_22346);
nand U22600 (N_22600,N_22368,N_22496);
nand U22601 (N_22601,N_22499,N_22444);
nor U22602 (N_22602,N_22394,N_22424);
and U22603 (N_22603,N_22252,N_22274);
and U22604 (N_22604,N_22310,N_22436);
or U22605 (N_22605,N_22473,N_22397);
or U22606 (N_22606,N_22400,N_22320);
nand U22607 (N_22607,N_22425,N_22410);
nand U22608 (N_22608,N_22464,N_22321);
or U22609 (N_22609,N_22332,N_22387);
or U22610 (N_22610,N_22315,N_22257);
xnor U22611 (N_22611,N_22469,N_22366);
nand U22612 (N_22612,N_22406,N_22395);
or U22613 (N_22613,N_22342,N_22416);
and U22614 (N_22614,N_22258,N_22339);
and U22615 (N_22615,N_22407,N_22432);
and U22616 (N_22616,N_22453,N_22309);
or U22617 (N_22617,N_22474,N_22354);
or U22618 (N_22618,N_22427,N_22450);
nand U22619 (N_22619,N_22434,N_22318);
nand U22620 (N_22620,N_22268,N_22490);
and U22621 (N_22621,N_22266,N_22493);
nand U22622 (N_22622,N_22488,N_22361);
or U22623 (N_22623,N_22364,N_22402);
or U22624 (N_22624,N_22291,N_22359);
nand U22625 (N_22625,N_22451,N_22412);
xnor U22626 (N_22626,N_22421,N_22397);
nor U22627 (N_22627,N_22362,N_22492);
xor U22628 (N_22628,N_22480,N_22342);
and U22629 (N_22629,N_22287,N_22432);
and U22630 (N_22630,N_22255,N_22424);
nor U22631 (N_22631,N_22413,N_22470);
and U22632 (N_22632,N_22322,N_22384);
nand U22633 (N_22633,N_22272,N_22409);
or U22634 (N_22634,N_22446,N_22329);
or U22635 (N_22635,N_22451,N_22380);
nand U22636 (N_22636,N_22295,N_22458);
nand U22637 (N_22637,N_22285,N_22287);
nand U22638 (N_22638,N_22324,N_22322);
nor U22639 (N_22639,N_22261,N_22384);
nand U22640 (N_22640,N_22281,N_22351);
or U22641 (N_22641,N_22299,N_22267);
and U22642 (N_22642,N_22299,N_22495);
and U22643 (N_22643,N_22357,N_22420);
and U22644 (N_22644,N_22473,N_22413);
and U22645 (N_22645,N_22433,N_22272);
nor U22646 (N_22646,N_22424,N_22381);
nand U22647 (N_22647,N_22327,N_22420);
or U22648 (N_22648,N_22372,N_22289);
nand U22649 (N_22649,N_22395,N_22498);
nor U22650 (N_22650,N_22326,N_22377);
nand U22651 (N_22651,N_22413,N_22293);
and U22652 (N_22652,N_22425,N_22339);
xnor U22653 (N_22653,N_22254,N_22316);
nor U22654 (N_22654,N_22446,N_22385);
and U22655 (N_22655,N_22458,N_22413);
xnor U22656 (N_22656,N_22325,N_22302);
xor U22657 (N_22657,N_22423,N_22266);
or U22658 (N_22658,N_22354,N_22417);
nand U22659 (N_22659,N_22418,N_22495);
nand U22660 (N_22660,N_22281,N_22395);
xor U22661 (N_22661,N_22434,N_22291);
and U22662 (N_22662,N_22435,N_22382);
nor U22663 (N_22663,N_22494,N_22460);
nand U22664 (N_22664,N_22297,N_22265);
nand U22665 (N_22665,N_22452,N_22259);
nand U22666 (N_22666,N_22376,N_22309);
xnor U22667 (N_22667,N_22372,N_22288);
xor U22668 (N_22668,N_22284,N_22463);
and U22669 (N_22669,N_22282,N_22356);
nand U22670 (N_22670,N_22303,N_22296);
nor U22671 (N_22671,N_22267,N_22416);
and U22672 (N_22672,N_22293,N_22271);
nand U22673 (N_22673,N_22292,N_22431);
nand U22674 (N_22674,N_22397,N_22444);
nand U22675 (N_22675,N_22396,N_22359);
xor U22676 (N_22676,N_22344,N_22491);
nand U22677 (N_22677,N_22457,N_22441);
and U22678 (N_22678,N_22469,N_22481);
or U22679 (N_22679,N_22433,N_22322);
xor U22680 (N_22680,N_22283,N_22264);
nor U22681 (N_22681,N_22426,N_22452);
nand U22682 (N_22682,N_22382,N_22419);
and U22683 (N_22683,N_22476,N_22305);
or U22684 (N_22684,N_22412,N_22480);
and U22685 (N_22685,N_22384,N_22368);
nand U22686 (N_22686,N_22433,N_22359);
or U22687 (N_22687,N_22298,N_22326);
xnor U22688 (N_22688,N_22380,N_22347);
xor U22689 (N_22689,N_22345,N_22276);
or U22690 (N_22690,N_22457,N_22305);
nor U22691 (N_22691,N_22258,N_22402);
nand U22692 (N_22692,N_22299,N_22319);
nand U22693 (N_22693,N_22419,N_22370);
or U22694 (N_22694,N_22312,N_22468);
xor U22695 (N_22695,N_22482,N_22415);
and U22696 (N_22696,N_22287,N_22414);
xnor U22697 (N_22697,N_22405,N_22488);
and U22698 (N_22698,N_22386,N_22453);
nor U22699 (N_22699,N_22475,N_22398);
or U22700 (N_22700,N_22387,N_22338);
or U22701 (N_22701,N_22365,N_22270);
or U22702 (N_22702,N_22487,N_22492);
xor U22703 (N_22703,N_22294,N_22398);
xnor U22704 (N_22704,N_22357,N_22262);
and U22705 (N_22705,N_22493,N_22407);
nand U22706 (N_22706,N_22371,N_22352);
xnor U22707 (N_22707,N_22417,N_22299);
xor U22708 (N_22708,N_22375,N_22466);
xnor U22709 (N_22709,N_22290,N_22420);
nand U22710 (N_22710,N_22433,N_22332);
nand U22711 (N_22711,N_22342,N_22368);
nand U22712 (N_22712,N_22471,N_22456);
nand U22713 (N_22713,N_22436,N_22322);
or U22714 (N_22714,N_22481,N_22383);
and U22715 (N_22715,N_22424,N_22375);
and U22716 (N_22716,N_22289,N_22470);
nand U22717 (N_22717,N_22304,N_22356);
and U22718 (N_22718,N_22392,N_22267);
xnor U22719 (N_22719,N_22377,N_22321);
xnor U22720 (N_22720,N_22497,N_22437);
xnor U22721 (N_22721,N_22434,N_22402);
xor U22722 (N_22722,N_22492,N_22454);
and U22723 (N_22723,N_22276,N_22339);
or U22724 (N_22724,N_22308,N_22262);
nand U22725 (N_22725,N_22407,N_22368);
nor U22726 (N_22726,N_22491,N_22403);
xnor U22727 (N_22727,N_22331,N_22374);
nor U22728 (N_22728,N_22455,N_22323);
nand U22729 (N_22729,N_22323,N_22429);
nand U22730 (N_22730,N_22407,N_22330);
and U22731 (N_22731,N_22327,N_22299);
nor U22732 (N_22732,N_22444,N_22269);
nor U22733 (N_22733,N_22323,N_22355);
and U22734 (N_22734,N_22477,N_22366);
nand U22735 (N_22735,N_22345,N_22295);
nor U22736 (N_22736,N_22319,N_22288);
xnor U22737 (N_22737,N_22286,N_22429);
xnor U22738 (N_22738,N_22445,N_22251);
nor U22739 (N_22739,N_22297,N_22252);
xnor U22740 (N_22740,N_22360,N_22460);
and U22741 (N_22741,N_22373,N_22370);
and U22742 (N_22742,N_22393,N_22256);
nor U22743 (N_22743,N_22425,N_22473);
or U22744 (N_22744,N_22484,N_22365);
xor U22745 (N_22745,N_22283,N_22455);
or U22746 (N_22746,N_22450,N_22322);
nor U22747 (N_22747,N_22313,N_22491);
nand U22748 (N_22748,N_22408,N_22309);
and U22749 (N_22749,N_22409,N_22474);
nand U22750 (N_22750,N_22583,N_22572);
or U22751 (N_22751,N_22587,N_22652);
and U22752 (N_22752,N_22631,N_22568);
xor U22753 (N_22753,N_22625,N_22501);
xor U22754 (N_22754,N_22681,N_22694);
or U22755 (N_22755,N_22669,N_22730);
xnor U22756 (N_22756,N_22748,N_22571);
nor U22757 (N_22757,N_22710,N_22645);
and U22758 (N_22758,N_22594,N_22584);
xor U22759 (N_22759,N_22680,N_22682);
or U22760 (N_22760,N_22524,N_22510);
nand U22761 (N_22761,N_22717,N_22707);
and U22762 (N_22762,N_22627,N_22527);
and U22763 (N_22763,N_22742,N_22693);
nor U22764 (N_22764,N_22605,N_22715);
nand U22765 (N_22765,N_22522,N_22678);
nor U22766 (N_22766,N_22606,N_22622);
xor U22767 (N_22767,N_22704,N_22667);
and U22768 (N_22768,N_22660,N_22567);
xor U22769 (N_22769,N_22604,N_22744);
xnor U22770 (N_22770,N_22609,N_22697);
nand U22771 (N_22771,N_22611,N_22502);
nand U22772 (N_22772,N_22560,N_22651);
and U22773 (N_22773,N_22559,N_22687);
nor U22774 (N_22774,N_22655,N_22732);
xnor U22775 (N_22775,N_22529,N_22671);
nand U22776 (N_22776,N_22500,N_22623);
or U22777 (N_22777,N_22614,N_22656);
nor U22778 (N_22778,N_22653,N_22679);
nor U22779 (N_22779,N_22506,N_22566);
nor U22780 (N_22780,N_22546,N_22558);
and U22781 (N_22781,N_22538,N_22722);
nand U22782 (N_22782,N_22716,N_22520);
or U22783 (N_22783,N_22507,N_22561);
nor U22784 (N_22784,N_22596,N_22737);
xor U22785 (N_22785,N_22613,N_22586);
xnor U22786 (N_22786,N_22509,N_22555);
and U22787 (N_22787,N_22602,N_22677);
nand U22788 (N_22788,N_22733,N_22521);
nor U22789 (N_22789,N_22731,N_22577);
and U22790 (N_22790,N_22540,N_22592);
and U22791 (N_22791,N_22570,N_22616);
nand U22792 (N_22792,N_22620,N_22535);
and U22793 (N_22793,N_22739,N_22600);
or U22794 (N_22794,N_22615,N_22564);
or U22795 (N_22795,N_22696,N_22557);
and U22796 (N_22796,N_22664,N_22593);
or U22797 (N_22797,N_22643,N_22536);
nor U22798 (N_22798,N_22741,N_22658);
xnor U22799 (N_22799,N_22565,N_22727);
nor U22800 (N_22800,N_22552,N_22576);
nand U22801 (N_22801,N_22612,N_22528);
xnor U22802 (N_22802,N_22665,N_22708);
nor U22803 (N_22803,N_22668,N_22513);
nand U22804 (N_22804,N_22673,N_22550);
or U22805 (N_22805,N_22738,N_22505);
or U22806 (N_22806,N_22712,N_22511);
or U22807 (N_22807,N_22698,N_22728);
nand U22808 (N_22808,N_22590,N_22688);
nand U22809 (N_22809,N_22661,N_22526);
or U22810 (N_22810,N_22556,N_22551);
or U22811 (N_22811,N_22736,N_22597);
xor U22812 (N_22812,N_22746,N_22640);
nor U22813 (N_22813,N_22543,N_22618);
or U22814 (N_22814,N_22735,N_22626);
xor U22815 (N_22815,N_22504,N_22603);
or U22816 (N_22816,N_22641,N_22686);
nand U22817 (N_22817,N_22699,N_22646);
xnor U22818 (N_22818,N_22726,N_22530);
nand U22819 (N_22819,N_22545,N_22749);
nor U22820 (N_22820,N_22537,N_22684);
nor U22821 (N_22821,N_22670,N_22523);
xor U22822 (N_22822,N_22666,N_22539);
or U22823 (N_22823,N_22674,N_22648);
xnor U22824 (N_22824,N_22654,N_22515);
and U22825 (N_22825,N_22619,N_22723);
or U22826 (N_22826,N_22542,N_22518);
and U22827 (N_22827,N_22599,N_22595);
nor U22828 (N_22828,N_22718,N_22553);
or U22829 (N_22829,N_22636,N_22598);
xor U22830 (N_22830,N_22709,N_22700);
or U22831 (N_22831,N_22676,N_22591);
nor U22832 (N_22832,N_22644,N_22548);
and U22833 (N_22833,N_22573,N_22706);
xnor U22834 (N_22834,N_22729,N_22649);
xnor U22835 (N_22835,N_22534,N_22743);
nand U22836 (N_22836,N_22705,N_22637);
nor U22837 (N_22837,N_22703,N_22547);
nand U22838 (N_22838,N_22563,N_22624);
and U22839 (N_22839,N_22634,N_22541);
xnor U22840 (N_22840,N_22662,N_22690);
and U22841 (N_22841,N_22663,N_22701);
nand U22842 (N_22842,N_22533,N_22579);
nor U22843 (N_22843,N_22711,N_22514);
xor U22844 (N_22844,N_22630,N_22585);
nor U22845 (N_22845,N_22517,N_22525);
xnor U22846 (N_22846,N_22647,N_22642);
and U22847 (N_22847,N_22608,N_22675);
xor U22848 (N_22848,N_22562,N_22601);
nor U22849 (N_22849,N_22569,N_22503);
or U22850 (N_22850,N_22531,N_22632);
and U22851 (N_22851,N_22578,N_22508);
and U22852 (N_22852,N_22532,N_22519);
nor U22853 (N_22853,N_22516,N_22740);
nor U22854 (N_22854,N_22685,N_22581);
nand U22855 (N_22855,N_22635,N_22720);
or U22856 (N_22856,N_22638,N_22639);
and U22857 (N_22857,N_22629,N_22607);
and U22858 (N_22858,N_22589,N_22725);
and U22859 (N_22859,N_22582,N_22695);
or U22860 (N_22860,N_22610,N_22734);
or U22861 (N_22861,N_22724,N_22713);
or U22862 (N_22862,N_22672,N_22574);
nor U22863 (N_22863,N_22580,N_22588);
xor U22864 (N_22864,N_22544,N_22512);
or U22865 (N_22865,N_22549,N_22721);
xnor U22866 (N_22866,N_22691,N_22747);
or U22867 (N_22867,N_22657,N_22692);
nor U22868 (N_22868,N_22683,N_22575);
nor U22869 (N_22869,N_22633,N_22714);
nand U22870 (N_22870,N_22650,N_22689);
nand U22871 (N_22871,N_22621,N_22617);
nor U22872 (N_22872,N_22628,N_22659);
nand U22873 (N_22873,N_22702,N_22554);
or U22874 (N_22874,N_22719,N_22745);
or U22875 (N_22875,N_22604,N_22532);
or U22876 (N_22876,N_22702,N_22531);
xor U22877 (N_22877,N_22544,N_22598);
nand U22878 (N_22878,N_22621,N_22720);
xor U22879 (N_22879,N_22711,N_22578);
or U22880 (N_22880,N_22671,N_22650);
nand U22881 (N_22881,N_22724,N_22648);
nand U22882 (N_22882,N_22623,N_22531);
or U22883 (N_22883,N_22682,N_22534);
and U22884 (N_22884,N_22735,N_22546);
or U22885 (N_22885,N_22573,N_22622);
and U22886 (N_22886,N_22616,N_22614);
and U22887 (N_22887,N_22698,N_22678);
and U22888 (N_22888,N_22737,N_22677);
nand U22889 (N_22889,N_22552,N_22559);
or U22890 (N_22890,N_22511,N_22620);
or U22891 (N_22891,N_22603,N_22748);
nor U22892 (N_22892,N_22713,N_22720);
or U22893 (N_22893,N_22562,N_22749);
or U22894 (N_22894,N_22585,N_22510);
or U22895 (N_22895,N_22606,N_22681);
nor U22896 (N_22896,N_22587,N_22659);
or U22897 (N_22897,N_22557,N_22657);
nor U22898 (N_22898,N_22667,N_22727);
and U22899 (N_22899,N_22660,N_22714);
or U22900 (N_22900,N_22669,N_22727);
and U22901 (N_22901,N_22681,N_22662);
nor U22902 (N_22902,N_22684,N_22600);
or U22903 (N_22903,N_22620,N_22581);
xor U22904 (N_22904,N_22556,N_22698);
xor U22905 (N_22905,N_22679,N_22697);
or U22906 (N_22906,N_22507,N_22744);
or U22907 (N_22907,N_22582,N_22600);
nand U22908 (N_22908,N_22618,N_22555);
nor U22909 (N_22909,N_22732,N_22645);
xor U22910 (N_22910,N_22692,N_22638);
nor U22911 (N_22911,N_22570,N_22666);
or U22912 (N_22912,N_22590,N_22671);
or U22913 (N_22913,N_22724,N_22613);
and U22914 (N_22914,N_22747,N_22556);
xnor U22915 (N_22915,N_22630,N_22623);
or U22916 (N_22916,N_22565,N_22532);
xnor U22917 (N_22917,N_22543,N_22501);
nor U22918 (N_22918,N_22570,N_22586);
nor U22919 (N_22919,N_22696,N_22566);
and U22920 (N_22920,N_22528,N_22744);
or U22921 (N_22921,N_22653,N_22590);
xor U22922 (N_22922,N_22693,N_22656);
nand U22923 (N_22923,N_22525,N_22705);
nand U22924 (N_22924,N_22537,N_22707);
nor U22925 (N_22925,N_22579,N_22640);
nor U22926 (N_22926,N_22525,N_22689);
or U22927 (N_22927,N_22610,N_22744);
xor U22928 (N_22928,N_22663,N_22721);
or U22929 (N_22929,N_22673,N_22551);
and U22930 (N_22930,N_22696,N_22600);
xnor U22931 (N_22931,N_22612,N_22566);
xor U22932 (N_22932,N_22700,N_22533);
and U22933 (N_22933,N_22707,N_22730);
xor U22934 (N_22934,N_22736,N_22741);
and U22935 (N_22935,N_22591,N_22720);
nor U22936 (N_22936,N_22644,N_22618);
and U22937 (N_22937,N_22641,N_22685);
or U22938 (N_22938,N_22627,N_22513);
xnor U22939 (N_22939,N_22528,N_22519);
nand U22940 (N_22940,N_22711,N_22616);
or U22941 (N_22941,N_22577,N_22726);
xor U22942 (N_22942,N_22722,N_22579);
or U22943 (N_22943,N_22581,N_22604);
and U22944 (N_22944,N_22661,N_22552);
xnor U22945 (N_22945,N_22746,N_22633);
or U22946 (N_22946,N_22749,N_22615);
nand U22947 (N_22947,N_22565,N_22508);
xnor U22948 (N_22948,N_22516,N_22674);
or U22949 (N_22949,N_22588,N_22728);
xor U22950 (N_22950,N_22580,N_22556);
xor U22951 (N_22951,N_22714,N_22540);
and U22952 (N_22952,N_22524,N_22523);
nand U22953 (N_22953,N_22541,N_22520);
and U22954 (N_22954,N_22697,N_22696);
and U22955 (N_22955,N_22621,N_22657);
and U22956 (N_22956,N_22638,N_22587);
nand U22957 (N_22957,N_22693,N_22629);
nor U22958 (N_22958,N_22527,N_22626);
nor U22959 (N_22959,N_22630,N_22731);
or U22960 (N_22960,N_22618,N_22656);
or U22961 (N_22961,N_22577,N_22668);
nor U22962 (N_22962,N_22697,N_22580);
or U22963 (N_22963,N_22618,N_22701);
nor U22964 (N_22964,N_22736,N_22502);
and U22965 (N_22965,N_22522,N_22543);
or U22966 (N_22966,N_22673,N_22602);
nand U22967 (N_22967,N_22538,N_22651);
nor U22968 (N_22968,N_22681,N_22536);
or U22969 (N_22969,N_22748,N_22725);
and U22970 (N_22970,N_22679,N_22568);
or U22971 (N_22971,N_22638,N_22598);
and U22972 (N_22972,N_22737,N_22509);
nand U22973 (N_22973,N_22593,N_22741);
nor U22974 (N_22974,N_22654,N_22701);
xor U22975 (N_22975,N_22601,N_22618);
xor U22976 (N_22976,N_22569,N_22590);
xor U22977 (N_22977,N_22540,N_22602);
xor U22978 (N_22978,N_22587,N_22612);
and U22979 (N_22979,N_22629,N_22502);
and U22980 (N_22980,N_22534,N_22609);
nand U22981 (N_22981,N_22637,N_22738);
nand U22982 (N_22982,N_22560,N_22674);
and U22983 (N_22983,N_22517,N_22523);
and U22984 (N_22984,N_22735,N_22624);
or U22985 (N_22985,N_22584,N_22574);
and U22986 (N_22986,N_22539,N_22559);
xnor U22987 (N_22987,N_22505,N_22724);
nor U22988 (N_22988,N_22606,N_22542);
xor U22989 (N_22989,N_22556,N_22567);
nand U22990 (N_22990,N_22537,N_22678);
nor U22991 (N_22991,N_22693,N_22744);
nor U22992 (N_22992,N_22698,N_22716);
nor U22993 (N_22993,N_22645,N_22639);
or U22994 (N_22994,N_22626,N_22724);
or U22995 (N_22995,N_22634,N_22667);
nor U22996 (N_22996,N_22582,N_22676);
and U22997 (N_22997,N_22744,N_22672);
and U22998 (N_22998,N_22597,N_22539);
nor U22999 (N_22999,N_22558,N_22697);
or U23000 (N_23000,N_22898,N_22809);
xnor U23001 (N_23001,N_22929,N_22866);
xor U23002 (N_23002,N_22807,N_22867);
nand U23003 (N_23003,N_22890,N_22893);
and U23004 (N_23004,N_22892,N_22824);
nor U23005 (N_23005,N_22934,N_22815);
or U23006 (N_23006,N_22774,N_22865);
or U23007 (N_23007,N_22902,N_22830);
or U23008 (N_23008,N_22861,N_22993);
nand U23009 (N_23009,N_22916,N_22833);
nand U23010 (N_23010,N_22941,N_22788);
xnor U23011 (N_23011,N_22996,N_22782);
and U23012 (N_23012,N_22918,N_22970);
and U23013 (N_23013,N_22963,N_22894);
and U23014 (N_23014,N_22797,N_22835);
and U23015 (N_23015,N_22876,N_22945);
and U23016 (N_23016,N_22755,N_22822);
or U23017 (N_23017,N_22883,N_22800);
nor U23018 (N_23018,N_22975,N_22956);
and U23019 (N_23019,N_22818,N_22864);
nor U23020 (N_23020,N_22952,N_22930);
or U23021 (N_23021,N_22966,N_22777);
nand U23022 (N_23022,N_22936,N_22753);
and U23023 (N_23023,N_22850,N_22926);
nor U23024 (N_23024,N_22968,N_22887);
xnor U23025 (N_23025,N_22779,N_22831);
and U23026 (N_23026,N_22816,N_22967);
xnor U23027 (N_23027,N_22962,N_22801);
or U23028 (N_23028,N_22857,N_22808);
and U23029 (N_23029,N_22954,N_22789);
nor U23030 (N_23030,N_22806,N_22879);
nor U23031 (N_23031,N_22812,N_22783);
or U23032 (N_23032,N_22889,N_22772);
nand U23033 (N_23033,N_22978,N_22798);
xor U23034 (N_23034,N_22762,N_22950);
or U23035 (N_23035,N_22886,N_22912);
nand U23036 (N_23036,N_22995,N_22903);
or U23037 (N_23037,N_22766,N_22776);
or U23038 (N_23038,N_22860,N_22919);
and U23039 (N_23039,N_22845,N_22829);
xnor U23040 (N_23040,N_22752,N_22909);
or U23041 (N_23041,N_22848,N_22947);
and U23042 (N_23042,N_22858,N_22870);
nor U23043 (N_23043,N_22946,N_22874);
or U23044 (N_23044,N_22884,N_22922);
or U23045 (N_23045,N_22924,N_22895);
xor U23046 (N_23046,N_22764,N_22820);
nand U23047 (N_23047,N_22986,N_22810);
nand U23048 (N_23048,N_22754,N_22940);
or U23049 (N_23049,N_22971,N_22997);
or U23050 (N_23050,N_22979,N_22759);
xnor U23051 (N_23051,N_22868,N_22969);
nor U23052 (N_23052,N_22987,N_22768);
nand U23053 (N_23053,N_22796,N_22852);
nor U23054 (N_23054,N_22790,N_22900);
nand U23055 (N_23055,N_22907,N_22972);
and U23056 (N_23056,N_22928,N_22836);
and U23057 (N_23057,N_22959,N_22942);
or U23058 (N_23058,N_22805,N_22990);
xor U23059 (N_23059,N_22846,N_22904);
nand U23060 (N_23060,N_22826,N_22957);
or U23061 (N_23061,N_22761,N_22856);
and U23062 (N_23062,N_22832,N_22961);
or U23063 (N_23063,N_22880,N_22758);
and U23064 (N_23064,N_22843,N_22825);
nor U23065 (N_23065,N_22778,N_22787);
xor U23066 (N_23066,N_22834,N_22780);
or U23067 (N_23067,N_22841,N_22877);
nand U23068 (N_23068,N_22793,N_22935);
or U23069 (N_23069,N_22974,N_22853);
xnor U23070 (N_23070,N_22786,N_22932);
or U23071 (N_23071,N_22844,N_22891);
nand U23072 (N_23072,N_22873,N_22765);
and U23073 (N_23073,N_22939,N_22994);
nor U23074 (N_23074,N_22855,N_22791);
xnor U23075 (N_23075,N_22985,N_22888);
nor U23076 (N_23076,N_22773,N_22803);
and U23077 (N_23077,N_22795,N_22821);
nand U23078 (N_23078,N_22911,N_22839);
nor U23079 (N_23079,N_22925,N_22785);
and U23080 (N_23080,N_22897,N_22794);
xor U23081 (N_23081,N_22770,N_22980);
and U23082 (N_23082,N_22988,N_22872);
xnor U23083 (N_23083,N_22944,N_22814);
nand U23084 (N_23084,N_22933,N_22854);
nor U23085 (N_23085,N_22949,N_22958);
and U23086 (N_23086,N_22955,N_22769);
and U23087 (N_23087,N_22960,N_22763);
xnor U23088 (N_23088,N_22869,N_22847);
nor U23089 (N_23089,N_22840,N_22849);
nor U23090 (N_23090,N_22842,N_22973);
xnor U23091 (N_23091,N_22981,N_22882);
nand U23092 (N_23092,N_22984,N_22906);
and U23093 (N_23093,N_22953,N_22965);
nand U23094 (N_23094,N_22998,N_22859);
nand U23095 (N_23095,N_22991,N_22863);
nor U23096 (N_23096,N_22784,N_22943);
nand U23097 (N_23097,N_22982,N_22781);
nand U23098 (N_23098,N_22823,N_22811);
xor U23099 (N_23099,N_22920,N_22802);
and U23100 (N_23100,N_22828,N_22751);
nand U23101 (N_23101,N_22771,N_22899);
or U23102 (N_23102,N_22804,N_22923);
or U23103 (N_23103,N_22896,N_22999);
or U23104 (N_23104,N_22851,N_22901);
nor U23105 (N_23105,N_22775,N_22976);
nor U23106 (N_23106,N_22827,N_22878);
and U23107 (N_23107,N_22819,N_22756);
nand U23108 (N_23108,N_22937,N_22799);
and U23109 (N_23109,N_22908,N_22910);
nand U23110 (N_23110,N_22917,N_22881);
nor U23111 (N_23111,N_22875,N_22767);
or U23112 (N_23112,N_22983,N_22905);
or U23113 (N_23113,N_22837,N_22792);
or U23114 (N_23114,N_22915,N_22862);
and U23115 (N_23115,N_22931,N_22989);
xnor U23116 (N_23116,N_22964,N_22951);
xnor U23117 (N_23117,N_22914,N_22760);
or U23118 (N_23118,N_22838,N_22992);
and U23119 (N_23119,N_22948,N_22871);
nor U23120 (N_23120,N_22813,N_22750);
xor U23121 (N_23121,N_22921,N_22757);
xor U23122 (N_23122,N_22913,N_22927);
and U23123 (N_23123,N_22885,N_22817);
or U23124 (N_23124,N_22938,N_22977);
xor U23125 (N_23125,N_22818,N_22829);
nor U23126 (N_23126,N_22986,N_22873);
nand U23127 (N_23127,N_22972,N_22750);
nand U23128 (N_23128,N_22791,N_22869);
nor U23129 (N_23129,N_22847,N_22812);
nor U23130 (N_23130,N_22829,N_22957);
or U23131 (N_23131,N_22911,N_22879);
and U23132 (N_23132,N_22854,N_22994);
and U23133 (N_23133,N_22874,N_22915);
nor U23134 (N_23134,N_22768,N_22841);
xnor U23135 (N_23135,N_22865,N_22810);
or U23136 (N_23136,N_22962,N_22763);
and U23137 (N_23137,N_22839,N_22822);
and U23138 (N_23138,N_22944,N_22841);
nor U23139 (N_23139,N_22768,N_22912);
xor U23140 (N_23140,N_22927,N_22844);
nand U23141 (N_23141,N_22930,N_22920);
xor U23142 (N_23142,N_22946,N_22997);
nand U23143 (N_23143,N_22800,N_22823);
and U23144 (N_23144,N_22787,N_22762);
and U23145 (N_23145,N_22944,N_22882);
xor U23146 (N_23146,N_22929,N_22860);
xnor U23147 (N_23147,N_22948,N_22908);
nor U23148 (N_23148,N_22783,N_22879);
or U23149 (N_23149,N_22845,N_22907);
or U23150 (N_23150,N_22838,N_22911);
xnor U23151 (N_23151,N_22900,N_22823);
nand U23152 (N_23152,N_22836,N_22876);
or U23153 (N_23153,N_22816,N_22819);
or U23154 (N_23154,N_22996,N_22979);
or U23155 (N_23155,N_22778,N_22757);
or U23156 (N_23156,N_22984,N_22932);
nand U23157 (N_23157,N_22848,N_22953);
nand U23158 (N_23158,N_22809,N_22967);
xnor U23159 (N_23159,N_22949,N_22960);
nor U23160 (N_23160,N_22983,N_22860);
nand U23161 (N_23161,N_22861,N_22777);
and U23162 (N_23162,N_22813,N_22904);
or U23163 (N_23163,N_22993,N_22840);
or U23164 (N_23164,N_22972,N_22904);
and U23165 (N_23165,N_22765,N_22941);
or U23166 (N_23166,N_22932,N_22804);
xor U23167 (N_23167,N_22764,N_22907);
or U23168 (N_23168,N_22870,N_22857);
xor U23169 (N_23169,N_22893,N_22915);
xor U23170 (N_23170,N_22968,N_22754);
nor U23171 (N_23171,N_22997,N_22757);
xnor U23172 (N_23172,N_22828,N_22939);
xnor U23173 (N_23173,N_22924,N_22859);
nand U23174 (N_23174,N_22932,N_22962);
nor U23175 (N_23175,N_22921,N_22832);
xnor U23176 (N_23176,N_22832,N_22779);
xor U23177 (N_23177,N_22886,N_22784);
xnor U23178 (N_23178,N_22756,N_22788);
or U23179 (N_23179,N_22834,N_22794);
nand U23180 (N_23180,N_22773,N_22825);
and U23181 (N_23181,N_22957,N_22981);
or U23182 (N_23182,N_22866,N_22923);
xor U23183 (N_23183,N_22919,N_22998);
and U23184 (N_23184,N_22956,N_22806);
xnor U23185 (N_23185,N_22789,N_22767);
or U23186 (N_23186,N_22967,N_22891);
xnor U23187 (N_23187,N_22975,N_22763);
xor U23188 (N_23188,N_22767,N_22896);
nand U23189 (N_23189,N_22939,N_22983);
xor U23190 (N_23190,N_22785,N_22949);
xor U23191 (N_23191,N_22948,N_22826);
nor U23192 (N_23192,N_22994,N_22933);
nor U23193 (N_23193,N_22958,N_22878);
or U23194 (N_23194,N_22936,N_22879);
and U23195 (N_23195,N_22902,N_22819);
or U23196 (N_23196,N_22976,N_22964);
nand U23197 (N_23197,N_22933,N_22819);
and U23198 (N_23198,N_22932,N_22787);
nand U23199 (N_23199,N_22936,N_22812);
and U23200 (N_23200,N_22950,N_22930);
or U23201 (N_23201,N_22859,N_22958);
xnor U23202 (N_23202,N_22915,N_22790);
and U23203 (N_23203,N_22776,N_22784);
nor U23204 (N_23204,N_22850,N_22811);
nand U23205 (N_23205,N_22940,N_22966);
and U23206 (N_23206,N_22885,N_22983);
nand U23207 (N_23207,N_22966,N_22830);
nand U23208 (N_23208,N_22813,N_22830);
and U23209 (N_23209,N_22965,N_22758);
nor U23210 (N_23210,N_22926,N_22762);
or U23211 (N_23211,N_22900,N_22906);
or U23212 (N_23212,N_22806,N_22779);
xor U23213 (N_23213,N_22902,N_22934);
nor U23214 (N_23214,N_22887,N_22816);
nand U23215 (N_23215,N_22830,N_22967);
xnor U23216 (N_23216,N_22865,N_22845);
and U23217 (N_23217,N_22756,N_22818);
xor U23218 (N_23218,N_22852,N_22813);
or U23219 (N_23219,N_22933,N_22936);
and U23220 (N_23220,N_22784,N_22845);
or U23221 (N_23221,N_22836,N_22884);
nand U23222 (N_23222,N_22890,N_22815);
xor U23223 (N_23223,N_22996,N_22826);
nor U23224 (N_23224,N_22916,N_22930);
nor U23225 (N_23225,N_22799,N_22869);
nor U23226 (N_23226,N_22832,N_22797);
nand U23227 (N_23227,N_22922,N_22779);
nand U23228 (N_23228,N_22897,N_22862);
or U23229 (N_23229,N_22882,N_22985);
and U23230 (N_23230,N_22785,N_22913);
and U23231 (N_23231,N_22914,N_22854);
xor U23232 (N_23232,N_22880,N_22839);
nand U23233 (N_23233,N_22820,N_22986);
xnor U23234 (N_23234,N_22880,N_22949);
nand U23235 (N_23235,N_22784,N_22887);
xnor U23236 (N_23236,N_22924,N_22813);
and U23237 (N_23237,N_22799,N_22806);
or U23238 (N_23238,N_22990,N_22825);
xor U23239 (N_23239,N_22789,N_22871);
nor U23240 (N_23240,N_22874,N_22994);
and U23241 (N_23241,N_22798,N_22785);
nand U23242 (N_23242,N_22792,N_22881);
nor U23243 (N_23243,N_22857,N_22929);
or U23244 (N_23244,N_22987,N_22946);
nand U23245 (N_23245,N_22893,N_22919);
and U23246 (N_23246,N_22787,N_22812);
xor U23247 (N_23247,N_22943,N_22874);
and U23248 (N_23248,N_22913,N_22948);
nand U23249 (N_23249,N_22928,N_22828);
xnor U23250 (N_23250,N_23235,N_23033);
or U23251 (N_23251,N_23016,N_23168);
xor U23252 (N_23252,N_23239,N_23194);
or U23253 (N_23253,N_23179,N_23096);
nand U23254 (N_23254,N_23025,N_23166);
xnor U23255 (N_23255,N_23092,N_23160);
or U23256 (N_23256,N_23066,N_23149);
or U23257 (N_23257,N_23020,N_23219);
and U23258 (N_23258,N_23228,N_23030);
and U23259 (N_23259,N_23104,N_23151);
or U23260 (N_23260,N_23086,N_23132);
nor U23261 (N_23261,N_23129,N_23039);
xor U23262 (N_23262,N_23084,N_23143);
and U23263 (N_23263,N_23165,N_23102);
nand U23264 (N_23264,N_23052,N_23050);
and U23265 (N_23265,N_23077,N_23126);
or U23266 (N_23266,N_23209,N_23237);
and U23267 (N_23267,N_23172,N_23090);
nor U23268 (N_23268,N_23138,N_23008);
and U23269 (N_23269,N_23013,N_23001);
nand U23270 (N_23270,N_23041,N_23247);
or U23271 (N_23271,N_23223,N_23206);
and U23272 (N_23272,N_23248,N_23245);
nor U23273 (N_23273,N_23007,N_23196);
nor U23274 (N_23274,N_23037,N_23119);
xnor U23275 (N_23275,N_23199,N_23024);
and U23276 (N_23276,N_23017,N_23015);
or U23277 (N_23277,N_23175,N_23216);
xor U23278 (N_23278,N_23082,N_23005);
xor U23279 (N_23279,N_23046,N_23002);
and U23280 (N_23280,N_23241,N_23061);
or U23281 (N_23281,N_23088,N_23014);
or U23282 (N_23282,N_23085,N_23230);
xor U23283 (N_23283,N_23226,N_23202);
xnor U23284 (N_23284,N_23079,N_23009);
nand U23285 (N_23285,N_23173,N_23038);
xor U23286 (N_23286,N_23064,N_23125);
xnor U23287 (N_23287,N_23070,N_23063);
xnor U23288 (N_23288,N_23011,N_23065);
or U23289 (N_23289,N_23116,N_23018);
or U23290 (N_23290,N_23184,N_23180);
xnor U23291 (N_23291,N_23191,N_23207);
nor U23292 (N_23292,N_23177,N_23128);
xor U23293 (N_23293,N_23100,N_23029);
nand U23294 (N_23294,N_23164,N_23000);
and U23295 (N_23295,N_23023,N_23187);
or U23296 (N_23296,N_23004,N_23112);
xor U23297 (N_23297,N_23130,N_23159);
nand U23298 (N_23298,N_23238,N_23121);
nand U23299 (N_23299,N_23019,N_23091);
or U23300 (N_23300,N_23156,N_23215);
or U23301 (N_23301,N_23072,N_23200);
or U23302 (N_23302,N_23056,N_23163);
nand U23303 (N_23303,N_23193,N_23081);
xnor U23304 (N_23304,N_23188,N_23148);
nand U23305 (N_23305,N_23097,N_23220);
nand U23306 (N_23306,N_23078,N_23227);
nor U23307 (N_23307,N_23040,N_23198);
and U23308 (N_23308,N_23074,N_23178);
and U23309 (N_23309,N_23221,N_23026);
or U23310 (N_23310,N_23089,N_23113);
nand U23311 (N_23311,N_23058,N_23045);
nor U23312 (N_23312,N_23076,N_23240);
and U23313 (N_23313,N_23003,N_23243);
nand U23314 (N_23314,N_23244,N_23242);
nor U23315 (N_23315,N_23142,N_23208);
nor U23316 (N_23316,N_23233,N_23204);
xnor U23317 (N_23317,N_23135,N_23028);
nand U23318 (N_23318,N_23152,N_23210);
nor U23319 (N_23319,N_23122,N_23162);
or U23320 (N_23320,N_23171,N_23048);
nand U23321 (N_23321,N_23150,N_23212);
xor U23322 (N_23322,N_23167,N_23186);
nor U23323 (N_23323,N_23010,N_23062);
or U23324 (N_23324,N_23139,N_23043);
and U23325 (N_23325,N_23176,N_23075);
nand U23326 (N_23326,N_23073,N_23124);
and U23327 (N_23327,N_23229,N_23140);
nand U23328 (N_23328,N_23211,N_23106);
nor U23329 (N_23329,N_23083,N_23021);
nand U23330 (N_23330,N_23114,N_23094);
nand U23331 (N_23331,N_23031,N_23236);
and U23332 (N_23332,N_23155,N_23141);
or U23333 (N_23333,N_23034,N_23055);
or U23334 (N_23334,N_23182,N_23123);
or U23335 (N_23335,N_23069,N_23190);
nand U23336 (N_23336,N_23195,N_23071);
xor U23337 (N_23337,N_23232,N_23225);
or U23338 (N_23338,N_23146,N_23203);
nor U23339 (N_23339,N_23117,N_23170);
xnor U23340 (N_23340,N_23214,N_23107);
or U23341 (N_23341,N_23218,N_23201);
and U23342 (N_23342,N_23153,N_23053);
or U23343 (N_23343,N_23067,N_23059);
xor U23344 (N_23344,N_23051,N_23012);
nand U23345 (N_23345,N_23099,N_23183);
or U23346 (N_23346,N_23246,N_23131);
nand U23347 (N_23347,N_23022,N_23103);
nor U23348 (N_23348,N_23093,N_23080);
nand U23349 (N_23349,N_23137,N_23049);
nand U23350 (N_23350,N_23042,N_23101);
nand U23351 (N_23351,N_23110,N_23205);
xnor U23352 (N_23352,N_23189,N_23127);
or U23353 (N_23353,N_23174,N_23234);
or U23354 (N_23354,N_23068,N_23098);
and U23355 (N_23355,N_23158,N_23027);
or U23356 (N_23356,N_23197,N_23036);
nand U23357 (N_23357,N_23109,N_23231);
nand U23358 (N_23358,N_23115,N_23136);
and U23359 (N_23359,N_23035,N_23144);
and U23360 (N_23360,N_23108,N_23032);
or U23361 (N_23361,N_23145,N_23185);
and U23362 (N_23362,N_23087,N_23105);
nand U23363 (N_23363,N_23120,N_23222);
and U23364 (N_23364,N_23224,N_23054);
nand U23365 (N_23365,N_23213,N_23154);
nor U23366 (N_23366,N_23192,N_23249);
nor U23367 (N_23367,N_23169,N_23047);
nand U23368 (N_23368,N_23157,N_23118);
xor U23369 (N_23369,N_23057,N_23134);
nor U23370 (N_23370,N_23133,N_23060);
xnor U23371 (N_23371,N_23217,N_23111);
nor U23372 (N_23372,N_23147,N_23044);
nor U23373 (N_23373,N_23006,N_23181);
and U23374 (N_23374,N_23161,N_23095);
and U23375 (N_23375,N_23021,N_23072);
and U23376 (N_23376,N_23027,N_23211);
xor U23377 (N_23377,N_23023,N_23165);
or U23378 (N_23378,N_23011,N_23189);
nand U23379 (N_23379,N_23123,N_23024);
and U23380 (N_23380,N_23021,N_23132);
nor U23381 (N_23381,N_23142,N_23141);
and U23382 (N_23382,N_23026,N_23124);
nor U23383 (N_23383,N_23038,N_23050);
nor U23384 (N_23384,N_23181,N_23038);
or U23385 (N_23385,N_23159,N_23212);
xor U23386 (N_23386,N_23110,N_23179);
or U23387 (N_23387,N_23135,N_23155);
and U23388 (N_23388,N_23058,N_23239);
xor U23389 (N_23389,N_23113,N_23041);
nor U23390 (N_23390,N_23027,N_23103);
and U23391 (N_23391,N_23209,N_23184);
or U23392 (N_23392,N_23150,N_23064);
nor U23393 (N_23393,N_23062,N_23232);
nor U23394 (N_23394,N_23246,N_23135);
nor U23395 (N_23395,N_23055,N_23038);
nand U23396 (N_23396,N_23038,N_23206);
xnor U23397 (N_23397,N_23183,N_23101);
or U23398 (N_23398,N_23064,N_23103);
nand U23399 (N_23399,N_23014,N_23214);
nand U23400 (N_23400,N_23005,N_23063);
nand U23401 (N_23401,N_23026,N_23102);
xnor U23402 (N_23402,N_23149,N_23174);
and U23403 (N_23403,N_23040,N_23025);
or U23404 (N_23404,N_23126,N_23018);
or U23405 (N_23405,N_23224,N_23070);
xor U23406 (N_23406,N_23113,N_23039);
and U23407 (N_23407,N_23171,N_23012);
and U23408 (N_23408,N_23179,N_23168);
or U23409 (N_23409,N_23046,N_23179);
nand U23410 (N_23410,N_23060,N_23208);
or U23411 (N_23411,N_23029,N_23230);
or U23412 (N_23412,N_23170,N_23004);
and U23413 (N_23413,N_23145,N_23162);
nand U23414 (N_23414,N_23108,N_23039);
nor U23415 (N_23415,N_23212,N_23146);
and U23416 (N_23416,N_23188,N_23130);
and U23417 (N_23417,N_23144,N_23125);
xor U23418 (N_23418,N_23006,N_23051);
and U23419 (N_23419,N_23049,N_23179);
or U23420 (N_23420,N_23224,N_23174);
or U23421 (N_23421,N_23029,N_23049);
nor U23422 (N_23422,N_23113,N_23025);
nand U23423 (N_23423,N_23202,N_23242);
xor U23424 (N_23424,N_23057,N_23053);
or U23425 (N_23425,N_23185,N_23000);
xnor U23426 (N_23426,N_23157,N_23111);
nand U23427 (N_23427,N_23157,N_23031);
and U23428 (N_23428,N_23227,N_23087);
xnor U23429 (N_23429,N_23004,N_23081);
nor U23430 (N_23430,N_23022,N_23045);
and U23431 (N_23431,N_23154,N_23095);
or U23432 (N_23432,N_23015,N_23111);
nor U23433 (N_23433,N_23076,N_23033);
xnor U23434 (N_23434,N_23143,N_23091);
xnor U23435 (N_23435,N_23045,N_23180);
nor U23436 (N_23436,N_23125,N_23182);
nor U23437 (N_23437,N_23153,N_23190);
and U23438 (N_23438,N_23191,N_23089);
nand U23439 (N_23439,N_23236,N_23123);
or U23440 (N_23440,N_23051,N_23035);
and U23441 (N_23441,N_23042,N_23178);
nor U23442 (N_23442,N_23141,N_23110);
nor U23443 (N_23443,N_23115,N_23202);
or U23444 (N_23444,N_23237,N_23116);
nor U23445 (N_23445,N_23031,N_23091);
and U23446 (N_23446,N_23175,N_23114);
and U23447 (N_23447,N_23166,N_23048);
or U23448 (N_23448,N_23179,N_23165);
nand U23449 (N_23449,N_23177,N_23166);
and U23450 (N_23450,N_23188,N_23027);
xor U23451 (N_23451,N_23241,N_23014);
and U23452 (N_23452,N_23123,N_23127);
xor U23453 (N_23453,N_23161,N_23076);
and U23454 (N_23454,N_23120,N_23067);
and U23455 (N_23455,N_23200,N_23146);
and U23456 (N_23456,N_23204,N_23169);
or U23457 (N_23457,N_23167,N_23200);
or U23458 (N_23458,N_23173,N_23014);
or U23459 (N_23459,N_23058,N_23067);
or U23460 (N_23460,N_23232,N_23212);
or U23461 (N_23461,N_23143,N_23111);
and U23462 (N_23462,N_23076,N_23039);
or U23463 (N_23463,N_23155,N_23090);
nand U23464 (N_23464,N_23240,N_23123);
or U23465 (N_23465,N_23133,N_23184);
xor U23466 (N_23466,N_23154,N_23124);
xor U23467 (N_23467,N_23155,N_23181);
nor U23468 (N_23468,N_23011,N_23124);
nor U23469 (N_23469,N_23123,N_23064);
nand U23470 (N_23470,N_23174,N_23191);
nand U23471 (N_23471,N_23220,N_23016);
and U23472 (N_23472,N_23186,N_23158);
xnor U23473 (N_23473,N_23009,N_23092);
and U23474 (N_23474,N_23157,N_23035);
nand U23475 (N_23475,N_23105,N_23186);
and U23476 (N_23476,N_23224,N_23097);
xnor U23477 (N_23477,N_23092,N_23152);
and U23478 (N_23478,N_23201,N_23150);
or U23479 (N_23479,N_23071,N_23144);
xor U23480 (N_23480,N_23146,N_23153);
or U23481 (N_23481,N_23134,N_23100);
and U23482 (N_23482,N_23223,N_23084);
and U23483 (N_23483,N_23041,N_23005);
nand U23484 (N_23484,N_23038,N_23095);
nand U23485 (N_23485,N_23203,N_23104);
and U23486 (N_23486,N_23012,N_23160);
nor U23487 (N_23487,N_23016,N_23177);
nand U23488 (N_23488,N_23122,N_23249);
or U23489 (N_23489,N_23079,N_23089);
and U23490 (N_23490,N_23205,N_23242);
xor U23491 (N_23491,N_23249,N_23038);
and U23492 (N_23492,N_23066,N_23185);
or U23493 (N_23493,N_23006,N_23088);
nand U23494 (N_23494,N_23171,N_23151);
nand U23495 (N_23495,N_23205,N_23215);
xnor U23496 (N_23496,N_23082,N_23175);
and U23497 (N_23497,N_23050,N_23235);
or U23498 (N_23498,N_23179,N_23198);
nand U23499 (N_23499,N_23190,N_23180);
nand U23500 (N_23500,N_23263,N_23494);
nand U23501 (N_23501,N_23471,N_23336);
or U23502 (N_23502,N_23309,N_23458);
xnor U23503 (N_23503,N_23372,N_23499);
xor U23504 (N_23504,N_23347,N_23270);
nor U23505 (N_23505,N_23370,N_23334);
nand U23506 (N_23506,N_23431,N_23492);
nor U23507 (N_23507,N_23386,N_23272);
nand U23508 (N_23508,N_23283,N_23444);
nor U23509 (N_23509,N_23475,N_23405);
nand U23510 (N_23510,N_23467,N_23424);
nor U23511 (N_23511,N_23407,N_23303);
nor U23512 (N_23512,N_23413,N_23310);
nand U23513 (N_23513,N_23417,N_23435);
nor U23514 (N_23514,N_23251,N_23432);
xor U23515 (N_23515,N_23252,N_23313);
xnor U23516 (N_23516,N_23394,N_23291);
or U23517 (N_23517,N_23393,N_23463);
and U23518 (N_23518,N_23285,N_23329);
xor U23519 (N_23519,N_23292,N_23462);
and U23520 (N_23520,N_23490,N_23275);
xnor U23521 (N_23521,N_23330,N_23469);
or U23522 (N_23522,N_23412,N_23383);
nand U23523 (N_23523,N_23367,N_23403);
nor U23524 (N_23524,N_23399,N_23437);
xnor U23525 (N_23525,N_23279,N_23489);
nor U23526 (N_23526,N_23306,N_23276);
nor U23527 (N_23527,N_23332,N_23409);
xnor U23528 (N_23528,N_23269,N_23391);
nor U23529 (N_23529,N_23355,N_23455);
nor U23530 (N_23530,N_23278,N_23398);
nand U23531 (N_23531,N_23449,N_23317);
nand U23532 (N_23532,N_23425,N_23316);
xnor U23533 (N_23533,N_23419,N_23312);
xor U23534 (N_23534,N_23302,N_23389);
and U23535 (N_23535,N_23408,N_23459);
and U23536 (N_23536,N_23445,N_23361);
nor U23537 (N_23537,N_23327,N_23268);
nand U23538 (N_23538,N_23371,N_23447);
nand U23539 (N_23539,N_23300,N_23356);
xnor U23540 (N_23540,N_23301,N_23296);
xor U23541 (N_23541,N_23480,N_23464);
xor U23542 (N_23542,N_23438,N_23323);
nor U23543 (N_23543,N_23390,N_23486);
nor U23544 (N_23544,N_23253,N_23457);
nor U23545 (N_23545,N_23271,N_23344);
or U23546 (N_23546,N_23274,N_23326);
and U23547 (N_23547,N_23456,N_23369);
xor U23548 (N_23548,N_23422,N_23363);
and U23549 (N_23549,N_23476,N_23266);
xor U23550 (N_23550,N_23345,N_23293);
or U23551 (N_23551,N_23428,N_23402);
nand U23552 (N_23552,N_23346,N_23325);
nor U23553 (N_23553,N_23396,N_23290);
xor U23554 (N_23554,N_23482,N_23477);
nand U23555 (N_23555,N_23374,N_23359);
xor U23556 (N_23556,N_23314,N_23453);
xor U23557 (N_23557,N_23362,N_23259);
nand U23558 (N_23558,N_23348,N_23255);
nand U23559 (N_23559,N_23380,N_23420);
xnor U23560 (N_23560,N_23258,N_23260);
nor U23561 (N_23561,N_23388,N_23441);
nor U23562 (N_23562,N_23448,N_23415);
and U23563 (N_23563,N_23440,N_23421);
xor U23564 (N_23564,N_23365,N_23339);
nand U23565 (N_23565,N_23395,N_23360);
xnor U23566 (N_23566,N_23442,N_23331);
xnor U23567 (N_23567,N_23351,N_23321);
nand U23568 (N_23568,N_23414,N_23354);
and U23569 (N_23569,N_23267,N_23304);
and U23570 (N_23570,N_23277,N_23384);
nor U23571 (N_23571,N_23335,N_23495);
and U23572 (N_23572,N_23484,N_23483);
nor U23573 (N_23573,N_23493,N_23400);
and U23574 (N_23574,N_23288,N_23257);
or U23575 (N_23575,N_23350,N_23311);
and U23576 (N_23576,N_23295,N_23443);
and U23577 (N_23577,N_23382,N_23468);
nor U23578 (N_23578,N_23377,N_23379);
nand U23579 (N_23579,N_23322,N_23397);
or U23580 (N_23580,N_23479,N_23284);
xor U23581 (N_23581,N_23299,N_23439);
and U23582 (N_23582,N_23433,N_23466);
xnor U23583 (N_23583,N_23411,N_23497);
nand U23584 (N_23584,N_23308,N_23488);
nor U23585 (N_23585,N_23423,N_23294);
nor U23586 (N_23586,N_23426,N_23446);
and U23587 (N_23587,N_23470,N_23474);
and U23588 (N_23588,N_23481,N_23373);
or U23589 (N_23589,N_23315,N_23385);
or U23590 (N_23590,N_23454,N_23282);
and U23591 (N_23591,N_23298,N_23320);
nor U23592 (N_23592,N_23496,N_23460);
and U23593 (N_23593,N_23485,N_23307);
nor U23594 (N_23594,N_23472,N_23436);
xor U23595 (N_23595,N_23429,N_23358);
or U23596 (N_23596,N_23392,N_23343);
xnor U23597 (N_23597,N_23498,N_23364);
or U23598 (N_23598,N_23450,N_23318);
nand U23599 (N_23599,N_23281,N_23319);
nand U23600 (N_23600,N_23262,N_23418);
or U23601 (N_23601,N_23340,N_23366);
and U23602 (N_23602,N_23341,N_23280);
nor U23603 (N_23603,N_23349,N_23461);
xnor U23604 (N_23604,N_23478,N_23376);
nor U23605 (N_23605,N_23297,N_23273);
and U23606 (N_23606,N_23451,N_23410);
nand U23607 (N_23607,N_23427,N_23491);
nor U23608 (N_23608,N_23256,N_23465);
or U23609 (N_23609,N_23342,N_23261);
xnor U23610 (N_23610,N_23254,N_23352);
or U23611 (N_23611,N_23406,N_23487);
xnor U23612 (N_23612,N_23324,N_23286);
nor U23613 (N_23613,N_23381,N_23401);
nand U23614 (N_23614,N_23264,N_23434);
or U23615 (N_23615,N_23473,N_23250);
and U23616 (N_23616,N_23375,N_23368);
or U23617 (N_23617,N_23378,N_23333);
and U23618 (N_23618,N_23337,N_23430);
xor U23619 (N_23619,N_23452,N_23387);
xnor U23620 (N_23620,N_23416,N_23338);
nand U23621 (N_23621,N_23265,N_23289);
nor U23622 (N_23622,N_23357,N_23353);
xnor U23623 (N_23623,N_23287,N_23328);
nor U23624 (N_23624,N_23305,N_23404);
nand U23625 (N_23625,N_23386,N_23349);
xor U23626 (N_23626,N_23255,N_23411);
xor U23627 (N_23627,N_23304,N_23385);
or U23628 (N_23628,N_23364,N_23400);
and U23629 (N_23629,N_23370,N_23300);
xnor U23630 (N_23630,N_23400,N_23376);
xnor U23631 (N_23631,N_23321,N_23350);
nand U23632 (N_23632,N_23272,N_23266);
and U23633 (N_23633,N_23344,N_23439);
nor U23634 (N_23634,N_23413,N_23438);
and U23635 (N_23635,N_23375,N_23304);
xnor U23636 (N_23636,N_23424,N_23356);
and U23637 (N_23637,N_23304,N_23423);
xor U23638 (N_23638,N_23426,N_23458);
or U23639 (N_23639,N_23329,N_23483);
nor U23640 (N_23640,N_23460,N_23469);
and U23641 (N_23641,N_23382,N_23346);
or U23642 (N_23642,N_23487,N_23400);
nor U23643 (N_23643,N_23359,N_23349);
and U23644 (N_23644,N_23289,N_23379);
or U23645 (N_23645,N_23341,N_23256);
xnor U23646 (N_23646,N_23326,N_23261);
nor U23647 (N_23647,N_23288,N_23432);
or U23648 (N_23648,N_23343,N_23407);
nor U23649 (N_23649,N_23484,N_23306);
nor U23650 (N_23650,N_23461,N_23454);
and U23651 (N_23651,N_23365,N_23276);
xor U23652 (N_23652,N_23360,N_23471);
xnor U23653 (N_23653,N_23381,N_23369);
or U23654 (N_23654,N_23404,N_23277);
and U23655 (N_23655,N_23347,N_23252);
xnor U23656 (N_23656,N_23376,N_23356);
nor U23657 (N_23657,N_23467,N_23445);
xnor U23658 (N_23658,N_23289,N_23433);
and U23659 (N_23659,N_23301,N_23318);
or U23660 (N_23660,N_23277,N_23431);
xor U23661 (N_23661,N_23332,N_23432);
nand U23662 (N_23662,N_23371,N_23423);
or U23663 (N_23663,N_23312,N_23281);
and U23664 (N_23664,N_23474,N_23413);
nand U23665 (N_23665,N_23480,N_23416);
or U23666 (N_23666,N_23420,N_23424);
nand U23667 (N_23667,N_23330,N_23304);
nand U23668 (N_23668,N_23289,N_23408);
or U23669 (N_23669,N_23278,N_23366);
and U23670 (N_23670,N_23344,N_23465);
and U23671 (N_23671,N_23489,N_23286);
and U23672 (N_23672,N_23335,N_23408);
nand U23673 (N_23673,N_23426,N_23414);
or U23674 (N_23674,N_23400,N_23465);
nand U23675 (N_23675,N_23296,N_23417);
and U23676 (N_23676,N_23391,N_23499);
and U23677 (N_23677,N_23415,N_23492);
and U23678 (N_23678,N_23274,N_23441);
or U23679 (N_23679,N_23375,N_23399);
nor U23680 (N_23680,N_23381,N_23483);
or U23681 (N_23681,N_23377,N_23472);
xnor U23682 (N_23682,N_23443,N_23394);
nand U23683 (N_23683,N_23265,N_23273);
xnor U23684 (N_23684,N_23384,N_23292);
nand U23685 (N_23685,N_23357,N_23286);
or U23686 (N_23686,N_23499,N_23440);
and U23687 (N_23687,N_23399,N_23310);
nand U23688 (N_23688,N_23440,N_23405);
or U23689 (N_23689,N_23492,N_23380);
and U23690 (N_23690,N_23450,N_23365);
and U23691 (N_23691,N_23396,N_23288);
or U23692 (N_23692,N_23397,N_23333);
and U23693 (N_23693,N_23254,N_23398);
and U23694 (N_23694,N_23347,N_23433);
or U23695 (N_23695,N_23425,N_23479);
xor U23696 (N_23696,N_23288,N_23301);
nor U23697 (N_23697,N_23439,N_23386);
nor U23698 (N_23698,N_23396,N_23374);
nor U23699 (N_23699,N_23405,N_23416);
nand U23700 (N_23700,N_23259,N_23272);
and U23701 (N_23701,N_23425,N_23267);
and U23702 (N_23702,N_23473,N_23477);
nor U23703 (N_23703,N_23253,N_23351);
or U23704 (N_23704,N_23370,N_23298);
nor U23705 (N_23705,N_23454,N_23253);
nor U23706 (N_23706,N_23255,N_23287);
nor U23707 (N_23707,N_23359,N_23446);
nor U23708 (N_23708,N_23340,N_23425);
nor U23709 (N_23709,N_23301,N_23260);
nor U23710 (N_23710,N_23398,N_23325);
nand U23711 (N_23711,N_23498,N_23414);
or U23712 (N_23712,N_23370,N_23254);
nand U23713 (N_23713,N_23476,N_23284);
or U23714 (N_23714,N_23459,N_23498);
nand U23715 (N_23715,N_23347,N_23457);
xnor U23716 (N_23716,N_23448,N_23450);
xnor U23717 (N_23717,N_23306,N_23263);
or U23718 (N_23718,N_23414,N_23298);
or U23719 (N_23719,N_23383,N_23334);
and U23720 (N_23720,N_23419,N_23250);
xor U23721 (N_23721,N_23337,N_23310);
or U23722 (N_23722,N_23359,N_23435);
xor U23723 (N_23723,N_23405,N_23337);
nand U23724 (N_23724,N_23362,N_23336);
nor U23725 (N_23725,N_23458,N_23386);
xor U23726 (N_23726,N_23269,N_23418);
nor U23727 (N_23727,N_23485,N_23368);
xor U23728 (N_23728,N_23452,N_23421);
or U23729 (N_23729,N_23264,N_23484);
nor U23730 (N_23730,N_23351,N_23435);
nand U23731 (N_23731,N_23292,N_23347);
or U23732 (N_23732,N_23413,N_23464);
xor U23733 (N_23733,N_23471,N_23252);
nand U23734 (N_23734,N_23291,N_23279);
or U23735 (N_23735,N_23436,N_23498);
nor U23736 (N_23736,N_23272,N_23310);
nand U23737 (N_23737,N_23437,N_23416);
nor U23738 (N_23738,N_23412,N_23469);
xnor U23739 (N_23739,N_23333,N_23254);
or U23740 (N_23740,N_23473,N_23335);
and U23741 (N_23741,N_23438,N_23338);
nand U23742 (N_23742,N_23290,N_23273);
nor U23743 (N_23743,N_23298,N_23312);
or U23744 (N_23744,N_23350,N_23291);
xor U23745 (N_23745,N_23323,N_23278);
and U23746 (N_23746,N_23409,N_23250);
xnor U23747 (N_23747,N_23335,N_23355);
or U23748 (N_23748,N_23384,N_23413);
nand U23749 (N_23749,N_23255,N_23297);
or U23750 (N_23750,N_23553,N_23652);
or U23751 (N_23751,N_23701,N_23632);
nor U23752 (N_23752,N_23559,N_23589);
and U23753 (N_23753,N_23562,N_23643);
and U23754 (N_23754,N_23548,N_23735);
and U23755 (N_23755,N_23619,N_23561);
or U23756 (N_23756,N_23539,N_23695);
nand U23757 (N_23757,N_23745,N_23663);
xor U23758 (N_23758,N_23637,N_23599);
nor U23759 (N_23759,N_23710,N_23697);
nand U23760 (N_23760,N_23602,N_23593);
xnor U23761 (N_23761,N_23542,N_23666);
nand U23762 (N_23762,N_23534,N_23521);
xnor U23763 (N_23763,N_23565,N_23721);
nor U23764 (N_23764,N_23596,N_23504);
or U23765 (N_23765,N_23597,N_23714);
or U23766 (N_23766,N_23635,N_23578);
or U23767 (N_23767,N_23513,N_23654);
or U23768 (N_23768,N_23517,N_23647);
and U23769 (N_23769,N_23516,N_23669);
nor U23770 (N_23770,N_23733,N_23744);
or U23771 (N_23771,N_23511,N_23688);
nor U23772 (N_23772,N_23625,N_23687);
nor U23773 (N_23773,N_23529,N_23698);
xnor U23774 (N_23774,N_23712,N_23560);
nor U23775 (N_23775,N_23677,N_23607);
xnor U23776 (N_23776,N_23732,N_23556);
or U23777 (N_23777,N_23684,N_23614);
and U23778 (N_23778,N_23613,N_23582);
or U23779 (N_23779,N_23685,N_23543);
and U23780 (N_23780,N_23609,N_23629);
and U23781 (N_23781,N_23734,N_23623);
or U23782 (N_23782,N_23700,N_23514);
nor U23783 (N_23783,N_23544,N_23610);
xor U23784 (N_23784,N_23678,N_23502);
nor U23785 (N_23785,N_23689,N_23691);
or U23786 (N_23786,N_23546,N_23527);
nand U23787 (N_23787,N_23672,N_23657);
nand U23788 (N_23788,N_23743,N_23645);
nand U23789 (N_23789,N_23603,N_23533);
or U23790 (N_23790,N_23665,N_23579);
xnor U23791 (N_23791,N_23711,N_23650);
and U23792 (N_23792,N_23584,N_23501);
nand U23793 (N_23793,N_23611,N_23592);
nand U23794 (N_23794,N_23523,N_23740);
nor U23795 (N_23795,N_23587,N_23670);
or U23796 (N_23796,N_23627,N_23616);
nand U23797 (N_23797,N_23736,N_23628);
nor U23798 (N_23798,N_23588,N_23651);
nor U23799 (N_23799,N_23550,N_23532);
or U23800 (N_23800,N_23633,N_23692);
and U23801 (N_23801,N_23737,N_23620);
xor U23802 (N_23802,N_23624,N_23617);
nor U23803 (N_23803,N_23601,N_23673);
and U23804 (N_23804,N_23549,N_23622);
or U23805 (N_23805,N_23715,N_23708);
and U23806 (N_23806,N_23634,N_23545);
nor U23807 (N_23807,N_23524,N_23717);
and U23808 (N_23808,N_23644,N_23720);
nor U23809 (N_23809,N_23705,N_23551);
or U23810 (N_23810,N_23581,N_23572);
and U23811 (N_23811,N_23640,N_23600);
and U23812 (N_23812,N_23509,N_23630);
xor U23813 (N_23813,N_23503,N_23659);
nor U23814 (N_23814,N_23646,N_23583);
or U23815 (N_23815,N_23585,N_23569);
and U23816 (N_23816,N_23727,N_23500);
xor U23817 (N_23817,N_23664,N_23703);
or U23818 (N_23818,N_23704,N_23515);
and U23819 (N_23819,N_23668,N_23571);
or U23820 (N_23820,N_23605,N_23580);
xnor U23821 (N_23821,N_23725,N_23508);
or U23822 (N_23822,N_23747,N_23591);
xor U23823 (N_23823,N_23731,N_23719);
nor U23824 (N_23824,N_23656,N_23618);
nand U23825 (N_23825,N_23739,N_23676);
and U23826 (N_23826,N_23520,N_23537);
nor U23827 (N_23827,N_23526,N_23575);
xnor U23828 (N_23828,N_23555,N_23748);
nand U23829 (N_23829,N_23730,N_23626);
or U23830 (N_23830,N_23648,N_23594);
or U23831 (N_23831,N_23638,N_23519);
xor U23832 (N_23832,N_23636,N_23577);
and U23833 (N_23833,N_23649,N_23686);
and U23834 (N_23834,N_23709,N_23724);
and U23835 (N_23835,N_23506,N_23671);
or U23836 (N_23836,N_23604,N_23749);
and U23837 (N_23837,N_23507,N_23612);
or U23838 (N_23838,N_23682,N_23696);
nand U23839 (N_23839,N_23718,N_23573);
or U23840 (N_23840,N_23655,N_23552);
xor U23841 (N_23841,N_23538,N_23512);
or U23842 (N_23842,N_23693,N_23510);
nor U23843 (N_23843,N_23570,N_23699);
and U23844 (N_23844,N_23590,N_23658);
xnor U23845 (N_23845,N_23707,N_23528);
nor U23846 (N_23846,N_23680,N_23728);
nand U23847 (N_23847,N_23631,N_23681);
nor U23848 (N_23848,N_23505,N_23729);
or U23849 (N_23849,N_23531,N_23536);
nand U23850 (N_23850,N_23621,N_23595);
xnor U23851 (N_23851,N_23530,N_23564);
or U23852 (N_23852,N_23726,N_23683);
nor U23853 (N_23853,N_23723,N_23547);
xor U23854 (N_23854,N_23706,N_23694);
xnor U23855 (N_23855,N_23557,N_23679);
xnor U23856 (N_23856,N_23674,N_23716);
nor U23857 (N_23857,N_23661,N_23522);
xor U23858 (N_23858,N_23525,N_23606);
and U23859 (N_23859,N_23642,N_23608);
xor U23860 (N_23860,N_23563,N_23574);
and U23861 (N_23861,N_23639,N_23566);
nand U23862 (N_23862,N_23518,N_23690);
nor U23863 (N_23863,N_23576,N_23702);
or U23864 (N_23864,N_23535,N_23586);
and U23865 (N_23865,N_23746,N_23660);
nand U23866 (N_23866,N_23741,N_23558);
xnor U23867 (N_23867,N_23641,N_23540);
and U23868 (N_23868,N_23738,N_23568);
or U23869 (N_23869,N_23653,N_23554);
or U23870 (N_23870,N_23667,N_23662);
xor U23871 (N_23871,N_23567,N_23742);
nor U23872 (N_23872,N_23675,N_23541);
nand U23873 (N_23873,N_23615,N_23722);
or U23874 (N_23874,N_23598,N_23713);
and U23875 (N_23875,N_23541,N_23587);
and U23876 (N_23876,N_23611,N_23541);
xnor U23877 (N_23877,N_23726,N_23678);
nor U23878 (N_23878,N_23682,N_23694);
or U23879 (N_23879,N_23511,N_23574);
nand U23880 (N_23880,N_23522,N_23602);
nand U23881 (N_23881,N_23598,N_23557);
xor U23882 (N_23882,N_23638,N_23575);
and U23883 (N_23883,N_23576,N_23581);
and U23884 (N_23884,N_23501,N_23717);
nor U23885 (N_23885,N_23693,N_23636);
nand U23886 (N_23886,N_23584,N_23574);
nor U23887 (N_23887,N_23540,N_23541);
xor U23888 (N_23888,N_23550,N_23580);
or U23889 (N_23889,N_23554,N_23647);
or U23890 (N_23890,N_23652,N_23544);
xor U23891 (N_23891,N_23582,N_23504);
nand U23892 (N_23892,N_23656,N_23568);
nand U23893 (N_23893,N_23638,N_23527);
nand U23894 (N_23894,N_23543,N_23638);
and U23895 (N_23895,N_23654,N_23649);
nand U23896 (N_23896,N_23744,N_23674);
xnor U23897 (N_23897,N_23513,N_23697);
and U23898 (N_23898,N_23683,N_23714);
and U23899 (N_23899,N_23572,N_23548);
nand U23900 (N_23900,N_23622,N_23621);
or U23901 (N_23901,N_23500,N_23618);
xor U23902 (N_23902,N_23573,N_23584);
xor U23903 (N_23903,N_23732,N_23688);
or U23904 (N_23904,N_23718,N_23523);
and U23905 (N_23905,N_23661,N_23533);
nor U23906 (N_23906,N_23626,N_23554);
or U23907 (N_23907,N_23504,N_23513);
nor U23908 (N_23908,N_23655,N_23536);
and U23909 (N_23909,N_23510,N_23644);
and U23910 (N_23910,N_23612,N_23666);
xnor U23911 (N_23911,N_23726,N_23665);
or U23912 (N_23912,N_23637,N_23530);
or U23913 (N_23913,N_23741,N_23573);
or U23914 (N_23914,N_23674,N_23649);
nand U23915 (N_23915,N_23679,N_23529);
and U23916 (N_23916,N_23671,N_23537);
xnor U23917 (N_23917,N_23724,N_23536);
xnor U23918 (N_23918,N_23612,N_23546);
nor U23919 (N_23919,N_23723,N_23552);
nor U23920 (N_23920,N_23649,N_23734);
nor U23921 (N_23921,N_23606,N_23696);
nor U23922 (N_23922,N_23515,N_23562);
nor U23923 (N_23923,N_23606,N_23592);
xnor U23924 (N_23924,N_23641,N_23716);
nand U23925 (N_23925,N_23743,N_23643);
xor U23926 (N_23926,N_23546,N_23736);
xnor U23927 (N_23927,N_23507,N_23531);
nand U23928 (N_23928,N_23542,N_23634);
nand U23929 (N_23929,N_23557,N_23670);
or U23930 (N_23930,N_23630,N_23530);
nand U23931 (N_23931,N_23743,N_23584);
or U23932 (N_23932,N_23656,N_23524);
nand U23933 (N_23933,N_23704,N_23666);
and U23934 (N_23934,N_23602,N_23647);
or U23935 (N_23935,N_23502,N_23650);
xor U23936 (N_23936,N_23646,N_23651);
and U23937 (N_23937,N_23645,N_23551);
nand U23938 (N_23938,N_23535,N_23645);
nand U23939 (N_23939,N_23737,N_23629);
nor U23940 (N_23940,N_23701,N_23593);
nand U23941 (N_23941,N_23741,N_23603);
or U23942 (N_23942,N_23668,N_23559);
nor U23943 (N_23943,N_23517,N_23549);
xnor U23944 (N_23944,N_23665,N_23706);
nand U23945 (N_23945,N_23553,N_23501);
or U23946 (N_23946,N_23615,N_23562);
nor U23947 (N_23947,N_23626,N_23597);
xor U23948 (N_23948,N_23716,N_23711);
xnor U23949 (N_23949,N_23604,N_23730);
xnor U23950 (N_23950,N_23515,N_23612);
xnor U23951 (N_23951,N_23679,N_23732);
nor U23952 (N_23952,N_23582,N_23554);
nor U23953 (N_23953,N_23505,N_23519);
nor U23954 (N_23954,N_23717,N_23515);
and U23955 (N_23955,N_23585,N_23509);
nor U23956 (N_23956,N_23594,N_23522);
nor U23957 (N_23957,N_23596,N_23539);
and U23958 (N_23958,N_23515,N_23623);
nand U23959 (N_23959,N_23584,N_23575);
or U23960 (N_23960,N_23608,N_23618);
xnor U23961 (N_23961,N_23583,N_23551);
or U23962 (N_23962,N_23504,N_23744);
and U23963 (N_23963,N_23518,N_23660);
and U23964 (N_23964,N_23501,N_23677);
or U23965 (N_23965,N_23535,N_23745);
and U23966 (N_23966,N_23594,N_23571);
nand U23967 (N_23967,N_23714,N_23572);
or U23968 (N_23968,N_23597,N_23573);
nand U23969 (N_23969,N_23654,N_23630);
nor U23970 (N_23970,N_23748,N_23558);
or U23971 (N_23971,N_23643,N_23651);
and U23972 (N_23972,N_23670,N_23654);
xnor U23973 (N_23973,N_23668,N_23591);
and U23974 (N_23974,N_23579,N_23642);
xnor U23975 (N_23975,N_23675,N_23515);
or U23976 (N_23976,N_23527,N_23681);
and U23977 (N_23977,N_23635,N_23667);
nor U23978 (N_23978,N_23736,N_23708);
nor U23979 (N_23979,N_23679,N_23692);
nand U23980 (N_23980,N_23686,N_23565);
nor U23981 (N_23981,N_23709,N_23690);
xor U23982 (N_23982,N_23587,N_23547);
or U23983 (N_23983,N_23612,N_23606);
nand U23984 (N_23984,N_23569,N_23579);
and U23985 (N_23985,N_23701,N_23665);
or U23986 (N_23986,N_23516,N_23539);
xor U23987 (N_23987,N_23640,N_23650);
xnor U23988 (N_23988,N_23740,N_23634);
nand U23989 (N_23989,N_23664,N_23636);
xor U23990 (N_23990,N_23636,N_23624);
xnor U23991 (N_23991,N_23728,N_23627);
and U23992 (N_23992,N_23665,N_23557);
xor U23993 (N_23993,N_23690,N_23512);
and U23994 (N_23994,N_23706,N_23581);
or U23995 (N_23995,N_23720,N_23705);
xor U23996 (N_23996,N_23536,N_23674);
or U23997 (N_23997,N_23726,N_23589);
nor U23998 (N_23998,N_23721,N_23638);
nor U23999 (N_23999,N_23636,N_23515);
or U24000 (N_24000,N_23786,N_23908);
or U24001 (N_24001,N_23923,N_23966);
nor U24002 (N_24002,N_23895,N_23911);
and U24003 (N_24003,N_23945,N_23819);
nor U24004 (N_24004,N_23858,N_23826);
or U24005 (N_24005,N_23791,N_23909);
nor U24006 (N_24006,N_23990,N_23825);
nor U24007 (N_24007,N_23868,N_23914);
xnor U24008 (N_24008,N_23934,N_23976);
xor U24009 (N_24009,N_23765,N_23827);
xor U24010 (N_24010,N_23770,N_23958);
xnor U24011 (N_24011,N_23939,N_23796);
or U24012 (N_24012,N_23954,N_23822);
xor U24013 (N_24013,N_23758,N_23899);
or U24014 (N_24014,N_23834,N_23871);
nand U24015 (N_24015,N_23855,N_23805);
and U24016 (N_24016,N_23901,N_23757);
and U24017 (N_24017,N_23982,N_23853);
and U24018 (N_24018,N_23836,N_23944);
and U24019 (N_24019,N_23813,N_23994);
nand U24020 (N_24020,N_23929,N_23949);
and U24021 (N_24021,N_23856,N_23927);
nand U24022 (N_24022,N_23861,N_23972);
nand U24023 (N_24023,N_23751,N_23788);
nand U24024 (N_24024,N_23832,N_23951);
or U24025 (N_24025,N_23844,N_23814);
xnor U24026 (N_24026,N_23970,N_23877);
nor U24027 (N_24027,N_23857,N_23953);
nor U24028 (N_24028,N_23969,N_23897);
or U24029 (N_24029,N_23938,N_23883);
xnor U24030 (N_24030,N_23917,N_23962);
nand U24031 (N_24031,N_23866,N_23925);
xor U24032 (N_24032,N_23991,N_23987);
and U24033 (N_24033,N_23816,N_23869);
and U24034 (N_24034,N_23759,N_23965);
nor U24035 (N_24035,N_23960,N_23766);
nor U24036 (N_24036,N_23879,N_23792);
nand U24037 (N_24037,N_23784,N_23957);
and U24038 (N_24038,N_23943,N_23946);
or U24039 (N_24039,N_23754,N_23812);
or U24040 (N_24040,N_23891,N_23961);
nand U24041 (N_24041,N_23886,N_23763);
or U24042 (N_24042,N_23829,N_23773);
xnor U24043 (N_24043,N_23959,N_23935);
nand U24044 (N_24044,N_23881,N_23806);
nand U24045 (N_24045,N_23797,N_23808);
nand U24046 (N_24046,N_23824,N_23838);
xor U24047 (N_24047,N_23867,N_23833);
nor U24048 (N_24048,N_23874,N_23811);
xnor U24049 (N_24049,N_23997,N_23980);
or U24050 (N_24050,N_23913,N_23842);
xor U24051 (N_24051,N_23892,N_23986);
and U24052 (N_24052,N_23907,N_23756);
nor U24053 (N_24053,N_23904,N_23978);
and U24054 (N_24054,N_23985,N_23801);
xor U24055 (N_24055,N_23890,N_23823);
or U24056 (N_24056,N_23998,N_23817);
and U24057 (N_24057,N_23936,N_23820);
xor U24058 (N_24058,N_23884,N_23903);
or U24059 (N_24059,N_23798,N_23835);
or U24060 (N_24060,N_23840,N_23989);
nor U24061 (N_24061,N_23768,N_23888);
nor U24062 (N_24062,N_23789,N_23984);
nand U24063 (N_24063,N_23956,N_23931);
xnor U24064 (N_24064,N_23849,N_23898);
nor U24065 (N_24065,N_23932,N_23963);
or U24066 (N_24066,N_23878,N_23782);
xor U24067 (N_24067,N_23802,N_23807);
nand U24068 (N_24068,N_23950,N_23981);
or U24069 (N_24069,N_23906,N_23947);
xor U24070 (N_24070,N_23865,N_23845);
and U24071 (N_24071,N_23780,N_23775);
or U24072 (N_24072,N_23771,N_23912);
xnor U24073 (N_24073,N_23922,N_23988);
xnor U24074 (N_24074,N_23772,N_23837);
nor U24075 (N_24075,N_23937,N_23755);
or U24076 (N_24076,N_23809,N_23921);
nor U24077 (N_24077,N_23841,N_23862);
and U24078 (N_24078,N_23785,N_23787);
nand U24079 (N_24079,N_23885,N_23804);
nor U24080 (N_24080,N_23769,N_23973);
xor U24081 (N_24081,N_23952,N_23762);
nor U24082 (N_24082,N_23752,N_23828);
xnor U24083 (N_24083,N_23900,N_23850);
nor U24084 (N_24084,N_23955,N_23974);
or U24085 (N_24085,N_23942,N_23760);
and U24086 (N_24086,N_23920,N_23778);
nor U24087 (N_24087,N_23859,N_23851);
and U24088 (N_24088,N_23876,N_23764);
xnor U24089 (N_24089,N_23777,N_23800);
xor U24090 (N_24090,N_23779,N_23873);
and U24091 (N_24091,N_23864,N_23846);
and U24092 (N_24092,N_23872,N_23848);
xor U24093 (N_24093,N_23926,N_23783);
and U24094 (N_24094,N_23894,N_23968);
nor U24095 (N_24095,N_23790,N_23983);
nor U24096 (N_24096,N_23933,N_23830);
nor U24097 (N_24097,N_23875,N_23928);
nor U24098 (N_24098,N_23948,N_23941);
nand U24099 (N_24099,N_23863,N_23967);
nor U24100 (N_24100,N_23880,N_23975);
nor U24101 (N_24101,N_23815,N_23839);
or U24102 (N_24102,N_23803,N_23860);
and U24103 (N_24103,N_23940,N_23887);
and U24104 (N_24104,N_23889,N_23767);
nand U24105 (N_24105,N_23795,N_23810);
and U24106 (N_24106,N_23776,N_23910);
xor U24107 (N_24107,N_23821,N_23902);
xor U24108 (N_24108,N_23870,N_23761);
nor U24109 (N_24109,N_23977,N_23993);
and U24110 (N_24110,N_23781,N_23847);
or U24111 (N_24111,N_23992,N_23893);
or U24112 (N_24112,N_23854,N_23930);
xor U24113 (N_24113,N_23916,N_23924);
nand U24114 (N_24114,N_23793,N_23852);
nor U24115 (N_24115,N_23818,N_23919);
nor U24116 (N_24116,N_23794,N_23896);
xor U24117 (N_24117,N_23996,N_23999);
or U24118 (N_24118,N_23843,N_23979);
and U24119 (N_24119,N_23831,N_23753);
nor U24120 (N_24120,N_23905,N_23750);
nand U24121 (N_24121,N_23774,N_23918);
nand U24122 (N_24122,N_23995,N_23971);
nor U24123 (N_24123,N_23915,N_23964);
nand U24124 (N_24124,N_23882,N_23799);
nand U24125 (N_24125,N_23857,N_23838);
xnor U24126 (N_24126,N_23760,N_23934);
and U24127 (N_24127,N_23945,N_23782);
nand U24128 (N_24128,N_23857,N_23915);
xnor U24129 (N_24129,N_23758,N_23805);
nor U24130 (N_24130,N_23861,N_23792);
xnor U24131 (N_24131,N_23789,N_23955);
nand U24132 (N_24132,N_23995,N_23938);
nand U24133 (N_24133,N_23990,N_23996);
and U24134 (N_24134,N_23969,N_23935);
and U24135 (N_24135,N_23990,N_23921);
nor U24136 (N_24136,N_23974,N_23798);
nand U24137 (N_24137,N_23821,N_23805);
or U24138 (N_24138,N_23750,N_23777);
and U24139 (N_24139,N_23968,N_23785);
and U24140 (N_24140,N_23846,N_23801);
and U24141 (N_24141,N_23756,N_23991);
and U24142 (N_24142,N_23912,N_23921);
nor U24143 (N_24143,N_23830,N_23883);
nor U24144 (N_24144,N_23919,N_23996);
nand U24145 (N_24145,N_23998,N_23823);
nor U24146 (N_24146,N_23945,N_23759);
and U24147 (N_24147,N_23991,N_23916);
nand U24148 (N_24148,N_23979,N_23975);
nand U24149 (N_24149,N_23868,N_23992);
and U24150 (N_24150,N_23889,N_23846);
xnor U24151 (N_24151,N_23777,N_23934);
xor U24152 (N_24152,N_23905,N_23783);
nand U24153 (N_24153,N_23980,N_23988);
and U24154 (N_24154,N_23846,N_23854);
nand U24155 (N_24155,N_23835,N_23990);
xnor U24156 (N_24156,N_23816,N_23852);
nor U24157 (N_24157,N_23877,N_23906);
nor U24158 (N_24158,N_23903,N_23963);
nor U24159 (N_24159,N_23998,N_23979);
and U24160 (N_24160,N_23789,N_23935);
nor U24161 (N_24161,N_23773,N_23953);
nand U24162 (N_24162,N_23972,N_23936);
xnor U24163 (N_24163,N_23826,N_23977);
nor U24164 (N_24164,N_23915,N_23755);
nand U24165 (N_24165,N_23937,N_23907);
nor U24166 (N_24166,N_23828,N_23949);
nand U24167 (N_24167,N_23998,N_23888);
nor U24168 (N_24168,N_23896,N_23952);
or U24169 (N_24169,N_23872,N_23904);
or U24170 (N_24170,N_23757,N_23952);
nand U24171 (N_24171,N_23912,N_23908);
and U24172 (N_24172,N_23915,N_23820);
and U24173 (N_24173,N_23801,N_23827);
xnor U24174 (N_24174,N_23984,N_23831);
and U24175 (N_24175,N_23968,N_23986);
and U24176 (N_24176,N_23799,N_23999);
nor U24177 (N_24177,N_23933,N_23977);
and U24178 (N_24178,N_23873,N_23986);
xor U24179 (N_24179,N_23847,N_23793);
nor U24180 (N_24180,N_23892,N_23879);
or U24181 (N_24181,N_23995,N_23887);
xor U24182 (N_24182,N_23751,N_23941);
xor U24183 (N_24183,N_23934,N_23874);
or U24184 (N_24184,N_23962,N_23972);
nand U24185 (N_24185,N_23973,N_23761);
nor U24186 (N_24186,N_23757,N_23880);
or U24187 (N_24187,N_23820,N_23882);
or U24188 (N_24188,N_23799,N_23991);
nand U24189 (N_24189,N_23936,N_23756);
and U24190 (N_24190,N_23971,N_23852);
or U24191 (N_24191,N_23908,N_23922);
nor U24192 (N_24192,N_23941,N_23942);
xor U24193 (N_24193,N_23770,N_23771);
and U24194 (N_24194,N_23846,N_23832);
and U24195 (N_24195,N_23857,N_23858);
xnor U24196 (N_24196,N_23766,N_23843);
xnor U24197 (N_24197,N_23864,N_23902);
and U24198 (N_24198,N_23904,N_23785);
nor U24199 (N_24199,N_23881,N_23821);
and U24200 (N_24200,N_23882,N_23911);
or U24201 (N_24201,N_23809,N_23924);
and U24202 (N_24202,N_23991,N_23944);
and U24203 (N_24203,N_23940,N_23955);
or U24204 (N_24204,N_23804,N_23893);
or U24205 (N_24205,N_23803,N_23788);
nor U24206 (N_24206,N_23937,N_23888);
or U24207 (N_24207,N_23801,N_23809);
xnor U24208 (N_24208,N_23757,N_23762);
xnor U24209 (N_24209,N_23892,N_23973);
xnor U24210 (N_24210,N_23902,N_23778);
and U24211 (N_24211,N_23852,N_23978);
nor U24212 (N_24212,N_23817,N_23819);
nor U24213 (N_24213,N_23851,N_23870);
nand U24214 (N_24214,N_23816,N_23930);
or U24215 (N_24215,N_23891,N_23845);
or U24216 (N_24216,N_23921,N_23966);
xor U24217 (N_24217,N_23929,N_23935);
xor U24218 (N_24218,N_23922,N_23944);
nor U24219 (N_24219,N_23907,N_23888);
nor U24220 (N_24220,N_23770,N_23959);
nand U24221 (N_24221,N_23803,N_23804);
nand U24222 (N_24222,N_23843,N_23886);
and U24223 (N_24223,N_23806,N_23932);
or U24224 (N_24224,N_23809,N_23926);
and U24225 (N_24225,N_23811,N_23797);
and U24226 (N_24226,N_23886,N_23798);
or U24227 (N_24227,N_23850,N_23997);
and U24228 (N_24228,N_23885,N_23972);
nand U24229 (N_24229,N_23883,N_23957);
nand U24230 (N_24230,N_23787,N_23751);
or U24231 (N_24231,N_23987,N_23979);
nor U24232 (N_24232,N_23831,N_23915);
or U24233 (N_24233,N_23939,N_23757);
xnor U24234 (N_24234,N_23838,N_23877);
and U24235 (N_24235,N_23919,N_23879);
nand U24236 (N_24236,N_23994,N_23836);
nand U24237 (N_24237,N_23935,N_23802);
nand U24238 (N_24238,N_23980,N_23839);
and U24239 (N_24239,N_23986,N_23764);
nand U24240 (N_24240,N_23838,N_23774);
xnor U24241 (N_24241,N_23980,N_23914);
nor U24242 (N_24242,N_23858,N_23947);
xor U24243 (N_24243,N_23834,N_23970);
and U24244 (N_24244,N_23898,N_23774);
and U24245 (N_24245,N_23922,N_23966);
or U24246 (N_24246,N_23964,N_23761);
or U24247 (N_24247,N_23925,N_23987);
and U24248 (N_24248,N_23975,N_23850);
xor U24249 (N_24249,N_23751,N_23802);
nand U24250 (N_24250,N_24133,N_24234);
nand U24251 (N_24251,N_24237,N_24117);
and U24252 (N_24252,N_24127,N_24174);
nor U24253 (N_24253,N_24111,N_24031);
and U24254 (N_24254,N_24204,N_24130);
nand U24255 (N_24255,N_24226,N_24187);
and U24256 (N_24256,N_24015,N_24057);
nor U24257 (N_24257,N_24188,N_24243);
xor U24258 (N_24258,N_24036,N_24217);
and U24259 (N_24259,N_24136,N_24148);
nand U24260 (N_24260,N_24227,N_24153);
nor U24261 (N_24261,N_24207,N_24211);
or U24262 (N_24262,N_24165,N_24197);
and U24263 (N_24263,N_24103,N_24132);
and U24264 (N_24264,N_24236,N_24199);
nor U24265 (N_24265,N_24116,N_24068);
or U24266 (N_24266,N_24198,N_24152);
xnor U24267 (N_24267,N_24105,N_24107);
nor U24268 (N_24268,N_24151,N_24225);
or U24269 (N_24269,N_24060,N_24238);
nor U24270 (N_24270,N_24195,N_24135);
xor U24271 (N_24271,N_24046,N_24129);
nor U24272 (N_24272,N_24182,N_24119);
and U24273 (N_24273,N_24069,N_24037);
or U24274 (N_24274,N_24168,N_24051);
and U24275 (N_24275,N_24139,N_24058);
nor U24276 (N_24276,N_24097,N_24241);
and U24277 (N_24277,N_24173,N_24170);
xnor U24278 (N_24278,N_24229,N_24184);
and U24279 (N_24279,N_24172,N_24162);
xor U24280 (N_24280,N_24218,N_24150);
nor U24281 (N_24281,N_24179,N_24235);
and U24282 (N_24282,N_24099,N_24002);
nand U24283 (N_24283,N_24093,N_24221);
or U24284 (N_24284,N_24045,N_24164);
or U24285 (N_24285,N_24048,N_24144);
nor U24286 (N_24286,N_24194,N_24185);
xor U24287 (N_24287,N_24055,N_24134);
xnor U24288 (N_24288,N_24191,N_24034);
nor U24289 (N_24289,N_24160,N_24104);
and U24290 (N_24290,N_24131,N_24120);
nor U24291 (N_24291,N_24040,N_24176);
nor U24292 (N_24292,N_24155,N_24163);
and U24293 (N_24293,N_24159,N_24074);
xor U24294 (N_24294,N_24017,N_24233);
nand U24295 (N_24295,N_24027,N_24011);
xnor U24296 (N_24296,N_24248,N_24030);
or U24297 (N_24297,N_24113,N_24213);
nand U24298 (N_24298,N_24154,N_24244);
and U24299 (N_24299,N_24047,N_24149);
or U24300 (N_24300,N_24114,N_24026);
nand U24301 (N_24301,N_24115,N_24169);
nor U24302 (N_24302,N_24084,N_24088);
xnor U24303 (N_24303,N_24006,N_24092);
nor U24304 (N_24304,N_24073,N_24110);
or U24305 (N_24305,N_24004,N_24224);
or U24306 (N_24306,N_24039,N_24106);
xnor U24307 (N_24307,N_24087,N_24021);
nand U24308 (N_24308,N_24167,N_24052);
nor U24309 (N_24309,N_24222,N_24050);
nor U24310 (N_24310,N_24071,N_24007);
or U24311 (N_24311,N_24090,N_24189);
and U24312 (N_24312,N_24082,N_24018);
xor U24313 (N_24313,N_24076,N_24249);
nand U24314 (N_24314,N_24231,N_24041);
or U24315 (N_24315,N_24064,N_24146);
xnor U24316 (N_24316,N_24206,N_24178);
nor U24317 (N_24317,N_24141,N_24008);
nor U24318 (N_24318,N_24022,N_24067);
nor U24319 (N_24319,N_24118,N_24247);
or U24320 (N_24320,N_24038,N_24072);
xnor U24321 (N_24321,N_24035,N_24020);
or U24322 (N_24322,N_24245,N_24053);
xor U24323 (N_24323,N_24089,N_24019);
and U24324 (N_24324,N_24059,N_24016);
nand U24325 (N_24325,N_24212,N_24142);
nor U24326 (N_24326,N_24230,N_24081);
or U24327 (N_24327,N_24171,N_24123);
nand U24328 (N_24328,N_24056,N_24078);
and U24329 (N_24329,N_24000,N_24175);
and U24330 (N_24330,N_24080,N_24143);
or U24331 (N_24331,N_24096,N_24102);
nor U24332 (N_24332,N_24158,N_24137);
nand U24333 (N_24333,N_24219,N_24042);
nor U24334 (N_24334,N_24140,N_24216);
xnor U24335 (N_24335,N_24192,N_24086);
nor U24336 (N_24336,N_24201,N_24023);
and U24337 (N_24337,N_24065,N_24083);
xnor U24338 (N_24338,N_24091,N_24145);
xnor U24339 (N_24339,N_24101,N_24157);
nor U24340 (N_24340,N_24240,N_24215);
nor U24341 (N_24341,N_24070,N_24125);
nor U24342 (N_24342,N_24239,N_24196);
nand U24343 (N_24343,N_24112,N_24223);
xnor U24344 (N_24344,N_24025,N_24161);
nor U24345 (N_24345,N_24109,N_24009);
or U24346 (N_24346,N_24177,N_24200);
nand U24347 (N_24347,N_24094,N_24032);
and U24348 (N_24348,N_24063,N_24180);
and U24349 (N_24349,N_24012,N_24066);
and U24350 (N_24350,N_24193,N_24054);
nand U24351 (N_24351,N_24095,N_24075);
nand U24352 (N_24352,N_24181,N_24098);
xnor U24353 (N_24353,N_24203,N_24029);
nor U24354 (N_24354,N_24079,N_24003);
xnor U24355 (N_24355,N_24156,N_24138);
nor U24356 (N_24356,N_24005,N_24043);
and U24357 (N_24357,N_24077,N_24033);
nand U24358 (N_24358,N_24242,N_24014);
nand U24359 (N_24359,N_24220,N_24190);
or U24360 (N_24360,N_24209,N_24202);
and U24361 (N_24361,N_24124,N_24166);
nor U24362 (N_24362,N_24013,N_24214);
nor U24363 (N_24363,N_24121,N_24186);
xnor U24364 (N_24364,N_24024,N_24205);
nor U24365 (N_24365,N_24044,N_24183);
or U24366 (N_24366,N_24126,N_24147);
nor U24367 (N_24367,N_24085,N_24100);
nor U24368 (N_24368,N_24228,N_24246);
and U24369 (N_24369,N_24010,N_24062);
and U24370 (N_24370,N_24061,N_24001);
or U24371 (N_24371,N_24208,N_24210);
nor U24372 (N_24372,N_24128,N_24049);
nor U24373 (N_24373,N_24028,N_24108);
and U24374 (N_24374,N_24232,N_24122);
nor U24375 (N_24375,N_24103,N_24010);
xnor U24376 (N_24376,N_24171,N_24202);
or U24377 (N_24377,N_24031,N_24055);
nand U24378 (N_24378,N_24082,N_24102);
xnor U24379 (N_24379,N_24113,N_24169);
nor U24380 (N_24380,N_24046,N_24048);
xor U24381 (N_24381,N_24101,N_24206);
xnor U24382 (N_24382,N_24126,N_24188);
and U24383 (N_24383,N_24243,N_24153);
nand U24384 (N_24384,N_24148,N_24187);
xnor U24385 (N_24385,N_24150,N_24199);
xor U24386 (N_24386,N_24244,N_24185);
nor U24387 (N_24387,N_24230,N_24196);
xor U24388 (N_24388,N_24004,N_24068);
or U24389 (N_24389,N_24078,N_24114);
or U24390 (N_24390,N_24225,N_24100);
or U24391 (N_24391,N_24159,N_24140);
xor U24392 (N_24392,N_24029,N_24026);
nand U24393 (N_24393,N_24199,N_24054);
nor U24394 (N_24394,N_24237,N_24073);
and U24395 (N_24395,N_24195,N_24030);
and U24396 (N_24396,N_24052,N_24223);
or U24397 (N_24397,N_24174,N_24060);
nand U24398 (N_24398,N_24240,N_24078);
nor U24399 (N_24399,N_24109,N_24161);
or U24400 (N_24400,N_24204,N_24119);
xnor U24401 (N_24401,N_24231,N_24158);
nor U24402 (N_24402,N_24204,N_24241);
and U24403 (N_24403,N_24054,N_24013);
nand U24404 (N_24404,N_24158,N_24047);
xnor U24405 (N_24405,N_24096,N_24101);
nand U24406 (N_24406,N_24157,N_24172);
and U24407 (N_24407,N_24190,N_24243);
or U24408 (N_24408,N_24141,N_24094);
nand U24409 (N_24409,N_24158,N_24006);
nand U24410 (N_24410,N_24174,N_24005);
nor U24411 (N_24411,N_24161,N_24246);
xnor U24412 (N_24412,N_24067,N_24072);
nor U24413 (N_24413,N_24192,N_24170);
nor U24414 (N_24414,N_24225,N_24007);
or U24415 (N_24415,N_24023,N_24076);
xor U24416 (N_24416,N_24212,N_24078);
xnor U24417 (N_24417,N_24041,N_24146);
nor U24418 (N_24418,N_24070,N_24186);
or U24419 (N_24419,N_24191,N_24228);
nor U24420 (N_24420,N_24243,N_24072);
nand U24421 (N_24421,N_24083,N_24085);
and U24422 (N_24422,N_24075,N_24160);
xor U24423 (N_24423,N_24069,N_24204);
nor U24424 (N_24424,N_24098,N_24045);
nand U24425 (N_24425,N_24210,N_24063);
and U24426 (N_24426,N_24051,N_24212);
nand U24427 (N_24427,N_24097,N_24099);
and U24428 (N_24428,N_24173,N_24208);
and U24429 (N_24429,N_24129,N_24071);
nor U24430 (N_24430,N_24219,N_24068);
and U24431 (N_24431,N_24171,N_24165);
nand U24432 (N_24432,N_24203,N_24155);
nor U24433 (N_24433,N_24150,N_24243);
and U24434 (N_24434,N_24055,N_24205);
or U24435 (N_24435,N_24128,N_24002);
xor U24436 (N_24436,N_24075,N_24073);
and U24437 (N_24437,N_24176,N_24170);
or U24438 (N_24438,N_24230,N_24002);
nand U24439 (N_24439,N_24150,N_24249);
xnor U24440 (N_24440,N_24128,N_24178);
nor U24441 (N_24441,N_24030,N_24104);
nor U24442 (N_24442,N_24177,N_24203);
nand U24443 (N_24443,N_24216,N_24008);
xor U24444 (N_24444,N_24038,N_24010);
nor U24445 (N_24445,N_24133,N_24210);
xor U24446 (N_24446,N_24144,N_24070);
and U24447 (N_24447,N_24218,N_24010);
nand U24448 (N_24448,N_24135,N_24120);
xor U24449 (N_24449,N_24029,N_24018);
xor U24450 (N_24450,N_24115,N_24082);
and U24451 (N_24451,N_24174,N_24230);
nand U24452 (N_24452,N_24151,N_24072);
nand U24453 (N_24453,N_24010,N_24226);
nand U24454 (N_24454,N_24137,N_24139);
and U24455 (N_24455,N_24174,N_24024);
and U24456 (N_24456,N_24020,N_24246);
nor U24457 (N_24457,N_24075,N_24210);
nand U24458 (N_24458,N_24114,N_24232);
and U24459 (N_24459,N_24074,N_24228);
and U24460 (N_24460,N_24203,N_24017);
nor U24461 (N_24461,N_24079,N_24210);
and U24462 (N_24462,N_24150,N_24101);
nand U24463 (N_24463,N_24015,N_24138);
nor U24464 (N_24464,N_24157,N_24008);
xor U24465 (N_24465,N_24070,N_24167);
and U24466 (N_24466,N_24205,N_24100);
xor U24467 (N_24467,N_24145,N_24061);
or U24468 (N_24468,N_24207,N_24026);
nand U24469 (N_24469,N_24101,N_24215);
or U24470 (N_24470,N_24226,N_24055);
nand U24471 (N_24471,N_24022,N_24085);
nor U24472 (N_24472,N_24165,N_24040);
nor U24473 (N_24473,N_24102,N_24208);
and U24474 (N_24474,N_24044,N_24094);
xnor U24475 (N_24475,N_24217,N_24224);
xor U24476 (N_24476,N_24175,N_24017);
or U24477 (N_24477,N_24195,N_24044);
xnor U24478 (N_24478,N_24204,N_24118);
and U24479 (N_24479,N_24152,N_24246);
xnor U24480 (N_24480,N_24197,N_24154);
xnor U24481 (N_24481,N_24052,N_24214);
or U24482 (N_24482,N_24026,N_24116);
or U24483 (N_24483,N_24141,N_24181);
nor U24484 (N_24484,N_24152,N_24098);
or U24485 (N_24485,N_24201,N_24237);
or U24486 (N_24486,N_24161,N_24057);
and U24487 (N_24487,N_24090,N_24186);
nor U24488 (N_24488,N_24005,N_24216);
and U24489 (N_24489,N_24191,N_24160);
or U24490 (N_24490,N_24107,N_24145);
and U24491 (N_24491,N_24182,N_24165);
and U24492 (N_24492,N_24146,N_24135);
xor U24493 (N_24493,N_24214,N_24047);
nand U24494 (N_24494,N_24223,N_24178);
and U24495 (N_24495,N_24029,N_24073);
or U24496 (N_24496,N_24040,N_24230);
xor U24497 (N_24497,N_24215,N_24199);
or U24498 (N_24498,N_24226,N_24016);
nand U24499 (N_24499,N_24130,N_24189);
nor U24500 (N_24500,N_24295,N_24258);
or U24501 (N_24501,N_24443,N_24406);
xnor U24502 (N_24502,N_24446,N_24429);
nor U24503 (N_24503,N_24250,N_24297);
nor U24504 (N_24504,N_24308,N_24356);
xnor U24505 (N_24505,N_24372,N_24405);
and U24506 (N_24506,N_24296,N_24408);
and U24507 (N_24507,N_24418,N_24457);
nor U24508 (N_24508,N_24345,N_24404);
xnor U24509 (N_24509,N_24423,N_24419);
nor U24510 (N_24510,N_24427,N_24390);
nand U24511 (N_24511,N_24333,N_24257);
and U24512 (N_24512,N_24319,N_24277);
nor U24513 (N_24513,N_24410,N_24252);
and U24514 (N_24514,N_24301,N_24344);
xnor U24515 (N_24515,N_24342,N_24335);
and U24516 (N_24516,N_24328,N_24445);
and U24517 (N_24517,N_24411,N_24477);
or U24518 (N_24518,N_24417,N_24306);
xor U24519 (N_24519,N_24375,N_24310);
nand U24520 (N_24520,N_24462,N_24331);
xnor U24521 (N_24521,N_24458,N_24270);
nor U24522 (N_24522,N_24413,N_24321);
or U24523 (N_24523,N_24431,N_24275);
and U24524 (N_24524,N_24386,N_24320);
xor U24525 (N_24525,N_24298,N_24414);
xor U24526 (N_24526,N_24271,N_24438);
nor U24527 (N_24527,N_24343,N_24387);
xor U24528 (N_24528,N_24430,N_24453);
or U24529 (N_24529,N_24373,N_24447);
nor U24530 (N_24530,N_24360,N_24384);
nor U24531 (N_24531,N_24374,N_24439);
nand U24532 (N_24532,N_24434,N_24341);
xnor U24533 (N_24533,N_24269,N_24428);
nand U24534 (N_24534,N_24440,N_24426);
and U24535 (N_24535,N_24432,N_24388);
xor U24536 (N_24536,N_24397,N_24288);
nand U24537 (N_24537,N_24379,N_24391);
nor U24538 (N_24538,N_24363,N_24433);
nand U24539 (N_24539,N_24484,N_24347);
or U24540 (N_24540,N_24272,N_24476);
nand U24541 (N_24541,N_24309,N_24380);
xnor U24542 (N_24542,N_24293,N_24437);
or U24543 (N_24543,N_24381,N_24354);
nor U24544 (N_24544,N_24496,N_24461);
xnor U24545 (N_24545,N_24316,N_24273);
nand U24546 (N_24546,N_24339,N_24268);
or U24547 (N_24547,N_24359,N_24338);
and U24548 (N_24548,N_24290,N_24324);
nand U24549 (N_24549,N_24256,N_24471);
nor U24550 (N_24550,N_24448,N_24402);
and U24551 (N_24551,N_24479,N_24409);
and U24552 (N_24552,N_24464,N_24436);
and U24553 (N_24553,N_24489,N_24400);
xnor U24554 (N_24554,N_24393,N_24420);
nand U24555 (N_24555,N_24425,N_24463);
or U24556 (N_24556,N_24253,N_24382);
nor U24557 (N_24557,N_24498,N_24467);
or U24558 (N_24558,N_24486,N_24480);
nor U24559 (N_24559,N_24281,N_24395);
xor U24560 (N_24560,N_24412,N_24455);
xor U24561 (N_24561,N_24350,N_24399);
and U24562 (N_24562,N_24473,N_24492);
xnor U24563 (N_24563,N_24407,N_24355);
nor U24564 (N_24564,N_24318,N_24483);
nor U24565 (N_24565,N_24452,N_24470);
xor U24566 (N_24566,N_24365,N_24317);
xor U24567 (N_24567,N_24330,N_24394);
nand U24568 (N_24568,N_24368,N_24322);
nor U24569 (N_24569,N_24361,N_24259);
nor U24570 (N_24570,N_24351,N_24282);
nand U24571 (N_24571,N_24422,N_24424);
xnor U24572 (N_24572,N_24370,N_24261);
and U24573 (N_24573,N_24490,N_24307);
xnor U24574 (N_24574,N_24475,N_24329);
or U24575 (N_24575,N_24495,N_24286);
xor U24576 (N_24576,N_24255,N_24442);
or U24577 (N_24577,N_24332,N_24369);
nor U24578 (N_24578,N_24289,N_24346);
nor U24579 (N_24579,N_24334,N_24357);
xor U24580 (N_24580,N_24260,N_24274);
xor U24581 (N_24581,N_24254,N_24352);
nor U24582 (N_24582,N_24469,N_24266);
xor U24583 (N_24583,N_24450,N_24385);
nand U24584 (N_24584,N_24314,N_24481);
or U24585 (N_24585,N_24313,N_24403);
nor U24586 (N_24586,N_24494,N_24364);
and U24587 (N_24587,N_24302,N_24396);
and U24588 (N_24588,N_24264,N_24465);
nor U24589 (N_24589,N_24284,N_24336);
nand U24590 (N_24590,N_24358,N_24415);
nor U24591 (N_24591,N_24327,N_24299);
nand U24592 (N_24592,N_24367,N_24278);
and U24593 (N_24593,N_24466,N_24305);
xor U24594 (N_24594,N_24392,N_24449);
or U24595 (N_24595,N_24340,N_24383);
nor U24596 (N_24596,N_24472,N_24487);
and U24597 (N_24597,N_24315,N_24497);
nand U24598 (N_24598,N_24416,N_24294);
nor U24599 (N_24599,N_24323,N_24499);
and U24600 (N_24600,N_24371,N_24304);
and U24601 (N_24601,N_24468,N_24325);
xor U24602 (N_24602,N_24267,N_24389);
or U24603 (N_24603,N_24362,N_24456);
or U24604 (N_24604,N_24353,N_24312);
and U24605 (N_24605,N_24482,N_24493);
or U24606 (N_24606,N_24376,N_24444);
nand U24607 (N_24607,N_24348,N_24292);
or U24608 (N_24608,N_24276,N_24377);
nand U24609 (N_24609,N_24285,N_24279);
or U24610 (N_24610,N_24441,N_24251);
or U24611 (N_24611,N_24488,N_24265);
or U24612 (N_24612,N_24349,N_24263);
xnor U24613 (N_24613,N_24326,N_24485);
nand U24614 (N_24614,N_24421,N_24491);
and U24615 (N_24615,N_24280,N_24454);
nor U24616 (N_24616,N_24459,N_24478);
xnor U24617 (N_24617,N_24451,N_24311);
and U24618 (N_24618,N_24398,N_24283);
and U24619 (N_24619,N_24401,N_24291);
nand U24620 (N_24620,N_24337,N_24303);
or U24621 (N_24621,N_24262,N_24474);
nor U24622 (N_24622,N_24287,N_24435);
xor U24623 (N_24623,N_24366,N_24300);
nand U24624 (N_24624,N_24460,N_24378);
nor U24625 (N_24625,N_24317,N_24419);
xnor U24626 (N_24626,N_24250,N_24301);
nand U24627 (N_24627,N_24304,N_24470);
nand U24628 (N_24628,N_24415,N_24351);
xor U24629 (N_24629,N_24289,N_24401);
nand U24630 (N_24630,N_24311,N_24256);
xor U24631 (N_24631,N_24353,N_24433);
xnor U24632 (N_24632,N_24404,N_24472);
nor U24633 (N_24633,N_24374,N_24481);
or U24634 (N_24634,N_24390,N_24267);
nor U24635 (N_24635,N_24293,N_24454);
xor U24636 (N_24636,N_24384,N_24336);
nand U24637 (N_24637,N_24340,N_24252);
or U24638 (N_24638,N_24332,N_24450);
and U24639 (N_24639,N_24423,N_24356);
xor U24640 (N_24640,N_24441,N_24324);
xor U24641 (N_24641,N_24252,N_24470);
nand U24642 (N_24642,N_24289,N_24292);
or U24643 (N_24643,N_24251,N_24453);
or U24644 (N_24644,N_24353,N_24488);
or U24645 (N_24645,N_24411,N_24387);
xnor U24646 (N_24646,N_24469,N_24490);
nor U24647 (N_24647,N_24489,N_24458);
nor U24648 (N_24648,N_24331,N_24436);
xor U24649 (N_24649,N_24352,N_24347);
nor U24650 (N_24650,N_24337,N_24387);
or U24651 (N_24651,N_24258,N_24275);
nor U24652 (N_24652,N_24388,N_24494);
nor U24653 (N_24653,N_24406,N_24433);
nand U24654 (N_24654,N_24319,N_24406);
nand U24655 (N_24655,N_24401,N_24468);
xnor U24656 (N_24656,N_24266,N_24305);
nor U24657 (N_24657,N_24285,N_24387);
and U24658 (N_24658,N_24358,N_24435);
nor U24659 (N_24659,N_24472,N_24412);
or U24660 (N_24660,N_24253,N_24266);
and U24661 (N_24661,N_24479,N_24338);
and U24662 (N_24662,N_24296,N_24307);
nand U24663 (N_24663,N_24357,N_24448);
nand U24664 (N_24664,N_24421,N_24305);
nand U24665 (N_24665,N_24428,N_24255);
and U24666 (N_24666,N_24352,N_24415);
xor U24667 (N_24667,N_24343,N_24355);
xor U24668 (N_24668,N_24458,N_24356);
nor U24669 (N_24669,N_24278,N_24454);
or U24670 (N_24670,N_24370,N_24398);
nor U24671 (N_24671,N_24368,N_24413);
xnor U24672 (N_24672,N_24376,N_24445);
nand U24673 (N_24673,N_24396,N_24468);
or U24674 (N_24674,N_24415,N_24280);
xnor U24675 (N_24675,N_24304,N_24319);
nand U24676 (N_24676,N_24309,N_24406);
or U24677 (N_24677,N_24339,N_24464);
and U24678 (N_24678,N_24422,N_24284);
and U24679 (N_24679,N_24361,N_24354);
nand U24680 (N_24680,N_24333,N_24277);
or U24681 (N_24681,N_24306,N_24484);
nand U24682 (N_24682,N_24459,N_24269);
and U24683 (N_24683,N_24432,N_24253);
nor U24684 (N_24684,N_24463,N_24451);
xor U24685 (N_24685,N_24307,N_24458);
nand U24686 (N_24686,N_24334,N_24377);
and U24687 (N_24687,N_24321,N_24391);
nand U24688 (N_24688,N_24397,N_24451);
xor U24689 (N_24689,N_24484,N_24313);
and U24690 (N_24690,N_24391,N_24353);
and U24691 (N_24691,N_24410,N_24284);
or U24692 (N_24692,N_24451,N_24303);
nor U24693 (N_24693,N_24485,N_24468);
or U24694 (N_24694,N_24276,N_24410);
and U24695 (N_24695,N_24391,N_24493);
and U24696 (N_24696,N_24377,N_24347);
and U24697 (N_24697,N_24396,N_24368);
and U24698 (N_24698,N_24293,N_24261);
xnor U24699 (N_24699,N_24318,N_24419);
nor U24700 (N_24700,N_24362,N_24495);
nor U24701 (N_24701,N_24499,N_24489);
nor U24702 (N_24702,N_24478,N_24449);
nor U24703 (N_24703,N_24328,N_24257);
xnor U24704 (N_24704,N_24310,N_24332);
xor U24705 (N_24705,N_24461,N_24382);
xnor U24706 (N_24706,N_24357,N_24408);
or U24707 (N_24707,N_24350,N_24375);
nor U24708 (N_24708,N_24316,N_24314);
nand U24709 (N_24709,N_24422,N_24363);
nor U24710 (N_24710,N_24493,N_24472);
nor U24711 (N_24711,N_24332,N_24425);
or U24712 (N_24712,N_24320,N_24290);
nand U24713 (N_24713,N_24296,N_24471);
or U24714 (N_24714,N_24489,N_24358);
xor U24715 (N_24715,N_24399,N_24309);
or U24716 (N_24716,N_24450,N_24454);
or U24717 (N_24717,N_24309,N_24376);
and U24718 (N_24718,N_24347,N_24345);
nor U24719 (N_24719,N_24464,N_24301);
xor U24720 (N_24720,N_24484,N_24499);
and U24721 (N_24721,N_24330,N_24375);
and U24722 (N_24722,N_24260,N_24312);
nor U24723 (N_24723,N_24344,N_24348);
or U24724 (N_24724,N_24266,N_24361);
or U24725 (N_24725,N_24365,N_24342);
nor U24726 (N_24726,N_24473,N_24324);
xnor U24727 (N_24727,N_24446,N_24271);
nand U24728 (N_24728,N_24386,N_24384);
xor U24729 (N_24729,N_24451,N_24328);
nor U24730 (N_24730,N_24318,N_24458);
nor U24731 (N_24731,N_24343,N_24468);
xnor U24732 (N_24732,N_24371,N_24390);
nor U24733 (N_24733,N_24293,N_24287);
and U24734 (N_24734,N_24344,N_24399);
nand U24735 (N_24735,N_24289,N_24322);
or U24736 (N_24736,N_24365,N_24448);
and U24737 (N_24737,N_24380,N_24441);
nand U24738 (N_24738,N_24381,N_24461);
nor U24739 (N_24739,N_24286,N_24418);
and U24740 (N_24740,N_24361,N_24309);
nor U24741 (N_24741,N_24282,N_24477);
xnor U24742 (N_24742,N_24276,N_24266);
or U24743 (N_24743,N_24364,N_24410);
nor U24744 (N_24744,N_24493,N_24392);
nand U24745 (N_24745,N_24445,N_24327);
or U24746 (N_24746,N_24429,N_24370);
xnor U24747 (N_24747,N_24368,N_24430);
xor U24748 (N_24748,N_24360,N_24434);
or U24749 (N_24749,N_24344,N_24390);
nand U24750 (N_24750,N_24653,N_24643);
or U24751 (N_24751,N_24713,N_24699);
nand U24752 (N_24752,N_24675,N_24531);
or U24753 (N_24753,N_24605,N_24682);
xor U24754 (N_24754,N_24632,N_24690);
and U24755 (N_24755,N_24734,N_24545);
nor U24756 (N_24756,N_24728,N_24748);
nor U24757 (N_24757,N_24564,N_24615);
and U24758 (N_24758,N_24530,N_24647);
xor U24759 (N_24759,N_24667,N_24627);
nand U24760 (N_24760,N_24689,N_24716);
nor U24761 (N_24761,N_24617,N_24718);
xor U24762 (N_24762,N_24630,N_24614);
xnor U24763 (N_24763,N_24612,N_24591);
or U24764 (N_24764,N_24693,N_24518);
or U24765 (N_24765,N_24576,N_24648);
xnor U24766 (N_24766,N_24574,N_24727);
and U24767 (N_24767,N_24532,N_24662);
nand U24768 (N_24768,N_24657,N_24714);
nand U24769 (N_24769,N_24580,N_24598);
and U24770 (N_24770,N_24676,N_24705);
and U24771 (N_24771,N_24749,N_24746);
or U24772 (N_24772,N_24568,N_24551);
and U24773 (N_24773,N_24700,N_24587);
and U24774 (N_24774,N_24540,N_24514);
nor U24775 (N_24775,N_24725,N_24679);
nor U24776 (N_24776,N_24560,N_24650);
xor U24777 (N_24777,N_24595,N_24736);
or U24778 (N_24778,N_24557,N_24507);
xor U24779 (N_24779,N_24552,N_24570);
or U24780 (N_24780,N_24542,N_24571);
or U24781 (N_24781,N_24585,N_24606);
nand U24782 (N_24782,N_24747,N_24546);
nand U24783 (N_24783,N_24593,N_24745);
nor U24784 (N_24784,N_24509,N_24629);
or U24785 (N_24785,N_24715,N_24502);
xor U24786 (N_24786,N_24534,N_24674);
nor U24787 (N_24787,N_24601,N_24695);
or U24788 (N_24788,N_24688,N_24516);
xnor U24789 (N_24789,N_24673,N_24635);
xor U24790 (N_24790,N_24521,N_24735);
nor U24791 (N_24791,N_24537,N_24651);
nor U24792 (N_24792,N_24737,N_24535);
nor U24793 (N_24793,N_24589,N_24661);
nand U24794 (N_24794,N_24555,N_24645);
xnor U24795 (N_24795,N_24513,N_24548);
nor U24796 (N_24796,N_24584,N_24694);
and U24797 (N_24797,N_24500,N_24594);
or U24798 (N_24798,N_24581,N_24644);
or U24799 (N_24799,N_24739,N_24708);
and U24800 (N_24800,N_24710,N_24603);
nand U24801 (N_24801,N_24717,N_24741);
xor U24802 (N_24802,N_24563,N_24697);
xnor U24803 (N_24803,N_24637,N_24670);
nor U24804 (N_24804,N_24533,N_24515);
nand U24805 (N_24805,N_24554,N_24719);
and U24806 (N_24806,N_24658,N_24639);
xnor U24807 (N_24807,N_24720,N_24582);
or U24808 (N_24808,N_24611,N_24501);
nand U24809 (N_24809,N_24671,N_24733);
nor U24810 (N_24810,N_24660,N_24562);
or U24811 (N_24811,N_24659,N_24723);
nand U24812 (N_24812,N_24698,N_24701);
nor U24813 (N_24813,N_24742,N_24663);
or U24814 (N_24814,N_24579,N_24613);
or U24815 (N_24815,N_24649,N_24508);
or U24816 (N_24816,N_24628,N_24622);
nor U24817 (N_24817,N_24512,N_24590);
xor U24818 (N_24818,N_24567,N_24634);
or U24819 (N_24819,N_24536,N_24550);
and U24820 (N_24820,N_24656,N_24619);
xor U24821 (N_24821,N_24706,N_24510);
nor U24822 (N_24822,N_24683,N_24556);
xnor U24823 (N_24823,N_24711,N_24607);
or U24824 (N_24824,N_24517,N_24539);
or U24825 (N_24825,N_24633,N_24588);
or U24826 (N_24826,N_24621,N_24505);
nor U24827 (N_24827,N_24573,N_24636);
and U24828 (N_24828,N_24744,N_24526);
xor U24829 (N_24829,N_24666,N_24704);
or U24830 (N_24830,N_24602,N_24609);
nand U24831 (N_24831,N_24655,N_24709);
nor U24832 (N_24832,N_24559,N_24672);
and U24833 (N_24833,N_24642,N_24712);
and U24834 (N_24834,N_24677,N_24641);
or U24835 (N_24835,N_24575,N_24681);
nand U24836 (N_24836,N_24625,N_24523);
or U24837 (N_24837,N_24566,N_24616);
nand U24838 (N_24838,N_24525,N_24558);
or U24839 (N_24839,N_24553,N_24604);
xor U24840 (N_24840,N_24686,N_24731);
or U24841 (N_24841,N_24569,N_24572);
xor U24842 (N_24842,N_24743,N_24583);
or U24843 (N_24843,N_24726,N_24664);
and U24844 (N_24844,N_24524,N_24600);
nor U24845 (N_24845,N_24610,N_24565);
nor U24846 (N_24846,N_24538,N_24687);
and U24847 (N_24847,N_24652,N_24640);
and U24848 (N_24848,N_24646,N_24597);
and U24849 (N_24849,N_24623,N_24586);
or U24850 (N_24850,N_24680,N_24504);
nand U24851 (N_24851,N_24503,N_24618);
nor U24852 (N_24852,N_24577,N_24654);
xnor U24853 (N_24853,N_24620,N_24678);
or U24854 (N_24854,N_24626,N_24543);
nand U24855 (N_24855,N_24520,N_24738);
or U24856 (N_24856,N_24696,N_24631);
nor U24857 (N_24857,N_24519,N_24740);
nand U24858 (N_24858,N_24561,N_24665);
xnor U24859 (N_24859,N_24522,N_24599);
or U24860 (N_24860,N_24707,N_24549);
xnor U24861 (N_24861,N_24692,N_24691);
and U24862 (N_24862,N_24528,N_24722);
nor U24863 (N_24863,N_24638,N_24669);
nor U24864 (N_24864,N_24592,N_24684);
xor U24865 (N_24865,N_24721,N_24578);
nor U24866 (N_24866,N_24608,N_24529);
or U24867 (N_24867,N_24527,N_24730);
xor U24868 (N_24868,N_24703,N_24596);
xor U24869 (N_24869,N_24685,N_24729);
nand U24870 (N_24870,N_24511,N_24544);
xnor U24871 (N_24871,N_24732,N_24547);
nand U24872 (N_24872,N_24668,N_24724);
nor U24873 (N_24873,N_24506,N_24624);
or U24874 (N_24874,N_24702,N_24541);
xor U24875 (N_24875,N_24651,N_24506);
or U24876 (N_24876,N_24649,N_24661);
or U24877 (N_24877,N_24572,N_24682);
nand U24878 (N_24878,N_24662,N_24607);
nand U24879 (N_24879,N_24746,N_24521);
xor U24880 (N_24880,N_24638,N_24536);
or U24881 (N_24881,N_24656,N_24726);
or U24882 (N_24882,N_24620,N_24612);
and U24883 (N_24883,N_24650,N_24519);
nand U24884 (N_24884,N_24585,N_24616);
or U24885 (N_24885,N_24581,N_24641);
nand U24886 (N_24886,N_24564,N_24737);
xor U24887 (N_24887,N_24525,N_24550);
xor U24888 (N_24888,N_24593,N_24619);
nor U24889 (N_24889,N_24606,N_24668);
xor U24890 (N_24890,N_24743,N_24519);
xor U24891 (N_24891,N_24524,N_24552);
xor U24892 (N_24892,N_24682,N_24514);
nand U24893 (N_24893,N_24604,N_24501);
or U24894 (N_24894,N_24612,N_24547);
and U24895 (N_24895,N_24741,N_24524);
nor U24896 (N_24896,N_24641,N_24637);
xnor U24897 (N_24897,N_24515,N_24527);
nor U24898 (N_24898,N_24576,N_24563);
or U24899 (N_24899,N_24640,N_24709);
and U24900 (N_24900,N_24609,N_24660);
xnor U24901 (N_24901,N_24592,N_24691);
nand U24902 (N_24902,N_24584,N_24718);
or U24903 (N_24903,N_24734,N_24532);
xor U24904 (N_24904,N_24568,N_24580);
xor U24905 (N_24905,N_24666,N_24699);
nor U24906 (N_24906,N_24677,N_24574);
xor U24907 (N_24907,N_24682,N_24533);
nor U24908 (N_24908,N_24662,N_24714);
or U24909 (N_24909,N_24655,N_24647);
and U24910 (N_24910,N_24630,N_24532);
and U24911 (N_24911,N_24643,N_24581);
nand U24912 (N_24912,N_24690,N_24652);
xor U24913 (N_24913,N_24676,N_24527);
or U24914 (N_24914,N_24556,N_24585);
and U24915 (N_24915,N_24595,N_24729);
nor U24916 (N_24916,N_24633,N_24563);
nor U24917 (N_24917,N_24572,N_24744);
or U24918 (N_24918,N_24626,N_24729);
xor U24919 (N_24919,N_24641,N_24616);
nor U24920 (N_24920,N_24747,N_24589);
nor U24921 (N_24921,N_24655,N_24568);
or U24922 (N_24922,N_24662,N_24571);
xor U24923 (N_24923,N_24701,N_24600);
and U24924 (N_24924,N_24657,N_24509);
or U24925 (N_24925,N_24697,N_24614);
or U24926 (N_24926,N_24675,N_24627);
and U24927 (N_24927,N_24510,N_24614);
or U24928 (N_24928,N_24545,N_24526);
xor U24929 (N_24929,N_24713,N_24556);
xnor U24930 (N_24930,N_24629,N_24556);
nor U24931 (N_24931,N_24599,N_24587);
and U24932 (N_24932,N_24675,N_24552);
xnor U24933 (N_24933,N_24504,N_24715);
nor U24934 (N_24934,N_24599,N_24697);
and U24935 (N_24935,N_24672,N_24682);
xor U24936 (N_24936,N_24632,N_24638);
xnor U24937 (N_24937,N_24524,N_24608);
nand U24938 (N_24938,N_24658,N_24597);
xor U24939 (N_24939,N_24616,N_24503);
xnor U24940 (N_24940,N_24530,N_24576);
xnor U24941 (N_24941,N_24578,N_24621);
nand U24942 (N_24942,N_24737,N_24745);
or U24943 (N_24943,N_24619,N_24520);
nor U24944 (N_24944,N_24520,N_24585);
or U24945 (N_24945,N_24598,N_24696);
or U24946 (N_24946,N_24525,N_24747);
nor U24947 (N_24947,N_24580,N_24711);
xor U24948 (N_24948,N_24602,N_24592);
and U24949 (N_24949,N_24576,N_24661);
and U24950 (N_24950,N_24668,N_24517);
or U24951 (N_24951,N_24746,N_24641);
and U24952 (N_24952,N_24703,N_24584);
and U24953 (N_24953,N_24626,N_24501);
or U24954 (N_24954,N_24627,N_24677);
nand U24955 (N_24955,N_24644,N_24624);
nand U24956 (N_24956,N_24644,N_24549);
xor U24957 (N_24957,N_24712,N_24540);
or U24958 (N_24958,N_24554,N_24581);
or U24959 (N_24959,N_24567,N_24625);
or U24960 (N_24960,N_24630,N_24522);
nor U24961 (N_24961,N_24501,N_24520);
and U24962 (N_24962,N_24528,N_24676);
and U24963 (N_24963,N_24734,N_24666);
nor U24964 (N_24964,N_24618,N_24614);
nor U24965 (N_24965,N_24670,N_24721);
xnor U24966 (N_24966,N_24571,N_24736);
nor U24967 (N_24967,N_24626,N_24589);
xnor U24968 (N_24968,N_24573,N_24682);
xnor U24969 (N_24969,N_24586,N_24524);
nor U24970 (N_24970,N_24742,N_24638);
nand U24971 (N_24971,N_24528,N_24525);
nor U24972 (N_24972,N_24707,N_24647);
nor U24973 (N_24973,N_24575,N_24550);
or U24974 (N_24974,N_24669,N_24687);
nand U24975 (N_24975,N_24522,N_24579);
or U24976 (N_24976,N_24572,N_24605);
xnor U24977 (N_24977,N_24637,N_24563);
nor U24978 (N_24978,N_24513,N_24501);
nand U24979 (N_24979,N_24521,N_24578);
and U24980 (N_24980,N_24582,N_24652);
nor U24981 (N_24981,N_24682,N_24602);
or U24982 (N_24982,N_24664,N_24626);
xnor U24983 (N_24983,N_24556,N_24688);
and U24984 (N_24984,N_24722,N_24686);
and U24985 (N_24985,N_24701,N_24603);
nand U24986 (N_24986,N_24648,N_24512);
xnor U24987 (N_24987,N_24537,N_24742);
nor U24988 (N_24988,N_24711,N_24635);
xnor U24989 (N_24989,N_24529,N_24586);
nor U24990 (N_24990,N_24664,N_24604);
or U24991 (N_24991,N_24665,N_24707);
xor U24992 (N_24992,N_24584,N_24697);
nor U24993 (N_24993,N_24577,N_24563);
nand U24994 (N_24994,N_24564,N_24502);
xnor U24995 (N_24995,N_24581,N_24712);
and U24996 (N_24996,N_24643,N_24620);
nor U24997 (N_24997,N_24627,N_24639);
or U24998 (N_24998,N_24544,N_24532);
or U24999 (N_24999,N_24599,N_24549);
nor U25000 (N_25000,N_24947,N_24771);
xnor U25001 (N_25001,N_24755,N_24820);
and U25002 (N_25002,N_24775,N_24783);
or U25003 (N_25003,N_24959,N_24971);
nand U25004 (N_25004,N_24919,N_24931);
or U25005 (N_25005,N_24798,N_24878);
xnor U25006 (N_25006,N_24757,N_24942);
nor U25007 (N_25007,N_24821,N_24850);
and U25008 (N_25008,N_24901,N_24984);
nor U25009 (N_25009,N_24992,N_24786);
xor U25010 (N_25010,N_24832,N_24787);
nor U25011 (N_25011,N_24792,N_24868);
or U25012 (N_25012,N_24814,N_24808);
nor U25013 (N_25013,N_24767,N_24855);
nor U25014 (N_25014,N_24918,N_24951);
or U25015 (N_25015,N_24988,N_24807);
nor U25016 (N_25016,N_24994,N_24773);
xnor U25017 (N_25017,N_24998,N_24817);
nand U25018 (N_25018,N_24888,N_24957);
or U25019 (N_25019,N_24754,N_24961);
and U25020 (N_25020,N_24964,N_24825);
nand U25021 (N_25021,N_24781,N_24811);
and U25022 (N_25022,N_24837,N_24860);
or U25023 (N_25023,N_24995,N_24910);
nand U25024 (N_25024,N_24803,N_24823);
xnor U25025 (N_25025,N_24851,N_24900);
nor U25026 (N_25026,N_24946,N_24899);
nor U25027 (N_25027,N_24960,N_24885);
nand U25028 (N_25028,N_24954,N_24785);
nor U25029 (N_25029,N_24768,N_24978);
xnor U25030 (N_25030,N_24914,N_24936);
or U25031 (N_25031,N_24893,N_24997);
and U25032 (N_25032,N_24943,N_24835);
nand U25033 (N_25033,N_24962,N_24782);
or U25034 (N_25034,N_24916,N_24970);
nand U25035 (N_25035,N_24751,N_24950);
or U25036 (N_25036,N_24898,N_24805);
nand U25037 (N_25037,N_24973,N_24913);
xnor U25038 (N_25038,N_24977,N_24818);
xnor U25039 (N_25039,N_24883,N_24897);
xnor U25040 (N_25040,N_24958,N_24846);
and U25041 (N_25041,N_24813,N_24908);
nor U25042 (N_25042,N_24812,N_24842);
nor U25043 (N_25043,N_24830,N_24765);
nand U25044 (N_25044,N_24933,N_24928);
xnor U25045 (N_25045,N_24866,N_24758);
nor U25046 (N_25046,N_24800,N_24774);
xnor U25047 (N_25047,N_24953,N_24856);
and U25048 (N_25048,N_24996,N_24780);
nor U25049 (N_25049,N_24819,N_24909);
nor U25050 (N_25050,N_24759,N_24865);
nand U25051 (N_25051,N_24956,N_24930);
or U25052 (N_25052,N_24922,N_24777);
or U25053 (N_25053,N_24874,N_24816);
nand U25054 (N_25054,N_24838,N_24831);
nor U25055 (N_25055,N_24940,N_24863);
nand U25056 (N_25056,N_24857,N_24779);
xnor U25057 (N_25057,N_24892,N_24806);
xnor U25058 (N_25058,N_24882,N_24766);
nor U25059 (N_25059,N_24829,N_24834);
or U25060 (N_25060,N_24797,N_24993);
and U25061 (N_25061,N_24881,N_24890);
xnor U25062 (N_25062,N_24969,N_24952);
nand U25063 (N_25063,N_24845,N_24778);
nor U25064 (N_25064,N_24836,N_24987);
nand U25065 (N_25065,N_24809,N_24979);
or U25066 (N_25066,N_24944,N_24871);
xnor U25067 (N_25067,N_24965,N_24986);
xnor U25068 (N_25068,N_24924,N_24861);
xor U25069 (N_25069,N_24945,N_24873);
nand U25070 (N_25070,N_24802,N_24886);
nand U25071 (N_25071,N_24891,N_24772);
and U25072 (N_25072,N_24905,N_24903);
and U25073 (N_25073,N_24848,N_24750);
nor U25074 (N_25074,N_24932,N_24815);
xnor U25075 (N_25075,N_24763,N_24833);
or U25076 (N_25076,N_24799,N_24912);
and U25077 (N_25077,N_24824,N_24841);
nand U25078 (N_25078,N_24966,N_24938);
and U25079 (N_25079,N_24975,N_24801);
nand U25080 (N_25080,N_24794,N_24769);
xnor U25081 (N_25081,N_24963,N_24972);
or U25082 (N_25082,N_24991,N_24847);
or U25083 (N_25083,N_24753,N_24875);
and U25084 (N_25084,N_24864,N_24926);
nand U25085 (N_25085,N_24982,N_24762);
and U25086 (N_25086,N_24793,N_24983);
xor U25087 (N_25087,N_24858,N_24862);
and U25088 (N_25088,N_24925,N_24929);
or U25089 (N_25089,N_24752,N_24789);
or U25090 (N_25090,N_24844,N_24826);
xnor U25091 (N_25091,N_24990,N_24917);
xor U25092 (N_25092,N_24976,N_24985);
nand U25093 (N_25093,N_24876,N_24915);
nor U25094 (N_25094,N_24859,N_24887);
or U25095 (N_25095,N_24828,N_24770);
and U25096 (N_25096,N_24853,N_24894);
nand U25097 (N_25097,N_24796,N_24840);
xnor U25098 (N_25098,N_24896,N_24921);
and U25099 (N_25099,N_24949,N_24804);
xor U25100 (N_25100,N_24904,N_24941);
or U25101 (N_25101,N_24923,N_24902);
and U25102 (N_25102,N_24884,N_24791);
nand U25103 (N_25103,N_24839,N_24872);
xnor U25104 (N_25104,N_24968,N_24906);
nand U25105 (N_25105,N_24967,N_24756);
and U25106 (N_25106,N_24869,N_24920);
and U25107 (N_25107,N_24760,N_24870);
xor U25108 (N_25108,N_24822,N_24939);
nor U25109 (N_25109,N_24776,N_24788);
or U25110 (N_25110,N_24790,N_24999);
or U25111 (N_25111,N_24843,N_24827);
xor U25112 (N_25112,N_24907,N_24974);
nand U25113 (N_25113,N_24877,N_24895);
or U25114 (N_25114,N_24852,N_24911);
and U25115 (N_25115,N_24889,N_24795);
or U25116 (N_25116,N_24810,N_24989);
nor U25117 (N_25117,N_24879,N_24784);
nor U25118 (N_25118,N_24981,N_24849);
nand U25119 (N_25119,N_24854,N_24935);
xnor U25120 (N_25120,N_24761,N_24955);
nor U25121 (N_25121,N_24948,N_24927);
nor U25122 (N_25122,N_24980,N_24937);
xnor U25123 (N_25123,N_24867,N_24934);
nor U25124 (N_25124,N_24764,N_24880);
nor U25125 (N_25125,N_24753,N_24968);
nand U25126 (N_25126,N_24866,N_24813);
and U25127 (N_25127,N_24992,N_24966);
or U25128 (N_25128,N_24837,N_24893);
nor U25129 (N_25129,N_24866,N_24801);
xnor U25130 (N_25130,N_24951,N_24911);
nor U25131 (N_25131,N_24820,N_24782);
nor U25132 (N_25132,N_24750,N_24773);
and U25133 (N_25133,N_24776,N_24866);
nor U25134 (N_25134,N_24937,N_24844);
xor U25135 (N_25135,N_24857,N_24958);
nand U25136 (N_25136,N_24987,N_24879);
and U25137 (N_25137,N_24877,N_24903);
xor U25138 (N_25138,N_24904,N_24920);
nand U25139 (N_25139,N_24982,N_24880);
nor U25140 (N_25140,N_24958,N_24810);
nand U25141 (N_25141,N_24882,N_24750);
nand U25142 (N_25142,N_24850,N_24852);
nor U25143 (N_25143,N_24782,N_24850);
nor U25144 (N_25144,N_24894,N_24912);
nor U25145 (N_25145,N_24783,N_24985);
nand U25146 (N_25146,N_24869,N_24848);
xor U25147 (N_25147,N_24783,N_24769);
or U25148 (N_25148,N_24966,N_24948);
nor U25149 (N_25149,N_24953,N_24834);
or U25150 (N_25150,N_24760,N_24904);
nor U25151 (N_25151,N_24914,N_24799);
xor U25152 (N_25152,N_24771,N_24892);
or U25153 (N_25153,N_24966,N_24805);
or U25154 (N_25154,N_24926,N_24923);
and U25155 (N_25155,N_24898,N_24873);
xnor U25156 (N_25156,N_24830,N_24834);
or U25157 (N_25157,N_24872,N_24936);
nand U25158 (N_25158,N_24755,N_24758);
nand U25159 (N_25159,N_24848,N_24817);
or U25160 (N_25160,N_24907,N_24934);
nor U25161 (N_25161,N_24843,N_24850);
or U25162 (N_25162,N_24937,N_24880);
nand U25163 (N_25163,N_24900,N_24778);
nand U25164 (N_25164,N_24861,N_24886);
xnor U25165 (N_25165,N_24861,N_24815);
nand U25166 (N_25166,N_24973,N_24907);
or U25167 (N_25167,N_24785,N_24797);
nor U25168 (N_25168,N_24898,N_24880);
nor U25169 (N_25169,N_24753,N_24850);
nand U25170 (N_25170,N_24800,N_24859);
xor U25171 (N_25171,N_24789,N_24978);
or U25172 (N_25172,N_24991,N_24776);
nand U25173 (N_25173,N_24986,N_24945);
nand U25174 (N_25174,N_24833,N_24759);
xor U25175 (N_25175,N_24950,N_24886);
nor U25176 (N_25176,N_24763,N_24993);
nand U25177 (N_25177,N_24944,N_24764);
or U25178 (N_25178,N_24763,N_24983);
or U25179 (N_25179,N_24755,N_24866);
or U25180 (N_25180,N_24947,N_24895);
and U25181 (N_25181,N_24869,N_24856);
xor U25182 (N_25182,N_24790,N_24816);
nor U25183 (N_25183,N_24929,N_24915);
nor U25184 (N_25184,N_24871,N_24949);
and U25185 (N_25185,N_24960,N_24959);
or U25186 (N_25186,N_24914,N_24802);
nand U25187 (N_25187,N_24868,N_24797);
or U25188 (N_25188,N_24930,N_24792);
nand U25189 (N_25189,N_24930,N_24831);
or U25190 (N_25190,N_24892,N_24889);
and U25191 (N_25191,N_24902,N_24805);
or U25192 (N_25192,N_24803,N_24774);
nor U25193 (N_25193,N_24902,N_24751);
nor U25194 (N_25194,N_24771,N_24924);
and U25195 (N_25195,N_24794,N_24932);
or U25196 (N_25196,N_24963,N_24804);
and U25197 (N_25197,N_24932,N_24887);
xor U25198 (N_25198,N_24986,N_24826);
nor U25199 (N_25199,N_24848,N_24853);
and U25200 (N_25200,N_24764,N_24992);
xor U25201 (N_25201,N_24933,N_24847);
nand U25202 (N_25202,N_24921,N_24821);
or U25203 (N_25203,N_24950,N_24758);
xor U25204 (N_25204,N_24759,N_24976);
xor U25205 (N_25205,N_24923,N_24799);
nand U25206 (N_25206,N_24835,N_24977);
nand U25207 (N_25207,N_24952,N_24770);
xor U25208 (N_25208,N_24933,N_24915);
and U25209 (N_25209,N_24846,N_24907);
nor U25210 (N_25210,N_24970,N_24880);
nor U25211 (N_25211,N_24987,N_24898);
or U25212 (N_25212,N_24848,N_24841);
nand U25213 (N_25213,N_24882,N_24821);
xor U25214 (N_25214,N_24931,N_24779);
and U25215 (N_25215,N_24905,N_24805);
and U25216 (N_25216,N_24913,N_24892);
xor U25217 (N_25217,N_24759,N_24819);
and U25218 (N_25218,N_24855,N_24948);
nor U25219 (N_25219,N_24959,N_24913);
nand U25220 (N_25220,N_24863,N_24822);
and U25221 (N_25221,N_24825,N_24871);
or U25222 (N_25222,N_24817,N_24912);
nor U25223 (N_25223,N_24819,N_24895);
nand U25224 (N_25224,N_24819,N_24893);
xor U25225 (N_25225,N_24784,N_24993);
nand U25226 (N_25226,N_24784,N_24826);
nand U25227 (N_25227,N_24783,N_24861);
or U25228 (N_25228,N_24772,N_24978);
xnor U25229 (N_25229,N_24944,N_24994);
nor U25230 (N_25230,N_24928,N_24782);
nand U25231 (N_25231,N_24890,N_24837);
and U25232 (N_25232,N_24784,N_24925);
xor U25233 (N_25233,N_24972,N_24772);
nand U25234 (N_25234,N_24926,N_24878);
or U25235 (N_25235,N_24976,N_24854);
and U25236 (N_25236,N_24851,N_24839);
or U25237 (N_25237,N_24906,N_24965);
and U25238 (N_25238,N_24960,N_24924);
and U25239 (N_25239,N_24798,N_24814);
xnor U25240 (N_25240,N_24798,N_24776);
nand U25241 (N_25241,N_24985,N_24997);
and U25242 (N_25242,N_24765,N_24853);
or U25243 (N_25243,N_24758,N_24912);
nand U25244 (N_25244,N_24942,N_24815);
xnor U25245 (N_25245,N_24846,N_24802);
or U25246 (N_25246,N_24944,N_24906);
nor U25247 (N_25247,N_24950,N_24966);
and U25248 (N_25248,N_24983,N_24972);
and U25249 (N_25249,N_24893,N_24758);
and U25250 (N_25250,N_25075,N_25083);
and U25251 (N_25251,N_25097,N_25094);
xnor U25252 (N_25252,N_25031,N_25203);
or U25253 (N_25253,N_25242,N_25139);
nand U25254 (N_25254,N_25046,N_25175);
nand U25255 (N_25255,N_25214,N_25130);
nand U25256 (N_25256,N_25199,N_25172);
and U25257 (N_25257,N_25190,N_25155);
nor U25258 (N_25258,N_25124,N_25115);
nor U25259 (N_25259,N_25174,N_25128);
or U25260 (N_25260,N_25148,N_25100);
and U25261 (N_25261,N_25068,N_25184);
nor U25262 (N_25262,N_25185,N_25222);
nor U25263 (N_25263,N_25099,N_25073);
nand U25264 (N_25264,N_25112,N_25229);
nor U25265 (N_25265,N_25240,N_25078);
xnor U25266 (N_25266,N_25061,N_25017);
and U25267 (N_25267,N_25035,N_25171);
nor U25268 (N_25268,N_25003,N_25197);
xnor U25269 (N_25269,N_25206,N_25062);
nor U25270 (N_25270,N_25117,N_25104);
or U25271 (N_25271,N_25110,N_25230);
and U25272 (N_25272,N_25109,N_25238);
nand U25273 (N_25273,N_25091,N_25137);
xor U25274 (N_25274,N_25015,N_25173);
and U25275 (N_25275,N_25058,N_25113);
nand U25276 (N_25276,N_25147,N_25038);
xor U25277 (N_25277,N_25131,N_25201);
nor U25278 (N_25278,N_25030,N_25223);
nand U25279 (N_25279,N_25055,N_25087);
nor U25280 (N_25280,N_25085,N_25237);
or U25281 (N_25281,N_25029,N_25162);
xnor U25282 (N_25282,N_25025,N_25165);
nor U25283 (N_25283,N_25052,N_25133);
and U25284 (N_25284,N_25111,N_25011);
xor U25285 (N_25285,N_25244,N_25006);
nand U25286 (N_25286,N_25157,N_25014);
nor U25287 (N_25287,N_25026,N_25040);
nand U25288 (N_25288,N_25243,N_25096);
nand U25289 (N_25289,N_25067,N_25121);
or U25290 (N_25290,N_25108,N_25146);
nand U25291 (N_25291,N_25063,N_25160);
or U25292 (N_25292,N_25123,N_25010);
or U25293 (N_25293,N_25178,N_25071);
xnor U25294 (N_25294,N_25141,N_25159);
xnor U25295 (N_25295,N_25004,N_25152);
or U25296 (N_25296,N_25008,N_25107);
and U25297 (N_25297,N_25034,N_25024);
nand U25298 (N_25298,N_25126,N_25013);
xnor U25299 (N_25299,N_25217,N_25050);
and U25300 (N_25300,N_25207,N_25216);
and U25301 (N_25301,N_25239,N_25150);
or U25302 (N_25302,N_25022,N_25151);
and U25303 (N_25303,N_25023,N_25249);
nand U25304 (N_25304,N_25009,N_25028);
and U25305 (N_25305,N_25154,N_25118);
and U25306 (N_25306,N_25079,N_25106);
xor U25307 (N_25307,N_25205,N_25166);
or U25308 (N_25308,N_25202,N_25248);
nand U25309 (N_25309,N_25226,N_25168);
or U25310 (N_25310,N_25236,N_25016);
xnor U25311 (N_25311,N_25192,N_25169);
nand U25312 (N_25312,N_25210,N_25057);
or U25313 (N_25313,N_25101,N_25233);
or U25314 (N_25314,N_25221,N_25156);
nand U25315 (N_25315,N_25225,N_25195);
nor U25316 (N_25316,N_25153,N_25065);
xor U25317 (N_25317,N_25129,N_25127);
or U25318 (N_25318,N_25098,N_25125);
nor U25319 (N_25319,N_25086,N_25018);
and U25320 (N_25320,N_25188,N_25218);
and U25321 (N_25321,N_25177,N_25180);
xnor U25322 (N_25322,N_25076,N_25183);
or U25323 (N_25323,N_25093,N_25163);
xnor U25324 (N_25324,N_25193,N_25000);
or U25325 (N_25325,N_25196,N_25039);
and U25326 (N_25326,N_25186,N_25005);
nor U25327 (N_25327,N_25212,N_25200);
or U25328 (N_25328,N_25103,N_25181);
and U25329 (N_25329,N_25092,N_25144);
or U25330 (N_25330,N_25102,N_25048);
or U25331 (N_25331,N_25082,N_25220);
nor U25332 (N_25332,N_25072,N_25161);
nor U25333 (N_25333,N_25081,N_25049);
and U25334 (N_25334,N_25158,N_25119);
and U25335 (N_25335,N_25051,N_25247);
xnor U25336 (N_25336,N_25043,N_25020);
and U25337 (N_25337,N_25135,N_25069);
and U25338 (N_25338,N_25044,N_25227);
or U25339 (N_25339,N_25234,N_25164);
xor U25340 (N_25340,N_25246,N_25047);
xor U25341 (N_25341,N_25027,N_25167);
and U25342 (N_25342,N_25002,N_25056);
nand U25343 (N_25343,N_25032,N_25036);
or U25344 (N_25344,N_25176,N_25089);
nor U25345 (N_25345,N_25149,N_25077);
or U25346 (N_25346,N_25066,N_25194);
nand U25347 (N_25347,N_25208,N_25136);
nor U25348 (N_25348,N_25215,N_25170);
or U25349 (N_25349,N_25187,N_25090);
xnor U25350 (N_25350,N_25142,N_25231);
nand U25351 (N_25351,N_25245,N_25224);
nand U25352 (N_25352,N_25211,N_25088);
and U25353 (N_25353,N_25198,N_25037);
nor U25354 (N_25354,N_25138,N_25191);
nor U25355 (N_25355,N_25122,N_25209);
and U25356 (N_25356,N_25189,N_25033);
and U25357 (N_25357,N_25095,N_25232);
xnor U25358 (N_25358,N_25143,N_25241);
nor U25359 (N_25359,N_25070,N_25213);
xnor U25360 (N_25360,N_25021,N_25105);
nor U25361 (N_25361,N_25064,N_25007);
and U25362 (N_25362,N_25001,N_25045);
xnor U25363 (N_25363,N_25219,N_25114);
or U25364 (N_25364,N_25074,N_25179);
and U25365 (N_25365,N_25060,N_25054);
xnor U25366 (N_25366,N_25053,N_25134);
and U25367 (N_25367,N_25084,N_25140);
and U25368 (N_25368,N_25204,N_25080);
nor U25369 (N_25369,N_25116,N_25182);
nor U25370 (N_25370,N_25120,N_25235);
nor U25371 (N_25371,N_25228,N_25012);
xnor U25372 (N_25372,N_25132,N_25041);
nor U25373 (N_25373,N_25059,N_25019);
and U25374 (N_25374,N_25145,N_25042);
xnor U25375 (N_25375,N_25130,N_25021);
nand U25376 (N_25376,N_25125,N_25119);
nor U25377 (N_25377,N_25025,N_25120);
nor U25378 (N_25378,N_25172,N_25205);
xor U25379 (N_25379,N_25063,N_25222);
xnor U25380 (N_25380,N_25108,N_25070);
or U25381 (N_25381,N_25178,N_25089);
nor U25382 (N_25382,N_25157,N_25171);
xor U25383 (N_25383,N_25175,N_25243);
or U25384 (N_25384,N_25244,N_25010);
or U25385 (N_25385,N_25221,N_25142);
nor U25386 (N_25386,N_25074,N_25137);
or U25387 (N_25387,N_25166,N_25121);
nand U25388 (N_25388,N_25106,N_25212);
or U25389 (N_25389,N_25049,N_25170);
or U25390 (N_25390,N_25228,N_25241);
nor U25391 (N_25391,N_25010,N_25183);
xnor U25392 (N_25392,N_25120,N_25115);
and U25393 (N_25393,N_25245,N_25227);
nor U25394 (N_25394,N_25198,N_25098);
xor U25395 (N_25395,N_25223,N_25003);
nor U25396 (N_25396,N_25125,N_25189);
xnor U25397 (N_25397,N_25245,N_25005);
or U25398 (N_25398,N_25222,N_25056);
or U25399 (N_25399,N_25147,N_25213);
nand U25400 (N_25400,N_25231,N_25075);
nor U25401 (N_25401,N_25022,N_25218);
and U25402 (N_25402,N_25072,N_25165);
and U25403 (N_25403,N_25023,N_25063);
xor U25404 (N_25404,N_25126,N_25237);
and U25405 (N_25405,N_25071,N_25161);
xor U25406 (N_25406,N_25158,N_25031);
and U25407 (N_25407,N_25180,N_25206);
nand U25408 (N_25408,N_25201,N_25024);
nand U25409 (N_25409,N_25234,N_25063);
nor U25410 (N_25410,N_25161,N_25100);
nor U25411 (N_25411,N_25179,N_25050);
and U25412 (N_25412,N_25097,N_25035);
nand U25413 (N_25413,N_25165,N_25202);
xnor U25414 (N_25414,N_25129,N_25235);
xnor U25415 (N_25415,N_25166,N_25206);
xnor U25416 (N_25416,N_25245,N_25203);
nor U25417 (N_25417,N_25151,N_25230);
and U25418 (N_25418,N_25079,N_25061);
and U25419 (N_25419,N_25187,N_25109);
xnor U25420 (N_25420,N_25123,N_25046);
xnor U25421 (N_25421,N_25164,N_25136);
nor U25422 (N_25422,N_25202,N_25221);
xor U25423 (N_25423,N_25151,N_25052);
and U25424 (N_25424,N_25153,N_25175);
nand U25425 (N_25425,N_25005,N_25223);
nor U25426 (N_25426,N_25180,N_25194);
nand U25427 (N_25427,N_25185,N_25113);
or U25428 (N_25428,N_25199,N_25069);
xor U25429 (N_25429,N_25228,N_25132);
and U25430 (N_25430,N_25185,N_25145);
and U25431 (N_25431,N_25205,N_25074);
nand U25432 (N_25432,N_25201,N_25186);
xor U25433 (N_25433,N_25082,N_25191);
or U25434 (N_25434,N_25031,N_25173);
nand U25435 (N_25435,N_25015,N_25231);
nor U25436 (N_25436,N_25017,N_25001);
xor U25437 (N_25437,N_25190,N_25023);
nor U25438 (N_25438,N_25174,N_25212);
xnor U25439 (N_25439,N_25209,N_25192);
nand U25440 (N_25440,N_25117,N_25076);
xnor U25441 (N_25441,N_25100,N_25233);
nand U25442 (N_25442,N_25143,N_25026);
or U25443 (N_25443,N_25158,N_25097);
nand U25444 (N_25444,N_25100,N_25137);
xnor U25445 (N_25445,N_25243,N_25074);
nand U25446 (N_25446,N_25243,N_25185);
nand U25447 (N_25447,N_25212,N_25157);
or U25448 (N_25448,N_25039,N_25031);
nand U25449 (N_25449,N_25220,N_25212);
nand U25450 (N_25450,N_25045,N_25154);
or U25451 (N_25451,N_25197,N_25247);
and U25452 (N_25452,N_25004,N_25094);
xnor U25453 (N_25453,N_25042,N_25062);
and U25454 (N_25454,N_25216,N_25228);
nand U25455 (N_25455,N_25239,N_25109);
nor U25456 (N_25456,N_25019,N_25148);
nor U25457 (N_25457,N_25060,N_25219);
or U25458 (N_25458,N_25003,N_25162);
or U25459 (N_25459,N_25103,N_25148);
or U25460 (N_25460,N_25133,N_25103);
xor U25461 (N_25461,N_25079,N_25111);
nand U25462 (N_25462,N_25209,N_25228);
nor U25463 (N_25463,N_25239,N_25211);
or U25464 (N_25464,N_25043,N_25045);
nand U25465 (N_25465,N_25232,N_25237);
and U25466 (N_25466,N_25031,N_25195);
nor U25467 (N_25467,N_25157,N_25085);
xnor U25468 (N_25468,N_25174,N_25224);
xor U25469 (N_25469,N_25037,N_25121);
and U25470 (N_25470,N_25161,N_25222);
nor U25471 (N_25471,N_25185,N_25072);
nor U25472 (N_25472,N_25018,N_25155);
or U25473 (N_25473,N_25017,N_25068);
or U25474 (N_25474,N_25068,N_25025);
and U25475 (N_25475,N_25033,N_25082);
and U25476 (N_25476,N_25020,N_25065);
or U25477 (N_25477,N_25249,N_25140);
or U25478 (N_25478,N_25225,N_25013);
nand U25479 (N_25479,N_25187,N_25020);
or U25480 (N_25480,N_25035,N_25220);
xor U25481 (N_25481,N_25055,N_25196);
nand U25482 (N_25482,N_25228,N_25182);
and U25483 (N_25483,N_25201,N_25046);
xnor U25484 (N_25484,N_25102,N_25154);
and U25485 (N_25485,N_25052,N_25041);
xor U25486 (N_25486,N_25104,N_25180);
nor U25487 (N_25487,N_25224,N_25118);
nand U25488 (N_25488,N_25224,N_25060);
nand U25489 (N_25489,N_25184,N_25244);
or U25490 (N_25490,N_25213,N_25172);
nor U25491 (N_25491,N_25209,N_25201);
or U25492 (N_25492,N_25028,N_25134);
or U25493 (N_25493,N_25219,N_25187);
xnor U25494 (N_25494,N_25105,N_25201);
nor U25495 (N_25495,N_25115,N_25188);
xnor U25496 (N_25496,N_25019,N_25130);
nand U25497 (N_25497,N_25196,N_25056);
or U25498 (N_25498,N_25159,N_25110);
xor U25499 (N_25499,N_25196,N_25159);
nand U25500 (N_25500,N_25488,N_25294);
xor U25501 (N_25501,N_25285,N_25478);
nand U25502 (N_25502,N_25305,N_25486);
nand U25503 (N_25503,N_25382,N_25466);
or U25504 (N_25504,N_25267,N_25359);
xor U25505 (N_25505,N_25341,N_25283);
and U25506 (N_25506,N_25268,N_25428);
nor U25507 (N_25507,N_25456,N_25462);
or U25508 (N_25508,N_25273,N_25314);
nand U25509 (N_25509,N_25331,N_25470);
or U25510 (N_25510,N_25260,N_25410);
nand U25511 (N_25511,N_25380,N_25265);
and U25512 (N_25512,N_25290,N_25460);
or U25513 (N_25513,N_25367,N_25439);
xnor U25514 (N_25514,N_25277,N_25477);
and U25515 (N_25515,N_25403,N_25333);
or U25516 (N_25516,N_25386,N_25459);
nand U25517 (N_25517,N_25446,N_25253);
xor U25518 (N_25518,N_25396,N_25490);
xor U25519 (N_25519,N_25276,N_25298);
xor U25520 (N_25520,N_25472,N_25362);
xor U25521 (N_25521,N_25479,N_25413);
and U25522 (N_25522,N_25339,N_25302);
nand U25523 (N_25523,N_25350,N_25385);
or U25524 (N_25524,N_25445,N_25296);
or U25525 (N_25525,N_25442,N_25360);
nand U25526 (N_25526,N_25322,N_25365);
or U25527 (N_25527,N_25419,N_25496);
and U25528 (N_25528,N_25356,N_25404);
or U25529 (N_25529,N_25480,N_25448);
or U25530 (N_25530,N_25420,N_25287);
or U25531 (N_25531,N_25414,N_25491);
or U25532 (N_25532,N_25266,N_25434);
xnor U25533 (N_25533,N_25402,N_25324);
or U25534 (N_25534,N_25361,N_25497);
nand U25535 (N_25535,N_25441,N_25326);
nand U25536 (N_25536,N_25433,N_25307);
nand U25537 (N_25537,N_25475,N_25429);
and U25538 (N_25538,N_25467,N_25259);
nor U25539 (N_25539,N_25288,N_25327);
or U25540 (N_25540,N_25257,N_25383);
nor U25541 (N_25541,N_25375,N_25281);
and U25542 (N_25542,N_25393,N_25256);
nor U25543 (N_25543,N_25476,N_25399);
nor U25544 (N_25544,N_25338,N_25292);
nor U25545 (N_25545,N_25318,N_25493);
nand U25546 (N_25546,N_25328,N_25309);
nand U25547 (N_25547,N_25251,N_25374);
nor U25548 (N_25548,N_25464,N_25443);
and U25549 (N_25549,N_25320,N_25368);
nand U25550 (N_25550,N_25263,N_25351);
xnor U25551 (N_25551,N_25310,N_25355);
and U25552 (N_25552,N_25492,N_25264);
xnor U25553 (N_25553,N_25358,N_25482);
or U25554 (N_25554,N_25494,N_25284);
and U25555 (N_25555,N_25395,N_25461);
xor U25556 (N_25556,N_25303,N_25406);
and U25557 (N_25557,N_25471,N_25408);
and U25558 (N_25558,N_25417,N_25463);
nor U25559 (N_25559,N_25437,N_25390);
or U25560 (N_25560,N_25407,N_25297);
nor U25561 (N_25561,N_25357,N_25495);
and U25562 (N_25562,N_25364,N_25376);
nor U25563 (N_25563,N_25308,N_25258);
nand U25564 (N_25564,N_25301,N_25340);
and U25565 (N_25565,N_25481,N_25261);
and U25566 (N_25566,N_25274,N_25421);
xnor U25567 (N_25567,N_25370,N_25325);
nand U25568 (N_25568,N_25312,N_25289);
nor U25569 (N_25569,N_25450,N_25432);
and U25570 (N_25570,N_25348,N_25352);
and U25571 (N_25571,N_25279,N_25425);
or U25572 (N_25572,N_25354,N_25498);
and U25573 (N_25573,N_25252,N_25342);
nand U25574 (N_25574,N_25405,N_25484);
and U25575 (N_25575,N_25457,N_25392);
nand U25576 (N_25576,N_25426,N_25270);
nor U25577 (N_25577,N_25334,N_25250);
nand U25578 (N_25578,N_25483,N_25391);
xor U25579 (N_25579,N_25424,N_25387);
and U25580 (N_25580,N_25254,N_25379);
nand U25581 (N_25581,N_25452,N_25317);
nand U25582 (N_25582,N_25313,N_25347);
nand U25583 (N_25583,N_25306,N_25409);
nor U25584 (N_25584,N_25344,N_25291);
or U25585 (N_25585,N_25278,N_25316);
nor U25586 (N_25586,N_25415,N_25400);
or U25587 (N_25587,N_25423,N_25311);
nor U25588 (N_25588,N_25373,N_25343);
xor U25589 (N_25589,N_25304,N_25451);
xor U25590 (N_25590,N_25458,N_25468);
nor U25591 (N_25591,N_25388,N_25293);
and U25592 (N_25592,N_25469,N_25438);
nand U25593 (N_25593,N_25431,N_25371);
xnor U25594 (N_25594,N_25394,N_25453);
or U25595 (N_25595,N_25384,N_25262);
nand U25596 (N_25596,N_25440,N_25353);
and U25597 (N_25597,N_25275,N_25455);
xor U25598 (N_25598,N_25282,N_25321);
and U25599 (N_25599,N_25255,N_25485);
nor U25600 (N_25600,N_25465,N_25319);
xnor U25601 (N_25601,N_25335,N_25487);
nor U25602 (N_25602,N_25332,N_25389);
or U25603 (N_25603,N_25418,N_25300);
and U25604 (N_25604,N_25280,N_25427);
nor U25605 (N_25605,N_25474,N_25447);
nor U25606 (N_25606,N_25422,N_25436);
or U25607 (N_25607,N_25416,N_25299);
nand U25608 (N_25608,N_25345,N_25411);
xnor U25609 (N_25609,N_25315,N_25369);
or U25610 (N_25610,N_25330,N_25329);
xor U25611 (N_25611,N_25272,N_25271);
or U25612 (N_25612,N_25366,N_25412);
nor U25613 (N_25613,N_25444,N_25295);
nor U25614 (N_25614,N_25449,N_25435);
or U25615 (N_25615,N_25372,N_25454);
nand U25616 (N_25616,N_25430,N_25397);
xor U25617 (N_25617,N_25378,N_25499);
nand U25618 (N_25618,N_25349,N_25286);
nand U25619 (N_25619,N_25363,N_25489);
xor U25620 (N_25620,N_25336,N_25323);
and U25621 (N_25621,N_25401,N_25473);
xnor U25622 (N_25622,N_25346,N_25398);
and U25623 (N_25623,N_25337,N_25269);
and U25624 (N_25624,N_25377,N_25381);
or U25625 (N_25625,N_25306,N_25312);
nand U25626 (N_25626,N_25466,N_25341);
nor U25627 (N_25627,N_25306,N_25429);
and U25628 (N_25628,N_25496,N_25420);
nand U25629 (N_25629,N_25352,N_25361);
nand U25630 (N_25630,N_25322,N_25484);
and U25631 (N_25631,N_25271,N_25464);
nor U25632 (N_25632,N_25274,N_25499);
or U25633 (N_25633,N_25395,N_25330);
nor U25634 (N_25634,N_25372,N_25417);
nand U25635 (N_25635,N_25306,N_25259);
nor U25636 (N_25636,N_25436,N_25377);
or U25637 (N_25637,N_25393,N_25439);
or U25638 (N_25638,N_25438,N_25387);
xnor U25639 (N_25639,N_25451,N_25375);
or U25640 (N_25640,N_25274,N_25324);
xor U25641 (N_25641,N_25286,N_25268);
and U25642 (N_25642,N_25409,N_25384);
nand U25643 (N_25643,N_25310,N_25309);
nand U25644 (N_25644,N_25356,N_25452);
or U25645 (N_25645,N_25315,N_25460);
nor U25646 (N_25646,N_25351,N_25404);
or U25647 (N_25647,N_25299,N_25435);
and U25648 (N_25648,N_25313,N_25474);
and U25649 (N_25649,N_25499,N_25496);
xnor U25650 (N_25650,N_25388,N_25338);
or U25651 (N_25651,N_25447,N_25286);
and U25652 (N_25652,N_25326,N_25386);
or U25653 (N_25653,N_25400,N_25302);
and U25654 (N_25654,N_25312,N_25277);
xnor U25655 (N_25655,N_25384,N_25414);
or U25656 (N_25656,N_25460,N_25285);
nor U25657 (N_25657,N_25353,N_25272);
nor U25658 (N_25658,N_25426,N_25482);
nand U25659 (N_25659,N_25385,N_25431);
or U25660 (N_25660,N_25435,N_25369);
nand U25661 (N_25661,N_25330,N_25483);
nand U25662 (N_25662,N_25252,N_25283);
nor U25663 (N_25663,N_25275,N_25427);
nand U25664 (N_25664,N_25282,N_25335);
nor U25665 (N_25665,N_25397,N_25440);
nand U25666 (N_25666,N_25370,N_25332);
xor U25667 (N_25667,N_25267,N_25266);
nor U25668 (N_25668,N_25394,N_25405);
nor U25669 (N_25669,N_25482,N_25254);
or U25670 (N_25670,N_25294,N_25296);
nor U25671 (N_25671,N_25362,N_25496);
xor U25672 (N_25672,N_25390,N_25343);
nor U25673 (N_25673,N_25344,N_25436);
and U25674 (N_25674,N_25322,N_25457);
nor U25675 (N_25675,N_25473,N_25317);
and U25676 (N_25676,N_25317,N_25422);
xor U25677 (N_25677,N_25351,N_25325);
xnor U25678 (N_25678,N_25349,N_25431);
and U25679 (N_25679,N_25421,N_25466);
nor U25680 (N_25680,N_25330,N_25301);
xnor U25681 (N_25681,N_25453,N_25498);
and U25682 (N_25682,N_25288,N_25362);
or U25683 (N_25683,N_25473,N_25445);
and U25684 (N_25684,N_25367,N_25349);
and U25685 (N_25685,N_25274,N_25341);
or U25686 (N_25686,N_25298,N_25370);
and U25687 (N_25687,N_25261,N_25404);
and U25688 (N_25688,N_25278,N_25265);
and U25689 (N_25689,N_25451,N_25464);
and U25690 (N_25690,N_25361,N_25473);
nand U25691 (N_25691,N_25458,N_25427);
xor U25692 (N_25692,N_25296,N_25348);
nand U25693 (N_25693,N_25386,N_25426);
nor U25694 (N_25694,N_25354,N_25342);
nor U25695 (N_25695,N_25419,N_25408);
xnor U25696 (N_25696,N_25276,N_25369);
or U25697 (N_25697,N_25311,N_25333);
xor U25698 (N_25698,N_25479,N_25293);
or U25699 (N_25699,N_25296,N_25494);
and U25700 (N_25700,N_25486,N_25378);
nor U25701 (N_25701,N_25443,N_25394);
xnor U25702 (N_25702,N_25453,N_25447);
nand U25703 (N_25703,N_25381,N_25364);
and U25704 (N_25704,N_25408,N_25266);
or U25705 (N_25705,N_25298,N_25300);
and U25706 (N_25706,N_25282,N_25271);
and U25707 (N_25707,N_25380,N_25363);
and U25708 (N_25708,N_25411,N_25420);
nand U25709 (N_25709,N_25398,N_25428);
nand U25710 (N_25710,N_25406,N_25379);
or U25711 (N_25711,N_25262,N_25305);
xor U25712 (N_25712,N_25335,N_25322);
or U25713 (N_25713,N_25373,N_25461);
nand U25714 (N_25714,N_25330,N_25384);
xnor U25715 (N_25715,N_25252,N_25425);
and U25716 (N_25716,N_25355,N_25266);
or U25717 (N_25717,N_25403,N_25269);
xor U25718 (N_25718,N_25488,N_25358);
nor U25719 (N_25719,N_25304,N_25373);
or U25720 (N_25720,N_25355,N_25255);
xor U25721 (N_25721,N_25403,N_25263);
or U25722 (N_25722,N_25265,N_25450);
nand U25723 (N_25723,N_25367,N_25250);
nand U25724 (N_25724,N_25488,N_25314);
and U25725 (N_25725,N_25376,N_25313);
or U25726 (N_25726,N_25394,N_25329);
nor U25727 (N_25727,N_25321,N_25495);
or U25728 (N_25728,N_25354,N_25297);
xor U25729 (N_25729,N_25385,N_25352);
or U25730 (N_25730,N_25268,N_25284);
or U25731 (N_25731,N_25353,N_25370);
nand U25732 (N_25732,N_25295,N_25346);
xnor U25733 (N_25733,N_25252,N_25419);
and U25734 (N_25734,N_25435,N_25474);
xor U25735 (N_25735,N_25300,N_25424);
xor U25736 (N_25736,N_25304,N_25372);
nor U25737 (N_25737,N_25312,N_25444);
xor U25738 (N_25738,N_25386,N_25353);
and U25739 (N_25739,N_25275,N_25443);
or U25740 (N_25740,N_25290,N_25320);
nand U25741 (N_25741,N_25469,N_25294);
nand U25742 (N_25742,N_25310,N_25302);
xor U25743 (N_25743,N_25440,N_25282);
nor U25744 (N_25744,N_25440,N_25403);
xnor U25745 (N_25745,N_25375,N_25363);
or U25746 (N_25746,N_25472,N_25486);
nor U25747 (N_25747,N_25304,N_25260);
nor U25748 (N_25748,N_25317,N_25290);
and U25749 (N_25749,N_25324,N_25252);
nand U25750 (N_25750,N_25693,N_25740);
nand U25751 (N_25751,N_25610,N_25551);
nand U25752 (N_25752,N_25627,N_25507);
and U25753 (N_25753,N_25748,N_25653);
and U25754 (N_25754,N_25588,N_25631);
nor U25755 (N_25755,N_25545,N_25594);
nor U25756 (N_25756,N_25669,N_25613);
or U25757 (N_25757,N_25719,N_25739);
nand U25758 (N_25758,N_25737,N_25646);
xor U25759 (N_25759,N_25640,N_25686);
and U25760 (N_25760,N_25515,N_25528);
nor U25761 (N_25761,N_25526,N_25622);
nor U25762 (N_25762,N_25616,N_25603);
and U25763 (N_25763,N_25662,N_25657);
nor U25764 (N_25764,N_25576,N_25654);
or U25765 (N_25765,N_25523,N_25505);
nand U25766 (N_25766,N_25604,N_25635);
and U25767 (N_25767,N_25517,N_25566);
and U25768 (N_25768,N_25597,N_25525);
nor U25769 (N_25769,N_25733,N_25655);
nor U25770 (N_25770,N_25673,N_25695);
nor U25771 (N_25771,N_25677,N_25735);
nor U25772 (N_25772,N_25641,N_25687);
nor U25773 (N_25773,N_25738,N_25659);
nor U25774 (N_25774,N_25547,N_25625);
and U25775 (N_25775,N_25674,N_25558);
xnor U25776 (N_25776,N_25514,N_25624);
nor U25777 (N_25777,N_25734,N_25516);
xor U25778 (N_25778,N_25581,N_25726);
or U25779 (N_25779,N_25632,N_25650);
and U25780 (N_25780,N_25549,N_25562);
or U25781 (N_25781,N_25591,N_25548);
nor U25782 (N_25782,N_25729,N_25745);
or U25783 (N_25783,N_25555,N_25690);
xor U25784 (N_25784,N_25592,N_25701);
xnor U25785 (N_25785,N_25556,N_25712);
nor U25786 (N_25786,N_25663,N_25533);
nor U25787 (N_25787,N_25511,N_25527);
nor U25788 (N_25788,N_25519,N_25544);
and U25789 (N_25789,N_25518,N_25723);
nor U25790 (N_25790,N_25658,N_25731);
nor U25791 (N_25791,N_25720,N_25552);
nor U25792 (N_25792,N_25721,N_25716);
nand U25793 (N_25793,N_25718,N_25570);
and U25794 (N_25794,N_25697,N_25599);
xor U25795 (N_25795,N_25500,N_25649);
nand U25796 (N_25796,N_25609,N_25602);
and U25797 (N_25797,N_25671,N_25578);
xor U25798 (N_25798,N_25684,N_25656);
nand U25799 (N_25799,N_25704,N_25676);
or U25800 (N_25800,N_25506,N_25584);
nand U25801 (N_25801,N_25681,N_25691);
xor U25802 (N_25802,N_25713,N_25502);
or U25803 (N_25803,N_25615,N_25727);
nand U25804 (N_25804,N_25696,N_25575);
or U25805 (N_25805,N_25543,N_25564);
nand U25806 (N_25806,N_25728,N_25619);
nand U25807 (N_25807,N_25736,N_25582);
nand U25808 (N_25808,N_25621,N_25563);
nor U25809 (N_25809,N_25577,N_25706);
nand U25810 (N_25810,N_25583,N_25538);
nand U25811 (N_25811,N_25705,N_25560);
xnor U25812 (N_25812,N_25611,N_25585);
or U25813 (N_25813,N_25537,N_25586);
xnor U25814 (N_25814,N_25553,N_25698);
xor U25815 (N_25815,N_25579,N_25699);
and U25816 (N_25816,N_25708,N_25521);
nand U25817 (N_25817,N_25541,N_25668);
or U25818 (N_25818,N_25666,N_25565);
and U25819 (N_25819,N_25652,N_25642);
and U25820 (N_25820,N_25638,N_25675);
and U25821 (N_25821,N_25568,N_25682);
xnor U25822 (N_25822,N_25651,N_25512);
nor U25823 (N_25823,N_25510,N_25747);
and U25824 (N_25824,N_25606,N_25680);
xor U25825 (N_25825,N_25571,N_25542);
and U25826 (N_25826,N_25741,N_25730);
or U25827 (N_25827,N_25629,N_25605);
xor U25828 (N_25828,N_25633,N_25614);
and U25829 (N_25829,N_25530,N_25679);
nor U25830 (N_25830,N_25744,N_25561);
or U25831 (N_25831,N_25643,N_25743);
or U25832 (N_25832,N_25531,N_25630);
nand U25833 (N_25833,N_25550,N_25574);
or U25834 (N_25834,N_25637,N_25535);
xor U25835 (N_25835,N_25540,N_25513);
or U25836 (N_25836,N_25539,N_25601);
nand U25837 (N_25837,N_25692,N_25580);
nand U25838 (N_25838,N_25694,N_25715);
and U25839 (N_25839,N_25636,N_25569);
nand U25840 (N_25840,N_25534,N_25532);
nand U25841 (N_25841,N_25714,N_25689);
xnor U25842 (N_25842,N_25522,N_25626);
nor U25843 (N_25843,N_25501,N_25702);
and U25844 (N_25844,N_25722,N_25725);
or U25845 (N_25845,N_25634,N_25648);
xnor U25846 (N_25846,N_25709,N_25710);
nand U25847 (N_25847,N_25700,N_25572);
nand U25848 (N_25848,N_25711,N_25639);
nor U25849 (N_25849,N_25593,N_25524);
or U25850 (N_25850,N_25667,N_25647);
xnor U25851 (N_25851,N_25504,N_25623);
xor U25852 (N_25852,N_25612,N_25595);
nor U25853 (N_25853,N_25587,N_25590);
nor U25854 (N_25854,N_25617,N_25685);
nor U25855 (N_25855,N_25546,N_25598);
and U25856 (N_25856,N_25664,N_25536);
xnor U25857 (N_25857,N_25670,N_25707);
nor U25858 (N_25858,N_25620,N_25559);
nor U25859 (N_25859,N_25672,N_25703);
and U25860 (N_25860,N_25520,N_25683);
nand U25861 (N_25861,N_25644,N_25554);
xnor U25862 (N_25862,N_25557,N_25618);
xor U25863 (N_25863,N_25607,N_25746);
xnor U25864 (N_25864,N_25503,N_25628);
and U25865 (N_25865,N_25742,N_25732);
and U25866 (N_25866,N_25717,N_25749);
xor U25867 (N_25867,N_25596,N_25688);
xnor U25868 (N_25868,N_25678,N_25567);
or U25869 (N_25869,N_25660,N_25600);
or U25870 (N_25870,N_25608,N_25509);
nor U25871 (N_25871,N_25529,N_25508);
nand U25872 (N_25872,N_25573,N_25645);
or U25873 (N_25873,N_25665,N_25589);
xnor U25874 (N_25874,N_25724,N_25661);
xor U25875 (N_25875,N_25547,N_25654);
xnor U25876 (N_25876,N_25543,N_25587);
nor U25877 (N_25877,N_25544,N_25734);
or U25878 (N_25878,N_25686,N_25501);
xor U25879 (N_25879,N_25508,N_25535);
xor U25880 (N_25880,N_25515,N_25581);
or U25881 (N_25881,N_25637,N_25501);
xor U25882 (N_25882,N_25516,N_25719);
or U25883 (N_25883,N_25530,N_25670);
or U25884 (N_25884,N_25563,N_25566);
and U25885 (N_25885,N_25628,N_25600);
and U25886 (N_25886,N_25592,N_25555);
nor U25887 (N_25887,N_25704,N_25521);
or U25888 (N_25888,N_25648,N_25618);
nor U25889 (N_25889,N_25567,N_25606);
xor U25890 (N_25890,N_25562,N_25616);
and U25891 (N_25891,N_25665,N_25606);
and U25892 (N_25892,N_25677,N_25531);
and U25893 (N_25893,N_25747,N_25647);
xor U25894 (N_25894,N_25741,N_25537);
or U25895 (N_25895,N_25560,N_25645);
xor U25896 (N_25896,N_25601,N_25735);
nor U25897 (N_25897,N_25713,N_25621);
nand U25898 (N_25898,N_25583,N_25522);
nor U25899 (N_25899,N_25678,N_25547);
nor U25900 (N_25900,N_25621,N_25607);
or U25901 (N_25901,N_25510,N_25581);
nor U25902 (N_25902,N_25579,N_25507);
xnor U25903 (N_25903,N_25512,N_25723);
or U25904 (N_25904,N_25737,N_25600);
xnor U25905 (N_25905,N_25736,N_25665);
xor U25906 (N_25906,N_25530,N_25745);
nor U25907 (N_25907,N_25553,N_25569);
xor U25908 (N_25908,N_25589,N_25696);
or U25909 (N_25909,N_25556,N_25653);
or U25910 (N_25910,N_25713,N_25566);
nand U25911 (N_25911,N_25632,N_25721);
nor U25912 (N_25912,N_25503,N_25658);
or U25913 (N_25913,N_25574,N_25535);
nor U25914 (N_25914,N_25724,N_25592);
xor U25915 (N_25915,N_25609,N_25575);
xnor U25916 (N_25916,N_25714,N_25586);
nor U25917 (N_25917,N_25746,N_25661);
xor U25918 (N_25918,N_25647,N_25668);
or U25919 (N_25919,N_25699,N_25739);
or U25920 (N_25920,N_25540,N_25667);
or U25921 (N_25921,N_25741,N_25584);
xnor U25922 (N_25922,N_25747,N_25676);
nand U25923 (N_25923,N_25512,N_25549);
nand U25924 (N_25924,N_25740,N_25615);
and U25925 (N_25925,N_25568,N_25604);
xnor U25926 (N_25926,N_25693,N_25622);
or U25927 (N_25927,N_25557,N_25710);
xor U25928 (N_25928,N_25708,N_25533);
xnor U25929 (N_25929,N_25723,N_25703);
nand U25930 (N_25930,N_25705,N_25662);
xor U25931 (N_25931,N_25560,N_25556);
xnor U25932 (N_25932,N_25621,N_25641);
nor U25933 (N_25933,N_25748,N_25660);
or U25934 (N_25934,N_25513,N_25708);
nor U25935 (N_25935,N_25541,N_25638);
and U25936 (N_25936,N_25590,N_25729);
nand U25937 (N_25937,N_25598,N_25682);
nand U25938 (N_25938,N_25624,N_25701);
and U25939 (N_25939,N_25615,N_25685);
and U25940 (N_25940,N_25647,N_25620);
and U25941 (N_25941,N_25711,N_25601);
and U25942 (N_25942,N_25610,N_25616);
and U25943 (N_25943,N_25717,N_25527);
nor U25944 (N_25944,N_25608,N_25564);
nor U25945 (N_25945,N_25704,N_25515);
or U25946 (N_25946,N_25698,N_25703);
nand U25947 (N_25947,N_25722,N_25624);
nor U25948 (N_25948,N_25595,N_25530);
or U25949 (N_25949,N_25543,N_25647);
xor U25950 (N_25950,N_25688,N_25601);
nor U25951 (N_25951,N_25697,N_25548);
nor U25952 (N_25952,N_25722,N_25720);
nor U25953 (N_25953,N_25530,N_25601);
nand U25954 (N_25954,N_25549,N_25578);
and U25955 (N_25955,N_25510,N_25573);
nand U25956 (N_25956,N_25734,N_25593);
xor U25957 (N_25957,N_25562,N_25600);
nor U25958 (N_25958,N_25537,N_25613);
xor U25959 (N_25959,N_25718,N_25661);
nand U25960 (N_25960,N_25732,N_25632);
or U25961 (N_25961,N_25551,N_25742);
nand U25962 (N_25962,N_25737,N_25653);
and U25963 (N_25963,N_25575,N_25671);
nor U25964 (N_25964,N_25606,N_25744);
or U25965 (N_25965,N_25556,N_25587);
nand U25966 (N_25966,N_25598,N_25712);
nand U25967 (N_25967,N_25667,N_25651);
nand U25968 (N_25968,N_25637,N_25728);
nor U25969 (N_25969,N_25605,N_25643);
nor U25970 (N_25970,N_25584,N_25541);
or U25971 (N_25971,N_25551,N_25719);
nor U25972 (N_25972,N_25564,N_25667);
nor U25973 (N_25973,N_25731,N_25746);
and U25974 (N_25974,N_25563,N_25723);
nand U25975 (N_25975,N_25540,N_25685);
and U25976 (N_25976,N_25678,N_25719);
xor U25977 (N_25977,N_25687,N_25576);
or U25978 (N_25978,N_25676,N_25656);
or U25979 (N_25979,N_25534,N_25531);
and U25980 (N_25980,N_25504,N_25635);
xnor U25981 (N_25981,N_25549,N_25722);
and U25982 (N_25982,N_25539,N_25697);
nand U25983 (N_25983,N_25528,N_25635);
nor U25984 (N_25984,N_25581,N_25735);
nand U25985 (N_25985,N_25539,N_25696);
nand U25986 (N_25986,N_25642,N_25664);
xor U25987 (N_25987,N_25616,N_25637);
or U25988 (N_25988,N_25655,N_25564);
nand U25989 (N_25989,N_25516,N_25693);
nand U25990 (N_25990,N_25660,N_25700);
nor U25991 (N_25991,N_25553,N_25643);
nor U25992 (N_25992,N_25604,N_25542);
nand U25993 (N_25993,N_25678,N_25597);
nor U25994 (N_25994,N_25650,N_25667);
nand U25995 (N_25995,N_25578,N_25705);
nand U25996 (N_25996,N_25594,N_25534);
and U25997 (N_25997,N_25508,N_25540);
nand U25998 (N_25998,N_25733,N_25702);
or U25999 (N_25999,N_25680,N_25676);
or U26000 (N_26000,N_25753,N_25864);
nor U26001 (N_26001,N_25893,N_25923);
or U26002 (N_26002,N_25922,N_25779);
nand U26003 (N_26003,N_25984,N_25994);
nor U26004 (N_26004,N_25979,N_25981);
nand U26005 (N_26005,N_25819,N_25868);
nand U26006 (N_26006,N_25803,N_25873);
nor U26007 (N_26007,N_25866,N_25825);
xor U26008 (N_26008,N_25885,N_25786);
nor U26009 (N_26009,N_25760,N_25863);
nand U26010 (N_26010,N_25821,N_25892);
and U26011 (N_26011,N_25982,N_25789);
xor U26012 (N_26012,N_25794,N_25816);
nand U26013 (N_26013,N_25845,N_25784);
nor U26014 (N_26014,N_25993,N_25764);
or U26015 (N_26015,N_25809,N_25822);
xor U26016 (N_26016,N_25995,N_25850);
nor U26017 (N_26017,N_25909,N_25962);
or U26018 (N_26018,N_25943,N_25990);
nand U26019 (N_26019,N_25769,N_25948);
nor U26020 (N_26020,N_25897,N_25757);
or U26021 (N_26021,N_25840,N_25793);
nand U26022 (N_26022,N_25936,N_25971);
and U26023 (N_26023,N_25901,N_25826);
nor U26024 (N_26024,N_25972,N_25991);
nand U26025 (N_26025,N_25983,N_25950);
or U26026 (N_26026,N_25841,N_25765);
nor U26027 (N_26027,N_25925,N_25961);
and U26028 (N_26028,N_25878,N_25859);
and U26029 (N_26029,N_25912,N_25951);
nand U26030 (N_26030,N_25785,N_25813);
or U26031 (N_26031,N_25879,N_25896);
nor U26032 (N_26032,N_25823,N_25883);
nor U26033 (N_26033,N_25906,N_25921);
and U26034 (N_26034,N_25941,N_25790);
nor U26035 (N_26035,N_25882,N_25932);
and U26036 (N_26036,N_25999,N_25768);
nor U26037 (N_26037,N_25829,N_25902);
xor U26038 (N_26038,N_25931,N_25774);
xnor U26039 (N_26039,N_25810,N_25988);
nor U26040 (N_26040,N_25942,N_25820);
xor U26041 (N_26041,N_25926,N_25792);
nand U26042 (N_26042,N_25959,N_25814);
xnor U26043 (N_26043,N_25875,N_25957);
nand U26044 (N_26044,N_25759,N_25857);
nand U26045 (N_26045,N_25937,N_25754);
nand U26046 (N_26046,N_25869,N_25985);
nand U26047 (N_26047,N_25751,N_25853);
nand U26048 (N_26048,N_25846,N_25976);
nand U26049 (N_26049,N_25838,N_25967);
xnor U26050 (N_26050,N_25817,N_25917);
or U26051 (N_26051,N_25977,N_25781);
and U26052 (N_26052,N_25904,N_25807);
nor U26053 (N_26053,N_25938,N_25755);
xor U26054 (N_26054,N_25954,N_25964);
or U26055 (N_26055,N_25911,N_25837);
or U26056 (N_26056,N_25916,N_25898);
nor U26057 (N_26057,N_25815,N_25812);
xnor U26058 (N_26058,N_25867,N_25858);
or U26059 (N_26059,N_25766,N_25920);
xnor U26060 (N_26060,N_25783,N_25870);
nand U26061 (N_26061,N_25918,N_25960);
nor U26062 (N_26062,N_25856,N_25796);
nand U26063 (N_26063,N_25855,N_25876);
nor U26064 (N_26064,N_25986,N_25861);
or U26065 (N_26065,N_25927,N_25787);
xor U26066 (N_26066,N_25848,N_25802);
nand U26067 (N_26067,N_25884,N_25992);
nand U26068 (N_26068,N_25956,N_25772);
nand U26069 (N_26069,N_25903,N_25890);
and U26070 (N_26070,N_25777,N_25928);
or U26071 (N_26071,N_25933,N_25804);
xor U26072 (N_26072,N_25862,N_25877);
xor U26073 (N_26073,N_25924,N_25907);
xnor U26074 (N_26074,N_25908,N_25805);
and U26075 (N_26075,N_25762,N_25778);
or U26076 (N_26076,N_25899,N_25895);
xor U26077 (N_26077,N_25914,N_25871);
nor U26078 (N_26078,N_25944,N_25860);
nand U26079 (N_26079,N_25808,N_25970);
nand U26080 (N_26080,N_25996,N_25974);
or U26081 (N_26081,N_25839,N_25791);
nand U26082 (N_26082,N_25797,N_25827);
and U26083 (N_26083,N_25763,N_25989);
and U26084 (N_26084,N_25750,N_25968);
and U26085 (N_26085,N_25780,N_25915);
and U26086 (N_26086,N_25872,N_25930);
nor U26087 (N_26087,N_25844,N_25886);
or U26088 (N_26088,N_25842,N_25946);
nor U26089 (N_26089,N_25913,N_25824);
nor U26090 (N_26090,N_25940,N_25900);
and U26091 (N_26091,N_25758,N_25880);
xor U26092 (N_26092,N_25929,N_25773);
and U26093 (N_26093,N_25831,N_25834);
or U26094 (N_26094,N_25767,N_25854);
xor U26095 (N_26095,N_25771,N_25800);
and U26096 (N_26096,N_25889,N_25836);
or U26097 (N_26097,N_25955,N_25828);
and U26098 (N_26098,N_25958,N_25756);
nor U26099 (N_26099,N_25953,N_25934);
nor U26100 (N_26100,N_25761,N_25833);
nor U26101 (N_26101,N_25752,N_25775);
nand U26102 (N_26102,N_25782,N_25947);
or U26103 (N_26103,N_25939,N_25806);
xor U26104 (N_26104,N_25949,N_25894);
nor U26105 (N_26105,N_25865,N_25965);
xnor U26106 (N_26106,N_25910,N_25818);
xor U26107 (N_26107,N_25966,N_25952);
and U26108 (N_26108,N_25776,N_25987);
nor U26109 (N_26109,N_25919,N_25835);
and U26110 (N_26110,N_25881,N_25830);
nand U26111 (N_26111,N_25935,N_25770);
xnor U26112 (N_26112,N_25851,N_25998);
nand U26113 (N_26113,N_25888,N_25795);
nor U26114 (N_26114,N_25973,N_25798);
xnor U26115 (N_26115,N_25975,N_25887);
or U26116 (N_26116,N_25978,N_25980);
nand U26117 (N_26117,N_25905,N_25849);
nand U26118 (N_26118,N_25832,N_25799);
xnor U26119 (N_26119,N_25997,N_25843);
and U26120 (N_26120,N_25847,N_25891);
xor U26121 (N_26121,N_25811,N_25963);
or U26122 (N_26122,N_25969,N_25945);
and U26123 (N_26123,N_25801,N_25788);
or U26124 (N_26124,N_25852,N_25874);
nor U26125 (N_26125,N_25912,N_25811);
xnor U26126 (N_26126,N_25880,N_25838);
nor U26127 (N_26127,N_25887,N_25906);
and U26128 (N_26128,N_25928,N_25903);
xnor U26129 (N_26129,N_25974,N_25795);
or U26130 (N_26130,N_25810,N_25872);
nand U26131 (N_26131,N_25766,N_25875);
or U26132 (N_26132,N_25983,N_25809);
or U26133 (N_26133,N_25899,N_25906);
and U26134 (N_26134,N_25853,N_25902);
xor U26135 (N_26135,N_25772,N_25862);
and U26136 (N_26136,N_25752,N_25973);
nor U26137 (N_26137,N_25914,N_25918);
and U26138 (N_26138,N_25865,N_25823);
xnor U26139 (N_26139,N_25941,N_25894);
nor U26140 (N_26140,N_25909,N_25903);
and U26141 (N_26141,N_25958,N_25776);
or U26142 (N_26142,N_25949,N_25846);
nor U26143 (N_26143,N_25859,N_25799);
nand U26144 (N_26144,N_25818,N_25756);
nor U26145 (N_26145,N_25780,N_25879);
and U26146 (N_26146,N_25839,N_25850);
and U26147 (N_26147,N_25752,N_25800);
nor U26148 (N_26148,N_25957,N_25894);
nand U26149 (N_26149,N_25828,N_25883);
nand U26150 (N_26150,N_25889,N_25941);
and U26151 (N_26151,N_25937,N_25901);
xor U26152 (N_26152,N_25933,N_25952);
and U26153 (N_26153,N_25810,N_25829);
and U26154 (N_26154,N_25961,N_25921);
xor U26155 (N_26155,N_25980,N_25891);
and U26156 (N_26156,N_25932,N_25910);
or U26157 (N_26157,N_25810,N_25769);
or U26158 (N_26158,N_25883,N_25965);
nand U26159 (N_26159,N_25930,N_25932);
nand U26160 (N_26160,N_25770,N_25857);
or U26161 (N_26161,N_25936,N_25796);
nand U26162 (N_26162,N_25832,N_25986);
nand U26163 (N_26163,N_25800,N_25893);
xnor U26164 (N_26164,N_25978,N_25841);
or U26165 (N_26165,N_25889,N_25939);
xnor U26166 (N_26166,N_25798,N_25882);
nand U26167 (N_26167,N_25877,N_25959);
xnor U26168 (N_26168,N_25835,N_25756);
or U26169 (N_26169,N_25843,N_25944);
xnor U26170 (N_26170,N_25924,N_25823);
xnor U26171 (N_26171,N_25879,N_25831);
nor U26172 (N_26172,N_25946,N_25897);
xnor U26173 (N_26173,N_25891,N_25821);
xnor U26174 (N_26174,N_25840,N_25974);
and U26175 (N_26175,N_25770,N_25751);
nand U26176 (N_26176,N_25770,N_25848);
xnor U26177 (N_26177,N_25998,N_25873);
nor U26178 (N_26178,N_25828,N_25942);
or U26179 (N_26179,N_25789,N_25807);
and U26180 (N_26180,N_25778,N_25819);
xor U26181 (N_26181,N_25801,N_25867);
or U26182 (N_26182,N_25834,N_25927);
or U26183 (N_26183,N_25807,N_25841);
nor U26184 (N_26184,N_25880,N_25853);
nand U26185 (N_26185,N_25804,N_25869);
xnor U26186 (N_26186,N_25877,N_25896);
xnor U26187 (N_26187,N_25793,N_25900);
or U26188 (N_26188,N_25862,N_25916);
or U26189 (N_26189,N_25785,N_25882);
or U26190 (N_26190,N_25786,N_25803);
nand U26191 (N_26191,N_25860,N_25927);
and U26192 (N_26192,N_25965,N_25768);
nor U26193 (N_26193,N_25902,N_25961);
and U26194 (N_26194,N_25920,N_25856);
xor U26195 (N_26195,N_25762,N_25921);
or U26196 (N_26196,N_25764,N_25958);
or U26197 (N_26197,N_25774,N_25972);
xnor U26198 (N_26198,N_25931,N_25896);
and U26199 (N_26199,N_25951,N_25930);
nand U26200 (N_26200,N_25826,N_25890);
xor U26201 (N_26201,N_25791,N_25975);
or U26202 (N_26202,N_25914,N_25770);
nor U26203 (N_26203,N_25794,N_25929);
or U26204 (N_26204,N_25945,N_25927);
nor U26205 (N_26205,N_25924,N_25880);
and U26206 (N_26206,N_25818,N_25783);
nand U26207 (N_26207,N_25800,N_25765);
and U26208 (N_26208,N_25898,N_25821);
xnor U26209 (N_26209,N_25904,N_25951);
or U26210 (N_26210,N_25843,N_25987);
or U26211 (N_26211,N_25833,N_25927);
or U26212 (N_26212,N_25750,N_25916);
nor U26213 (N_26213,N_25851,N_25911);
nand U26214 (N_26214,N_25880,N_25852);
or U26215 (N_26215,N_25999,N_25857);
and U26216 (N_26216,N_25989,N_25972);
xnor U26217 (N_26217,N_25912,N_25958);
xnor U26218 (N_26218,N_25928,N_25943);
nand U26219 (N_26219,N_25927,N_25795);
or U26220 (N_26220,N_25877,N_25863);
nand U26221 (N_26221,N_25851,N_25790);
nand U26222 (N_26222,N_25933,N_25795);
nand U26223 (N_26223,N_25844,N_25977);
nor U26224 (N_26224,N_25944,N_25857);
or U26225 (N_26225,N_25757,N_25830);
nor U26226 (N_26226,N_25973,N_25876);
xor U26227 (N_26227,N_25914,N_25840);
nand U26228 (N_26228,N_25818,N_25949);
or U26229 (N_26229,N_25878,N_25996);
or U26230 (N_26230,N_25871,N_25937);
nand U26231 (N_26231,N_25841,N_25917);
xor U26232 (N_26232,N_25775,N_25846);
or U26233 (N_26233,N_25937,N_25858);
nand U26234 (N_26234,N_25798,N_25788);
xor U26235 (N_26235,N_25781,N_25921);
xor U26236 (N_26236,N_25859,N_25873);
and U26237 (N_26237,N_25860,N_25851);
or U26238 (N_26238,N_25812,N_25963);
or U26239 (N_26239,N_25799,N_25803);
or U26240 (N_26240,N_25910,N_25751);
and U26241 (N_26241,N_25948,N_25845);
xor U26242 (N_26242,N_25820,N_25841);
nand U26243 (N_26243,N_25963,N_25896);
nor U26244 (N_26244,N_25759,N_25836);
nor U26245 (N_26245,N_25978,N_25893);
nor U26246 (N_26246,N_25888,N_25931);
nand U26247 (N_26247,N_25983,N_25915);
xor U26248 (N_26248,N_25764,N_25938);
nor U26249 (N_26249,N_25977,N_25975);
nor U26250 (N_26250,N_26223,N_26081);
and U26251 (N_26251,N_26002,N_26117);
and U26252 (N_26252,N_26077,N_26134);
and U26253 (N_26253,N_26114,N_26218);
nor U26254 (N_26254,N_26057,N_26173);
and U26255 (N_26255,N_26084,N_26155);
or U26256 (N_26256,N_26040,N_26124);
xor U26257 (N_26257,N_26188,N_26098);
nand U26258 (N_26258,N_26185,N_26079);
nand U26259 (N_26259,N_26242,N_26176);
nor U26260 (N_26260,N_26201,N_26128);
or U26261 (N_26261,N_26133,N_26142);
nor U26262 (N_26262,N_26145,N_26011);
xnor U26263 (N_26263,N_26249,N_26052);
xor U26264 (N_26264,N_26048,N_26206);
xor U26265 (N_26265,N_26127,N_26065);
or U26266 (N_26266,N_26049,N_26154);
and U26267 (N_26267,N_26225,N_26097);
nor U26268 (N_26268,N_26083,N_26119);
and U26269 (N_26269,N_26203,N_26181);
or U26270 (N_26270,N_26168,N_26159);
nand U26271 (N_26271,N_26023,N_26056);
xor U26272 (N_26272,N_26208,N_26088);
nand U26273 (N_26273,N_26004,N_26059);
and U26274 (N_26274,N_26175,N_26042);
and U26275 (N_26275,N_26003,N_26073);
nand U26276 (N_26276,N_26019,N_26179);
nor U26277 (N_26277,N_26246,N_26021);
nor U26278 (N_26278,N_26099,N_26162);
nand U26279 (N_26279,N_26029,N_26227);
and U26280 (N_26280,N_26146,N_26041);
xor U26281 (N_26281,N_26123,N_26122);
nor U26282 (N_26282,N_26207,N_26110);
nand U26283 (N_26283,N_26091,N_26007);
and U26284 (N_26284,N_26180,N_26022);
or U26285 (N_26285,N_26060,N_26183);
or U26286 (N_26286,N_26095,N_26116);
nand U26287 (N_26287,N_26164,N_26093);
nor U26288 (N_26288,N_26037,N_26047);
nand U26289 (N_26289,N_26121,N_26141);
nand U26290 (N_26290,N_26221,N_26213);
xnor U26291 (N_26291,N_26120,N_26187);
xnor U26292 (N_26292,N_26070,N_26196);
and U26293 (N_26293,N_26232,N_26131);
xor U26294 (N_26294,N_26100,N_26222);
or U26295 (N_26295,N_26241,N_26199);
or U26296 (N_26296,N_26171,N_26076);
xnor U26297 (N_26297,N_26143,N_26158);
nand U26298 (N_26298,N_26036,N_26032);
nor U26299 (N_26299,N_26126,N_26205);
nor U26300 (N_26300,N_26184,N_26226);
nor U26301 (N_26301,N_26139,N_26054);
xnor U26302 (N_26302,N_26072,N_26028);
xor U26303 (N_26303,N_26010,N_26229);
nand U26304 (N_26304,N_26062,N_26166);
xnor U26305 (N_26305,N_26024,N_26220);
nand U26306 (N_26306,N_26151,N_26216);
or U26307 (N_26307,N_26219,N_26129);
nor U26308 (N_26308,N_26152,N_26160);
nor U26309 (N_26309,N_26106,N_26174);
xnor U26310 (N_26310,N_26027,N_26058);
or U26311 (N_26311,N_26214,N_26016);
nor U26312 (N_26312,N_26140,N_26005);
xor U26313 (N_26313,N_26061,N_26118);
nor U26314 (N_26314,N_26192,N_26104);
nor U26315 (N_26315,N_26244,N_26012);
and U26316 (N_26316,N_26115,N_26069);
and U26317 (N_26317,N_26045,N_26235);
nand U26318 (N_26318,N_26228,N_26063);
and U26319 (N_26319,N_26215,N_26148);
nor U26320 (N_26320,N_26243,N_26178);
xor U26321 (N_26321,N_26198,N_26210);
or U26322 (N_26322,N_26038,N_26013);
and U26323 (N_26323,N_26245,N_26092);
nor U26324 (N_26324,N_26169,N_26202);
or U26325 (N_26325,N_26177,N_26138);
nor U26326 (N_26326,N_26051,N_26043);
and U26327 (N_26327,N_26066,N_26186);
and U26328 (N_26328,N_26111,N_26153);
nand U26329 (N_26329,N_26240,N_26071);
nand U26330 (N_26330,N_26087,N_26195);
and U26331 (N_26331,N_26105,N_26033);
nand U26332 (N_26332,N_26014,N_26086);
or U26333 (N_26333,N_26191,N_26112);
and U26334 (N_26334,N_26020,N_26034);
xor U26335 (N_26335,N_26064,N_26094);
nor U26336 (N_26336,N_26035,N_26075);
or U26337 (N_26337,N_26082,N_26046);
nor U26338 (N_26338,N_26090,N_26039);
nor U26339 (N_26339,N_26190,N_26130);
and U26340 (N_26340,N_26247,N_26231);
or U26341 (N_26341,N_26103,N_26108);
or U26342 (N_26342,N_26006,N_26189);
or U26343 (N_26343,N_26053,N_26001);
nor U26344 (N_26344,N_26209,N_26074);
or U26345 (N_26345,N_26211,N_26167);
nor U26346 (N_26346,N_26236,N_26136);
nor U26347 (N_26347,N_26101,N_26015);
nor U26348 (N_26348,N_26234,N_26200);
nand U26349 (N_26349,N_26217,N_26239);
nand U26350 (N_26350,N_26031,N_26237);
nand U26351 (N_26351,N_26067,N_26080);
nand U26352 (N_26352,N_26147,N_26050);
and U26353 (N_26353,N_26044,N_26230);
or U26354 (N_26354,N_26156,N_26085);
xnor U26355 (N_26355,N_26165,N_26089);
xnor U26356 (N_26356,N_26248,N_26204);
or U26357 (N_26357,N_26030,N_26163);
nand U26358 (N_26358,N_26132,N_26008);
nand U26359 (N_26359,N_26157,N_26233);
and U26360 (N_26360,N_26068,N_26144);
nor U26361 (N_26361,N_26170,N_26212);
or U26362 (N_26362,N_26137,N_26000);
and U26363 (N_26363,N_26009,N_26135);
or U26364 (N_26364,N_26238,N_26182);
nand U26365 (N_26365,N_26025,N_26107);
nor U26366 (N_26366,N_26078,N_26109);
nor U26367 (N_26367,N_26125,N_26017);
nand U26368 (N_26368,N_26102,N_26197);
or U26369 (N_26369,N_26172,N_26193);
or U26370 (N_26370,N_26113,N_26194);
xnor U26371 (N_26371,N_26161,N_26150);
or U26372 (N_26372,N_26149,N_26096);
xnor U26373 (N_26373,N_26018,N_26224);
xor U26374 (N_26374,N_26055,N_26026);
xor U26375 (N_26375,N_26017,N_26208);
xnor U26376 (N_26376,N_26219,N_26153);
or U26377 (N_26377,N_26169,N_26143);
or U26378 (N_26378,N_26154,N_26209);
xor U26379 (N_26379,N_26152,N_26148);
or U26380 (N_26380,N_26155,N_26154);
or U26381 (N_26381,N_26071,N_26160);
nor U26382 (N_26382,N_26160,N_26211);
or U26383 (N_26383,N_26176,N_26212);
xnor U26384 (N_26384,N_26056,N_26008);
nand U26385 (N_26385,N_26145,N_26240);
nand U26386 (N_26386,N_26229,N_26066);
xor U26387 (N_26387,N_26005,N_26241);
xnor U26388 (N_26388,N_26061,N_26192);
nor U26389 (N_26389,N_26222,N_26121);
nor U26390 (N_26390,N_26207,N_26225);
or U26391 (N_26391,N_26092,N_26176);
nor U26392 (N_26392,N_26204,N_26067);
nand U26393 (N_26393,N_26090,N_26117);
xnor U26394 (N_26394,N_26172,N_26213);
and U26395 (N_26395,N_26126,N_26219);
nand U26396 (N_26396,N_26010,N_26149);
or U26397 (N_26397,N_26034,N_26075);
or U26398 (N_26398,N_26037,N_26019);
nand U26399 (N_26399,N_26241,N_26245);
nand U26400 (N_26400,N_26153,N_26186);
nand U26401 (N_26401,N_26187,N_26049);
xor U26402 (N_26402,N_26133,N_26022);
nor U26403 (N_26403,N_26171,N_26035);
and U26404 (N_26404,N_26206,N_26140);
nor U26405 (N_26405,N_26136,N_26065);
xor U26406 (N_26406,N_26042,N_26236);
nand U26407 (N_26407,N_26151,N_26093);
and U26408 (N_26408,N_26053,N_26232);
nor U26409 (N_26409,N_26117,N_26100);
and U26410 (N_26410,N_26125,N_26048);
and U26411 (N_26411,N_26055,N_26221);
nor U26412 (N_26412,N_26066,N_26033);
or U26413 (N_26413,N_26077,N_26167);
nand U26414 (N_26414,N_26073,N_26055);
xor U26415 (N_26415,N_26016,N_26150);
or U26416 (N_26416,N_26165,N_26031);
nand U26417 (N_26417,N_26096,N_26022);
nor U26418 (N_26418,N_26207,N_26178);
nor U26419 (N_26419,N_26241,N_26034);
xnor U26420 (N_26420,N_26230,N_26040);
nand U26421 (N_26421,N_26078,N_26240);
and U26422 (N_26422,N_26130,N_26024);
and U26423 (N_26423,N_26031,N_26064);
xor U26424 (N_26424,N_26000,N_26050);
nand U26425 (N_26425,N_26007,N_26068);
or U26426 (N_26426,N_26119,N_26195);
nor U26427 (N_26427,N_26073,N_26029);
and U26428 (N_26428,N_26203,N_26129);
and U26429 (N_26429,N_26149,N_26204);
xnor U26430 (N_26430,N_26083,N_26100);
xnor U26431 (N_26431,N_26101,N_26137);
nor U26432 (N_26432,N_26152,N_26103);
xor U26433 (N_26433,N_26127,N_26149);
nand U26434 (N_26434,N_26049,N_26081);
nor U26435 (N_26435,N_26168,N_26127);
nor U26436 (N_26436,N_26211,N_26030);
and U26437 (N_26437,N_26157,N_26062);
nand U26438 (N_26438,N_26146,N_26004);
xor U26439 (N_26439,N_26162,N_26001);
nor U26440 (N_26440,N_26148,N_26153);
or U26441 (N_26441,N_26090,N_26142);
and U26442 (N_26442,N_26175,N_26151);
or U26443 (N_26443,N_26043,N_26235);
nor U26444 (N_26444,N_26007,N_26174);
nand U26445 (N_26445,N_26124,N_26041);
or U26446 (N_26446,N_26003,N_26199);
and U26447 (N_26447,N_26028,N_26119);
xor U26448 (N_26448,N_26002,N_26009);
nand U26449 (N_26449,N_26178,N_26142);
or U26450 (N_26450,N_26049,N_26038);
and U26451 (N_26451,N_26082,N_26203);
xor U26452 (N_26452,N_26153,N_26197);
and U26453 (N_26453,N_26102,N_26097);
or U26454 (N_26454,N_26152,N_26094);
xnor U26455 (N_26455,N_26119,N_26045);
and U26456 (N_26456,N_26063,N_26180);
and U26457 (N_26457,N_26085,N_26135);
nor U26458 (N_26458,N_26049,N_26134);
nand U26459 (N_26459,N_26190,N_26067);
or U26460 (N_26460,N_26226,N_26157);
or U26461 (N_26461,N_26226,N_26098);
or U26462 (N_26462,N_26202,N_26117);
nand U26463 (N_26463,N_26114,N_26051);
and U26464 (N_26464,N_26023,N_26155);
and U26465 (N_26465,N_26149,N_26153);
and U26466 (N_26466,N_26018,N_26077);
xor U26467 (N_26467,N_26150,N_26097);
and U26468 (N_26468,N_26077,N_26080);
and U26469 (N_26469,N_26018,N_26045);
nor U26470 (N_26470,N_26045,N_26216);
and U26471 (N_26471,N_26114,N_26084);
xnor U26472 (N_26472,N_26147,N_26064);
xor U26473 (N_26473,N_26014,N_26031);
and U26474 (N_26474,N_26156,N_26225);
xor U26475 (N_26475,N_26212,N_26049);
and U26476 (N_26476,N_26197,N_26041);
and U26477 (N_26477,N_26115,N_26174);
xor U26478 (N_26478,N_26070,N_26135);
and U26479 (N_26479,N_26224,N_26240);
nand U26480 (N_26480,N_26095,N_26167);
nand U26481 (N_26481,N_26114,N_26060);
nand U26482 (N_26482,N_26084,N_26206);
xnor U26483 (N_26483,N_26169,N_26168);
nand U26484 (N_26484,N_26024,N_26171);
and U26485 (N_26485,N_26172,N_26114);
and U26486 (N_26486,N_26224,N_26112);
and U26487 (N_26487,N_26174,N_26000);
nor U26488 (N_26488,N_26058,N_26020);
nand U26489 (N_26489,N_26089,N_26001);
xor U26490 (N_26490,N_26242,N_26222);
nor U26491 (N_26491,N_26104,N_26206);
or U26492 (N_26492,N_26249,N_26107);
nand U26493 (N_26493,N_26172,N_26014);
xor U26494 (N_26494,N_26046,N_26110);
or U26495 (N_26495,N_26085,N_26086);
nor U26496 (N_26496,N_26122,N_26164);
nor U26497 (N_26497,N_26047,N_26098);
xor U26498 (N_26498,N_26094,N_26070);
nand U26499 (N_26499,N_26134,N_26217);
or U26500 (N_26500,N_26380,N_26493);
nor U26501 (N_26501,N_26338,N_26487);
and U26502 (N_26502,N_26444,N_26401);
xor U26503 (N_26503,N_26461,N_26426);
and U26504 (N_26504,N_26397,N_26387);
nor U26505 (N_26505,N_26396,N_26381);
and U26506 (N_26506,N_26349,N_26368);
and U26507 (N_26507,N_26433,N_26436);
nor U26508 (N_26508,N_26498,N_26364);
xor U26509 (N_26509,N_26463,N_26253);
or U26510 (N_26510,N_26298,N_26252);
nand U26511 (N_26511,N_26443,N_26317);
and U26512 (N_26512,N_26475,N_26330);
and U26513 (N_26513,N_26263,N_26371);
or U26514 (N_26514,N_26407,N_26250);
nor U26515 (N_26515,N_26499,N_26476);
and U26516 (N_26516,N_26469,N_26313);
or U26517 (N_26517,N_26315,N_26255);
and U26518 (N_26518,N_26382,N_26296);
nor U26519 (N_26519,N_26425,N_26442);
or U26520 (N_26520,N_26483,N_26404);
nand U26521 (N_26521,N_26405,N_26283);
and U26522 (N_26522,N_26366,N_26266);
and U26523 (N_26523,N_26280,N_26327);
and U26524 (N_26524,N_26299,N_26354);
xor U26525 (N_26525,N_26282,N_26312);
xor U26526 (N_26526,N_26441,N_26251);
and U26527 (N_26527,N_26448,N_26357);
nand U26528 (N_26528,N_26489,N_26383);
nand U26529 (N_26529,N_26309,N_26413);
nor U26530 (N_26530,N_26390,N_26477);
or U26531 (N_26531,N_26468,N_26272);
xnor U26532 (N_26532,N_26496,N_26322);
nand U26533 (N_26533,N_26286,N_26486);
or U26534 (N_26534,N_26423,N_26437);
or U26535 (N_26535,N_26325,N_26321);
nor U26536 (N_26536,N_26399,N_26347);
and U26537 (N_26537,N_26302,N_26395);
nor U26538 (N_26538,N_26379,N_26361);
xnor U26539 (N_26539,N_26278,N_26454);
and U26540 (N_26540,N_26424,N_26478);
nand U26541 (N_26541,N_26398,N_26301);
or U26542 (N_26542,N_26481,N_26440);
nand U26543 (N_26543,N_26324,N_26473);
xnor U26544 (N_26544,N_26400,N_26447);
xnor U26545 (N_26545,N_26259,N_26377);
nand U26546 (N_26546,N_26295,N_26284);
or U26547 (N_26547,N_26258,N_26374);
nor U26548 (N_26548,N_26262,N_26351);
xnor U26549 (N_26549,N_26432,N_26455);
or U26550 (N_26550,N_26288,N_26488);
and U26551 (N_26551,N_26445,N_26466);
xor U26552 (N_26552,N_26328,N_26406);
nand U26553 (N_26553,N_26453,N_26431);
nor U26554 (N_26554,N_26345,N_26450);
or U26555 (N_26555,N_26305,N_26490);
nor U26556 (N_26556,N_26464,N_26402);
or U26557 (N_26557,N_26269,N_26342);
nand U26558 (N_26558,N_26416,N_26427);
nand U26559 (N_26559,N_26409,N_26285);
nand U26560 (N_26560,N_26316,N_26393);
xor U26561 (N_26561,N_26287,N_26429);
nand U26562 (N_26562,N_26273,N_26420);
and U26563 (N_26563,N_26408,N_26438);
nand U26564 (N_26564,N_26360,N_26430);
nand U26565 (N_26565,N_26276,N_26449);
or U26566 (N_26566,N_26497,N_26365);
nand U26567 (N_26567,N_26257,N_26358);
xor U26568 (N_26568,N_26419,N_26310);
nand U26569 (N_26569,N_26293,N_26378);
nand U26570 (N_26570,N_26352,N_26465);
nor U26571 (N_26571,N_26462,N_26350);
xor U26572 (N_26572,N_26346,N_26412);
nor U26573 (N_26573,N_26271,N_26275);
xnor U26574 (N_26574,N_26318,N_26484);
and U26575 (N_26575,N_26292,N_26434);
nand U26576 (N_26576,N_26332,N_26348);
nor U26577 (N_26577,N_26356,N_26392);
nand U26578 (N_26578,N_26491,N_26308);
nor U26579 (N_26579,N_26362,N_26270);
or U26580 (N_26580,N_26485,N_26474);
xor U26581 (N_26581,N_26303,N_26341);
nand U26582 (N_26582,N_26254,N_26337);
nand U26583 (N_26583,N_26300,N_26331);
nor U26584 (N_26584,N_26319,N_26470);
xor U26585 (N_26585,N_26297,N_26479);
xnor U26586 (N_26586,N_26394,N_26385);
and U26587 (N_26587,N_26265,N_26334);
and U26588 (N_26588,N_26472,N_26340);
and U26589 (N_26589,N_26304,N_26267);
nor U26590 (N_26590,N_26333,N_26277);
and U26591 (N_26591,N_26320,N_26307);
nor U26592 (N_26592,N_26290,N_26281);
nand U26593 (N_26593,N_26375,N_26311);
and U26594 (N_26594,N_26494,N_26336);
and U26595 (N_26595,N_26435,N_26456);
and U26596 (N_26596,N_26482,N_26480);
nand U26597 (N_26597,N_26384,N_26274);
or U26598 (N_26598,N_26422,N_26471);
or U26599 (N_26599,N_26289,N_26355);
nor U26600 (N_26600,N_26344,N_26264);
and U26601 (N_26601,N_26467,N_26411);
and U26602 (N_26602,N_26373,N_26279);
or U26603 (N_26603,N_26459,N_26326);
nand U26604 (N_26604,N_26268,N_26415);
xor U26605 (N_26605,N_26460,N_26495);
nor U26606 (N_26606,N_26446,N_26359);
xnor U26607 (N_26607,N_26391,N_26418);
nor U26608 (N_26608,N_26372,N_26389);
xnor U26609 (N_26609,N_26439,N_26329);
and U26610 (N_26610,N_26291,N_26335);
xor U26611 (N_26611,N_26451,N_26370);
nand U26612 (N_26612,N_26410,N_26256);
and U26613 (N_26613,N_26492,N_26369);
and U26614 (N_26614,N_26417,N_26386);
and U26615 (N_26615,N_26428,N_26452);
and U26616 (N_26616,N_26414,N_26339);
or U26617 (N_26617,N_26294,N_26363);
nand U26618 (N_26618,N_26403,N_26458);
nor U26619 (N_26619,N_26343,N_26376);
xnor U26620 (N_26620,N_26314,N_26388);
or U26621 (N_26621,N_26306,N_26457);
or U26622 (N_26622,N_26367,N_26421);
xor U26623 (N_26623,N_26261,N_26353);
and U26624 (N_26624,N_26323,N_26260);
and U26625 (N_26625,N_26346,N_26409);
nor U26626 (N_26626,N_26364,N_26291);
xnor U26627 (N_26627,N_26412,N_26275);
nor U26628 (N_26628,N_26344,N_26266);
or U26629 (N_26629,N_26324,N_26361);
and U26630 (N_26630,N_26395,N_26320);
nand U26631 (N_26631,N_26315,N_26325);
xnor U26632 (N_26632,N_26332,N_26377);
nor U26633 (N_26633,N_26355,N_26331);
or U26634 (N_26634,N_26401,N_26426);
or U26635 (N_26635,N_26403,N_26456);
or U26636 (N_26636,N_26291,N_26338);
and U26637 (N_26637,N_26277,N_26258);
nand U26638 (N_26638,N_26482,N_26464);
and U26639 (N_26639,N_26296,N_26284);
or U26640 (N_26640,N_26390,N_26452);
nor U26641 (N_26641,N_26321,N_26412);
and U26642 (N_26642,N_26373,N_26437);
and U26643 (N_26643,N_26418,N_26443);
nor U26644 (N_26644,N_26385,N_26474);
and U26645 (N_26645,N_26350,N_26405);
nand U26646 (N_26646,N_26276,N_26382);
nor U26647 (N_26647,N_26405,N_26495);
nor U26648 (N_26648,N_26453,N_26417);
or U26649 (N_26649,N_26274,N_26480);
nor U26650 (N_26650,N_26418,N_26289);
xor U26651 (N_26651,N_26259,N_26408);
and U26652 (N_26652,N_26314,N_26382);
and U26653 (N_26653,N_26424,N_26301);
nor U26654 (N_26654,N_26301,N_26346);
nand U26655 (N_26655,N_26420,N_26473);
nand U26656 (N_26656,N_26452,N_26404);
xnor U26657 (N_26657,N_26363,N_26461);
nand U26658 (N_26658,N_26312,N_26319);
or U26659 (N_26659,N_26307,N_26482);
and U26660 (N_26660,N_26311,N_26371);
or U26661 (N_26661,N_26363,N_26484);
nor U26662 (N_26662,N_26344,N_26276);
xor U26663 (N_26663,N_26445,N_26290);
xor U26664 (N_26664,N_26374,N_26250);
nor U26665 (N_26665,N_26410,N_26317);
nor U26666 (N_26666,N_26285,N_26326);
nor U26667 (N_26667,N_26364,N_26377);
and U26668 (N_26668,N_26272,N_26374);
nor U26669 (N_26669,N_26397,N_26280);
and U26670 (N_26670,N_26443,N_26377);
or U26671 (N_26671,N_26254,N_26308);
and U26672 (N_26672,N_26263,N_26412);
xor U26673 (N_26673,N_26326,N_26291);
nand U26674 (N_26674,N_26341,N_26429);
and U26675 (N_26675,N_26467,N_26489);
or U26676 (N_26676,N_26337,N_26387);
and U26677 (N_26677,N_26370,N_26312);
xor U26678 (N_26678,N_26402,N_26468);
or U26679 (N_26679,N_26263,N_26433);
or U26680 (N_26680,N_26326,N_26396);
and U26681 (N_26681,N_26414,N_26400);
xor U26682 (N_26682,N_26349,N_26432);
xnor U26683 (N_26683,N_26343,N_26434);
nor U26684 (N_26684,N_26325,N_26473);
nor U26685 (N_26685,N_26490,N_26404);
or U26686 (N_26686,N_26405,N_26472);
or U26687 (N_26687,N_26409,N_26380);
nor U26688 (N_26688,N_26462,N_26481);
xnor U26689 (N_26689,N_26429,N_26264);
xnor U26690 (N_26690,N_26401,N_26433);
or U26691 (N_26691,N_26347,N_26411);
and U26692 (N_26692,N_26261,N_26379);
nor U26693 (N_26693,N_26338,N_26383);
and U26694 (N_26694,N_26461,N_26290);
xnor U26695 (N_26695,N_26404,N_26432);
or U26696 (N_26696,N_26376,N_26288);
nor U26697 (N_26697,N_26422,N_26459);
xnor U26698 (N_26698,N_26310,N_26339);
and U26699 (N_26699,N_26418,N_26264);
and U26700 (N_26700,N_26350,N_26364);
or U26701 (N_26701,N_26277,N_26407);
xnor U26702 (N_26702,N_26292,N_26420);
nand U26703 (N_26703,N_26494,N_26388);
or U26704 (N_26704,N_26263,N_26280);
xor U26705 (N_26705,N_26378,N_26298);
or U26706 (N_26706,N_26297,N_26443);
nor U26707 (N_26707,N_26382,N_26451);
nor U26708 (N_26708,N_26436,N_26274);
or U26709 (N_26709,N_26360,N_26274);
and U26710 (N_26710,N_26301,N_26349);
nand U26711 (N_26711,N_26344,N_26466);
nand U26712 (N_26712,N_26396,N_26316);
xnor U26713 (N_26713,N_26486,N_26480);
and U26714 (N_26714,N_26255,N_26281);
and U26715 (N_26715,N_26448,N_26435);
xnor U26716 (N_26716,N_26492,N_26286);
nor U26717 (N_26717,N_26332,N_26318);
and U26718 (N_26718,N_26438,N_26483);
and U26719 (N_26719,N_26340,N_26385);
or U26720 (N_26720,N_26402,N_26385);
nand U26721 (N_26721,N_26339,N_26404);
nor U26722 (N_26722,N_26493,N_26272);
nand U26723 (N_26723,N_26369,N_26331);
nor U26724 (N_26724,N_26412,N_26341);
or U26725 (N_26725,N_26285,N_26310);
and U26726 (N_26726,N_26453,N_26307);
and U26727 (N_26727,N_26341,N_26466);
or U26728 (N_26728,N_26328,N_26414);
nand U26729 (N_26729,N_26289,N_26303);
nor U26730 (N_26730,N_26282,N_26281);
nor U26731 (N_26731,N_26283,N_26330);
nor U26732 (N_26732,N_26348,N_26450);
nor U26733 (N_26733,N_26317,N_26313);
xnor U26734 (N_26734,N_26382,N_26265);
or U26735 (N_26735,N_26318,N_26489);
nor U26736 (N_26736,N_26269,N_26433);
nor U26737 (N_26737,N_26497,N_26330);
xnor U26738 (N_26738,N_26268,N_26485);
and U26739 (N_26739,N_26277,N_26323);
nor U26740 (N_26740,N_26339,N_26436);
nor U26741 (N_26741,N_26358,N_26454);
nand U26742 (N_26742,N_26426,N_26266);
and U26743 (N_26743,N_26275,N_26425);
nand U26744 (N_26744,N_26430,N_26397);
xor U26745 (N_26745,N_26373,N_26267);
xor U26746 (N_26746,N_26318,N_26398);
or U26747 (N_26747,N_26267,N_26292);
nand U26748 (N_26748,N_26458,N_26296);
nand U26749 (N_26749,N_26306,N_26263);
and U26750 (N_26750,N_26731,N_26587);
nand U26751 (N_26751,N_26685,N_26526);
nand U26752 (N_26752,N_26675,N_26539);
nand U26753 (N_26753,N_26681,N_26656);
nor U26754 (N_26754,N_26729,N_26704);
or U26755 (N_26755,N_26670,N_26691);
or U26756 (N_26756,N_26650,N_26728);
nor U26757 (N_26757,N_26665,N_26624);
or U26758 (N_26758,N_26623,N_26727);
nand U26759 (N_26759,N_26601,N_26513);
and U26760 (N_26760,N_26648,N_26611);
or U26761 (N_26761,N_26600,N_26719);
xnor U26762 (N_26762,N_26563,N_26747);
and U26763 (N_26763,N_26643,N_26524);
xnor U26764 (N_26764,N_26636,N_26516);
xor U26765 (N_26765,N_26703,N_26680);
xor U26766 (N_26766,N_26720,N_26541);
nand U26767 (N_26767,N_26741,N_26535);
xnor U26768 (N_26768,N_26620,N_26594);
nand U26769 (N_26769,N_26617,N_26613);
xnor U26770 (N_26770,N_26560,N_26511);
nand U26771 (N_26771,N_26626,N_26637);
xor U26772 (N_26772,N_26736,N_26544);
xnor U26773 (N_26773,N_26548,N_26644);
or U26774 (N_26774,N_26553,N_26669);
nor U26775 (N_26775,N_26674,N_26602);
and U26776 (N_26776,N_26571,N_26507);
and U26777 (N_26777,N_26604,N_26706);
or U26778 (N_26778,N_26708,N_26559);
and U26779 (N_26779,N_26520,N_26584);
xnor U26780 (N_26780,N_26501,N_26543);
and U26781 (N_26781,N_26562,N_26567);
or U26782 (N_26782,N_26523,N_26663);
and U26783 (N_26783,N_26676,N_26672);
nor U26784 (N_26784,N_26597,N_26595);
nor U26785 (N_26785,N_26531,N_26661);
or U26786 (N_26786,N_26692,N_26723);
xor U26787 (N_26787,N_26694,N_26590);
nand U26788 (N_26788,N_26538,N_26622);
nor U26789 (N_26789,N_26546,N_26558);
nand U26790 (N_26790,N_26629,N_26709);
or U26791 (N_26791,N_26577,N_26688);
nor U26792 (N_26792,N_26696,N_26514);
xor U26793 (N_26793,N_26625,N_26651);
xor U26794 (N_26794,N_26545,N_26642);
and U26795 (N_26795,N_26542,N_26592);
nand U26796 (N_26796,N_26666,N_26618);
or U26797 (N_26797,N_26653,N_26698);
nand U26798 (N_26798,N_26660,N_26646);
or U26799 (N_26799,N_26671,N_26677);
or U26800 (N_26800,N_26735,N_26655);
or U26801 (N_26801,N_26580,N_26515);
xnor U26802 (N_26802,N_26599,N_26683);
xnor U26803 (N_26803,N_26621,N_26667);
nand U26804 (N_26804,N_26537,N_26554);
or U26805 (N_26805,N_26525,N_26569);
xor U26806 (N_26806,N_26589,N_26603);
or U26807 (N_26807,N_26512,N_26519);
nand U26808 (N_26808,N_26722,N_26639);
and U26809 (N_26809,N_26596,N_26712);
nor U26810 (N_26810,N_26641,N_26588);
xnor U26811 (N_26811,N_26557,N_26575);
and U26812 (N_26812,N_26744,N_26693);
nand U26813 (N_26813,N_26565,N_26573);
or U26814 (N_26814,N_26730,N_26609);
nand U26815 (N_26815,N_26534,N_26508);
and U26816 (N_26816,N_26732,N_26724);
xor U26817 (N_26817,N_26555,N_26605);
or U26818 (N_26818,N_26522,N_26654);
and U26819 (N_26819,N_26586,N_26549);
and U26820 (N_26820,N_26689,N_26570);
xnor U26821 (N_26821,N_26579,N_26610);
and U26822 (N_26822,N_26711,N_26566);
and U26823 (N_26823,N_26721,N_26733);
nand U26824 (N_26824,N_26614,N_26608);
or U26825 (N_26825,N_26628,N_26657);
and U26826 (N_26826,N_26506,N_26556);
or U26827 (N_26827,N_26568,N_26699);
nand U26828 (N_26828,N_26726,N_26503);
xor U26829 (N_26829,N_26690,N_26528);
or U26830 (N_26830,N_26630,N_26632);
xnor U26831 (N_26831,N_26529,N_26710);
nor U26832 (N_26832,N_26518,N_26734);
nand U26833 (N_26833,N_26684,N_26737);
xor U26834 (N_26834,N_26612,N_26662);
nor U26835 (N_26835,N_26504,N_26619);
xor U26836 (N_26836,N_26500,N_26550);
or U26837 (N_26837,N_26582,N_26743);
nand U26838 (N_26838,N_26510,N_26527);
and U26839 (N_26839,N_26673,N_26572);
nor U26840 (N_26840,N_26717,N_26581);
xor U26841 (N_26841,N_26532,N_26606);
and U26842 (N_26842,N_26713,N_26725);
and U26843 (N_26843,N_26749,N_26718);
or U26844 (N_26844,N_26705,N_26649);
and U26845 (N_26845,N_26634,N_26607);
xor U26846 (N_26846,N_26576,N_26578);
and U26847 (N_26847,N_26640,N_26533);
nor U26848 (N_26848,N_26745,N_26687);
and U26849 (N_26849,N_26695,N_26739);
xor U26850 (N_26850,N_26505,N_26682);
or U26851 (N_26851,N_26716,N_26652);
nor U26852 (N_26852,N_26638,N_26686);
xnor U26853 (N_26853,N_26658,N_26530);
nand U26854 (N_26854,N_26659,N_26521);
nand U26855 (N_26855,N_26707,N_26502);
or U26856 (N_26856,N_26748,N_26540);
and U26857 (N_26857,N_26678,N_26700);
or U26858 (N_26858,N_26664,N_26746);
nand U26859 (N_26859,N_26679,N_26645);
nand U26860 (N_26860,N_26536,N_26627);
and U26861 (N_26861,N_26702,N_26701);
xnor U26862 (N_26862,N_26574,N_26552);
and U26863 (N_26863,N_26635,N_26714);
and U26864 (N_26864,N_26593,N_26615);
and U26865 (N_26865,N_26697,N_26631);
and U26866 (N_26866,N_26561,N_26547);
and U26867 (N_26867,N_26509,N_26738);
xnor U26868 (N_26868,N_26517,N_26583);
xor U26869 (N_26869,N_26598,N_26591);
xnor U26870 (N_26870,N_26668,N_26616);
or U26871 (N_26871,N_26647,N_26585);
and U26872 (N_26872,N_26564,N_26551);
nand U26873 (N_26873,N_26633,N_26715);
or U26874 (N_26874,N_26742,N_26740);
nand U26875 (N_26875,N_26553,N_26676);
and U26876 (N_26876,N_26509,N_26584);
nand U26877 (N_26877,N_26580,N_26708);
nor U26878 (N_26878,N_26680,N_26627);
or U26879 (N_26879,N_26645,N_26657);
xnor U26880 (N_26880,N_26674,N_26661);
xor U26881 (N_26881,N_26553,N_26749);
nand U26882 (N_26882,N_26734,N_26733);
nor U26883 (N_26883,N_26517,N_26669);
and U26884 (N_26884,N_26715,N_26726);
nor U26885 (N_26885,N_26573,N_26650);
nor U26886 (N_26886,N_26523,N_26653);
and U26887 (N_26887,N_26628,N_26700);
or U26888 (N_26888,N_26624,N_26638);
nor U26889 (N_26889,N_26665,N_26592);
or U26890 (N_26890,N_26590,N_26595);
and U26891 (N_26891,N_26741,N_26577);
nor U26892 (N_26892,N_26557,N_26633);
or U26893 (N_26893,N_26698,N_26673);
xor U26894 (N_26894,N_26727,N_26680);
and U26895 (N_26895,N_26671,N_26503);
and U26896 (N_26896,N_26512,N_26611);
or U26897 (N_26897,N_26557,N_26586);
nor U26898 (N_26898,N_26581,N_26504);
nor U26899 (N_26899,N_26581,N_26574);
or U26900 (N_26900,N_26734,N_26594);
nand U26901 (N_26901,N_26661,N_26589);
or U26902 (N_26902,N_26618,N_26688);
nor U26903 (N_26903,N_26575,N_26668);
xnor U26904 (N_26904,N_26598,N_26652);
nor U26905 (N_26905,N_26727,N_26731);
xnor U26906 (N_26906,N_26643,N_26635);
or U26907 (N_26907,N_26668,N_26701);
or U26908 (N_26908,N_26687,N_26717);
xnor U26909 (N_26909,N_26669,N_26644);
or U26910 (N_26910,N_26504,N_26630);
xnor U26911 (N_26911,N_26574,N_26543);
nor U26912 (N_26912,N_26723,N_26679);
nor U26913 (N_26913,N_26689,N_26514);
xor U26914 (N_26914,N_26732,N_26733);
nor U26915 (N_26915,N_26647,N_26537);
nand U26916 (N_26916,N_26709,N_26634);
xor U26917 (N_26917,N_26746,N_26621);
nor U26918 (N_26918,N_26583,N_26703);
and U26919 (N_26919,N_26668,N_26663);
xor U26920 (N_26920,N_26647,N_26629);
nand U26921 (N_26921,N_26693,N_26737);
or U26922 (N_26922,N_26682,N_26526);
xnor U26923 (N_26923,N_26509,N_26525);
nor U26924 (N_26924,N_26558,N_26736);
nand U26925 (N_26925,N_26744,N_26629);
or U26926 (N_26926,N_26707,N_26686);
nor U26927 (N_26927,N_26516,N_26718);
nor U26928 (N_26928,N_26662,N_26505);
nor U26929 (N_26929,N_26711,N_26700);
or U26930 (N_26930,N_26675,N_26676);
nand U26931 (N_26931,N_26603,N_26534);
xnor U26932 (N_26932,N_26704,N_26747);
nand U26933 (N_26933,N_26522,N_26588);
nor U26934 (N_26934,N_26743,N_26520);
xor U26935 (N_26935,N_26618,N_26585);
nand U26936 (N_26936,N_26597,N_26704);
or U26937 (N_26937,N_26708,N_26515);
or U26938 (N_26938,N_26558,N_26557);
nand U26939 (N_26939,N_26702,N_26705);
nand U26940 (N_26940,N_26604,N_26717);
nor U26941 (N_26941,N_26737,N_26698);
and U26942 (N_26942,N_26579,N_26614);
nor U26943 (N_26943,N_26544,N_26551);
nand U26944 (N_26944,N_26712,N_26711);
nand U26945 (N_26945,N_26737,N_26645);
and U26946 (N_26946,N_26609,N_26592);
or U26947 (N_26947,N_26691,N_26663);
nor U26948 (N_26948,N_26720,N_26713);
nand U26949 (N_26949,N_26737,N_26720);
or U26950 (N_26950,N_26532,N_26609);
xor U26951 (N_26951,N_26656,N_26648);
xor U26952 (N_26952,N_26561,N_26731);
nand U26953 (N_26953,N_26636,N_26555);
xor U26954 (N_26954,N_26554,N_26685);
xnor U26955 (N_26955,N_26748,N_26727);
nand U26956 (N_26956,N_26607,N_26708);
nor U26957 (N_26957,N_26693,N_26697);
nand U26958 (N_26958,N_26637,N_26548);
nand U26959 (N_26959,N_26640,N_26525);
or U26960 (N_26960,N_26678,N_26685);
or U26961 (N_26961,N_26524,N_26599);
and U26962 (N_26962,N_26673,N_26544);
xnor U26963 (N_26963,N_26666,N_26507);
and U26964 (N_26964,N_26518,N_26659);
and U26965 (N_26965,N_26642,N_26553);
xor U26966 (N_26966,N_26518,N_26575);
or U26967 (N_26967,N_26550,N_26518);
xor U26968 (N_26968,N_26508,N_26686);
nor U26969 (N_26969,N_26734,N_26633);
xnor U26970 (N_26970,N_26523,N_26669);
xor U26971 (N_26971,N_26645,N_26732);
nor U26972 (N_26972,N_26680,N_26658);
xnor U26973 (N_26973,N_26683,N_26623);
xnor U26974 (N_26974,N_26589,N_26730);
and U26975 (N_26975,N_26596,N_26605);
and U26976 (N_26976,N_26628,N_26549);
and U26977 (N_26977,N_26573,N_26542);
or U26978 (N_26978,N_26667,N_26735);
or U26979 (N_26979,N_26654,N_26624);
nor U26980 (N_26980,N_26511,N_26566);
and U26981 (N_26981,N_26630,N_26654);
and U26982 (N_26982,N_26524,N_26507);
nand U26983 (N_26983,N_26723,N_26580);
or U26984 (N_26984,N_26583,N_26577);
nor U26985 (N_26985,N_26500,N_26540);
nor U26986 (N_26986,N_26713,N_26639);
nor U26987 (N_26987,N_26570,N_26571);
nand U26988 (N_26988,N_26665,N_26654);
nor U26989 (N_26989,N_26553,N_26601);
or U26990 (N_26990,N_26729,N_26535);
nor U26991 (N_26991,N_26501,N_26506);
nor U26992 (N_26992,N_26590,N_26558);
and U26993 (N_26993,N_26525,N_26576);
or U26994 (N_26994,N_26748,N_26643);
or U26995 (N_26995,N_26523,N_26704);
nand U26996 (N_26996,N_26516,N_26536);
nor U26997 (N_26997,N_26614,N_26545);
nor U26998 (N_26998,N_26572,N_26582);
xnor U26999 (N_26999,N_26539,N_26546);
nand U27000 (N_27000,N_26987,N_26802);
and U27001 (N_27001,N_26874,N_26875);
or U27002 (N_27002,N_26837,N_26867);
xnor U27003 (N_27003,N_26855,N_26955);
or U27004 (N_27004,N_26806,N_26765);
nand U27005 (N_27005,N_26941,N_26981);
and U27006 (N_27006,N_26872,N_26887);
or U27007 (N_27007,N_26804,N_26933);
and U27008 (N_27008,N_26970,N_26779);
and U27009 (N_27009,N_26992,N_26935);
nor U27010 (N_27010,N_26852,N_26936);
or U27011 (N_27011,N_26972,N_26807);
xnor U27012 (N_27012,N_26861,N_26750);
or U27013 (N_27013,N_26991,N_26897);
xor U27014 (N_27014,N_26790,N_26838);
or U27015 (N_27015,N_26982,N_26884);
or U27016 (N_27016,N_26752,N_26915);
or U27017 (N_27017,N_26766,N_26853);
or U27018 (N_27018,N_26929,N_26953);
or U27019 (N_27019,N_26883,N_26793);
nor U27020 (N_27020,N_26858,N_26985);
and U27021 (N_27021,N_26785,N_26866);
nand U27022 (N_27022,N_26820,N_26873);
xnor U27023 (N_27023,N_26946,N_26836);
and U27024 (N_27024,N_26845,N_26794);
or U27025 (N_27025,N_26879,N_26817);
and U27026 (N_27026,N_26797,N_26956);
nand U27027 (N_27027,N_26840,N_26942);
nor U27028 (N_27028,N_26975,N_26823);
nor U27029 (N_27029,N_26847,N_26977);
nand U27030 (N_27030,N_26891,N_26893);
or U27031 (N_27031,N_26792,N_26940);
nor U27032 (N_27032,N_26918,N_26895);
nand U27033 (N_27033,N_26880,N_26831);
or U27034 (N_27034,N_26833,N_26950);
nor U27035 (N_27035,N_26908,N_26938);
nand U27036 (N_27036,N_26778,N_26978);
and U27037 (N_27037,N_26799,N_26967);
and U27038 (N_27038,N_26890,N_26815);
xnor U27039 (N_27039,N_26851,N_26782);
or U27040 (N_27040,N_26767,N_26812);
or U27041 (N_27041,N_26926,N_26800);
or U27042 (N_27042,N_26772,N_26993);
nor U27043 (N_27043,N_26882,N_26819);
nor U27044 (N_27044,N_26943,N_26829);
and U27045 (N_27045,N_26796,N_26934);
nand U27046 (N_27046,N_26760,N_26947);
and U27047 (N_27047,N_26911,N_26763);
nand U27048 (N_27048,N_26900,N_26770);
nor U27049 (N_27049,N_26921,N_26924);
nor U27050 (N_27050,N_26920,N_26775);
and U27051 (N_27051,N_26835,N_26962);
nand U27052 (N_27052,N_26907,N_26986);
xnor U27053 (N_27053,N_26951,N_26830);
xor U27054 (N_27054,N_26885,N_26832);
nor U27055 (N_27055,N_26821,N_26808);
nand U27056 (N_27056,N_26974,N_26944);
xnor U27057 (N_27057,N_26754,N_26904);
and U27058 (N_27058,N_26932,N_26959);
nor U27059 (N_27059,N_26860,N_26759);
nand U27060 (N_27060,N_26958,N_26769);
nor U27061 (N_27061,N_26862,N_26989);
xnor U27062 (N_27062,N_26863,N_26898);
nand U27063 (N_27063,N_26952,N_26839);
or U27064 (N_27064,N_26798,N_26922);
or U27065 (N_27065,N_26780,N_26859);
nor U27066 (N_27066,N_26865,N_26979);
and U27067 (N_27067,N_26937,N_26996);
and U27068 (N_27068,N_26966,N_26886);
xor U27069 (N_27069,N_26927,N_26814);
xor U27070 (N_27070,N_26939,N_26773);
or U27071 (N_27071,N_26856,N_26925);
and U27072 (N_27072,N_26916,N_26849);
xor U27073 (N_27073,N_26784,N_26818);
xnor U27074 (N_27074,N_26848,N_26810);
or U27075 (N_27075,N_26795,N_26999);
and U27076 (N_27076,N_26764,N_26758);
and U27077 (N_27077,N_26843,N_26917);
and U27078 (N_27078,N_26816,N_26998);
or U27079 (N_27079,N_26954,N_26828);
and U27080 (N_27080,N_26803,N_26968);
or U27081 (N_27081,N_26903,N_26976);
nor U27082 (N_27082,N_26961,N_26930);
or U27083 (N_27083,N_26870,N_26871);
and U27084 (N_27084,N_26902,N_26827);
nor U27085 (N_27085,N_26912,N_26751);
or U27086 (N_27086,N_26825,N_26757);
nand U27087 (N_27087,N_26896,N_26761);
nor U27088 (N_27088,N_26864,N_26997);
or U27089 (N_27089,N_26777,N_26931);
nand U27090 (N_27090,N_26980,N_26877);
nor U27091 (N_27091,N_26841,N_26994);
nand U27092 (N_27092,N_26771,N_26973);
nor U27093 (N_27093,N_26949,N_26945);
nor U27094 (N_27094,N_26957,N_26755);
xor U27095 (N_27095,N_26846,N_26786);
nand U27096 (N_27096,N_26789,N_26850);
or U27097 (N_27097,N_26756,N_26905);
or U27098 (N_27098,N_26854,N_26801);
nand U27099 (N_27099,N_26842,N_26913);
nand U27100 (N_27100,N_26984,N_26844);
nand U27101 (N_27101,N_26813,N_26811);
nor U27102 (N_27102,N_26868,N_26888);
or U27103 (N_27103,N_26928,N_26781);
xnor U27104 (N_27104,N_26768,N_26788);
and U27105 (N_27105,N_26923,N_26990);
nand U27106 (N_27106,N_26889,N_26948);
and U27107 (N_27107,N_26901,N_26960);
nand U27108 (N_27108,N_26878,N_26965);
and U27109 (N_27109,N_26787,N_26909);
nor U27110 (N_27110,N_26894,N_26881);
nand U27111 (N_27111,N_26914,N_26892);
nor U27112 (N_27112,N_26876,N_26762);
or U27113 (N_27113,N_26963,N_26809);
xnor U27114 (N_27114,N_26869,N_26783);
xor U27115 (N_27115,N_26971,N_26919);
or U27116 (N_27116,N_26910,N_26964);
or U27117 (N_27117,N_26906,N_26834);
xnor U27118 (N_27118,N_26969,N_26899);
nand U27119 (N_27119,N_26826,N_26995);
nand U27120 (N_27120,N_26791,N_26857);
xnor U27121 (N_27121,N_26753,N_26805);
nand U27122 (N_27122,N_26822,N_26988);
or U27123 (N_27123,N_26824,N_26774);
xnor U27124 (N_27124,N_26776,N_26983);
xor U27125 (N_27125,N_26781,N_26765);
nor U27126 (N_27126,N_26822,N_26897);
nand U27127 (N_27127,N_26959,N_26832);
nand U27128 (N_27128,N_26938,N_26964);
xor U27129 (N_27129,N_26985,N_26774);
xnor U27130 (N_27130,N_26918,N_26766);
nand U27131 (N_27131,N_26940,N_26753);
xor U27132 (N_27132,N_26930,N_26819);
nor U27133 (N_27133,N_26794,N_26979);
and U27134 (N_27134,N_26953,N_26786);
nand U27135 (N_27135,N_26985,N_26845);
and U27136 (N_27136,N_26885,N_26976);
nor U27137 (N_27137,N_26965,N_26953);
xnor U27138 (N_27138,N_26805,N_26750);
xor U27139 (N_27139,N_26997,N_26973);
nor U27140 (N_27140,N_26804,N_26772);
or U27141 (N_27141,N_26927,N_26910);
nand U27142 (N_27142,N_26883,N_26986);
and U27143 (N_27143,N_26888,N_26789);
nor U27144 (N_27144,N_26812,N_26881);
nand U27145 (N_27145,N_26896,N_26777);
and U27146 (N_27146,N_26908,N_26779);
nor U27147 (N_27147,N_26799,N_26770);
nor U27148 (N_27148,N_26966,N_26787);
xnor U27149 (N_27149,N_26968,N_26892);
and U27150 (N_27150,N_26791,N_26967);
nand U27151 (N_27151,N_26859,N_26817);
xnor U27152 (N_27152,N_26962,N_26785);
nand U27153 (N_27153,N_26992,N_26973);
xnor U27154 (N_27154,N_26957,N_26969);
nor U27155 (N_27155,N_26930,N_26887);
and U27156 (N_27156,N_26960,N_26981);
or U27157 (N_27157,N_26868,N_26815);
nor U27158 (N_27158,N_26879,N_26904);
nand U27159 (N_27159,N_26832,N_26886);
xor U27160 (N_27160,N_26931,N_26844);
or U27161 (N_27161,N_26801,N_26932);
and U27162 (N_27162,N_26860,N_26875);
and U27163 (N_27163,N_26796,N_26958);
nand U27164 (N_27164,N_26967,N_26784);
xor U27165 (N_27165,N_26953,N_26827);
xnor U27166 (N_27166,N_26938,N_26927);
or U27167 (N_27167,N_26955,N_26896);
or U27168 (N_27168,N_26953,N_26810);
and U27169 (N_27169,N_26885,N_26929);
nand U27170 (N_27170,N_26921,N_26827);
nor U27171 (N_27171,N_26777,N_26861);
and U27172 (N_27172,N_26932,N_26879);
or U27173 (N_27173,N_26775,N_26818);
xor U27174 (N_27174,N_26978,N_26835);
or U27175 (N_27175,N_26789,N_26812);
xor U27176 (N_27176,N_26875,N_26978);
nor U27177 (N_27177,N_26933,N_26837);
xnor U27178 (N_27178,N_26863,N_26913);
nand U27179 (N_27179,N_26819,N_26949);
and U27180 (N_27180,N_26779,N_26759);
xnor U27181 (N_27181,N_26767,N_26985);
nor U27182 (N_27182,N_26961,N_26815);
and U27183 (N_27183,N_26790,N_26827);
xor U27184 (N_27184,N_26842,N_26755);
or U27185 (N_27185,N_26887,N_26904);
nand U27186 (N_27186,N_26801,N_26751);
or U27187 (N_27187,N_26904,N_26771);
xor U27188 (N_27188,N_26917,N_26750);
xor U27189 (N_27189,N_26755,N_26967);
and U27190 (N_27190,N_26875,N_26954);
nand U27191 (N_27191,N_26826,N_26864);
nand U27192 (N_27192,N_26941,N_26903);
xor U27193 (N_27193,N_26952,N_26911);
nand U27194 (N_27194,N_26770,N_26913);
nand U27195 (N_27195,N_26891,N_26795);
nor U27196 (N_27196,N_26900,N_26934);
or U27197 (N_27197,N_26958,N_26798);
and U27198 (N_27198,N_26836,N_26943);
nand U27199 (N_27199,N_26960,N_26839);
nor U27200 (N_27200,N_26797,N_26919);
nand U27201 (N_27201,N_26803,N_26872);
nor U27202 (N_27202,N_26798,N_26909);
xor U27203 (N_27203,N_26939,N_26893);
or U27204 (N_27204,N_26912,N_26940);
nor U27205 (N_27205,N_26990,N_26975);
nand U27206 (N_27206,N_26872,N_26864);
nand U27207 (N_27207,N_26928,N_26882);
and U27208 (N_27208,N_26781,N_26906);
nand U27209 (N_27209,N_26874,N_26825);
and U27210 (N_27210,N_26829,N_26991);
nor U27211 (N_27211,N_26940,N_26896);
and U27212 (N_27212,N_26984,N_26848);
nor U27213 (N_27213,N_26826,N_26883);
or U27214 (N_27214,N_26949,N_26794);
and U27215 (N_27215,N_26778,N_26793);
or U27216 (N_27216,N_26910,N_26785);
nor U27217 (N_27217,N_26813,N_26775);
nor U27218 (N_27218,N_26871,N_26848);
nor U27219 (N_27219,N_26837,N_26943);
nand U27220 (N_27220,N_26984,N_26770);
and U27221 (N_27221,N_26969,N_26820);
and U27222 (N_27222,N_26798,N_26817);
nor U27223 (N_27223,N_26779,N_26987);
or U27224 (N_27224,N_26798,N_26937);
and U27225 (N_27225,N_26966,N_26988);
xnor U27226 (N_27226,N_26998,N_26964);
xnor U27227 (N_27227,N_26845,N_26953);
and U27228 (N_27228,N_26968,N_26800);
xor U27229 (N_27229,N_26972,N_26956);
xor U27230 (N_27230,N_26874,N_26856);
and U27231 (N_27231,N_26941,N_26778);
xor U27232 (N_27232,N_26852,N_26752);
nor U27233 (N_27233,N_26756,N_26779);
xor U27234 (N_27234,N_26890,N_26950);
nand U27235 (N_27235,N_26944,N_26933);
xor U27236 (N_27236,N_26823,N_26948);
or U27237 (N_27237,N_26775,N_26842);
nor U27238 (N_27238,N_26913,N_26911);
xnor U27239 (N_27239,N_26957,N_26805);
xor U27240 (N_27240,N_26997,N_26984);
xnor U27241 (N_27241,N_26833,N_26870);
nand U27242 (N_27242,N_26839,N_26842);
nand U27243 (N_27243,N_26759,N_26840);
and U27244 (N_27244,N_26972,N_26801);
or U27245 (N_27245,N_26933,N_26970);
nor U27246 (N_27246,N_26994,N_26759);
nand U27247 (N_27247,N_26840,N_26900);
xor U27248 (N_27248,N_26828,N_26799);
and U27249 (N_27249,N_26776,N_26954);
or U27250 (N_27250,N_27213,N_27215);
and U27251 (N_27251,N_27010,N_27121);
xnor U27252 (N_27252,N_27074,N_27205);
nand U27253 (N_27253,N_27037,N_27005);
xor U27254 (N_27254,N_27170,N_27241);
or U27255 (N_27255,N_27052,N_27111);
xnor U27256 (N_27256,N_27050,N_27163);
or U27257 (N_27257,N_27176,N_27200);
and U27258 (N_27258,N_27027,N_27187);
xnor U27259 (N_27259,N_27230,N_27222);
and U27260 (N_27260,N_27044,N_27247);
and U27261 (N_27261,N_27218,N_27133);
or U27262 (N_27262,N_27207,N_27029);
or U27263 (N_27263,N_27234,N_27165);
nor U27264 (N_27264,N_27212,N_27235);
or U27265 (N_27265,N_27020,N_27203);
nand U27266 (N_27266,N_27167,N_27179);
xnor U27267 (N_27267,N_27184,N_27102);
and U27268 (N_27268,N_27047,N_27124);
nor U27269 (N_27269,N_27156,N_27064);
xor U27270 (N_27270,N_27002,N_27028);
xor U27271 (N_27271,N_27033,N_27195);
or U27272 (N_27272,N_27245,N_27058);
nor U27273 (N_27273,N_27243,N_27211);
xnor U27274 (N_27274,N_27060,N_27105);
nand U27275 (N_27275,N_27104,N_27189);
and U27276 (N_27276,N_27001,N_27079);
nor U27277 (N_27277,N_27128,N_27022);
xor U27278 (N_27278,N_27127,N_27084);
xnor U27279 (N_27279,N_27070,N_27065);
nand U27280 (N_27280,N_27067,N_27173);
and U27281 (N_27281,N_27095,N_27039);
xnor U27282 (N_27282,N_27016,N_27197);
nand U27283 (N_27283,N_27154,N_27149);
nand U27284 (N_27284,N_27181,N_27003);
or U27285 (N_27285,N_27096,N_27069);
nand U27286 (N_27286,N_27026,N_27140);
nor U27287 (N_27287,N_27150,N_27158);
nor U27288 (N_27288,N_27106,N_27209);
nor U27289 (N_27289,N_27094,N_27248);
nor U27290 (N_27290,N_27071,N_27024);
nor U27291 (N_27291,N_27025,N_27093);
nand U27292 (N_27292,N_27151,N_27119);
nand U27293 (N_27293,N_27108,N_27118);
nand U27294 (N_27294,N_27145,N_27092);
xor U27295 (N_27295,N_27110,N_27030);
nor U27296 (N_27296,N_27204,N_27055);
and U27297 (N_27297,N_27198,N_27068);
xor U27298 (N_27298,N_27229,N_27148);
and U27299 (N_27299,N_27099,N_27136);
nor U27300 (N_27300,N_27143,N_27240);
or U27301 (N_27301,N_27122,N_27153);
nand U27302 (N_27302,N_27043,N_27159);
nand U27303 (N_27303,N_27138,N_27238);
xor U27304 (N_27304,N_27009,N_27123);
nand U27305 (N_27305,N_27196,N_27112);
xor U27306 (N_27306,N_27171,N_27000);
nand U27307 (N_27307,N_27107,N_27019);
and U27308 (N_27308,N_27188,N_27226);
nand U27309 (N_27309,N_27134,N_27076);
xnor U27310 (N_27310,N_27178,N_27223);
and U27311 (N_27311,N_27175,N_27054);
nand U27312 (N_27312,N_27088,N_27168);
and U27313 (N_27313,N_27103,N_27081);
xor U27314 (N_27314,N_27157,N_27172);
nand U27315 (N_27315,N_27042,N_27014);
nand U27316 (N_27316,N_27186,N_27021);
nor U27317 (N_27317,N_27046,N_27051);
nor U27318 (N_27318,N_27169,N_27210);
or U27319 (N_27319,N_27221,N_27225);
or U27320 (N_27320,N_27155,N_27164);
nor U27321 (N_27321,N_27078,N_27237);
nand U27322 (N_27322,N_27032,N_27183);
nor U27323 (N_27323,N_27182,N_27089);
and U27324 (N_27324,N_27048,N_27090);
or U27325 (N_27325,N_27036,N_27227);
or U27326 (N_27326,N_27233,N_27246);
nand U27327 (N_27327,N_27201,N_27132);
and U27328 (N_27328,N_27049,N_27015);
and U27329 (N_27329,N_27012,N_27142);
or U27330 (N_27330,N_27082,N_27100);
or U27331 (N_27331,N_27144,N_27086);
nor U27332 (N_27332,N_27077,N_27031);
xor U27333 (N_27333,N_27113,N_27115);
or U27334 (N_27334,N_27053,N_27017);
nand U27335 (N_27335,N_27109,N_27066);
xnor U27336 (N_27336,N_27162,N_27097);
nand U27337 (N_27337,N_27177,N_27116);
or U27338 (N_27338,N_27041,N_27125);
and U27339 (N_27339,N_27057,N_27220);
or U27340 (N_27340,N_27152,N_27004);
nand U27341 (N_27341,N_27061,N_27190);
or U27342 (N_27342,N_27219,N_27034);
nand U27343 (N_27343,N_27007,N_27087);
nor U27344 (N_27344,N_27231,N_27141);
and U27345 (N_27345,N_27239,N_27192);
xor U27346 (N_27346,N_27193,N_27045);
nor U27347 (N_27347,N_27035,N_27101);
and U27348 (N_27348,N_27008,N_27147);
nand U27349 (N_27349,N_27202,N_27117);
or U27350 (N_27350,N_27146,N_27180);
nor U27351 (N_27351,N_27040,N_27139);
xnor U27352 (N_27352,N_27206,N_27135);
or U27353 (N_27353,N_27161,N_27080);
and U27354 (N_27354,N_27208,N_27006);
or U27355 (N_27355,N_27174,N_27137);
or U27356 (N_27356,N_27018,N_27214);
nand U27357 (N_27357,N_27085,N_27194);
nor U27358 (N_27358,N_27199,N_27236);
and U27359 (N_27359,N_27075,N_27228);
xor U27360 (N_27360,N_27062,N_27126);
or U27361 (N_27361,N_27191,N_27249);
and U27362 (N_27362,N_27120,N_27224);
nand U27363 (N_27363,N_27185,N_27242);
and U27364 (N_27364,N_27056,N_27072);
nor U27365 (N_27365,N_27023,N_27244);
and U27366 (N_27366,N_27073,N_27059);
nand U27367 (N_27367,N_27098,N_27129);
xnor U27368 (N_27368,N_27114,N_27091);
or U27369 (N_27369,N_27232,N_27160);
nor U27370 (N_27370,N_27216,N_27130);
and U27371 (N_27371,N_27131,N_27011);
xor U27372 (N_27372,N_27063,N_27013);
nand U27373 (N_27373,N_27166,N_27083);
xor U27374 (N_27374,N_27038,N_27217);
nand U27375 (N_27375,N_27175,N_27108);
and U27376 (N_27376,N_27158,N_27030);
and U27377 (N_27377,N_27106,N_27024);
xor U27378 (N_27378,N_27205,N_27043);
and U27379 (N_27379,N_27013,N_27026);
xor U27380 (N_27380,N_27044,N_27129);
nand U27381 (N_27381,N_27212,N_27050);
xor U27382 (N_27382,N_27026,N_27095);
or U27383 (N_27383,N_27126,N_27070);
nor U27384 (N_27384,N_27018,N_27243);
nand U27385 (N_27385,N_27049,N_27247);
xnor U27386 (N_27386,N_27183,N_27148);
nor U27387 (N_27387,N_27103,N_27187);
nand U27388 (N_27388,N_27177,N_27052);
nand U27389 (N_27389,N_27208,N_27102);
or U27390 (N_27390,N_27126,N_27051);
nor U27391 (N_27391,N_27203,N_27003);
and U27392 (N_27392,N_27136,N_27244);
and U27393 (N_27393,N_27023,N_27094);
or U27394 (N_27394,N_27110,N_27187);
or U27395 (N_27395,N_27072,N_27202);
nand U27396 (N_27396,N_27073,N_27164);
nand U27397 (N_27397,N_27067,N_27084);
or U27398 (N_27398,N_27170,N_27224);
or U27399 (N_27399,N_27130,N_27248);
nand U27400 (N_27400,N_27207,N_27174);
xnor U27401 (N_27401,N_27013,N_27048);
nand U27402 (N_27402,N_27233,N_27070);
or U27403 (N_27403,N_27163,N_27074);
nand U27404 (N_27404,N_27128,N_27236);
xor U27405 (N_27405,N_27244,N_27056);
and U27406 (N_27406,N_27106,N_27188);
nand U27407 (N_27407,N_27204,N_27196);
nand U27408 (N_27408,N_27058,N_27102);
or U27409 (N_27409,N_27160,N_27200);
xor U27410 (N_27410,N_27054,N_27079);
nand U27411 (N_27411,N_27232,N_27139);
or U27412 (N_27412,N_27029,N_27221);
or U27413 (N_27413,N_27197,N_27053);
nand U27414 (N_27414,N_27220,N_27200);
and U27415 (N_27415,N_27220,N_27052);
or U27416 (N_27416,N_27010,N_27162);
or U27417 (N_27417,N_27198,N_27246);
or U27418 (N_27418,N_27142,N_27049);
nand U27419 (N_27419,N_27165,N_27013);
nand U27420 (N_27420,N_27138,N_27053);
nor U27421 (N_27421,N_27169,N_27011);
and U27422 (N_27422,N_27056,N_27119);
xor U27423 (N_27423,N_27205,N_27044);
or U27424 (N_27424,N_27161,N_27122);
and U27425 (N_27425,N_27193,N_27164);
nand U27426 (N_27426,N_27112,N_27227);
nand U27427 (N_27427,N_27058,N_27108);
or U27428 (N_27428,N_27159,N_27197);
nor U27429 (N_27429,N_27208,N_27010);
and U27430 (N_27430,N_27214,N_27234);
nor U27431 (N_27431,N_27149,N_27110);
or U27432 (N_27432,N_27020,N_27041);
or U27433 (N_27433,N_27033,N_27129);
or U27434 (N_27434,N_27051,N_27013);
and U27435 (N_27435,N_27118,N_27067);
nand U27436 (N_27436,N_27195,N_27203);
nand U27437 (N_27437,N_27183,N_27143);
and U27438 (N_27438,N_27129,N_27039);
or U27439 (N_27439,N_27049,N_27025);
xor U27440 (N_27440,N_27110,N_27014);
xor U27441 (N_27441,N_27225,N_27187);
or U27442 (N_27442,N_27083,N_27192);
xnor U27443 (N_27443,N_27211,N_27183);
nor U27444 (N_27444,N_27123,N_27075);
nand U27445 (N_27445,N_27066,N_27242);
nor U27446 (N_27446,N_27121,N_27106);
or U27447 (N_27447,N_27099,N_27048);
xnor U27448 (N_27448,N_27155,N_27147);
and U27449 (N_27449,N_27011,N_27100);
or U27450 (N_27450,N_27241,N_27008);
and U27451 (N_27451,N_27183,N_27073);
xnor U27452 (N_27452,N_27144,N_27173);
and U27453 (N_27453,N_27083,N_27214);
or U27454 (N_27454,N_27020,N_27233);
nor U27455 (N_27455,N_27053,N_27179);
nor U27456 (N_27456,N_27173,N_27033);
xnor U27457 (N_27457,N_27021,N_27116);
xnor U27458 (N_27458,N_27119,N_27026);
xor U27459 (N_27459,N_27232,N_27036);
or U27460 (N_27460,N_27246,N_27053);
and U27461 (N_27461,N_27011,N_27108);
and U27462 (N_27462,N_27231,N_27120);
and U27463 (N_27463,N_27088,N_27217);
nor U27464 (N_27464,N_27175,N_27132);
nand U27465 (N_27465,N_27058,N_27127);
or U27466 (N_27466,N_27061,N_27215);
xnor U27467 (N_27467,N_27077,N_27167);
xnor U27468 (N_27468,N_27192,N_27215);
or U27469 (N_27469,N_27076,N_27196);
nand U27470 (N_27470,N_27011,N_27015);
or U27471 (N_27471,N_27105,N_27000);
and U27472 (N_27472,N_27166,N_27174);
and U27473 (N_27473,N_27171,N_27087);
nand U27474 (N_27474,N_27189,N_27158);
nand U27475 (N_27475,N_27132,N_27163);
nor U27476 (N_27476,N_27174,N_27222);
nand U27477 (N_27477,N_27008,N_27167);
nor U27478 (N_27478,N_27108,N_27007);
or U27479 (N_27479,N_27190,N_27029);
nor U27480 (N_27480,N_27013,N_27043);
and U27481 (N_27481,N_27068,N_27151);
nor U27482 (N_27482,N_27031,N_27148);
and U27483 (N_27483,N_27071,N_27096);
nand U27484 (N_27484,N_27135,N_27090);
nor U27485 (N_27485,N_27172,N_27116);
and U27486 (N_27486,N_27219,N_27132);
nor U27487 (N_27487,N_27024,N_27030);
nand U27488 (N_27488,N_27007,N_27122);
nor U27489 (N_27489,N_27023,N_27068);
nand U27490 (N_27490,N_27195,N_27041);
xor U27491 (N_27491,N_27076,N_27005);
or U27492 (N_27492,N_27243,N_27163);
xor U27493 (N_27493,N_27099,N_27107);
or U27494 (N_27494,N_27185,N_27208);
xor U27495 (N_27495,N_27013,N_27093);
and U27496 (N_27496,N_27244,N_27091);
and U27497 (N_27497,N_27078,N_27165);
or U27498 (N_27498,N_27225,N_27195);
nor U27499 (N_27499,N_27209,N_27003);
nand U27500 (N_27500,N_27455,N_27490);
nor U27501 (N_27501,N_27399,N_27457);
nor U27502 (N_27502,N_27341,N_27293);
nor U27503 (N_27503,N_27424,N_27398);
xnor U27504 (N_27504,N_27284,N_27252);
or U27505 (N_27505,N_27414,N_27335);
nor U27506 (N_27506,N_27297,N_27357);
and U27507 (N_27507,N_27267,N_27401);
or U27508 (N_27508,N_27380,N_27323);
nand U27509 (N_27509,N_27411,N_27409);
nor U27510 (N_27510,N_27333,N_27389);
or U27511 (N_27511,N_27382,N_27445);
xor U27512 (N_27512,N_27425,N_27459);
xnor U27513 (N_27513,N_27319,N_27487);
xnor U27514 (N_27514,N_27353,N_27478);
or U27515 (N_27515,N_27447,N_27273);
nand U27516 (N_27516,N_27493,N_27289);
nand U27517 (N_27517,N_27363,N_27268);
nand U27518 (N_27518,N_27430,N_27436);
or U27519 (N_27519,N_27471,N_27486);
nor U27520 (N_27520,N_27264,N_27317);
nand U27521 (N_27521,N_27279,N_27352);
and U27522 (N_27522,N_27361,N_27371);
nor U27523 (N_27523,N_27451,N_27497);
and U27524 (N_27524,N_27294,N_27467);
xor U27525 (N_27525,N_27378,N_27310);
nand U27526 (N_27526,N_27379,N_27390);
nand U27527 (N_27527,N_27412,N_27265);
nand U27528 (N_27528,N_27391,N_27368);
nand U27529 (N_27529,N_27427,N_27438);
nor U27530 (N_27530,N_27444,N_27448);
nand U27531 (N_27531,N_27304,N_27301);
and U27532 (N_27532,N_27359,N_27303);
xor U27533 (N_27533,N_27324,N_27278);
nand U27534 (N_27534,N_27462,N_27491);
xnor U27535 (N_27535,N_27376,N_27407);
xor U27536 (N_27536,N_27282,N_27292);
and U27537 (N_27537,N_27394,N_27452);
or U27538 (N_27538,N_27350,N_27277);
nand U27539 (N_27539,N_27388,N_27271);
and U27540 (N_27540,N_27318,N_27302);
nand U27541 (N_27541,N_27375,N_27251);
xnor U27542 (N_27542,N_27449,N_27494);
or U27543 (N_27543,N_27336,N_27463);
and U27544 (N_27544,N_27315,N_27370);
xor U27545 (N_27545,N_27320,N_27281);
or U27546 (N_27546,N_27299,N_27434);
or U27547 (N_27547,N_27440,N_27443);
xnor U27548 (N_27548,N_27280,N_27385);
or U27549 (N_27549,N_27495,N_27311);
and U27550 (N_27550,N_27396,N_27499);
and U27551 (N_27551,N_27377,N_27314);
nand U27552 (N_27552,N_27306,N_27477);
or U27553 (N_27553,N_27256,N_27488);
nor U27554 (N_27554,N_27461,N_27386);
nand U27555 (N_27555,N_27261,N_27288);
xor U27556 (N_27556,N_27383,N_27365);
nor U27557 (N_27557,N_27484,N_27250);
xor U27558 (N_27558,N_27332,N_27473);
and U27559 (N_27559,N_27367,N_27272);
or U27560 (N_27560,N_27309,N_27421);
nor U27561 (N_27561,N_27397,N_27330);
xor U27562 (N_27562,N_27441,N_27329);
nand U27563 (N_27563,N_27472,N_27348);
nand U27564 (N_27564,N_27358,N_27392);
or U27565 (N_27565,N_27346,N_27283);
xnor U27566 (N_27566,N_27454,N_27432);
and U27567 (N_27567,N_27415,N_27381);
and U27568 (N_27568,N_27465,N_27485);
or U27569 (N_27569,N_27402,N_27469);
and U27570 (N_27570,N_27433,N_27428);
or U27571 (N_27571,N_27468,N_27285);
or U27572 (N_27572,N_27286,N_27426);
xnor U27573 (N_27573,N_27287,N_27347);
nand U27574 (N_27574,N_27270,N_27258);
nor U27575 (N_27575,N_27260,N_27372);
xnor U27576 (N_27576,N_27429,N_27450);
nor U27577 (N_27577,N_27345,N_27431);
and U27578 (N_27578,N_27321,N_27254);
or U27579 (N_27579,N_27307,N_27422);
and U27580 (N_27580,N_27274,N_27437);
xnor U27581 (N_27581,N_27400,N_27366);
or U27582 (N_27582,N_27395,N_27325);
nand U27583 (N_27583,N_27470,N_27334);
xor U27584 (N_27584,N_27253,N_27364);
nand U27585 (N_27585,N_27263,N_27404);
and U27586 (N_27586,N_27354,N_27328);
or U27587 (N_27587,N_27356,N_27413);
or U27588 (N_27588,N_27344,N_27387);
nor U27589 (N_27589,N_27298,N_27410);
nand U27590 (N_27590,N_27393,N_27313);
or U27591 (N_27591,N_27498,N_27355);
and U27592 (N_27592,N_27349,N_27269);
xnor U27593 (N_27593,N_27339,N_27300);
and U27594 (N_27594,N_27464,N_27374);
and U27595 (N_27595,N_27316,N_27403);
nand U27596 (N_27596,N_27419,N_27420);
nand U27597 (N_27597,N_27305,N_27351);
nand U27598 (N_27598,N_27456,N_27369);
xor U27599 (N_27599,N_27373,N_27475);
nor U27600 (N_27600,N_27442,N_27466);
and U27601 (N_27601,N_27474,N_27257);
and U27602 (N_27602,N_27295,N_27262);
and U27603 (N_27603,N_27322,N_27331);
and U27604 (N_27604,N_27435,N_27259);
nor U27605 (N_27605,N_27418,N_27360);
nor U27606 (N_27606,N_27362,N_27308);
nand U27607 (N_27607,N_27312,N_27439);
or U27608 (N_27608,N_27275,N_27406);
nand U27609 (N_27609,N_27496,N_27276);
nor U27610 (N_27610,N_27492,N_27384);
or U27611 (N_27611,N_27476,N_27338);
or U27612 (N_27612,N_27483,N_27291);
nand U27613 (N_27613,N_27290,N_27340);
and U27614 (N_27614,N_27296,N_27423);
nor U27615 (N_27615,N_27326,N_27266);
and U27616 (N_27616,N_27343,N_27255);
and U27617 (N_27617,N_27327,N_27417);
or U27618 (N_27618,N_27460,N_27481);
nand U27619 (N_27619,N_27408,N_27337);
xor U27620 (N_27620,N_27342,N_27479);
xor U27621 (N_27621,N_27489,N_27446);
nor U27622 (N_27622,N_27405,N_27453);
nor U27623 (N_27623,N_27480,N_27458);
or U27624 (N_27624,N_27482,N_27416);
xnor U27625 (N_27625,N_27281,N_27353);
nor U27626 (N_27626,N_27475,N_27493);
or U27627 (N_27627,N_27464,N_27466);
xnor U27628 (N_27628,N_27320,N_27471);
nand U27629 (N_27629,N_27274,N_27486);
nand U27630 (N_27630,N_27363,N_27330);
or U27631 (N_27631,N_27264,N_27397);
and U27632 (N_27632,N_27356,N_27446);
and U27633 (N_27633,N_27389,N_27270);
xor U27634 (N_27634,N_27448,N_27291);
nor U27635 (N_27635,N_27460,N_27377);
nor U27636 (N_27636,N_27424,N_27336);
and U27637 (N_27637,N_27286,N_27407);
and U27638 (N_27638,N_27303,N_27485);
xnor U27639 (N_27639,N_27491,N_27254);
nor U27640 (N_27640,N_27436,N_27255);
or U27641 (N_27641,N_27411,N_27450);
and U27642 (N_27642,N_27283,N_27292);
and U27643 (N_27643,N_27269,N_27467);
and U27644 (N_27644,N_27259,N_27312);
xnor U27645 (N_27645,N_27256,N_27335);
xor U27646 (N_27646,N_27351,N_27309);
nand U27647 (N_27647,N_27436,N_27372);
and U27648 (N_27648,N_27436,N_27309);
nor U27649 (N_27649,N_27394,N_27326);
nand U27650 (N_27650,N_27298,N_27394);
nor U27651 (N_27651,N_27253,N_27403);
xor U27652 (N_27652,N_27340,N_27361);
nand U27653 (N_27653,N_27457,N_27416);
nor U27654 (N_27654,N_27284,N_27429);
or U27655 (N_27655,N_27490,N_27284);
or U27656 (N_27656,N_27351,N_27386);
and U27657 (N_27657,N_27355,N_27327);
xor U27658 (N_27658,N_27302,N_27269);
or U27659 (N_27659,N_27359,N_27356);
nand U27660 (N_27660,N_27423,N_27431);
nor U27661 (N_27661,N_27311,N_27450);
and U27662 (N_27662,N_27494,N_27362);
xnor U27663 (N_27663,N_27465,N_27284);
and U27664 (N_27664,N_27491,N_27350);
nand U27665 (N_27665,N_27443,N_27325);
or U27666 (N_27666,N_27373,N_27255);
nand U27667 (N_27667,N_27325,N_27474);
and U27668 (N_27668,N_27409,N_27381);
and U27669 (N_27669,N_27479,N_27475);
xor U27670 (N_27670,N_27378,N_27408);
nand U27671 (N_27671,N_27277,N_27293);
nor U27672 (N_27672,N_27322,N_27480);
nor U27673 (N_27673,N_27416,N_27341);
nand U27674 (N_27674,N_27489,N_27271);
nand U27675 (N_27675,N_27466,N_27432);
nand U27676 (N_27676,N_27358,N_27443);
xnor U27677 (N_27677,N_27390,N_27435);
xnor U27678 (N_27678,N_27359,N_27270);
and U27679 (N_27679,N_27410,N_27476);
nor U27680 (N_27680,N_27489,N_27332);
nand U27681 (N_27681,N_27457,N_27405);
nand U27682 (N_27682,N_27388,N_27384);
nand U27683 (N_27683,N_27478,N_27422);
nand U27684 (N_27684,N_27371,N_27319);
or U27685 (N_27685,N_27444,N_27309);
and U27686 (N_27686,N_27339,N_27325);
or U27687 (N_27687,N_27453,N_27332);
nand U27688 (N_27688,N_27367,N_27274);
nor U27689 (N_27689,N_27471,N_27255);
xnor U27690 (N_27690,N_27308,N_27446);
and U27691 (N_27691,N_27450,N_27457);
and U27692 (N_27692,N_27348,N_27441);
or U27693 (N_27693,N_27317,N_27362);
nand U27694 (N_27694,N_27421,N_27397);
or U27695 (N_27695,N_27267,N_27423);
and U27696 (N_27696,N_27422,N_27485);
or U27697 (N_27697,N_27446,N_27457);
xnor U27698 (N_27698,N_27383,N_27302);
xnor U27699 (N_27699,N_27304,N_27289);
and U27700 (N_27700,N_27428,N_27418);
and U27701 (N_27701,N_27318,N_27474);
nand U27702 (N_27702,N_27284,N_27479);
nor U27703 (N_27703,N_27304,N_27375);
nand U27704 (N_27704,N_27330,N_27408);
xnor U27705 (N_27705,N_27250,N_27497);
nand U27706 (N_27706,N_27325,N_27354);
or U27707 (N_27707,N_27327,N_27254);
nor U27708 (N_27708,N_27343,N_27274);
nor U27709 (N_27709,N_27428,N_27261);
nand U27710 (N_27710,N_27311,N_27444);
xor U27711 (N_27711,N_27477,N_27494);
nor U27712 (N_27712,N_27385,N_27452);
and U27713 (N_27713,N_27305,N_27332);
nand U27714 (N_27714,N_27314,N_27440);
or U27715 (N_27715,N_27265,N_27274);
nand U27716 (N_27716,N_27330,N_27474);
nor U27717 (N_27717,N_27338,N_27319);
xnor U27718 (N_27718,N_27259,N_27495);
xnor U27719 (N_27719,N_27417,N_27279);
or U27720 (N_27720,N_27369,N_27372);
xor U27721 (N_27721,N_27497,N_27382);
xor U27722 (N_27722,N_27433,N_27345);
xnor U27723 (N_27723,N_27401,N_27415);
nand U27724 (N_27724,N_27410,N_27297);
nor U27725 (N_27725,N_27419,N_27349);
nand U27726 (N_27726,N_27262,N_27420);
or U27727 (N_27727,N_27468,N_27341);
nand U27728 (N_27728,N_27410,N_27381);
and U27729 (N_27729,N_27402,N_27369);
and U27730 (N_27730,N_27349,N_27288);
nor U27731 (N_27731,N_27392,N_27409);
nand U27732 (N_27732,N_27334,N_27446);
xnor U27733 (N_27733,N_27257,N_27344);
or U27734 (N_27734,N_27385,N_27364);
nor U27735 (N_27735,N_27278,N_27339);
nor U27736 (N_27736,N_27298,N_27282);
nor U27737 (N_27737,N_27496,N_27354);
or U27738 (N_27738,N_27347,N_27377);
or U27739 (N_27739,N_27359,N_27304);
nand U27740 (N_27740,N_27459,N_27368);
xor U27741 (N_27741,N_27415,N_27272);
or U27742 (N_27742,N_27427,N_27439);
or U27743 (N_27743,N_27355,N_27475);
and U27744 (N_27744,N_27427,N_27311);
xor U27745 (N_27745,N_27282,N_27347);
nand U27746 (N_27746,N_27420,N_27410);
and U27747 (N_27747,N_27364,N_27304);
and U27748 (N_27748,N_27265,N_27307);
nor U27749 (N_27749,N_27274,N_27474);
or U27750 (N_27750,N_27604,N_27621);
nand U27751 (N_27751,N_27585,N_27592);
or U27752 (N_27752,N_27561,N_27703);
and U27753 (N_27753,N_27669,N_27686);
xor U27754 (N_27754,N_27603,N_27724);
and U27755 (N_27755,N_27682,N_27583);
nor U27756 (N_27756,N_27729,N_27627);
nor U27757 (N_27757,N_27602,N_27638);
or U27758 (N_27758,N_27720,N_27689);
nor U27759 (N_27759,N_27578,N_27513);
or U27760 (N_27760,N_27529,N_27524);
or U27761 (N_27761,N_27625,N_27635);
nand U27762 (N_27762,N_27525,N_27545);
or U27763 (N_27763,N_27519,N_27630);
and U27764 (N_27764,N_27553,N_27556);
nor U27765 (N_27765,N_27607,N_27721);
or U27766 (N_27766,N_27574,N_27537);
or U27767 (N_27767,N_27615,N_27712);
nor U27768 (N_27768,N_27503,N_27582);
and U27769 (N_27769,N_27555,N_27659);
and U27770 (N_27770,N_27610,N_27523);
nor U27771 (N_27771,N_27613,N_27534);
xnor U27772 (N_27772,N_27748,N_27741);
nor U27773 (N_27773,N_27586,N_27678);
and U27774 (N_27774,N_27532,N_27535);
xnor U27775 (N_27775,N_27598,N_27710);
or U27776 (N_27776,N_27623,N_27601);
or U27777 (N_27777,N_27747,N_27652);
and U27778 (N_27778,N_27629,N_27709);
nand U27779 (N_27779,N_27732,N_27714);
nand U27780 (N_27780,N_27707,N_27501);
or U27781 (N_27781,N_27569,N_27699);
and U27782 (N_27782,N_27677,N_27527);
nand U27783 (N_27783,N_27595,N_27565);
xor U27784 (N_27784,N_27536,N_27609);
and U27785 (N_27785,N_27684,N_27673);
xnor U27786 (N_27786,N_27606,N_27551);
and U27787 (N_27787,N_27576,N_27666);
xor U27788 (N_27788,N_27514,N_27680);
nand U27789 (N_27789,N_27575,N_27508);
nor U27790 (N_27790,N_27530,N_27691);
or U27791 (N_27791,N_27730,N_27579);
or U27792 (N_27792,N_27634,N_27648);
or U27793 (N_27793,N_27599,N_27591);
nand U27794 (N_27794,N_27675,N_27521);
and U27795 (N_27795,N_27653,N_27560);
or U27796 (N_27796,N_27676,N_27628);
nor U27797 (N_27797,N_27716,N_27708);
or U27798 (N_27798,N_27517,N_27564);
or U27799 (N_27799,N_27507,N_27559);
xnor U27800 (N_27800,N_27624,N_27643);
xnor U27801 (N_27801,N_27695,N_27512);
nand U27802 (N_27802,N_27528,N_27506);
xnor U27803 (N_27803,N_27644,N_27738);
or U27804 (N_27804,N_27726,N_27661);
or U27805 (N_27805,N_27672,N_27723);
nand U27806 (N_27806,N_27735,N_27660);
and U27807 (N_27807,N_27704,N_27746);
and U27808 (N_27808,N_27505,N_27745);
and U27809 (N_27809,N_27650,N_27500);
nand U27810 (N_27810,N_27719,N_27737);
nor U27811 (N_27811,N_27566,N_27674);
nand U27812 (N_27812,N_27740,N_27550);
xnor U27813 (N_27813,N_27544,N_27557);
nor U27814 (N_27814,N_27612,N_27611);
and U27815 (N_27815,N_27587,N_27725);
xor U27816 (N_27816,N_27522,N_27706);
nor U27817 (N_27817,N_27614,N_27731);
nand U27818 (N_27818,N_27580,N_27697);
nor U27819 (N_27819,N_27552,N_27665);
xnor U27820 (N_27820,N_27681,N_27640);
and U27821 (N_27821,N_27558,N_27713);
nand U27822 (N_27822,N_27663,N_27571);
nor U27823 (N_27823,N_27705,N_27533);
nor U27824 (N_27824,N_27633,N_27619);
or U27825 (N_27825,N_27562,N_27588);
xnor U27826 (N_27826,N_27538,N_27657);
or U27827 (N_27827,N_27670,N_27518);
xor U27828 (N_27828,N_27594,N_27700);
and U27829 (N_27829,N_27549,N_27547);
nand U27830 (N_27830,N_27687,N_27509);
nor U27831 (N_27831,N_27520,N_27671);
xor U27832 (N_27832,N_27698,N_27693);
xor U27833 (N_27833,N_27722,N_27502);
nand U27834 (N_27834,N_27543,N_27694);
and U27835 (N_27835,N_27637,N_27516);
nor U27836 (N_27836,N_27651,N_27742);
nor U27837 (N_27837,N_27642,N_27541);
xor U27838 (N_27838,N_27743,N_27540);
or U27839 (N_27839,N_27616,N_27542);
nor U27840 (N_27840,N_27656,N_27510);
nand U27841 (N_27841,N_27739,N_27734);
nor U27842 (N_27842,N_27662,N_27620);
nand U27843 (N_27843,N_27539,N_27622);
nor U27844 (N_27844,N_27526,N_27572);
nor U27845 (N_27845,N_27626,N_27573);
xnor U27846 (N_27846,N_27727,N_27679);
or U27847 (N_27847,N_27664,N_27702);
nand U27848 (N_27848,N_27744,N_27728);
xnor U27849 (N_27849,N_27584,N_27717);
nor U27850 (N_27850,N_27596,N_27617);
nand U27851 (N_27851,N_27568,N_27639);
nand U27852 (N_27852,N_27593,N_27641);
nand U27853 (N_27853,N_27692,N_27711);
nor U27854 (N_27854,N_27655,N_27589);
and U27855 (N_27855,N_27688,N_27701);
and U27856 (N_27856,N_27733,N_27600);
nor U27857 (N_27857,N_27597,N_27683);
nor U27858 (N_27858,N_27567,N_27647);
and U27859 (N_27859,N_27636,N_27715);
nand U27860 (N_27860,N_27581,N_27577);
nor U27861 (N_27861,N_27531,N_27654);
or U27862 (N_27862,N_27696,N_27548);
and U27863 (N_27863,N_27736,N_27618);
xor U27864 (N_27864,N_27632,N_27667);
nor U27865 (N_27865,N_27668,N_27690);
nand U27866 (N_27866,N_27554,N_27570);
nor U27867 (N_27867,N_27515,N_27718);
nand U27868 (N_27868,N_27631,N_27605);
nor U27869 (N_27869,N_27590,N_27563);
xnor U27870 (N_27870,N_27504,N_27645);
nand U27871 (N_27871,N_27649,N_27511);
nand U27872 (N_27872,N_27685,N_27749);
and U27873 (N_27873,N_27608,N_27646);
nor U27874 (N_27874,N_27658,N_27546);
xor U27875 (N_27875,N_27660,N_27644);
and U27876 (N_27876,N_27574,N_27566);
and U27877 (N_27877,N_27687,N_27636);
nand U27878 (N_27878,N_27684,N_27657);
or U27879 (N_27879,N_27710,N_27622);
xor U27880 (N_27880,N_27744,N_27517);
or U27881 (N_27881,N_27687,N_27557);
or U27882 (N_27882,N_27557,N_27595);
xnor U27883 (N_27883,N_27514,N_27633);
xnor U27884 (N_27884,N_27612,N_27702);
xnor U27885 (N_27885,N_27594,N_27502);
or U27886 (N_27886,N_27606,N_27731);
xnor U27887 (N_27887,N_27712,N_27503);
and U27888 (N_27888,N_27534,N_27566);
nor U27889 (N_27889,N_27674,N_27559);
xnor U27890 (N_27890,N_27612,N_27680);
or U27891 (N_27891,N_27644,N_27745);
and U27892 (N_27892,N_27676,N_27577);
xor U27893 (N_27893,N_27688,N_27656);
xor U27894 (N_27894,N_27646,N_27704);
or U27895 (N_27895,N_27540,N_27551);
nor U27896 (N_27896,N_27600,N_27628);
nor U27897 (N_27897,N_27729,N_27685);
nand U27898 (N_27898,N_27573,N_27675);
nand U27899 (N_27899,N_27589,N_27695);
and U27900 (N_27900,N_27611,N_27639);
nor U27901 (N_27901,N_27710,N_27587);
nor U27902 (N_27902,N_27665,N_27601);
or U27903 (N_27903,N_27730,N_27740);
xnor U27904 (N_27904,N_27730,N_27639);
nand U27905 (N_27905,N_27748,N_27705);
nand U27906 (N_27906,N_27701,N_27587);
xor U27907 (N_27907,N_27644,N_27564);
or U27908 (N_27908,N_27616,N_27647);
and U27909 (N_27909,N_27528,N_27726);
xnor U27910 (N_27910,N_27619,N_27500);
and U27911 (N_27911,N_27576,N_27577);
nand U27912 (N_27912,N_27526,N_27575);
nand U27913 (N_27913,N_27651,N_27623);
and U27914 (N_27914,N_27614,N_27651);
or U27915 (N_27915,N_27548,N_27646);
or U27916 (N_27916,N_27566,N_27668);
and U27917 (N_27917,N_27570,N_27628);
and U27918 (N_27918,N_27586,N_27684);
and U27919 (N_27919,N_27744,N_27543);
nand U27920 (N_27920,N_27652,N_27623);
nand U27921 (N_27921,N_27511,N_27527);
nor U27922 (N_27922,N_27645,N_27522);
nand U27923 (N_27923,N_27519,N_27672);
nand U27924 (N_27924,N_27530,N_27581);
nand U27925 (N_27925,N_27679,N_27677);
nand U27926 (N_27926,N_27688,N_27642);
nand U27927 (N_27927,N_27662,N_27532);
xnor U27928 (N_27928,N_27538,N_27521);
nand U27929 (N_27929,N_27617,N_27502);
and U27930 (N_27930,N_27513,N_27704);
or U27931 (N_27931,N_27537,N_27638);
nand U27932 (N_27932,N_27562,N_27749);
nor U27933 (N_27933,N_27670,N_27602);
nor U27934 (N_27934,N_27707,N_27708);
xnor U27935 (N_27935,N_27525,N_27696);
or U27936 (N_27936,N_27566,N_27723);
nor U27937 (N_27937,N_27676,N_27565);
and U27938 (N_27938,N_27700,N_27607);
and U27939 (N_27939,N_27660,N_27739);
nor U27940 (N_27940,N_27726,N_27654);
nor U27941 (N_27941,N_27700,N_27547);
nand U27942 (N_27942,N_27654,N_27547);
xnor U27943 (N_27943,N_27659,N_27736);
nand U27944 (N_27944,N_27604,N_27602);
and U27945 (N_27945,N_27540,N_27595);
nor U27946 (N_27946,N_27624,N_27533);
nand U27947 (N_27947,N_27508,N_27660);
nand U27948 (N_27948,N_27606,N_27737);
or U27949 (N_27949,N_27569,N_27539);
nand U27950 (N_27950,N_27638,N_27730);
nor U27951 (N_27951,N_27565,N_27682);
nor U27952 (N_27952,N_27709,N_27712);
or U27953 (N_27953,N_27551,N_27680);
and U27954 (N_27954,N_27527,N_27664);
nand U27955 (N_27955,N_27518,N_27668);
or U27956 (N_27956,N_27548,N_27607);
or U27957 (N_27957,N_27603,N_27612);
xnor U27958 (N_27958,N_27631,N_27667);
xor U27959 (N_27959,N_27685,N_27594);
or U27960 (N_27960,N_27743,N_27607);
xnor U27961 (N_27961,N_27591,N_27606);
nor U27962 (N_27962,N_27716,N_27513);
and U27963 (N_27963,N_27665,N_27658);
and U27964 (N_27964,N_27727,N_27644);
nand U27965 (N_27965,N_27565,N_27599);
nor U27966 (N_27966,N_27513,N_27549);
nor U27967 (N_27967,N_27622,N_27521);
nand U27968 (N_27968,N_27734,N_27539);
xor U27969 (N_27969,N_27502,N_27673);
nor U27970 (N_27970,N_27673,N_27524);
or U27971 (N_27971,N_27510,N_27720);
and U27972 (N_27972,N_27626,N_27514);
nand U27973 (N_27973,N_27733,N_27624);
xnor U27974 (N_27974,N_27508,N_27747);
nand U27975 (N_27975,N_27585,N_27536);
xnor U27976 (N_27976,N_27601,N_27535);
nor U27977 (N_27977,N_27625,N_27697);
or U27978 (N_27978,N_27575,N_27584);
nand U27979 (N_27979,N_27692,N_27736);
and U27980 (N_27980,N_27728,N_27709);
xnor U27981 (N_27981,N_27505,N_27533);
or U27982 (N_27982,N_27712,N_27501);
xor U27983 (N_27983,N_27650,N_27528);
xnor U27984 (N_27984,N_27635,N_27566);
and U27985 (N_27985,N_27660,N_27729);
nand U27986 (N_27986,N_27700,N_27562);
xor U27987 (N_27987,N_27653,N_27725);
nor U27988 (N_27988,N_27556,N_27712);
nand U27989 (N_27989,N_27640,N_27532);
nor U27990 (N_27990,N_27525,N_27702);
nor U27991 (N_27991,N_27646,N_27663);
and U27992 (N_27992,N_27570,N_27669);
nor U27993 (N_27993,N_27572,N_27662);
nand U27994 (N_27994,N_27549,N_27504);
or U27995 (N_27995,N_27610,N_27693);
and U27996 (N_27996,N_27593,N_27583);
xnor U27997 (N_27997,N_27573,N_27582);
nor U27998 (N_27998,N_27564,N_27727);
or U27999 (N_27999,N_27682,N_27536);
nor U28000 (N_28000,N_27931,N_27924);
and U28001 (N_28001,N_27886,N_27879);
xor U28002 (N_28002,N_27949,N_27938);
nor U28003 (N_28003,N_27772,N_27920);
xor U28004 (N_28004,N_27795,N_27853);
and U28005 (N_28005,N_27894,N_27956);
and U28006 (N_28006,N_27843,N_27836);
or U28007 (N_28007,N_27875,N_27874);
nand U28008 (N_28008,N_27842,N_27887);
and U28009 (N_28009,N_27932,N_27757);
or U28010 (N_28010,N_27979,N_27776);
or U28011 (N_28011,N_27935,N_27806);
or U28012 (N_28012,N_27813,N_27933);
xor U28013 (N_28013,N_27777,N_27865);
xor U28014 (N_28014,N_27943,N_27810);
nand U28015 (N_28015,N_27761,N_27906);
and U28016 (N_28016,N_27889,N_27974);
or U28017 (N_28017,N_27944,N_27860);
xnor U28018 (N_28018,N_27996,N_27845);
nor U28019 (N_28019,N_27922,N_27814);
nor U28020 (N_28020,N_27780,N_27873);
xor U28021 (N_28021,N_27970,N_27818);
or U28022 (N_28022,N_27800,N_27997);
nand U28023 (N_28023,N_27785,N_27982);
nand U28024 (N_28024,N_27815,N_27969);
nor U28025 (N_28025,N_27820,N_27902);
and U28026 (N_28026,N_27768,N_27835);
nand U28027 (N_28027,N_27939,N_27866);
and U28028 (N_28028,N_27999,N_27963);
and U28029 (N_28029,N_27833,N_27802);
nand U28030 (N_28030,N_27913,N_27799);
nand U28031 (N_28031,N_27900,N_27980);
xnor U28032 (N_28032,N_27872,N_27793);
xor U28033 (N_28033,N_27832,N_27888);
or U28034 (N_28034,N_27909,N_27891);
or U28035 (N_28035,N_27918,N_27990);
xor U28036 (N_28036,N_27767,N_27822);
xnor U28037 (N_28037,N_27798,N_27985);
xnor U28038 (N_28038,N_27998,N_27779);
nand U28039 (N_28039,N_27880,N_27801);
xor U28040 (N_28040,N_27870,N_27773);
xnor U28041 (N_28041,N_27829,N_27828);
or U28042 (N_28042,N_27796,N_27992);
or U28043 (N_28043,N_27946,N_27750);
and U28044 (N_28044,N_27912,N_27993);
nand U28045 (N_28045,N_27923,N_27821);
and U28046 (N_28046,N_27981,N_27781);
or U28047 (N_28047,N_27753,N_27751);
or U28048 (N_28048,N_27991,N_27859);
nand U28049 (N_28049,N_27819,N_27823);
xor U28050 (N_28050,N_27890,N_27864);
nor U28051 (N_28051,N_27910,N_27862);
xnor U28052 (N_28052,N_27968,N_27883);
nand U28053 (N_28053,N_27976,N_27987);
nand U28054 (N_28054,N_27812,N_27847);
xnor U28055 (N_28055,N_27966,N_27953);
or U28056 (N_28056,N_27774,N_27841);
nor U28057 (N_28057,N_27848,N_27811);
nor U28058 (N_28058,N_27789,N_27762);
xor U28059 (N_28059,N_27867,N_27892);
and U28060 (N_28060,N_27770,N_27878);
nand U28061 (N_28061,N_27784,N_27827);
xor U28062 (N_28062,N_27831,N_27852);
nor U28063 (N_28063,N_27755,N_27857);
xor U28064 (N_28064,N_27917,N_27834);
nor U28065 (N_28065,N_27901,N_27927);
and U28066 (N_28066,N_27948,N_27763);
xor U28067 (N_28067,N_27903,N_27915);
and U28068 (N_28068,N_27817,N_27805);
and U28069 (N_28069,N_27964,N_27790);
and U28070 (N_28070,N_27965,N_27850);
nand U28071 (N_28071,N_27881,N_27995);
xnor U28072 (N_28072,N_27911,N_27925);
nor U28073 (N_28073,N_27758,N_27752);
and U28074 (N_28074,N_27807,N_27869);
xnor U28075 (N_28075,N_27786,N_27914);
xor U28076 (N_28076,N_27861,N_27921);
or U28077 (N_28077,N_27849,N_27989);
and U28078 (N_28078,N_27816,N_27942);
nand U28079 (N_28079,N_27765,N_27788);
xor U28080 (N_28080,N_27830,N_27945);
or U28081 (N_28081,N_27895,N_27898);
and U28082 (N_28082,N_27754,N_27897);
xor U28083 (N_28083,N_27855,N_27856);
nand U28084 (N_28084,N_27958,N_27764);
nand U28085 (N_28085,N_27804,N_27908);
or U28086 (N_28086,N_27794,N_27947);
xor U28087 (N_28087,N_27882,N_27839);
and U28088 (N_28088,N_27775,N_27826);
xor U28089 (N_28089,N_27863,N_27904);
and U28090 (N_28090,N_27941,N_27936);
xor U28091 (N_28091,N_27871,N_27926);
or U28092 (N_28092,N_27957,N_27782);
or U28093 (N_28093,N_27824,N_27907);
xor U28094 (N_28094,N_27928,N_27846);
nor U28095 (N_28095,N_27838,N_27759);
xor U28096 (N_28096,N_27962,N_27986);
nand U28097 (N_28097,N_27988,N_27971);
and U28098 (N_28098,N_27837,N_27916);
or U28099 (N_28099,N_27978,N_27929);
nand U28100 (N_28100,N_27955,N_27950);
nand U28101 (N_28101,N_27972,N_27877);
and U28102 (N_28102,N_27803,N_27851);
nor U28103 (N_28103,N_27951,N_27919);
or U28104 (N_28104,N_27876,N_27899);
or U28105 (N_28105,N_27791,N_27896);
or U28106 (N_28106,N_27934,N_27960);
xnor U28107 (N_28107,N_27961,N_27959);
or U28108 (N_28108,N_27937,N_27769);
xor U28109 (N_28109,N_27973,N_27930);
and U28110 (N_28110,N_27858,N_27808);
and U28111 (N_28111,N_27797,N_27756);
and U28112 (N_28112,N_27885,N_27787);
or U28113 (N_28113,N_27854,N_27940);
nand U28114 (N_28114,N_27809,N_27844);
or U28115 (N_28115,N_27771,N_27954);
and U28116 (N_28116,N_27983,N_27792);
or U28117 (N_28117,N_27984,N_27952);
nor U28118 (N_28118,N_27893,N_27766);
nand U28119 (N_28119,N_27840,N_27868);
xor U28120 (N_28120,N_27967,N_27977);
and U28121 (N_28121,N_27778,N_27760);
nor U28122 (N_28122,N_27825,N_27905);
xor U28123 (N_28123,N_27884,N_27783);
nor U28124 (N_28124,N_27994,N_27975);
or U28125 (N_28125,N_27853,N_27974);
nor U28126 (N_28126,N_27887,N_27900);
and U28127 (N_28127,N_27928,N_27973);
or U28128 (N_28128,N_27771,N_27884);
nor U28129 (N_28129,N_27769,N_27975);
or U28130 (N_28130,N_27953,N_27772);
xnor U28131 (N_28131,N_27851,N_27912);
nor U28132 (N_28132,N_27757,N_27981);
nor U28133 (N_28133,N_27935,N_27843);
and U28134 (N_28134,N_27931,N_27821);
and U28135 (N_28135,N_27924,N_27870);
and U28136 (N_28136,N_27776,N_27845);
xor U28137 (N_28137,N_27990,N_27871);
nand U28138 (N_28138,N_27881,N_27994);
xnor U28139 (N_28139,N_27886,N_27806);
nor U28140 (N_28140,N_27780,N_27996);
or U28141 (N_28141,N_27854,N_27974);
and U28142 (N_28142,N_27983,N_27886);
nand U28143 (N_28143,N_27969,N_27911);
or U28144 (N_28144,N_27827,N_27794);
nand U28145 (N_28145,N_27909,N_27979);
and U28146 (N_28146,N_27956,N_27966);
or U28147 (N_28147,N_27887,N_27793);
nand U28148 (N_28148,N_27872,N_27797);
xnor U28149 (N_28149,N_27917,N_27905);
nand U28150 (N_28150,N_27896,N_27852);
and U28151 (N_28151,N_27785,N_27940);
nor U28152 (N_28152,N_27863,N_27857);
or U28153 (N_28153,N_27841,N_27940);
nor U28154 (N_28154,N_27791,N_27822);
xor U28155 (N_28155,N_27848,N_27915);
nor U28156 (N_28156,N_27833,N_27785);
or U28157 (N_28157,N_27812,N_27803);
nor U28158 (N_28158,N_27837,N_27801);
and U28159 (N_28159,N_27837,N_27759);
nand U28160 (N_28160,N_27963,N_27817);
nor U28161 (N_28161,N_27979,N_27931);
or U28162 (N_28162,N_27960,N_27814);
nand U28163 (N_28163,N_27917,N_27908);
or U28164 (N_28164,N_27889,N_27988);
or U28165 (N_28165,N_27838,N_27867);
and U28166 (N_28166,N_27970,N_27964);
xor U28167 (N_28167,N_27896,N_27799);
nor U28168 (N_28168,N_27956,N_27979);
and U28169 (N_28169,N_27884,N_27774);
nand U28170 (N_28170,N_27787,N_27785);
and U28171 (N_28171,N_27820,N_27872);
nor U28172 (N_28172,N_27969,N_27910);
nand U28173 (N_28173,N_27778,N_27939);
and U28174 (N_28174,N_27861,N_27862);
nor U28175 (N_28175,N_27885,N_27886);
xor U28176 (N_28176,N_27944,N_27847);
nand U28177 (N_28177,N_27957,N_27868);
and U28178 (N_28178,N_27787,N_27968);
xor U28179 (N_28179,N_27850,N_27849);
nand U28180 (N_28180,N_27809,N_27879);
nand U28181 (N_28181,N_27885,N_27868);
and U28182 (N_28182,N_27792,N_27978);
nand U28183 (N_28183,N_27866,N_27769);
and U28184 (N_28184,N_27973,N_27913);
nand U28185 (N_28185,N_27880,N_27815);
nor U28186 (N_28186,N_27917,N_27998);
and U28187 (N_28187,N_27944,N_27880);
nand U28188 (N_28188,N_27833,N_27767);
nand U28189 (N_28189,N_27811,N_27763);
or U28190 (N_28190,N_27932,N_27859);
and U28191 (N_28191,N_27832,N_27810);
nand U28192 (N_28192,N_27971,N_27908);
nor U28193 (N_28193,N_27813,N_27914);
nand U28194 (N_28194,N_27853,N_27811);
nand U28195 (N_28195,N_27778,N_27777);
nor U28196 (N_28196,N_27811,N_27884);
and U28197 (N_28197,N_27804,N_27981);
and U28198 (N_28198,N_27872,N_27831);
nand U28199 (N_28199,N_27829,N_27812);
or U28200 (N_28200,N_27787,N_27883);
and U28201 (N_28201,N_27777,N_27923);
or U28202 (N_28202,N_27804,N_27780);
nor U28203 (N_28203,N_27934,N_27834);
or U28204 (N_28204,N_27863,N_27921);
nor U28205 (N_28205,N_27770,N_27877);
or U28206 (N_28206,N_27861,N_27940);
xor U28207 (N_28207,N_27860,N_27968);
xor U28208 (N_28208,N_27953,N_27959);
and U28209 (N_28209,N_27895,N_27750);
or U28210 (N_28210,N_27782,N_27789);
and U28211 (N_28211,N_27808,N_27879);
nand U28212 (N_28212,N_27905,N_27860);
nand U28213 (N_28213,N_27901,N_27852);
nand U28214 (N_28214,N_27803,N_27976);
or U28215 (N_28215,N_27928,N_27867);
or U28216 (N_28216,N_27938,N_27816);
nand U28217 (N_28217,N_27984,N_27809);
nand U28218 (N_28218,N_27977,N_27832);
nand U28219 (N_28219,N_27989,N_27902);
or U28220 (N_28220,N_27941,N_27773);
xnor U28221 (N_28221,N_27840,N_27796);
nand U28222 (N_28222,N_27808,N_27884);
and U28223 (N_28223,N_27957,N_27788);
and U28224 (N_28224,N_27849,N_27892);
or U28225 (N_28225,N_27821,N_27901);
nor U28226 (N_28226,N_27814,N_27842);
xnor U28227 (N_28227,N_27835,N_27920);
nor U28228 (N_28228,N_27784,N_27929);
or U28229 (N_28229,N_27928,N_27915);
xnor U28230 (N_28230,N_27759,N_27921);
or U28231 (N_28231,N_27971,N_27812);
xor U28232 (N_28232,N_27929,N_27980);
nand U28233 (N_28233,N_27850,N_27877);
and U28234 (N_28234,N_27777,N_27996);
xnor U28235 (N_28235,N_27998,N_27988);
or U28236 (N_28236,N_27949,N_27855);
or U28237 (N_28237,N_27842,N_27974);
nor U28238 (N_28238,N_27802,N_27845);
nor U28239 (N_28239,N_27931,N_27879);
xnor U28240 (N_28240,N_27813,N_27765);
nand U28241 (N_28241,N_27886,N_27919);
nand U28242 (N_28242,N_27871,N_27806);
or U28243 (N_28243,N_27845,N_27816);
nand U28244 (N_28244,N_27830,N_27890);
xnor U28245 (N_28245,N_27920,N_27889);
or U28246 (N_28246,N_27810,N_27945);
and U28247 (N_28247,N_27790,N_27801);
xnor U28248 (N_28248,N_27776,N_27910);
or U28249 (N_28249,N_27817,N_27975);
nand U28250 (N_28250,N_28163,N_28136);
and U28251 (N_28251,N_28213,N_28248);
nand U28252 (N_28252,N_28041,N_28177);
nand U28253 (N_28253,N_28190,N_28245);
or U28254 (N_28254,N_28153,N_28031);
and U28255 (N_28255,N_28077,N_28064);
xnor U28256 (N_28256,N_28139,N_28197);
xor U28257 (N_28257,N_28036,N_28236);
and U28258 (N_28258,N_28210,N_28060);
or U28259 (N_28259,N_28212,N_28174);
or U28260 (N_28260,N_28241,N_28067);
nor U28261 (N_28261,N_28111,N_28232);
nor U28262 (N_28262,N_28164,N_28166);
and U28263 (N_28263,N_28070,N_28135);
xnor U28264 (N_28264,N_28222,N_28238);
xor U28265 (N_28265,N_28081,N_28157);
nand U28266 (N_28266,N_28184,N_28161);
and U28267 (N_28267,N_28209,N_28114);
nor U28268 (N_28268,N_28019,N_28040);
or U28269 (N_28269,N_28100,N_28092);
and U28270 (N_28270,N_28030,N_28078);
nor U28271 (N_28271,N_28089,N_28194);
and U28272 (N_28272,N_28009,N_28086);
or U28273 (N_28273,N_28096,N_28144);
xor U28274 (N_28274,N_28000,N_28120);
nor U28275 (N_28275,N_28215,N_28221);
and U28276 (N_28276,N_28061,N_28039);
nand U28277 (N_28277,N_28090,N_28156);
nor U28278 (N_28278,N_28199,N_28196);
or U28279 (N_28279,N_28165,N_28017);
nand U28280 (N_28280,N_28066,N_28071);
or U28281 (N_28281,N_28116,N_28047);
or U28282 (N_28282,N_28079,N_28002);
and U28283 (N_28283,N_28006,N_28219);
or U28284 (N_28284,N_28237,N_28140);
xor U28285 (N_28285,N_28158,N_28082);
xnor U28286 (N_28286,N_28138,N_28247);
xor U28287 (N_28287,N_28118,N_28123);
nor U28288 (N_28288,N_28110,N_28033);
and U28289 (N_28289,N_28011,N_28159);
nand U28290 (N_28290,N_28147,N_28054);
nand U28291 (N_28291,N_28091,N_28132);
xor U28292 (N_28292,N_28207,N_28173);
xor U28293 (N_28293,N_28239,N_28201);
and U28294 (N_28294,N_28169,N_28130);
or U28295 (N_28295,N_28024,N_28018);
and U28296 (N_28296,N_28073,N_28103);
nand U28297 (N_28297,N_28225,N_28171);
nor U28298 (N_28298,N_28023,N_28063);
nor U28299 (N_28299,N_28227,N_28125);
or U28300 (N_28300,N_28020,N_28108);
or U28301 (N_28301,N_28065,N_28029);
xor U28302 (N_28302,N_28145,N_28059);
nand U28303 (N_28303,N_28034,N_28128);
and U28304 (N_28304,N_28050,N_28137);
nor U28305 (N_28305,N_28014,N_28055);
or U28306 (N_28306,N_28240,N_28187);
and U28307 (N_28307,N_28220,N_28142);
or U28308 (N_28308,N_28022,N_28141);
xnor U28309 (N_28309,N_28188,N_28013);
or U28310 (N_28310,N_28037,N_28146);
and U28311 (N_28311,N_28233,N_28151);
or U28312 (N_28312,N_28057,N_28095);
xnor U28313 (N_28313,N_28226,N_28170);
nand U28314 (N_28314,N_28203,N_28074);
or U28315 (N_28315,N_28216,N_28122);
nor U28316 (N_28316,N_28104,N_28056);
xnor U28317 (N_28317,N_28053,N_28175);
nor U28318 (N_28318,N_28004,N_28242);
nand U28319 (N_28319,N_28133,N_28026);
nor U28320 (N_28320,N_28234,N_28032);
nor U28321 (N_28321,N_28246,N_28243);
nor U28322 (N_28322,N_28195,N_28223);
and U28323 (N_28323,N_28115,N_28178);
nor U28324 (N_28324,N_28102,N_28044);
nor U28325 (N_28325,N_28016,N_28205);
xor U28326 (N_28326,N_28183,N_28181);
xnor U28327 (N_28327,N_28154,N_28072);
nor U28328 (N_28328,N_28126,N_28167);
nand U28329 (N_28329,N_28107,N_28109);
nand U28330 (N_28330,N_28008,N_28075);
nor U28331 (N_28331,N_28021,N_28168);
nor U28332 (N_28332,N_28012,N_28204);
nand U28333 (N_28333,N_28069,N_28049);
nand U28334 (N_28334,N_28098,N_28080);
nor U28335 (N_28335,N_28228,N_28076);
and U28336 (N_28336,N_28121,N_28083);
nor U28337 (N_28337,N_28150,N_28099);
nor U28338 (N_28338,N_28087,N_28229);
nand U28339 (N_28339,N_28106,N_28206);
nor U28340 (N_28340,N_28200,N_28186);
and U28341 (N_28341,N_28027,N_28224);
or U28342 (N_28342,N_28045,N_28062);
and U28343 (N_28343,N_28113,N_28043);
nand U28344 (N_28344,N_28112,N_28172);
xor U28345 (N_28345,N_28231,N_28211);
xnor U28346 (N_28346,N_28155,N_28084);
and U28347 (N_28347,N_28025,N_28001);
nand U28348 (N_28348,N_28117,N_28218);
or U28349 (N_28349,N_28143,N_28244);
xor U28350 (N_28350,N_28176,N_28149);
or U28351 (N_28351,N_28189,N_28129);
nor U28352 (N_28352,N_28042,N_28068);
or U28353 (N_28353,N_28179,N_28124);
nor U28354 (N_28354,N_28005,N_28119);
nor U28355 (N_28355,N_28191,N_28185);
or U28356 (N_28356,N_28028,N_28198);
and U28357 (N_28357,N_28131,N_28003);
nor U28358 (N_28358,N_28134,N_28127);
and U28359 (N_28359,N_28180,N_28249);
and U28360 (N_28360,N_28007,N_28097);
or U28361 (N_28361,N_28182,N_28093);
nor U28362 (N_28362,N_28052,N_28235);
xor U28363 (N_28363,N_28105,N_28152);
or U28364 (N_28364,N_28214,N_28217);
xor U28365 (N_28365,N_28160,N_28010);
nand U28366 (N_28366,N_28202,N_28046);
xor U28367 (N_28367,N_28085,N_28058);
and U28368 (N_28368,N_28048,N_28094);
or U28369 (N_28369,N_28038,N_28051);
or U28370 (N_28370,N_28015,N_28148);
nand U28371 (N_28371,N_28208,N_28101);
xor U28372 (N_28372,N_28192,N_28035);
nor U28373 (N_28373,N_28162,N_28088);
nand U28374 (N_28374,N_28193,N_28230);
and U28375 (N_28375,N_28005,N_28186);
xnor U28376 (N_28376,N_28051,N_28184);
xnor U28377 (N_28377,N_28164,N_28070);
nor U28378 (N_28378,N_28207,N_28131);
or U28379 (N_28379,N_28216,N_28024);
xnor U28380 (N_28380,N_28119,N_28154);
nand U28381 (N_28381,N_28221,N_28152);
or U28382 (N_28382,N_28203,N_28192);
nand U28383 (N_28383,N_28190,N_28176);
or U28384 (N_28384,N_28159,N_28179);
and U28385 (N_28385,N_28056,N_28153);
or U28386 (N_28386,N_28179,N_28170);
nand U28387 (N_28387,N_28186,N_28020);
xnor U28388 (N_28388,N_28193,N_28208);
nand U28389 (N_28389,N_28235,N_28171);
and U28390 (N_28390,N_28080,N_28111);
xor U28391 (N_28391,N_28247,N_28044);
nand U28392 (N_28392,N_28159,N_28052);
or U28393 (N_28393,N_28101,N_28224);
or U28394 (N_28394,N_28142,N_28067);
nor U28395 (N_28395,N_28031,N_28072);
xor U28396 (N_28396,N_28142,N_28198);
xor U28397 (N_28397,N_28099,N_28229);
and U28398 (N_28398,N_28238,N_28105);
or U28399 (N_28399,N_28160,N_28167);
or U28400 (N_28400,N_28207,N_28227);
xnor U28401 (N_28401,N_28203,N_28029);
nor U28402 (N_28402,N_28159,N_28028);
nand U28403 (N_28403,N_28184,N_28202);
nand U28404 (N_28404,N_28103,N_28056);
or U28405 (N_28405,N_28200,N_28204);
nand U28406 (N_28406,N_28086,N_28084);
or U28407 (N_28407,N_28012,N_28207);
or U28408 (N_28408,N_28181,N_28240);
or U28409 (N_28409,N_28043,N_28154);
and U28410 (N_28410,N_28122,N_28157);
and U28411 (N_28411,N_28048,N_28078);
xnor U28412 (N_28412,N_28149,N_28096);
nor U28413 (N_28413,N_28142,N_28090);
nor U28414 (N_28414,N_28069,N_28244);
xor U28415 (N_28415,N_28126,N_28004);
xor U28416 (N_28416,N_28105,N_28022);
xnor U28417 (N_28417,N_28106,N_28016);
or U28418 (N_28418,N_28044,N_28188);
and U28419 (N_28419,N_28196,N_28243);
xnor U28420 (N_28420,N_28035,N_28082);
nor U28421 (N_28421,N_28124,N_28040);
and U28422 (N_28422,N_28162,N_28005);
nand U28423 (N_28423,N_28166,N_28203);
xor U28424 (N_28424,N_28188,N_28233);
nor U28425 (N_28425,N_28036,N_28138);
xnor U28426 (N_28426,N_28123,N_28225);
or U28427 (N_28427,N_28024,N_28164);
xor U28428 (N_28428,N_28076,N_28095);
xor U28429 (N_28429,N_28171,N_28249);
nand U28430 (N_28430,N_28130,N_28099);
or U28431 (N_28431,N_28024,N_28097);
nand U28432 (N_28432,N_28019,N_28199);
and U28433 (N_28433,N_28167,N_28024);
nor U28434 (N_28434,N_28065,N_28226);
and U28435 (N_28435,N_28222,N_28247);
nand U28436 (N_28436,N_28164,N_28169);
or U28437 (N_28437,N_28186,N_28233);
nand U28438 (N_28438,N_28226,N_28207);
xnor U28439 (N_28439,N_28129,N_28034);
nand U28440 (N_28440,N_28178,N_28150);
xor U28441 (N_28441,N_28193,N_28083);
or U28442 (N_28442,N_28064,N_28040);
nor U28443 (N_28443,N_28202,N_28142);
or U28444 (N_28444,N_28098,N_28226);
or U28445 (N_28445,N_28074,N_28027);
nand U28446 (N_28446,N_28146,N_28059);
nand U28447 (N_28447,N_28182,N_28181);
nand U28448 (N_28448,N_28027,N_28076);
xor U28449 (N_28449,N_28091,N_28184);
and U28450 (N_28450,N_28194,N_28161);
nand U28451 (N_28451,N_28178,N_28041);
and U28452 (N_28452,N_28239,N_28161);
xor U28453 (N_28453,N_28072,N_28020);
nor U28454 (N_28454,N_28158,N_28021);
nor U28455 (N_28455,N_28050,N_28041);
xor U28456 (N_28456,N_28013,N_28097);
nand U28457 (N_28457,N_28044,N_28189);
xnor U28458 (N_28458,N_28234,N_28002);
or U28459 (N_28459,N_28191,N_28047);
nor U28460 (N_28460,N_28162,N_28227);
nand U28461 (N_28461,N_28234,N_28091);
nor U28462 (N_28462,N_28194,N_28232);
nand U28463 (N_28463,N_28095,N_28039);
nand U28464 (N_28464,N_28010,N_28051);
or U28465 (N_28465,N_28006,N_28192);
or U28466 (N_28466,N_28203,N_28048);
and U28467 (N_28467,N_28069,N_28193);
or U28468 (N_28468,N_28132,N_28033);
and U28469 (N_28469,N_28018,N_28046);
or U28470 (N_28470,N_28215,N_28077);
and U28471 (N_28471,N_28017,N_28223);
nor U28472 (N_28472,N_28240,N_28232);
nand U28473 (N_28473,N_28023,N_28124);
and U28474 (N_28474,N_28038,N_28021);
and U28475 (N_28475,N_28206,N_28119);
or U28476 (N_28476,N_28193,N_28073);
or U28477 (N_28477,N_28061,N_28198);
nand U28478 (N_28478,N_28132,N_28061);
xnor U28479 (N_28479,N_28106,N_28130);
nor U28480 (N_28480,N_28089,N_28216);
and U28481 (N_28481,N_28011,N_28140);
nor U28482 (N_28482,N_28123,N_28000);
nand U28483 (N_28483,N_28107,N_28182);
xor U28484 (N_28484,N_28019,N_28062);
nand U28485 (N_28485,N_28210,N_28124);
xnor U28486 (N_28486,N_28238,N_28042);
xnor U28487 (N_28487,N_28121,N_28190);
and U28488 (N_28488,N_28033,N_28071);
nor U28489 (N_28489,N_28231,N_28089);
nand U28490 (N_28490,N_28086,N_28157);
and U28491 (N_28491,N_28047,N_28161);
nor U28492 (N_28492,N_28025,N_28160);
or U28493 (N_28493,N_28109,N_28189);
nand U28494 (N_28494,N_28174,N_28198);
or U28495 (N_28495,N_28120,N_28042);
nor U28496 (N_28496,N_28011,N_28150);
or U28497 (N_28497,N_28105,N_28227);
xor U28498 (N_28498,N_28135,N_28011);
nor U28499 (N_28499,N_28140,N_28002);
nor U28500 (N_28500,N_28443,N_28267);
nor U28501 (N_28501,N_28365,N_28408);
nand U28502 (N_28502,N_28265,N_28341);
or U28503 (N_28503,N_28407,N_28380);
or U28504 (N_28504,N_28378,N_28471);
and U28505 (N_28505,N_28421,N_28426);
or U28506 (N_28506,N_28262,N_28384);
nor U28507 (N_28507,N_28453,N_28311);
or U28508 (N_28508,N_28442,N_28395);
nand U28509 (N_28509,N_28431,N_28418);
and U28510 (N_28510,N_28400,N_28279);
nor U28511 (N_28511,N_28413,N_28417);
nor U28512 (N_28512,N_28349,N_28329);
nor U28513 (N_28513,N_28363,N_28324);
nand U28514 (N_28514,N_28332,N_28405);
xor U28515 (N_28515,N_28483,N_28458);
and U28516 (N_28516,N_28444,N_28312);
nor U28517 (N_28517,N_28411,N_28399);
nand U28518 (N_28518,N_28290,N_28364);
nand U28519 (N_28519,N_28331,N_28354);
and U28520 (N_28520,N_28278,N_28455);
and U28521 (N_28521,N_28414,N_28465);
or U28522 (N_28522,N_28422,N_28284);
or U28523 (N_28523,N_28445,N_28448);
nor U28524 (N_28524,N_28327,N_28469);
or U28525 (N_28525,N_28498,N_28462);
or U28526 (N_28526,N_28306,N_28253);
xor U28527 (N_28527,N_28438,N_28492);
nor U28528 (N_28528,N_28352,N_28261);
nand U28529 (N_28529,N_28360,N_28270);
nor U28530 (N_28530,N_28314,N_28266);
nand U28531 (N_28531,N_28372,N_28355);
or U28532 (N_28532,N_28348,N_28477);
nor U28533 (N_28533,N_28404,N_28346);
or U28534 (N_28534,N_28330,N_28376);
nor U28535 (N_28535,N_28291,N_28467);
nor U28536 (N_28536,N_28283,N_28379);
xnor U28537 (N_28537,N_28373,N_28474);
and U28538 (N_28538,N_28416,N_28464);
xnor U28539 (N_28539,N_28287,N_28293);
nor U28540 (N_28540,N_28487,N_28370);
nand U28541 (N_28541,N_28440,N_28401);
nand U28542 (N_28542,N_28361,N_28495);
xor U28543 (N_28543,N_28398,N_28402);
or U28544 (N_28544,N_28430,N_28494);
nor U28545 (N_28545,N_28297,N_28308);
nor U28546 (N_28546,N_28396,N_28454);
or U28547 (N_28547,N_28470,N_28480);
nand U28548 (N_28548,N_28432,N_28436);
xor U28549 (N_28549,N_28473,N_28461);
or U28550 (N_28550,N_28298,N_28450);
and U28551 (N_28551,N_28320,N_28342);
or U28552 (N_28552,N_28449,N_28447);
nor U28553 (N_28553,N_28446,N_28264);
or U28554 (N_28554,N_28280,N_28328);
nor U28555 (N_28555,N_28345,N_28351);
nand U28556 (N_28556,N_28389,N_28456);
nor U28557 (N_28557,N_28285,N_28313);
xor U28558 (N_28558,N_28323,N_28488);
nand U28559 (N_28559,N_28325,N_28309);
or U28560 (N_28560,N_28282,N_28250);
nand U28561 (N_28561,N_28254,N_28321);
or U28562 (N_28562,N_28335,N_28347);
nand U28563 (N_28563,N_28392,N_28307);
nand U28564 (N_28564,N_28319,N_28434);
xnor U28565 (N_28565,N_28344,N_28472);
nand U28566 (N_28566,N_28326,N_28459);
nand U28567 (N_28567,N_28423,N_28394);
nand U28568 (N_28568,N_28486,N_28439);
xnor U28569 (N_28569,N_28252,N_28371);
nor U28570 (N_28570,N_28268,N_28356);
nor U28571 (N_28571,N_28369,N_28419);
xor U28572 (N_28572,N_28499,N_28479);
xor U28573 (N_28573,N_28271,N_28412);
nor U28574 (N_28574,N_28476,N_28468);
xnor U28575 (N_28575,N_28385,N_28334);
or U28576 (N_28576,N_28391,N_28263);
nor U28577 (N_28577,N_28481,N_28463);
nor U28578 (N_28578,N_28318,N_28466);
xnor U28579 (N_28579,N_28343,N_28420);
and U28580 (N_28580,N_28485,N_28299);
nor U28581 (N_28581,N_28409,N_28286);
xor U28582 (N_28582,N_28415,N_28359);
and U28583 (N_28583,N_28457,N_28353);
or U28584 (N_28584,N_28338,N_28386);
xor U28585 (N_28585,N_28269,N_28295);
xnor U28586 (N_28586,N_28382,N_28281);
nand U28587 (N_28587,N_28301,N_28489);
xnor U28588 (N_28588,N_28437,N_28251);
and U28589 (N_28589,N_28393,N_28336);
and U28590 (N_28590,N_28397,N_28429);
xor U28591 (N_28591,N_28358,N_28460);
nand U28592 (N_28592,N_28497,N_28340);
or U28593 (N_28593,N_28478,N_28406);
xnor U28594 (N_28594,N_28337,N_28303);
and U28595 (N_28595,N_28357,N_28333);
or U28596 (N_28596,N_28275,N_28367);
nor U28597 (N_28597,N_28491,N_28375);
nor U28598 (N_28598,N_28339,N_28294);
nand U28599 (N_28599,N_28315,N_28259);
and U28600 (N_28600,N_28322,N_28289);
and U28601 (N_28601,N_28484,N_28272);
or U28602 (N_28602,N_28255,N_28362);
nand U28603 (N_28603,N_28276,N_28435);
nor U28604 (N_28604,N_28258,N_28377);
and U28605 (N_28605,N_28451,N_28425);
xnor U28606 (N_28606,N_28427,N_28433);
xnor U28607 (N_28607,N_28296,N_28305);
xnor U28608 (N_28608,N_28424,N_28496);
or U28609 (N_28609,N_28388,N_28441);
nand U28610 (N_28610,N_28475,N_28260);
and U28611 (N_28611,N_28310,N_28410);
nor U28612 (N_28612,N_28381,N_28273);
nand U28613 (N_28613,N_28292,N_28302);
and U28614 (N_28614,N_28493,N_28383);
xnor U28615 (N_28615,N_28403,N_28428);
nand U28616 (N_28616,N_28300,N_28387);
and U28617 (N_28617,N_28374,N_28366);
or U28618 (N_28618,N_28288,N_28482);
xnor U28619 (N_28619,N_28274,N_28390);
or U28620 (N_28620,N_28490,N_28350);
or U28621 (N_28621,N_28368,N_28316);
and U28622 (N_28622,N_28257,N_28256);
nand U28623 (N_28623,N_28452,N_28317);
nand U28624 (N_28624,N_28304,N_28277);
and U28625 (N_28625,N_28318,N_28397);
and U28626 (N_28626,N_28358,N_28262);
and U28627 (N_28627,N_28433,N_28407);
xnor U28628 (N_28628,N_28292,N_28464);
or U28629 (N_28629,N_28376,N_28473);
or U28630 (N_28630,N_28410,N_28390);
nand U28631 (N_28631,N_28352,N_28334);
nor U28632 (N_28632,N_28411,N_28371);
nor U28633 (N_28633,N_28332,N_28255);
and U28634 (N_28634,N_28488,N_28312);
and U28635 (N_28635,N_28280,N_28299);
or U28636 (N_28636,N_28310,N_28392);
nand U28637 (N_28637,N_28383,N_28324);
or U28638 (N_28638,N_28290,N_28388);
nand U28639 (N_28639,N_28307,N_28268);
and U28640 (N_28640,N_28483,N_28251);
xnor U28641 (N_28641,N_28252,N_28477);
nor U28642 (N_28642,N_28387,N_28301);
or U28643 (N_28643,N_28477,N_28461);
nand U28644 (N_28644,N_28343,N_28259);
xnor U28645 (N_28645,N_28338,N_28347);
and U28646 (N_28646,N_28255,N_28318);
xor U28647 (N_28647,N_28326,N_28458);
or U28648 (N_28648,N_28361,N_28295);
xor U28649 (N_28649,N_28494,N_28303);
or U28650 (N_28650,N_28371,N_28299);
and U28651 (N_28651,N_28439,N_28491);
and U28652 (N_28652,N_28298,N_28387);
nand U28653 (N_28653,N_28378,N_28379);
and U28654 (N_28654,N_28425,N_28386);
xor U28655 (N_28655,N_28399,N_28388);
and U28656 (N_28656,N_28467,N_28255);
and U28657 (N_28657,N_28365,N_28410);
xnor U28658 (N_28658,N_28401,N_28329);
or U28659 (N_28659,N_28355,N_28486);
nor U28660 (N_28660,N_28309,N_28455);
nand U28661 (N_28661,N_28426,N_28417);
and U28662 (N_28662,N_28298,N_28287);
or U28663 (N_28663,N_28319,N_28339);
or U28664 (N_28664,N_28383,N_28266);
nand U28665 (N_28665,N_28347,N_28292);
nand U28666 (N_28666,N_28292,N_28356);
nand U28667 (N_28667,N_28492,N_28386);
nor U28668 (N_28668,N_28397,N_28320);
nor U28669 (N_28669,N_28474,N_28407);
nor U28670 (N_28670,N_28486,N_28454);
xnor U28671 (N_28671,N_28444,N_28261);
nor U28672 (N_28672,N_28359,N_28258);
xnor U28673 (N_28673,N_28445,N_28277);
nor U28674 (N_28674,N_28493,N_28358);
xor U28675 (N_28675,N_28393,N_28469);
and U28676 (N_28676,N_28331,N_28446);
or U28677 (N_28677,N_28254,N_28476);
or U28678 (N_28678,N_28321,N_28355);
nor U28679 (N_28679,N_28297,N_28466);
and U28680 (N_28680,N_28267,N_28382);
xor U28681 (N_28681,N_28452,N_28354);
or U28682 (N_28682,N_28487,N_28323);
nand U28683 (N_28683,N_28256,N_28251);
nor U28684 (N_28684,N_28492,N_28372);
nand U28685 (N_28685,N_28354,N_28276);
or U28686 (N_28686,N_28415,N_28331);
xnor U28687 (N_28687,N_28317,N_28267);
nand U28688 (N_28688,N_28332,N_28271);
or U28689 (N_28689,N_28489,N_28317);
nor U28690 (N_28690,N_28497,N_28287);
xnor U28691 (N_28691,N_28499,N_28473);
or U28692 (N_28692,N_28391,N_28357);
nand U28693 (N_28693,N_28291,N_28457);
nand U28694 (N_28694,N_28452,N_28391);
nand U28695 (N_28695,N_28263,N_28433);
nor U28696 (N_28696,N_28414,N_28397);
nor U28697 (N_28697,N_28299,N_28378);
and U28698 (N_28698,N_28479,N_28496);
nand U28699 (N_28699,N_28311,N_28295);
nor U28700 (N_28700,N_28283,N_28302);
or U28701 (N_28701,N_28357,N_28419);
and U28702 (N_28702,N_28295,N_28322);
or U28703 (N_28703,N_28375,N_28487);
nand U28704 (N_28704,N_28428,N_28418);
nor U28705 (N_28705,N_28336,N_28457);
nor U28706 (N_28706,N_28438,N_28365);
nor U28707 (N_28707,N_28400,N_28326);
nor U28708 (N_28708,N_28463,N_28368);
and U28709 (N_28709,N_28277,N_28490);
nor U28710 (N_28710,N_28359,N_28493);
or U28711 (N_28711,N_28296,N_28449);
xnor U28712 (N_28712,N_28301,N_28257);
xnor U28713 (N_28713,N_28373,N_28492);
xnor U28714 (N_28714,N_28267,N_28476);
nor U28715 (N_28715,N_28433,N_28477);
nand U28716 (N_28716,N_28493,N_28270);
nor U28717 (N_28717,N_28332,N_28299);
xnor U28718 (N_28718,N_28404,N_28430);
or U28719 (N_28719,N_28454,N_28465);
xor U28720 (N_28720,N_28365,N_28256);
xnor U28721 (N_28721,N_28372,N_28296);
and U28722 (N_28722,N_28482,N_28314);
xnor U28723 (N_28723,N_28356,N_28379);
xor U28724 (N_28724,N_28285,N_28461);
and U28725 (N_28725,N_28452,N_28263);
xnor U28726 (N_28726,N_28347,N_28342);
nor U28727 (N_28727,N_28362,N_28290);
xor U28728 (N_28728,N_28481,N_28303);
nor U28729 (N_28729,N_28405,N_28400);
or U28730 (N_28730,N_28351,N_28443);
nor U28731 (N_28731,N_28476,N_28354);
and U28732 (N_28732,N_28386,N_28481);
nand U28733 (N_28733,N_28409,N_28357);
or U28734 (N_28734,N_28479,N_28270);
nand U28735 (N_28735,N_28390,N_28475);
nor U28736 (N_28736,N_28357,N_28396);
and U28737 (N_28737,N_28436,N_28358);
nor U28738 (N_28738,N_28388,N_28324);
and U28739 (N_28739,N_28253,N_28485);
xor U28740 (N_28740,N_28307,N_28414);
xor U28741 (N_28741,N_28418,N_28379);
and U28742 (N_28742,N_28272,N_28475);
nand U28743 (N_28743,N_28470,N_28398);
xor U28744 (N_28744,N_28460,N_28310);
nor U28745 (N_28745,N_28429,N_28287);
and U28746 (N_28746,N_28283,N_28451);
xor U28747 (N_28747,N_28309,N_28362);
nor U28748 (N_28748,N_28368,N_28497);
and U28749 (N_28749,N_28432,N_28297);
xor U28750 (N_28750,N_28749,N_28554);
or U28751 (N_28751,N_28703,N_28654);
nand U28752 (N_28752,N_28687,N_28607);
nand U28753 (N_28753,N_28680,N_28747);
xnor U28754 (N_28754,N_28558,N_28727);
or U28755 (N_28755,N_28663,N_28579);
and U28756 (N_28756,N_28596,N_28633);
xnor U28757 (N_28757,N_28668,N_28734);
nand U28758 (N_28758,N_28737,N_28603);
nand U28759 (N_28759,N_28677,N_28748);
xor U28760 (N_28760,N_28635,N_28509);
nand U28761 (N_28761,N_28672,N_28524);
nor U28762 (N_28762,N_28643,N_28627);
nor U28763 (N_28763,N_28743,N_28656);
nor U28764 (N_28764,N_28523,N_28712);
and U28765 (N_28765,N_28662,N_28539);
nor U28766 (N_28766,N_28546,N_28729);
or U28767 (N_28767,N_28665,N_28700);
or U28768 (N_28768,N_28718,N_28527);
nor U28769 (N_28769,N_28653,N_28659);
or U28770 (N_28770,N_28536,N_28722);
and U28771 (N_28771,N_28642,N_28544);
and U28772 (N_28772,N_28724,N_28689);
and U28773 (N_28773,N_28738,N_28549);
or U28774 (N_28774,N_28624,N_28726);
xnor U28775 (N_28775,N_28553,N_28531);
nand U28776 (N_28776,N_28513,N_28664);
or U28777 (N_28777,N_28696,N_28593);
nor U28778 (N_28778,N_28719,N_28511);
xnor U28779 (N_28779,N_28508,N_28715);
nand U28780 (N_28780,N_28601,N_28552);
nor U28781 (N_28781,N_28728,N_28503);
nor U28782 (N_28782,N_28604,N_28615);
and U28783 (N_28783,N_28500,N_28583);
nor U28784 (N_28784,N_28555,N_28660);
nor U28785 (N_28785,N_28651,N_28564);
nand U28786 (N_28786,N_28745,N_28620);
nor U28787 (N_28787,N_28691,N_28530);
or U28788 (N_28788,N_28534,N_28688);
nand U28789 (N_28789,N_28697,N_28577);
or U28790 (N_28790,N_28504,N_28704);
and U28791 (N_28791,N_28512,N_28515);
xor U28792 (N_28792,N_28517,N_28600);
nand U28793 (N_28793,N_28637,N_28625);
nor U28794 (N_28794,N_28505,N_28575);
nor U28795 (N_28795,N_28709,N_28641);
and U28796 (N_28796,N_28667,N_28639);
xor U28797 (N_28797,N_28671,N_28721);
and U28798 (N_28798,N_28645,N_28650);
and U28799 (N_28799,N_28739,N_28613);
or U28800 (N_28800,N_28649,N_28580);
or U28801 (N_28801,N_28698,N_28661);
xor U28802 (N_28802,N_28655,N_28589);
xor U28803 (N_28803,N_28547,N_28699);
nand U28804 (N_28804,N_28587,N_28540);
nor U28805 (N_28805,N_28702,N_28548);
and U28806 (N_28806,N_28638,N_28507);
xor U28807 (N_28807,N_28675,N_28502);
and U28808 (N_28808,N_28629,N_28525);
nor U28809 (N_28809,N_28682,N_28679);
xor U28810 (N_28810,N_28520,N_28740);
and U28811 (N_28811,N_28588,N_28717);
nand U28812 (N_28812,N_28622,N_28658);
nor U28813 (N_28813,N_28632,N_28617);
nand U28814 (N_28814,N_28648,N_28529);
nand U28815 (N_28815,N_28666,N_28736);
nand U28816 (N_28816,N_28640,N_28652);
xnor U28817 (N_28817,N_28605,N_28646);
and U28818 (N_28818,N_28518,N_28621);
and U28819 (N_28819,N_28686,N_28674);
nor U28820 (N_28820,N_28541,N_28570);
xnor U28821 (N_28821,N_28574,N_28537);
xor U28822 (N_28822,N_28506,N_28522);
or U28823 (N_28823,N_28733,N_28744);
or U28824 (N_28824,N_28619,N_28592);
and U28825 (N_28825,N_28708,N_28731);
or U28826 (N_28826,N_28562,N_28521);
or U28827 (N_28827,N_28669,N_28628);
xnor U28828 (N_28828,N_28705,N_28578);
nand U28829 (N_28829,N_28585,N_28647);
and U28830 (N_28830,N_28586,N_28706);
or U28831 (N_28831,N_28730,N_28673);
and U28832 (N_28832,N_28742,N_28636);
and U28833 (N_28833,N_28678,N_28519);
nand U28834 (N_28834,N_28543,N_28631);
and U28835 (N_28835,N_28685,N_28538);
nor U28836 (N_28836,N_28701,N_28606);
xnor U28837 (N_28837,N_28569,N_28514);
nand U28838 (N_28838,N_28550,N_28532);
xor U28839 (N_28839,N_28535,N_28657);
xnor U28840 (N_28840,N_28608,N_28609);
and U28841 (N_28841,N_28713,N_28711);
and U28842 (N_28842,N_28746,N_28741);
or U28843 (N_28843,N_28557,N_28723);
xnor U28844 (N_28844,N_28732,N_28611);
and U28845 (N_28845,N_28567,N_28581);
nand U28846 (N_28846,N_28681,N_28510);
xor U28847 (N_28847,N_28714,N_28594);
xor U28848 (N_28848,N_28602,N_28599);
xnor U28849 (N_28849,N_28610,N_28568);
or U28850 (N_28850,N_28571,N_28695);
xor U28851 (N_28851,N_28551,N_28556);
and U28852 (N_28852,N_28725,N_28693);
nor U28853 (N_28853,N_28612,N_28683);
nand U28854 (N_28854,N_28545,N_28584);
nor U28855 (N_28855,N_28563,N_28566);
nand U28856 (N_28856,N_28501,N_28684);
and U28857 (N_28857,N_28533,N_28644);
xor U28858 (N_28858,N_28630,N_28526);
nand U28859 (N_28859,N_28735,N_28720);
nand U28860 (N_28860,N_28626,N_28670);
nand U28861 (N_28861,N_28516,N_28710);
nand U28862 (N_28862,N_28561,N_28576);
nand U28863 (N_28863,N_28676,N_28559);
nand U28864 (N_28864,N_28595,N_28565);
nor U28865 (N_28865,N_28528,N_28694);
or U28866 (N_28866,N_28692,N_28618);
xnor U28867 (N_28867,N_28634,N_28597);
or U28868 (N_28868,N_28572,N_28690);
or U28869 (N_28869,N_28542,N_28560);
nor U28870 (N_28870,N_28582,N_28573);
and U28871 (N_28871,N_28591,N_28707);
and U28872 (N_28872,N_28716,N_28598);
xnor U28873 (N_28873,N_28623,N_28616);
nand U28874 (N_28874,N_28614,N_28590);
and U28875 (N_28875,N_28533,N_28601);
nor U28876 (N_28876,N_28587,N_28518);
and U28877 (N_28877,N_28713,N_28594);
xnor U28878 (N_28878,N_28627,N_28748);
and U28879 (N_28879,N_28546,N_28723);
nor U28880 (N_28880,N_28721,N_28550);
nor U28881 (N_28881,N_28636,N_28587);
nor U28882 (N_28882,N_28745,N_28689);
nor U28883 (N_28883,N_28519,N_28732);
xnor U28884 (N_28884,N_28515,N_28712);
xor U28885 (N_28885,N_28643,N_28673);
nand U28886 (N_28886,N_28590,N_28588);
nand U28887 (N_28887,N_28658,N_28703);
and U28888 (N_28888,N_28505,N_28600);
nor U28889 (N_28889,N_28734,N_28566);
or U28890 (N_28890,N_28711,N_28525);
nor U28891 (N_28891,N_28505,N_28725);
nand U28892 (N_28892,N_28714,N_28510);
xor U28893 (N_28893,N_28500,N_28698);
nand U28894 (N_28894,N_28569,N_28528);
nand U28895 (N_28895,N_28544,N_28603);
or U28896 (N_28896,N_28680,N_28655);
xor U28897 (N_28897,N_28599,N_28640);
and U28898 (N_28898,N_28611,N_28575);
nand U28899 (N_28899,N_28679,N_28720);
or U28900 (N_28900,N_28533,N_28661);
and U28901 (N_28901,N_28669,N_28577);
nand U28902 (N_28902,N_28703,N_28517);
or U28903 (N_28903,N_28679,N_28604);
or U28904 (N_28904,N_28539,N_28554);
xor U28905 (N_28905,N_28719,N_28622);
nor U28906 (N_28906,N_28639,N_28532);
or U28907 (N_28907,N_28550,N_28656);
and U28908 (N_28908,N_28715,N_28647);
nor U28909 (N_28909,N_28541,N_28537);
xor U28910 (N_28910,N_28551,N_28723);
nor U28911 (N_28911,N_28539,N_28727);
or U28912 (N_28912,N_28638,N_28541);
nand U28913 (N_28913,N_28568,N_28533);
xor U28914 (N_28914,N_28719,N_28720);
and U28915 (N_28915,N_28725,N_28740);
or U28916 (N_28916,N_28586,N_28730);
xor U28917 (N_28917,N_28725,N_28728);
nor U28918 (N_28918,N_28501,N_28517);
nor U28919 (N_28919,N_28742,N_28550);
or U28920 (N_28920,N_28546,N_28610);
nor U28921 (N_28921,N_28652,N_28728);
or U28922 (N_28922,N_28673,N_28690);
or U28923 (N_28923,N_28549,N_28719);
and U28924 (N_28924,N_28740,N_28733);
or U28925 (N_28925,N_28639,N_28518);
nand U28926 (N_28926,N_28548,N_28647);
and U28927 (N_28927,N_28680,N_28693);
and U28928 (N_28928,N_28727,N_28593);
nand U28929 (N_28929,N_28703,N_28522);
nor U28930 (N_28930,N_28500,N_28577);
and U28931 (N_28931,N_28725,N_28684);
and U28932 (N_28932,N_28504,N_28536);
xor U28933 (N_28933,N_28564,N_28740);
xor U28934 (N_28934,N_28690,N_28611);
nand U28935 (N_28935,N_28717,N_28678);
xor U28936 (N_28936,N_28608,N_28590);
nor U28937 (N_28937,N_28546,N_28531);
nor U28938 (N_28938,N_28749,N_28716);
and U28939 (N_28939,N_28600,N_28576);
nand U28940 (N_28940,N_28647,N_28529);
and U28941 (N_28941,N_28656,N_28664);
or U28942 (N_28942,N_28664,N_28658);
or U28943 (N_28943,N_28728,N_28568);
or U28944 (N_28944,N_28723,N_28545);
or U28945 (N_28945,N_28587,N_28728);
xor U28946 (N_28946,N_28596,N_28505);
and U28947 (N_28947,N_28730,N_28569);
nand U28948 (N_28948,N_28529,N_28506);
and U28949 (N_28949,N_28547,N_28600);
xor U28950 (N_28950,N_28638,N_28608);
xor U28951 (N_28951,N_28624,N_28676);
xor U28952 (N_28952,N_28719,N_28739);
xnor U28953 (N_28953,N_28602,N_28686);
nor U28954 (N_28954,N_28581,N_28668);
xor U28955 (N_28955,N_28701,N_28739);
and U28956 (N_28956,N_28578,N_28582);
and U28957 (N_28957,N_28707,N_28509);
nor U28958 (N_28958,N_28707,N_28729);
and U28959 (N_28959,N_28743,N_28556);
and U28960 (N_28960,N_28650,N_28552);
or U28961 (N_28961,N_28523,N_28643);
xnor U28962 (N_28962,N_28699,N_28559);
nand U28963 (N_28963,N_28539,N_28588);
nand U28964 (N_28964,N_28747,N_28596);
xnor U28965 (N_28965,N_28642,N_28598);
and U28966 (N_28966,N_28677,N_28663);
and U28967 (N_28967,N_28642,N_28639);
or U28968 (N_28968,N_28613,N_28730);
and U28969 (N_28969,N_28719,N_28502);
nor U28970 (N_28970,N_28540,N_28523);
nand U28971 (N_28971,N_28561,N_28625);
nor U28972 (N_28972,N_28572,N_28621);
nand U28973 (N_28973,N_28623,N_28558);
and U28974 (N_28974,N_28649,N_28733);
xor U28975 (N_28975,N_28737,N_28728);
and U28976 (N_28976,N_28526,N_28712);
nor U28977 (N_28977,N_28582,N_28629);
nand U28978 (N_28978,N_28676,N_28625);
nor U28979 (N_28979,N_28581,N_28584);
or U28980 (N_28980,N_28513,N_28531);
nor U28981 (N_28981,N_28673,N_28747);
nand U28982 (N_28982,N_28727,N_28677);
xor U28983 (N_28983,N_28586,N_28721);
nor U28984 (N_28984,N_28734,N_28535);
xnor U28985 (N_28985,N_28688,N_28693);
xnor U28986 (N_28986,N_28657,N_28687);
or U28987 (N_28987,N_28669,N_28518);
nor U28988 (N_28988,N_28526,N_28663);
nand U28989 (N_28989,N_28659,N_28635);
and U28990 (N_28990,N_28724,N_28648);
nor U28991 (N_28991,N_28622,N_28536);
and U28992 (N_28992,N_28745,N_28748);
nor U28993 (N_28993,N_28706,N_28527);
xnor U28994 (N_28994,N_28598,N_28685);
xnor U28995 (N_28995,N_28546,N_28722);
nand U28996 (N_28996,N_28580,N_28698);
nand U28997 (N_28997,N_28694,N_28555);
or U28998 (N_28998,N_28714,N_28538);
nand U28999 (N_28999,N_28585,N_28668);
and U29000 (N_29000,N_28917,N_28884);
and U29001 (N_29001,N_28873,N_28838);
xor U29002 (N_29002,N_28781,N_28812);
xor U29003 (N_29003,N_28948,N_28989);
or U29004 (N_29004,N_28936,N_28877);
xnor U29005 (N_29005,N_28758,N_28777);
xor U29006 (N_29006,N_28928,N_28864);
and U29007 (N_29007,N_28831,N_28800);
and U29008 (N_29008,N_28760,N_28820);
nand U29009 (N_29009,N_28931,N_28938);
xor U29010 (N_29010,N_28910,N_28954);
nor U29011 (N_29011,N_28755,N_28809);
or U29012 (N_29012,N_28813,N_28814);
nand U29013 (N_29013,N_28801,N_28834);
nand U29014 (N_29014,N_28935,N_28966);
xnor U29015 (N_29015,N_28985,N_28793);
and U29016 (N_29016,N_28836,N_28763);
or U29017 (N_29017,N_28778,N_28904);
nor U29018 (N_29018,N_28851,N_28880);
nor U29019 (N_29019,N_28789,N_28782);
nand U29020 (N_29020,N_28824,N_28762);
nor U29021 (N_29021,N_28891,N_28817);
nor U29022 (N_29022,N_28912,N_28811);
nor U29023 (N_29023,N_28840,N_28772);
nand U29024 (N_29024,N_28861,N_28850);
nand U29025 (N_29025,N_28988,N_28855);
xnor U29026 (N_29026,N_28771,N_28906);
xnor U29027 (N_29027,N_28983,N_28788);
xnor U29028 (N_29028,N_28865,N_28862);
or U29029 (N_29029,N_28879,N_28795);
nor U29030 (N_29030,N_28815,N_28791);
xor U29031 (N_29031,N_28960,N_28892);
nor U29032 (N_29032,N_28970,N_28952);
or U29033 (N_29033,N_28962,N_28969);
xnor U29034 (N_29034,N_28830,N_28909);
or U29035 (N_29035,N_28900,N_28914);
xnor U29036 (N_29036,N_28926,N_28981);
or U29037 (N_29037,N_28849,N_28802);
nor U29038 (N_29038,N_28869,N_28991);
nand U29039 (N_29039,N_28761,N_28959);
nor U29040 (N_29040,N_28887,N_28816);
nand U29041 (N_29041,N_28833,N_28986);
xnor U29042 (N_29042,N_28907,N_28957);
xnor U29043 (N_29043,N_28796,N_28965);
and U29044 (N_29044,N_28876,N_28823);
or U29045 (N_29045,N_28799,N_28953);
or U29046 (N_29046,N_28947,N_28921);
and U29047 (N_29047,N_28895,N_28845);
nor U29048 (N_29048,N_28896,N_28951);
nor U29049 (N_29049,N_28908,N_28803);
xnor U29050 (N_29050,N_28774,N_28916);
or U29051 (N_29051,N_28819,N_28930);
or U29052 (N_29052,N_28770,N_28806);
nor U29053 (N_29053,N_28842,N_28853);
xor U29054 (N_29054,N_28955,N_28792);
nor U29055 (N_29055,N_28786,N_28958);
nor U29056 (N_29056,N_28875,N_28751);
nand U29057 (N_29057,N_28808,N_28780);
nor U29058 (N_29058,N_28797,N_28994);
xor U29059 (N_29059,N_28956,N_28856);
nor U29060 (N_29060,N_28943,N_28881);
and U29061 (N_29061,N_28848,N_28868);
nand U29062 (N_29062,N_28903,N_28934);
nor U29063 (N_29063,N_28753,N_28790);
or U29064 (N_29064,N_28993,N_28882);
nand U29065 (N_29065,N_28978,N_28854);
nor U29066 (N_29066,N_28911,N_28996);
nor U29067 (N_29067,N_28886,N_28852);
xor U29068 (N_29068,N_28870,N_28963);
xor U29069 (N_29069,N_28804,N_28915);
nor U29070 (N_29070,N_28843,N_28967);
or U29071 (N_29071,N_28999,N_28920);
nand U29072 (N_29072,N_28766,N_28929);
and U29073 (N_29073,N_28961,N_28807);
nor U29074 (N_29074,N_28767,N_28764);
or U29075 (N_29075,N_28905,N_28773);
nand U29076 (N_29076,N_28899,N_28769);
and U29077 (N_29077,N_28940,N_28894);
xor U29078 (N_29078,N_28827,N_28846);
nor U29079 (N_29079,N_28982,N_28984);
and U29080 (N_29080,N_28998,N_28902);
and U29081 (N_29081,N_28839,N_28810);
nand U29082 (N_29082,N_28874,N_28942);
nand U29083 (N_29083,N_28979,N_28866);
xnor U29084 (N_29084,N_28941,N_28901);
xnor U29085 (N_29085,N_28923,N_28785);
and U29086 (N_29086,N_28784,N_28939);
nand U29087 (N_29087,N_28997,N_28783);
xor U29088 (N_29088,N_28835,N_28925);
xor U29089 (N_29089,N_28933,N_28837);
and U29090 (N_29090,N_28847,N_28757);
nand U29091 (N_29091,N_28898,N_28768);
or U29092 (N_29092,N_28752,N_28924);
nor U29093 (N_29093,N_28945,N_28859);
nor U29094 (N_29094,N_28756,N_28841);
and U29095 (N_29095,N_28974,N_28971);
nand U29096 (N_29096,N_28775,N_28821);
and U29097 (N_29097,N_28828,N_28822);
and U29098 (N_29098,N_28950,N_28863);
xnor U29099 (N_29099,N_28949,N_28867);
xor U29100 (N_29100,N_28826,N_28975);
or U29101 (N_29101,N_28890,N_28832);
or U29102 (N_29102,N_28927,N_28829);
nand U29103 (N_29103,N_28992,N_28977);
and U29104 (N_29104,N_28932,N_28897);
nor U29105 (N_29105,N_28976,N_28919);
or U29106 (N_29106,N_28765,N_28787);
nor U29107 (N_29107,N_28871,N_28922);
nand U29108 (N_29108,N_28878,N_28858);
nor U29109 (N_29109,N_28779,N_28805);
nand U29110 (N_29110,N_28759,N_28844);
xnor U29111 (N_29111,N_28825,N_28995);
nand U29112 (N_29112,N_28937,N_28972);
nand U29113 (N_29113,N_28990,N_28980);
xor U29114 (N_29114,N_28885,N_28860);
nor U29115 (N_29115,N_28893,N_28883);
nor U29116 (N_29116,N_28776,N_28794);
xnor U29117 (N_29117,N_28872,N_28818);
or U29118 (N_29118,N_28913,N_28918);
nor U29119 (N_29119,N_28964,N_28946);
and U29120 (N_29120,N_28754,N_28889);
xnor U29121 (N_29121,N_28973,N_28857);
nand U29122 (N_29122,N_28798,N_28944);
or U29123 (N_29123,N_28750,N_28888);
nand U29124 (N_29124,N_28968,N_28987);
nand U29125 (N_29125,N_28921,N_28848);
xnor U29126 (N_29126,N_28832,N_28824);
nand U29127 (N_29127,N_28876,N_28834);
nor U29128 (N_29128,N_28886,N_28795);
and U29129 (N_29129,N_28915,N_28907);
nor U29130 (N_29130,N_28787,N_28994);
nor U29131 (N_29131,N_28947,N_28784);
nand U29132 (N_29132,N_28928,N_28808);
or U29133 (N_29133,N_28852,N_28959);
or U29134 (N_29134,N_28788,N_28996);
or U29135 (N_29135,N_28826,N_28995);
or U29136 (N_29136,N_28975,N_28941);
or U29137 (N_29137,N_28931,N_28791);
and U29138 (N_29138,N_28814,N_28865);
nand U29139 (N_29139,N_28915,N_28862);
nand U29140 (N_29140,N_28903,N_28806);
and U29141 (N_29141,N_28908,N_28884);
nand U29142 (N_29142,N_28952,N_28785);
and U29143 (N_29143,N_28965,N_28945);
nand U29144 (N_29144,N_28989,N_28992);
or U29145 (N_29145,N_28831,N_28757);
xor U29146 (N_29146,N_28866,N_28940);
and U29147 (N_29147,N_28804,N_28837);
nand U29148 (N_29148,N_28801,N_28794);
nor U29149 (N_29149,N_28953,N_28998);
nand U29150 (N_29150,N_28949,N_28766);
and U29151 (N_29151,N_28758,N_28877);
xnor U29152 (N_29152,N_28791,N_28909);
nor U29153 (N_29153,N_28844,N_28908);
or U29154 (N_29154,N_28751,N_28985);
and U29155 (N_29155,N_28811,N_28851);
and U29156 (N_29156,N_28862,N_28947);
nand U29157 (N_29157,N_28937,N_28985);
nor U29158 (N_29158,N_28898,N_28925);
or U29159 (N_29159,N_28804,N_28836);
nor U29160 (N_29160,N_28878,N_28991);
and U29161 (N_29161,N_28994,N_28798);
nand U29162 (N_29162,N_28905,N_28853);
and U29163 (N_29163,N_28947,N_28804);
xor U29164 (N_29164,N_28805,N_28839);
xor U29165 (N_29165,N_28762,N_28893);
nand U29166 (N_29166,N_28768,N_28851);
or U29167 (N_29167,N_28919,N_28859);
and U29168 (N_29168,N_28983,N_28923);
nand U29169 (N_29169,N_28826,N_28893);
xor U29170 (N_29170,N_28911,N_28990);
or U29171 (N_29171,N_28761,N_28767);
nor U29172 (N_29172,N_28820,N_28789);
nand U29173 (N_29173,N_28816,N_28810);
xnor U29174 (N_29174,N_28845,N_28890);
nor U29175 (N_29175,N_28872,N_28959);
or U29176 (N_29176,N_28992,N_28803);
xor U29177 (N_29177,N_28844,N_28770);
nand U29178 (N_29178,N_28863,N_28916);
nand U29179 (N_29179,N_28902,N_28949);
or U29180 (N_29180,N_28772,N_28905);
nand U29181 (N_29181,N_28997,N_28857);
xnor U29182 (N_29182,N_28823,N_28814);
or U29183 (N_29183,N_28794,N_28800);
and U29184 (N_29184,N_28772,N_28876);
nand U29185 (N_29185,N_28972,N_28951);
or U29186 (N_29186,N_28795,N_28831);
or U29187 (N_29187,N_28817,N_28828);
or U29188 (N_29188,N_28848,N_28873);
nor U29189 (N_29189,N_28937,N_28761);
and U29190 (N_29190,N_28951,N_28803);
xnor U29191 (N_29191,N_28856,N_28914);
xnor U29192 (N_29192,N_28809,N_28876);
and U29193 (N_29193,N_28971,N_28940);
xnor U29194 (N_29194,N_28929,N_28975);
nand U29195 (N_29195,N_28778,N_28831);
and U29196 (N_29196,N_28790,N_28997);
nand U29197 (N_29197,N_28989,N_28969);
nand U29198 (N_29198,N_28823,N_28779);
xor U29199 (N_29199,N_28778,N_28788);
nand U29200 (N_29200,N_28789,N_28923);
nor U29201 (N_29201,N_28948,N_28782);
or U29202 (N_29202,N_28840,N_28934);
nand U29203 (N_29203,N_28996,N_28771);
xor U29204 (N_29204,N_28995,N_28781);
nand U29205 (N_29205,N_28945,N_28761);
and U29206 (N_29206,N_28920,N_28965);
and U29207 (N_29207,N_28911,N_28770);
xnor U29208 (N_29208,N_28945,N_28924);
xnor U29209 (N_29209,N_28858,N_28880);
nand U29210 (N_29210,N_28946,N_28836);
or U29211 (N_29211,N_28845,N_28903);
nand U29212 (N_29212,N_28937,N_28844);
nand U29213 (N_29213,N_28795,N_28976);
xnor U29214 (N_29214,N_28938,N_28859);
or U29215 (N_29215,N_28896,N_28925);
xnor U29216 (N_29216,N_28913,N_28800);
nand U29217 (N_29217,N_28865,N_28939);
or U29218 (N_29218,N_28772,N_28958);
nor U29219 (N_29219,N_28919,N_28931);
or U29220 (N_29220,N_28979,N_28767);
nand U29221 (N_29221,N_28793,N_28821);
xor U29222 (N_29222,N_28788,N_28941);
or U29223 (N_29223,N_28799,N_28965);
xor U29224 (N_29224,N_28971,N_28818);
nor U29225 (N_29225,N_28903,N_28933);
nand U29226 (N_29226,N_28989,N_28877);
and U29227 (N_29227,N_28863,N_28898);
and U29228 (N_29228,N_28870,N_28860);
nor U29229 (N_29229,N_28874,N_28987);
nand U29230 (N_29230,N_28998,N_28791);
nand U29231 (N_29231,N_28925,N_28998);
nand U29232 (N_29232,N_28858,N_28786);
nand U29233 (N_29233,N_28800,N_28919);
or U29234 (N_29234,N_28767,N_28822);
xnor U29235 (N_29235,N_28881,N_28909);
xor U29236 (N_29236,N_28910,N_28879);
or U29237 (N_29237,N_28988,N_28984);
xnor U29238 (N_29238,N_28783,N_28931);
xor U29239 (N_29239,N_28818,N_28951);
or U29240 (N_29240,N_28977,N_28978);
or U29241 (N_29241,N_28762,N_28915);
xnor U29242 (N_29242,N_28824,N_28863);
or U29243 (N_29243,N_28894,N_28911);
nand U29244 (N_29244,N_28909,N_28847);
nor U29245 (N_29245,N_28756,N_28821);
nand U29246 (N_29246,N_28959,N_28886);
xor U29247 (N_29247,N_28899,N_28996);
nand U29248 (N_29248,N_28922,N_28931);
xnor U29249 (N_29249,N_28851,N_28817);
and U29250 (N_29250,N_29192,N_29026);
nand U29251 (N_29251,N_29220,N_29193);
nor U29252 (N_29252,N_29178,N_29175);
nand U29253 (N_29253,N_29049,N_29002);
and U29254 (N_29254,N_29007,N_29188);
nand U29255 (N_29255,N_29203,N_29060);
nand U29256 (N_29256,N_29215,N_29098);
nor U29257 (N_29257,N_29083,N_29216);
or U29258 (N_29258,N_29079,N_29039);
or U29259 (N_29259,N_29074,N_29071);
nand U29260 (N_29260,N_29237,N_29044);
or U29261 (N_29261,N_29020,N_29173);
and U29262 (N_29262,N_29244,N_29110);
and U29263 (N_29263,N_29148,N_29003);
xnor U29264 (N_29264,N_29134,N_29153);
or U29265 (N_29265,N_29191,N_29056);
xnor U29266 (N_29266,N_29092,N_29009);
or U29267 (N_29267,N_29243,N_29105);
xnor U29268 (N_29268,N_29168,N_29189);
nand U29269 (N_29269,N_29167,N_29067);
and U29270 (N_29270,N_29053,N_29101);
xnor U29271 (N_29271,N_29121,N_29027);
and U29272 (N_29272,N_29036,N_29024);
xor U29273 (N_29273,N_29022,N_29000);
nor U29274 (N_29274,N_29095,N_29096);
xnor U29275 (N_29275,N_29217,N_29238);
nand U29276 (N_29276,N_29031,N_29144);
and U29277 (N_29277,N_29010,N_29051);
nand U29278 (N_29278,N_29113,N_29207);
xnor U29279 (N_29279,N_29186,N_29120);
nor U29280 (N_29280,N_29091,N_29038);
nand U29281 (N_29281,N_29107,N_29073);
and U29282 (N_29282,N_29177,N_29205);
nand U29283 (N_29283,N_29248,N_29058);
xnor U29284 (N_29284,N_29155,N_29075);
or U29285 (N_29285,N_29057,N_29145);
nand U29286 (N_29286,N_29076,N_29240);
nor U29287 (N_29287,N_29185,N_29055);
and U29288 (N_29288,N_29179,N_29149);
or U29289 (N_29289,N_29032,N_29159);
xnor U29290 (N_29290,N_29034,N_29204);
nor U29291 (N_29291,N_29208,N_29019);
and U29292 (N_29292,N_29194,N_29046);
and U29293 (N_29293,N_29218,N_29233);
xor U29294 (N_29294,N_29234,N_29090);
xnor U29295 (N_29295,N_29164,N_29061);
and U29296 (N_29296,N_29198,N_29135);
xnor U29297 (N_29297,N_29078,N_29229);
and U29298 (N_29298,N_29236,N_29050);
and U29299 (N_29299,N_29176,N_29059);
or U29300 (N_29300,N_29231,N_29108);
and U29301 (N_29301,N_29142,N_29152);
xor U29302 (N_29302,N_29130,N_29085);
nand U29303 (N_29303,N_29111,N_29102);
xnor U29304 (N_29304,N_29161,N_29162);
and U29305 (N_29305,N_29040,N_29239);
or U29306 (N_29306,N_29210,N_29171);
xnor U29307 (N_29307,N_29143,N_29170);
nor U29308 (N_29308,N_29064,N_29223);
or U29309 (N_29309,N_29160,N_29005);
xor U29310 (N_29310,N_29242,N_29147);
nor U29311 (N_29311,N_29118,N_29213);
nand U29312 (N_29312,N_29048,N_29246);
and U29313 (N_29313,N_29077,N_29131);
xnor U29314 (N_29314,N_29182,N_29156);
and U29315 (N_29315,N_29225,N_29140);
nand U29316 (N_29316,N_29114,N_29163);
nor U29317 (N_29317,N_29109,N_29094);
or U29318 (N_29318,N_29137,N_29219);
xnor U29319 (N_29319,N_29212,N_29211);
or U29320 (N_29320,N_29139,N_29017);
nand U29321 (N_29321,N_29041,N_29169);
and U29322 (N_29322,N_29087,N_29070);
and U29323 (N_29323,N_29172,N_29089);
and U29324 (N_29324,N_29245,N_29206);
nor U29325 (N_29325,N_29021,N_29062);
nor U29326 (N_29326,N_29063,N_29150);
nand U29327 (N_29327,N_29069,N_29013);
or U29328 (N_29328,N_29247,N_29081);
or U29329 (N_29329,N_29112,N_29197);
nand U29330 (N_29330,N_29001,N_29146);
xor U29331 (N_29331,N_29093,N_29023);
xnor U29332 (N_29332,N_29209,N_29228);
nand U29333 (N_29333,N_29004,N_29184);
and U29334 (N_29334,N_29099,N_29116);
nand U29335 (N_29335,N_29128,N_29066);
and U29336 (N_29336,N_29181,N_29025);
and U29337 (N_29337,N_29249,N_29086);
nand U29338 (N_29338,N_29043,N_29030);
nor U29339 (N_29339,N_29035,N_29080);
xor U29340 (N_29340,N_29068,N_29084);
nand U29341 (N_29341,N_29166,N_29174);
nor U29342 (N_29342,N_29200,N_29201);
nor U29343 (N_29343,N_29126,N_29119);
or U29344 (N_29344,N_29011,N_29014);
nor U29345 (N_29345,N_29042,N_29065);
and U29346 (N_29346,N_29124,N_29117);
nand U29347 (N_29347,N_29037,N_29227);
and U29348 (N_29348,N_29136,N_29138);
or U29349 (N_29349,N_29052,N_29154);
and U29350 (N_29350,N_29106,N_29100);
and U29351 (N_29351,N_29125,N_29195);
nor U29352 (N_29352,N_29151,N_29123);
nand U29353 (N_29353,N_29006,N_29012);
or U29354 (N_29354,N_29196,N_29033);
or U29355 (N_29355,N_29224,N_29115);
nand U29356 (N_29356,N_29127,N_29104);
nand U29357 (N_29357,N_29157,N_29232);
nor U29358 (N_29358,N_29103,N_29047);
and U29359 (N_29359,N_29190,N_29180);
nand U29360 (N_29360,N_29082,N_29008);
and U29361 (N_29361,N_29018,N_29015);
or U29362 (N_29362,N_29029,N_29214);
and U29363 (N_29363,N_29129,N_29222);
and U29364 (N_29364,N_29165,N_29202);
nor U29365 (N_29365,N_29183,N_29235);
or U29366 (N_29366,N_29221,N_29133);
nand U29367 (N_29367,N_29016,N_29097);
xor U29368 (N_29368,N_29122,N_29132);
or U29369 (N_29369,N_29054,N_29230);
nand U29370 (N_29370,N_29072,N_29028);
nor U29371 (N_29371,N_29158,N_29226);
and U29372 (N_29372,N_29088,N_29187);
or U29373 (N_29373,N_29199,N_29141);
and U29374 (N_29374,N_29241,N_29045);
nor U29375 (N_29375,N_29010,N_29221);
xnor U29376 (N_29376,N_29203,N_29221);
nand U29377 (N_29377,N_29197,N_29068);
or U29378 (N_29378,N_29008,N_29166);
nor U29379 (N_29379,N_29124,N_29157);
or U29380 (N_29380,N_29127,N_29100);
and U29381 (N_29381,N_29119,N_29156);
or U29382 (N_29382,N_29035,N_29205);
nand U29383 (N_29383,N_29226,N_29084);
nand U29384 (N_29384,N_29149,N_29048);
or U29385 (N_29385,N_29120,N_29167);
nor U29386 (N_29386,N_29156,N_29160);
nand U29387 (N_29387,N_29127,N_29077);
and U29388 (N_29388,N_29019,N_29098);
and U29389 (N_29389,N_29003,N_29138);
xor U29390 (N_29390,N_29018,N_29074);
nor U29391 (N_29391,N_29226,N_29065);
xor U29392 (N_29392,N_29170,N_29190);
and U29393 (N_29393,N_29225,N_29072);
or U29394 (N_29394,N_29021,N_29121);
or U29395 (N_29395,N_29039,N_29204);
nor U29396 (N_29396,N_29040,N_29088);
nor U29397 (N_29397,N_29030,N_29135);
nor U29398 (N_29398,N_29176,N_29194);
nor U29399 (N_29399,N_29106,N_29228);
nand U29400 (N_29400,N_29003,N_29036);
nor U29401 (N_29401,N_29168,N_29214);
and U29402 (N_29402,N_29005,N_29068);
nor U29403 (N_29403,N_29192,N_29075);
and U29404 (N_29404,N_29063,N_29082);
and U29405 (N_29405,N_29158,N_29089);
nand U29406 (N_29406,N_29122,N_29041);
nand U29407 (N_29407,N_29100,N_29212);
nor U29408 (N_29408,N_29199,N_29225);
xnor U29409 (N_29409,N_29126,N_29060);
or U29410 (N_29410,N_29202,N_29174);
and U29411 (N_29411,N_29111,N_29246);
or U29412 (N_29412,N_29241,N_29059);
xor U29413 (N_29413,N_29049,N_29095);
or U29414 (N_29414,N_29219,N_29249);
xor U29415 (N_29415,N_29065,N_29228);
or U29416 (N_29416,N_29085,N_29013);
and U29417 (N_29417,N_29062,N_29075);
and U29418 (N_29418,N_29163,N_29165);
or U29419 (N_29419,N_29240,N_29242);
nand U29420 (N_29420,N_29018,N_29019);
xor U29421 (N_29421,N_29101,N_29241);
nor U29422 (N_29422,N_29234,N_29038);
nor U29423 (N_29423,N_29025,N_29018);
or U29424 (N_29424,N_29012,N_29247);
and U29425 (N_29425,N_29041,N_29247);
or U29426 (N_29426,N_29067,N_29106);
nor U29427 (N_29427,N_29224,N_29235);
and U29428 (N_29428,N_29214,N_29244);
nand U29429 (N_29429,N_29242,N_29095);
nand U29430 (N_29430,N_29109,N_29058);
nor U29431 (N_29431,N_29071,N_29007);
and U29432 (N_29432,N_29114,N_29039);
nand U29433 (N_29433,N_29104,N_29016);
xor U29434 (N_29434,N_29100,N_29172);
nor U29435 (N_29435,N_29077,N_29004);
and U29436 (N_29436,N_29186,N_29066);
nand U29437 (N_29437,N_29109,N_29153);
and U29438 (N_29438,N_29007,N_29238);
nor U29439 (N_29439,N_29198,N_29212);
or U29440 (N_29440,N_29134,N_29073);
and U29441 (N_29441,N_29169,N_29060);
and U29442 (N_29442,N_29028,N_29048);
and U29443 (N_29443,N_29181,N_29023);
and U29444 (N_29444,N_29170,N_29020);
nor U29445 (N_29445,N_29243,N_29024);
nor U29446 (N_29446,N_29242,N_29224);
and U29447 (N_29447,N_29105,N_29196);
and U29448 (N_29448,N_29116,N_29179);
nor U29449 (N_29449,N_29107,N_29034);
nor U29450 (N_29450,N_29248,N_29080);
or U29451 (N_29451,N_29087,N_29016);
nor U29452 (N_29452,N_29019,N_29074);
or U29453 (N_29453,N_29036,N_29028);
nand U29454 (N_29454,N_29219,N_29079);
and U29455 (N_29455,N_29236,N_29185);
or U29456 (N_29456,N_29046,N_29037);
or U29457 (N_29457,N_29215,N_29205);
xor U29458 (N_29458,N_29227,N_29061);
nor U29459 (N_29459,N_29131,N_29110);
nand U29460 (N_29460,N_29065,N_29170);
xor U29461 (N_29461,N_29160,N_29100);
nand U29462 (N_29462,N_29155,N_29234);
xor U29463 (N_29463,N_29191,N_29024);
nor U29464 (N_29464,N_29115,N_29133);
nand U29465 (N_29465,N_29159,N_29230);
or U29466 (N_29466,N_29037,N_29172);
and U29467 (N_29467,N_29184,N_29190);
xnor U29468 (N_29468,N_29188,N_29034);
nor U29469 (N_29469,N_29044,N_29083);
nor U29470 (N_29470,N_29123,N_29156);
xnor U29471 (N_29471,N_29079,N_29152);
nand U29472 (N_29472,N_29053,N_29153);
and U29473 (N_29473,N_29247,N_29227);
nor U29474 (N_29474,N_29156,N_29109);
xor U29475 (N_29475,N_29205,N_29187);
nor U29476 (N_29476,N_29147,N_29247);
xnor U29477 (N_29477,N_29202,N_29111);
nand U29478 (N_29478,N_29082,N_29238);
and U29479 (N_29479,N_29069,N_29219);
nand U29480 (N_29480,N_29044,N_29154);
xnor U29481 (N_29481,N_29200,N_29170);
nor U29482 (N_29482,N_29246,N_29134);
nor U29483 (N_29483,N_29046,N_29138);
and U29484 (N_29484,N_29227,N_29029);
nor U29485 (N_29485,N_29093,N_29099);
nor U29486 (N_29486,N_29023,N_29183);
nor U29487 (N_29487,N_29231,N_29076);
xnor U29488 (N_29488,N_29102,N_29020);
nor U29489 (N_29489,N_29126,N_29160);
or U29490 (N_29490,N_29213,N_29026);
nor U29491 (N_29491,N_29168,N_29096);
nor U29492 (N_29492,N_29018,N_29006);
xor U29493 (N_29493,N_29240,N_29078);
xnor U29494 (N_29494,N_29006,N_29204);
xnor U29495 (N_29495,N_29223,N_29128);
nor U29496 (N_29496,N_29189,N_29163);
and U29497 (N_29497,N_29182,N_29145);
nor U29498 (N_29498,N_29189,N_29207);
nor U29499 (N_29499,N_29061,N_29003);
and U29500 (N_29500,N_29343,N_29256);
and U29501 (N_29501,N_29496,N_29362);
or U29502 (N_29502,N_29383,N_29366);
nand U29503 (N_29503,N_29375,N_29292);
nor U29504 (N_29504,N_29363,N_29364);
and U29505 (N_29505,N_29463,N_29277);
nand U29506 (N_29506,N_29324,N_29272);
nor U29507 (N_29507,N_29438,N_29384);
nor U29508 (N_29508,N_29333,N_29477);
or U29509 (N_29509,N_29259,N_29453);
nor U29510 (N_29510,N_29287,N_29318);
xnor U29511 (N_29511,N_29422,N_29392);
or U29512 (N_29512,N_29421,N_29338);
nand U29513 (N_29513,N_29388,N_29452);
xor U29514 (N_29514,N_29491,N_29300);
nand U29515 (N_29515,N_29447,N_29429);
and U29516 (N_29516,N_29327,N_29393);
and U29517 (N_29517,N_29252,N_29387);
nor U29518 (N_29518,N_29400,N_29328);
or U29519 (N_29519,N_29341,N_29346);
nor U29520 (N_29520,N_29270,N_29374);
nor U29521 (N_29521,N_29345,N_29425);
nand U29522 (N_29522,N_29329,N_29444);
and U29523 (N_29523,N_29445,N_29416);
nand U29524 (N_29524,N_29258,N_29257);
nand U29525 (N_29525,N_29320,N_29390);
or U29526 (N_29526,N_29412,N_29464);
and U29527 (N_29527,N_29316,N_29386);
or U29528 (N_29528,N_29378,N_29373);
nand U29529 (N_29529,N_29289,N_29401);
and U29530 (N_29530,N_29462,N_29409);
nand U29531 (N_29531,N_29391,N_29474);
and U29532 (N_29532,N_29467,N_29295);
and U29533 (N_29533,N_29399,N_29377);
xor U29534 (N_29534,N_29348,N_29303);
xnor U29535 (N_29535,N_29396,N_29282);
nor U29536 (N_29536,N_29269,N_29475);
nor U29537 (N_29537,N_29385,N_29273);
or U29538 (N_29538,N_29321,N_29296);
and U29539 (N_29539,N_29441,N_29492);
nand U29540 (N_29540,N_29479,N_29294);
nand U29541 (N_29541,N_29290,N_29426);
and U29542 (N_29542,N_29405,N_29472);
xor U29543 (N_29543,N_29334,N_29495);
and U29544 (N_29544,N_29288,N_29481);
nor U29545 (N_29545,N_29353,N_29354);
or U29546 (N_29546,N_29417,N_29356);
nor U29547 (N_29547,N_29323,N_29315);
nand U29548 (N_29548,N_29434,N_29278);
nor U29549 (N_29549,N_29424,N_29418);
and U29550 (N_29550,N_29493,N_29461);
and U29551 (N_29551,N_29478,N_29284);
nor U29552 (N_29552,N_29326,N_29430);
nor U29553 (N_29553,N_29250,N_29261);
nand U29554 (N_29554,N_29466,N_29442);
xor U29555 (N_29555,N_29439,N_29254);
xor U29556 (N_29556,N_29266,N_29370);
nor U29557 (N_29557,N_29420,N_29317);
nor U29558 (N_29558,N_29280,N_29480);
xor U29559 (N_29559,N_29402,N_29361);
or U29560 (N_29560,N_29360,N_29293);
and U29561 (N_29561,N_29379,N_29414);
nand U29562 (N_29562,N_29415,N_29298);
and U29563 (N_29563,N_29423,N_29313);
xnor U29564 (N_29564,N_29301,N_29335);
nand U29565 (N_29565,N_29260,N_29494);
nand U29566 (N_29566,N_29302,N_29286);
nand U29567 (N_29567,N_29365,N_29397);
nor U29568 (N_29568,N_29368,N_29428);
xnor U29569 (N_29569,N_29465,N_29433);
and U29570 (N_29570,N_29271,N_29275);
nor U29571 (N_29571,N_29255,N_29413);
and U29572 (N_29572,N_29497,N_29331);
and U29573 (N_29573,N_29499,N_29469);
nand U29574 (N_29574,N_29352,N_29304);
and U29575 (N_29575,N_29340,N_29455);
or U29576 (N_29576,N_29406,N_29431);
and U29577 (N_29577,N_29404,N_29367);
or U29578 (N_29578,N_29251,N_29263);
and U29579 (N_29579,N_29344,N_29371);
or U29580 (N_29580,N_29471,N_29468);
nand U29581 (N_29581,N_29381,N_29389);
nand U29582 (N_29582,N_29336,N_29411);
nor U29583 (N_29583,N_29482,N_29395);
nand U29584 (N_29584,N_29299,N_29319);
or U29585 (N_29585,N_29312,N_29274);
or U29586 (N_29586,N_29487,N_29484);
nor U29587 (N_29587,N_29470,N_29349);
nor U29588 (N_29588,N_29262,N_29459);
nor U29589 (N_29589,N_29337,N_29435);
and U29590 (N_29590,N_29398,N_29454);
xnor U29591 (N_29591,N_29253,N_29419);
and U29592 (N_29592,N_29440,N_29308);
or U29593 (N_29593,N_29443,N_29325);
nor U29594 (N_29594,N_29305,N_29486);
nand U29595 (N_29595,N_29460,N_29372);
or U29596 (N_29596,N_29394,N_29357);
nand U29597 (N_29597,N_29490,N_29332);
xnor U29598 (N_29598,N_29279,N_29451);
nor U29599 (N_29599,N_29458,N_29473);
nor U29600 (N_29600,N_29359,N_29285);
or U29601 (N_29601,N_29347,N_29264);
or U29602 (N_29602,N_29498,N_29265);
xor U29603 (N_29603,N_29355,N_29427);
xnor U29604 (N_29604,N_29457,N_29322);
nor U29605 (N_29605,N_29382,N_29488);
nand U29606 (N_29606,N_29310,N_29267);
nand U29607 (N_29607,N_29309,N_29369);
xor U29608 (N_29608,N_29450,N_29403);
xnor U29609 (N_29609,N_29283,N_29483);
nor U29610 (N_29610,N_29311,N_29436);
or U29611 (N_29611,N_29437,N_29485);
nand U29612 (N_29612,N_29276,N_29446);
nand U29613 (N_29613,N_29351,N_29281);
nand U29614 (N_29614,N_29432,N_29268);
or U29615 (N_29615,N_29297,N_29307);
or U29616 (N_29616,N_29407,N_29358);
nor U29617 (N_29617,N_29449,N_29350);
nor U29618 (N_29618,N_29339,N_29314);
nand U29619 (N_29619,N_29410,N_29376);
and U29620 (N_29620,N_29476,N_29456);
nor U29621 (N_29621,N_29291,N_29342);
and U29622 (N_29622,N_29408,N_29330);
xnor U29623 (N_29623,N_29489,N_29306);
and U29624 (N_29624,N_29448,N_29380);
xor U29625 (N_29625,N_29357,N_29408);
nand U29626 (N_29626,N_29270,N_29252);
and U29627 (N_29627,N_29473,N_29409);
xnor U29628 (N_29628,N_29327,N_29445);
nand U29629 (N_29629,N_29426,N_29482);
nor U29630 (N_29630,N_29439,N_29334);
and U29631 (N_29631,N_29370,N_29375);
or U29632 (N_29632,N_29316,N_29320);
or U29633 (N_29633,N_29287,N_29381);
nand U29634 (N_29634,N_29338,N_29405);
nand U29635 (N_29635,N_29416,N_29335);
or U29636 (N_29636,N_29408,N_29399);
nor U29637 (N_29637,N_29297,N_29458);
or U29638 (N_29638,N_29283,N_29355);
xnor U29639 (N_29639,N_29316,N_29407);
nand U29640 (N_29640,N_29297,N_29369);
and U29641 (N_29641,N_29415,N_29346);
or U29642 (N_29642,N_29367,N_29306);
or U29643 (N_29643,N_29409,N_29376);
nor U29644 (N_29644,N_29449,N_29262);
nor U29645 (N_29645,N_29329,N_29436);
or U29646 (N_29646,N_29471,N_29332);
nor U29647 (N_29647,N_29275,N_29417);
xor U29648 (N_29648,N_29404,N_29471);
xor U29649 (N_29649,N_29270,N_29394);
xnor U29650 (N_29650,N_29386,N_29389);
xor U29651 (N_29651,N_29304,N_29254);
or U29652 (N_29652,N_29460,N_29481);
nand U29653 (N_29653,N_29316,N_29450);
or U29654 (N_29654,N_29353,N_29474);
nand U29655 (N_29655,N_29379,N_29354);
nor U29656 (N_29656,N_29430,N_29352);
xnor U29657 (N_29657,N_29486,N_29324);
nor U29658 (N_29658,N_29378,N_29407);
nand U29659 (N_29659,N_29258,N_29297);
nand U29660 (N_29660,N_29488,N_29346);
or U29661 (N_29661,N_29317,N_29254);
nand U29662 (N_29662,N_29280,N_29436);
and U29663 (N_29663,N_29347,N_29478);
nor U29664 (N_29664,N_29426,N_29275);
nor U29665 (N_29665,N_29440,N_29473);
nor U29666 (N_29666,N_29455,N_29445);
nor U29667 (N_29667,N_29396,N_29265);
xnor U29668 (N_29668,N_29286,N_29319);
and U29669 (N_29669,N_29309,N_29261);
xor U29670 (N_29670,N_29269,N_29327);
or U29671 (N_29671,N_29420,N_29414);
xnor U29672 (N_29672,N_29312,N_29421);
nand U29673 (N_29673,N_29413,N_29349);
xor U29674 (N_29674,N_29342,N_29491);
nand U29675 (N_29675,N_29351,N_29324);
and U29676 (N_29676,N_29322,N_29409);
xor U29677 (N_29677,N_29497,N_29255);
nand U29678 (N_29678,N_29318,N_29468);
nor U29679 (N_29679,N_29384,N_29380);
or U29680 (N_29680,N_29404,N_29311);
and U29681 (N_29681,N_29311,N_29486);
nor U29682 (N_29682,N_29306,N_29338);
or U29683 (N_29683,N_29379,N_29385);
or U29684 (N_29684,N_29285,N_29459);
nand U29685 (N_29685,N_29457,N_29295);
xnor U29686 (N_29686,N_29273,N_29397);
xnor U29687 (N_29687,N_29326,N_29280);
nand U29688 (N_29688,N_29487,N_29270);
nor U29689 (N_29689,N_29350,N_29426);
nor U29690 (N_29690,N_29426,N_29252);
or U29691 (N_29691,N_29374,N_29366);
and U29692 (N_29692,N_29274,N_29355);
xor U29693 (N_29693,N_29262,N_29474);
nand U29694 (N_29694,N_29453,N_29350);
or U29695 (N_29695,N_29267,N_29283);
nor U29696 (N_29696,N_29462,N_29304);
nor U29697 (N_29697,N_29332,N_29437);
nor U29698 (N_29698,N_29395,N_29404);
nor U29699 (N_29699,N_29473,N_29489);
nor U29700 (N_29700,N_29340,N_29461);
nand U29701 (N_29701,N_29362,N_29435);
nor U29702 (N_29702,N_29351,N_29403);
nand U29703 (N_29703,N_29350,N_29304);
nor U29704 (N_29704,N_29314,N_29311);
nand U29705 (N_29705,N_29299,N_29255);
nand U29706 (N_29706,N_29453,N_29253);
or U29707 (N_29707,N_29252,N_29473);
and U29708 (N_29708,N_29252,N_29407);
or U29709 (N_29709,N_29467,N_29326);
xor U29710 (N_29710,N_29366,N_29361);
and U29711 (N_29711,N_29368,N_29388);
xor U29712 (N_29712,N_29339,N_29327);
and U29713 (N_29713,N_29437,N_29322);
nand U29714 (N_29714,N_29330,N_29424);
and U29715 (N_29715,N_29404,N_29430);
nand U29716 (N_29716,N_29318,N_29480);
and U29717 (N_29717,N_29301,N_29490);
nor U29718 (N_29718,N_29292,N_29452);
and U29719 (N_29719,N_29279,N_29477);
or U29720 (N_29720,N_29342,N_29348);
nor U29721 (N_29721,N_29412,N_29295);
nor U29722 (N_29722,N_29260,N_29295);
xor U29723 (N_29723,N_29328,N_29435);
and U29724 (N_29724,N_29276,N_29338);
and U29725 (N_29725,N_29298,N_29372);
or U29726 (N_29726,N_29468,N_29326);
and U29727 (N_29727,N_29277,N_29372);
xor U29728 (N_29728,N_29340,N_29419);
xor U29729 (N_29729,N_29481,N_29257);
nand U29730 (N_29730,N_29424,N_29367);
and U29731 (N_29731,N_29301,N_29430);
nor U29732 (N_29732,N_29465,N_29254);
nand U29733 (N_29733,N_29475,N_29406);
nor U29734 (N_29734,N_29253,N_29438);
xor U29735 (N_29735,N_29349,N_29317);
xor U29736 (N_29736,N_29326,N_29477);
xnor U29737 (N_29737,N_29359,N_29257);
xor U29738 (N_29738,N_29390,N_29475);
and U29739 (N_29739,N_29444,N_29333);
nor U29740 (N_29740,N_29354,N_29450);
xor U29741 (N_29741,N_29394,N_29323);
xnor U29742 (N_29742,N_29353,N_29441);
xor U29743 (N_29743,N_29414,N_29467);
nand U29744 (N_29744,N_29308,N_29475);
nor U29745 (N_29745,N_29491,N_29318);
or U29746 (N_29746,N_29292,N_29388);
nor U29747 (N_29747,N_29350,N_29473);
or U29748 (N_29748,N_29328,N_29369);
nand U29749 (N_29749,N_29321,N_29272);
xor U29750 (N_29750,N_29722,N_29587);
nor U29751 (N_29751,N_29634,N_29504);
or U29752 (N_29752,N_29542,N_29683);
nor U29753 (N_29753,N_29738,N_29643);
and U29754 (N_29754,N_29729,N_29638);
xnor U29755 (N_29755,N_29655,N_29585);
and U29756 (N_29756,N_29582,N_29615);
and U29757 (N_29757,N_29574,N_29592);
xor U29758 (N_29758,N_29706,N_29691);
xnor U29759 (N_29759,N_29593,N_29690);
xnor U29760 (N_29760,N_29561,N_29700);
and U29761 (N_29761,N_29596,N_29598);
or U29762 (N_29762,N_29518,N_29631);
xor U29763 (N_29763,N_29676,N_29624);
xor U29764 (N_29764,N_29563,N_29679);
and U29765 (N_29765,N_29603,N_29703);
or U29766 (N_29766,N_29663,N_29580);
and U29767 (N_29767,N_29583,N_29550);
nor U29768 (N_29768,N_29526,N_29695);
nor U29769 (N_29769,N_29599,N_29726);
nor U29770 (N_29770,N_29567,N_29513);
and U29771 (N_29771,N_29537,N_29607);
xor U29772 (N_29772,N_29616,N_29736);
and U29773 (N_29773,N_29519,N_29648);
nand U29774 (N_29774,N_29571,N_29669);
and U29775 (N_29775,N_29512,N_29739);
nor U29776 (N_29776,N_29556,N_29613);
and U29777 (N_29777,N_29697,N_29584);
and U29778 (N_29778,N_29680,N_29650);
or U29779 (N_29779,N_29654,N_29621);
xnor U29780 (N_29780,N_29578,N_29713);
or U29781 (N_29781,N_29701,N_29731);
or U29782 (N_29782,N_29595,N_29741);
xnor U29783 (N_29783,N_29533,N_29590);
xor U29784 (N_29784,N_29649,N_29536);
nand U29785 (N_29785,N_29732,N_29678);
and U29786 (N_29786,N_29544,N_29594);
nand U29787 (N_29787,N_29558,N_29699);
or U29788 (N_29788,N_29619,N_29721);
and U29789 (N_29789,N_29562,N_29747);
nor U29790 (N_29790,N_29687,N_29605);
and U29791 (N_29791,N_29671,N_29517);
nor U29792 (N_29792,N_29646,N_29746);
xnor U29793 (N_29793,N_29627,N_29591);
or U29794 (N_29794,N_29659,N_29724);
or U29795 (N_29795,N_29626,N_29538);
nor U29796 (N_29796,N_29652,N_29610);
or U29797 (N_29797,N_29614,N_29718);
nor U29798 (N_29798,N_29532,N_29704);
and U29799 (N_29799,N_29508,N_29639);
and U29800 (N_29800,N_29712,N_29541);
nor U29801 (N_29801,N_29623,N_29633);
nand U29802 (N_29802,N_29743,N_29727);
or U29803 (N_29803,N_29682,N_29534);
xnor U29804 (N_29804,N_29716,N_29637);
nand U29805 (N_29805,N_29662,N_29719);
nor U29806 (N_29806,N_29546,N_29612);
nand U29807 (N_29807,N_29658,N_29507);
xnor U29808 (N_29808,N_29653,N_29503);
or U29809 (N_29809,N_29539,N_29730);
or U29810 (N_29810,N_29608,N_29674);
xnor U29811 (N_29811,N_29696,N_29566);
xnor U29812 (N_29812,N_29600,N_29501);
nor U29813 (N_29813,N_29636,N_29577);
or U29814 (N_29814,N_29656,N_29548);
or U29815 (N_29815,N_29640,N_29549);
or U29816 (N_29816,N_29715,N_29564);
nand U29817 (N_29817,N_29723,N_29557);
xor U29818 (N_29818,N_29688,N_29661);
nor U29819 (N_29819,N_29581,N_29728);
xnor U29820 (N_29820,N_29569,N_29510);
or U29821 (N_29821,N_29606,N_29515);
xor U29822 (N_29822,N_29657,N_29588);
nor U29823 (N_29823,N_29524,N_29622);
xnor U29824 (N_29824,N_29735,N_29745);
nor U29825 (N_29825,N_29714,N_29570);
xor U29826 (N_29826,N_29660,N_29673);
and U29827 (N_29827,N_29500,N_29672);
nor U29828 (N_29828,N_29547,N_29568);
nor U29829 (N_29829,N_29514,N_29529);
nand U29830 (N_29830,N_29651,N_29665);
nor U29831 (N_29831,N_29545,N_29520);
nand U29832 (N_29832,N_29744,N_29677);
and U29833 (N_29833,N_29565,N_29552);
nor U29834 (N_29834,N_29611,N_29628);
or U29835 (N_29835,N_29711,N_29632);
and U29836 (N_29836,N_29642,N_29685);
nand U29837 (N_29837,N_29670,N_29586);
nand U29838 (N_29838,N_29647,N_29681);
and U29839 (N_29839,N_29630,N_29551);
nor U29840 (N_29840,N_29625,N_29579);
nor U29841 (N_29841,N_29749,N_29693);
or U29842 (N_29842,N_29516,N_29528);
or U29843 (N_29843,N_29573,N_29531);
nand U29844 (N_29844,N_29609,N_29604);
or U29845 (N_29845,N_29527,N_29509);
nand U29846 (N_29846,N_29620,N_29692);
or U29847 (N_29847,N_29684,N_29530);
and U29848 (N_29848,N_29572,N_29748);
and U29849 (N_29849,N_29702,N_29686);
and U29850 (N_29850,N_29733,N_29720);
nor U29851 (N_29851,N_29725,N_29717);
nor U29852 (N_29852,N_29505,N_29559);
and U29853 (N_29853,N_29740,N_29602);
and U29854 (N_29854,N_29635,N_29575);
or U29855 (N_29855,N_29668,N_29707);
or U29856 (N_29856,N_29664,N_29553);
nand U29857 (N_29857,N_29737,N_29698);
and U29858 (N_29858,N_29523,N_29502);
xor U29859 (N_29859,N_29705,N_29666);
nand U29860 (N_29860,N_29589,N_29641);
nor U29861 (N_29861,N_29511,N_29540);
nand U29862 (N_29862,N_29554,N_29708);
xor U29863 (N_29863,N_29543,N_29597);
xnor U29864 (N_29864,N_29525,N_29522);
nor U29865 (N_29865,N_29601,N_29576);
or U29866 (N_29866,N_29734,N_29667);
xor U29867 (N_29867,N_29645,N_29675);
and U29868 (N_29868,N_29644,N_29689);
or U29869 (N_29869,N_29618,N_29617);
xnor U29870 (N_29870,N_29555,N_29629);
nand U29871 (N_29871,N_29521,N_29694);
xor U29872 (N_29872,N_29535,N_29560);
xor U29873 (N_29873,N_29710,N_29506);
xnor U29874 (N_29874,N_29742,N_29709);
nor U29875 (N_29875,N_29583,N_29605);
xnor U29876 (N_29876,N_29631,N_29513);
nor U29877 (N_29877,N_29670,N_29631);
or U29878 (N_29878,N_29505,N_29595);
and U29879 (N_29879,N_29730,N_29571);
nor U29880 (N_29880,N_29527,N_29670);
xnor U29881 (N_29881,N_29575,N_29722);
and U29882 (N_29882,N_29604,N_29613);
or U29883 (N_29883,N_29637,N_29602);
or U29884 (N_29884,N_29578,N_29513);
nand U29885 (N_29885,N_29550,N_29564);
or U29886 (N_29886,N_29661,N_29646);
xnor U29887 (N_29887,N_29585,N_29725);
nor U29888 (N_29888,N_29599,N_29713);
or U29889 (N_29889,N_29601,N_29589);
xnor U29890 (N_29890,N_29748,N_29596);
nor U29891 (N_29891,N_29661,N_29719);
nand U29892 (N_29892,N_29678,N_29680);
xor U29893 (N_29893,N_29623,N_29732);
nor U29894 (N_29894,N_29738,N_29648);
xor U29895 (N_29895,N_29661,N_29622);
xnor U29896 (N_29896,N_29654,N_29709);
nor U29897 (N_29897,N_29526,N_29684);
xor U29898 (N_29898,N_29653,N_29587);
xor U29899 (N_29899,N_29621,N_29715);
xnor U29900 (N_29900,N_29583,N_29699);
or U29901 (N_29901,N_29691,N_29740);
xnor U29902 (N_29902,N_29610,N_29589);
nor U29903 (N_29903,N_29716,N_29502);
nand U29904 (N_29904,N_29708,N_29721);
nand U29905 (N_29905,N_29550,N_29715);
nand U29906 (N_29906,N_29747,N_29661);
xor U29907 (N_29907,N_29705,N_29672);
or U29908 (N_29908,N_29697,N_29665);
xnor U29909 (N_29909,N_29516,N_29733);
and U29910 (N_29910,N_29556,N_29510);
nor U29911 (N_29911,N_29734,N_29722);
or U29912 (N_29912,N_29721,N_29620);
nor U29913 (N_29913,N_29510,N_29531);
or U29914 (N_29914,N_29674,N_29543);
or U29915 (N_29915,N_29681,N_29640);
nor U29916 (N_29916,N_29523,N_29710);
or U29917 (N_29917,N_29505,N_29552);
and U29918 (N_29918,N_29748,N_29736);
nand U29919 (N_29919,N_29713,N_29715);
xor U29920 (N_29920,N_29641,N_29676);
nor U29921 (N_29921,N_29705,N_29634);
and U29922 (N_29922,N_29672,N_29612);
nor U29923 (N_29923,N_29735,N_29696);
nor U29924 (N_29924,N_29577,N_29665);
or U29925 (N_29925,N_29612,N_29507);
nor U29926 (N_29926,N_29688,N_29562);
or U29927 (N_29927,N_29676,N_29630);
nand U29928 (N_29928,N_29604,N_29709);
xor U29929 (N_29929,N_29717,N_29599);
or U29930 (N_29930,N_29599,N_29715);
nand U29931 (N_29931,N_29518,N_29656);
nand U29932 (N_29932,N_29643,N_29669);
nand U29933 (N_29933,N_29709,N_29744);
xnor U29934 (N_29934,N_29615,N_29543);
nor U29935 (N_29935,N_29513,N_29549);
nand U29936 (N_29936,N_29623,N_29577);
and U29937 (N_29937,N_29740,N_29510);
and U29938 (N_29938,N_29585,N_29584);
nor U29939 (N_29939,N_29718,N_29601);
and U29940 (N_29940,N_29564,N_29649);
and U29941 (N_29941,N_29697,N_29708);
nor U29942 (N_29942,N_29548,N_29726);
nor U29943 (N_29943,N_29731,N_29578);
nor U29944 (N_29944,N_29676,N_29606);
xor U29945 (N_29945,N_29521,N_29616);
xnor U29946 (N_29946,N_29711,N_29634);
nor U29947 (N_29947,N_29684,N_29642);
or U29948 (N_29948,N_29596,N_29530);
nand U29949 (N_29949,N_29543,N_29539);
and U29950 (N_29950,N_29711,N_29510);
or U29951 (N_29951,N_29578,N_29541);
nand U29952 (N_29952,N_29629,N_29721);
xnor U29953 (N_29953,N_29724,N_29537);
xnor U29954 (N_29954,N_29736,N_29738);
or U29955 (N_29955,N_29524,N_29666);
xor U29956 (N_29956,N_29568,N_29675);
xor U29957 (N_29957,N_29594,N_29639);
nand U29958 (N_29958,N_29590,N_29723);
nor U29959 (N_29959,N_29699,N_29636);
and U29960 (N_29960,N_29735,N_29730);
nor U29961 (N_29961,N_29530,N_29652);
and U29962 (N_29962,N_29530,N_29547);
or U29963 (N_29963,N_29585,N_29529);
or U29964 (N_29964,N_29634,N_29540);
xor U29965 (N_29965,N_29691,N_29634);
nand U29966 (N_29966,N_29651,N_29658);
and U29967 (N_29967,N_29650,N_29526);
xor U29968 (N_29968,N_29675,N_29692);
xor U29969 (N_29969,N_29746,N_29538);
nand U29970 (N_29970,N_29702,N_29717);
nand U29971 (N_29971,N_29512,N_29684);
nand U29972 (N_29972,N_29670,N_29552);
nor U29973 (N_29973,N_29715,N_29744);
or U29974 (N_29974,N_29699,N_29709);
and U29975 (N_29975,N_29523,N_29723);
and U29976 (N_29976,N_29620,N_29707);
or U29977 (N_29977,N_29605,N_29659);
xnor U29978 (N_29978,N_29527,N_29743);
or U29979 (N_29979,N_29543,N_29733);
and U29980 (N_29980,N_29731,N_29573);
xnor U29981 (N_29981,N_29614,N_29739);
xor U29982 (N_29982,N_29504,N_29521);
xnor U29983 (N_29983,N_29504,N_29732);
and U29984 (N_29984,N_29641,N_29682);
xnor U29985 (N_29985,N_29647,N_29622);
or U29986 (N_29986,N_29536,N_29681);
nor U29987 (N_29987,N_29630,N_29531);
and U29988 (N_29988,N_29507,N_29649);
nand U29989 (N_29989,N_29526,N_29657);
and U29990 (N_29990,N_29618,N_29530);
or U29991 (N_29991,N_29539,N_29542);
or U29992 (N_29992,N_29652,N_29654);
or U29993 (N_29993,N_29705,N_29712);
nand U29994 (N_29994,N_29551,N_29545);
nand U29995 (N_29995,N_29504,N_29567);
nor U29996 (N_29996,N_29636,N_29525);
or U29997 (N_29997,N_29622,N_29554);
and U29998 (N_29998,N_29610,N_29530);
and U29999 (N_29999,N_29569,N_29736);
nor U30000 (N_30000,N_29772,N_29759);
xor U30001 (N_30001,N_29837,N_29815);
nor U30002 (N_30002,N_29895,N_29765);
and U30003 (N_30003,N_29926,N_29891);
nand U30004 (N_30004,N_29954,N_29885);
nor U30005 (N_30005,N_29915,N_29822);
nand U30006 (N_30006,N_29816,N_29857);
and U30007 (N_30007,N_29909,N_29861);
nor U30008 (N_30008,N_29862,N_29897);
and U30009 (N_30009,N_29940,N_29876);
nor U30010 (N_30010,N_29943,N_29997);
nand U30011 (N_30011,N_29889,N_29786);
xnor U30012 (N_30012,N_29869,N_29824);
nor U30013 (N_30013,N_29910,N_29911);
xnor U30014 (N_30014,N_29965,N_29966);
nor U30015 (N_30015,N_29963,N_29987);
xor U30016 (N_30016,N_29769,N_29797);
nand U30017 (N_30017,N_29778,N_29863);
and U30018 (N_30018,N_29962,N_29764);
nor U30019 (N_30019,N_29931,N_29901);
or U30020 (N_30020,N_29848,N_29866);
nand U30021 (N_30021,N_29974,N_29828);
xnor U30022 (N_30022,N_29917,N_29920);
and U30023 (N_30023,N_29996,N_29750);
or U30024 (N_30024,N_29957,N_29827);
xor U30025 (N_30025,N_29930,N_29896);
nand U30026 (N_30026,N_29975,N_29958);
or U30027 (N_30027,N_29875,N_29913);
xnor U30028 (N_30028,N_29807,N_29880);
and U30029 (N_30029,N_29798,N_29868);
nand U30030 (N_30030,N_29884,N_29841);
nor U30031 (N_30031,N_29933,N_29960);
nand U30032 (N_30032,N_29938,N_29886);
nand U30033 (N_30033,N_29903,N_29919);
nand U30034 (N_30034,N_29838,N_29927);
or U30035 (N_30035,N_29937,N_29916);
nor U30036 (N_30036,N_29834,N_29760);
and U30037 (N_30037,N_29792,N_29860);
nor U30038 (N_30038,N_29844,N_29936);
and U30039 (N_30039,N_29979,N_29755);
nand U30040 (N_30040,N_29887,N_29907);
and U30041 (N_30041,N_29809,N_29766);
nor U30042 (N_30042,N_29808,N_29758);
xnor U30043 (N_30043,N_29795,N_29984);
or U30044 (N_30044,N_29802,N_29825);
and U30045 (N_30045,N_29817,N_29977);
and U30046 (N_30046,N_29770,N_29780);
xnor U30047 (N_30047,N_29908,N_29925);
nor U30048 (N_30048,N_29900,N_29971);
xor U30049 (N_30049,N_29973,N_29921);
or U30050 (N_30050,N_29964,N_29843);
nand U30051 (N_30051,N_29976,N_29883);
xnor U30052 (N_30052,N_29835,N_29773);
or U30053 (N_30053,N_29830,N_29948);
or U30054 (N_30054,N_29801,N_29810);
and U30055 (N_30055,N_29912,N_29849);
and U30056 (N_30056,N_29774,N_29946);
xnor U30057 (N_30057,N_29864,N_29820);
nor U30058 (N_30058,N_29782,N_29829);
or U30059 (N_30059,N_29893,N_29767);
nor U30060 (N_30060,N_29871,N_29995);
nand U30061 (N_30061,N_29804,N_29942);
nor U30062 (N_30062,N_29776,N_29836);
and U30063 (N_30063,N_29865,N_29986);
xor U30064 (N_30064,N_29941,N_29847);
xnor U30065 (N_30065,N_29981,N_29929);
nor U30066 (N_30066,N_29881,N_29842);
or U30067 (N_30067,N_29888,N_29821);
or U30068 (N_30068,N_29906,N_29856);
nand U30069 (N_30069,N_29793,N_29879);
and U30070 (N_30070,N_29787,N_29935);
nor U30071 (N_30071,N_29831,N_29819);
and U30072 (N_30072,N_29784,N_29813);
nor U30073 (N_30073,N_29763,N_29854);
and U30074 (N_30074,N_29999,N_29989);
nor U30075 (N_30075,N_29753,N_29898);
nor U30076 (N_30076,N_29811,N_29994);
nand U30077 (N_30077,N_29902,N_29823);
and U30078 (N_30078,N_29923,N_29761);
nand U30079 (N_30079,N_29762,N_29968);
xor U30080 (N_30080,N_29882,N_29991);
nor U30081 (N_30081,N_29905,N_29928);
xor U30082 (N_30082,N_29990,N_29833);
xor U30083 (N_30083,N_29771,N_29982);
nor U30084 (N_30084,N_29805,N_29945);
xor U30085 (N_30085,N_29947,N_29873);
nor U30086 (N_30086,N_29877,N_29794);
nand U30087 (N_30087,N_29799,N_29899);
xnor U30088 (N_30088,N_29939,N_29754);
and U30089 (N_30089,N_29949,N_29988);
and U30090 (N_30090,N_29790,N_29972);
xor U30091 (N_30091,N_29992,N_29914);
and U30092 (N_30092,N_29918,N_29785);
xor U30093 (N_30093,N_29969,N_29852);
xnor U30094 (N_30094,N_29956,N_29924);
or U30095 (N_30095,N_29985,N_29845);
or U30096 (N_30096,N_29840,N_29832);
nand U30097 (N_30097,N_29789,N_29783);
xnor U30098 (N_30098,N_29967,N_29993);
or U30099 (N_30099,N_29955,N_29850);
nor U30100 (N_30100,N_29777,N_29998);
xor U30101 (N_30101,N_29892,N_29814);
nor U30102 (N_30102,N_29768,N_29751);
or U30103 (N_30103,N_29800,N_29894);
and U30104 (N_30104,N_29779,N_29978);
xor U30105 (N_30105,N_29878,N_29961);
xor U30106 (N_30106,N_29781,N_29970);
or U30107 (N_30107,N_29846,N_29952);
xor U30108 (N_30108,N_29757,N_29904);
or U30109 (N_30109,N_29796,N_29752);
nand U30110 (N_30110,N_29775,N_29855);
and U30111 (N_30111,N_29791,N_29953);
and U30112 (N_30112,N_29870,N_29803);
and U30113 (N_30113,N_29853,N_29867);
nand U30114 (N_30114,N_29818,N_29980);
nor U30115 (N_30115,N_29890,N_29872);
nor U30116 (N_30116,N_29806,N_29983);
nor U30117 (N_30117,N_29826,N_29922);
and U30118 (N_30118,N_29788,N_29839);
and U30119 (N_30119,N_29874,N_29756);
and U30120 (N_30120,N_29812,N_29959);
nand U30121 (N_30121,N_29859,N_29851);
nand U30122 (N_30122,N_29934,N_29932);
nor U30123 (N_30123,N_29944,N_29950);
nand U30124 (N_30124,N_29951,N_29858);
or U30125 (N_30125,N_29910,N_29924);
nor U30126 (N_30126,N_29964,N_29793);
and U30127 (N_30127,N_29939,N_29813);
nand U30128 (N_30128,N_29765,N_29932);
nand U30129 (N_30129,N_29931,N_29976);
and U30130 (N_30130,N_29915,N_29770);
or U30131 (N_30131,N_29797,N_29955);
xor U30132 (N_30132,N_29813,N_29974);
nor U30133 (N_30133,N_29794,N_29780);
and U30134 (N_30134,N_29875,N_29901);
nand U30135 (N_30135,N_29780,N_29855);
or U30136 (N_30136,N_29800,N_29864);
or U30137 (N_30137,N_29762,N_29924);
or U30138 (N_30138,N_29940,N_29944);
and U30139 (N_30139,N_29935,N_29821);
xor U30140 (N_30140,N_29940,N_29803);
or U30141 (N_30141,N_29781,N_29928);
nand U30142 (N_30142,N_29947,N_29991);
xor U30143 (N_30143,N_29969,N_29894);
nand U30144 (N_30144,N_29910,N_29976);
nor U30145 (N_30145,N_29880,N_29874);
or U30146 (N_30146,N_29991,N_29822);
xnor U30147 (N_30147,N_29814,N_29801);
xnor U30148 (N_30148,N_29990,N_29920);
xnor U30149 (N_30149,N_29868,N_29946);
xor U30150 (N_30150,N_29951,N_29886);
or U30151 (N_30151,N_29771,N_29966);
xor U30152 (N_30152,N_29779,N_29754);
nor U30153 (N_30153,N_29751,N_29916);
nor U30154 (N_30154,N_29962,N_29814);
nor U30155 (N_30155,N_29991,N_29970);
nor U30156 (N_30156,N_29771,N_29905);
and U30157 (N_30157,N_29838,N_29824);
or U30158 (N_30158,N_29918,N_29872);
nor U30159 (N_30159,N_29759,N_29986);
nor U30160 (N_30160,N_29836,N_29866);
xnor U30161 (N_30161,N_29891,N_29918);
and U30162 (N_30162,N_29926,N_29956);
or U30163 (N_30163,N_29767,N_29863);
or U30164 (N_30164,N_29932,N_29953);
nor U30165 (N_30165,N_29829,N_29933);
or U30166 (N_30166,N_29801,N_29796);
or U30167 (N_30167,N_29952,N_29776);
or U30168 (N_30168,N_29976,N_29943);
and U30169 (N_30169,N_29896,N_29883);
xor U30170 (N_30170,N_29984,N_29820);
nand U30171 (N_30171,N_29963,N_29841);
and U30172 (N_30172,N_29919,N_29758);
and U30173 (N_30173,N_29762,N_29783);
or U30174 (N_30174,N_29956,N_29992);
xor U30175 (N_30175,N_29872,N_29844);
and U30176 (N_30176,N_29911,N_29899);
and U30177 (N_30177,N_29911,N_29859);
nand U30178 (N_30178,N_29954,N_29806);
xor U30179 (N_30179,N_29992,N_29857);
and U30180 (N_30180,N_29933,N_29861);
or U30181 (N_30181,N_29893,N_29774);
nor U30182 (N_30182,N_29921,N_29861);
nor U30183 (N_30183,N_29756,N_29900);
nor U30184 (N_30184,N_29884,N_29878);
and U30185 (N_30185,N_29763,N_29852);
and U30186 (N_30186,N_29833,N_29830);
nor U30187 (N_30187,N_29950,N_29887);
nor U30188 (N_30188,N_29818,N_29784);
nand U30189 (N_30189,N_29945,N_29934);
nor U30190 (N_30190,N_29790,N_29884);
nor U30191 (N_30191,N_29913,N_29885);
nor U30192 (N_30192,N_29934,N_29821);
and U30193 (N_30193,N_29774,N_29903);
nor U30194 (N_30194,N_29882,N_29811);
nor U30195 (N_30195,N_29892,N_29996);
nand U30196 (N_30196,N_29799,N_29832);
nor U30197 (N_30197,N_29842,N_29814);
nand U30198 (N_30198,N_29876,N_29822);
nand U30199 (N_30199,N_29938,N_29937);
or U30200 (N_30200,N_29819,N_29798);
or U30201 (N_30201,N_29997,N_29908);
and U30202 (N_30202,N_29758,N_29795);
xnor U30203 (N_30203,N_29777,N_29783);
and U30204 (N_30204,N_29877,N_29791);
or U30205 (N_30205,N_29851,N_29832);
and U30206 (N_30206,N_29793,N_29821);
nor U30207 (N_30207,N_29950,N_29959);
xor U30208 (N_30208,N_29816,N_29942);
nand U30209 (N_30209,N_29895,N_29762);
or U30210 (N_30210,N_29780,N_29799);
or U30211 (N_30211,N_29958,N_29842);
or U30212 (N_30212,N_29867,N_29849);
or U30213 (N_30213,N_29904,N_29814);
and U30214 (N_30214,N_29839,N_29863);
nor U30215 (N_30215,N_29800,N_29765);
nand U30216 (N_30216,N_29776,N_29800);
nor U30217 (N_30217,N_29988,N_29910);
xor U30218 (N_30218,N_29780,N_29789);
nor U30219 (N_30219,N_29961,N_29992);
and U30220 (N_30220,N_29832,N_29830);
or U30221 (N_30221,N_29862,N_29873);
nor U30222 (N_30222,N_29956,N_29873);
nor U30223 (N_30223,N_29783,N_29888);
nand U30224 (N_30224,N_29919,N_29871);
xnor U30225 (N_30225,N_29936,N_29890);
or U30226 (N_30226,N_29967,N_29839);
xnor U30227 (N_30227,N_29813,N_29835);
and U30228 (N_30228,N_29835,N_29981);
nor U30229 (N_30229,N_29807,N_29982);
nand U30230 (N_30230,N_29864,N_29964);
or U30231 (N_30231,N_29860,N_29867);
nand U30232 (N_30232,N_29758,N_29857);
xor U30233 (N_30233,N_29947,N_29850);
and U30234 (N_30234,N_29885,N_29824);
xnor U30235 (N_30235,N_29941,N_29780);
or U30236 (N_30236,N_29761,N_29929);
or U30237 (N_30237,N_29809,N_29836);
xor U30238 (N_30238,N_29991,N_29799);
nand U30239 (N_30239,N_29934,N_29908);
and U30240 (N_30240,N_29753,N_29947);
xnor U30241 (N_30241,N_29837,N_29904);
and U30242 (N_30242,N_29987,N_29788);
and U30243 (N_30243,N_29876,N_29834);
or U30244 (N_30244,N_29812,N_29774);
nand U30245 (N_30245,N_29942,N_29974);
and U30246 (N_30246,N_29944,N_29946);
xor U30247 (N_30247,N_29938,N_29966);
nor U30248 (N_30248,N_29775,N_29947);
or U30249 (N_30249,N_29861,N_29811);
and U30250 (N_30250,N_30211,N_30055);
nand U30251 (N_30251,N_30185,N_30130);
or U30252 (N_30252,N_30120,N_30115);
nor U30253 (N_30253,N_30000,N_30033);
and U30254 (N_30254,N_30192,N_30140);
or U30255 (N_30255,N_30020,N_30005);
or U30256 (N_30256,N_30056,N_30248);
or U30257 (N_30257,N_30219,N_30008);
nor U30258 (N_30258,N_30068,N_30046);
xor U30259 (N_30259,N_30154,N_30016);
and U30260 (N_30260,N_30070,N_30222);
and U30261 (N_30261,N_30039,N_30143);
and U30262 (N_30262,N_30190,N_30137);
nand U30263 (N_30263,N_30009,N_30221);
nand U30264 (N_30264,N_30026,N_30158);
or U30265 (N_30265,N_30196,N_30215);
nor U30266 (N_30266,N_30231,N_30146);
xnor U30267 (N_30267,N_30091,N_30133);
xnor U30268 (N_30268,N_30167,N_30142);
xnor U30269 (N_30269,N_30060,N_30191);
and U30270 (N_30270,N_30187,N_30225);
nor U30271 (N_30271,N_30013,N_30004);
nor U30272 (N_30272,N_30012,N_30122);
and U30273 (N_30273,N_30199,N_30245);
nor U30274 (N_30274,N_30031,N_30178);
and U30275 (N_30275,N_30049,N_30010);
or U30276 (N_30276,N_30123,N_30236);
nand U30277 (N_30277,N_30220,N_30007);
xor U30278 (N_30278,N_30134,N_30181);
nand U30279 (N_30279,N_30200,N_30213);
nand U30280 (N_30280,N_30080,N_30088);
or U30281 (N_30281,N_30112,N_30011);
nor U30282 (N_30282,N_30223,N_30081);
nand U30283 (N_30283,N_30125,N_30210);
or U30284 (N_30284,N_30038,N_30212);
nand U30285 (N_30285,N_30179,N_30239);
nor U30286 (N_30286,N_30157,N_30066);
and U30287 (N_30287,N_30111,N_30232);
xnor U30288 (N_30288,N_30205,N_30052);
and U30289 (N_30289,N_30147,N_30144);
xnor U30290 (N_30290,N_30131,N_30023);
or U30291 (N_30291,N_30092,N_30006);
or U30292 (N_30292,N_30103,N_30109);
or U30293 (N_30293,N_30022,N_30107);
or U30294 (N_30294,N_30160,N_30098);
or U30295 (N_30295,N_30176,N_30214);
nor U30296 (N_30296,N_30030,N_30128);
and U30297 (N_30297,N_30175,N_30044);
nand U30298 (N_30298,N_30047,N_30036);
nand U30299 (N_30299,N_30201,N_30186);
or U30300 (N_30300,N_30065,N_30105);
nand U30301 (N_30301,N_30209,N_30169);
nand U30302 (N_30302,N_30099,N_30184);
and U30303 (N_30303,N_30193,N_30182);
and U30304 (N_30304,N_30230,N_30249);
nand U30305 (N_30305,N_30173,N_30108);
and U30306 (N_30306,N_30162,N_30048);
or U30307 (N_30307,N_30207,N_30101);
xnor U30308 (N_30308,N_30166,N_30024);
nor U30309 (N_30309,N_30089,N_30235);
nor U30310 (N_30310,N_30136,N_30233);
xnor U30311 (N_30311,N_30029,N_30145);
nand U30312 (N_30312,N_30096,N_30014);
nand U30313 (N_30313,N_30238,N_30153);
nor U30314 (N_30314,N_30085,N_30135);
and U30315 (N_30315,N_30204,N_30246);
and U30316 (N_30316,N_30077,N_30102);
xnor U30317 (N_30317,N_30206,N_30198);
and U30318 (N_30318,N_30124,N_30054);
and U30319 (N_30319,N_30119,N_30063);
nand U30320 (N_30320,N_30188,N_30003);
nand U30321 (N_30321,N_30218,N_30171);
xnor U30322 (N_30322,N_30161,N_30095);
and U30323 (N_30323,N_30094,N_30129);
nor U30324 (N_30324,N_30229,N_30069);
and U30325 (N_30325,N_30168,N_30164);
or U30326 (N_30326,N_30138,N_30126);
and U30327 (N_30327,N_30180,N_30165);
xor U30328 (N_30328,N_30035,N_30072);
nor U30329 (N_30329,N_30104,N_30139);
or U30330 (N_30330,N_30058,N_30183);
nor U30331 (N_30331,N_30018,N_30032);
and U30332 (N_30332,N_30019,N_30045);
nand U30333 (N_30333,N_30106,N_30244);
nand U30334 (N_30334,N_30028,N_30127);
or U30335 (N_30335,N_30148,N_30237);
or U30336 (N_30336,N_30062,N_30226);
nand U30337 (N_30337,N_30110,N_30202);
or U30338 (N_30338,N_30240,N_30057);
xor U30339 (N_30339,N_30170,N_30017);
and U30340 (N_30340,N_30041,N_30216);
xor U30341 (N_30341,N_30097,N_30079);
and U30342 (N_30342,N_30243,N_30197);
and U30343 (N_30343,N_30224,N_30163);
xor U30344 (N_30344,N_30040,N_30189);
nand U30345 (N_30345,N_30076,N_30172);
nand U30346 (N_30346,N_30093,N_30247);
xor U30347 (N_30347,N_30050,N_30121);
nor U30348 (N_30348,N_30234,N_30087);
and U30349 (N_30349,N_30150,N_30071);
nor U30350 (N_30350,N_30151,N_30042);
nand U30351 (N_30351,N_30116,N_30113);
xor U30352 (N_30352,N_30132,N_30053);
or U30353 (N_30353,N_30059,N_30195);
nand U30354 (N_30354,N_30067,N_30217);
nor U30355 (N_30355,N_30001,N_30082);
nand U30356 (N_30356,N_30086,N_30002);
nand U30357 (N_30357,N_30037,N_30015);
nand U30358 (N_30358,N_30078,N_30156);
and U30359 (N_30359,N_30025,N_30064);
nand U30360 (N_30360,N_30155,N_30149);
or U30361 (N_30361,N_30100,N_30027);
xnor U30362 (N_30362,N_30075,N_30174);
xnor U30363 (N_30363,N_30177,N_30073);
nor U30364 (N_30364,N_30034,N_30241);
xnor U30365 (N_30365,N_30203,N_30141);
and U30366 (N_30366,N_30061,N_30194);
nor U30367 (N_30367,N_30152,N_30208);
xnor U30368 (N_30368,N_30043,N_30242);
and U30369 (N_30369,N_30051,N_30084);
and U30370 (N_30370,N_30074,N_30228);
xnor U30371 (N_30371,N_30117,N_30114);
and U30372 (N_30372,N_30083,N_30090);
xnor U30373 (N_30373,N_30021,N_30159);
xor U30374 (N_30374,N_30118,N_30227);
xor U30375 (N_30375,N_30046,N_30157);
and U30376 (N_30376,N_30198,N_30142);
xnor U30377 (N_30377,N_30040,N_30215);
xor U30378 (N_30378,N_30238,N_30161);
nand U30379 (N_30379,N_30077,N_30113);
or U30380 (N_30380,N_30193,N_30003);
and U30381 (N_30381,N_30070,N_30246);
and U30382 (N_30382,N_30182,N_30122);
xnor U30383 (N_30383,N_30165,N_30022);
and U30384 (N_30384,N_30222,N_30111);
nor U30385 (N_30385,N_30069,N_30243);
or U30386 (N_30386,N_30103,N_30243);
xor U30387 (N_30387,N_30051,N_30221);
nand U30388 (N_30388,N_30085,N_30065);
and U30389 (N_30389,N_30022,N_30228);
xor U30390 (N_30390,N_30105,N_30190);
nor U30391 (N_30391,N_30034,N_30172);
nor U30392 (N_30392,N_30043,N_30118);
xnor U30393 (N_30393,N_30007,N_30115);
and U30394 (N_30394,N_30043,N_30055);
nor U30395 (N_30395,N_30002,N_30231);
and U30396 (N_30396,N_30191,N_30086);
nand U30397 (N_30397,N_30164,N_30206);
nand U30398 (N_30398,N_30008,N_30116);
and U30399 (N_30399,N_30089,N_30071);
nor U30400 (N_30400,N_30030,N_30182);
xnor U30401 (N_30401,N_30222,N_30036);
nand U30402 (N_30402,N_30209,N_30130);
nor U30403 (N_30403,N_30176,N_30014);
and U30404 (N_30404,N_30249,N_30186);
xnor U30405 (N_30405,N_30093,N_30241);
xnor U30406 (N_30406,N_30182,N_30018);
or U30407 (N_30407,N_30211,N_30093);
and U30408 (N_30408,N_30013,N_30093);
xnor U30409 (N_30409,N_30072,N_30198);
and U30410 (N_30410,N_30017,N_30198);
nand U30411 (N_30411,N_30187,N_30027);
or U30412 (N_30412,N_30021,N_30132);
xor U30413 (N_30413,N_30201,N_30075);
nand U30414 (N_30414,N_30106,N_30047);
xor U30415 (N_30415,N_30170,N_30162);
nand U30416 (N_30416,N_30029,N_30215);
nand U30417 (N_30417,N_30201,N_30030);
nand U30418 (N_30418,N_30084,N_30119);
and U30419 (N_30419,N_30180,N_30109);
nand U30420 (N_30420,N_30180,N_30114);
nor U30421 (N_30421,N_30238,N_30241);
xor U30422 (N_30422,N_30164,N_30228);
nor U30423 (N_30423,N_30227,N_30197);
nor U30424 (N_30424,N_30213,N_30105);
and U30425 (N_30425,N_30132,N_30015);
and U30426 (N_30426,N_30249,N_30218);
nor U30427 (N_30427,N_30088,N_30043);
nand U30428 (N_30428,N_30047,N_30151);
nor U30429 (N_30429,N_30001,N_30000);
nand U30430 (N_30430,N_30244,N_30194);
and U30431 (N_30431,N_30136,N_30145);
and U30432 (N_30432,N_30064,N_30054);
xor U30433 (N_30433,N_30247,N_30050);
nand U30434 (N_30434,N_30207,N_30190);
and U30435 (N_30435,N_30057,N_30031);
or U30436 (N_30436,N_30188,N_30161);
and U30437 (N_30437,N_30148,N_30144);
xnor U30438 (N_30438,N_30047,N_30037);
or U30439 (N_30439,N_30212,N_30111);
xor U30440 (N_30440,N_30168,N_30047);
and U30441 (N_30441,N_30015,N_30055);
or U30442 (N_30442,N_30137,N_30107);
or U30443 (N_30443,N_30135,N_30195);
xnor U30444 (N_30444,N_30122,N_30070);
or U30445 (N_30445,N_30068,N_30143);
and U30446 (N_30446,N_30073,N_30235);
xor U30447 (N_30447,N_30223,N_30107);
and U30448 (N_30448,N_30179,N_30103);
or U30449 (N_30449,N_30203,N_30031);
nor U30450 (N_30450,N_30062,N_30129);
nor U30451 (N_30451,N_30179,N_30119);
xor U30452 (N_30452,N_30167,N_30043);
and U30453 (N_30453,N_30208,N_30141);
nand U30454 (N_30454,N_30239,N_30094);
nor U30455 (N_30455,N_30143,N_30244);
xor U30456 (N_30456,N_30078,N_30013);
xor U30457 (N_30457,N_30179,N_30046);
and U30458 (N_30458,N_30034,N_30068);
xnor U30459 (N_30459,N_30049,N_30105);
xnor U30460 (N_30460,N_30017,N_30201);
xnor U30461 (N_30461,N_30135,N_30152);
and U30462 (N_30462,N_30173,N_30166);
xnor U30463 (N_30463,N_30178,N_30119);
nand U30464 (N_30464,N_30139,N_30217);
nand U30465 (N_30465,N_30072,N_30163);
nand U30466 (N_30466,N_30152,N_30138);
xor U30467 (N_30467,N_30242,N_30151);
nor U30468 (N_30468,N_30075,N_30074);
or U30469 (N_30469,N_30071,N_30218);
xnor U30470 (N_30470,N_30153,N_30087);
xor U30471 (N_30471,N_30069,N_30044);
and U30472 (N_30472,N_30230,N_30058);
nor U30473 (N_30473,N_30042,N_30160);
and U30474 (N_30474,N_30085,N_30222);
nor U30475 (N_30475,N_30151,N_30119);
nand U30476 (N_30476,N_30067,N_30113);
or U30477 (N_30477,N_30060,N_30193);
nor U30478 (N_30478,N_30109,N_30185);
nor U30479 (N_30479,N_30227,N_30138);
or U30480 (N_30480,N_30198,N_30153);
xor U30481 (N_30481,N_30001,N_30095);
nand U30482 (N_30482,N_30240,N_30018);
or U30483 (N_30483,N_30041,N_30148);
nor U30484 (N_30484,N_30124,N_30059);
or U30485 (N_30485,N_30083,N_30206);
and U30486 (N_30486,N_30126,N_30025);
nor U30487 (N_30487,N_30139,N_30211);
and U30488 (N_30488,N_30039,N_30053);
xor U30489 (N_30489,N_30208,N_30160);
nor U30490 (N_30490,N_30041,N_30036);
xnor U30491 (N_30491,N_30190,N_30092);
xor U30492 (N_30492,N_30138,N_30217);
or U30493 (N_30493,N_30084,N_30126);
xor U30494 (N_30494,N_30210,N_30039);
nand U30495 (N_30495,N_30021,N_30074);
and U30496 (N_30496,N_30070,N_30128);
xor U30497 (N_30497,N_30137,N_30192);
nor U30498 (N_30498,N_30159,N_30240);
or U30499 (N_30499,N_30002,N_30220);
nor U30500 (N_30500,N_30274,N_30412);
xor U30501 (N_30501,N_30260,N_30476);
and U30502 (N_30502,N_30268,N_30487);
xor U30503 (N_30503,N_30266,N_30416);
nand U30504 (N_30504,N_30371,N_30373);
nor U30505 (N_30505,N_30300,N_30454);
xnor U30506 (N_30506,N_30491,N_30307);
or U30507 (N_30507,N_30286,N_30308);
nor U30508 (N_30508,N_30409,N_30346);
and U30509 (N_30509,N_30320,N_30343);
and U30510 (N_30510,N_30313,N_30348);
and U30511 (N_30511,N_30361,N_30332);
and U30512 (N_30512,N_30468,N_30380);
xnor U30513 (N_30513,N_30276,N_30338);
nor U30514 (N_30514,N_30334,N_30292);
or U30515 (N_30515,N_30422,N_30493);
nand U30516 (N_30516,N_30404,N_30426);
or U30517 (N_30517,N_30494,N_30317);
or U30518 (N_30518,N_30467,N_30269);
nand U30519 (N_30519,N_30324,N_30363);
xnor U30520 (N_30520,N_30263,N_30367);
nor U30521 (N_30521,N_30377,N_30295);
or U30522 (N_30522,N_30403,N_30273);
nand U30523 (N_30523,N_30433,N_30424);
nand U30524 (N_30524,N_30453,N_30462);
nor U30525 (N_30525,N_30452,N_30392);
nor U30526 (N_30526,N_30482,N_30279);
nand U30527 (N_30527,N_30470,N_30486);
xor U30528 (N_30528,N_30396,N_30285);
or U30529 (N_30529,N_30407,N_30335);
or U30530 (N_30530,N_30459,N_30379);
nor U30531 (N_30531,N_30288,N_30417);
and U30532 (N_30532,N_30496,N_30302);
xor U30533 (N_30533,N_30387,N_30289);
or U30534 (N_30534,N_30419,N_30305);
nor U30535 (N_30535,N_30441,N_30333);
xnor U30536 (N_30536,N_30410,N_30431);
nand U30537 (N_30537,N_30388,N_30329);
and U30538 (N_30538,N_30282,N_30397);
or U30539 (N_30539,N_30341,N_30378);
xor U30540 (N_30540,N_30314,N_30303);
nor U30541 (N_30541,N_30406,N_30429);
or U30542 (N_30542,N_30370,N_30366);
and U30543 (N_30543,N_30306,N_30258);
and U30544 (N_30544,N_30278,N_30428);
or U30545 (N_30545,N_30349,N_30290);
nor U30546 (N_30546,N_30461,N_30298);
xnor U30547 (N_30547,N_30336,N_30451);
xor U30548 (N_30548,N_30294,N_30345);
xnor U30549 (N_30549,N_30430,N_30492);
nor U30550 (N_30550,N_30434,N_30411);
or U30551 (N_30551,N_30251,N_30259);
nand U30552 (N_30552,N_30400,N_30497);
xor U30553 (N_30553,N_30472,N_30479);
xor U30554 (N_30554,N_30254,N_30483);
nand U30555 (N_30555,N_30331,N_30287);
nor U30556 (N_30556,N_30337,N_30464);
and U30557 (N_30557,N_30401,N_30484);
nor U30558 (N_30558,N_30339,N_30393);
or U30559 (N_30559,N_30425,N_30421);
and U30560 (N_30560,N_30359,N_30374);
xor U30561 (N_30561,N_30382,N_30304);
and U30562 (N_30562,N_30437,N_30385);
and U30563 (N_30563,N_30328,N_30267);
and U30564 (N_30564,N_30321,N_30465);
and U30565 (N_30565,N_30384,N_30443);
xnor U30566 (N_30566,N_30394,N_30347);
or U30567 (N_30567,N_30466,N_30478);
nor U30568 (N_30568,N_30275,N_30488);
or U30569 (N_30569,N_30365,N_30391);
nor U30570 (N_30570,N_30499,N_30398);
xnor U30571 (N_30571,N_30327,N_30284);
or U30572 (N_30572,N_30253,N_30311);
xnor U30573 (N_30573,N_30360,N_30418);
and U30574 (N_30574,N_30460,N_30322);
and U30575 (N_30575,N_30475,N_30390);
nand U30576 (N_30576,N_30312,N_30455);
and U30577 (N_30577,N_30442,N_30458);
xor U30578 (N_30578,N_30480,N_30271);
or U30579 (N_30579,N_30261,N_30381);
xor U30580 (N_30580,N_30344,N_30323);
nor U30581 (N_30581,N_30456,N_30356);
or U30582 (N_30582,N_30265,N_30427);
nand U30583 (N_30583,N_30474,N_30296);
nand U30584 (N_30584,N_30402,N_30355);
and U30585 (N_30585,N_30330,N_30293);
and U30586 (N_30586,N_30301,N_30450);
or U30587 (N_30587,N_30250,N_30357);
nor U30588 (N_30588,N_30389,N_30316);
and U30589 (N_30589,N_30299,N_30297);
or U30590 (N_30590,N_30383,N_30256);
nor U30591 (N_30591,N_30440,N_30375);
or U30592 (N_30592,N_30272,N_30291);
nor U30593 (N_30593,N_30352,N_30354);
and U30594 (N_30594,N_30358,N_30477);
or U30595 (N_30595,N_30340,N_30376);
or U30596 (N_30596,N_30469,N_30318);
or U30597 (N_30597,N_30444,N_30264);
nand U30598 (N_30598,N_30257,N_30489);
or U30599 (N_30599,N_30435,N_30423);
nand U30600 (N_30600,N_30414,N_30309);
xor U30601 (N_30601,N_30315,N_30325);
or U30602 (N_30602,N_30395,N_30310);
nor U30603 (N_30603,N_30405,N_30445);
or U30604 (N_30604,N_30319,N_30471);
nor U30605 (N_30605,N_30364,N_30342);
or U30606 (N_30606,N_30368,N_30447);
or U30607 (N_30607,N_30326,N_30351);
nand U30608 (N_30608,N_30420,N_30473);
and U30609 (N_30609,N_30270,N_30372);
and U30610 (N_30610,N_30386,N_30277);
nor U30611 (N_30611,N_30457,N_30350);
or U30612 (N_30612,N_30280,N_30436);
or U30613 (N_30613,N_30408,N_30413);
nor U30614 (N_30614,N_30463,N_30448);
or U30615 (N_30615,N_30353,N_30262);
or U30616 (N_30616,N_30490,N_30485);
or U30617 (N_30617,N_30438,N_30362);
nor U30618 (N_30618,N_30281,N_30439);
nor U30619 (N_30619,N_30415,N_30446);
xnor U30620 (N_30620,N_30399,N_30481);
or U30621 (N_30621,N_30252,N_30495);
xnor U30622 (N_30622,N_30449,N_30283);
and U30623 (N_30623,N_30255,N_30432);
nand U30624 (N_30624,N_30369,N_30498);
xor U30625 (N_30625,N_30387,N_30362);
or U30626 (N_30626,N_30496,N_30426);
or U30627 (N_30627,N_30273,N_30430);
nand U30628 (N_30628,N_30425,N_30263);
nor U30629 (N_30629,N_30305,N_30438);
or U30630 (N_30630,N_30490,N_30453);
nor U30631 (N_30631,N_30266,N_30411);
and U30632 (N_30632,N_30274,N_30295);
or U30633 (N_30633,N_30418,N_30335);
xor U30634 (N_30634,N_30367,N_30323);
or U30635 (N_30635,N_30291,N_30376);
or U30636 (N_30636,N_30431,N_30421);
or U30637 (N_30637,N_30286,N_30294);
and U30638 (N_30638,N_30470,N_30288);
xnor U30639 (N_30639,N_30261,N_30433);
xor U30640 (N_30640,N_30265,N_30466);
nor U30641 (N_30641,N_30483,N_30390);
or U30642 (N_30642,N_30488,N_30411);
and U30643 (N_30643,N_30439,N_30370);
nand U30644 (N_30644,N_30467,N_30395);
xnor U30645 (N_30645,N_30259,N_30265);
nand U30646 (N_30646,N_30468,N_30464);
or U30647 (N_30647,N_30316,N_30318);
nand U30648 (N_30648,N_30307,N_30347);
and U30649 (N_30649,N_30326,N_30308);
xnor U30650 (N_30650,N_30485,N_30326);
and U30651 (N_30651,N_30258,N_30380);
xor U30652 (N_30652,N_30484,N_30450);
nand U30653 (N_30653,N_30386,N_30411);
nand U30654 (N_30654,N_30388,N_30289);
or U30655 (N_30655,N_30311,N_30438);
nand U30656 (N_30656,N_30318,N_30272);
and U30657 (N_30657,N_30302,N_30487);
nand U30658 (N_30658,N_30295,N_30300);
and U30659 (N_30659,N_30404,N_30271);
and U30660 (N_30660,N_30437,N_30432);
and U30661 (N_30661,N_30280,N_30438);
nor U30662 (N_30662,N_30345,N_30254);
and U30663 (N_30663,N_30462,N_30396);
nor U30664 (N_30664,N_30499,N_30444);
or U30665 (N_30665,N_30416,N_30434);
and U30666 (N_30666,N_30324,N_30471);
and U30667 (N_30667,N_30469,N_30356);
and U30668 (N_30668,N_30300,N_30259);
nor U30669 (N_30669,N_30394,N_30497);
xor U30670 (N_30670,N_30313,N_30454);
nor U30671 (N_30671,N_30314,N_30318);
and U30672 (N_30672,N_30268,N_30333);
and U30673 (N_30673,N_30346,N_30440);
nand U30674 (N_30674,N_30252,N_30387);
xor U30675 (N_30675,N_30466,N_30302);
xnor U30676 (N_30676,N_30293,N_30464);
nand U30677 (N_30677,N_30413,N_30344);
nor U30678 (N_30678,N_30300,N_30286);
xor U30679 (N_30679,N_30353,N_30382);
nand U30680 (N_30680,N_30250,N_30377);
nand U30681 (N_30681,N_30463,N_30399);
nor U30682 (N_30682,N_30458,N_30293);
nor U30683 (N_30683,N_30493,N_30309);
nand U30684 (N_30684,N_30392,N_30347);
xor U30685 (N_30685,N_30458,N_30372);
or U30686 (N_30686,N_30460,N_30461);
xor U30687 (N_30687,N_30441,N_30278);
nor U30688 (N_30688,N_30464,N_30371);
or U30689 (N_30689,N_30452,N_30403);
nor U30690 (N_30690,N_30428,N_30465);
xor U30691 (N_30691,N_30321,N_30328);
xor U30692 (N_30692,N_30263,N_30270);
and U30693 (N_30693,N_30377,N_30453);
and U30694 (N_30694,N_30352,N_30419);
nand U30695 (N_30695,N_30325,N_30281);
or U30696 (N_30696,N_30329,N_30454);
xnor U30697 (N_30697,N_30391,N_30424);
xor U30698 (N_30698,N_30278,N_30357);
and U30699 (N_30699,N_30287,N_30261);
nand U30700 (N_30700,N_30490,N_30380);
and U30701 (N_30701,N_30499,N_30414);
or U30702 (N_30702,N_30480,N_30318);
xnor U30703 (N_30703,N_30326,N_30353);
xor U30704 (N_30704,N_30498,N_30443);
nand U30705 (N_30705,N_30289,N_30458);
and U30706 (N_30706,N_30432,N_30331);
or U30707 (N_30707,N_30388,N_30497);
and U30708 (N_30708,N_30395,N_30451);
xnor U30709 (N_30709,N_30482,N_30353);
or U30710 (N_30710,N_30418,N_30338);
or U30711 (N_30711,N_30406,N_30422);
xnor U30712 (N_30712,N_30475,N_30477);
and U30713 (N_30713,N_30435,N_30383);
nand U30714 (N_30714,N_30356,N_30492);
or U30715 (N_30715,N_30490,N_30280);
and U30716 (N_30716,N_30477,N_30479);
nand U30717 (N_30717,N_30378,N_30445);
or U30718 (N_30718,N_30328,N_30483);
or U30719 (N_30719,N_30271,N_30410);
or U30720 (N_30720,N_30429,N_30333);
nand U30721 (N_30721,N_30337,N_30491);
nor U30722 (N_30722,N_30338,N_30425);
and U30723 (N_30723,N_30349,N_30419);
or U30724 (N_30724,N_30304,N_30422);
nor U30725 (N_30725,N_30425,N_30436);
xor U30726 (N_30726,N_30482,N_30449);
nand U30727 (N_30727,N_30432,N_30485);
nor U30728 (N_30728,N_30365,N_30323);
nor U30729 (N_30729,N_30432,N_30314);
xor U30730 (N_30730,N_30350,N_30465);
nor U30731 (N_30731,N_30421,N_30354);
or U30732 (N_30732,N_30339,N_30396);
and U30733 (N_30733,N_30481,N_30257);
nor U30734 (N_30734,N_30303,N_30481);
or U30735 (N_30735,N_30318,N_30417);
nor U30736 (N_30736,N_30426,N_30303);
or U30737 (N_30737,N_30457,N_30491);
nor U30738 (N_30738,N_30302,N_30384);
xnor U30739 (N_30739,N_30258,N_30482);
xnor U30740 (N_30740,N_30268,N_30391);
and U30741 (N_30741,N_30265,N_30382);
nor U30742 (N_30742,N_30325,N_30474);
or U30743 (N_30743,N_30251,N_30415);
and U30744 (N_30744,N_30443,N_30471);
or U30745 (N_30745,N_30392,N_30271);
and U30746 (N_30746,N_30350,N_30347);
or U30747 (N_30747,N_30408,N_30444);
xnor U30748 (N_30748,N_30265,N_30394);
nor U30749 (N_30749,N_30273,N_30429);
and U30750 (N_30750,N_30623,N_30507);
xor U30751 (N_30751,N_30521,N_30617);
and U30752 (N_30752,N_30519,N_30523);
nand U30753 (N_30753,N_30604,N_30555);
nor U30754 (N_30754,N_30537,N_30638);
nand U30755 (N_30755,N_30731,N_30657);
xor U30756 (N_30756,N_30634,N_30746);
and U30757 (N_30757,N_30679,N_30533);
and U30758 (N_30758,N_30571,N_30705);
nor U30759 (N_30759,N_30573,N_30696);
and U30760 (N_30760,N_30745,N_30618);
nand U30761 (N_30761,N_30671,N_30632);
and U30762 (N_30762,N_30620,N_30644);
and U30763 (N_30763,N_30697,N_30504);
nand U30764 (N_30764,N_30542,N_30683);
xnor U30765 (N_30765,N_30538,N_30730);
xor U30766 (N_30766,N_30599,N_30548);
nor U30767 (N_30767,N_30635,N_30695);
nand U30768 (N_30768,N_30564,N_30626);
nand U30769 (N_30769,N_30596,N_30574);
and U30770 (N_30770,N_30743,N_30526);
nand U30771 (N_30771,N_30576,N_30556);
nand U30772 (N_30772,N_30649,N_30560);
and U30773 (N_30773,N_30744,N_30647);
nand U30774 (N_30774,N_30566,N_30678);
xor U30775 (N_30775,N_30568,N_30653);
xor U30776 (N_30776,N_30600,N_30723);
nand U30777 (N_30777,N_30546,N_30630);
xnor U30778 (N_30778,N_30572,N_30561);
nor U30779 (N_30779,N_30656,N_30606);
xnor U30780 (N_30780,N_30510,N_30633);
or U30781 (N_30781,N_30550,N_30693);
xnor U30782 (N_30782,N_30625,N_30524);
or U30783 (N_30783,N_30581,N_30684);
nand U30784 (N_30784,N_30594,N_30514);
or U30785 (N_30785,N_30607,N_30652);
or U30786 (N_30786,N_30513,N_30582);
and U30787 (N_30787,N_30502,N_30710);
nor U30788 (N_30788,N_30616,N_30639);
xnor U30789 (N_30789,N_30536,N_30569);
and U30790 (N_30790,N_30609,N_30682);
or U30791 (N_30791,N_30670,N_30545);
xor U30792 (N_30792,N_30528,N_30725);
nand U30793 (N_30793,N_30714,N_30559);
or U30794 (N_30794,N_30665,N_30651);
or U30795 (N_30795,N_30702,N_30701);
nor U30796 (N_30796,N_30552,N_30674);
nand U30797 (N_30797,N_30636,N_30584);
or U30798 (N_30798,N_30643,N_30726);
nand U30799 (N_30799,N_30516,N_30689);
or U30800 (N_30800,N_30578,N_30640);
nand U30801 (N_30801,N_30694,N_30722);
or U30802 (N_30802,N_30707,N_30737);
xnor U30803 (N_30803,N_30738,N_30704);
and U30804 (N_30804,N_30691,N_30733);
or U30805 (N_30805,N_30716,N_30668);
nor U30806 (N_30806,N_30642,N_30551);
or U30807 (N_30807,N_30512,N_30585);
xor U30808 (N_30808,N_30724,N_30655);
or U30809 (N_30809,N_30715,N_30648);
or U30810 (N_30810,N_30531,N_30747);
or U30811 (N_30811,N_30517,N_30669);
or U30812 (N_30812,N_30540,N_30699);
nand U30813 (N_30813,N_30590,N_30610);
or U30814 (N_30814,N_30698,N_30592);
or U30815 (N_30815,N_30562,N_30720);
xor U30816 (N_30816,N_30681,N_30664);
nand U30817 (N_30817,N_30565,N_30739);
and U30818 (N_30818,N_30660,N_30591);
and U30819 (N_30819,N_30532,N_30518);
nand U30820 (N_30820,N_30557,N_30709);
or U30821 (N_30821,N_30575,N_30735);
or U30822 (N_30822,N_30688,N_30577);
nand U30823 (N_30823,N_30719,N_30749);
and U30824 (N_30824,N_30692,N_30598);
and U30825 (N_30825,N_30520,N_30654);
nor U30826 (N_30826,N_30646,N_30666);
nand U30827 (N_30827,N_30706,N_30522);
nand U30828 (N_30828,N_30663,N_30621);
xor U30829 (N_30829,N_30718,N_30727);
nand U30830 (N_30830,N_30511,N_30658);
nand U30831 (N_30831,N_30586,N_30567);
nor U30832 (N_30832,N_30515,N_30539);
and U30833 (N_30833,N_30700,N_30662);
or U30834 (N_30834,N_30619,N_30628);
nand U30835 (N_30835,N_30506,N_30741);
xor U30836 (N_30836,N_30712,N_30736);
and U30837 (N_30837,N_30588,N_30641);
and U30838 (N_30838,N_30608,N_30593);
and U30839 (N_30839,N_30605,N_30602);
nor U30840 (N_30840,N_30535,N_30675);
xor U30841 (N_30841,N_30615,N_30583);
xor U30842 (N_30842,N_30614,N_30686);
and U30843 (N_30843,N_30547,N_30587);
or U30844 (N_30844,N_30673,N_30685);
and U30845 (N_30845,N_30589,N_30711);
nor U30846 (N_30846,N_30554,N_30627);
nor U30847 (N_30847,N_30734,N_30624);
xnor U30848 (N_30848,N_30612,N_30508);
xnor U30849 (N_30849,N_30509,N_30680);
nand U30850 (N_30850,N_30580,N_30717);
or U30851 (N_30851,N_30613,N_30611);
nor U30852 (N_30852,N_30553,N_30645);
or U30853 (N_30853,N_30687,N_30563);
nor U30854 (N_30854,N_30543,N_30534);
nor U30855 (N_30855,N_30558,N_30672);
xnor U30856 (N_30856,N_30505,N_30740);
nand U30857 (N_30857,N_30742,N_30661);
xnor U30858 (N_30858,N_30570,N_30597);
and U30859 (N_30859,N_30713,N_30622);
xnor U30860 (N_30860,N_30732,N_30650);
xor U30861 (N_30861,N_30629,N_30729);
or U30862 (N_30862,N_30541,N_30637);
nand U30863 (N_30863,N_30703,N_30708);
and U30864 (N_30864,N_30667,N_30527);
nand U30865 (N_30865,N_30525,N_30631);
xnor U30866 (N_30866,N_30530,N_30728);
and U30867 (N_30867,N_30676,N_30529);
nor U30868 (N_30868,N_30748,N_30579);
nand U30869 (N_30869,N_30603,N_30549);
xnor U30870 (N_30870,N_30690,N_30544);
and U30871 (N_30871,N_30601,N_30500);
xnor U30872 (N_30872,N_30501,N_30659);
xor U30873 (N_30873,N_30503,N_30677);
nand U30874 (N_30874,N_30721,N_30595);
or U30875 (N_30875,N_30637,N_30652);
or U30876 (N_30876,N_30685,N_30696);
nor U30877 (N_30877,N_30677,N_30572);
nor U30878 (N_30878,N_30569,N_30675);
and U30879 (N_30879,N_30621,N_30639);
and U30880 (N_30880,N_30743,N_30564);
nor U30881 (N_30881,N_30568,N_30586);
and U30882 (N_30882,N_30647,N_30728);
xnor U30883 (N_30883,N_30731,N_30728);
nand U30884 (N_30884,N_30715,N_30555);
and U30885 (N_30885,N_30588,N_30547);
or U30886 (N_30886,N_30652,N_30615);
nor U30887 (N_30887,N_30585,N_30679);
and U30888 (N_30888,N_30552,N_30691);
nor U30889 (N_30889,N_30558,N_30641);
nand U30890 (N_30890,N_30638,N_30741);
and U30891 (N_30891,N_30605,N_30690);
and U30892 (N_30892,N_30711,N_30648);
nor U30893 (N_30893,N_30563,N_30551);
nor U30894 (N_30894,N_30704,N_30713);
and U30895 (N_30895,N_30633,N_30570);
nor U30896 (N_30896,N_30594,N_30510);
xnor U30897 (N_30897,N_30611,N_30504);
nor U30898 (N_30898,N_30609,N_30630);
nand U30899 (N_30899,N_30584,N_30635);
nand U30900 (N_30900,N_30517,N_30691);
nand U30901 (N_30901,N_30518,N_30671);
xnor U30902 (N_30902,N_30556,N_30608);
xor U30903 (N_30903,N_30511,N_30581);
and U30904 (N_30904,N_30740,N_30624);
or U30905 (N_30905,N_30670,N_30746);
nand U30906 (N_30906,N_30508,N_30662);
nand U30907 (N_30907,N_30742,N_30709);
or U30908 (N_30908,N_30696,N_30676);
nand U30909 (N_30909,N_30699,N_30501);
and U30910 (N_30910,N_30532,N_30593);
and U30911 (N_30911,N_30515,N_30645);
and U30912 (N_30912,N_30519,N_30632);
nand U30913 (N_30913,N_30502,N_30520);
nand U30914 (N_30914,N_30504,N_30599);
xor U30915 (N_30915,N_30635,N_30702);
nor U30916 (N_30916,N_30730,N_30615);
nor U30917 (N_30917,N_30548,N_30740);
nor U30918 (N_30918,N_30561,N_30690);
and U30919 (N_30919,N_30580,N_30675);
xor U30920 (N_30920,N_30654,N_30556);
xor U30921 (N_30921,N_30574,N_30606);
and U30922 (N_30922,N_30704,N_30687);
nor U30923 (N_30923,N_30615,N_30739);
or U30924 (N_30924,N_30731,N_30627);
nor U30925 (N_30925,N_30575,N_30718);
nor U30926 (N_30926,N_30578,N_30528);
and U30927 (N_30927,N_30531,N_30629);
or U30928 (N_30928,N_30619,N_30504);
nand U30929 (N_30929,N_30591,N_30720);
and U30930 (N_30930,N_30575,N_30736);
or U30931 (N_30931,N_30661,N_30511);
xnor U30932 (N_30932,N_30544,N_30662);
or U30933 (N_30933,N_30532,N_30667);
xor U30934 (N_30934,N_30649,N_30653);
xnor U30935 (N_30935,N_30576,N_30590);
nand U30936 (N_30936,N_30542,N_30557);
nor U30937 (N_30937,N_30673,N_30552);
or U30938 (N_30938,N_30711,N_30630);
nor U30939 (N_30939,N_30590,N_30559);
xor U30940 (N_30940,N_30520,N_30507);
and U30941 (N_30941,N_30518,N_30574);
nand U30942 (N_30942,N_30722,N_30523);
xor U30943 (N_30943,N_30719,N_30568);
xor U30944 (N_30944,N_30707,N_30518);
nor U30945 (N_30945,N_30654,N_30512);
or U30946 (N_30946,N_30608,N_30665);
and U30947 (N_30947,N_30571,N_30600);
or U30948 (N_30948,N_30656,N_30660);
or U30949 (N_30949,N_30521,N_30594);
xnor U30950 (N_30950,N_30615,N_30509);
xor U30951 (N_30951,N_30705,N_30674);
and U30952 (N_30952,N_30733,N_30537);
nand U30953 (N_30953,N_30743,N_30745);
and U30954 (N_30954,N_30539,N_30744);
nand U30955 (N_30955,N_30700,N_30603);
nand U30956 (N_30956,N_30697,N_30659);
nor U30957 (N_30957,N_30562,N_30527);
xor U30958 (N_30958,N_30722,N_30690);
xor U30959 (N_30959,N_30539,N_30694);
or U30960 (N_30960,N_30615,N_30610);
or U30961 (N_30961,N_30605,N_30536);
xnor U30962 (N_30962,N_30576,N_30675);
nor U30963 (N_30963,N_30720,N_30595);
xnor U30964 (N_30964,N_30533,N_30691);
nor U30965 (N_30965,N_30688,N_30749);
xnor U30966 (N_30966,N_30586,N_30540);
and U30967 (N_30967,N_30663,N_30694);
or U30968 (N_30968,N_30622,N_30510);
nand U30969 (N_30969,N_30742,N_30685);
and U30970 (N_30970,N_30721,N_30502);
xnor U30971 (N_30971,N_30653,N_30535);
or U30972 (N_30972,N_30558,N_30737);
nor U30973 (N_30973,N_30511,N_30652);
and U30974 (N_30974,N_30687,N_30711);
nor U30975 (N_30975,N_30526,N_30562);
and U30976 (N_30976,N_30747,N_30603);
xnor U30977 (N_30977,N_30510,N_30602);
nand U30978 (N_30978,N_30511,N_30623);
or U30979 (N_30979,N_30726,N_30565);
and U30980 (N_30980,N_30573,N_30543);
and U30981 (N_30981,N_30587,N_30647);
or U30982 (N_30982,N_30633,N_30516);
xor U30983 (N_30983,N_30532,N_30665);
nand U30984 (N_30984,N_30681,N_30554);
nor U30985 (N_30985,N_30520,N_30634);
and U30986 (N_30986,N_30568,N_30699);
nor U30987 (N_30987,N_30515,N_30682);
nand U30988 (N_30988,N_30580,N_30695);
xnor U30989 (N_30989,N_30536,N_30730);
and U30990 (N_30990,N_30533,N_30588);
nor U30991 (N_30991,N_30502,N_30641);
nand U30992 (N_30992,N_30689,N_30737);
nand U30993 (N_30993,N_30643,N_30665);
nand U30994 (N_30994,N_30528,N_30712);
xnor U30995 (N_30995,N_30641,N_30672);
and U30996 (N_30996,N_30612,N_30630);
nand U30997 (N_30997,N_30646,N_30524);
or U30998 (N_30998,N_30699,N_30688);
and U30999 (N_30999,N_30526,N_30558);
and U31000 (N_31000,N_30804,N_30895);
nand U31001 (N_31001,N_30979,N_30763);
or U31002 (N_31002,N_30995,N_30867);
nand U31003 (N_31003,N_30816,N_30886);
nor U31004 (N_31004,N_30957,N_30925);
or U31005 (N_31005,N_30948,N_30938);
or U31006 (N_31006,N_30776,N_30965);
nor U31007 (N_31007,N_30836,N_30917);
or U31008 (N_31008,N_30906,N_30767);
or U31009 (N_31009,N_30978,N_30779);
nand U31010 (N_31010,N_30774,N_30819);
xor U31011 (N_31011,N_30991,N_30947);
or U31012 (N_31012,N_30857,N_30870);
nand U31013 (N_31013,N_30987,N_30798);
nand U31014 (N_31014,N_30990,N_30962);
nor U31015 (N_31015,N_30958,N_30810);
and U31016 (N_31016,N_30791,N_30863);
and U31017 (N_31017,N_30815,N_30828);
xnor U31018 (N_31018,N_30869,N_30770);
xor U31019 (N_31019,N_30854,N_30818);
and U31020 (N_31020,N_30907,N_30915);
nand U31021 (N_31021,N_30799,N_30797);
nor U31022 (N_31022,N_30878,N_30865);
xnor U31023 (N_31023,N_30795,N_30789);
nor U31024 (N_31024,N_30758,N_30927);
or U31025 (N_31025,N_30993,N_30902);
nand U31026 (N_31026,N_30899,N_30811);
xnor U31027 (N_31027,N_30900,N_30859);
and U31028 (N_31028,N_30998,N_30773);
and U31029 (N_31029,N_30969,N_30766);
and U31030 (N_31030,N_30997,N_30922);
xor U31031 (N_31031,N_30768,N_30891);
or U31032 (N_31032,N_30783,N_30796);
nand U31033 (N_31033,N_30834,N_30950);
nor U31034 (N_31034,N_30853,N_30762);
and U31035 (N_31035,N_30826,N_30806);
xnor U31036 (N_31036,N_30981,N_30843);
nor U31037 (N_31037,N_30982,N_30890);
and U31038 (N_31038,N_30793,N_30924);
nor U31039 (N_31039,N_30944,N_30866);
nor U31040 (N_31040,N_30852,N_30939);
nand U31041 (N_31041,N_30956,N_30802);
xor U31042 (N_31042,N_30999,N_30928);
nand U31043 (N_31043,N_30817,N_30889);
xnor U31044 (N_31044,N_30835,N_30918);
or U31045 (N_31045,N_30919,N_30750);
and U31046 (N_31046,N_30887,N_30970);
xnor U31047 (N_31047,N_30936,N_30851);
or U31048 (N_31048,N_30986,N_30864);
xor U31049 (N_31049,N_30967,N_30755);
and U31050 (N_31050,N_30882,N_30805);
xor U31051 (N_31051,N_30757,N_30841);
nand U31052 (N_31052,N_30908,N_30792);
and U31053 (N_31053,N_30959,N_30894);
nand U31054 (N_31054,N_30777,N_30976);
xor U31055 (N_31055,N_30994,N_30787);
nand U31056 (N_31056,N_30868,N_30881);
xor U31057 (N_31057,N_30984,N_30931);
nand U31058 (N_31058,N_30801,N_30973);
and U31059 (N_31059,N_30752,N_30814);
or U31060 (N_31060,N_30992,N_30856);
nand U31061 (N_31061,N_30808,N_30850);
nor U31062 (N_31062,N_30825,N_30968);
xor U31063 (N_31063,N_30892,N_30782);
nor U31064 (N_31064,N_30955,N_30842);
and U31065 (N_31065,N_30812,N_30961);
and U31066 (N_31066,N_30753,N_30830);
nand U31067 (N_31067,N_30897,N_30871);
or U31068 (N_31068,N_30769,N_30914);
xor U31069 (N_31069,N_30880,N_30831);
nand U31070 (N_31070,N_30949,N_30921);
xnor U31071 (N_31071,N_30858,N_30832);
nand U31072 (N_31072,N_30951,N_30775);
and U31073 (N_31073,N_30974,N_30874);
or U31074 (N_31074,N_30885,N_30855);
and U31075 (N_31075,N_30913,N_30904);
or U31076 (N_31076,N_30788,N_30903);
or U31077 (N_31077,N_30964,N_30943);
nor U31078 (N_31078,N_30821,N_30785);
nand U31079 (N_31079,N_30963,N_30909);
xnor U31080 (N_31080,N_30980,N_30920);
nand U31081 (N_31081,N_30960,N_30876);
nor U31082 (N_31082,N_30940,N_30946);
nand U31083 (N_31083,N_30845,N_30759);
xnor U31084 (N_31084,N_30778,N_30977);
nor U31085 (N_31085,N_30937,N_30760);
nor U31086 (N_31086,N_30846,N_30823);
or U31087 (N_31087,N_30942,N_30756);
nor U31088 (N_31088,N_30844,N_30848);
nand U31089 (N_31089,N_30875,N_30988);
xor U31090 (N_31090,N_30934,N_30790);
nor U31091 (N_31091,N_30879,N_30838);
nand U31092 (N_31092,N_30803,N_30829);
or U31093 (N_31093,N_30911,N_30923);
nand U31094 (N_31094,N_30824,N_30813);
xnor U31095 (N_31095,N_30954,N_30884);
and U31096 (N_31096,N_30784,N_30861);
nand U31097 (N_31097,N_30912,N_30833);
nor U31098 (N_31098,N_30972,N_30772);
and U31099 (N_31099,N_30771,N_30847);
or U31100 (N_31100,N_30765,N_30800);
or U31101 (N_31101,N_30929,N_30751);
xor U31102 (N_31102,N_30761,N_30933);
nand U31103 (N_31103,N_30985,N_30996);
or U31104 (N_31104,N_30860,N_30781);
nor U31105 (N_31105,N_30901,N_30935);
nand U31106 (N_31106,N_30820,N_30873);
nor U31107 (N_31107,N_30941,N_30893);
and U31108 (N_31108,N_30862,N_30827);
nor U31109 (N_31109,N_30930,N_30910);
and U31110 (N_31110,N_30898,N_30794);
nor U31111 (N_31111,N_30780,N_30809);
nor U31112 (N_31112,N_30849,N_30822);
nand U31113 (N_31113,N_30872,N_30926);
nand U31114 (N_31114,N_30952,N_30945);
nand U31115 (N_31115,N_30837,N_30989);
xor U31116 (N_31116,N_30786,N_30754);
and U31117 (N_31117,N_30905,N_30953);
xor U31118 (N_31118,N_30883,N_30839);
xnor U31119 (N_31119,N_30877,N_30896);
or U31120 (N_31120,N_30807,N_30975);
and U31121 (N_31121,N_30840,N_30966);
and U31122 (N_31122,N_30932,N_30971);
nand U31123 (N_31123,N_30888,N_30764);
nand U31124 (N_31124,N_30916,N_30983);
or U31125 (N_31125,N_30906,N_30770);
nor U31126 (N_31126,N_30907,N_30979);
nor U31127 (N_31127,N_30970,N_30808);
xor U31128 (N_31128,N_30867,N_30939);
xor U31129 (N_31129,N_30774,N_30914);
nor U31130 (N_31130,N_30977,N_30898);
and U31131 (N_31131,N_30884,N_30828);
and U31132 (N_31132,N_30956,N_30754);
and U31133 (N_31133,N_30865,N_30853);
nand U31134 (N_31134,N_30894,N_30987);
xor U31135 (N_31135,N_30756,N_30759);
or U31136 (N_31136,N_30882,N_30849);
nand U31137 (N_31137,N_30890,N_30964);
or U31138 (N_31138,N_30818,N_30796);
or U31139 (N_31139,N_30861,N_30947);
nor U31140 (N_31140,N_30876,N_30924);
nand U31141 (N_31141,N_30802,N_30794);
xnor U31142 (N_31142,N_30898,N_30833);
or U31143 (N_31143,N_30888,N_30984);
nor U31144 (N_31144,N_30770,N_30994);
and U31145 (N_31145,N_30947,N_30752);
xnor U31146 (N_31146,N_30755,N_30930);
xor U31147 (N_31147,N_30969,N_30802);
or U31148 (N_31148,N_30955,N_30823);
nand U31149 (N_31149,N_30921,N_30915);
nand U31150 (N_31150,N_30875,N_30884);
nand U31151 (N_31151,N_30772,N_30787);
or U31152 (N_31152,N_30860,N_30962);
nand U31153 (N_31153,N_30832,N_30878);
nand U31154 (N_31154,N_30790,N_30975);
xor U31155 (N_31155,N_30850,N_30821);
or U31156 (N_31156,N_30823,N_30917);
xnor U31157 (N_31157,N_30838,N_30804);
nor U31158 (N_31158,N_30937,N_30831);
and U31159 (N_31159,N_30965,N_30761);
nor U31160 (N_31160,N_30805,N_30990);
nor U31161 (N_31161,N_30976,N_30956);
and U31162 (N_31162,N_30802,N_30762);
and U31163 (N_31163,N_30863,N_30775);
or U31164 (N_31164,N_30759,N_30786);
nor U31165 (N_31165,N_30798,N_30923);
nor U31166 (N_31166,N_30820,N_30778);
or U31167 (N_31167,N_30915,N_30790);
nand U31168 (N_31168,N_30867,N_30889);
nand U31169 (N_31169,N_30920,N_30795);
xnor U31170 (N_31170,N_30934,N_30899);
and U31171 (N_31171,N_30911,N_30822);
nand U31172 (N_31172,N_30814,N_30945);
or U31173 (N_31173,N_30919,N_30867);
nand U31174 (N_31174,N_30789,N_30836);
and U31175 (N_31175,N_30972,N_30790);
xnor U31176 (N_31176,N_30761,N_30952);
xnor U31177 (N_31177,N_30839,N_30888);
or U31178 (N_31178,N_30861,N_30844);
and U31179 (N_31179,N_30881,N_30981);
or U31180 (N_31180,N_30838,N_30793);
or U31181 (N_31181,N_30958,N_30766);
or U31182 (N_31182,N_30844,N_30913);
nand U31183 (N_31183,N_30967,N_30819);
or U31184 (N_31184,N_30797,N_30814);
nor U31185 (N_31185,N_30996,N_30886);
nand U31186 (N_31186,N_30802,N_30861);
nand U31187 (N_31187,N_30772,N_30862);
nand U31188 (N_31188,N_30826,N_30797);
nand U31189 (N_31189,N_30972,N_30828);
or U31190 (N_31190,N_30943,N_30821);
xor U31191 (N_31191,N_30879,N_30798);
xor U31192 (N_31192,N_30804,N_30930);
and U31193 (N_31193,N_30889,N_30892);
and U31194 (N_31194,N_30885,N_30790);
and U31195 (N_31195,N_30967,N_30811);
nor U31196 (N_31196,N_30911,N_30818);
nor U31197 (N_31197,N_30941,N_30812);
or U31198 (N_31198,N_30912,N_30887);
nand U31199 (N_31199,N_30957,N_30818);
and U31200 (N_31200,N_30915,N_30901);
nor U31201 (N_31201,N_30855,N_30810);
nand U31202 (N_31202,N_30895,N_30878);
and U31203 (N_31203,N_30767,N_30916);
and U31204 (N_31204,N_30867,N_30763);
and U31205 (N_31205,N_30934,N_30788);
and U31206 (N_31206,N_30831,N_30950);
and U31207 (N_31207,N_30955,N_30757);
or U31208 (N_31208,N_30932,N_30875);
nand U31209 (N_31209,N_30973,N_30956);
nand U31210 (N_31210,N_30798,N_30836);
nor U31211 (N_31211,N_30981,N_30854);
nand U31212 (N_31212,N_30777,N_30871);
nor U31213 (N_31213,N_30876,N_30969);
nor U31214 (N_31214,N_30764,N_30865);
nand U31215 (N_31215,N_30804,N_30873);
nand U31216 (N_31216,N_30965,N_30925);
nand U31217 (N_31217,N_30810,N_30943);
xnor U31218 (N_31218,N_30932,N_30970);
xor U31219 (N_31219,N_30821,N_30927);
xnor U31220 (N_31220,N_30991,N_30945);
nand U31221 (N_31221,N_30891,N_30930);
xor U31222 (N_31222,N_30878,N_30945);
nand U31223 (N_31223,N_30982,N_30768);
xnor U31224 (N_31224,N_30954,N_30965);
or U31225 (N_31225,N_30821,N_30981);
and U31226 (N_31226,N_30906,N_30804);
nor U31227 (N_31227,N_30843,N_30806);
xor U31228 (N_31228,N_30926,N_30766);
or U31229 (N_31229,N_30761,N_30879);
nand U31230 (N_31230,N_30808,N_30904);
nand U31231 (N_31231,N_30990,N_30856);
and U31232 (N_31232,N_30798,N_30824);
or U31233 (N_31233,N_30839,N_30911);
or U31234 (N_31234,N_30754,N_30757);
nor U31235 (N_31235,N_30998,N_30865);
nand U31236 (N_31236,N_30811,N_30904);
xnor U31237 (N_31237,N_30753,N_30939);
and U31238 (N_31238,N_30935,N_30825);
or U31239 (N_31239,N_30877,N_30756);
nor U31240 (N_31240,N_30863,N_30954);
xor U31241 (N_31241,N_30975,N_30942);
and U31242 (N_31242,N_30808,N_30964);
and U31243 (N_31243,N_30757,N_30921);
and U31244 (N_31244,N_30853,N_30891);
nand U31245 (N_31245,N_30976,N_30792);
or U31246 (N_31246,N_30893,N_30755);
or U31247 (N_31247,N_30881,N_30899);
or U31248 (N_31248,N_30827,N_30905);
nor U31249 (N_31249,N_30965,N_30876);
and U31250 (N_31250,N_31059,N_31058);
nand U31251 (N_31251,N_31225,N_31229);
xnor U31252 (N_31252,N_31136,N_31205);
nand U31253 (N_31253,N_31184,N_31186);
nor U31254 (N_31254,N_31129,N_31192);
xor U31255 (N_31255,N_31240,N_31210);
and U31256 (N_31256,N_31032,N_31172);
or U31257 (N_31257,N_31090,N_31103);
nor U31258 (N_31258,N_31170,N_31246);
nor U31259 (N_31259,N_31006,N_31138);
nand U31260 (N_31260,N_31010,N_31015);
and U31261 (N_31261,N_31099,N_31197);
xnor U31262 (N_31262,N_31011,N_31101);
or U31263 (N_31263,N_31089,N_31017);
nor U31264 (N_31264,N_31004,N_31014);
nand U31265 (N_31265,N_31024,N_31031);
nand U31266 (N_31266,N_31143,N_31112);
xnor U31267 (N_31267,N_31066,N_31231);
nand U31268 (N_31268,N_31071,N_31209);
nor U31269 (N_31269,N_31007,N_31203);
nor U31270 (N_31270,N_31008,N_31081);
and U31271 (N_31271,N_31052,N_31030);
or U31272 (N_31272,N_31221,N_31181);
nor U31273 (N_31273,N_31086,N_31216);
and U31274 (N_31274,N_31085,N_31022);
nor U31275 (N_31275,N_31188,N_31061);
nor U31276 (N_31276,N_31135,N_31202);
nor U31277 (N_31277,N_31056,N_31185);
and U31278 (N_31278,N_31041,N_31180);
xor U31279 (N_31279,N_31157,N_31235);
nor U31280 (N_31280,N_31219,N_31005);
nor U31281 (N_31281,N_31106,N_31223);
or U31282 (N_31282,N_31070,N_31088);
xnor U31283 (N_31283,N_31108,N_31001);
xnor U31284 (N_31284,N_31177,N_31069);
nand U31285 (N_31285,N_31049,N_31153);
nor U31286 (N_31286,N_31207,N_31043);
nand U31287 (N_31287,N_31140,N_31206);
nand U31288 (N_31288,N_31178,N_31147);
and U31289 (N_31289,N_31174,N_31020);
and U31290 (N_31290,N_31166,N_31018);
nor U31291 (N_31291,N_31191,N_31169);
nand U31292 (N_31292,N_31176,N_31038);
and U31293 (N_31293,N_31104,N_31168);
nand U31294 (N_31294,N_31114,N_31167);
xnor U31295 (N_31295,N_31098,N_31237);
or U31296 (N_31296,N_31121,N_31062);
nand U31297 (N_31297,N_31116,N_31244);
nand U31298 (N_31298,N_31165,N_31187);
nand U31299 (N_31299,N_31164,N_31193);
xor U31300 (N_31300,N_31080,N_31072);
nand U31301 (N_31301,N_31123,N_31047);
nand U31302 (N_31302,N_31171,N_31033);
nor U31303 (N_31303,N_31087,N_31247);
and U31304 (N_31304,N_31236,N_31190);
nor U31305 (N_31305,N_31021,N_31074);
nand U31306 (N_31306,N_31002,N_31064);
and U31307 (N_31307,N_31162,N_31034);
nor U31308 (N_31308,N_31023,N_31084);
nand U31309 (N_31309,N_31158,N_31077);
nor U31310 (N_31310,N_31243,N_31012);
nand U31311 (N_31311,N_31161,N_31105);
nor U31312 (N_31312,N_31109,N_31128);
nor U31313 (N_31313,N_31029,N_31159);
nand U31314 (N_31314,N_31095,N_31196);
xnor U31315 (N_31315,N_31068,N_31051);
and U31316 (N_31316,N_31044,N_31218);
xnor U31317 (N_31317,N_31217,N_31226);
and U31318 (N_31318,N_31173,N_31242);
nand U31319 (N_31319,N_31097,N_31079);
nand U31320 (N_31320,N_31073,N_31233);
xnor U31321 (N_31321,N_31152,N_31137);
nor U31322 (N_31322,N_31125,N_31189);
nor U31323 (N_31323,N_31115,N_31148);
nand U31324 (N_31324,N_31102,N_31037);
nand U31325 (N_31325,N_31096,N_31027);
nand U31326 (N_31326,N_31025,N_31230);
nor U31327 (N_31327,N_31245,N_31139);
or U31328 (N_31328,N_31124,N_31026);
and U31329 (N_31329,N_31215,N_31212);
nand U31330 (N_31330,N_31144,N_31036);
xnor U31331 (N_31331,N_31122,N_31040);
nor U31332 (N_31332,N_31195,N_31057);
nor U31333 (N_31333,N_31042,N_31130);
or U31334 (N_31334,N_31100,N_31119);
nand U31335 (N_31335,N_31238,N_31228);
nor U31336 (N_31336,N_31082,N_31045);
nor U31337 (N_31337,N_31213,N_31076);
or U31338 (N_31338,N_31000,N_31132);
xnor U31339 (N_31339,N_31134,N_31151);
nor U31340 (N_31340,N_31232,N_31133);
xor U31341 (N_31341,N_31053,N_31118);
or U31342 (N_31342,N_31063,N_31019);
xnor U31343 (N_31343,N_31204,N_31046);
or U31344 (N_31344,N_31092,N_31039);
nand U31345 (N_31345,N_31055,N_31199);
xnor U31346 (N_31346,N_31003,N_31145);
and U31347 (N_31347,N_31150,N_31146);
xnor U31348 (N_31348,N_31198,N_31155);
and U31349 (N_31349,N_31160,N_31009);
xor U31350 (N_31350,N_31126,N_31141);
and U31351 (N_31351,N_31227,N_31175);
nand U31352 (N_31352,N_31065,N_31183);
nor U31353 (N_31353,N_31156,N_31094);
and U31354 (N_31354,N_31028,N_31163);
nor U31355 (N_31355,N_31013,N_31127);
and U31356 (N_31356,N_31016,N_31110);
or U31357 (N_31357,N_31054,N_31201);
nor U31358 (N_31358,N_31241,N_31200);
or U31359 (N_31359,N_31222,N_31208);
or U31360 (N_31360,N_31131,N_31067);
and U31361 (N_31361,N_31111,N_31220);
nor U31362 (N_31362,N_31249,N_31182);
nor U31363 (N_31363,N_31179,N_31048);
xor U31364 (N_31364,N_31075,N_31078);
and U31365 (N_31365,N_31060,N_31194);
nand U31366 (N_31366,N_31107,N_31211);
or U31367 (N_31367,N_31083,N_31239);
xor U31368 (N_31368,N_31234,N_31149);
xor U31369 (N_31369,N_31154,N_31050);
and U31370 (N_31370,N_31224,N_31120);
nand U31371 (N_31371,N_31093,N_31091);
xor U31372 (N_31372,N_31142,N_31035);
or U31373 (N_31373,N_31113,N_31214);
nor U31374 (N_31374,N_31117,N_31248);
nor U31375 (N_31375,N_31141,N_31086);
nor U31376 (N_31376,N_31027,N_31225);
and U31377 (N_31377,N_31015,N_31190);
nor U31378 (N_31378,N_31007,N_31118);
nand U31379 (N_31379,N_31124,N_31074);
and U31380 (N_31380,N_31244,N_31146);
nor U31381 (N_31381,N_31032,N_31223);
or U31382 (N_31382,N_31034,N_31128);
or U31383 (N_31383,N_31192,N_31064);
or U31384 (N_31384,N_31185,N_31183);
xnor U31385 (N_31385,N_31233,N_31038);
xnor U31386 (N_31386,N_31169,N_31038);
and U31387 (N_31387,N_31052,N_31057);
or U31388 (N_31388,N_31168,N_31006);
nor U31389 (N_31389,N_31242,N_31160);
nor U31390 (N_31390,N_31066,N_31071);
or U31391 (N_31391,N_31107,N_31060);
and U31392 (N_31392,N_31087,N_31126);
and U31393 (N_31393,N_31165,N_31201);
nand U31394 (N_31394,N_31195,N_31122);
or U31395 (N_31395,N_31222,N_31057);
or U31396 (N_31396,N_31059,N_31227);
nor U31397 (N_31397,N_31153,N_31224);
and U31398 (N_31398,N_31037,N_31223);
and U31399 (N_31399,N_31071,N_31141);
xnor U31400 (N_31400,N_31068,N_31202);
nand U31401 (N_31401,N_31106,N_31127);
or U31402 (N_31402,N_31017,N_31069);
nand U31403 (N_31403,N_31150,N_31023);
xnor U31404 (N_31404,N_31074,N_31116);
or U31405 (N_31405,N_31071,N_31038);
nand U31406 (N_31406,N_31056,N_31208);
nand U31407 (N_31407,N_31067,N_31208);
nor U31408 (N_31408,N_31220,N_31227);
nor U31409 (N_31409,N_31030,N_31059);
nor U31410 (N_31410,N_31036,N_31043);
xnor U31411 (N_31411,N_31181,N_31223);
and U31412 (N_31412,N_31002,N_31151);
xor U31413 (N_31413,N_31001,N_31220);
xor U31414 (N_31414,N_31116,N_31032);
xor U31415 (N_31415,N_31106,N_31030);
or U31416 (N_31416,N_31234,N_31187);
nor U31417 (N_31417,N_31003,N_31158);
nor U31418 (N_31418,N_31045,N_31140);
nor U31419 (N_31419,N_31115,N_31090);
xnor U31420 (N_31420,N_31131,N_31147);
nand U31421 (N_31421,N_31141,N_31093);
xor U31422 (N_31422,N_31120,N_31218);
nor U31423 (N_31423,N_31195,N_31168);
xnor U31424 (N_31424,N_31019,N_31043);
and U31425 (N_31425,N_31074,N_31203);
and U31426 (N_31426,N_31236,N_31037);
or U31427 (N_31427,N_31191,N_31185);
nand U31428 (N_31428,N_31108,N_31007);
and U31429 (N_31429,N_31081,N_31103);
and U31430 (N_31430,N_31151,N_31249);
and U31431 (N_31431,N_31133,N_31149);
xnor U31432 (N_31432,N_31110,N_31001);
nor U31433 (N_31433,N_31176,N_31173);
or U31434 (N_31434,N_31045,N_31179);
nand U31435 (N_31435,N_31008,N_31087);
nor U31436 (N_31436,N_31092,N_31233);
and U31437 (N_31437,N_31032,N_31171);
nand U31438 (N_31438,N_31119,N_31087);
nand U31439 (N_31439,N_31093,N_31235);
xnor U31440 (N_31440,N_31114,N_31008);
or U31441 (N_31441,N_31208,N_31098);
nor U31442 (N_31442,N_31228,N_31173);
and U31443 (N_31443,N_31209,N_31164);
nand U31444 (N_31444,N_31166,N_31004);
xnor U31445 (N_31445,N_31008,N_31174);
or U31446 (N_31446,N_31171,N_31246);
or U31447 (N_31447,N_31157,N_31045);
and U31448 (N_31448,N_31141,N_31103);
xnor U31449 (N_31449,N_31006,N_31102);
xor U31450 (N_31450,N_31015,N_31171);
xnor U31451 (N_31451,N_31106,N_31243);
and U31452 (N_31452,N_31139,N_31088);
or U31453 (N_31453,N_31068,N_31114);
xor U31454 (N_31454,N_31202,N_31065);
or U31455 (N_31455,N_31094,N_31245);
and U31456 (N_31456,N_31071,N_31188);
nand U31457 (N_31457,N_31241,N_31126);
or U31458 (N_31458,N_31198,N_31208);
nand U31459 (N_31459,N_31232,N_31131);
and U31460 (N_31460,N_31162,N_31059);
xor U31461 (N_31461,N_31160,N_31130);
and U31462 (N_31462,N_31203,N_31084);
nand U31463 (N_31463,N_31022,N_31001);
nor U31464 (N_31464,N_31117,N_31024);
or U31465 (N_31465,N_31064,N_31093);
or U31466 (N_31466,N_31140,N_31177);
nor U31467 (N_31467,N_31208,N_31152);
and U31468 (N_31468,N_31126,N_31027);
nand U31469 (N_31469,N_31053,N_31037);
or U31470 (N_31470,N_31159,N_31209);
nand U31471 (N_31471,N_31160,N_31039);
xor U31472 (N_31472,N_31075,N_31090);
xor U31473 (N_31473,N_31175,N_31033);
xnor U31474 (N_31474,N_31165,N_31067);
and U31475 (N_31475,N_31209,N_31009);
or U31476 (N_31476,N_31033,N_31060);
nand U31477 (N_31477,N_31210,N_31198);
or U31478 (N_31478,N_31130,N_31022);
nand U31479 (N_31479,N_31131,N_31231);
and U31480 (N_31480,N_31244,N_31016);
xor U31481 (N_31481,N_31059,N_31118);
and U31482 (N_31482,N_31103,N_31232);
nor U31483 (N_31483,N_31167,N_31146);
and U31484 (N_31484,N_31071,N_31146);
nand U31485 (N_31485,N_31111,N_31022);
xnor U31486 (N_31486,N_31087,N_31201);
xor U31487 (N_31487,N_31238,N_31236);
nor U31488 (N_31488,N_31070,N_31193);
nor U31489 (N_31489,N_31173,N_31245);
nand U31490 (N_31490,N_31148,N_31072);
nand U31491 (N_31491,N_31029,N_31061);
or U31492 (N_31492,N_31106,N_31099);
and U31493 (N_31493,N_31228,N_31172);
xor U31494 (N_31494,N_31007,N_31182);
and U31495 (N_31495,N_31198,N_31021);
or U31496 (N_31496,N_31002,N_31183);
nor U31497 (N_31497,N_31111,N_31148);
or U31498 (N_31498,N_31175,N_31055);
nor U31499 (N_31499,N_31241,N_31128);
and U31500 (N_31500,N_31446,N_31370);
or U31501 (N_31501,N_31336,N_31260);
xnor U31502 (N_31502,N_31478,N_31393);
and U31503 (N_31503,N_31359,N_31316);
xnor U31504 (N_31504,N_31412,N_31258);
nor U31505 (N_31505,N_31279,N_31272);
nand U31506 (N_31506,N_31474,N_31396);
xnor U31507 (N_31507,N_31318,N_31292);
and U31508 (N_31508,N_31368,N_31353);
nor U31509 (N_31509,N_31486,N_31466);
nor U31510 (N_31510,N_31265,N_31257);
or U31511 (N_31511,N_31340,N_31250);
or U31512 (N_31512,N_31496,N_31369);
xnor U31513 (N_31513,N_31358,N_31497);
nand U31514 (N_31514,N_31282,N_31286);
xor U31515 (N_31515,N_31442,N_31350);
xor U31516 (N_31516,N_31490,N_31306);
or U31517 (N_31517,N_31263,N_31410);
nand U31518 (N_31518,N_31295,N_31430);
nor U31519 (N_31519,N_31420,N_31328);
xnor U31520 (N_31520,N_31448,N_31329);
and U31521 (N_31521,N_31473,N_31348);
and U31522 (N_31522,N_31277,N_31366);
xnor U31523 (N_31523,N_31499,N_31262);
and U31524 (N_31524,N_31355,N_31480);
nor U31525 (N_31525,N_31450,N_31376);
or U31526 (N_31526,N_31371,N_31301);
nand U31527 (N_31527,N_31409,N_31281);
and U31528 (N_31528,N_31274,N_31352);
and U31529 (N_31529,N_31290,N_31303);
or U31530 (N_31530,N_31287,N_31405);
xnor U31531 (N_31531,N_31342,N_31417);
xor U31532 (N_31532,N_31307,N_31337);
nand U31533 (N_31533,N_31383,N_31331);
or U31534 (N_31534,N_31347,N_31462);
and U31535 (N_31535,N_31289,N_31382);
and U31536 (N_31536,N_31264,N_31300);
xnor U31537 (N_31537,N_31384,N_31381);
or U31538 (N_31538,N_31457,N_31404);
or U31539 (N_31539,N_31333,N_31356);
nand U31540 (N_31540,N_31275,N_31465);
and U31541 (N_31541,N_31492,N_31327);
or U31542 (N_31542,N_31406,N_31440);
and U31543 (N_31543,N_31494,N_31387);
or U31544 (N_31544,N_31380,N_31429);
or U31545 (N_31545,N_31471,N_31438);
xnor U31546 (N_31546,N_31373,N_31426);
nand U31547 (N_31547,N_31269,N_31365);
nor U31548 (N_31548,N_31361,N_31310);
and U31549 (N_31549,N_31447,N_31401);
nand U31550 (N_31550,N_31319,N_31255);
nand U31551 (N_31551,N_31425,N_31271);
nand U31552 (N_31552,N_31297,N_31252);
nor U31553 (N_31553,N_31311,N_31268);
xnor U31554 (N_31554,N_31345,N_31386);
nand U31555 (N_31555,N_31259,N_31445);
and U31556 (N_31556,N_31493,N_31253);
nor U31557 (N_31557,N_31360,N_31481);
and U31558 (N_31558,N_31304,N_31293);
xnor U31559 (N_31559,N_31283,N_31487);
xnor U31560 (N_31560,N_31472,N_31276);
nor U31561 (N_31561,N_31312,N_31285);
xnor U31562 (N_31562,N_31498,N_31261);
nor U31563 (N_31563,N_31408,N_31424);
nand U31564 (N_31564,N_31305,N_31362);
nor U31565 (N_31565,N_31294,N_31273);
and U31566 (N_31566,N_31339,N_31455);
xnor U31567 (N_31567,N_31431,N_31251);
xor U31568 (N_31568,N_31291,N_31334);
xor U31569 (N_31569,N_31418,N_31364);
or U31570 (N_31570,N_31313,N_31278);
nor U31571 (N_31571,N_31484,N_31254);
or U31572 (N_31572,N_31391,N_31323);
xor U31573 (N_31573,N_31256,N_31346);
nor U31574 (N_31574,N_31296,N_31476);
xor U31575 (N_31575,N_31422,N_31454);
or U31576 (N_31576,N_31439,N_31351);
or U31577 (N_31577,N_31437,N_31385);
xnor U31578 (N_31578,N_31427,N_31309);
nand U31579 (N_31579,N_31458,N_31389);
xor U31580 (N_31580,N_31357,N_31325);
nand U31581 (N_31581,N_31453,N_31320);
nand U31582 (N_31582,N_31392,N_31299);
xnor U31583 (N_31583,N_31367,N_31460);
nand U31584 (N_31584,N_31341,N_31267);
nor U31585 (N_31585,N_31374,N_31363);
nor U31586 (N_31586,N_31372,N_31449);
nand U31587 (N_31587,N_31379,N_31326);
nor U31588 (N_31588,N_31441,N_31377);
xnor U31589 (N_31589,N_31402,N_31475);
xnor U31590 (N_31590,N_31338,N_31403);
nor U31591 (N_31591,N_31280,N_31395);
and U31592 (N_31592,N_31324,N_31433);
or U31593 (N_31593,N_31332,N_31464);
or U31594 (N_31594,N_31467,N_31421);
xnor U31595 (N_31595,N_31321,N_31469);
and U31596 (N_31596,N_31463,N_31423);
nor U31597 (N_31597,N_31416,N_31399);
or U31598 (N_31598,N_31451,N_31468);
nor U31599 (N_31599,N_31434,N_31452);
nand U31600 (N_31600,N_31308,N_31398);
and U31601 (N_31601,N_31343,N_31270);
and U31602 (N_31602,N_31435,N_31488);
and U31603 (N_31603,N_31284,N_31495);
nor U31604 (N_31604,N_31335,N_31459);
or U31605 (N_31605,N_31428,N_31397);
xor U31606 (N_31606,N_31432,N_31477);
nand U31607 (N_31607,N_31436,N_31354);
xor U31608 (N_31608,N_31413,N_31411);
xor U31609 (N_31609,N_31414,N_31479);
and U31610 (N_31610,N_31407,N_31266);
or U31611 (N_31611,N_31317,N_31322);
nand U31612 (N_31612,N_31415,N_31444);
and U31613 (N_31613,N_31394,N_31344);
nor U31614 (N_31614,N_31314,N_31315);
nand U31615 (N_31615,N_31489,N_31470);
or U31616 (N_31616,N_31330,N_31375);
and U31617 (N_31617,N_31390,N_31482);
and U31618 (N_31618,N_31302,N_31456);
xor U31619 (N_31619,N_31400,N_31349);
xnor U31620 (N_31620,N_31485,N_31483);
nand U31621 (N_31621,N_31388,N_31288);
or U31622 (N_31622,N_31461,N_31298);
and U31623 (N_31623,N_31491,N_31443);
and U31624 (N_31624,N_31419,N_31378);
and U31625 (N_31625,N_31397,N_31394);
xnor U31626 (N_31626,N_31345,N_31319);
and U31627 (N_31627,N_31308,N_31315);
xor U31628 (N_31628,N_31386,N_31479);
nor U31629 (N_31629,N_31471,N_31262);
or U31630 (N_31630,N_31450,N_31356);
nor U31631 (N_31631,N_31450,N_31378);
nor U31632 (N_31632,N_31311,N_31341);
xor U31633 (N_31633,N_31260,N_31416);
xor U31634 (N_31634,N_31438,N_31363);
nand U31635 (N_31635,N_31288,N_31331);
nor U31636 (N_31636,N_31489,N_31252);
or U31637 (N_31637,N_31436,N_31386);
and U31638 (N_31638,N_31417,N_31498);
and U31639 (N_31639,N_31311,N_31449);
nand U31640 (N_31640,N_31387,N_31309);
xor U31641 (N_31641,N_31258,N_31395);
or U31642 (N_31642,N_31465,N_31497);
nand U31643 (N_31643,N_31303,N_31316);
nor U31644 (N_31644,N_31318,N_31335);
and U31645 (N_31645,N_31344,N_31325);
nor U31646 (N_31646,N_31314,N_31417);
nor U31647 (N_31647,N_31257,N_31423);
nand U31648 (N_31648,N_31494,N_31424);
or U31649 (N_31649,N_31446,N_31460);
or U31650 (N_31650,N_31305,N_31277);
xor U31651 (N_31651,N_31466,N_31311);
nor U31652 (N_31652,N_31257,N_31305);
nand U31653 (N_31653,N_31368,N_31310);
or U31654 (N_31654,N_31471,N_31338);
and U31655 (N_31655,N_31271,N_31459);
and U31656 (N_31656,N_31483,N_31452);
or U31657 (N_31657,N_31290,N_31398);
and U31658 (N_31658,N_31352,N_31439);
nand U31659 (N_31659,N_31490,N_31276);
and U31660 (N_31660,N_31387,N_31325);
and U31661 (N_31661,N_31468,N_31449);
or U31662 (N_31662,N_31310,N_31389);
nor U31663 (N_31663,N_31478,N_31301);
xnor U31664 (N_31664,N_31352,N_31495);
nor U31665 (N_31665,N_31339,N_31315);
or U31666 (N_31666,N_31329,N_31425);
and U31667 (N_31667,N_31494,N_31486);
or U31668 (N_31668,N_31499,N_31454);
and U31669 (N_31669,N_31304,N_31407);
and U31670 (N_31670,N_31415,N_31361);
nor U31671 (N_31671,N_31281,N_31282);
xnor U31672 (N_31672,N_31379,N_31408);
xnor U31673 (N_31673,N_31426,N_31423);
nor U31674 (N_31674,N_31340,N_31288);
nor U31675 (N_31675,N_31377,N_31298);
nor U31676 (N_31676,N_31257,N_31330);
nand U31677 (N_31677,N_31456,N_31478);
nand U31678 (N_31678,N_31436,N_31314);
nand U31679 (N_31679,N_31425,N_31306);
or U31680 (N_31680,N_31418,N_31440);
and U31681 (N_31681,N_31437,N_31446);
nor U31682 (N_31682,N_31270,N_31384);
xor U31683 (N_31683,N_31447,N_31264);
nor U31684 (N_31684,N_31290,N_31449);
nand U31685 (N_31685,N_31481,N_31469);
xor U31686 (N_31686,N_31351,N_31273);
or U31687 (N_31687,N_31280,N_31387);
and U31688 (N_31688,N_31452,N_31311);
and U31689 (N_31689,N_31451,N_31388);
or U31690 (N_31690,N_31326,N_31293);
or U31691 (N_31691,N_31313,N_31293);
nor U31692 (N_31692,N_31293,N_31266);
nand U31693 (N_31693,N_31380,N_31412);
or U31694 (N_31694,N_31357,N_31356);
or U31695 (N_31695,N_31401,N_31477);
nor U31696 (N_31696,N_31441,N_31406);
and U31697 (N_31697,N_31462,N_31291);
and U31698 (N_31698,N_31360,N_31413);
or U31699 (N_31699,N_31378,N_31322);
xnor U31700 (N_31700,N_31368,N_31347);
or U31701 (N_31701,N_31252,N_31303);
nor U31702 (N_31702,N_31350,N_31317);
or U31703 (N_31703,N_31377,N_31255);
nor U31704 (N_31704,N_31470,N_31325);
nor U31705 (N_31705,N_31372,N_31499);
nor U31706 (N_31706,N_31484,N_31401);
nand U31707 (N_31707,N_31377,N_31301);
nand U31708 (N_31708,N_31408,N_31321);
xor U31709 (N_31709,N_31401,N_31387);
and U31710 (N_31710,N_31316,N_31288);
and U31711 (N_31711,N_31474,N_31427);
or U31712 (N_31712,N_31407,N_31436);
xnor U31713 (N_31713,N_31416,N_31452);
and U31714 (N_31714,N_31409,N_31454);
or U31715 (N_31715,N_31435,N_31483);
nand U31716 (N_31716,N_31428,N_31284);
xnor U31717 (N_31717,N_31389,N_31288);
xnor U31718 (N_31718,N_31356,N_31329);
nand U31719 (N_31719,N_31371,N_31359);
nor U31720 (N_31720,N_31487,N_31424);
and U31721 (N_31721,N_31342,N_31402);
and U31722 (N_31722,N_31452,N_31463);
nand U31723 (N_31723,N_31493,N_31385);
xnor U31724 (N_31724,N_31326,N_31378);
nand U31725 (N_31725,N_31323,N_31435);
and U31726 (N_31726,N_31486,N_31328);
nand U31727 (N_31727,N_31494,N_31422);
and U31728 (N_31728,N_31262,N_31459);
xor U31729 (N_31729,N_31324,N_31355);
or U31730 (N_31730,N_31324,N_31440);
nand U31731 (N_31731,N_31320,N_31386);
nand U31732 (N_31732,N_31321,N_31430);
xor U31733 (N_31733,N_31295,N_31330);
or U31734 (N_31734,N_31477,N_31342);
nor U31735 (N_31735,N_31401,N_31437);
nand U31736 (N_31736,N_31344,N_31426);
nand U31737 (N_31737,N_31444,N_31331);
and U31738 (N_31738,N_31283,N_31426);
and U31739 (N_31739,N_31353,N_31335);
and U31740 (N_31740,N_31322,N_31274);
xnor U31741 (N_31741,N_31310,N_31423);
nor U31742 (N_31742,N_31368,N_31433);
or U31743 (N_31743,N_31398,N_31370);
nand U31744 (N_31744,N_31435,N_31450);
and U31745 (N_31745,N_31402,N_31318);
or U31746 (N_31746,N_31350,N_31289);
or U31747 (N_31747,N_31405,N_31462);
and U31748 (N_31748,N_31483,N_31252);
xor U31749 (N_31749,N_31415,N_31348);
or U31750 (N_31750,N_31645,N_31582);
nand U31751 (N_31751,N_31749,N_31660);
or U31752 (N_31752,N_31705,N_31644);
nor U31753 (N_31753,N_31630,N_31536);
and U31754 (N_31754,N_31597,N_31663);
nor U31755 (N_31755,N_31545,N_31509);
nand U31756 (N_31756,N_31659,N_31616);
and U31757 (N_31757,N_31642,N_31621);
or U31758 (N_31758,N_31599,N_31504);
nor U31759 (N_31759,N_31626,N_31500);
and U31760 (N_31760,N_31503,N_31627);
or U31761 (N_31761,N_31712,N_31513);
and U31762 (N_31762,N_31528,N_31638);
and U31763 (N_31763,N_31566,N_31696);
nor U31764 (N_31764,N_31611,N_31707);
nand U31765 (N_31765,N_31567,N_31591);
or U31766 (N_31766,N_31640,N_31649);
nand U31767 (N_31767,N_31550,N_31635);
and U31768 (N_31768,N_31526,N_31514);
nand U31769 (N_31769,N_31710,N_31547);
nor U31770 (N_31770,N_31537,N_31704);
nand U31771 (N_31771,N_31632,N_31676);
nand U31772 (N_31772,N_31685,N_31628);
xnor U31773 (N_31773,N_31650,N_31601);
nand U31774 (N_31774,N_31727,N_31714);
nor U31775 (N_31775,N_31581,N_31655);
and U31776 (N_31776,N_31561,N_31523);
nor U31777 (N_31777,N_31729,N_31680);
and U31778 (N_31778,N_31682,N_31726);
nor U31779 (N_31779,N_31706,N_31636);
nor U31780 (N_31780,N_31716,N_31665);
or U31781 (N_31781,N_31653,N_31548);
or U31782 (N_31782,N_31671,N_31595);
nand U31783 (N_31783,N_31607,N_31745);
nand U31784 (N_31784,N_31505,N_31692);
xor U31785 (N_31785,N_31613,N_31738);
or U31786 (N_31786,N_31694,N_31647);
and U31787 (N_31787,N_31715,N_31584);
and U31788 (N_31788,N_31546,N_31569);
xnor U31789 (N_31789,N_31551,N_31713);
and U31790 (N_31790,N_31560,N_31718);
or U31791 (N_31791,N_31512,N_31557);
nand U31792 (N_31792,N_31587,N_31668);
xnor U31793 (N_31793,N_31697,N_31717);
or U31794 (N_31794,N_31744,N_31552);
and U31795 (N_31795,N_31625,N_31728);
nor U31796 (N_31796,N_31686,N_31516);
and U31797 (N_31797,N_31565,N_31748);
nand U31798 (N_31798,N_31612,N_31579);
or U31799 (N_31799,N_31590,N_31593);
nor U31800 (N_31800,N_31654,N_31538);
xor U31801 (N_31801,N_31646,N_31652);
or U31802 (N_31802,N_31577,N_31656);
and U31803 (N_31803,N_31734,N_31708);
nor U31804 (N_31804,N_31699,N_31634);
nand U31805 (N_31805,N_31605,N_31604);
and U31806 (N_31806,N_31502,N_31598);
xnor U31807 (N_31807,N_31510,N_31683);
and U31808 (N_31808,N_31735,N_31633);
nor U31809 (N_31809,N_31639,N_31730);
and U31810 (N_31810,N_31690,N_31725);
or U31811 (N_31811,N_31622,N_31556);
nand U31812 (N_31812,N_31606,N_31583);
and U31813 (N_31813,N_31703,N_31677);
xnor U31814 (N_31814,N_31691,N_31662);
nand U31815 (N_31815,N_31602,N_31524);
nor U31816 (N_31816,N_31643,N_31614);
or U31817 (N_31817,N_31721,N_31506);
and U31818 (N_31818,N_31554,N_31670);
and U31819 (N_31819,N_31539,N_31520);
nand U31820 (N_31820,N_31501,N_31533);
and U31821 (N_31821,N_31573,N_31740);
nor U31822 (N_31822,N_31666,N_31674);
nand U31823 (N_31823,N_31511,N_31519);
and U31824 (N_31824,N_31742,N_31529);
nand U31825 (N_31825,N_31540,N_31555);
nor U31826 (N_31826,N_31518,N_31695);
xor U31827 (N_31827,N_31688,N_31578);
and U31828 (N_31828,N_31594,N_31693);
nand U31829 (N_31829,N_31631,N_31572);
nor U31830 (N_31830,N_31571,N_31576);
xnor U31831 (N_31831,N_31570,N_31684);
nand U31832 (N_31832,N_31617,N_31711);
xor U31833 (N_31833,N_31563,N_31574);
nor U31834 (N_31834,N_31553,N_31589);
xor U31835 (N_31835,N_31722,N_31673);
and U31836 (N_31836,N_31702,N_31596);
nor U31837 (N_31837,N_31619,N_31580);
xor U31838 (N_31838,N_31588,N_31736);
and U31839 (N_31839,N_31681,N_31527);
and U31840 (N_31840,N_31568,N_31618);
and U31841 (N_31841,N_31507,N_31603);
xnor U31842 (N_31842,N_31530,N_31562);
xor U31843 (N_31843,N_31532,N_31542);
xor U31844 (N_31844,N_31575,N_31531);
xnor U31845 (N_31845,N_31737,N_31675);
or U31846 (N_31846,N_31623,N_31741);
and U31847 (N_31847,N_31664,N_31658);
nor U31848 (N_31848,N_31661,N_31610);
nand U31849 (N_31849,N_31672,N_31641);
xor U31850 (N_31850,N_31558,N_31564);
nand U31851 (N_31851,N_31657,N_31586);
nor U31852 (N_31852,N_31678,N_31667);
nor U31853 (N_31853,N_31620,N_31600);
or U31854 (N_31854,N_31508,N_31709);
and U31855 (N_31855,N_31534,N_31747);
or U31856 (N_31856,N_31525,N_31651);
and U31857 (N_31857,N_31723,N_31535);
and U31858 (N_31858,N_31592,N_31724);
or U31859 (N_31859,N_31698,N_31544);
or U31860 (N_31860,N_31637,N_31746);
xor U31861 (N_31861,N_31541,N_31549);
and U31862 (N_31862,N_31732,N_31719);
nor U31863 (N_31863,N_31739,N_31624);
and U31864 (N_31864,N_31733,N_31720);
nor U31865 (N_31865,N_31700,N_31689);
xnor U31866 (N_31866,N_31669,N_31629);
xnor U31867 (N_31867,N_31521,N_31679);
nand U31868 (N_31868,N_31522,N_31543);
and U31869 (N_31869,N_31731,N_31517);
nand U31870 (N_31870,N_31687,N_31609);
xor U31871 (N_31871,N_31559,N_31743);
or U31872 (N_31872,N_31608,N_31585);
and U31873 (N_31873,N_31615,N_31515);
nor U31874 (N_31874,N_31648,N_31701);
nor U31875 (N_31875,N_31656,N_31645);
or U31876 (N_31876,N_31594,N_31548);
nand U31877 (N_31877,N_31715,N_31573);
or U31878 (N_31878,N_31681,N_31715);
and U31879 (N_31879,N_31533,N_31704);
nand U31880 (N_31880,N_31616,N_31518);
nand U31881 (N_31881,N_31699,N_31721);
xor U31882 (N_31882,N_31721,N_31653);
xor U31883 (N_31883,N_31652,N_31749);
or U31884 (N_31884,N_31729,N_31547);
and U31885 (N_31885,N_31735,N_31609);
or U31886 (N_31886,N_31571,N_31575);
or U31887 (N_31887,N_31600,N_31647);
nand U31888 (N_31888,N_31745,N_31682);
nor U31889 (N_31889,N_31631,N_31640);
nor U31890 (N_31890,N_31500,N_31525);
or U31891 (N_31891,N_31639,N_31638);
and U31892 (N_31892,N_31510,N_31578);
nand U31893 (N_31893,N_31728,N_31597);
or U31894 (N_31894,N_31648,N_31611);
xnor U31895 (N_31895,N_31671,N_31545);
and U31896 (N_31896,N_31745,N_31533);
or U31897 (N_31897,N_31594,N_31589);
and U31898 (N_31898,N_31724,N_31738);
or U31899 (N_31899,N_31662,N_31616);
and U31900 (N_31900,N_31586,N_31700);
or U31901 (N_31901,N_31592,N_31630);
xor U31902 (N_31902,N_31681,N_31638);
xor U31903 (N_31903,N_31629,N_31607);
nand U31904 (N_31904,N_31713,N_31702);
xnor U31905 (N_31905,N_31703,N_31639);
xor U31906 (N_31906,N_31541,N_31565);
nand U31907 (N_31907,N_31735,N_31727);
xor U31908 (N_31908,N_31728,N_31563);
or U31909 (N_31909,N_31638,N_31660);
xor U31910 (N_31910,N_31687,N_31676);
nand U31911 (N_31911,N_31738,N_31585);
or U31912 (N_31912,N_31657,N_31585);
xnor U31913 (N_31913,N_31706,N_31733);
or U31914 (N_31914,N_31585,N_31710);
nor U31915 (N_31915,N_31701,N_31675);
nand U31916 (N_31916,N_31591,N_31629);
or U31917 (N_31917,N_31647,N_31538);
xnor U31918 (N_31918,N_31556,N_31506);
nor U31919 (N_31919,N_31548,N_31725);
or U31920 (N_31920,N_31745,N_31690);
xnor U31921 (N_31921,N_31524,N_31732);
or U31922 (N_31922,N_31727,N_31649);
nor U31923 (N_31923,N_31598,N_31703);
xnor U31924 (N_31924,N_31605,N_31540);
or U31925 (N_31925,N_31648,N_31695);
nor U31926 (N_31926,N_31598,N_31530);
or U31927 (N_31927,N_31607,N_31581);
or U31928 (N_31928,N_31662,N_31557);
xnor U31929 (N_31929,N_31607,N_31675);
or U31930 (N_31930,N_31589,N_31501);
nor U31931 (N_31931,N_31588,N_31712);
or U31932 (N_31932,N_31554,N_31563);
nor U31933 (N_31933,N_31703,N_31671);
nor U31934 (N_31934,N_31659,N_31539);
nor U31935 (N_31935,N_31725,N_31702);
nand U31936 (N_31936,N_31714,N_31624);
nand U31937 (N_31937,N_31606,N_31730);
and U31938 (N_31938,N_31580,N_31550);
nand U31939 (N_31939,N_31721,N_31739);
nand U31940 (N_31940,N_31620,N_31554);
and U31941 (N_31941,N_31642,N_31559);
and U31942 (N_31942,N_31718,N_31644);
xnor U31943 (N_31943,N_31595,N_31602);
and U31944 (N_31944,N_31581,N_31707);
or U31945 (N_31945,N_31683,N_31574);
nand U31946 (N_31946,N_31634,N_31524);
and U31947 (N_31947,N_31644,N_31716);
xor U31948 (N_31948,N_31561,N_31535);
and U31949 (N_31949,N_31746,N_31587);
xor U31950 (N_31950,N_31562,N_31547);
or U31951 (N_31951,N_31614,N_31717);
or U31952 (N_31952,N_31670,N_31726);
and U31953 (N_31953,N_31726,N_31504);
and U31954 (N_31954,N_31562,N_31594);
nor U31955 (N_31955,N_31559,N_31689);
and U31956 (N_31956,N_31748,N_31734);
nand U31957 (N_31957,N_31634,N_31630);
xnor U31958 (N_31958,N_31517,N_31563);
and U31959 (N_31959,N_31503,N_31704);
xor U31960 (N_31960,N_31593,N_31592);
xnor U31961 (N_31961,N_31628,N_31647);
nor U31962 (N_31962,N_31733,N_31509);
nor U31963 (N_31963,N_31502,N_31693);
nand U31964 (N_31964,N_31747,N_31630);
and U31965 (N_31965,N_31514,N_31635);
nor U31966 (N_31966,N_31531,N_31706);
nor U31967 (N_31967,N_31706,N_31612);
or U31968 (N_31968,N_31515,N_31653);
nor U31969 (N_31969,N_31705,N_31538);
or U31970 (N_31970,N_31663,N_31522);
nor U31971 (N_31971,N_31631,N_31526);
and U31972 (N_31972,N_31596,N_31600);
or U31973 (N_31973,N_31686,N_31713);
nand U31974 (N_31974,N_31607,N_31662);
or U31975 (N_31975,N_31664,N_31656);
nand U31976 (N_31976,N_31645,N_31686);
and U31977 (N_31977,N_31746,N_31594);
nor U31978 (N_31978,N_31730,N_31705);
and U31979 (N_31979,N_31704,N_31640);
xor U31980 (N_31980,N_31601,N_31715);
nor U31981 (N_31981,N_31659,N_31526);
or U31982 (N_31982,N_31673,N_31671);
nor U31983 (N_31983,N_31572,N_31548);
nor U31984 (N_31984,N_31522,N_31534);
or U31985 (N_31985,N_31526,N_31551);
or U31986 (N_31986,N_31731,N_31509);
xnor U31987 (N_31987,N_31632,N_31505);
nand U31988 (N_31988,N_31743,N_31710);
xor U31989 (N_31989,N_31589,N_31710);
xor U31990 (N_31990,N_31613,N_31699);
and U31991 (N_31991,N_31643,N_31715);
and U31992 (N_31992,N_31510,N_31678);
xnor U31993 (N_31993,N_31536,N_31551);
and U31994 (N_31994,N_31513,N_31683);
xor U31995 (N_31995,N_31693,N_31556);
and U31996 (N_31996,N_31698,N_31722);
nand U31997 (N_31997,N_31547,N_31516);
or U31998 (N_31998,N_31512,N_31521);
xor U31999 (N_31999,N_31708,N_31632);
or U32000 (N_32000,N_31967,N_31753);
nor U32001 (N_32001,N_31974,N_31867);
nand U32002 (N_32002,N_31861,N_31751);
nor U32003 (N_32003,N_31863,N_31977);
and U32004 (N_32004,N_31781,N_31878);
nand U32005 (N_32005,N_31814,N_31813);
xor U32006 (N_32006,N_31903,N_31824);
nand U32007 (N_32007,N_31833,N_31957);
xnor U32008 (N_32008,N_31775,N_31979);
xor U32009 (N_32009,N_31800,N_31755);
or U32010 (N_32010,N_31963,N_31951);
xnor U32011 (N_32011,N_31795,N_31921);
nand U32012 (N_32012,N_31966,N_31990);
nor U32013 (N_32013,N_31865,N_31986);
or U32014 (N_32014,N_31890,N_31831);
nand U32015 (N_32015,N_31932,N_31756);
or U32016 (N_32016,N_31772,N_31952);
or U32017 (N_32017,N_31891,N_31776);
nand U32018 (N_32018,N_31931,N_31823);
xor U32019 (N_32019,N_31994,N_31939);
nor U32020 (N_32020,N_31774,N_31769);
nand U32021 (N_32021,N_31857,N_31782);
and U32022 (N_32022,N_31898,N_31873);
nor U32023 (N_32023,N_31999,N_31911);
nand U32024 (N_32024,N_31920,N_31950);
xor U32025 (N_32025,N_31914,N_31760);
xnor U32026 (N_32026,N_31758,N_31810);
or U32027 (N_32027,N_31848,N_31837);
and U32028 (N_32028,N_31777,N_31991);
nand U32029 (N_32029,N_31997,N_31959);
nand U32030 (N_32030,N_31904,N_31993);
and U32031 (N_32031,N_31802,N_31875);
and U32032 (N_32032,N_31825,N_31801);
nor U32033 (N_32033,N_31841,N_31763);
nand U32034 (N_32034,N_31757,N_31944);
or U32035 (N_32035,N_31815,N_31936);
nor U32036 (N_32036,N_31754,N_31877);
and U32037 (N_32037,N_31830,N_31962);
nand U32038 (N_32038,N_31924,N_31874);
or U32039 (N_32039,N_31826,N_31960);
and U32040 (N_32040,N_31850,N_31956);
nand U32041 (N_32041,N_31893,N_31886);
and U32042 (N_32042,N_31807,N_31929);
nor U32043 (N_32043,N_31750,N_31858);
or U32044 (N_32044,N_31928,N_31766);
nor U32045 (N_32045,N_31840,N_31899);
xnor U32046 (N_32046,N_31786,N_31803);
nor U32047 (N_32047,N_31905,N_31768);
nand U32048 (N_32048,N_31938,N_31771);
nand U32049 (N_32049,N_31976,N_31883);
nand U32050 (N_32050,N_31853,N_31933);
nand U32051 (N_32051,N_31918,N_31934);
nand U32052 (N_32052,N_31961,N_31971);
xnor U32053 (N_32053,N_31852,N_31790);
nand U32054 (N_32054,N_31995,N_31972);
nand U32055 (N_32055,N_31925,N_31882);
xnor U32056 (N_32056,N_31985,N_31779);
nand U32057 (N_32057,N_31909,N_31799);
nand U32058 (N_32058,N_31923,N_31838);
nand U32059 (N_32059,N_31855,N_31888);
xor U32060 (N_32060,N_31998,N_31992);
nand U32061 (N_32061,N_31770,N_31884);
nand U32062 (N_32062,N_31780,N_31839);
xor U32063 (N_32063,N_31922,N_31806);
and U32064 (N_32064,N_31989,N_31844);
or U32065 (N_32065,N_31942,N_31968);
and U32066 (N_32066,N_31879,N_31902);
nand U32067 (N_32067,N_31940,N_31819);
and U32068 (N_32068,N_31864,N_31761);
or U32069 (N_32069,N_31881,N_31862);
nand U32070 (N_32070,N_31788,N_31785);
or U32071 (N_32071,N_31906,N_31912);
and U32072 (N_32072,N_31842,N_31859);
or U32073 (N_32073,N_31870,N_31797);
or U32074 (N_32074,N_31953,N_31818);
or U32075 (N_32075,N_31847,N_31869);
nand U32076 (N_32076,N_31856,N_31835);
nand U32077 (N_32077,N_31778,N_31773);
nor U32078 (N_32078,N_31901,N_31954);
nand U32079 (N_32079,N_31783,N_31964);
xnor U32080 (N_32080,N_31784,N_31871);
and U32081 (N_32081,N_31948,N_31913);
nand U32082 (N_32082,N_31980,N_31908);
or U32083 (N_32083,N_31987,N_31935);
nor U32084 (N_32084,N_31759,N_31827);
nand U32085 (N_32085,N_31880,N_31836);
or U32086 (N_32086,N_31941,N_31981);
xor U32087 (N_32087,N_31868,N_31793);
nor U32088 (N_32088,N_31876,N_31970);
and U32089 (N_32089,N_31958,N_31927);
nand U32090 (N_32090,N_31812,N_31787);
nor U32091 (N_32091,N_31791,N_31820);
or U32092 (N_32092,N_31907,N_31796);
xnor U32093 (N_32093,N_31817,N_31765);
and U32094 (N_32094,N_31917,N_31764);
xnor U32095 (N_32095,N_31860,N_31792);
nand U32096 (N_32096,N_31984,N_31866);
nand U32097 (N_32097,N_31829,N_31965);
nor U32098 (N_32098,N_31804,N_31975);
or U32099 (N_32099,N_31849,N_31798);
or U32100 (N_32100,N_31910,N_31762);
xor U32101 (N_32101,N_31794,N_31955);
xnor U32102 (N_32102,N_31892,N_31937);
xor U32103 (N_32103,N_31843,N_31816);
and U32104 (N_32104,N_31809,N_31752);
or U32105 (N_32105,N_31945,N_31943);
nor U32106 (N_32106,N_31811,N_31854);
and U32107 (N_32107,N_31789,N_31919);
or U32108 (N_32108,N_31805,N_31808);
nor U32109 (N_32109,N_31885,N_31900);
nand U32110 (N_32110,N_31983,N_31851);
and U32111 (N_32111,N_31828,N_31988);
and U32112 (N_32112,N_31889,N_31846);
and U32113 (N_32113,N_31896,N_31996);
xnor U32114 (N_32114,N_31832,N_31821);
nor U32115 (N_32115,N_31915,N_31895);
xor U32116 (N_32116,N_31916,N_31946);
xnor U32117 (N_32117,N_31887,N_31947);
nor U32118 (N_32118,N_31872,N_31845);
nor U32119 (N_32119,N_31982,N_31949);
nand U32120 (N_32120,N_31834,N_31897);
xor U32121 (N_32121,N_31767,N_31822);
and U32122 (N_32122,N_31973,N_31926);
nand U32123 (N_32123,N_31978,N_31930);
nand U32124 (N_32124,N_31894,N_31969);
and U32125 (N_32125,N_31753,N_31758);
nand U32126 (N_32126,N_31798,N_31954);
and U32127 (N_32127,N_31932,N_31905);
nand U32128 (N_32128,N_31936,N_31821);
nand U32129 (N_32129,N_31916,N_31776);
and U32130 (N_32130,N_31781,N_31893);
and U32131 (N_32131,N_31947,N_31776);
xor U32132 (N_32132,N_31901,N_31849);
or U32133 (N_32133,N_31832,N_31967);
xor U32134 (N_32134,N_31982,N_31954);
xnor U32135 (N_32135,N_31794,N_31861);
nor U32136 (N_32136,N_31790,N_31886);
nand U32137 (N_32137,N_31900,N_31909);
and U32138 (N_32138,N_31919,N_31821);
xnor U32139 (N_32139,N_31754,N_31912);
nor U32140 (N_32140,N_31964,N_31860);
nand U32141 (N_32141,N_31883,N_31974);
or U32142 (N_32142,N_31843,N_31951);
nor U32143 (N_32143,N_31948,N_31971);
or U32144 (N_32144,N_31857,N_31886);
and U32145 (N_32145,N_31996,N_31831);
nor U32146 (N_32146,N_31959,N_31777);
and U32147 (N_32147,N_31972,N_31752);
xnor U32148 (N_32148,N_31789,N_31873);
nor U32149 (N_32149,N_31850,N_31994);
nor U32150 (N_32150,N_31836,N_31814);
nand U32151 (N_32151,N_31970,N_31828);
or U32152 (N_32152,N_31779,N_31963);
and U32153 (N_32153,N_31866,N_31851);
nand U32154 (N_32154,N_31805,N_31832);
xor U32155 (N_32155,N_31999,N_31754);
nor U32156 (N_32156,N_31973,N_31852);
nor U32157 (N_32157,N_31840,N_31761);
nand U32158 (N_32158,N_31957,N_31988);
xor U32159 (N_32159,N_31923,N_31882);
and U32160 (N_32160,N_31901,N_31810);
xnor U32161 (N_32161,N_31918,N_31971);
nand U32162 (N_32162,N_31806,N_31811);
nand U32163 (N_32163,N_31922,N_31991);
nor U32164 (N_32164,N_31959,N_31895);
nand U32165 (N_32165,N_31825,N_31938);
nor U32166 (N_32166,N_31799,N_31805);
or U32167 (N_32167,N_31758,N_31822);
nand U32168 (N_32168,N_31876,N_31751);
nand U32169 (N_32169,N_31866,N_31827);
and U32170 (N_32170,N_31937,N_31925);
nand U32171 (N_32171,N_31754,N_31783);
nor U32172 (N_32172,N_31777,N_31846);
or U32173 (N_32173,N_31816,N_31915);
nand U32174 (N_32174,N_31990,N_31978);
xor U32175 (N_32175,N_31989,N_31869);
nor U32176 (N_32176,N_31856,N_31892);
nor U32177 (N_32177,N_31949,N_31777);
xnor U32178 (N_32178,N_31756,N_31918);
or U32179 (N_32179,N_31842,N_31780);
and U32180 (N_32180,N_31915,N_31952);
xor U32181 (N_32181,N_31948,N_31979);
xor U32182 (N_32182,N_31814,N_31848);
nor U32183 (N_32183,N_31794,N_31773);
nor U32184 (N_32184,N_31767,N_31789);
or U32185 (N_32185,N_31874,N_31798);
nor U32186 (N_32186,N_31976,N_31979);
nor U32187 (N_32187,N_31876,N_31804);
xnor U32188 (N_32188,N_31840,N_31998);
and U32189 (N_32189,N_31770,N_31949);
nand U32190 (N_32190,N_31839,N_31835);
or U32191 (N_32191,N_31816,N_31811);
nand U32192 (N_32192,N_31877,N_31885);
xor U32193 (N_32193,N_31866,N_31928);
nand U32194 (N_32194,N_31793,N_31936);
nor U32195 (N_32195,N_31792,N_31968);
xnor U32196 (N_32196,N_31857,N_31751);
and U32197 (N_32197,N_31760,N_31826);
or U32198 (N_32198,N_31957,N_31862);
nand U32199 (N_32199,N_31926,N_31823);
nand U32200 (N_32200,N_31989,N_31915);
xor U32201 (N_32201,N_31981,N_31810);
xnor U32202 (N_32202,N_31966,N_31916);
xor U32203 (N_32203,N_31790,N_31770);
nor U32204 (N_32204,N_31760,N_31968);
and U32205 (N_32205,N_31780,N_31962);
nor U32206 (N_32206,N_31822,N_31933);
xor U32207 (N_32207,N_31798,N_31987);
or U32208 (N_32208,N_31806,N_31973);
and U32209 (N_32209,N_31912,N_31848);
or U32210 (N_32210,N_31905,N_31815);
nor U32211 (N_32211,N_31859,N_31852);
or U32212 (N_32212,N_31826,N_31955);
and U32213 (N_32213,N_31884,N_31896);
or U32214 (N_32214,N_31929,N_31966);
xor U32215 (N_32215,N_31905,N_31756);
nand U32216 (N_32216,N_31790,N_31813);
nand U32217 (N_32217,N_31798,N_31820);
nand U32218 (N_32218,N_31762,N_31872);
nor U32219 (N_32219,N_31846,N_31866);
xor U32220 (N_32220,N_31949,N_31771);
nor U32221 (N_32221,N_31961,N_31889);
nor U32222 (N_32222,N_31922,N_31977);
or U32223 (N_32223,N_31805,N_31931);
nor U32224 (N_32224,N_31912,N_31828);
and U32225 (N_32225,N_31869,N_31985);
and U32226 (N_32226,N_31807,N_31816);
xnor U32227 (N_32227,N_31976,N_31836);
nor U32228 (N_32228,N_31797,N_31783);
and U32229 (N_32229,N_31928,N_31969);
nand U32230 (N_32230,N_31976,N_31782);
xnor U32231 (N_32231,N_31769,N_31972);
and U32232 (N_32232,N_31867,N_31812);
and U32233 (N_32233,N_31808,N_31900);
nor U32234 (N_32234,N_31798,N_31770);
nor U32235 (N_32235,N_31875,N_31969);
nor U32236 (N_32236,N_31872,N_31967);
xnor U32237 (N_32237,N_31944,N_31766);
and U32238 (N_32238,N_31752,N_31909);
xnor U32239 (N_32239,N_31779,N_31893);
and U32240 (N_32240,N_31907,N_31797);
nand U32241 (N_32241,N_31813,N_31967);
nand U32242 (N_32242,N_31899,N_31856);
or U32243 (N_32243,N_31782,N_31833);
and U32244 (N_32244,N_31764,N_31778);
or U32245 (N_32245,N_31822,N_31871);
nand U32246 (N_32246,N_31803,N_31922);
or U32247 (N_32247,N_31950,N_31875);
and U32248 (N_32248,N_31812,N_31800);
xnor U32249 (N_32249,N_31815,N_31897);
nand U32250 (N_32250,N_32198,N_32174);
xor U32251 (N_32251,N_32177,N_32175);
nor U32252 (N_32252,N_32041,N_32133);
nand U32253 (N_32253,N_32124,N_32022);
nor U32254 (N_32254,N_32094,N_32084);
and U32255 (N_32255,N_32113,N_32005);
nand U32256 (N_32256,N_32248,N_32233);
and U32257 (N_32257,N_32047,N_32123);
nor U32258 (N_32258,N_32031,N_32105);
nor U32259 (N_32259,N_32002,N_32213);
nand U32260 (N_32260,N_32115,N_32180);
or U32261 (N_32261,N_32048,N_32173);
and U32262 (N_32262,N_32239,N_32228);
and U32263 (N_32263,N_32076,N_32219);
xor U32264 (N_32264,N_32044,N_32040);
and U32265 (N_32265,N_32085,N_32082);
xor U32266 (N_32266,N_32011,N_32195);
or U32267 (N_32267,N_32103,N_32057);
and U32268 (N_32268,N_32038,N_32088);
nor U32269 (N_32269,N_32182,N_32054);
nand U32270 (N_32270,N_32142,N_32194);
or U32271 (N_32271,N_32092,N_32083);
nand U32272 (N_32272,N_32167,N_32091);
or U32273 (N_32273,N_32161,N_32197);
nor U32274 (N_32274,N_32018,N_32151);
or U32275 (N_32275,N_32106,N_32014);
nor U32276 (N_32276,N_32117,N_32023);
and U32277 (N_32277,N_32099,N_32237);
or U32278 (N_32278,N_32086,N_32060);
xnor U32279 (N_32279,N_32140,N_32049);
nor U32280 (N_32280,N_32216,N_32052);
nand U32281 (N_32281,N_32095,N_32164);
and U32282 (N_32282,N_32204,N_32203);
xor U32283 (N_32283,N_32053,N_32241);
and U32284 (N_32284,N_32129,N_32127);
or U32285 (N_32285,N_32035,N_32188);
xnor U32286 (N_32286,N_32070,N_32066);
or U32287 (N_32287,N_32171,N_32007);
nand U32288 (N_32288,N_32163,N_32074);
and U32289 (N_32289,N_32102,N_32062);
and U32290 (N_32290,N_32211,N_32075);
and U32291 (N_32291,N_32021,N_32242);
or U32292 (N_32292,N_32169,N_32073);
and U32293 (N_32293,N_32110,N_32186);
and U32294 (N_32294,N_32148,N_32134);
nor U32295 (N_32295,N_32019,N_32145);
nor U32296 (N_32296,N_32027,N_32227);
xnor U32297 (N_32297,N_32111,N_32050);
or U32298 (N_32298,N_32039,N_32139);
nor U32299 (N_32299,N_32064,N_32236);
and U32300 (N_32300,N_32138,N_32225);
nand U32301 (N_32301,N_32008,N_32166);
nand U32302 (N_32302,N_32191,N_32079);
and U32303 (N_32303,N_32029,N_32135);
nor U32304 (N_32304,N_32187,N_32012);
nor U32305 (N_32305,N_32097,N_32162);
nand U32306 (N_32306,N_32063,N_32184);
xnor U32307 (N_32307,N_32077,N_32034);
xnor U32308 (N_32308,N_32033,N_32235);
or U32309 (N_32309,N_32128,N_32179);
xor U32310 (N_32310,N_32212,N_32221);
nor U32311 (N_32311,N_32026,N_32232);
xnor U32312 (N_32312,N_32231,N_32156);
or U32313 (N_32313,N_32016,N_32058);
nand U32314 (N_32314,N_32207,N_32183);
and U32315 (N_32315,N_32042,N_32223);
or U32316 (N_32316,N_32116,N_32199);
and U32317 (N_32317,N_32229,N_32065);
xnor U32318 (N_32318,N_32080,N_32037);
nor U32319 (N_32319,N_32176,N_32246);
nand U32320 (N_32320,N_32020,N_32108);
nand U32321 (N_32321,N_32032,N_32170);
nand U32322 (N_32322,N_32205,N_32132);
nand U32323 (N_32323,N_32172,N_32240);
or U32324 (N_32324,N_32004,N_32093);
or U32325 (N_32325,N_32067,N_32226);
xnor U32326 (N_32326,N_32131,N_32192);
and U32327 (N_32327,N_32160,N_32210);
nor U32328 (N_32328,N_32015,N_32071);
and U32329 (N_32329,N_32159,N_32030);
or U32330 (N_32330,N_32100,N_32181);
nand U32331 (N_32331,N_32104,N_32081);
and U32332 (N_32332,N_32096,N_32118);
nand U32333 (N_32333,N_32051,N_32112);
nand U32334 (N_32334,N_32178,N_32234);
nand U32335 (N_32335,N_32120,N_32245);
or U32336 (N_32336,N_32158,N_32013);
or U32337 (N_32337,N_32137,N_32059);
and U32338 (N_32338,N_32168,N_32025);
nand U32339 (N_32339,N_32209,N_32003);
and U32340 (N_32340,N_32202,N_32006);
nor U32341 (N_32341,N_32214,N_32107);
nand U32342 (N_32342,N_32201,N_32153);
nor U32343 (N_32343,N_32024,N_32017);
nor U32344 (N_32344,N_32222,N_32220);
xnor U32345 (N_32345,N_32119,N_32218);
or U32346 (N_32346,N_32149,N_32224);
nor U32347 (N_32347,N_32193,N_32244);
nor U32348 (N_32348,N_32238,N_32101);
xor U32349 (N_32349,N_32001,N_32150);
nand U32350 (N_32350,N_32190,N_32061);
or U32351 (N_32351,N_32185,N_32249);
nor U32352 (N_32352,N_32055,N_32072);
or U32353 (N_32353,N_32230,N_32208);
nor U32354 (N_32354,N_32200,N_32144);
and U32355 (N_32355,N_32068,N_32114);
and U32356 (N_32356,N_32247,N_32165);
and U32357 (N_32357,N_32069,N_32157);
nor U32358 (N_32358,N_32136,N_32109);
nor U32359 (N_32359,N_32056,N_32010);
or U32360 (N_32360,N_32155,N_32146);
and U32361 (N_32361,N_32125,N_32089);
and U32362 (N_32362,N_32215,N_32028);
xnor U32363 (N_32363,N_32098,N_32141);
nand U32364 (N_32364,N_32043,N_32087);
and U32365 (N_32365,N_32130,N_32046);
xnor U32366 (N_32366,N_32143,N_32121);
and U32367 (N_32367,N_32078,N_32122);
nand U32368 (N_32368,N_32152,N_32036);
nor U32369 (N_32369,N_32154,N_32206);
and U32370 (N_32370,N_32090,N_32217);
nor U32371 (N_32371,N_32189,N_32147);
and U32372 (N_32372,N_32000,N_32243);
xor U32373 (N_32373,N_32009,N_32126);
nor U32374 (N_32374,N_32196,N_32045);
or U32375 (N_32375,N_32152,N_32092);
and U32376 (N_32376,N_32091,N_32080);
xor U32377 (N_32377,N_32220,N_32024);
or U32378 (N_32378,N_32148,N_32010);
nand U32379 (N_32379,N_32050,N_32015);
and U32380 (N_32380,N_32002,N_32204);
and U32381 (N_32381,N_32165,N_32112);
or U32382 (N_32382,N_32023,N_32119);
xnor U32383 (N_32383,N_32129,N_32086);
nand U32384 (N_32384,N_32190,N_32068);
and U32385 (N_32385,N_32151,N_32125);
nand U32386 (N_32386,N_32045,N_32028);
nor U32387 (N_32387,N_32216,N_32011);
nor U32388 (N_32388,N_32008,N_32161);
nand U32389 (N_32389,N_32020,N_32062);
or U32390 (N_32390,N_32062,N_32004);
xor U32391 (N_32391,N_32006,N_32100);
or U32392 (N_32392,N_32112,N_32007);
xnor U32393 (N_32393,N_32063,N_32005);
nand U32394 (N_32394,N_32128,N_32184);
xor U32395 (N_32395,N_32203,N_32038);
nor U32396 (N_32396,N_32152,N_32153);
or U32397 (N_32397,N_32130,N_32071);
nand U32398 (N_32398,N_32003,N_32083);
or U32399 (N_32399,N_32067,N_32136);
or U32400 (N_32400,N_32203,N_32003);
and U32401 (N_32401,N_32026,N_32007);
xor U32402 (N_32402,N_32006,N_32086);
nand U32403 (N_32403,N_32104,N_32064);
nor U32404 (N_32404,N_32020,N_32175);
xnor U32405 (N_32405,N_32225,N_32018);
xnor U32406 (N_32406,N_32038,N_32037);
nand U32407 (N_32407,N_32205,N_32173);
xnor U32408 (N_32408,N_32033,N_32068);
nand U32409 (N_32409,N_32149,N_32001);
nor U32410 (N_32410,N_32188,N_32215);
and U32411 (N_32411,N_32046,N_32067);
or U32412 (N_32412,N_32114,N_32205);
or U32413 (N_32413,N_32078,N_32160);
nor U32414 (N_32414,N_32138,N_32093);
nor U32415 (N_32415,N_32239,N_32144);
nand U32416 (N_32416,N_32058,N_32209);
or U32417 (N_32417,N_32153,N_32159);
nand U32418 (N_32418,N_32170,N_32104);
xnor U32419 (N_32419,N_32106,N_32249);
nor U32420 (N_32420,N_32197,N_32244);
nor U32421 (N_32421,N_32221,N_32229);
nand U32422 (N_32422,N_32007,N_32228);
and U32423 (N_32423,N_32224,N_32046);
xor U32424 (N_32424,N_32083,N_32020);
xor U32425 (N_32425,N_32219,N_32174);
xnor U32426 (N_32426,N_32070,N_32203);
xor U32427 (N_32427,N_32198,N_32085);
nor U32428 (N_32428,N_32235,N_32112);
nor U32429 (N_32429,N_32163,N_32245);
or U32430 (N_32430,N_32114,N_32043);
or U32431 (N_32431,N_32115,N_32158);
nand U32432 (N_32432,N_32079,N_32216);
nand U32433 (N_32433,N_32223,N_32017);
and U32434 (N_32434,N_32191,N_32023);
xnor U32435 (N_32435,N_32070,N_32041);
and U32436 (N_32436,N_32208,N_32142);
or U32437 (N_32437,N_32099,N_32112);
and U32438 (N_32438,N_32144,N_32059);
and U32439 (N_32439,N_32014,N_32118);
nand U32440 (N_32440,N_32042,N_32219);
or U32441 (N_32441,N_32015,N_32221);
and U32442 (N_32442,N_32173,N_32054);
xnor U32443 (N_32443,N_32207,N_32177);
xnor U32444 (N_32444,N_32102,N_32034);
nor U32445 (N_32445,N_32148,N_32000);
or U32446 (N_32446,N_32159,N_32051);
and U32447 (N_32447,N_32120,N_32121);
xor U32448 (N_32448,N_32114,N_32169);
nor U32449 (N_32449,N_32022,N_32044);
nand U32450 (N_32450,N_32085,N_32062);
nand U32451 (N_32451,N_32141,N_32111);
nand U32452 (N_32452,N_32217,N_32221);
nor U32453 (N_32453,N_32017,N_32034);
and U32454 (N_32454,N_32024,N_32211);
nor U32455 (N_32455,N_32156,N_32013);
or U32456 (N_32456,N_32031,N_32132);
nor U32457 (N_32457,N_32177,N_32097);
nor U32458 (N_32458,N_32171,N_32137);
nor U32459 (N_32459,N_32194,N_32009);
nand U32460 (N_32460,N_32247,N_32016);
and U32461 (N_32461,N_32169,N_32242);
or U32462 (N_32462,N_32068,N_32184);
nand U32463 (N_32463,N_32086,N_32083);
and U32464 (N_32464,N_32105,N_32171);
xor U32465 (N_32465,N_32047,N_32240);
nor U32466 (N_32466,N_32043,N_32191);
and U32467 (N_32467,N_32088,N_32007);
xnor U32468 (N_32468,N_32167,N_32201);
nor U32469 (N_32469,N_32069,N_32152);
and U32470 (N_32470,N_32079,N_32055);
or U32471 (N_32471,N_32090,N_32035);
nor U32472 (N_32472,N_32172,N_32035);
and U32473 (N_32473,N_32246,N_32111);
or U32474 (N_32474,N_32011,N_32024);
xor U32475 (N_32475,N_32044,N_32204);
nor U32476 (N_32476,N_32247,N_32121);
nand U32477 (N_32477,N_32226,N_32214);
nand U32478 (N_32478,N_32222,N_32079);
nor U32479 (N_32479,N_32041,N_32207);
nand U32480 (N_32480,N_32019,N_32245);
nor U32481 (N_32481,N_32234,N_32035);
xnor U32482 (N_32482,N_32193,N_32202);
and U32483 (N_32483,N_32174,N_32181);
nand U32484 (N_32484,N_32227,N_32057);
nor U32485 (N_32485,N_32141,N_32177);
or U32486 (N_32486,N_32025,N_32046);
or U32487 (N_32487,N_32241,N_32166);
nand U32488 (N_32488,N_32003,N_32031);
xnor U32489 (N_32489,N_32061,N_32154);
xnor U32490 (N_32490,N_32137,N_32181);
xnor U32491 (N_32491,N_32238,N_32047);
xor U32492 (N_32492,N_32050,N_32181);
and U32493 (N_32493,N_32167,N_32171);
nand U32494 (N_32494,N_32199,N_32033);
nand U32495 (N_32495,N_32106,N_32241);
nor U32496 (N_32496,N_32020,N_32070);
nor U32497 (N_32497,N_32061,N_32032);
xor U32498 (N_32498,N_32019,N_32170);
nand U32499 (N_32499,N_32203,N_32000);
or U32500 (N_32500,N_32315,N_32488);
nor U32501 (N_32501,N_32314,N_32265);
or U32502 (N_32502,N_32405,N_32348);
nand U32503 (N_32503,N_32481,N_32310);
nor U32504 (N_32504,N_32261,N_32357);
or U32505 (N_32505,N_32392,N_32394);
or U32506 (N_32506,N_32296,N_32430);
xnor U32507 (N_32507,N_32473,N_32294);
or U32508 (N_32508,N_32479,N_32331);
nor U32509 (N_32509,N_32306,N_32309);
or U32510 (N_32510,N_32381,N_32312);
nor U32511 (N_32511,N_32330,N_32271);
and U32512 (N_32512,N_32295,N_32283);
or U32513 (N_32513,N_32487,N_32354);
and U32514 (N_32514,N_32484,N_32421);
or U32515 (N_32515,N_32439,N_32422);
nand U32516 (N_32516,N_32474,N_32260);
or U32517 (N_32517,N_32471,N_32253);
and U32518 (N_32518,N_32391,N_32403);
and U32519 (N_32519,N_32377,N_32436);
and U32520 (N_32520,N_32302,N_32397);
nand U32521 (N_32521,N_32255,N_32413);
or U32522 (N_32522,N_32390,N_32389);
nand U32523 (N_32523,N_32333,N_32353);
nand U32524 (N_32524,N_32328,N_32399);
nor U32525 (N_32525,N_32451,N_32276);
nand U32526 (N_32526,N_32461,N_32466);
and U32527 (N_32527,N_32257,N_32297);
and U32528 (N_32528,N_32300,N_32457);
xor U32529 (N_32529,N_32303,N_32356);
or U32530 (N_32530,N_32441,N_32432);
nor U32531 (N_32531,N_32320,N_32376);
nand U32532 (N_32532,N_32456,N_32398);
nor U32533 (N_32533,N_32401,N_32367);
xnor U32534 (N_32534,N_32370,N_32292);
nor U32535 (N_32535,N_32277,N_32337);
or U32536 (N_32536,N_32378,N_32339);
and U32537 (N_32537,N_32323,N_32465);
nor U32538 (N_32538,N_32402,N_32268);
xnor U32539 (N_32539,N_32251,N_32485);
and U32540 (N_32540,N_32284,N_32287);
xor U32541 (N_32541,N_32365,N_32388);
xor U32542 (N_32542,N_32301,N_32344);
nor U32543 (N_32543,N_32368,N_32346);
xnor U32544 (N_32544,N_32498,N_32351);
or U32545 (N_32545,N_32273,N_32419);
and U32546 (N_32546,N_32270,N_32290);
and U32547 (N_32547,N_32272,N_32263);
and U32548 (N_32548,N_32431,N_32472);
xor U32549 (N_32549,N_32410,N_32322);
nand U32550 (N_32550,N_32486,N_32452);
xor U32551 (N_32551,N_32293,N_32429);
xnor U32552 (N_32552,N_32475,N_32495);
and U32553 (N_32553,N_32406,N_32454);
xor U32554 (N_32554,N_32449,N_32445);
xnor U32555 (N_32555,N_32308,N_32395);
or U32556 (N_32556,N_32307,N_32332);
xnor U32557 (N_32557,N_32369,N_32400);
xor U32558 (N_32558,N_32476,N_32264);
and U32559 (N_32559,N_32453,N_32443);
or U32560 (N_32560,N_32267,N_32254);
nand U32561 (N_32561,N_32345,N_32349);
nor U32562 (N_32562,N_32440,N_32298);
nor U32563 (N_32563,N_32286,N_32408);
and U32564 (N_32564,N_32380,N_32375);
xnor U32565 (N_32565,N_32499,N_32256);
nor U32566 (N_32566,N_32489,N_32482);
and U32567 (N_32567,N_32359,N_32278);
and U32568 (N_32568,N_32329,N_32347);
nor U32569 (N_32569,N_32423,N_32258);
xor U32570 (N_32570,N_32438,N_32463);
and U32571 (N_32571,N_32496,N_32411);
or U32572 (N_32572,N_32469,N_32478);
nor U32573 (N_32573,N_32274,N_32319);
nand U32574 (N_32574,N_32490,N_32352);
and U32575 (N_32575,N_32424,N_32280);
and U32576 (N_32576,N_32316,N_32304);
nand U32577 (N_32577,N_32382,N_32313);
or U32578 (N_32578,N_32426,N_32363);
xnor U32579 (N_32579,N_32384,N_32420);
or U32580 (N_32580,N_32464,N_32336);
and U32581 (N_32581,N_32358,N_32266);
or U32582 (N_32582,N_32433,N_32362);
nand U32583 (N_32583,N_32493,N_32418);
nand U32584 (N_32584,N_32448,N_32435);
nor U32585 (N_32585,N_32428,N_32317);
xnor U32586 (N_32586,N_32386,N_32415);
nand U32587 (N_32587,N_32447,N_32262);
nor U32588 (N_32588,N_32412,N_32467);
nand U32589 (N_32589,N_32350,N_32446);
and U32590 (N_32590,N_32318,N_32462);
and U32591 (N_32591,N_32342,N_32442);
nor U32592 (N_32592,N_32250,N_32480);
and U32593 (N_32593,N_32355,N_32414);
nor U32594 (N_32594,N_32327,N_32444);
nor U32595 (N_32595,N_32393,N_32364);
nor U32596 (N_32596,N_32379,N_32494);
nand U32597 (N_32597,N_32324,N_32282);
and U32598 (N_32598,N_32477,N_32491);
xor U32599 (N_32599,N_32326,N_32459);
nand U32600 (N_32600,N_32360,N_32468);
and U32601 (N_32601,N_32409,N_32416);
nand U32602 (N_32602,N_32404,N_32299);
nand U32603 (N_32603,N_32269,N_32374);
or U32604 (N_32604,N_32366,N_32483);
nor U32605 (N_32605,N_32334,N_32455);
xnor U32606 (N_32606,N_32281,N_32259);
or U32607 (N_32607,N_32458,N_32371);
nor U32608 (N_32608,N_32289,N_32437);
xor U32609 (N_32609,N_32450,N_32288);
nor U32610 (N_32610,N_32275,N_32372);
and U32611 (N_32611,N_32387,N_32492);
nor U32612 (N_32612,N_32373,N_32341);
nor U32613 (N_32613,N_32252,N_32470);
xor U32614 (N_32614,N_32385,N_32407);
and U32615 (N_32615,N_32335,N_32427);
xor U32616 (N_32616,N_32325,N_32383);
nand U32617 (N_32617,N_32434,N_32305);
or U32618 (N_32618,N_32343,N_32425);
nand U32619 (N_32619,N_32361,N_32497);
and U32620 (N_32620,N_32311,N_32340);
nand U32621 (N_32621,N_32279,N_32285);
or U32622 (N_32622,N_32396,N_32417);
and U32623 (N_32623,N_32338,N_32321);
and U32624 (N_32624,N_32460,N_32291);
and U32625 (N_32625,N_32338,N_32340);
and U32626 (N_32626,N_32315,N_32396);
nor U32627 (N_32627,N_32351,N_32271);
or U32628 (N_32628,N_32457,N_32368);
and U32629 (N_32629,N_32436,N_32472);
xor U32630 (N_32630,N_32379,N_32394);
and U32631 (N_32631,N_32466,N_32460);
xnor U32632 (N_32632,N_32342,N_32447);
and U32633 (N_32633,N_32427,N_32322);
and U32634 (N_32634,N_32338,N_32347);
and U32635 (N_32635,N_32476,N_32326);
or U32636 (N_32636,N_32336,N_32321);
xor U32637 (N_32637,N_32479,N_32334);
nand U32638 (N_32638,N_32376,N_32386);
xor U32639 (N_32639,N_32341,N_32424);
nor U32640 (N_32640,N_32427,N_32413);
nor U32641 (N_32641,N_32334,N_32489);
nand U32642 (N_32642,N_32392,N_32391);
nor U32643 (N_32643,N_32320,N_32299);
or U32644 (N_32644,N_32489,N_32476);
and U32645 (N_32645,N_32262,N_32485);
nand U32646 (N_32646,N_32459,N_32445);
nand U32647 (N_32647,N_32354,N_32453);
xor U32648 (N_32648,N_32436,N_32491);
or U32649 (N_32649,N_32469,N_32382);
and U32650 (N_32650,N_32490,N_32442);
nor U32651 (N_32651,N_32335,N_32479);
or U32652 (N_32652,N_32364,N_32409);
and U32653 (N_32653,N_32386,N_32481);
nor U32654 (N_32654,N_32283,N_32433);
xnor U32655 (N_32655,N_32474,N_32427);
and U32656 (N_32656,N_32451,N_32350);
or U32657 (N_32657,N_32259,N_32492);
nor U32658 (N_32658,N_32397,N_32380);
nor U32659 (N_32659,N_32443,N_32446);
and U32660 (N_32660,N_32310,N_32461);
or U32661 (N_32661,N_32324,N_32394);
or U32662 (N_32662,N_32363,N_32471);
nor U32663 (N_32663,N_32326,N_32253);
and U32664 (N_32664,N_32418,N_32487);
or U32665 (N_32665,N_32412,N_32446);
nand U32666 (N_32666,N_32346,N_32423);
nor U32667 (N_32667,N_32414,N_32426);
xnor U32668 (N_32668,N_32361,N_32481);
or U32669 (N_32669,N_32480,N_32295);
nand U32670 (N_32670,N_32291,N_32317);
or U32671 (N_32671,N_32394,N_32495);
or U32672 (N_32672,N_32494,N_32421);
and U32673 (N_32673,N_32315,N_32348);
and U32674 (N_32674,N_32318,N_32302);
xnor U32675 (N_32675,N_32398,N_32386);
or U32676 (N_32676,N_32352,N_32258);
nor U32677 (N_32677,N_32426,N_32464);
nand U32678 (N_32678,N_32379,N_32332);
and U32679 (N_32679,N_32285,N_32452);
xor U32680 (N_32680,N_32352,N_32457);
nor U32681 (N_32681,N_32331,N_32357);
and U32682 (N_32682,N_32316,N_32496);
nand U32683 (N_32683,N_32284,N_32331);
and U32684 (N_32684,N_32446,N_32307);
nand U32685 (N_32685,N_32489,N_32314);
or U32686 (N_32686,N_32437,N_32287);
nand U32687 (N_32687,N_32419,N_32305);
xnor U32688 (N_32688,N_32457,N_32334);
xor U32689 (N_32689,N_32338,N_32438);
or U32690 (N_32690,N_32347,N_32282);
nor U32691 (N_32691,N_32471,N_32372);
xor U32692 (N_32692,N_32454,N_32305);
nand U32693 (N_32693,N_32410,N_32483);
xor U32694 (N_32694,N_32288,N_32267);
nand U32695 (N_32695,N_32407,N_32337);
or U32696 (N_32696,N_32491,N_32360);
nor U32697 (N_32697,N_32286,N_32297);
and U32698 (N_32698,N_32325,N_32470);
nor U32699 (N_32699,N_32269,N_32372);
nand U32700 (N_32700,N_32441,N_32326);
or U32701 (N_32701,N_32431,N_32434);
xor U32702 (N_32702,N_32316,N_32469);
xor U32703 (N_32703,N_32269,N_32420);
nor U32704 (N_32704,N_32458,N_32465);
and U32705 (N_32705,N_32417,N_32437);
or U32706 (N_32706,N_32284,N_32487);
and U32707 (N_32707,N_32431,N_32267);
nor U32708 (N_32708,N_32279,N_32411);
nand U32709 (N_32709,N_32257,N_32295);
or U32710 (N_32710,N_32345,N_32311);
xnor U32711 (N_32711,N_32383,N_32449);
or U32712 (N_32712,N_32321,N_32320);
nand U32713 (N_32713,N_32284,N_32457);
or U32714 (N_32714,N_32314,N_32289);
nor U32715 (N_32715,N_32396,N_32306);
xor U32716 (N_32716,N_32285,N_32293);
nand U32717 (N_32717,N_32339,N_32372);
xnor U32718 (N_32718,N_32468,N_32382);
xnor U32719 (N_32719,N_32259,N_32316);
nor U32720 (N_32720,N_32488,N_32446);
or U32721 (N_32721,N_32367,N_32393);
or U32722 (N_32722,N_32462,N_32362);
nor U32723 (N_32723,N_32377,N_32467);
or U32724 (N_32724,N_32385,N_32340);
or U32725 (N_32725,N_32268,N_32337);
nor U32726 (N_32726,N_32301,N_32434);
xnor U32727 (N_32727,N_32360,N_32442);
nor U32728 (N_32728,N_32321,N_32385);
or U32729 (N_32729,N_32409,N_32456);
and U32730 (N_32730,N_32462,N_32405);
nand U32731 (N_32731,N_32458,N_32415);
or U32732 (N_32732,N_32252,N_32294);
nand U32733 (N_32733,N_32377,N_32346);
nand U32734 (N_32734,N_32270,N_32288);
and U32735 (N_32735,N_32346,N_32373);
or U32736 (N_32736,N_32310,N_32250);
xor U32737 (N_32737,N_32318,N_32402);
xor U32738 (N_32738,N_32397,N_32342);
nand U32739 (N_32739,N_32328,N_32262);
nor U32740 (N_32740,N_32466,N_32307);
or U32741 (N_32741,N_32411,N_32499);
xor U32742 (N_32742,N_32298,N_32410);
xnor U32743 (N_32743,N_32261,N_32372);
nor U32744 (N_32744,N_32402,N_32380);
nor U32745 (N_32745,N_32383,N_32343);
nor U32746 (N_32746,N_32375,N_32269);
xor U32747 (N_32747,N_32315,N_32394);
or U32748 (N_32748,N_32399,N_32451);
and U32749 (N_32749,N_32358,N_32342);
xnor U32750 (N_32750,N_32560,N_32648);
nand U32751 (N_32751,N_32680,N_32519);
nor U32752 (N_32752,N_32702,N_32599);
and U32753 (N_32753,N_32646,N_32624);
and U32754 (N_32754,N_32647,N_32704);
or U32755 (N_32755,N_32693,N_32654);
and U32756 (N_32756,N_32507,N_32721);
nand U32757 (N_32757,N_32649,N_32720);
nor U32758 (N_32758,N_32736,N_32516);
nor U32759 (N_32759,N_32617,N_32746);
and U32760 (N_32760,N_32522,N_32542);
nand U32761 (N_32761,N_32668,N_32568);
or U32762 (N_32762,N_32638,N_32745);
nand U32763 (N_32763,N_32734,N_32643);
and U32764 (N_32764,N_32652,N_32714);
and U32765 (N_32765,N_32558,N_32637);
or U32766 (N_32766,N_32500,N_32656);
and U32767 (N_32767,N_32641,N_32605);
and U32768 (N_32768,N_32583,N_32505);
xor U32769 (N_32769,N_32604,N_32608);
nor U32770 (N_32770,N_32689,N_32694);
nand U32771 (N_32771,N_32596,N_32703);
nand U32772 (N_32772,N_32574,N_32582);
or U32773 (N_32773,N_32743,N_32662);
xor U32774 (N_32774,N_32576,N_32666);
nor U32775 (N_32775,N_32545,N_32547);
nor U32776 (N_32776,N_32521,N_32747);
nand U32777 (N_32777,N_32523,N_32526);
nand U32778 (N_32778,N_32731,N_32667);
nor U32779 (N_32779,N_32612,N_32715);
and U32780 (N_32780,N_32629,N_32534);
nor U32781 (N_32781,N_32517,N_32506);
or U32782 (N_32782,N_32735,N_32711);
and U32783 (N_32783,N_32592,N_32581);
nand U32784 (N_32784,N_32690,N_32630);
and U32785 (N_32785,N_32540,N_32595);
nor U32786 (N_32786,N_32676,N_32537);
xnor U32787 (N_32787,N_32564,N_32511);
xnor U32788 (N_32788,N_32586,N_32610);
and U32789 (N_32789,N_32679,N_32525);
nor U32790 (N_32790,N_32509,N_32644);
nor U32791 (N_32791,N_32744,N_32632);
or U32792 (N_32792,N_32673,N_32544);
nor U32793 (N_32793,N_32614,N_32728);
xnor U32794 (N_32794,N_32657,N_32520);
nand U32795 (N_32795,N_32688,N_32619);
or U32796 (N_32796,N_32636,N_32671);
nor U32797 (N_32797,N_32699,N_32645);
nor U32798 (N_32798,N_32623,N_32600);
xor U32799 (N_32799,N_32672,N_32732);
nand U32800 (N_32800,N_32561,N_32513);
xnor U32801 (N_32801,N_32567,N_32719);
xor U32802 (N_32802,N_32741,N_32627);
nor U32803 (N_32803,N_32527,N_32712);
nor U32804 (N_32804,N_32682,N_32551);
nand U32805 (N_32805,N_32524,N_32669);
nor U32806 (N_32806,N_32572,N_32622);
xnor U32807 (N_32807,N_32691,N_32543);
nor U32808 (N_32808,N_32739,N_32661);
and U32809 (N_32809,N_32740,N_32510);
or U32810 (N_32810,N_32615,N_32569);
and U32811 (N_32811,N_32594,N_32566);
nand U32812 (N_32812,N_32609,N_32503);
or U32813 (N_32813,N_32579,N_32707);
and U32814 (N_32814,N_32722,N_32737);
nand U32815 (N_32815,N_32665,N_32738);
nor U32816 (N_32816,N_32710,N_32742);
nor U32817 (N_32817,N_32642,N_32628);
xor U32818 (N_32818,N_32531,N_32607);
nand U32819 (N_32819,N_32602,N_32724);
nor U32820 (N_32820,N_32550,N_32723);
nor U32821 (N_32821,N_32621,N_32611);
nor U32822 (N_32822,N_32591,N_32650);
or U32823 (N_32823,N_32530,N_32613);
nand U32824 (N_32824,N_32683,N_32565);
nor U32825 (N_32825,N_32557,N_32634);
nor U32826 (N_32826,N_32539,N_32589);
and U32827 (N_32827,N_32580,N_32549);
and U32828 (N_32828,N_32559,N_32606);
nor U32829 (N_32829,N_32562,N_32555);
or U32830 (N_32830,N_32514,N_32696);
nand U32831 (N_32831,N_32501,N_32651);
nor U32832 (N_32832,N_32515,N_32546);
xnor U32833 (N_32833,N_32705,N_32674);
and U32834 (N_32834,N_32571,N_32620);
and U32835 (N_32835,N_32697,N_32670);
nor U32836 (N_32836,N_32508,N_32590);
nor U32837 (N_32837,N_32597,N_32664);
xnor U32838 (N_32838,N_32512,N_32584);
or U32839 (N_32839,N_32686,N_32631);
xnor U32840 (N_32840,N_32533,N_32716);
nor U32841 (N_32841,N_32718,N_32626);
or U32842 (N_32842,N_32733,N_32535);
nor U32843 (N_32843,N_32695,N_32577);
nand U32844 (N_32844,N_32563,N_32726);
and U32845 (N_32845,N_32659,N_32598);
xor U32846 (N_32846,N_32625,N_32633);
nand U32847 (N_32847,N_32713,N_32504);
xor U32848 (N_32848,N_32616,N_32552);
nor U32849 (N_32849,N_32677,N_32655);
or U32850 (N_32850,N_32529,N_32685);
nand U32851 (N_32851,N_32578,N_32587);
and U32852 (N_32852,N_32681,N_32729);
or U32853 (N_32853,N_32725,N_32556);
nor U32854 (N_32854,N_32570,N_32502);
or U32855 (N_32855,N_32692,N_32640);
xor U32856 (N_32856,N_32687,N_32698);
xnor U32857 (N_32857,N_32554,N_32678);
nand U32858 (N_32858,N_32749,N_32575);
xor U32859 (N_32859,N_32585,N_32553);
nor U32860 (N_32860,N_32730,N_32601);
xor U32861 (N_32861,N_32708,N_32588);
nand U32862 (N_32862,N_32701,N_32675);
and U32863 (N_32863,N_32536,N_32573);
and U32864 (N_32864,N_32653,N_32700);
xor U32865 (N_32865,N_32603,N_32639);
and U32866 (N_32866,N_32541,N_32727);
and U32867 (N_32867,N_32717,N_32706);
and U32868 (N_32868,N_32548,N_32618);
nor U32869 (N_32869,N_32684,N_32660);
nor U32870 (N_32870,N_32663,N_32593);
nor U32871 (N_32871,N_32748,N_32538);
and U32872 (N_32872,N_32532,N_32518);
and U32873 (N_32873,N_32528,N_32709);
xnor U32874 (N_32874,N_32658,N_32635);
nor U32875 (N_32875,N_32642,N_32612);
nand U32876 (N_32876,N_32732,N_32638);
xnor U32877 (N_32877,N_32650,N_32526);
and U32878 (N_32878,N_32652,N_32684);
nor U32879 (N_32879,N_32637,N_32510);
nand U32880 (N_32880,N_32671,N_32723);
xnor U32881 (N_32881,N_32708,N_32729);
or U32882 (N_32882,N_32680,N_32510);
nor U32883 (N_32883,N_32606,N_32508);
nand U32884 (N_32884,N_32668,N_32717);
nand U32885 (N_32885,N_32500,N_32601);
xnor U32886 (N_32886,N_32547,N_32520);
nand U32887 (N_32887,N_32561,N_32607);
and U32888 (N_32888,N_32656,N_32629);
nor U32889 (N_32889,N_32540,N_32656);
xnor U32890 (N_32890,N_32647,N_32678);
nor U32891 (N_32891,N_32540,N_32747);
nor U32892 (N_32892,N_32613,N_32575);
or U32893 (N_32893,N_32691,N_32722);
xnor U32894 (N_32894,N_32708,N_32630);
and U32895 (N_32895,N_32573,N_32643);
nor U32896 (N_32896,N_32617,N_32640);
or U32897 (N_32897,N_32735,N_32639);
nand U32898 (N_32898,N_32588,N_32628);
xnor U32899 (N_32899,N_32512,N_32549);
nor U32900 (N_32900,N_32593,N_32517);
nor U32901 (N_32901,N_32641,N_32579);
nand U32902 (N_32902,N_32663,N_32665);
xor U32903 (N_32903,N_32745,N_32711);
xnor U32904 (N_32904,N_32730,N_32693);
or U32905 (N_32905,N_32650,N_32642);
or U32906 (N_32906,N_32610,N_32612);
or U32907 (N_32907,N_32569,N_32590);
nor U32908 (N_32908,N_32683,N_32525);
and U32909 (N_32909,N_32654,N_32675);
or U32910 (N_32910,N_32718,N_32577);
nand U32911 (N_32911,N_32541,N_32637);
and U32912 (N_32912,N_32536,N_32694);
nor U32913 (N_32913,N_32606,N_32634);
xor U32914 (N_32914,N_32634,N_32625);
or U32915 (N_32915,N_32529,N_32520);
nor U32916 (N_32916,N_32592,N_32593);
and U32917 (N_32917,N_32623,N_32687);
or U32918 (N_32918,N_32527,N_32550);
nor U32919 (N_32919,N_32731,N_32714);
xnor U32920 (N_32920,N_32515,N_32675);
or U32921 (N_32921,N_32591,N_32523);
nor U32922 (N_32922,N_32639,N_32510);
and U32923 (N_32923,N_32528,N_32727);
xnor U32924 (N_32924,N_32672,N_32529);
or U32925 (N_32925,N_32714,N_32738);
or U32926 (N_32926,N_32690,N_32564);
nor U32927 (N_32927,N_32671,N_32725);
nand U32928 (N_32928,N_32581,N_32727);
and U32929 (N_32929,N_32651,N_32645);
and U32930 (N_32930,N_32554,N_32616);
nor U32931 (N_32931,N_32591,N_32534);
xnor U32932 (N_32932,N_32580,N_32519);
xnor U32933 (N_32933,N_32688,N_32506);
nand U32934 (N_32934,N_32618,N_32579);
nor U32935 (N_32935,N_32706,N_32740);
nor U32936 (N_32936,N_32530,N_32722);
nor U32937 (N_32937,N_32653,N_32642);
xnor U32938 (N_32938,N_32623,N_32564);
nand U32939 (N_32939,N_32627,N_32636);
and U32940 (N_32940,N_32639,N_32517);
nand U32941 (N_32941,N_32631,N_32521);
and U32942 (N_32942,N_32682,N_32704);
nor U32943 (N_32943,N_32635,N_32598);
xor U32944 (N_32944,N_32666,N_32522);
nor U32945 (N_32945,N_32681,N_32573);
and U32946 (N_32946,N_32651,N_32731);
nor U32947 (N_32947,N_32508,N_32540);
nor U32948 (N_32948,N_32529,N_32648);
or U32949 (N_32949,N_32744,N_32739);
nor U32950 (N_32950,N_32516,N_32680);
nor U32951 (N_32951,N_32547,N_32706);
xnor U32952 (N_32952,N_32656,N_32534);
and U32953 (N_32953,N_32640,N_32508);
nand U32954 (N_32954,N_32742,N_32642);
nand U32955 (N_32955,N_32690,N_32738);
and U32956 (N_32956,N_32567,N_32594);
or U32957 (N_32957,N_32637,N_32703);
nand U32958 (N_32958,N_32576,N_32536);
nand U32959 (N_32959,N_32633,N_32686);
xor U32960 (N_32960,N_32639,N_32702);
xnor U32961 (N_32961,N_32560,N_32659);
xnor U32962 (N_32962,N_32544,N_32583);
nor U32963 (N_32963,N_32693,N_32586);
nor U32964 (N_32964,N_32561,N_32695);
nor U32965 (N_32965,N_32591,N_32611);
xnor U32966 (N_32966,N_32647,N_32608);
xor U32967 (N_32967,N_32597,N_32530);
and U32968 (N_32968,N_32707,N_32534);
nand U32969 (N_32969,N_32679,N_32528);
nor U32970 (N_32970,N_32513,N_32666);
xnor U32971 (N_32971,N_32739,N_32627);
xor U32972 (N_32972,N_32681,N_32627);
nand U32973 (N_32973,N_32557,N_32514);
xnor U32974 (N_32974,N_32680,N_32545);
xor U32975 (N_32975,N_32513,N_32738);
xor U32976 (N_32976,N_32720,N_32665);
and U32977 (N_32977,N_32519,N_32740);
and U32978 (N_32978,N_32535,N_32718);
nand U32979 (N_32979,N_32580,N_32633);
nor U32980 (N_32980,N_32592,N_32702);
nand U32981 (N_32981,N_32599,N_32584);
xnor U32982 (N_32982,N_32536,N_32607);
nand U32983 (N_32983,N_32547,N_32742);
nand U32984 (N_32984,N_32698,N_32601);
xnor U32985 (N_32985,N_32738,N_32510);
nor U32986 (N_32986,N_32513,N_32720);
and U32987 (N_32987,N_32511,N_32589);
or U32988 (N_32988,N_32571,N_32608);
nor U32989 (N_32989,N_32562,N_32680);
nor U32990 (N_32990,N_32526,N_32715);
nor U32991 (N_32991,N_32615,N_32643);
xor U32992 (N_32992,N_32703,N_32554);
or U32993 (N_32993,N_32741,N_32691);
or U32994 (N_32994,N_32537,N_32732);
nor U32995 (N_32995,N_32501,N_32524);
xor U32996 (N_32996,N_32591,N_32726);
and U32997 (N_32997,N_32522,N_32738);
nor U32998 (N_32998,N_32549,N_32710);
nand U32999 (N_32999,N_32720,N_32700);
nand U33000 (N_33000,N_32792,N_32922);
or U33001 (N_33001,N_32951,N_32848);
xnor U33002 (N_33002,N_32941,N_32911);
xor U33003 (N_33003,N_32884,N_32919);
xor U33004 (N_33004,N_32791,N_32956);
xnor U33005 (N_33005,N_32770,N_32809);
nand U33006 (N_33006,N_32962,N_32855);
nor U33007 (N_33007,N_32983,N_32984);
nor U33008 (N_33008,N_32771,N_32873);
xor U33009 (N_33009,N_32830,N_32868);
nand U33010 (N_33010,N_32981,N_32892);
and U33011 (N_33011,N_32938,N_32969);
nor U33012 (N_33012,N_32876,N_32939);
xnor U33013 (N_33013,N_32993,N_32977);
xor U33014 (N_33014,N_32942,N_32944);
nand U33015 (N_33015,N_32997,N_32880);
xor U33016 (N_33016,N_32856,N_32989);
nor U33017 (N_33017,N_32865,N_32821);
xnor U33018 (N_33018,N_32839,N_32979);
xor U33019 (N_33019,N_32841,N_32847);
or U33020 (N_33020,N_32998,N_32804);
or U33021 (N_33021,N_32886,N_32846);
nand U33022 (N_33022,N_32808,N_32759);
xnor U33023 (N_33023,N_32888,N_32843);
or U33024 (N_33024,N_32751,N_32796);
nor U33025 (N_33025,N_32906,N_32964);
nor U33026 (N_33026,N_32899,N_32769);
or U33027 (N_33027,N_32918,N_32940);
xnor U33028 (N_33028,N_32845,N_32913);
nor U33029 (N_33029,N_32975,N_32974);
nand U33030 (N_33030,N_32858,N_32932);
nand U33031 (N_33031,N_32812,N_32823);
nand U33032 (N_33032,N_32836,N_32768);
and U33033 (N_33033,N_32915,N_32774);
nor U33034 (N_33034,N_32953,N_32832);
and U33035 (N_33035,N_32773,N_32948);
and U33036 (N_33036,N_32816,N_32784);
or U33037 (N_33037,N_32766,N_32959);
xnor U33038 (N_33038,N_32780,N_32863);
nand U33039 (N_33039,N_32963,N_32924);
or U33040 (N_33040,N_32966,N_32870);
or U33041 (N_33041,N_32897,N_32807);
nand U33042 (N_33042,N_32752,N_32901);
nand U33043 (N_33043,N_32793,N_32782);
and U33044 (N_33044,N_32900,N_32970);
nor U33045 (N_33045,N_32840,N_32801);
and U33046 (N_33046,N_32795,N_32775);
nand U33047 (N_33047,N_32799,N_32838);
nand U33048 (N_33048,N_32849,N_32937);
xor U33049 (N_33049,N_32862,N_32947);
and U33050 (N_33050,N_32776,N_32827);
and U33051 (N_33051,N_32869,N_32824);
xor U33052 (N_33052,N_32999,N_32767);
xor U33053 (N_33053,N_32916,N_32786);
and U33054 (N_33054,N_32788,N_32810);
and U33055 (N_33055,N_32905,N_32831);
or U33056 (N_33056,N_32995,N_32756);
nor U33057 (N_33057,N_32978,N_32930);
nand U33058 (N_33058,N_32850,N_32898);
or U33059 (N_33059,N_32936,N_32895);
nand U33060 (N_33060,N_32835,N_32760);
nand U33061 (N_33061,N_32990,N_32802);
and U33062 (N_33062,N_32750,N_32933);
or U33063 (N_33063,N_32829,N_32887);
and U33064 (N_33064,N_32891,N_32878);
and U33065 (N_33065,N_32864,N_32777);
or U33066 (N_33066,N_32958,N_32928);
or U33067 (N_33067,N_32822,N_32935);
nand U33068 (N_33068,N_32991,N_32967);
nand U33069 (N_33069,N_32996,N_32971);
nand U33070 (N_33070,N_32753,N_32787);
nand U33071 (N_33071,N_32805,N_32894);
and U33072 (N_33072,N_32762,N_32818);
nand U33073 (N_33073,N_32949,N_32854);
or U33074 (N_33074,N_32893,N_32754);
nand U33075 (N_33075,N_32968,N_32857);
or U33076 (N_33076,N_32778,N_32833);
xor U33077 (N_33077,N_32758,N_32817);
nand U33078 (N_33078,N_32955,N_32912);
or U33079 (N_33079,N_32772,N_32851);
and U33080 (N_33080,N_32881,N_32992);
nor U33081 (N_33081,N_32779,N_32790);
or U33082 (N_33082,N_32903,N_32781);
xor U33083 (N_33083,N_32965,N_32844);
and U33084 (N_33084,N_32837,N_32872);
nor U33085 (N_33085,N_32946,N_32934);
xor U33086 (N_33086,N_32755,N_32879);
and U33087 (N_33087,N_32976,N_32763);
and U33088 (N_33088,N_32877,N_32811);
and U33089 (N_33089,N_32890,N_32828);
nor U33090 (N_33090,N_32859,N_32907);
or U33091 (N_33091,N_32757,N_32783);
xor U33092 (N_33092,N_32853,N_32961);
and U33093 (N_33093,N_32874,N_32798);
or U33094 (N_33094,N_32943,N_32926);
and U33095 (N_33095,N_32909,N_32960);
xnor U33096 (N_33096,N_32794,N_32819);
and U33097 (N_33097,N_32925,N_32931);
or U33098 (N_33098,N_32866,N_32908);
nand U33099 (N_33099,N_32834,N_32914);
xor U33100 (N_33100,N_32885,N_32950);
xnor U33101 (N_33101,N_32921,N_32761);
nand U33102 (N_33102,N_32987,N_32883);
or U33103 (N_33103,N_32986,N_32882);
nand U33104 (N_33104,N_32871,N_32860);
or U33105 (N_33105,N_32826,N_32972);
nor U33106 (N_33106,N_32957,N_32952);
or U33107 (N_33107,N_32994,N_32789);
xnor U33108 (N_33108,N_32896,N_32889);
nor U33109 (N_33109,N_32814,N_32927);
nand U33110 (N_33110,N_32980,N_32920);
xnor U33111 (N_33111,N_32945,N_32797);
nand U33112 (N_33112,N_32875,N_32813);
nand U33113 (N_33113,N_32815,N_32867);
or U33114 (N_33114,N_32764,N_32954);
nand U33115 (N_33115,N_32910,N_32803);
nand U33116 (N_33116,N_32806,N_32785);
nand U33117 (N_33117,N_32825,N_32985);
or U33118 (N_33118,N_32904,N_32861);
or U33119 (N_33119,N_32917,N_32800);
and U33120 (N_33120,N_32929,N_32973);
and U33121 (N_33121,N_32902,N_32852);
nor U33122 (N_33122,N_32923,N_32842);
nor U33123 (N_33123,N_32982,N_32765);
nand U33124 (N_33124,N_32820,N_32988);
nor U33125 (N_33125,N_32984,N_32919);
nand U33126 (N_33126,N_32984,N_32900);
nand U33127 (N_33127,N_32938,N_32984);
nor U33128 (N_33128,N_32977,N_32953);
nor U33129 (N_33129,N_32833,N_32931);
xnor U33130 (N_33130,N_32857,N_32805);
nand U33131 (N_33131,N_32995,N_32963);
nand U33132 (N_33132,N_32783,N_32981);
xor U33133 (N_33133,N_32956,N_32977);
and U33134 (N_33134,N_32892,N_32818);
xnor U33135 (N_33135,N_32888,N_32976);
or U33136 (N_33136,N_32874,N_32773);
nor U33137 (N_33137,N_32901,N_32974);
nor U33138 (N_33138,N_32765,N_32971);
and U33139 (N_33139,N_32948,N_32821);
xnor U33140 (N_33140,N_32754,N_32976);
and U33141 (N_33141,N_32906,N_32938);
or U33142 (N_33142,N_32811,N_32999);
and U33143 (N_33143,N_32758,N_32829);
or U33144 (N_33144,N_32994,N_32981);
nor U33145 (N_33145,N_32795,N_32894);
xor U33146 (N_33146,N_32813,N_32897);
xnor U33147 (N_33147,N_32877,N_32879);
and U33148 (N_33148,N_32794,N_32915);
or U33149 (N_33149,N_32770,N_32757);
nand U33150 (N_33150,N_32870,N_32903);
and U33151 (N_33151,N_32870,N_32934);
nor U33152 (N_33152,N_32994,N_32946);
or U33153 (N_33153,N_32978,N_32795);
xnor U33154 (N_33154,N_32812,N_32863);
nor U33155 (N_33155,N_32884,N_32860);
nor U33156 (N_33156,N_32765,N_32831);
nand U33157 (N_33157,N_32922,N_32942);
nor U33158 (N_33158,N_32783,N_32884);
xnor U33159 (N_33159,N_32855,N_32845);
nor U33160 (N_33160,N_32941,N_32810);
and U33161 (N_33161,N_32832,N_32840);
or U33162 (N_33162,N_32932,N_32865);
xnor U33163 (N_33163,N_32784,N_32915);
or U33164 (N_33164,N_32957,N_32961);
or U33165 (N_33165,N_32768,N_32881);
and U33166 (N_33166,N_32992,N_32951);
or U33167 (N_33167,N_32982,N_32862);
nor U33168 (N_33168,N_32826,N_32996);
nand U33169 (N_33169,N_32988,N_32911);
xnor U33170 (N_33170,N_32800,N_32781);
xor U33171 (N_33171,N_32901,N_32996);
nor U33172 (N_33172,N_32793,N_32873);
nand U33173 (N_33173,N_32939,N_32947);
and U33174 (N_33174,N_32963,N_32951);
or U33175 (N_33175,N_32806,N_32862);
nor U33176 (N_33176,N_32981,N_32922);
xor U33177 (N_33177,N_32994,N_32885);
nor U33178 (N_33178,N_32863,N_32883);
nand U33179 (N_33179,N_32757,N_32812);
nor U33180 (N_33180,N_32757,N_32971);
nor U33181 (N_33181,N_32903,N_32794);
and U33182 (N_33182,N_32992,N_32910);
nor U33183 (N_33183,N_32919,N_32777);
nand U33184 (N_33184,N_32943,N_32973);
xor U33185 (N_33185,N_32979,N_32755);
nor U33186 (N_33186,N_32943,N_32778);
and U33187 (N_33187,N_32963,N_32803);
and U33188 (N_33188,N_32946,N_32849);
xor U33189 (N_33189,N_32924,N_32758);
nand U33190 (N_33190,N_32839,N_32973);
and U33191 (N_33191,N_32964,N_32819);
nor U33192 (N_33192,N_32799,N_32919);
xor U33193 (N_33193,N_32942,N_32798);
nand U33194 (N_33194,N_32807,N_32923);
nand U33195 (N_33195,N_32923,N_32870);
xor U33196 (N_33196,N_32904,N_32752);
xor U33197 (N_33197,N_32874,N_32964);
nand U33198 (N_33198,N_32840,N_32816);
nand U33199 (N_33199,N_32977,N_32859);
xor U33200 (N_33200,N_32903,N_32890);
or U33201 (N_33201,N_32836,N_32770);
or U33202 (N_33202,N_32801,N_32861);
nand U33203 (N_33203,N_32882,N_32889);
and U33204 (N_33204,N_32884,N_32990);
and U33205 (N_33205,N_32865,N_32909);
nand U33206 (N_33206,N_32839,N_32898);
or U33207 (N_33207,N_32958,N_32813);
nand U33208 (N_33208,N_32865,N_32809);
nand U33209 (N_33209,N_32996,N_32995);
xnor U33210 (N_33210,N_32997,N_32965);
nand U33211 (N_33211,N_32904,N_32766);
nand U33212 (N_33212,N_32780,N_32966);
xnor U33213 (N_33213,N_32920,N_32869);
xnor U33214 (N_33214,N_32786,N_32854);
nor U33215 (N_33215,N_32978,N_32840);
nor U33216 (N_33216,N_32883,N_32791);
xnor U33217 (N_33217,N_32839,N_32910);
and U33218 (N_33218,N_32778,N_32869);
nor U33219 (N_33219,N_32847,N_32797);
or U33220 (N_33220,N_32767,N_32923);
or U33221 (N_33221,N_32829,N_32855);
and U33222 (N_33222,N_32846,N_32773);
xnor U33223 (N_33223,N_32786,N_32904);
nand U33224 (N_33224,N_32845,N_32812);
or U33225 (N_33225,N_32848,N_32900);
nor U33226 (N_33226,N_32930,N_32778);
nor U33227 (N_33227,N_32809,N_32861);
and U33228 (N_33228,N_32987,N_32972);
nor U33229 (N_33229,N_32973,N_32887);
xnor U33230 (N_33230,N_32913,N_32811);
nor U33231 (N_33231,N_32756,N_32855);
xor U33232 (N_33232,N_32773,N_32822);
nand U33233 (N_33233,N_32944,N_32830);
nand U33234 (N_33234,N_32818,N_32810);
nand U33235 (N_33235,N_32800,N_32970);
and U33236 (N_33236,N_32912,N_32882);
nor U33237 (N_33237,N_32932,N_32761);
xnor U33238 (N_33238,N_32930,N_32843);
nand U33239 (N_33239,N_32782,N_32778);
or U33240 (N_33240,N_32754,N_32899);
or U33241 (N_33241,N_32923,N_32941);
nor U33242 (N_33242,N_32991,N_32868);
xor U33243 (N_33243,N_32864,N_32984);
and U33244 (N_33244,N_32975,N_32966);
or U33245 (N_33245,N_32774,N_32839);
nand U33246 (N_33246,N_32896,N_32916);
and U33247 (N_33247,N_32793,N_32822);
and U33248 (N_33248,N_32908,N_32752);
and U33249 (N_33249,N_32995,N_32899);
nand U33250 (N_33250,N_33244,N_33228);
nand U33251 (N_33251,N_33160,N_33157);
nor U33252 (N_33252,N_33084,N_33122);
xor U33253 (N_33253,N_33167,N_33012);
nand U33254 (N_33254,N_33184,N_33159);
or U33255 (N_33255,N_33227,N_33182);
nor U33256 (N_33256,N_33105,N_33110);
nand U33257 (N_33257,N_33223,N_33241);
nand U33258 (N_33258,N_33156,N_33007);
xor U33259 (N_33259,N_33031,N_33002);
and U33260 (N_33260,N_33225,N_33240);
nor U33261 (N_33261,N_33090,N_33045);
nor U33262 (N_33262,N_33044,N_33246);
nand U33263 (N_33263,N_33153,N_33216);
nand U33264 (N_33264,N_33163,N_33118);
nand U33265 (N_33265,N_33239,N_33181);
xor U33266 (N_33266,N_33088,N_33172);
or U33267 (N_33267,N_33024,N_33069);
or U33268 (N_33268,N_33248,N_33104);
nand U33269 (N_33269,N_33029,N_33186);
or U33270 (N_33270,N_33130,N_33095);
nor U33271 (N_33271,N_33131,N_33132);
nor U33272 (N_33272,N_33196,N_33198);
nor U33273 (N_33273,N_33036,N_33112);
and U33274 (N_33274,N_33201,N_33193);
xor U33275 (N_33275,N_33176,N_33058);
or U33276 (N_33276,N_33151,N_33059);
nor U33277 (N_33277,N_33200,N_33143);
nand U33278 (N_33278,N_33134,N_33203);
nand U33279 (N_33279,N_33195,N_33065);
nor U33280 (N_33280,N_33048,N_33042);
xor U33281 (N_33281,N_33206,N_33073);
or U33282 (N_33282,N_33019,N_33004);
nand U33283 (N_33283,N_33202,N_33215);
xor U33284 (N_33284,N_33117,N_33078);
xor U33285 (N_33285,N_33179,N_33071);
and U33286 (N_33286,N_33124,N_33094);
and U33287 (N_33287,N_33141,N_33079);
nand U33288 (N_33288,N_33210,N_33187);
nor U33289 (N_33289,N_33098,N_33076);
nand U33290 (N_33290,N_33115,N_33154);
xor U33291 (N_33291,N_33204,N_33113);
xor U33292 (N_33292,N_33052,N_33020);
xnor U33293 (N_33293,N_33218,N_33224);
or U33294 (N_33294,N_33017,N_33233);
and U33295 (N_33295,N_33234,N_33074);
nor U33296 (N_33296,N_33043,N_33089);
nand U33297 (N_33297,N_33022,N_33023);
nor U33298 (N_33298,N_33190,N_33070);
nor U33299 (N_33299,N_33180,N_33080);
and U33300 (N_33300,N_33014,N_33140);
xor U33301 (N_33301,N_33238,N_33136);
nor U33302 (N_33302,N_33082,N_33231);
xnor U33303 (N_33303,N_33108,N_33050);
and U33304 (N_33304,N_33035,N_33162);
and U33305 (N_33305,N_33101,N_33057);
nor U33306 (N_33306,N_33145,N_33054);
or U33307 (N_33307,N_33123,N_33120);
xor U33308 (N_33308,N_33194,N_33211);
nand U33309 (N_33309,N_33041,N_33232);
xnor U33310 (N_33310,N_33128,N_33009);
nor U33311 (N_33311,N_33107,N_33243);
and U33312 (N_33312,N_33064,N_33011);
or U33313 (N_33313,N_33013,N_33099);
or U33314 (N_33314,N_33125,N_33165);
nand U33315 (N_33315,N_33142,N_33191);
xor U33316 (N_33316,N_33226,N_33005);
or U33317 (N_33317,N_33209,N_33106);
or U33318 (N_33318,N_33235,N_33055);
or U33319 (N_33319,N_33039,N_33249);
xnor U33320 (N_33320,N_33060,N_33021);
or U33321 (N_33321,N_33062,N_33129);
nor U33322 (N_33322,N_33150,N_33168);
xor U33323 (N_33323,N_33192,N_33018);
nand U33324 (N_33324,N_33247,N_33083);
nor U33325 (N_33325,N_33199,N_33103);
and U33326 (N_33326,N_33146,N_33010);
and U33327 (N_33327,N_33028,N_33026);
or U33328 (N_33328,N_33032,N_33087);
nand U33329 (N_33329,N_33075,N_33015);
or U33330 (N_33330,N_33027,N_33147);
or U33331 (N_33331,N_33207,N_33063);
nand U33332 (N_33332,N_33222,N_33100);
and U33333 (N_33333,N_33178,N_33111);
nand U33334 (N_33334,N_33096,N_33205);
nand U33335 (N_33335,N_33164,N_33102);
and U33336 (N_33336,N_33008,N_33229);
nor U33337 (N_33337,N_33174,N_33137);
xnor U33338 (N_33338,N_33220,N_33169);
nand U33339 (N_33339,N_33093,N_33046);
xor U33340 (N_33340,N_33072,N_33236);
nand U33341 (N_33341,N_33189,N_33126);
nor U33342 (N_33342,N_33171,N_33242);
and U33343 (N_33343,N_33030,N_33208);
nor U33344 (N_33344,N_33038,N_33034);
xor U33345 (N_33345,N_33016,N_33212);
and U33346 (N_33346,N_33149,N_33025);
xnor U33347 (N_33347,N_33047,N_33139);
nand U33348 (N_33348,N_33214,N_33053);
or U33349 (N_33349,N_33185,N_33109);
nor U33350 (N_33350,N_33219,N_33188);
or U33351 (N_33351,N_33086,N_33091);
and U33352 (N_33352,N_33245,N_33197);
xor U33353 (N_33353,N_33068,N_33135);
nor U33354 (N_33354,N_33003,N_33092);
and U33355 (N_33355,N_33237,N_33213);
nor U33356 (N_33356,N_33177,N_33127);
and U33357 (N_33357,N_33173,N_33056);
nor U33358 (N_33358,N_33170,N_33175);
and U33359 (N_33359,N_33217,N_33152);
nor U33360 (N_33360,N_33006,N_33067);
or U33361 (N_33361,N_33221,N_33085);
nand U33362 (N_33362,N_33037,N_33133);
xnor U33363 (N_33363,N_33183,N_33049);
nand U33364 (N_33364,N_33001,N_33040);
or U33365 (N_33365,N_33138,N_33066);
xor U33366 (N_33366,N_33158,N_33166);
and U33367 (N_33367,N_33161,N_33114);
xnor U33368 (N_33368,N_33144,N_33230);
nor U33369 (N_33369,N_33061,N_33000);
nand U33370 (N_33370,N_33155,N_33116);
and U33371 (N_33371,N_33097,N_33033);
or U33372 (N_33372,N_33119,N_33121);
and U33373 (N_33373,N_33081,N_33148);
and U33374 (N_33374,N_33077,N_33051);
nand U33375 (N_33375,N_33199,N_33106);
or U33376 (N_33376,N_33062,N_33046);
and U33377 (N_33377,N_33128,N_33075);
and U33378 (N_33378,N_33182,N_33150);
nor U33379 (N_33379,N_33009,N_33145);
nand U33380 (N_33380,N_33095,N_33101);
nand U33381 (N_33381,N_33231,N_33137);
and U33382 (N_33382,N_33138,N_33201);
nand U33383 (N_33383,N_33052,N_33131);
nor U33384 (N_33384,N_33191,N_33044);
nor U33385 (N_33385,N_33237,N_33035);
xnor U33386 (N_33386,N_33127,N_33032);
nor U33387 (N_33387,N_33065,N_33062);
and U33388 (N_33388,N_33085,N_33242);
or U33389 (N_33389,N_33246,N_33223);
xnor U33390 (N_33390,N_33135,N_33204);
nor U33391 (N_33391,N_33207,N_33106);
nand U33392 (N_33392,N_33234,N_33136);
xnor U33393 (N_33393,N_33128,N_33148);
xor U33394 (N_33394,N_33043,N_33157);
nor U33395 (N_33395,N_33016,N_33040);
and U33396 (N_33396,N_33170,N_33057);
and U33397 (N_33397,N_33036,N_33157);
nand U33398 (N_33398,N_33067,N_33247);
and U33399 (N_33399,N_33088,N_33028);
xnor U33400 (N_33400,N_33221,N_33074);
and U33401 (N_33401,N_33119,N_33023);
and U33402 (N_33402,N_33188,N_33127);
nand U33403 (N_33403,N_33206,N_33099);
or U33404 (N_33404,N_33174,N_33176);
or U33405 (N_33405,N_33060,N_33019);
xnor U33406 (N_33406,N_33044,N_33042);
and U33407 (N_33407,N_33204,N_33053);
or U33408 (N_33408,N_33097,N_33165);
and U33409 (N_33409,N_33124,N_33131);
and U33410 (N_33410,N_33067,N_33156);
nor U33411 (N_33411,N_33143,N_33083);
or U33412 (N_33412,N_33043,N_33185);
xor U33413 (N_33413,N_33067,N_33229);
and U33414 (N_33414,N_33023,N_33170);
or U33415 (N_33415,N_33024,N_33140);
or U33416 (N_33416,N_33115,N_33112);
and U33417 (N_33417,N_33217,N_33179);
nand U33418 (N_33418,N_33128,N_33034);
nand U33419 (N_33419,N_33006,N_33200);
nand U33420 (N_33420,N_33070,N_33108);
nor U33421 (N_33421,N_33023,N_33008);
or U33422 (N_33422,N_33023,N_33211);
nor U33423 (N_33423,N_33224,N_33014);
and U33424 (N_33424,N_33131,N_33061);
and U33425 (N_33425,N_33126,N_33029);
and U33426 (N_33426,N_33068,N_33167);
and U33427 (N_33427,N_33180,N_33185);
or U33428 (N_33428,N_33141,N_33145);
and U33429 (N_33429,N_33223,N_33093);
and U33430 (N_33430,N_33119,N_33022);
xor U33431 (N_33431,N_33143,N_33152);
and U33432 (N_33432,N_33192,N_33109);
or U33433 (N_33433,N_33014,N_33078);
and U33434 (N_33434,N_33068,N_33152);
or U33435 (N_33435,N_33030,N_33201);
nor U33436 (N_33436,N_33151,N_33170);
nand U33437 (N_33437,N_33064,N_33167);
nor U33438 (N_33438,N_33077,N_33122);
xnor U33439 (N_33439,N_33098,N_33052);
nand U33440 (N_33440,N_33214,N_33179);
nor U33441 (N_33441,N_33163,N_33130);
xor U33442 (N_33442,N_33120,N_33035);
nand U33443 (N_33443,N_33040,N_33075);
nor U33444 (N_33444,N_33018,N_33213);
and U33445 (N_33445,N_33130,N_33216);
xnor U33446 (N_33446,N_33132,N_33216);
xor U33447 (N_33447,N_33005,N_33222);
nor U33448 (N_33448,N_33108,N_33217);
nand U33449 (N_33449,N_33085,N_33039);
nor U33450 (N_33450,N_33123,N_33137);
nor U33451 (N_33451,N_33030,N_33016);
and U33452 (N_33452,N_33225,N_33052);
nand U33453 (N_33453,N_33226,N_33147);
and U33454 (N_33454,N_33107,N_33174);
nand U33455 (N_33455,N_33080,N_33160);
xor U33456 (N_33456,N_33222,N_33239);
nand U33457 (N_33457,N_33089,N_33030);
or U33458 (N_33458,N_33021,N_33153);
nand U33459 (N_33459,N_33065,N_33045);
nor U33460 (N_33460,N_33214,N_33177);
xor U33461 (N_33461,N_33091,N_33012);
xnor U33462 (N_33462,N_33151,N_33056);
nor U33463 (N_33463,N_33179,N_33105);
and U33464 (N_33464,N_33069,N_33044);
and U33465 (N_33465,N_33087,N_33019);
nand U33466 (N_33466,N_33016,N_33008);
and U33467 (N_33467,N_33163,N_33209);
or U33468 (N_33468,N_33111,N_33124);
or U33469 (N_33469,N_33053,N_33093);
nor U33470 (N_33470,N_33151,N_33120);
xor U33471 (N_33471,N_33186,N_33006);
xor U33472 (N_33472,N_33163,N_33210);
xor U33473 (N_33473,N_33041,N_33144);
xor U33474 (N_33474,N_33151,N_33179);
or U33475 (N_33475,N_33174,N_33119);
nand U33476 (N_33476,N_33147,N_33227);
or U33477 (N_33477,N_33019,N_33148);
nand U33478 (N_33478,N_33056,N_33236);
nor U33479 (N_33479,N_33177,N_33161);
and U33480 (N_33480,N_33171,N_33205);
and U33481 (N_33481,N_33119,N_33008);
and U33482 (N_33482,N_33220,N_33177);
or U33483 (N_33483,N_33219,N_33172);
nand U33484 (N_33484,N_33154,N_33156);
and U33485 (N_33485,N_33130,N_33066);
or U33486 (N_33486,N_33131,N_33200);
or U33487 (N_33487,N_33047,N_33224);
nand U33488 (N_33488,N_33240,N_33215);
nor U33489 (N_33489,N_33225,N_33145);
nor U33490 (N_33490,N_33049,N_33069);
or U33491 (N_33491,N_33103,N_33044);
or U33492 (N_33492,N_33156,N_33147);
nand U33493 (N_33493,N_33057,N_33185);
xnor U33494 (N_33494,N_33214,N_33118);
nand U33495 (N_33495,N_33182,N_33185);
xnor U33496 (N_33496,N_33061,N_33006);
nor U33497 (N_33497,N_33173,N_33183);
or U33498 (N_33498,N_33023,N_33130);
or U33499 (N_33499,N_33227,N_33156);
and U33500 (N_33500,N_33398,N_33486);
nor U33501 (N_33501,N_33386,N_33351);
and U33502 (N_33502,N_33495,N_33280);
and U33503 (N_33503,N_33261,N_33355);
nand U33504 (N_33504,N_33291,N_33372);
or U33505 (N_33505,N_33388,N_33327);
nand U33506 (N_33506,N_33407,N_33316);
and U33507 (N_33507,N_33473,N_33286);
or U33508 (N_33508,N_33290,N_33496);
nand U33509 (N_33509,N_33406,N_33455);
nor U33510 (N_33510,N_33384,N_33418);
or U33511 (N_33511,N_33449,N_33461);
nand U33512 (N_33512,N_33471,N_33399);
nor U33513 (N_33513,N_33416,N_33266);
nor U33514 (N_33514,N_33250,N_33448);
nor U33515 (N_33515,N_33382,N_33335);
or U33516 (N_33516,N_33295,N_33324);
nand U33517 (N_33517,N_33320,N_33370);
or U33518 (N_33518,N_33282,N_33492);
or U33519 (N_33519,N_33307,N_33332);
xnor U33520 (N_33520,N_33367,N_33312);
nor U33521 (N_33521,N_33342,N_33442);
and U33522 (N_33522,N_33293,N_33334);
nand U33523 (N_33523,N_33402,N_33333);
and U33524 (N_33524,N_33365,N_33460);
xnor U33525 (N_33525,N_33287,N_33321);
nor U33526 (N_33526,N_33452,N_33408);
and U33527 (N_33527,N_33410,N_33468);
xor U33528 (N_33528,N_33356,N_33259);
xor U33529 (N_33529,N_33318,N_33270);
nand U33530 (N_33530,N_33257,N_33437);
nand U33531 (N_33531,N_33359,N_33499);
nand U33532 (N_33532,N_33337,N_33456);
nand U33533 (N_33533,N_33268,N_33255);
nor U33534 (N_33534,N_33276,N_33360);
or U33535 (N_33535,N_33443,N_33381);
nor U33536 (N_33536,N_33436,N_33278);
xnor U33537 (N_33537,N_33353,N_33273);
nand U33538 (N_33538,N_33385,N_33378);
xnor U33539 (N_33539,N_33485,N_33390);
or U33540 (N_33540,N_33413,N_33432);
nand U33541 (N_33541,N_33440,N_33404);
nor U33542 (N_33542,N_33349,N_33377);
nor U33543 (N_33543,N_33325,N_33271);
xnor U33544 (N_33544,N_33348,N_33412);
or U33545 (N_33545,N_33454,N_33279);
or U33546 (N_33546,N_33379,N_33256);
and U33547 (N_33547,N_33415,N_33306);
xnor U33548 (N_33548,N_33441,N_33314);
and U33549 (N_33549,N_33414,N_33426);
and U33550 (N_33550,N_33393,N_33474);
nor U33551 (N_33551,N_33338,N_33345);
and U33552 (N_33552,N_33470,N_33429);
nor U33553 (N_33553,N_33310,N_33478);
nand U33554 (N_33554,N_33395,N_33258);
nand U33555 (N_33555,N_33430,N_33444);
nor U33556 (N_33556,N_33357,N_33420);
xor U33557 (N_33557,N_33482,N_33313);
and U33558 (N_33558,N_33494,N_33262);
or U33559 (N_33559,N_33435,N_33422);
or U33560 (N_33560,N_33469,N_33284);
nand U33561 (N_33561,N_33301,N_33303);
or U33562 (N_33562,N_33376,N_33308);
xor U33563 (N_33563,N_33375,N_33425);
xor U33564 (N_33564,N_33343,N_33267);
nand U33565 (N_33565,N_33341,N_33297);
nor U33566 (N_33566,N_33464,N_33401);
xor U33567 (N_33567,N_33383,N_33362);
or U33568 (N_33568,N_33354,N_33392);
or U33569 (N_33569,N_33487,N_33299);
or U33570 (N_33570,N_33264,N_33403);
or U33571 (N_33571,N_33329,N_33467);
xor U33572 (N_33572,N_33491,N_33305);
xor U33573 (N_33573,N_33380,N_33366);
nand U33574 (N_33574,N_33447,N_33364);
and U33575 (N_33575,N_33319,N_33445);
xor U33576 (N_33576,N_33277,N_33389);
xor U33577 (N_33577,N_33302,N_33328);
and U33578 (N_33578,N_33330,N_33252);
and U33579 (N_33579,N_33311,N_33427);
xor U33580 (N_33580,N_33344,N_33433);
xnor U33581 (N_33581,N_33394,N_33405);
and U33582 (N_33582,N_33417,N_33331);
and U33583 (N_33583,N_33304,N_33446);
and U33584 (N_33584,N_33275,N_33409);
nor U33585 (N_33585,N_33490,N_33371);
nor U33586 (N_33586,N_33397,N_33350);
xnor U33587 (N_33587,N_33493,N_33373);
nand U33588 (N_33588,N_33438,N_33477);
or U33589 (N_33589,N_33481,N_33260);
xnor U33590 (N_33590,N_33281,N_33358);
nand U33591 (N_33591,N_33439,N_33497);
nand U33592 (N_33592,N_33484,N_33480);
or U33593 (N_33593,N_33346,N_33488);
or U33594 (N_33594,N_33483,N_33434);
nor U33595 (N_33595,N_33254,N_33352);
xor U33596 (N_33596,N_33466,N_33457);
or U33597 (N_33597,N_33451,N_33315);
nor U33598 (N_33598,N_33400,N_33296);
or U33599 (N_33599,N_33453,N_33272);
and U33600 (N_33600,N_33472,N_33475);
nor U33601 (N_33601,N_33323,N_33462);
and U33602 (N_33602,N_33263,N_33489);
xnor U33603 (N_33603,N_33391,N_33411);
nand U33604 (N_33604,N_33431,N_33465);
or U33605 (N_33605,N_33428,N_33300);
nor U33606 (N_33606,N_33476,N_33265);
nor U33607 (N_33607,N_33336,N_33396);
and U33608 (N_33608,N_33274,N_33361);
and U33609 (N_33609,N_33283,N_33326);
and U33610 (N_33610,N_33309,N_33387);
or U33611 (N_33611,N_33423,N_33424);
xnor U33612 (N_33612,N_33340,N_33288);
xor U33613 (N_33613,N_33298,N_33369);
nand U33614 (N_33614,N_33294,N_33269);
and U33615 (N_33615,N_33479,N_33253);
or U33616 (N_33616,N_33450,N_33322);
xor U33617 (N_33617,N_33419,N_33421);
or U33618 (N_33618,N_33292,N_33347);
nand U33619 (N_33619,N_33251,N_33317);
nor U33620 (N_33620,N_33458,N_33285);
and U33621 (N_33621,N_33289,N_33459);
nor U33622 (N_33622,N_33463,N_33368);
and U33623 (N_33623,N_33339,N_33363);
and U33624 (N_33624,N_33498,N_33374);
nor U33625 (N_33625,N_33465,N_33414);
nand U33626 (N_33626,N_33327,N_33481);
nor U33627 (N_33627,N_33321,N_33265);
nand U33628 (N_33628,N_33341,N_33370);
nor U33629 (N_33629,N_33422,N_33252);
nand U33630 (N_33630,N_33374,N_33289);
xnor U33631 (N_33631,N_33279,N_33283);
nand U33632 (N_33632,N_33435,N_33478);
xor U33633 (N_33633,N_33253,N_33283);
and U33634 (N_33634,N_33494,N_33453);
nand U33635 (N_33635,N_33283,N_33344);
nand U33636 (N_33636,N_33449,N_33457);
xnor U33637 (N_33637,N_33434,N_33383);
nand U33638 (N_33638,N_33442,N_33370);
nor U33639 (N_33639,N_33467,N_33452);
xor U33640 (N_33640,N_33441,N_33494);
xnor U33641 (N_33641,N_33418,N_33424);
xor U33642 (N_33642,N_33381,N_33384);
or U33643 (N_33643,N_33429,N_33371);
nand U33644 (N_33644,N_33381,N_33267);
and U33645 (N_33645,N_33480,N_33314);
nand U33646 (N_33646,N_33499,N_33332);
or U33647 (N_33647,N_33286,N_33409);
and U33648 (N_33648,N_33423,N_33455);
xor U33649 (N_33649,N_33273,N_33493);
and U33650 (N_33650,N_33353,N_33346);
nand U33651 (N_33651,N_33295,N_33473);
nand U33652 (N_33652,N_33395,N_33498);
or U33653 (N_33653,N_33410,N_33386);
or U33654 (N_33654,N_33472,N_33453);
or U33655 (N_33655,N_33268,N_33330);
xnor U33656 (N_33656,N_33318,N_33391);
or U33657 (N_33657,N_33346,N_33416);
nor U33658 (N_33658,N_33433,N_33350);
or U33659 (N_33659,N_33323,N_33319);
nand U33660 (N_33660,N_33263,N_33461);
or U33661 (N_33661,N_33480,N_33391);
or U33662 (N_33662,N_33481,N_33468);
or U33663 (N_33663,N_33462,N_33381);
nand U33664 (N_33664,N_33311,N_33382);
nor U33665 (N_33665,N_33464,N_33379);
xor U33666 (N_33666,N_33330,N_33454);
or U33667 (N_33667,N_33414,N_33314);
xor U33668 (N_33668,N_33398,N_33412);
xor U33669 (N_33669,N_33417,N_33266);
nand U33670 (N_33670,N_33382,N_33273);
xor U33671 (N_33671,N_33360,N_33444);
nand U33672 (N_33672,N_33273,N_33342);
and U33673 (N_33673,N_33447,N_33256);
or U33674 (N_33674,N_33393,N_33438);
nor U33675 (N_33675,N_33259,N_33293);
nor U33676 (N_33676,N_33324,N_33417);
and U33677 (N_33677,N_33250,N_33457);
or U33678 (N_33678,N_33339,N_33483);
xnor U33679 (N_33679,N_33483,N_33472);
nor U33680 (N_33680,N_33442,N_33325);
or U33681 (N_33681,N_33403,N_33407);
xor U33682 (N_33682,N_33489,N_33451);
nand U33683 (N_33683,N_33439,N_33436);
or U33684 (N_33684,N_33303,N_33340);
nor U33685 (N_33685,N_33313,N_33373);
and U33686 (N_33686,N_33487,N_33279);
and U33687 (N_33687,N_33347,N_33407);
and U33688 (N_33688,N_33491,N_33475);
nor U33689 (N_33689,N_33273,N_33475);
or U33690 (N_33690,N_33414,N_33378);
or U33691 (N_33691,N_33421,N_33307);
nand U33692 (N_33692,N_33454,N_33443);
and U33693 (N_33693,N_33329,N_33356);
nor U33694 (N_33694,N_33437,N_33444);
nand U33695 (N_33695,N_33461,N_33439);
and U33696 (N_33696,N_33289,N_33293);
nor U33697 (N_33697,N_33491,N_33296);
xor U33698 (N_33698,N_33340,N_33314);
nor U33699 (N_33699,N_33431,N_33299);
or U33700 (N_33700,N_33347,N_33360);
and U33701 (N_33701,N_33300,N_33383);
xor U33702 (N_33702,N_33326,N_33456);
xnor U33703 (N_33703,N_33315,N_33314);
and U33704 (N_33704,N_33278,N_33429);
or U33705 (N_33705,N_33397,N_33365);
or U33706 (N_33706,N_33411,N_33401);
nand U33707 (N_33707,N_33484,N_33451);
or U33708 (N_33708,N_33310,N_33385);
or U33709 (N_33709,N_33425,N_33457);
nor U33710 (N_33710,N_33327,N_33395);
or U33711 (N_33711,N_33291,N_33286);
and U33712 (N_33712,N_33279,N_33438);
nand U33713 (N_33713,N_33491,N_33251);
nand U33714 (N_33714,N_33279,N_33259);
and U33715 (N_33715,N_33432,N_33275);
nor U33716 (N_33716,N_33410,N_33375);
nor U33717 (N_33717,N_33476,N_33414);
or U33718 (N_33718,N_33404,N_33461);
nor U33719 (N_33719,N_33306,N_33298);
or U33720 (N_33720,N_33481,N_33275);
nor U33721 (N_33721,N_33272,N_33392);
nor U33722 (N_33722,N_33379,N_33408);
xor U33723 (N_33723,N_33457,N_33372);
nand U33724 (N_33724,N_33459,N_33299);
or U33725 (N_33725,N_33267,N_33284);
or U33726 (N_33726,N_33365,N_33329);
nand U33727 (N_33727,N_33463,N_33370);
xor U33728 (N_33728,N_33491,N_33383);
xnor U33729 (N_33729,N_33476,N_33397);
nor U33730 (N_33730,N_33433,N_33365);
xnor U33731 (N_33731,N_33326,N_33483);
nand U33732 (N_33732,N_33476,N_33254);
nor U33733 (N_33733,N_33482,N_33376);
or U33734 (N_33734,N_33422,N_33285);
nand U33735 (N_33735,N_33404,N_33294);
or U33736 (N_33736,N_33281,N_33426);
nor U33737 (N_33737,N_33314,N_33271);
nand U33738 (N_33738,N_33357,N_33483);
nor U33739 (N_33739,N_33287,N_33254);
or U33740 (N_33740,N_33399,N_33303);
nand U33741 (N_33741,N_33294,N_33356);
xnor U33742 (N_33742,N_33257,N_33391);
nor U33743 (N_33743,N_33483,N_33389);
or U33744 (N_33744,N_33412,N_33434);
xnor U33745 (N_33745,N_33383,N_33468);
nand U33746 (N_33746,N_33493,N_33277);
or U33747 (N_33747,N_33297,N_33366);
nor U33748 (N_33748,N_33336,N_33438);
nor U33749 (N_33749,N_33488,N_33414);
or U33750 (N_33750,N_33613,N_33640);
or U33751 (N_33751,N_33503,N_33642);
and U33752 (N_33752,N_33687,N_33649);
or U33753 (N_33753,N_33666,N_33522);
nand U33754 (N_33754,N_33736,N_33507);
or U33755 (N_33755,N_33623,N_33715);
xnor U33756 (N_33756,N_33703,N_33568);
xnor U33757 (N_33757,N_33545,N_33609);
or U33758 (N_33758,N_33717,N_33583);
nand U33759 (N_33759,N_33725,N_33721);
and U33760 (N_33760,N_33540,N_33551);
or U33761 (N_33761,N_33657,N_33636);
xnor U33762 (N_33762,N_33719,N_33589);
xnor U33763 (N_33763,N_33709,N_33704);
xor U33764 (N_33764,N_33580,N_33518);
xnor U33765 (N_33765,N_33677,N_33711);
and U33766 (N_33766,N_33607,N_33734);
or U33767 (N_33767,N_33556,N_33651);
or U33768 (N_33768,N_33534,N_33602);
and U33769 (N_33769,N_33587,N_33659);
or U33770 (N_33770,N_33630,N_33614);
nor U33771 (N_33771,N_33696,N_33653);
or U33772 (N_33772,N_33591,N_33529);
nand U33773 (N_33773,N_33596,N_33532);
and U33774 (N_33774,N_33673,N_33627);
nand U33775 (N_33775,N_33552,N_33645);
and U33776 (N_33776,N_33575,N_33533);
nor U33777 (N_33777,N_33699,N_33537);
or U33778 (N_33778,N_33694,N_33650);
or U33779 (N_33779,N_33510,N_33678);
or U33780 (N_33780,N_33606,N_33512);
nand U33781 (N_33781,N_33595,N_33599);
xnor U33782 (N_33782,N_33557,N_33565);
or U33783 (N_33783,N_33726,N_33601);
or U33784 (N_33784,N_33558,N_33712);
and U33785 (N_33785,N_33670,N_33621);
xnor U33786 (N_33786,N_33585,N_33646);
or U33787 (N_33787,N_33631,N_33598);
nor U33788 (N_33788,N_33597,N_33735);
nand U33789 (N_33789,N_33626,N_33740);
and U33790 (N_33790,N_33539,N_33722);
xnor U33791 (N_33791,N_33577,N_33662);
xnor U33792 (N_33792,N_33641,N_33643);
nand U33793 (N_33793,N_33502,N_33586);
or U33794 (N_33794,N_33652,N_33701);
xor U33795 (N_33795,N_33560,N_33569);
xnor U33796 (N_33796,N_33618,N_33679);
nor U33797 (N_33797,N_33525,N_33689);
or U33798 (N_33798,N_33566,N_33654);
or U33799 (N_33799,N_33676,N_33690);
nor U33800 (N_33800,N_33706,N_33663);
or U33801 (N_33801,N_33655,N_33672);
xnor U33802 (N_33802,N_33521,N_33548);
and U33803 (N_33803,N_33691,N_33592);
and U33804 (N_33804,N_33695,N_33553);
and U33805 (N_33805,N_33682,N_33504);
or U33806 (N_33806,N_33674,N_33500);
nor U33807 (N_33807,N_33612,N_33702);
or U33808 (N_33808,N_33634,N_33671);
nand U33809 (N_33809,N_33505,N_33541);
or U33810 (N_33810,N_33698,N_33629);
xnor U33811 (N_33811,N_33668,N_33747);
nor U33812 (N_33812,N_33675,N_33658);
and U33813 (N_33813,N_33531,N_33543);
or U33814 (N_33814,N_33608,N_33620);
or U33815 (N_33815,N_33574,N_33624);
nor U33816 (N_33816,N_33547,N_33632);
or U33817 (N_33817,N_33637,N_33564);
xnor U33818 (N_33818,N_33737,N_33661);
or U33819 (N_33819,N_33563,N_33544);
nor U33820 (N_33820,N_33588,N_33524);
nand U33821 (N_33821,N_33604,N_33710);
or U33822 (N_33822,N_33688,N_33559);
nand U33823 (N_33823,N_33681,N_33680);
nand U33824 (N_33824,N_33693,N_33526);
nor U33825 (N_33825,N_33733,N_33656);
nand U33826 (N_33826,N_33714,N_33605);
nor U33827 (N_33827,N_33619,N_33600);
xnor U33828 (N_33828,N_33576,N_33667);
or U33829 (N_33829,N_33514,N_33684);
xor U33830 (N_33830,N_33508,N_33622);
xor U33831 (N_33831,N_33542,N_33509);
and U33832 (N_33832,N_33616,N_33648);
xnor U33833 (N_33833,N_33546,N_33579);
or U33834 (N_33834,N_33728,N_33665);
or U33835 (N_33835,N_33549,N_33732);
or U33836 (N_33836,N_33692,N_33581);
nor U33837 (N_33837,N_33615,N_33535);
nor U33838 (N_33838,N_33685,N_33724);
xnor U33839 (N_33839,N_33749,N_33707);
nor U33840 (N_33840,N_33567,N_33515);
or U33841 (N_33841,N_33748,N_33571);
or U33842 (N_33842,N_33570,N_33530);
or U33843 (N_33843,N_33603,N_33572);
nor U33844 (N_33844,N_33669,N_33538);
nor U33845 (N_33845,N_33617,N_33644);
or U33846 (N_33846,N_33729,N_33639);
or U33847 (N_33847,N_33511,N_33705);
and U33848 (N_33848,N_33516,N_33611);
nor U33849 (N_33849,N_33519,N_33700);
nand U33850 (N_33850,N_33550,N_33561);
and U33851 (N_33851,N_33501,N_33686);
and U33852 (N_33852,N_33730,N_33746);
or U33853 (N_33853,N_33513,N_33520);
xnor U33854 (N_33854,N_33744,N_33720);
nand U33855 (N_33855,N_33697,N_33554);
and U33856 (N_33856,N_33523,N_33517);
and U33857 (N_33857,N_33638,N_33723);
xnor U33858 (N_33858,N_33708,N_33590);
xnor U33859 (N_33859,N_33664,N_33506);
nor U33860 (N_33860,N_33628,N_33584);
nor U33861 (N_33861,N_33555,N_33633);
nand U33862 (N_33862,N_33716,N_33742);
and U33863 (N_33863,N_33562,N_33660);
xnor U33864 (N_33864,N_33738,N_33713);
or U33865 (N_33865,N_33739,N_33718);
and U33866 (N_33866,N_33745,N_33582);
or U33867 (N_33867,N_33625,N_33741);
nand U33868 (N_33868,N_33683,N_33743);
xor U33869 (N_33869,N_33527,N_33635);
nand U33870 (N_33870,N_33647,N_33528);
nor U33871 (N_33871,N_33536,N_33731);
nand U33872 (N_33872,N_33593,N_33594);
nor U33873 (N_33873,N_33727,N_33573);
nand U33874 (N_33874,N_33610,N_33578);
and U33875 (N_33875,N_33667,N_33731);
xor U33876 (N_33876,N_33693,N_33551);
nor U33877 (N_33877,N_33711,N_33543);
nor U33878 (N_33878,N_33714,N_33704);
and U33879 (N_33879,N_33724,N_33707);
nor U33880 (N_33880,N_33619,N_33653);
nor U33881 (N_33881,N_33569,N_33686);
and U33882 (N_33882,N_33613,N_33556);
and U33883 (N_33883,N_33685,N_33717);
xnor U33884 (N_33884,N_33541,N_33653);
nor U33885 (N_33885,N_33639,N_33535);
or U33886 (N_33886,N_33635,N_33663);
xor U33887 (N_33887,N_33666,N_33573);
or U33888 (N_33888,N_33546,N_33628);
xor U33889 (N_33889,N_33722,N_33619);
nor U33890 (N_33890,N_33674,N_33570);
and U33891 (N_33891,N_33590,N_33739);
and U33892 (N_33892,N_33657,N_33594);
nor U33893 (N_33893,N_33719,N_33562);
and U33894 (N_33894,N_33693,N_33516);
xor U33895 (N_33895,N_33637,N_33710);
nor U33896 (N_33896,N_33716,N_33724);
and U33897 (N_33897,N_33547,N_33568);
or U33898 (N_33898,N_33582,N_33591);
xor U33899 (N_33899,N_33514,N_33587);
nor U33900 (N_33900,N_33645,N_33553);
nor U33901 (N_33901,N_33526,N_33633);
and U33902 (N_33902,N_33597,N_33695);
xnor U33903 (N_33903,N_33545,N_33706);
or U33904 (N_33904,N_33535,N_33516);
and U33905 (N_33905,N_33680,N_33655);
and U33906 (N_33906,N_33506,N_33589);
nor U33907 (N_33907,N_33683,N_33672);
nand U33908 (N_33908,N_33637,N_33659);
nand U33909 (N_33909,N_33571,N_33680);
xor U33910 (N_33910,N_33709,N_33713);
or U33911 (N_33911,N_33562,N_33716);
or U33912 (N_33912,N_33633,N_33583);
and U33913 (N_33913,N_33713,N_33575);
or U33914 (N_33914,N_33555,N_33648);
or U33915 (N_33915,N_33706,N_33737);
nand U33916 (N_33916,N_33527,N_33516);
and U33917 (N_33917,N_33571,N_33578);
xor U33918 (N_33918,N_33692,N_33672);
and U33919 (N_33919,N_33568,N_33718);
and U33920 (N_33920,N_33705,N_33724);
xnor U33921 (N_33921,N_33612,N_33685);
nand U33922 (N_33922,N_33682,N_33647);
and U33923 (N_33923,N_33593,N_33630);
or U33924 (N_33924,N_33599,N_33638);
and U33925 (N_33925,N_33536,N_33523);
or U33926 (N_33926,N_33665,N_33689);
or U33927 (N_33927,N_33521,N_33606);
xor U33928 (N_33928,N_33558,N_33568);
nand U33929 (N_33929,N_33639,N_33713);
nand U33930 (N_33930,N_33660,N_33697);
nor U33931 (N_33931,N_33623,N_33576);
xor U33932 (N_33932,N_33576,N_33591);
and U33933 (N_33933,N_33678,N_33522);
nand U33934 (N_33934,N_33719,N_33724);
or U33935 (N_33935,N_33570,N_33645);
nor U33936 (N_33936,N_33618,N_33627);
nor U33937 (N_33937,N_33595,N_33530);
nand U33938 (N_33938,N_33510,N_33616);
nor U33939 (N_33939,N_33576,N_33505);
nand U33940 (N_33940,N_33708,N_33525);
or U33941 (N_33941,N_33749,N_33569);
nor U33942 (N_33942,N_33677,N_33509);
and U33943 (N_33943,N_33706,N_33625);
nand U33944 (N_33944,N_33681,N_33662);
xor U33945 (N_33945,N_33528,N_33501);
nand U33946 (N_33946,N_33596,N_33559);
nor U33947 (N_33947,N_33623,N_33653);
nand U33948 (N_33948,N_33742,N_33659);
xnor U33949 (N_33949,N_33656,N_33547);
nand U33950 (N_33950,N_33502,N_33563);
nor U33951 (N_33951,N_33506,N_33706);
and U33952 (N_33952,N_33666,N_33702);
nand U33953 (N_33953,N_33663,N_33626);
or U33954 (N_33954,N_33660,N_33692);
nor U33955 (N_33955,N_33685,N_33737);
and U33956 (N_33956,N_33728,N_33541);
nand U33957 (N_33957,N_33571,N_33550);
nor U33958 (N_33958,N_33682,N_33609);
or U33959 (N_33959,N_33732,N_33589);
or U33960 (N_33960,N_33550,N_33568);
xor U33961 (N_33961,N_33569,N_33728);
nor U33962 (N_33962,N_33500,N_33649);
nand U33963 (N_33963,N_33593,N_33555);
and U33964 (N_33964,N_33671,N_33654);
and U33965 (N_33965,N_33552,N_33710);
nand U33966 (N_33966,N_33675,N_33681);
and U33967 (N_33967,N_33591,N_33717);
and U33968 (N_33968,N_33596,N_33692);
and U33969 (N_33969,N_33587,N_33581);
nand U33970 (N_33970,N_33590,N_33674);
or U33971 (N_33971,N_33587,N_33692);
xnor U33972 (N_33972,N_33665,N_33632);
nor U33973 (N_33973,N_33698,N_33643);
nor U33974 (N_33974,N_33575,N_33548);
nand U33975 (N_33975,N_33598,N_33615);
or U33976 (N_33976,N_33533,N_33530);
nor U33977 (N_33977,N_33616,N_33643);
or U33978 (N_33978,N_33585,N_33552);
xnor U33979 (N_33979,N_33599,N_33649);
nor U33980 (N_33980,N_33640,N_33641);
and U33981 (N_33981,N_33525,N_33550);
nand U33982 (N_33982,N_33668,N_33576);
and U33983 (N_33983,N_33526,N_33580);
and U33984 (N_33984,N_33575,N_33746);
and U33985 (N_33985,N_33689,N_33732);
or U33986 (N_33986,N_33712,N_33618);
or U33987 (N_33987,N_33694,N_33516);
xnor U33988 (N_33988,N_33538,N_33734);
nand U33989 (N_33989,N_33560,N_33538);
and U33990 (N_33990,N_33602,N_33696);
nand U33991 (N_33991,N_33600,N_33734);
and U33992 (N_33992,N_33718,N_33521);
and U33993 (N_33993,N_33695,N_33620);
nor U33994 (N_33994,N_33603,N_33641);
and U33995 (N_33995,N_33552,N_33600);
xnor U33996 (N_33996,N_33609,N_33622);
xnor U33997 (N_33997,N_33591,N_33533);
and U33998 (N_33998,N_33535,N_33594);
xor U33999 (N_33999,N_33736,N_33739);
nor U34000 (N_34000,N_33919,N_33865);
nor U34001 (N_34001,N_33913,N_33896);
xor U34002 (N_34002,N_33916,N_33862);
xnor U34003 (N_34003,N_33992,N_33923);
and U34004 (N_34004,N_33835,N_33817);
and U34005 (N_34005,N_33824,N_33974);
xnor U34006 (N_34006,N_33796,N_33864);
nor U34007 (N_34007,N_33965,N_33950);
and U34008 (N_34008,N_33931,N_33845);
nand U34009 (N_34009,N_33847,N_33907);
nor U34010 (N_34010,N_33764,N_33832);
or U34011 (N_34011,N_33932,N_33980);
or U34012 (N_34012,N_33902,N_33802);
or U34013 (N_34013,N_33883,N_33823);
nand U34014 (N_34014,N_33828,N_33952);
nor U34015 (N_34015,N_33971,N_33797);
nor U34016 (N_34016,N_33782,N_33921);
and U34017 (N_34017,N_33788,N_33898);
nor U34018 (N_34018,N_33861,N_33936);
xnor U34019 (N_34019,N_33754,N_33978);
or U34020 (N_34020,N_33994,N_33996);
nor U34021 (N_34021,N_33777,N_33818);
nor U34022 (N_34022,N_33860,N_33998);
nand U34023 (N_34023,N_33810,N_33918);
xnor U34024 (N_34024,N_33838,N_33939);
nor U34025 (N_34025,N_33816,N_33943);
nand U34026 (N_34026,N_33956,N_33868);
or U34027 (N_34027,N_33842,N_33758);
and U34028 (N_34028,N_33927,N_33922);
xor U34029 (N_34029,N_33881,N_33890);
xnor U34030 (N_34030,N_33787,N_33848);
or U34031 (N_34031,N_33946,N_33940);
nand U34032 (N_34032,N_33806,N_33933);
or U34033 (N_34033,N_33834,N_33803);
nor U34034 (N_34034,N_33863,N_33964);
xor U34035 (N_34035,N_33867,N_33825);
or U34036 (N_34036,N_33768,N_33779);
or U34037 (N_34037,N_33814,N_33856);
or U34038 (N_34038,N_33853,N_33947);
and U34039 (N_34039,N_33770,N_33973);
nand U34040 (N_34040,N_33905,N_33910);
nand U34041 (N_34041,N_33988,N_33897);
nand U34042 (N_34042,N_33794,N_33953);
nand U34043 (N_34043,N_33786,N_33789);
nand U34044 (N_34044,N_33977,N_33908);
and U34045 (N_34045,N_33986,N_33780);
nor U34046 (N_34046,N_33813,N_33804);
nand U34047 (N_34047,N_33761,N_33812);
or U34048 (N_34048,N_33801,N_33850);
nand U34049 (N_34049,N_33886,N_33773);
nand U34050 (N_34050,N_33982,N_33903);
xnor U34051 (N_34051,N_33869,N_33955);
nand U34052 (N_34052,N_33799,N_33901);
xnor U34053 (N_34053,N_33917,N_33769);
nand U34054 (N_34054,N_33959,N_33962);
nand U34055 (N_34055,N_33873,N_33885);
or U34056 (N_34056,N_33819,N_33876);
or U34057 (N_34057,N_33987,N_33808);
nor U34058 (N_34058,N_33822,N_33878);
and U34059 (N_34059,N_33963,N_33830);
nor U34060 (N_34060,N_33846,N_33843);
and U34061 (N_34061,N_33763,N_33870);
and U34062 (N_34062,N_33859,N_33957);
and U34063 (N_34063,N_33985,N_33841);
nor U34064 (N_34064,N_33800,N_33821);
xnor U34065 (N_34065,N_33968,N_33925);
nand U34066 (N_34066,N_33755,N_33831);
nand U34067 (N_34067,N_33972,N_33990);
nand U34068 (N_34068,N_33894,N_33944);
nand U34069 (N_34069,N_33766,N_33966);
nor U34070 (N_34070,N_33776,N_33900);
nor U34071 (N_34071,N_33760,N_33951);
or U34072 (N_34072,N_33983,N_33899);
and U34073 (N_34073,N_33945,N_33854);
and U34074 (N_34074,N_33781,N_33938);
nand U34075 (N_34075,N_33887,N_33941);
and U34076 (N_34076,N_33807,N_33997);
nand U34077 (N_34077,N_33879,N_33991);
nor U34078 (N_34078,N_33995,N_33874);
or U34079 (N_34079,N_33904,N_33970);
nand U34080 (N_34080,N_33771,N_33911);
xnor U34081 (N_34081,N_33820,N_33811);
nand U34082 (N_34082,N_33915,N_33750);
or U34083 (N_34083,N_33993,N_33891);
xnor U34084 (N_34084,N_33937,N_33778);
nand U34085 (N_34085,N_33912,N_33979);
xnor U34086 (N_34086,N_33767,N_33762);
and U34087 (N_34087,N_33774,N_33790);
nor U34088 (N_34088,N_33976,N_33772);
nor U34089 (N_34089,N_33928,N_33948);
nor U34090 (N_34090,N_33960,N_33893);
and U34091 (N_34091,N_33866,N_33858);
and U34092 (N_34092,N_33975,N_33969);
xnor U34093 (N_34093,N_33929,N_33884);
xor U34094 (N_34094,N_33989,N_33775);
nand U34095 (N_34095,N_33880,N_33815);
and U34096 (N_34096,N_33935,N_33827);
nand U34097 (N_34097,N_33914,N_33920);
nor U34098 (N_34098,N_33855,N_33954);
or U34099 (N_34099,N_33829,N_33967);
and U34100 (N_34100,N_33999,N_33909);
or U34101 (N_34101,N_33833,N_33759);
and U34102 (N_34102,N_33872,N_33751);
or U34103 (N_34103,N_33882,N_33753);
nor U34104 (N_34104,N_33958,N_33852);
nor U34105 (N_34105,N_33840,N_33857);
nor U34106 (N_34106,N_33984,N_33934);
and U34107 (N_34107,N_33906,N_33877);
nand U34108 (N_34108,N_33851,N_33875);
or U34109 (N_34109,N_33791,N_33809);
and U34110 (N_34110,N_33844,N_33805);
nand U34111 (N_34111,N_33924,N_33849);
and U34112 (N_34112,N_33756,N_33981);
xor U34113 (N_34113,N_33783,N_33793);
nand U34114 (N_34114,N_33949,N_33792);
xnor U34115 (N_34115,N_33871,N_33895);
nand U34116 (N_34116,N_33961,N_33930);
xnor U34117 (N_34117,N_33892,N_33888);
nand U34118 (N_34118,N_33837,N_33826);
xor U34119 (N_34119,N_33784,N_33836);
xor U34120 (N_34120,N_33785,N_33942);
and U34121 (N_34121,N_33798,N_33889);
nand U34122 (N_34122,N_33752,N_33795);
or U34123 (N_34123,N_33757,N_33926);
and U34124 (N_34124,N_33839,N_33765);
or U34125 (N_34125,N_33795,N_33841);
xor U34126 (N_34126,N_33812,N_33991);
nor U34127 (N_34127,N_33922,N_33850);
nor U34128 (N_34128,N_33998,N_33892);
and U34129 (N_34129,N_33949,N_33861);
or U34130 (N_34130,N_33793,N_33828);
nor U34131 (N_34131,N_33879,N_33881);
nor U34132 (N_34132,N_33910,N_33972);
xnor U34133 (N_34133,N_33902,N_33954);
and U34134 (N_34134,N_33902,N_33912);
nor U34135 (N_34135,N_33775,N_33876);
nand U34136 (N_34136,N_33906,N_33812);
and U34137 (N_34137,N_33769,N_33999);
nand U34138 (N_34138,N_33782,N_33826);
nand U34139 (N_34139,N_33922,N_33844);
nor U34140 (N_34140,N_33968,N_33911);
or U34141 (N_34141,N_33994,N_33995);
and U34142 (N_34142,N_33757,N_33922);
or U34143 (N_34143,N_33814,N_33825);
and U34144 (N_34144,N_33761,N_33973);
and U34145 (N_34145,N_33785,N_33974);
or U34146 (N_34146,N_33938,N_33817);
and U34147 (N_34147,N_33851,N_33860);
xnor U34148 (N_34148,N_33997,N_33963);
nor U34149 (N_34149,N_33778,N_33795);
nand U34150 (N_34150,N_33925,N_33980);
nor U34151 (N_34151,N_33895,N_33945);
xor U34152 (N_34152,N_33932,N_33952);
xor U34153 (N_34153,N_33972,N_33939);
xor U34154 (N_34154,N_33826,N_33821);
or U34155 (N_34155,N_33928,N_33862);
and U34156 (N_34156,N_33918,N_33814);
xor U34157 (N_34157,N_33866,N_33924);
and U34158 (N_34158,N_33937,N_33812);
nand U34159 (N_34159,N_33795,N_33921);
nand U34160 (N_34160,N_33875,N_33863);
xnor U34161 (N_34161,N_33858,N_33790);
or U34162 (N_34162,N_33774,N_33779);
nor U34163 (N_34163,N_33832,N_33923);
nand U34164 (N_34164,N_33838,N_33858);
nor U34165 (N_34165,N_33819,N_33945);
nor U34166 (N_34166,N_33877,N_33781);
or U34167 (N_34167,N_33938,N_33841);
nand U34168 (N_34168,N_33917,N_33767);
nand U34169 (N_34169,N_33990,N_33906);
nor U34170 (N_34170,N_33771,N_33921);
nor U34171 (N_34171,N_33917,N_33971);
nand U34172 (N_34172,N_33911,N_33765);
xnor U34173 (N_34173,N_33965,N_33993);
and U34174 (N_34174,N_33888,N_33785);
nor U34175 (N_34175,N_33779,N_33974);
and U34176 (N_34176,N_33792,N_33842);
or U34177 (N_34177,N_33904,N_33979);
nor U34178 (N_34178,N_33842,N_33955);
nand U34179 (N_34179,N_33955,N_33896);
and U34180 (N_34180,N_33966,N_33775);
or U34181 (N_34181,N_33765,N_33881);
or U34182 (N_34182,N_33882,N_33838);
nor U34183 (N_34183,N_33869,N_33805);
nor U34184 (N_34184,N_33788,N_33873);
nor U34185 (N_34185,N_33763,N_33904);
xor U34186 (N_34186,N_33912,N_33841);
nand U34187 (N_34187,N_33799,N_33928);
or U34188 (N_34188,N_33871,N_33894);
xnor U34189 (N_34189,N_33972,N_33779);
xnor U34190 (N_34190,N_33892,N_33813);
nor U34191 (N_34191,N_33856,N_33753);
nand U34192 (N_34192,N_33890,N_33844);
and U34193 (N_34193,N_33959,N_33778);
nor U34194 (N_34194,N_33957,N_33872);
and U34195 (N_34195,N_33781,N_33942);
or U34196 (N_34196,N_33860,N_33824);
nor U34197 (N_34197,N_33758,N_33963);
nand U34198 (N_34198,N_33964,N_33801);
xor U34199 (N_34199,N_33929,N_33824);
and U34200 (N_34200,N_33902,N_33899);
and U34201 (N_34201,N_33924,N_33828);
xnor U34202 (N_34202,N_33957,N_33911);
nand U34203 (N_34203,N_33781,N_33843);
or U34204 (N_34204,N_33771,N_33961);
xor U34205 (N_34205,N_33919,N_33778);
xnor U34206 (N_34206,N_33875,N_33850);
xor U34207 (N_34207,N_33876,N_33859);
nor U34208 (N_34208,N_33982,N_33964);
nand U34209 (N_34209,N_33972,N_33937);
nor U34210 (N_34210,N_33932,N_33968);
xor U34211 (N_34211,N_33774,N_33888);
or U34212 (N_34212,N_33779,N_33827);
xor U34213 (N_34213,N_33869,N_33811);
or U34214 (N_34214,N_33771,N_33832);
xnor U34215 (N_34215,N_33931,N_33994);
nand U34216 (N_34216,N_33805,N_33976);
nor U34217 (N_34217,N_33917,N_33885);
and U34218 (N_34218,N_33966,N_33839);
and U34219 (N_34219,N_33915,N_33988);
nor U34220 (N_34220,N_33828,N_33808);
nor U34221 (N_34221,N_33785,N_33875);
or U34222 (N_34222,N_33839,N_33819);
and U34223 (N_34223,N_33853,N_33860);
or U34224 (N_34224,N_33913,N_33895);
nor U34225 (N_34225,N_33827,N_33821);
or U34226 (N_34226,N_33862,N_33880);
nand U34227 (N_34227,N_33989,N_33860);
xor U34228 (N_34228,N_33905,N_33780);
or U34229 (N_34229,N_33959,N_33916);
nor U34230 (N_34230,N_33774,N_33791);
or U34231 (N_34231,N_33944,N_33969);
and U34232 (N_34232,N_33932,N_33914);
nand U34233 (N_34233,N_33900,N_33858);
nor U34234 (N_34234,N_33790,N_33761);
and U34235 (N_34235,N_33979,N_33864);
nor U34236 (N_34236,N_33775,N_33947);
xor U34237 (N_34237,N_33800,N_33778);
and U34238 (N_34238,N_33887,N_33918);
and U34239 (N_34239,N_33904,N_33797);
xnor U34240 (N_34240,N_33939,N_33915);
nor U34241 (N_34241,N_33983,N_33910);
nand U34242 (N_34242,N_33846,N_33989);
or U34243 (N_34243,N_33935,N_33957);
and U34244 (N_34244,N_33824,N_33918);
or U34245 (N_34245,N_33921,N_33767);
nor U34246 (N_34246,N_33934,N_33794);
xor U34247 (N_34247,N_33834,N_33773);
or U34248 (N_34248,N_33981,N_33874);
nor U34249 (N_34249,N_33797,N_33783);
and U34250 (N_34250,N_34008,N_34147);
and U34251 (N_34251,N_34100,N_34024);
nand U34252 (N_34252,N_34212,N_34188);
xnor U34253 (N_34253,N_34187,N_34145);
nor U34254 (N_34254,N_34151,N_34082);
or U34255 (N_34255,N_34184,N_34055);
xnor U34256 (N_34256,N_34016,N_34172);
nor U34257 (N_34257,N_34009,N_34171);
nor U34258 (N_34258,N_34164,N_34070);
nand U34259 (N_34259,N_34032,N_34037);
nand U34260 (N_34260,N_34051,N_34226);
and U34261 (N_34261,N_34074,N_34192);
and U34262 (N_34262,N_34246,N_34219);
and U34263 (N_34263,N_34213,N_34177);
xor U34264 (N_34264,N_34231,N_34058);
or U34265 (N_34265,N_34097,N_34129);
or U34266 (N_34266,N_34143,N_34191);
xnor U34267 (N_34267,N_34222,N_34110);
nor U34268 (N_34268,N_34133,N_34062);
nor U34269 (N_34269,N_34022,N_34241);
nand U34270 (N_34270,N_34175,N_34002);
and U34271 (N_34271,N_34190,N_34098);
xor U34272 (N_34272,N_34088,N_34208);
nor U34273 (N_34273,N_34076,N_34033);
nor U34274 (N_34274,N_34113,N_34056);
or U34275 (N_34275,N_34077,N_34013);
and U34276 (N_34276,N_34135,N_34047);
xnor U34277 (N_34277,N_34180,N_34085);
and U34278 (N_34278,N_34214,N_34039);
nand U34279 (N_34279,N_34007,N_34029);
nand U34280 (N_34280,N_34086,N_34115);
xnor U34281 (N_34281,N_34136,N_34216);
and U34282 (N_34282,N_34126,N_34099);
or U34283 (N_34283,N_34227,N_34026);
xnor U34284 (N_34284,N_34018,N_34153);
and U34285 (N_34285,N_34131,N_34069);
xnor U34286 (N_34286,N_34004,N_34163);
nor U34287 (N_34287,N_34064,N_34057);
and U34288 (N_34288,N_34108,N_34049);
and U34289 (N_34289,N_34244,N_34050);
xnor U34290 (N_34290,N_34193,N_34146);
or U34291 (N_34291,N_34228,N_34245);
nor U34292 (N_34292,N_34243,N_34234);
xnor U34293 (N_34293,N_34122,N_34158);
nor U34294 (N_34294,N_34091,N_34040);
xor U34295 (N_34295,N_34090,N_34152);
nor U34296 (N_34296,N_34137,N_34157);
nor U34297 (N_34297,N_34217,N_34201);
nor U34298 (N_34298,N_34112,N_34053);
xnor U34299 (N_34299,N_34169,N_34023);
xor U34300 (N_34300,N_34041,N_34239);
and U34301 (N_34301,N_34148,N_34198);
xnor U34302 (N_34302,N_34149,N_34215);
xor U34303 (N_34303,N_34031,N_34012);
nor U34304 (N_34304,N_34144,N_34087);
xnor U34305 (N_34305,N_34078,N_34107);
or U34306 (N_34306,N_34165,N_34142);
nor U34307 (N_34307,N_34189,N_34210);
nand U34308 (N_34308,N_34025,N_34066);
xnor U34309 (N_34309,N_34200,N_34006);
nor U34310 (N_34310,N_34072,N_34068);
nor U34311 (N_34311,N_34242,N_34178);
and U34312 (N_34312,N_34170,N_34119);
nor U34313 (N_34313,N_34020,N_34003);
nand U34314 (N_34314,N_34046,N_34038);
nand U34315 (N_34315,N_34204,N_34125);
nor U34316 (N_34316,N_34124,N_34060);
xnor U34317 (N_34317,N_34021,N_34205);
nand U34318 (N_34318,N_34159,N_34238);
and U34319 (N_34319,N_34156,N_34073);
and U34320 (N_34320,N_34127,N_34120);
or U34321 (N_34321,N_34042,N_34117);
xnor U34322 (N_34322,N_34236,N_34011);
nand U34323 (N_34323,N_34017,N_34092);
nor U34324 (N_34324,N_34209,N_34247);
and U34325 (N_34325,N_34045,N_34161);
nand U34326 (N_34326,N_34221,N_34054);
nand U34327 (N_34327,N_34207,N_34083);
and U34328 (N_34328,N_34063,N_34116);
nor U34329 (N_34329,N_34181,N_34123);
and U34330 (N_34330,N_34089,N_34102);
nor U34331 (N_34331,N_34220,N_34202);
and U34332 (N_34332,N_34197,N_34035);
or U34333 (N_34333,N_34121,N_34196);
nor U34334 (N_34334,N_34248,N_34139);
or U34335 (N_34335,N_34109,N_34150);
or U34336 (N_34336,N_34095,N_34075);
and U34337 (N_34337,N_34103,N_34176);
or U34338 (N_34338,N_34182,N_34138);
xnor U34339 (N_34339,N_34067,N_34154);
xnor U34340 (N_34340,N_34130,N_34030);
nand U34341 (N_34341,N_34093,N_34014);
and U34342 (N_34342,N_34132,N_34101);
nand U34343 (N_34343,N_34174,N_34104);
xor U34344 (N_34344,N_34114,N_34167);
nand U34345 (N_34345,N_34000,N_34223);
nor U34346 (N_34346,N_34128,N_34015);
nor U34347 (N_34347,N_34010,N_34036);
nor U34348 (N_34348,N_34160,N_34061);
nand U34349 (N_34349,N_34183,N_34218);
or U34350 (N_34350,N_34229,N_34168);
nand U34351 (N_34351,N_34225,N_34195);
xor U34352 (N_34352,N_34179,N_34203);
and U34353 (N_34353,N_34166,N_34237);
or U34354 (N_34354,N_34048,N_34211);
nand U34355 (N_34355,N_34059,N_34079);
and U34356 (N_34356,N_34094,N_34162);
and U34357 (N_34357,N_34235,N_34194);
and U34358 (N_34358,N_34173,N_34233);
nand U34359 (N_34359,N_34106,N_34186);
and U34360 (N_34360,N_34034,N_34096);
nand U34361 (N_34361,N_34044,N_34065);
or U34362 (N_34362,N_34027,N_34118);
nor U34363 (N_34363,N_34005,N_34249);
xor U34364 (N_34364,N_34111,N_34043);
or U34365 (N_34365,N_34206,N_34081);
xor U34366 (N_34366,N_34232,N_34141);
or U34367 (N_34367,N_34071,N_34140);
or U34368 (N_34368,N_34019,N_34001);
nor U34369 (N_34369,N_34105,N_34084);
nor U34370 (N_34370,N_34080,N_34230);
and U34371 (N_34371,N_34199,N_34155);
or U34372 (N_34372,N_34028,N_34134);
xor U34373 (N_34373,N_34224,N_34185);
nand U34374 (N_34374,N_34240,N_34052);
or U34375 (N_34375,N_34050,N_34034);
nand U34376 (N_34376,N_34183,N_34225);
nor U34377 (N_34377,N_34209,N_34170);
nand U34378 (N_34378,N_34112,N_34066);
nand U34379 (N_34379,N_34029,N_34002);
xnor U34380 (N_34380,N_34240,N_34155);
or U34381 (N_34381,N_34100,N_34172);
or U34382 (N_34382,N_34014,N_34133);
nand U34383 (N_34383,N_34105,N_34163);
nor U34384 (N_34384,N_34033,N_34013);
xor U34385 (N_34385,N_34019,N_34021);
nor U34386 (N_34386,N_34144,N_34165);
nand U34387 (N_34387,N_34118,N_34125);
xor U34388 (N_34388,N_34174,N_34040);
nor U34389 (N_34389,N_34086,N_34060);
and U34390 (N_34390,N_34188,N_34133);
or U34391 (N_34391,N_34234,N_34069);
and U34392 (N_34392,N_34079,N_34072);
or U34393 (N_34393,N_34055,N_34210);
or U34394 (N_34394,N_34080,N_34003);
nor U34395 (N_34395,N_34173,N_34231);
nand U34396 (N_34396,N_34117,N_34093);
nor U34397 (N_34397,N_34054,N_34076);
or U34398 (N_34398,N_34145,N_34070);
nand U34399 (N_34399,N_34211,N_34075);
nor U34400 (N_34400,N_34150,N_34160);
and U34401 (N_34401,N_34124,N_34243);
nor U34402 (N_34402,N_34182,N_34028);
xnor U34403 (N_34403,N_34228,N_34229);
nand U34404 (N_34404,N_34224,N_34032);
nor U34405 (N_34405,N_34041,N_34020);
and U34406 (N_34406,N_34226,N_34196);
nor U34407 (N_34407,N_34065,N_34013);
xor U34408 (N_34408,N_34229,N_34237);
nand U34409 (N_34409,N_34047,N_34201);
nand U34410 (N_34410,N_34109,N_34110);
nor U34411 (N_34411,N_34132,N_34151);
nand U34412 (N_34412,N_34186,N_34033);
nor U34413 (N_34413,N_34040,N_34104);
or U34414 (N_34414,N_34161,N_34121);
or U34415 (N_34415,N_34107,N_34190);
nand U34416 (N_34416,N_34053,N_34136);
nor U34417 (N_34417,N_34014,N_34162);
xnor U34418 (N_34418,N_34201,N_34023);
nand U34419 (N_34419,N_34210,N_34129);
and U34420 (N_34420,N_34093,N_34151);
nor U34421 (N_34421,N_34193,N_34052);
and U34422 (N_34422,N_34215,N_34243);
or U34423 (N_34423,N_34073,N_34001);
nand U34424 (N_34424,N_34131,N_34205);
or U34425 (N_34425,N_34168,N_34234);
nor U34426 (N_34426,N_34104,N_34056);
nor U34427 (N_34427,N_34246,N_34126);
xnor U34428 (N_34428,N_34205,N_34122);
nand U34429 (N_34429,N_34201,N_34016);
and U34430 (N_34430,N_34211,N_34173);
or U34431 (N_34431,N_34192,N_34014);
nor U34432 (N_34432,N_34185,N_34154);
and U34433 (N_34433,N_34120,N_34198);
xnor U34434 (N_34434,N_34057,N_34248);
and U34435 (N_34435,N_34197,N_34027);
xnor U34436 (N_34436,N_34012,N_34048);
or U34437 (N_34437,N_34067,N_34155);
nor U34438 (N_34438,N_34120,N_34045);
nor U34439 (N_34439,N_34018,N_34170);
nand U34440 (N_34440,N_34162,N_34025);
and U34441 (N_34441,N_34062,N_34117);
nand U34442 (N_34442,N_34014,N_34114);
xor U34443 (N_34443,N_34229,N_34192);
nor U34444 (N_34444,N_34046,N_34096);
nor U34445 (N_34445,N_34182,N_34104);
nor U34446 (N_34446,N_34044,N_34142);
and U34447 (N_34447,N_34039,N_34036);
or U34448 (N_34448,N_34186,N_34146);
xor U34449 (N_34449,N_34171,N_34227);
nor U34450 (N_34450,N_34088,N_34145);
xor U34451 (N_34451,N_34160,N_34025);
nand U34452 (N_34452,N_34219,N_34171);
or U34453 (N_34453,N_34147,N_34025);
or U34454 (N_34454,N_34228,N_34014);
and U34455 (N_34455,N_34080,N_34118);
and U34456 (N_34456,N_34076,N_34072);
and U34457 (N_34457,N_34132,N_34119);
xnor U34458 (N_34458,N_34012,N_34155);
or U34459 (N_34459,N_34096,N_34081);
nand U34460 (N_34460,N_34058,N_34069);
xnor U34461 (N_34461,N_34133,N_34234);
and U34462 (N_34462,N_34002,N_34121);
xnor U34463 (N_34463,N_34174,N_34169);
or U34464 (N_34464,N_34144,N_34199);
nor U34465 (N_34465,N_34159,N_34083);
and U34466 (N_34466,N_34032,N_34015);
xnor U34467 (N_34467,N_34157,N_34112);
or U34468 (N_34468,N_34034,N_34206);
xnor U34469 (N_34469,N_34030,N_34089);
nand U34470 (N_34470,N_34004,N_34081);
and U34471 (N_34471,N_34046,N_34127);
or U34472 (N_34472,N_34194,N_34071);
nand U34473 (N_34473,N_34237,N_34065);
nand U34474 (N_34474,N_34228,N_34102);
nor U34475 (N_34475,N_34092,N_34099);
and U34476 (N_34476,N_34132,N_34060);
xor U34477 (N_34477,N_34239,N_34211);
xnor U34478 (N_34478,N_34176,N_34006);
and U34479 (N_34479,N_34103,N_34009);
or U34480 (N_34480,N_34016,N_34244);
nor U34481 (N_34481,N_34159,N_34124);
and U34482 (N_34482,N_34197,N_34034);
xor U34483 (N_34483,N_34169,N_34017);
xnor U34484 (N_34484,N_34165,N_34180);
xor U34485 (N_34485,N_34061,N_34207);
nor U34486 (N_34486,N_34089,N_34196);
and U34487 (N_34487,N_34238,N_34094);
nor U34488 (N_34488,N_34235,N_34198);
nor U34489 (N_34489,N_34079,N_34122);
or U34490 (N_34490,N_34072,N_34181);
xor U34491 (N_34491,N_34169,N_34126);
nor U34492 (N_34492,N_34245,N_34199);
xor U34493 (N_34493,N_34188,N_34192);
nand U34494 (N_34494,N_34134,N_34160);
xor U34495 (N_34495,N_34184,N_34021);
and U34496 (N_34496,N_34095,N_34168);
and U34497 (N_34497,N_34122,N_34046);
nand U34498 (N_34498,N_34059,N_34056);
xor U34499 (N_34499,N_34163,N_34153);
nor U34500 (N_34500,N_34303,N_34493);
and U34501 (N_34501,N_34250,N_34308);
or U34502 (N_34502,N_34352,N_34478);
or U34503 (N_34503,N_34460,N_34466);
nand U34504 (N_34504,N_34347,N_34394);
xnor U34505 (N_34505,N_34360,N_34376);
nand U34506 (N_34506,N_34265,N_34491);
nor U34507 (N_34507,N_34314,N_34477);
or U34508 (N_34508,N_34448,N_34307);
or U34509 (N_34509,N_34404,N_34298);
or U34510 (N_34510,N_34379,N_34356);
xor U34511 (N_34511,N_34328,N_34251);
and U34512 (N_34512,N_34371,N_34320);
and U34513 (N_34513,N_34452,N_34361);
or U34514 (N_34514,N_34351,N_34438);
xor U34515 (N_34515,N_34369,N_34412);
or U34516 (N_34516,N_34313,N_34468);
and U34517 (N_34517,N_34318,N_34278);
nor U34518 (N_34518,N_34373,N_34286);
and U34519 (N_34519,N_34301,N_34464);
and U34520 (N_34520,N_34324,N_34270);
nor U34521 (N_34521,N_34476,N_34386);
nor U34522 (N_34522,N_34305,N_34323);
nand U34523 (N_34523,N_34418,N_34421);
or U34524 (N_34524,N_34381,N_34341);
and U34525 (N_34525,N_34374,N_34490);
and U34526 (N_34526,N_34327,N_34433);
or U34527 (N_34527,N_34407,N_34330);
or U34528 (N_34528,N_34322,N_34456);
or U34529 (N_34529,N_34359,N_34435);
nor U34530 (N_34530,N_34484,N_34317);
nand U34531 (N_34531,N_34387,N_34362);
nand U34532 (N_34532,N_34295,N_34403);
xnor U34533 (N_34533,N_34469,N_34299);
nor U34534 (N_34534,N_34385,N_34419);
nor U34535 (N_34535,N_34431,N_34458);
nor U34536 (N_34536,N_34336,N_34259);
and U34537 (N_34537,N_34400,N_34416);
nand U34538 (N_34538,N_34329,N_34348);
nand U34539 (N_34539,N_34480,N_34276);
xor U34540 (N_34540,N_34346,N_34335);
nor U34541 (N_34541,N_34383,N_34428);
and U34542 (N_34542,N_34410,N_34391);
or U34543 (N_34543,N_34274,N_34300);
nand U34544 (N_34544,N_34446,N_34289);
nand U34545 (N_34545,N_34257,N_34414);
or U34546 (N_34546,N_34467,N_34309);
or U34547 (N_34547,N_34424,N_34425);
xor U34548 (N_34548,N_34349,N_34364);
xnor U34549 (N_34549,N_34311,N_34304);
xor U34550 (N_34550,N_34489,N_34337);
and U34551 (N_34551,N_34273,N_34302);
and U34552 (N_34552,N_34409,N_34481);
xor U34553 (N_34553,N_34280,N_34454);
nand U34554 (N_34554,N_34363,N_34366);
nand U34555 (N_34555,N_34397,N_34389);
xnor U34556 (N_34556,N_34262,N_34267);
or U34557 (N_34557,N_34258,N_34457);
or U34558 (N_34558,N_34427,N_34287);
xor U34559 (N_34559,N_34297,N_34358);
and U34560 (N_34560,N_34392,N_34312);
and U34561 (N_34561,N_34370,N_34382);
or U34562 (N_34562,N_34253,N_34310);
and U34563 (N_34563,N_34332,N_34378);
or U34564 (N_34564,N_34401,N_34473);
nand U34565 (N_34565,N_34475,N_34380);
nor U34566 (N_34566,N_34499,N_34252);
xor U34567 (N_34567,N_34406,N_34331);
or U34568 (N_34568,N_34474,N_34293);
nor U34569 (N_34569,N_34461,N_34354);
nand U34570 (N_34570,N_34453,N_34445);
nor U34571 (N_34571,N_34447,N_34268);
and U34572 (N_34572,N_34260,N_34437);
and U34573 (N_34573,N_34344,N_34355);
xnor U34574 (N_34574,N_34462,N_34430);
or U34575 (N_34575,N_34282,N_34319);
xor U34576 (N_34576,N_34345,N_34256);
xnor U34577 (N_34577,N_34368,N_34492);
and U34578 (N_34578,N_34441,N_34390);
and U34579 (N_34579,N_34277,N_34488);
or U34580 (N_34580,N_34494,N_34479);
nand U34581 (N_34581,N_34439,N_34496);
nor U34582 (N_34582,N_34291,N_34316);
and U34583 (N_34583,N_34285,N_34423);
xnor U34584 (N_34584,N_34396,N_34275);
nor U34585 (N_34585,N_34436,N_34384);
nor U34586 (N_34586,N_34377,N_34372);
or U34587 (N_34587,N_34459,N_34271);
and U34588 (N_34588,N_34342,N_34325);
nand U34589 (N_34589,N_34255,N_34279);
nor U34590 (N_34590,N_34444,N_34411);
or U34591 (N_34591,N_34306,N_34450);
or U34592 (N_34592,N_34413,N_34426);
nand U34593 (N_34593,N_34284,N_34395);
xnor U34594 (N_34594,N_34497,N_34367);
nor U34595 (N_34595,N_34470,N_34290);
nand U34596 (N_34596,N_34451,N_34338);
nand U34597 (N_34597,N_34442,N_34422);
and U34598 (N_34598,N_34315,N_34402);
nand U34599 (N_34599,N_34272,N_34449);
and U34600 (N_34600,N_34487,N_34288);
nand U34601 (N_34601,N_34294,N_34333);
xor U34602 (N_34602,N_34483,N_34292);
and U34603 (N_34603,N_34440,N_34398);
nand U34604 (N_34604,N_34486,N_34434);
or U34605 (N_34605,N_34393,N_34405);
nand U34606 (N_34606,N_34485,N_34498);
nand U34607 (N_34607,N_34417,N_34388);
nand U34608 (N_34608,N_34357,N_34296);
nor U34609 (N_34609,N_34482,N_34350);
nor U34610 (N_34610,N_34334,N_34455);
nand U34611 (N_34611,N_34463,N_34415);
nor U34612 (N_34612,N_34266,N_34261);
xnor U34613 (N_34613,N_34399,N_34443);
nand U34614 (N_34614,N_34408,N_34321);
nand U34615 (N_34615,N_34429,N_34420);
and U34616 (N_34616,N_34281,N_34495);
xor U34617 (N_34617,N_34269,N_34465);
xnor U34618 (N_34618,N_34254,N_34264);
or U34619 (N_34619,N_34471,N_34339);
or U34620 (N_34620,N_34340,N_34263);
nand U34621 (N_34621,N_34472,N_34365);
and U34622 (N_34622,N_34353,N_34375);
and U34623 (N_34623,N_34343,N_34326);
xor U34624 (N_34624,N_34432,N_34283);
nand U34625 (N_34625,N_34399,N_34485);
nand U34626 (N_34626,N_34404,N_34375);
or U34627 (N_34627,N_34488,N_34377);
or U34628 (N_34628,N_34404,N_34428);
or U34629 (N_34629,N_34456,N_34403);
nand U34630 (N_34630,N_34289,N_34328);
nand U34631 (N_34631,N_34415,N_34348);
or U34632 (N_34632,N_34268,N_34408);
and U34633 (N_34633,N_34401,N_34299);
or U34634 (N_34634,N_34299,N_34460);
nor U34635 (N_34635,N_34291,N_34487);
or U34636 (N_34636,N_34494,N_34424);
or U34637 (N_34637,N_34264,N_34313);
nand U34638 (N_34638,N_34395,N_34342);
nand U34639 (N_34639,N_34320,N_34324);
xor U34640 (N_34640,N_34375,N_34293);
nand U34641 (N_34641,N_34285,N_34370);
nor U34642 (N_34642,N_34463,N_34497);
or U34643 (N_34643,N_34342,N_34483);
or U34644 (N_34644,N_34372,N_34276);
and U34645 (N_34645,N_34405,N_34429);
or U34646 (N_34646,N_34459,N_34477);
nor U34647 (N_34647,N_34475,N_34354);
or U34648 (N_34648,N_34377,N_34481);
or U34649 (N_34649,N_34260,N_34496);
nor U34650 (N_34650,N_34427,N_34344);
xor U34651 (N_34651,N_34357,N_34459);
xnor U34652 (N_34652,N_34443,N_34476);
xor U34653 (N_34653,N_34488,N_34405);
nor U34654 (N_34654,N_34338,N_34402);
nand U34655 (N_34655,N_34475,N_34366);
nand U34656 (N_34656,N_34363,N_34307);
nor U34657 (N_34657,N_34291,N_34393);
or U34658 (N_34658,N_34357,N_34276);
nor U34659 (N_34659,N_34446,N_34480);
xnor U34660 (N_34660,N_34387,N_34446);
and U34661 (N_34661,N_34422,N_34282);
or U34662 (N_34662,N_34491,N_34329);
nor U34663 (N_34663,N_34317,N_34373);
and U34664 (N_34664,N_34272,N_34419);
and U34665 (N_34665,N_34407,N_34408);
xnor U34666 (N_34666,N_34469,N_34468);
xnor U34667 (N_34667,N_34439,N_34283);
and U34668 (N_34668,N_34467,N_34438);
xor U34669 (N_34669,N_34360,N_34394);
nand U34670 (N_34670,N_34478,N_34315);
nor U34671 (N_34671,N_34355,N_34366);
and U34672 (N_34672,N_34391,N_34286);
or U34673 (N_34673,N_34307,N_34438);
nand U34674 (N_34674,N_34296,N_34431);
and U34675 (N_34675,N_34466,N_34269);
and U34676 (N_34676,N_34252,N_34390);
nand U34677 (N_34677,N_34396,N_34492);
xor U34678 (N_34678,N_34358,N_34463);
and U34679 (N_34679,N_34426,N_34330);
nand U34680 (N_34680,N_34370,N_34392);
nor U34681 (N_34681,N_34335,N_34305);
nor U34682 (N_34682,N_34266,N_34341);
or U34683 (N_34683,N_34374,N_34313);
nor U34684 (N_34684,N_34428,N_34385);
xnor U34685 (N_34685,N_34279,N_34342);
or U34686 (N_34686,N_34434,N_34326);
and U34687 (N_34687,N_34333,N_34399);
or U34688 (N_34688,N_34370,N_34380);
xor U34689 (N_34689,N_34357,N_34356);
and U34690 (N_34690,N_34295,N_34483);
nand U34691 (N_34691,N_34445,N_34438);
xor U34692 (N_34692,N_34291,N_34335);
or U34693 (N_34693,N_34414,N_34453);
nor U34694 (N_34694,N_34302,N_34437);
nor U34695 (N_34695,N_34423,N_34481);
and U34696 (N_34696,N_34491,N_34311);
or U34697 (N_34697,N_34265,N_34253);
or U34698 (N_34698,N_34297,N_34483);
nand U34699 (N_34699,N_34273,N_34438);
and U34700 (N_34700,N_34412,N_34450);
xor U34701 (N_34701,N_34303,N_34389);
and U34702 (N_34702,N_34434,N_34296);
nand U34703 (N_34703,N_34293,N_34464);
nand U34704 (N_34704,N_34350,N_34476);
and U34705 (N_34705,N_34473,N_34323);
nand U34706 (N_34706,N_34368,N_34384);
and U34707 (N_34707,N_34356,N_34304);
or U34708 (N_34708,N_34308,N_34263);
or U34709 (N_34709,N_34322,N_34371);
or U34710 (N_34710,N_34461,N_34313);
or U34711 (N_34711,N_34275,N_34317);
nor U34712 (N_34712,N_34259,N_34452);
and U34713 (N_34713,N_34377,N_34335);
and U34714 (N_34714,N_34379,N_34426);
or U34715 (N_34715,N_34425,N_34348);
or U34716 (N_34716,N_34429,N_34398);
xor U34717 (N_34717,N_34294,N_34405);
nand U34718 (N_34718,N_34431,N_34285);
and U34719 (N_34719,N_34321,N_34370);
nor U34720 (N_34720,N_34334,N_34437);
or U34721 (N_34721,N_34262,N_34391);
or U34722 (N_34722,N_34303,N_34428);
nor U34723 (N_34723,N_34316,N_34448);
nor U34724 (N_34724,N_34469,N_34496);
and U34725 (N_34725,N_34262,N_34411);
xnor U34726 (N_34726,N_34287,N_34275);
or U34727 (N_34727,N_34429,N_34356);
nor U34728 (N_34728,N_34369,N_34301);
nor U34729 (N_34729,N_34412,N_34286);
and U34730 (N_34730,N_34321,N_34300);
xnor U34731 (N_34731,N_34334,N_34294);
xnor U34732 (N_34732,N_34284,N_34291);
nor U34733 (N_34733,N_34387,N_34276);
or U34734 (N_34734,N_34482,N_34333);
xor U34735 (N_34735,N_34438,N_34490);
xor U34736 (N_34736,N_34431,N_34356);
nor U34737 (N_34737,N_34347,N_34476);
xor U34738 (N_34738,N_34377,N_34317);
xor U34739 (N_34739,N_34373,N_34293);
and U34740 (N_34740,N_34315,N_34346);
xnor U34741 (N_34741,N_34428,N_34250);
nor U34742 (N_34742,N_34364,N_34490);
xnor U34743 (N_34743,N_34448,N_34317);
and U34744 (N_34744,N_34278,N_34369);
xor U34745 (N_34745,N_34347,N_34257);
nand U34746 (N_34746,N_34298,N_34398);
and U34747 (N_34747,N_34384,N_34265);
and U34748 (N_34748,N_34342,N_34346);
or U34749 (N_34749,N_34373,N_34494);
nor U34750 (N_34750,N_34589,N_34699);
xor U34751 (N_34751,N_34576,N_34512);
and U34752 (N_34752,N_34708,N_34640);
and U34753 (N_34753,N_34710,N_34529);
nand U34754 (N_34754,N_34530,N_34527);
xor U34755 (N_34755,N_34545,N_34656);
nand U34756 (N_34756,N_34606,N_34607);
or U34757 (N_34757,N_34565,N_34732);
nand U34758 (N_34758,N_34548,N_34654);
nor U34759 (N_34759,N_34525,N_34514);
nor U34760 (N_34760,N_34676,N_34690);
and U34761 (N_34761,N_34588,N_34633);
xnor U34762 (N_34762,N_34646,N_34661);
xnor U34763 (N_34763,N_34601,N_34531);
and U34764 (N_34764,N_34556,N_34683);
nand U34765 (N_34765,N_34526,N_34700);
nor U34766 (N_34766,N_34585,N_34534);
nand U34767 (N_34767,N_34593,N_34731);
nand U34768 (N_34768,N_34546,N_34692);
and U34769 (N_34769,N_34738,N_34668);
and U34770 (N_34770,N_34521,N_34575);
or U34771 (N_34771,N_34631,N_34608);
nor U34772 (N_34772,N_34518,N_34622);
and U34773 (N_34773,N_34509,N_34727);
nand U34774 (N_34774,N_34619,N_34703);
nor U34775 (N_34775,N_34628,N_34729);
xor U34776 (N_34776,N_34748,N_34670);
xnor U34777 (N_34777,N_34691,N_34539);
nor U34778 (N_34778,N_34501,N_34567);
nand U34779 (N_34779,N_34583,N_34663);
and U34780 (N_34780,N_34693,N_34744);
nand U34781 (N_34781,N_34747,N_34624);
nor U34782 (N_34782,N_34644,N_34702);
xor U34783 (N_34783,N_34511,N_34544);
xor U34784 (N_34784,N_34714,N_34687);
xor U34785 (N_34785,N_34560,N_34620);
nor U34786 (N_34786,N_34503,N_34659);
nand U34787 (N_34787,N_34645,N_34552);
nand U34788 (N_34788,N_34508,N_34581);
xnor U34789 (N_34789,N_34516,N_34558);
nor U34790 (N_34790,N_34559,N_34502);
nor U34791 (N_34791,N_34706,N_34600);
nand U34792 (N_34792,N_34627,N_34647);
and U34793 (N_34793,N_34557,N_34705);
nor U34794 (N_34794,N_34681,N_34648);
xnor U34795 (N_34795,N_34726,N_34639);
nor U34796 (N_34796,N_34655,N_34614);
nor U34797 (N_34797,N_34717,N_34740);
xor U34798 (N_34798,N_34635,N_34570);
and U34799 (N_34799,N_34610,N_34604);
or U34800 (N_34800,N_34533,N_34672);
nor U34801 (N_34801,N_34746,N_34505);
nand U34802 (N_34802,N_34718,N_34742);
and U34803 (N_34803,N_34697,N_34674);
nand U34804 (N_34804,N_34617,N_34666);
xnor U34805 (N_34805,N_34615,N_34554);
nor U34806 (N_34806,N_34569,N_34743);
nand U34807 (N_34807,N_34724,N_34555);
nor U34808 (N_34808,N_34671,N_34688);
and U34809 (N_34809,N_34713,N_34566);
or U34810 (N_34810,N_34568,N_34586);
nor U34811 (N_34811,N_34719,N_34701);
nand U34812 (N_34812,N_34673,N_34540);
nor U34813 (N_34813,N_34504,N_34741);
nor U34814 (N_34814,N_34599,N_34720);
nor U34815 (N_34815,N_34587,N_34550);
xor U34816 (N_34816,N_34597,N_34641);
nand U34817 (N_34817,N_34669,N_34618);
xnor U34818 (N_34818,N_34651,N_34519);
nand U34819 (N_34819,N_34632,N_34577);
nor U34820 (N_34820,N_34621,N_34634);
xnor U34821 (N_34821,N_34520,N_34590);
nor U34822 (N_34822,N_34605,N_34667);
xor U34823 (N_34823,N_34517,N_34715);
xor U34824 (N_34824,N_34698,N_34513);
xnor U34825 (N_34825,N_34580,N_34642);
and U34826 (N_34826,N_34528,N_34594);
nor U34827 (N_34827,N_34596,N_34716);
xor U34828 (N_34828,N_34745,N_34660);
nand U34829 (N_34829,N_34584,N_34572);
or U34830 (N_34830,N_34707,N_34680);
nand U34831 (N_34831,N_34536,N_34662);
nand U34832 (N_34832,N_34723,N_34609);
and U34833 (N_34833,N_34679,N_34629);
nand U34834 (N_34834,N_34682,N_34562);
nand U34835 (N_34835,N_34595,N_34626);
and U34836 (N_34836,N_34721,N_34573);
or U34837 (N_34837,N_34695,N_34664);
nand U34838 (N_34838,N_34598,N_34657);
nor U34839 (N_34839,N_34563,N_34709);
nand U34840 (N_34840,N_34522,N_34547);
and U34841 (N_34841,N_34678,N_34638);
and U34842 (N_34842,N_34571,N_34650);
and U34843 (N_34843,N_34652,N_34665);
nand U34844 (N_34844,N_34549,N_34643);
and U34845 (N_34845,N_34574,N_34675);
nand U34846 (N_34846,N_34739,N_34524);
xnor U34847 (N_34847,N_34613,N_34737);
and U34848 (N_34848,N_34579,N_34735);
and U34849 (N_34849,N_34616,N_34561);
nor U34850 (N_34850,N_34553,N_34736);
nor U34851 (N_34851,N_34684,N_34612);
nor U34852 (N_34852,N_34538,N_34542);
xnor U34853 (N_34853,N_34734,N_34677);
and U34854 (N_34854,N_34686,N_34722);
xor U34855 (N_34855,N_34515,N_34653);
and U34856 (N_34856,N_34537,N_34733);
and U34857 (N_34857,N_34611,N_34535);
nor U34858 (N_34858,N_34603,N_34541);
xor U34859 (N_34859,N_34730,N_34564);
nor U34860 (N_34860,N_34532,N_34712);
xor U34861 (N_34861,N_34500,N_34704);
and U34862 (N_34862,N_34749,N_34510);
xor U34863 (N_34863,N_34592,N_34694);
nand U34864 (N_34864,N_34637,N_34506);
xor U34865 (N_34865,N_34658,N_34685);
and U34866 (N_34866,N_34689,N_34551);
and U34867 (N_34867,N_34696,N_34625);
nor U34868 (N_34868,N_34636,N_34725);
nand U34869 (N_34869,N_34649,N_34523);
xor U34870 (N_34870,N_34591,N_34507);
nor U34871 (N_34871,N_34623,N_34543);
xnor U34872 (N_34872,N_34578,N_34582);
or U34873 (N_34873,N_34728,N_34630);
or U34874 (N_34874,N_34711,N_34602);
nor U34875 (N_34875,N_34606,N_34609);
xor U34876 (N_34876,N_34679,N_34545);
nor U34877 (N_34877,N_34736,N_34709);
and U34878 (N_34878,N_34735,N_34669);
and U34879 (N_34879,N_34606,N_34526);
nor U34880 (N_34880,N_34539,N_34538);
nand U34881 (N_34881,N_34628,N_34690);
nand U34882 (N_34882,N_34535,N_34515);
nand U34883 (N_34883,N_34624,N_34556);
or U34884 (N_34884,N_34594,N_34687);
xnor U34885 (N_34885,N_34703,N_34554);
or U34886 (N_34886,N_34500,N_34610);
nor U34887 (N_34887,N_34500,N_34640);
nor U34888 (N_34888,N_34534,N_34500);
xnor U34889 (N_34889,N_34698,N_34701);
nand U34890 (N_34890,N_34742,N_34568);
xnor U34891 (N_34891,N_34537,N_34737);
nand U34892 (N_34892,N_34585,N_34616);
nor U34893 (N_34893,N_34704,N_34692);
nand U34894 (N_34894,N_34641,N_34721);
or U34895 (N_34895,N_34562,N_34667);
and U34896 (N_34896,N_34548,N_34526);
or U34897 (N_34897,N_34717,N_34635);
and U34898 (N_34898,N_34589,N_34707);
nor U34899 (N_34899,N_34625,N_34526);
or U34900 (N_34900,N_34739,N_34713);
xor U34901 (N_34901,N_34663,N_34609);
or U34902 (N_34902,N_34692,N_34586);
nand U34903 (N_34903,N_34613,N_34533);
nor U34904 (N_34904,N_34537,N_34605);
nand U34905 (N_34905,N_34639,N_34550);
nand U34906 (N_34906,N_34613,N_34749);
nand U34907 (N_34907,N_34599,N_34593);
nor U34908 (N_34908,N_34592,N_34702);
nand U34909 (N_34909,N_34662,N_34712);
nor U34910 (N_34910,N_34653,N_34621);
xnor U34911 (N_34911,N_34733,N_34633);
nor U34912 (N_34912,N_34747,N_34686);
and U34913 (N_34913,N_34627,N_34745);
xor U34914 (N_34914,N_34594,N_34616);
and U34915 (N_34915,N_34567,N_34564);
or U34916 (N_34916,N_34672,N_34709);
nor U34917 (N_34917,N_34733,N_34611);
nor U34918 (N_34918,N_34738,N_34725);
xnor U34919 (N_34919,N_34634,N_34581);
and U34920 (N_34920,N_34632,N_34736);
and U34921 (N_34921,N_34659,N_34715);
or U34922 (N_34922,N_34681,N_34527);
or U34923 (N_34923,N_34639,N_34585);
and U34924 (N_34924,N_34748,N_34677);
xor U34925 (N_34925,N_34666,N_34736);
or U34926 (N_34926,N_34643,N_34587);
xnor U34927 (N_34927,N_34582,N_34657);
or U34928 (N_34928,N_34689,N_34695);
nand U34929 (N_34929,N_34565,N_34536);
or U34930 (N_34930,N_34638,N_34597);
or U34931 (N_34931,N_34678,N_34582);
xnor U34932 (N_34932,N_34735,N_34596);
or U34933 (N_34933,N_34683,N_34689);
xnor U34934 (N_34934,N_34667,N_34549);
nor U34935 (N_34935,N_34729,N_34509);
xor U34936 (N_34936,N_34564,N_34714);
nor U34937 (N_34937,N_34611,N_34742);
nor U34938 (N_34938,N_34705,N_34505);
or U34939 (N_34939,N_34518,N_34546);
and U34940 (N_34940,N_34699,N_34605);
nand U34941 (N_34941,N_34663,N_34568);
nor U34942 (N_34942,N_34716,N_34669);
nand U34943 (N_34943,N_34534,N_34647);
nand U34944 (N_34944,N_34512,N_34589);
nand U34945 (N_34945,N_34717,N_34603);
xor U34946 (N_34946,N_34680,N_34668);
and U34947 (N_34947,N_34722,N_34683);
nand U34948 (N_34948,N_34526,N_34600);
xnor U34949 (N_34949,N_34736,N_34611);
nand U34950 (N_34950,N_34611,N_34565);
xor U34951 (N_34951,N_34583,N_34660);
or U34952 (N_34952,N_34604,N_34587);
nor U34953 (N_34953,N_34737,N_34579);
nand U34954 (N_34954,N_34583,N_34504);
xnor U34955 (N_34955,N_34559,N_34614);
nand U34956 (N_34956,N_34524,N_34605);
and U34957 (N_34957,N_34620,N_34604);
and U34958 (N_34958,N_34680,N_34500);
nand U34959 (N_34959,N_34688,N_34716);
or U34960 (N_34960,N_34742,N_34580);
and U34961 (N_34961,N_34642,N_34582);
and U34962 (N_34962,N_34568,N_34602);
nor U34963 (N_34963,N_34559,N_34582);
or U34964 (N_34964,N_34546,N_34648);
or U34965 (N_34965,N_34549,N_34642);
xnor U34966 (N_34966,N_34577,N_34560);
and U34967 (N_34967,N_34515,N_34615);
nor U34968 (N_34968,N_34637,N_34596);
nand U34969 (N_34969,N_34677,N_34700);
and U34970 (N_34970,N_34561,N_34647);
xnor U34971 (N_34971,N_34612,N_34575);
nand U34972 (N_34972,N_34544,N_34509);
xor U34973 (N_34973,N_34749,N_34692);
xnor U34974 (N_34974,N_34745,N_34515);
nor U34975 (N_34975,N_34713,N_34529);
nor U34976 (N_34976,N_34593,N_34640);
or U34977 (N_34977,N_34628,N_34700);
xor U34978 (N_34978,N_34607,N_34608);
and U34979 (N_34979,N_34628,N_34592);
and U34980 (N_34980,N_34742,N_34625);
xnor U34981 (N_34981,N_34693,N_34517);
or U34982 (N_34982,N_34574,N_34535);
nor U34983 (N_34983,N_34656,N_34668);
xor U34984 (N_34984,N_34558,N_34694);
and U34985 (N_34985,N_34607,N_34541);
xor U34986 (N_34986,N_34620,N_34719);
nor U34987 (N_34987,N_34747,N_34597);
nand U34988 (N_34988,N_34509,N_34656);
nor U34989 (N_34989,N_34639,N_34692);
nand U34990 (N_34990,N_34570,N_34551);
nor U34991 (N_34991,N_34513,N_34655);
xnor U34992 (N_34992,N_34503,N_34686);
xor U34993 (N_34993,N_34713,N_34621);
or U34994 (N_34994,N_34673,N_34618);
nand U34995 (N_34995,N_34720,N_34592);
and U34996 (N_34996,N_34701,N_34517);
nand U34997 (N_34997,N_34502,N_34673);
nor U34998 (N_34998,N_34601,N_34542);
or U34999 (N_34999,N_34731,N_34685);
or U35000 (N_35000,N_34998,N_34898);
or U35001 (N_35001,N_34844,N_34897);
nand U35002 (N_35002,N_34801,N_34896);
or U35003 (N_35003,N_34935,N_34957);
or U35004 (N_35004,N_34759,N_34977);
or U35005 (N_35005,N_34785,N_34754);
nand U35006 (N_35006,N_34944,N_34925);
and U35007 (N_35007,N_34988,N_34903);
nand U35008 (N_35008,N_34871,N_34763);
xor U35009 (N_35009,N_34830,N_34956);
xor U35010 (N_35010,N_34932,N_34953);
nand U35011 (N_35011,N_34765,N_34908);
or U35012 (N_35012,N_34824,N_34779);
nand U35013 (N_35013,N_34979,N_34974);
nand U35014 (N_35014,N_34773,N_34946);
xor U35015 (N_35015,N_34873,N_34997);
nor U35016 (N_35016,N_34943,N_34876);
xor U35017 (N_35017,N_34942,N_34808);
nand U35018 (N_35018,N_34756,N_34975);
or U35019 (N_35019,N_34955,N_34827);
and U35020 (N_35020,N_34775,N_34973);
nand U35021 (N_35021,N_34845,N_34854);
nand U35022 (N_35022,N_34926,N_34774);
nor U35023 (N_35023,N_34812,N_34852);
nand U35024 (N_35024,N_34762,N_34848);
xor U35025 (N_35025,N_34869,N_34795);
or U35026 (N_35026,N_34923,N_34856);
nand U35027 (N_35027,N_34823,N_34863);
nand U35028 (N_35028,N_34888,N_34833);
and U35029 (N_35029,N_34770,N_34791);
or U35030 (N_35030,N_34821,N_34790);
and U35031 (N_35031,N_34799,N_34987);
nor U35032 (N_35032,N_34906,N_34950);
or U35033 (N_35033,N_34877,N_34990);
or U35034 (N_35034,N_34834,N_34940);
or U35035 (N_35035,N_34776,N_34855);
nand U35036 (N_35036,N_34819,N_34794);
nor U35037 (N_35037,N_34996,N_34914);
or U35038 (N_35038,N_34933,N_34802);
or U35039 (N_35039,N_34798,N_34969);
nor U35040 (N_35040,N_34899,N_34751);
xnor U35041 (N_35041,N_34951,N_34980);
and U35042 (N_35042,N_34900,N_34894);
or U35043 (N_35043,N_34954,N_34864);
xor U35044 (N_35044,N_34850,N_34991);
xor U35045 (N_35045,N_34915,N_34804);
nand U35046 (N_35046,N_34928,N_34966);
nor U35047 (N_35047,N_34868,N_34766);
nand U35048 (N_35048,N_34875,N_34931);
nand U35049 (N_35049,N_34919,N_34921);
xnor U35050 (N_35050,N_34971,N_34891);
or U35051 (N_35051,N_34916,N_34907);
or U35052 (N_35052,N_34853,N_34828);
nand U35053 (N_35053,N_34889,N_34959);
or U35054 (N_35054,N_34930,N_34994);
or U35055 (N_35055,N_34968,N_34895);
nand U35056 (N_35056,N_34836,N_34878);
nor U35057 (N_35057,N_34870,N_34818);
xor U35058 (N_35058,N_34769,N_34961);
xor U35059 (N_35059,N_34885,N_34767);
xor U35060 (N_35060,N_34781,N_34780);
xnor U35061 (N_35061,N_34841,N_34913);
or U35062 (N_35062,N_34760,N_34901);
nor U35063 (N_35063,N_34874,N_34938);
or U35064 (N_35064,N_34814,N_34800);
and U35065 (N_35065,N_34792,N_34811);
and U35066 (N_35066,N_34945,N_34887);
and U35067 (N_35067,N_34832,N_34934);
nor U35068 (N_35068,N_34886,N_34796);
nand U35069 (N_35069,N_34778,N_34866);
nand U35070 (N_35070,N_34872,N_34829);
and U35071 (N_35071,N_34839,N_34806);
nand U35072 (N_35072,N_34840,N_34793);
xnor U35073 (N_35073,N_34993,N_34985);
and U35074 (N_35074,N_34826,N_34999);
or U35075 (N_35075,N_34758,N_34964);
nand U35076 (N_35076,N_34947,N_34761);
nand U35077 (N_35077,N_34882,N_34904);
nor U35078 (N_35078,N_34797,N_34861);
nor U35079 (N_35079,N_34867,N_34757);
or U35080 (N_35080,N_34843,N_34958);
nor U35081 (N_35081,N_34965,N_34883);
nor U35082 (N_35082,N_34936,N_34815);
nand U35083 (N_35083,N_34817,N_34978);
nand U35084 (N_35084,N_34851,N_34929);
nand U35085 (N_35085,N_34807,N_34948);
nor U35086 (N_35086,N_34995,N_34847);
xor U35087 (N_35087,N_34941,N_34949);
and U35088 (N_35088,N_34838,N_34837);
nand U35089 (N_35089,N_34820,N_34983);
nand U35090 (N_35090,N_34859,N_34918);
or U35091 (N_35091,N_34816,N_34972);
nand U35092 (N_35092,N_34805,N_34772);
or U35093 (N_35093,N_34911,N_34777);
xor U35094 (N_35094,N_34976,N_34917);
nand U35095 (N_35095,N_34902,N_34753);
nand U35096 (N_35096,N_34784,N_34989);
nor U35097 (N_35097,N_34860,N_34842);
nand U35098 (N_35098,N_34884,N_34986);
nor U35099 (N_35099,N_34835,N_34893);
and U35100 (N_35100,N_34825,N_34822);
and U35101 (N_35101,N_34922,N_34831);
xnor U35102 (N_35102,N_34771,N_34857);
and U35103 (N_35103,N_34892,N_34810);
xor U35104 (N_35104,N_34879,N_34984);
or U35105 (N_35105,N_34755,N_34960);
xnor U35106 (N_35106,N_34786,N_34783);
xnor U35107 (N_35107,N_34937,N_34846);
or U35108 (N_35108,N_34813,N_34880);
xor U35109 (N_35109,N_34768,N_34858);
nor U35110 (N_35110,N_34962,N_34981);
xnor U35111 (N_35111,N_34803,N_34782);
xnor U35112 (N_35112,N_34912,N_34952);
nand U35113 (N_35113,N_34924,N_34927);
and U35114 (N_35114,N_34909,N_34920);
nand U35115 (N_35115,N_34881,N_34849);
nand U35116 (N_35116,N_34764,N_34890);
xor U35117 (N_35117,N_34865,N_34862);
nand U35118 (N_35118,N_34789,N_34982);
nor U35119 (N_35119,N_34809,N_34963);
nor U35120 (N_35120,N_34905,N_34787);
and U35121 (N_35121,N_34750,N_34970);
and U35122 (N_35122,N_34992,N_34910);
xor U35123 (N_35123,N_34752,N_34788);
xnor U35124 (N_35124,N_34967,N_34939);
and U35125 (N_35125,N_34900,N_34973);
and U35126 (N_35126,N_34898,N_34892);
and U35127 (N_35127,N_34789,N_34814);
and U35128 (N_35128,N_34924,N_34790);
or U35129 (N_35129,N_34762,N_34992);
or U35130 (N_35130,N_34806,N_34753);
nand U35131 (N_35131,N_34804,N_34765);
and U35132 (N_35132,N_34872,N_34851);
nor U35133 (N_35133,N_34944,N_34993);
xor U35134 (N_35134,N_34773,N_34890);
nand U35135 (N_35135,N_34821,N_34916);
nand U35136 (N_35136,N_34790,N_34777);
and U35137 (N_35137,N_34939,N_34799);
xor U35138 (N_35138,N_34895,N_34773);
and U35139 (N_35139,N_34885,N_34810);
nand U35140 (N_35140,N_34960,N_34933);
or U35141 (N_35141,N_34924,N_34831);
xnor U35142 (N_35142,N_34888,N_34889);
or U35143 (N_35143,N_34864,N_34817);
nand U35144 (N_35144,N_34820,N_34779);
nor U35145 (N_35145,N_34772,N_34798);
nor U35146 (N_35146,N_34936,N_34779);
and U35147 (N_35147,N_34978,N_34823);
or U35148 (N_35148,N_34920,N_34767);
or U35149 (N_35149,N_34853,N_34894);
xnor U35150 (N_35150,N_34756,N_34842);
or U35151 (N_35151,N_34758,N_34875);
nor U35152 (N_35152,N_34905,N_34853);
or U35153 (N_35153,N_34823,N_34801);
or U35154 (N_35154,N_34888,N_34890);
nand U35155 (N_35155,N_34781,N_34816);
or U35156 (N_35156,N_34981,N_34761);
nor U35157 (N_35157,N_34836,N_34819);
xor U35158 (N_35158,N_34918,N_34952);
nor U35159 (N_35159,N_34933,N_34983);
nor U35160 (N_35160,N_34778,N_34895);
nor U35161 (N_35161,N_34929,N_34801);
nand U35162 (N_35162,N_34818,N_34813);
or U35163 (N_35163,N_34996,N_34811);
nor U35164 (N_35164,N_34979,N_34999);
xor U35165 (N_35165,N_34824,N_34759);
xnor U35166 (N_35166,N_34957,N_34971);
or U35167 (N_35167,N_34897,N_34946);
xor U35168 (N_35168,N_34843,N_34828);
nor U35169 (N_35169,N_34909,N_34810);
and U35170 (N_35170,N_34893,N_34856);
nor U35171 (N_35171,N_34899,N_34880);
xnor U35172 (N_35172,N_34815,N_34846);
xnor U35173 (N_35173,N_34890,N_34820);
nor U35174 (N_35174,N_34982,N_34983);
nor U35175 (N_35175,N_34835,N_34770);
nand U35176 (N_35176,N_34881,N_34950);
nor U35177 (N_35177,N_34959,N_34963);
or U35178 (N_35178,N_34814,N_34909);
nand U35179 (N_35179,N_34807,N_34816);
and U35180 (N_35180,N_34760,N_34959);
nor U35181 (N_35181,N_34884,N_34843);
nand U35182 (N_35182,N_34837,N_34955);
nor U35183 (N_35183,N_34868,N_34768);
and U35184 (N_35184,N_34774,N_34798);
nor U35185 (N_35185,N_34988,N_34927);
or U35186 (N_35186,N_34974,N_34934);
nand U35187 (N_35187,N_34895,N_34906);
or U35188 (N_35188,N_34803,N_34770);
or U35189 (N_35189,N_34988,N_34965);
and U35190 (N_35190,N_34908,N_34805);
nand U35191 (N_35191,N_34761,N_34915);
and U35192 (N_35192,N_34999,N_34905);
nor U35193 (N_35193,N_34768,N_34767);
nor U35194 (N_35194,N_34788,N_34960);
xor U35195 (N_35195,N_34937,N_34887);
nand U35196 (N_35196,N_34764,N_34875);
or U35197 (N_35197,N_34891,N_34963);
xor U35198 (N_35198,N_34805,N_34794);
nand U35199 (N_35199,N_34838,N_34984);
nand U35200 (N_35200,N_34816,N_34856);
nand U35201 (N_35201,N_34996,N_34772);
nor U35202 (N_35202,N_34867,N_34927);
or U35203 (N_35203,N_34841,N_34842);
and U35204 (N_35204,N_34977,N_34984);
xor U35205 (N_35205,N_34946,N_34909);
and U35206 (N_35206,N_34881,N_34934);
nor U35207 (N_35207,N_34915,N_34842);
and U35208 (N_35208,N_34981,N_34853);
and U35209 (N_35209,N_34950,N_34980);
nor U35210 (N_35210,N_34780,N_34811);
xor U35211 (N_35211,N_34910,N_34950);
nand U35212 (N_35212,N_34802,N_34841);
xnor U35213 (N_35213,N_34959,N_34770);
and U35214 (N_35214,N_34923,N_34917);
nand U35215 (N_35215,N_34955,N_34788);
and U35216 (N_35216,N_34896,N_34780);
xor U35217 (N_35217,N_34962,N_34895);
xnor U35218 (N_35218,N_34825,N_34931);
and U35219 (N_35219,N_34931,N_34841);
nor U35220 (N_35220,N_34981,N_34910);
nor U35221 (N_35221,N_34983,N_34763);
and U35222 (N_35222,N_34859,N_34929);
xor U35223 (N_35223,N_34773,N_34889);
nor U35224 (N_35224,N_34919,N_34838);
nand U35225 (N_35225,N_34845,N_34918);
nand U35226 (N_35226,N_34771,N_34942);
and U35227 (N_35227,N_34813,N_34781);
xnor U35228 (N_35228,N_34800,N_34774);
xnor U35229 (N_35229,N_34794,N_34849);
and U35230 (N_35230,N_34918,N_34837);
xnor U35231 (N_35231,N_34963,N_34987);
and U35232 (N_35232,N_34793,N_34785);
nand U35233 (N_35233,N_34833,N_34794);
or U35234 (N_35234,N_34885,N_34796);
nand U35235 (N_35235,N_34857,N_34886);
nor U35236 (N_35236,N_34893,N_34956);
nor U35237 (N_35237,N_34805,N_34776);
nand U35238 (N_35238,N_34864,N_34994);
and U35239 (N_35239,N_34771,N_34900);
or U35240 (N_35240,N_34943,N_34890);
nand U35241 (N_35241,N_34870,N_34918);
and U35242 (N_35242,N_34961,N_34872);
or U35243 (N_35243,N_34981,N_34803);
and U35244 (N_35244,N_34997,N_34853);
and U35245 (N_35245,N_34945,N_34818);
nor U35246 (N_35246,N_34876,N_34924);
or U35247 (N_35247,N_34869,N_34959);
nand U35248 (N_35248,N_34870,N_34788);
nor U35249 (N_35249,N_34775,N_34948);
and U35250 (N_35250,N_35182,N_35049);
nor U35251 (N_35251,N_35026,N_35162);
nand U35252 (N_35252,N_35186,N_35230);
or U35253 (N_35253,N_35236,N_35194);
or U35254 (N_35254,N_35138,N_35040);
or U35255 (N_35255,N_35094,N_35000);
nor U35256 (N_35256,N_35131,N_35222);
nand U35257 (N_35257,N_35060,N_35013);
or U35258 (N_35258,N_35238,N_35103);
or U35259 (N_35259,N_35037,N_35050);
or U35260 (N_35260,N_35226,N_35036);
nand U35261 (N_35261,N_35132,N_35052);
nor U35262 (N_35262,N_35201,N_35137);
nor U35263 (N_35263,N_35108,N_35122);
or U35264 (N_35264,N_35002,N_35027);
or U35265 (N_35265,N_35213,N_35224);
xnor U35266 (N_35266,N_35187,N_35214);
nand U35267 (N_35267,N_35078,N_35051);
nor U35268 (N_35268,N_35090,N_35130);
nand U35269 (N_35269,N_35133,N_35202);
xnor U35270 (N_35270,N_35030,N_35123);
nor U35271 (N_35271,N_35128,N_35159);
xor U35272 (N_35272,N_35129,N_35047);
xnor U35273 (N_35273,N_35173,N_35117);
and U35274 (N_35274,N_35001,N_35134);
xnor U35275 (N_35275,N_35121,N_35168);
nand U35276 (N_35276,N_35033,N_35032);
or U35277 (N_35277,N_35116,N_35160);
nor U35278 (N_35278,N_35124,N_35091);
nor U35279 (N_35279,N_35196,N_35095);
nand U35280 (N_35280,N_35198,N_35206);
nand U35281 (N_35281,N_35003,N_35061);
and U35282 (N_35282,N_35241,N_35034);
and U35283 (N_35283,N_35158,N_35176);
and U35284 (N_35284,N_35195,N_35055);
and U35285 (N_35285,N_35208,N_35150);
and U35286 (N_35286,N_35164,N_35125);
and U35287 (N_35287,N_35192,N_35212);
and U35288 (N_35288,N_35197,N_35035);
nor U35289 (N_35289,N_35139,N_35245);
nor U35290 (N_35290,N_35070,N_35081);
xor U35291 (N_35291,N_35048,N_35063);
and U35292 (N_35292,N_35087,N_35244);
xnor U35293 (N_35293,N_35011,N_35009);
and U35294 (N_35294,N_35235,N_35025);
or U35295 (N_35295,N_35233,N_35210);
nand U35296 (N_35296,N_35079,N_35056);
nor U35297 (N_35297,N_35120,N_35215);
nor U35298 (N_35298,N_35046,N_35077);
nand U35299 (N_35299,N_35080,N_35172);
and U35300 (N_35300,N_35118,N_35152);
nor U35301 (N_35301,N_35200,N_35175);
nor U35302 (N_35302,N_35086,N_35064);
and U35303 (N_35303,N_35005,N_35031);
xnor U35304 (N_35304,N_35219,N_35184);
xor U35305 (N_35305,N_35004,N_35098);
or U35306 (N_35306,N_35107,N_35148);
or U35307 (N_35307,N_35045,N_35190);
xnor U35308 (N_35308,N_35147,N_35217);
xnor U35309 (N_35309,N_35240,N_35113);
nand U35310 (N_35310,N_35069,N_35073);
nor U35311 (N_35311,N_35163,N_35075);
and U35312 (N_35312,N_35178,N_35015);
xor U35313 (N_35313,N_35022,N_35119);
or U35314 (N_35314,N_35174,N_35211);
nand U35315 (N_35315,N_35010,N_35221);
nor U35316 (N_35316,N_35074,N_35076);
or U35317 (N_35317,N_35191,N_35145);
and U35318 (N_35318,N_35024,N_35223);
and U35319 (N_35319,N_35023,N_35249);
xor U35320 (N_35320,N_35006,N_35007);
xnor U35321 (N_35321,N_35114,N_35171);
nor U35322 (N_35322,N_35154,N_35146);
and U35323 (N_35323,N_35029,N_35089);
and U35324 (N_35324,N_35067,N_35109);
and U35325 (N_35325,N_35209,N_35143);
or U35326 (N_35326,N_35066,N_35220);
nor U35327 (N_35327,N_35115,N_35028);
or U35328 (N_35328,N_35068,N_35096);
xnor U35329 (N_35329,N_35093,N_35082);
or U35330 (N_35330,N_35232,N_35228);
and U35331 (N_35331,N_35016,N_35084);
or U35332 (N_35332,N_35193,N_35019);
or U35333 (N_35333,N_35088,N_35183);
xnor U35334 (N_35334,N_35065,N_35097);
and U35335 (N_35335,N_35042,N_35207);
nand U35336 (N_35336,N_35165,N_35179);
nor U35337 (N_35337,N_35057,N_35083);
nor U35338 (N_35338,N_35018,N_35218);
and U35339 (N_35339,N_35140,N_35099);
nor U35340 (N_35340,N_35041,N_35169);
nor U35341 (N_35341,N_35038,N_35102);
nor U35342 (N_35342,N_35092,N_35141);
nand U35343 (N_35343,N_35151,N_35106);
xnor U35344 (N_35344,N_35177,N_35142);
xnor U35345 (N_35345,N_35237,N_35020);
nor U35346 (N_35346,N_35216,N_35021);
nand U35347 (N_35347,N_35144,N_35100);
or U35348 (N_35348,N_35242,N_35110);
nor U35349 (N_35349,N_35205,N_35234);
or U35350 (N_35350,N_35204,N_35229);
xor U35351 (N_35351,N_35188,N_35085);
nand U35352 (N_35352,N_35246,N_35185);
and U35353 (N_35353,N_35072,N_35062);
or U35354 (N_35354,N_35059,N_35227);
and U35355 (N_35355,N_35112,N_35189);
or U35356 (N_35356,N_35135,N_35149);
nor U35357 (N_35357,N_35156,N_35231);
nand U35358 (N_35358,N_35039,N_35225);
xnor U35359 (N_35359,N_35105,N_35111);
and U35360 (N_35360,N_35053,N_35248);
nor U35361 (N_35361,N_35180,N_35104);
and U35362 (N_35362,N_35199,N_35181);
or U35363 (N_35363,N_35044,N_35167);
nand U35364 (N_35364,N_35170,N_35126);
or U35365 (N_35365,N_35043,N_35136);
and U35366 (N_35366,N_35054,N_35012);
or U35367 (N_35367,N_35157,N_35008);
and U35368 (N_35368,N_35101,N_35014);
nor U35369 (N_35369,N_35058,N_35071);
xnor U35370 (N_35370,N_35239,N_35017);
and U35371 (N_35371,N_35127,N_35247);
nand U35372 (N_35372,N_35153,N_35203);
nor U35373 (N_35373,N_35161,N_35166);
nor U35374 (N_35374,N_35155,N_35243);
nor U35375 (N_35375,N_35228,N_35155);
or U35376 (N_35376,N_35042,N_35118);
nor U35377 (N_35377,N_35101,N_35194);
or U35378 (N_35378,N_35226,N_35139);
nor U35379 (N_35379,N_35216,N_35186);
xor U35380 (N_35380,N_35247,N_35091);
xor U35381 (N_35381,N_35187,N_35062);
xnor U35382 (N_35382,N_35231,N_35061);
nand U35383 (N_35383,N_35066,N_35075);
nand U35384 (N_35384,N_35228,N_35082);
and U35385 (N_35385,N_35040,N_35046);
nand U35386 (N_35386,N_35142,N_35147);
and U35387 (N_35387,N_35243,N_35134);
xor U35388 (N_35388,N_35027,N_35188);
xor U35389 (N_35389,N_35232,N_35086);
nor U35390 (N_35390,N_35048,N_35169);
xnor U35391 (N_35391,N_35063,N_35031);
and U35392 (N_35392,N_35177,N_35156);
nor U35393 (N_35393,N_35026,N_35014);
or U35394 (N_35394,N_35129,N_35113);
or U35395 (N_35395,N_35186,N_35183);
xnor U35396 (N_35396,N_35205,N_35089);
nand U35397 (N_35397,N_35199,N_35042);
nand U35398 (N_35398,N_35106,N_35038);
and U35399 (N_35399,N_35108,N_35199);
or U35400 (N_35400,N_35123,N_35216);
or U35401 (N_35401,N_35196,N_35014);
nor U35402 (N_35402,N_35097,N_35124);
nand U35403 (N_35403,N_35166,N_35234);
or U35404 (N_35404,N_35207,N_35194);
nand U35405 (N_35405,N_35212,N_35175);
nand U35406 (N_35406,N_35173,N_35062);
xor U35407 (N_35407,N_35136,N_35091);
nor U35408 (N_35408,N_35214,N_35210);
nand U35409 (N_35409,N_35245,N_35132);
nor U35410 (N_35410,N_35056,N_35147);
nor U35411 (N_35411,N_35210,N_35149);
or U35412 (N_35412,N_35219,N_35202);
xor U35413 (N_35413,N_35222,N_35091);
nor U35414 (N_35414,N_35090,N_35122);
nand U35415 (N_35415,N_35132,N_35107);
and U35416 (N_35416,N_35142,N_35018);
nor U35417 (N_35417,N_35064,N_35101);
nand U35418 (N_35418,N_35238,N_35015);
and U35419 (N_35419,N_35137,N_35195);
or U35420 (N_35420,N_35204,N_35238);
or U35421 (N_35421,N_35225,N_35246);
xnor U35422 (N_35422,N_35085,N_35121);
or U35423 (N_35423,N_35096,N_35217);
or U35424 (N_35424,N_35231,N_35027);
or U35425 (N_35425,N_35078,N_35034);
nor U35426 (N_35426,N_35016,N_35135);
or U35427 (N_35427,N_35116,N_35220);
nor U35428 (N_35428,N_35193,N_35101);
nand U35429 (N_35429,N_35235,N_35073);
xor U35430 (N_35430,N_35080,N_35191);
and U35431 (N_35431,N_35143,N_35142);
and U35432 (N_35432,N_35037,N_35129);
nor U35433 (N_35433,N_35091,N_35180);
nand U35434 (N_35434,N_35017,N_35059);
nor U35435 (N_35435,N_35120,N_35007);
nor U35436 (N_35436,N_35189,N_35160);
or U35437 (N_35437,N_35039,N_35230);
xnor U35438 (N_35438,N_35243,N_35028);
nand U35439 (N_35439,N_35238,N_35003);
and U35440 (N_35440,N_35047,N_35148);
or U35441 (N_35441,N_35157,N_35147);
xnor U35442 (N_35442,N_35083,N_35149);
or U35443 (N_35443,N_35027,N_35222);
nor U35444 (N_35444,N_35147,N_35213);
xnor U35445 (N_35445,N_35037,N_35008);
and U35446 (N_35446,N_35040,N_35025);
nor U35447 (N_35447,N_35148,N_35109);
or U35448 (N_35448,N_35234,N_35035);
nand U35449 (N_35449,N_35028,N_35187);
nand U35450 (N_35450,N_35069,N_35136);
nor U35451 (N_35451,N_35159,N_35165);
or U35452 (N_35452,N_35230,N_35018);
nand U35453 (N_35453,N_35092,N_35080);
nor U35454 (N_35454,N_35247,N_35171);
xnor U35455 (N_35455,N_35026,N_35088);
nand U35456 (N_35456,N_35189,N_35222);
nor U35457 (N_35457,N_35246,N_35180);
and U35458 (N_35458,N_35222,N_35144);
nand U35459 (N_35459,N_35064,N_35239);
xor U35460 (N_35460,N_35023,N_35025);
or U35461 (N_35461,N_35167,N_35151);
or U35462 (N_35462,N_35065,N_35158);
nand U35463 (N_35463,N_35095,N_35159);
and U35464 (N_35464,N_35047,N_35178);
xor U35465 (N_35465,N_35227,N_35237);
or U35466 (N_35466,N_35009,N_35031);
or U35467 (N_35467,N_35002,N_35105);
nor U35468 (N_35468,N_35020,N_35184);
xnor U35469 (N_35469,N_35027,N_35169);
nand U35470 (N_35470,N_35028,N_35058);
or U35471 (N_35471,N_35168,N_35058);
nor U35472 (N_35472,N_35214,N_35085);
nor U35473 (N_35473,N_35070,N_35079);
xnor U35474 (N_35474,N_35232,N_35236);
nor U35475 (N_35475,N_35186,N_35247);
nor U35476 (N_35476,N_35038,N_35126);
xor U35477 (N_35477,N_35233,N_35216);
xnor U35478 (N_35478,N_35083,N_35198);
nor U35479 (N_35479,N_35226,N_35076);
or U35480 (N_35480,N_35034,N_35011);
nor U35481 (N_35481,N_35237,N_35126);
and U35482 (N_35482,N_35107,N_35207);
xnor U35483 (N_35483,N_35050,N_35109);
xor U35484 (N_35484,N_35228,N_35075);
and U35485 (N_35485,N_35192,N_35165);
xnor U35486 (N_35486,N_35046,N_35130);
xor U35487 (N_35487,N_35121,N_35166);
xor U35488 (N_35488,N_35086,N_35012);
and U35489 (N_35489,N_35174,N_35129);
nand U35490 (N_35490,N_35109,N_35203);
nor U35491 (N_35491,N_35033,N_35135);
and U35492 (N_35492,N_35089,N_35007);
nor U35493 (N_35493,N_35046,N_35179);
or U35494 (N_35494,N_35233,N_35120);
or U35495 (N_35495,N_35151,N_35233);
nor U35496 (N_35496,N_35012,N_35221);
or U35497 (N_35497,N_35162,N_35078);
xor U35498 (N_35498,N_35116,N_35015);
or U35499 (N_35499,N_35023,N_35014);
or U35500 (N_35500,N_35343,N_35283);
or U35501 (N_35501,N_35375,N_35323);
or U35502 (N_35502,N_35463,N_35392);
or U35503 (N_35503,N_35475,N_35439);
or U35504 (N_35504,N_35272,N_35423);
and U35505 (N_35505,N_35438,N_35450);
and U35506 (N_35506,N_35326,N_35321);
nand U35507 (N_35507,N_35490,N_35338);
or U35508 (N_35508,N_35266,N_35270);
or U35509 (N_35509,N_35268,N_35496);
or U35510 (N_35510,N_35421,N_35355);
and U35511 (N_35511,N_35431,N_35377);
and U35512 (N_35512,N_35342,N_35444);
nand U35513 (N_35513,N_35498,N_35330);
xor U35514 (N_35514,N_35310,N_35406);
or U35515 (N_35515,N_35373,N_35331);
and U35516 (N_35516,N_35484,N_35488);
or U35517 (N_35517,N_35411,N_35339);
or U35518 (N_35518,N_35404,N_35472);
and U35519 (N_35519,N_35297,N_35401);
nor U35520 (N_35520,N_35288,N_35362);
or U35521 (N_35521,N_35378,N_35263);
nand U35522 (N_35522,N_35400,N_35491);
or U35523 (N_35523,N_35391,N_35478);
or U35524 (N_35524,N_35258,N_35264);
nor U35525 (N_35525,N_35482,N_35437);
or U35526 (N_35526,N_35398,N_35254);
and U35527 (N_35527,N_35471,N_35273);
nand U35528 (N_35528,N_35267,N_35379);
nor U35529 (N_35529,N_35269,N_35413);
nand U35530 (N_35530,N_35376,N_35418);
nor U35531 (N_35531,N_35280,N_35356);
or U35532 (N_35532,N_35306,N_35276);
xor U35533 (N_35533,N_35260,N_35299);
or U35534 (N_35534,N_35345,N_35485);
nor U35535 (N_35535,N_35460,N_35387);
nor U35536 (N_35536,N_35317,N_35452);
xor U35537 (N_35537,N_35352,N_35464);
nand U35538 (N_35538,N_35459,N_35319);
xor U35539 (N_35539,N_35434,N_35477);
nand U35540 (N_35540,N_35493,N_35315);
nor U35541 (N_35541,N_35346,N_35429);
nor U35542 (N_35542,N_35279,N_35415);
nand U35543 (N_35543,N_35255,N_35422);
nor U35544 (N_35544,N_35403,N_35298);
or U35545 (N_35545,N_35430,N_35402);
and U35546 (N_35546,N_35369,N_35448);
xnor U35547 (N_35547,N_35282,N_35489);
or U35548 (N_35548,N_35311,N_35292);
nor U35549 (N_35549,N_35433,N_35337);
xnor U35550 (N_35550,N_35256,N_35494);
nor U35551 (N_35551,N_35293,N_35347);
xor U35552 (N_35552,N_35394,N_35259);
nand U35553 (N_35553,N_35351,N_35388);
nand U35554 (N_35554,N_35252,N_35316);
and U35555 (N_35555,N_35302,N_35476);
xor U35556 (N_35556,N_35449,N_35405);
nand U35557 (N_35557,N_35446,N_35286);
xnor U35558 (N_35558,N_35251,N_35416);
or U35559 (N_35559,N_35363,N_35275);
and U35560 (N_35560,N_35305,N_35495);
nand U35561 (N_35561,N_35281,N_35468);
nand U35562 (N_35562,N_35357,N_35397);
nand U35563 (N_35563,N_35350,N_35480);
nand U35564 (N_35564,N_35469,N_35349);
and U35565 (N_35565,N_35483,N_35334);
nand U35566 (N_35566,N_35271,N_35265);
xnor U35567 (N_35567,N_35412,N_35370);
and U35568 (N_35568,N_35408,N_35367);
or U35569 (N_35569,N_35312,N_35424);
and U35570 (N_35570,N_35274,N_35294);
xor U35571 (N_35571,N_35365,N_35389);
nor U35572 (N_35572,N_35257,N_35348);
nand U35573 (N_35573,N_35497,N_35486);
or U35574 (N_35574,N_35462,N_35301);
or U35575 (N_35575,N_35327,N_35360);
nor U35576 (N_35576,N_35427,N_35396);
nor U35577 (N_35577,N_35407,N_35278);
xnor U35578 (N_35578,N_35341,N_35436);
nand U35579 (N_35579,N_35332,N_35390);
nand U35580 (N_35580,N_35435,N_35313);
nor U35581 (N_35581,N_35465,N_35300);
or U35582 (N_35582,N_35290,N_35284);
nand U35583 (N_35583,N_35457,N_35304);
or U35584 (N_35584,N_35374,N_35393);
and U35585 (N_35585,N_35303,N_35382);
or U35586 (N_35586,N_35428,N_35442);
and U35587 (N_35587,N_35320,N_35336);
nand U35588 (N_35588,N_35340,N_35368);
nor U35589 (N_35589,N_35353,N_35420);
nor U35590 (N_35590,N_35383,N_35333);
or U35591 (N_35591,N_35443,N_35386);
xnor U35592 (N_35592,N_35467,N_35470);
xor U35593 (N_35593,N_35440,N_35287);
and U35594 (N_35594,N_35291,N_35487);
xor U35595 (N_35595,N_35395,N_35318);
or U35596 (N_35596,N_35324,N_35344);
nor U35597 (N_35597,N_35414,N_35454);
and U35598 (N_35598,N_35250,N_35458);
nand U35599 (N_35599,N_35455,N_35441);
xor U35600 (N_35600,N_35372,N_35445);
nand U35601 (N_35601,N_35314,N_35410);
and U35602 (N_35602,N_35432,N_35447);
nor U35603 (N_35603,N_35361,N_35253);
nand U35604 (N_35604,N_35453,N_35426);
nor U35605 (N_35605,N_35277,N_35262);
xor U35606 (N_35606,N_35322,N_35499);
or U35607 (N_35607,N_35481,N_35417);
nor U35608 (N_35608,N_35456,N_35409);
or U35609 (N_35609,N_35451,N_35425);
or U35610 (N_35610,N_35364,N_35492);
and U35611 (N_35611,N_35385,N_35335);
and U35612 (N_35612,N_35307,N_35308);
nand U35613 (N_35613,N_35359,N_35461);
or U35614 (N_35614,N_35371,N_35329);
nand U35615 (N_35615,N_35419,N_35474);
or U35616 (N_35616,N_35354,N_35296);
xnor U35617 (N_35617,N_35473,N_35380);
or U35618 (N_35618,N_35325,N_35466);
xnor U35619 (N_35619,N_35479,N_35309);
or U35620 (N_35620,N_35289,N_35358);
and U35621 (N_35621,N_35399,N_35328);
and U35622 (N_35622,N_35381,N_35285);
and U35623 (N_35623,N_35261,N_35295);
or U35624 (N_35624,N_35384,N_35366);
nor U35625 (N_35625,N_35259,N_35456);
xnor U35626 (N_35626,N_35321,N_35462);
nor U35627 (N_35627,N_35453,N_35339);
or U35628 (N_35628,N_35280,N_35346);
nand U35629 (N_35629,N_35473,N_35365);
xor U35630 (N_35630,N_35468,N_35276);
nand U35631 (N_35631,N_35320,N_35283);
xor U35632 (N_35632,N_35289,N_35404);
nand U35633 (N_35633,N_35278,N_35430);
xor U35634 (N_35634,N_35351,N_35398);
and U35635 (N_35635,N_35357,N_35367);
or U35636 (N_35636,N_35307,N_35371);
nand U35637 (N_35637,N_35315,N_35481);
nor U35638 (N_35638,N_35421,N_35459);
nand U35639 (N_35639,N_35310,N_35351);
nand U35640 (N_35640,N_35436,N_35355);
and U35641 (N_35641,N_35483,N_35434);
nand U35642 (N_35642,N_35494,N_35288);
nand U35643 (N_35643,N_35276,N_35328);
xor U35644 (N_35644,N_35499,N_35264);
nor U35645 (N_35645,N_35398,N_35278);
or U35646 (N_35646,N_35435,N_35328);
nand U35647 (N_35647,N_35390,N_35297);
and U35648 (N_35648,N_35337,N_35293);
xnor U35649 (N_35649,N_35470,N_35323);
nand U35650 (N_35650,N_35458,N_35373);
and U35651 (N_35651,N_35403,N_35397);
and U35652 (N_35652,N_35436,N_35332);
nor U35653 (N_35653,N_35363,N_35312);
xnor U35654 (N_35654,N_35436,N_35300);
nor U35655 (N_35655,N_35362,N_35373);
nand U35656 (N_35656,N_35258,N_35359);
xor U35657 (N_35657,N_35430,N_35424);
nand U35658 (N_35658,N_35498,N_35316);
or U35659 (N_35659,N_35252,N_35496);
nand U35660 (N_35660,N_35266,N_35355);
and U35661 (N_35661,N_35386,N_35395);
or U35662 (N_35662,N_35348,N_35400);
xor U35663 (N_35663,N_35420,N_35463);
nor U35664 (N_35664,N_35489,N_35498);
nor U35665 (N_35665,N_35393,N_35253);
xnor U35666 (N_35666,N_35419,N_35270);
nor U35667 (N_35667,N_35482,N_35444);
nor U35668 (N_35668,N_35438,N_35363);
or U35669 (N_35669,N_35276,N_35465);
xnor U35670 (N_35670,N_35496,N_35336);
xnor U35671 (N_35671,N_35381,N_35272);
nor U35672 (N_35672,N_35474,N_35445);
nand U35673 (N_35673,N_35444,N_35497);
nor U35674 (N_35674,N_35358,N_35320);
or U35675 (N_35675,N_35338,N_35358);
nor U35676 (N_35676,N_35378,N_35382);
or U35677 (N_35677,N_35321,N_35391);
nor U35678 (N_35678,N_35292,N_35455);
nor U35679 (N_35679,N_35460,N_35311);
xnor U35680 (N_35680,N_35296,N_35480);
and U35681 (N_35681,N_35397,N_35376);
xnor U35682 (N_35682,N_35470,N_35430);
and U35683 (N_35683,N_35305,N_35341);
and U35684 (N_35684,N_35298,N_35290);
xnor U35685 (N_35685,N_35386,N_35352);
nor U35686 (N_35686,N_35422,N_35437);
and U35687 (N_35687,N_35355,N_35462);
or U35688 (N_35688,N_35348,N_35443);
and U35689 (N_35689,N_35271,N_35365);
nand U35690 (N_35690,N_35261,N_35496);
nand U35691 (N_35691,N_35266,N_35251);
nand U35692 (N_35692,N_35364,N_35453);
nand U35693 (N_35693,N_35413,N_35451);
or U35694 (N_35694,N_35381,N_35389);
nor U35695 (N_35695,N_35424,N_35290);
or U35696 (N_35696,N_35395,N_35376);
nor U35697 (N_35697,N_35285,N_35488);
nand U35698 (N_35698,N_35324,N_35414);
nor U35699 (N_35699,N_35467,N_35358);
and U35700 (N_35700,N_35463,N_35298);
or U35701 (N_35701,N_35444,N_35339);
nand U35702 (N_35702,N_35287,N_35312);
nor U35703 (N_35703,N_35496,N_35446);
and U35704 (N_35704,N_35375,N_35341);
or U35705 (N_35705,N_35284,N_35452);
and U35706 (N_35706,N_35350,N_35309);
nor U35707 (N_35707,N_35336,N_35254);
or U35708 (N_35708,N_35271,N_35410);
xnor U35709 (N_35709,N_35421,N_35305);
and U35710 (N_35710,N_35259,N_35403);
xor U35711 (N_35711,N_35263,N_35391);
xnor U35712 (N_35712,N_35337,N_35437);
xnor U35713 (N_35713,N_35343,N_35346);
xor U35714 (N_35714,N_35344,N_35447);
or U35715 (N_35715,N_35418,N_35334);
nor U35716 (N_35716,N_35319,N_35295);
or U35717 (N_35717,N_35424,N_35415);
or U35718 (N_35718,N_35269,N_35457);
xnor U35719 (N_35719,N_35445,N_35333);
and U35720 (N_35720,N_35426,N_35444);
nand U35721 (N_35721,N_35470,N_35347);
nand U35722 (N_35722,N_35379,N_35317);
xor U35723 (N_35723,N_35368,N_35471);
nand U35724 (N_35724,N_35359,N_35442);
nand U35725 (N_35725,N_35253,N_35354);
or U35726 (N_35726,N_35434,N_35491);
xnor U35727 (N_35727,N_35457,N_35498);
xor U35728 (N_35728,N_35445,N_35331);
nor U35729 (N_35729,N_35485,N_35404);
nor U35730 (N_35730,N_35319,N_35485);
nor U35731 (N_35731,N_35461,N_35491);
nor U35732 (N_35732,N_35482,N_35276);
or U35733 (N_35733,N_35306,N_35311);
and U35734 (N_35734,N_35412,N_35343);
and U35735 (N_35735,N_35306,N_35478);
xor U35736 (N_35736,N_35274,N_35275);
nand U35737 (N_35737,N_35485,N_35497);
or U35738 (N_35738,N_35257,N_35288);
xnor U35739 (N_35739,N_35323,N_35287);
xor U35740 (N_35740,N_35467,N_35320);
nand U35741 (N_35741,N_35311,N_35477);
nand U35742 (N_35742,N_35337,N_35384);
or U35743 (N_35743,N_35480,N_35407);
nor U35744 (N_35744,N_35479,N_35368);
nand U35745 (N_35745,N_35320,N_35384);
xor U35746 (N_35746,N_35381,N_35447);
nor U35747 (N_35747,N_35492,N_35304);
nor U35748 (N_35748,N_35351,N_35475);
and U35749 (N_35749,N_35341,N_35361);
xor U35750 (N_35750,N_35670,N_35671);
and U35751 (N_35751,N_35654,N_35558);
or U35752 (N_35752,N_35608,N_35629);
nand U35753 (N_35753,N_35655,N_35618);
and U35754 (N_35754,N_35692,N_35650);
xnor U35755 (N_35755,N_35602,N_35640);
or U35756 (N_35756,N_35611,N_35663);
nand U35757 (N_35757,N_35567,N_35570);
nor U35758 (N_35758,N_35565,N_35635);
nor U35759 (N_35759,N_35623,N_35519);
nor U35760 (N_35760,N_35507,N_35702);
nand U35761 (N_35761,N_35660,N_35545);
nand U35762 (N_35762,N_35676,N_35564);
or U35763 (N_35763,N_35693,N_35546);
nor U35764 (N_35764,N_35607,N_35636);
nand U35765 (N_35765,N_35733,N_35522);
and U35766 (N_35766,N_35684,N_35529);
or U35767 (N_35767,N_35613,N_35728);
and U35768 (N_35768,N_35646,N_35617);
xnor U35769 (N_35769,N_35738,N_35606);
and U35770 (N_35770,N_35632,N_35593);
nor U35771 (N_35771,N_35615,N_35642);
or U35772 (N_35772,N_35595,N_35683);
xor U35773 (N_35773,N_35509,N_35644);
xor U35774 (N_35774,N_35737,N_35614);
or U35775 (N_35775,N_35555,N_35708);
and U35776 (N_35776,N_35572,N_35552);
nor U35777 (N_35777,N_35664,N_35600);
xnor U35778 (N_35778,N_35645,N_35543);
nor U35779 (N_35779,N_35575,N_35707);
xnor U35780 (N_35780,N_35513,N_35719);
and U35781 (N_35781,N_35682,N_35704);
nand U35782 (N_35782,N_35537,N_35511);
or U35783 (N_35783,N_35594,N_35508);
or U35784 (N_35784,N_35582,N_35727);
nor U35785 (N_35785,N_35599,N_35667);
nand U35786 (N_35786,N_35621,N_35603);
nand U35787 (N_35787,N_35514,N_35518);
nor U35788 (N_35788,N_35515,N_35540);
or U35789 (N_35789,N_35605,N_35542);
nor U35790 (N_35790,N_35681,N_35528);
nor U35791 (N_35791,N_35643,N_35685);
nand U35792 (N_35792,N_35633,N_35557);
xnor U35793 (N_35793,N_35731,N_35745);
nand U35794 (N_35794,N_35674,N_35724);
or U35795 (N_35795,N_35679,N_35740);
and U35796 (N_35796,N_35686,N_35657);
nand U35797 (N_35797,N_35656,N_35673);
nor U35798 (N_35798,N_35627,N_35585);
xnor U35799 (N_35799,N_35604,N_35649);
or U35800 (N_35800,N_35701,N_35639);
xor U35801 (N_35801,N_35678,N_35736);
xnor U35802 (N_35802,N_35730,N_35566);
xor U35803 (N_35803,N_35574,N_35717);
xnor U35804 (N_35804,N_35510,N_35732);
xnor U35805 (N_35805,N_35699,N_35536);
nand U35806 (N_35806,N_35535,N_35666);
and U35807 (N_35807,N_35662,N_35541);
and U35808 (N_35808,N_35722,N_35501);
and U35809 (N_35809,N_35652,N_35549);
nor U35810 (N_35810,N_35577,N_35583);
and U35811 (N_35811,N_35601,N_35700);
xor U35812 (N_35812,N_35573,N_35556);
or U35813 (N_35813,N_35742,N_35616);
or U35814 (N_35814,N_35533,N_35721);
nor U35815 (N_35815,N_35591,N_35677);
or U35816 (N_35816,N_35581,N_35739);
nor U35817 (N_35817,N_35539,N_35622);
nor U35818 (N_35818,N_35697,N_35687);
xor U35819 (N_35819,N_35505,N_35610);
nor U35820 (N_35820,N_35688,N_35560);
and U35821 (N_35821,N_35587,N_35512);
or U35822 (N_35822,N_35626,N_35590);
nand U35823 (N_35823,N_35553,N_35744);
xor U35824 (N_35824,N_35711,N_35520);
nand U35825 (N_35825,N_35516,N_35709);
nand U35826 (N_35826,N_35638,N_35524);
xor U35827 (N_35827,N_35713,N_35694);
or U35828 (N_35828,N_35706,N_35571);
and U35829 (N_35829,N_35538,N_35691);
or U35830 (N_35830,N_35741,N_35658);
xor U35831 (N_35831,N_35672,N_35743);
nor U35832 (N_35832,N_35548,N_35689);
or U35833 (N_35833,N_35661,N_35716);
nor U35834 (N_35834,N_35747,N_35503);
and U35835 (N_35835,N_35550,N_35668);
and U35836 (N_35836,N_35637,N_35584);
nor U35837 (N_35837,N_35559,N_35597);
xnor U35838 (N_35838,N_35675,N_35589);
or U35839 (N_35839,N_35586,N_35576);
nor U35840 (N_35840,N_35554,N_35746);
and U35841 (N_35841,N_35718,N_35517);
and U35842 (N_35842,N_35547,N_35705);
and U35843 (N_35843,N_35562,N_35612);
nand U35844 (N_35844,N_35530,N_35648);
xnor U35845 (N_35845,N_35710,N_35609);
nor U35846 (N_35846,N_35561,N_35715);
nor U35847 (N_35847,N_35659,N_35544);
xnor U35848 (N_35848,N_35653,N_35620);
nand U35849 (N_35849,N_35563,N_35748);
and U35850 (N_35850,N_35631,N_35502);
xor U35851 (N_35851,N_35569,N_35624);
nand U35852 (N_35852,N_35647,N_35696);
nor U35853 (N_35853,N_35641,N_35531);
nor U35854 (N_35854,N_35527,N_35729);
or U35855 (N_35855,N_35588,N_35506);
nand U35856 (N_35856,N_35534,N_35714);
nand U35857 (N_35857,N_35726,N_35598);
nor U35858 (N_35858,N_35625,N_35532);
xor U35859 (N_35859,N_35500,N_35579);
nor U35860 (N_35860,N_35525,N_35712);
or U35861 (N_35861,N_35735,N_35680);
or U35862 (N_35862,N_35665,N_35734);
or U35863 (N_35863,N_35749,N_35619);
nand U35864 (N_35864,N_35703,N_35723);
xnor U35865 (N_35865,N_35630,N_35698);
and U35866 (N_35866,N_35596,N_35669);
nand U35867 (N_35867,N_35720,N_35695);
xnor U35868 (N_35868,N_35551,N_35526);
nor U35869 (N_35869,N_35521,N_35628);
nor U35870 (N_35870,N_35690,N_35568);
nand U35871 (N_35871,N_35592,N_35504);
nand U35872 (N_35872,N_35725,N_35634);
or U35873 (N_35873,N_35523,N_35580);
nor U35874 (N_35874,N_35651,N_35578);
nand U35875 (N_35875,N_35713,N_35646);
xnor U35876 (N_35876,N_35630,N_35562);
or U35877 (N_35877,N_35672,N_35706);
nor U35878 (N_35878,N_35542,N_35675);
nand U35879 (N_35879,N_35701,N_35529);
and U35880 (N_35880,N_35626,N_35676);
nor U35881 (N_35881,N_35579,N_35706);
nand U35882 (N_35882,N_35710,N_35582);
or U35883 (N_35883,N_35668,N_35735);
nor U35884 (N_35884,N_35593,N_35711);
or U35885 (N_35885,N_35542,N_35621);
or U35886 (N_35886,N_35574,N_35563);
nor U35887 (N_35887,N_35531,N_35689);
nor U35888 (N_35888,N_35577,N_35645);
xnor U35889 (N_35889,N_35696,N_35651);
xnor U35890 (N_35890,N_35597,N_35695);
and U35891 (N_35891,N_35604,N_35602);
nand U35892 (N_35892,N_35550,N_35514);
nor U35893 (N_35893,N_35650,N_35634);
or U35894 (N_35894,N_35708,N_35528);
or U35895 (N_35895,N_35701,N_35628);
xor U35896 (N_35896,N_35679,N_35630);
xor U35897 (N_35897,N_35741,N_35659);
xnor U35898 (N_35898,N_35684,N_35527);
or U35899 (N_35899,N_35651,N_35535);
xor U35900 (N_35900,N_35528,N_35581);
xnor U35901 (N_35901,N_35634,N_35544);
and U35902 (N_35902,N_35618,N_35600);
xnor U35903 (N_35903,N_35711,N_35654);
nor U35904 (N_35904,N_35632,N_35653);
or U35905 (N_35905,N_35711,N_35736);
xnor U35906 (N_35906,N_35686,N_35574);
nand U35907 (N_35907,N_35552,N_35568);
or U35908 (N_35908,N_35612,N_35602);
or U35909 (N_35909,N_35747,N_35570);
nor U35910 (N_35910,N_35561,N_35509);
or U35911 (N_35911,N_35713,N_35613);
nor U35912 (N_35912,N_35503,N_35728);
or U35913 (N_35913,N_35711,N_35535);
nor U35914 (N_35914,N_35580,N_35720);
nand U35915 (N_35915,N_35675,N_35725);
xnor U35916 (N_35916,N_35558,N_35729);
xnor U35917 (N_35917,N_35610,N_35652);
and U35918 (N_35918,N_35651,N_35640);
nor U35919 (N_35919,N_35706,N_35626);
xnor U35920 (N_35920,N_35560,N_35600);
nand U35921 (N_35921,N_35553,N_35629);
xnor U35922 (N_35922,N_35687,N_35675);
xor U35923 (N_35923,N_35550,N_35568);
and U35924 (N_35924,N_35685,N_35642);
and U35925 (N_35925,N_35688,N_35700);
nand U35926 (N_35926,N_35644,N_35551);
and U35927 (N_35927,N_35564,N_35735);
nand U35928 (N_35928,N_35623,N_35612);
nor U35929 (N_35929,N_35652,N_35683);
nand U35930 (N_35930,N_35593,N_35545);
or U35931 (N_35931,N_35607,N_35722);
xor U35932 (N_35932,N_35681,N_35621);
nor U35933 (N_35933,N_35642,N_35580);
nor U35934 (N_35934,N_35523,N_35558);
and U35935 (N_35935,N_35504,N_35613);
and U35936 (N_35936,N_35505,N_35643);
or U35937 (N_35937,N_35611,N_35590);
or U35938 (N_35938,N_35502,N_35702);
xnor U35939 (N_35939,N_35626,N_35605);
or U35940 (N_35940,N_35673,N_35643);
nand U35941 (N_35941,N_35664,N_35606);
xor U35942 (N_35942,N_35598,N_35694);
xnor U35943 (N_35943,N_35541,N_35661);
or U35944 (N_35944,N_35575,N_35721);
xnor U35945 (N_35945,N_35583,N_35568);
nand U35946 (N_35946,N_35515,N_35576);
xor U35947 (N_35947,N_35691,N_35661);
nand U35948 (N_35948,N_35656,N_35603);
nand U35949 (N_35949,N_35577,N_35629);
or U35950 (N_35950,N_35517,N_35735);
xnor U35951 (N_35951,N_35670,N_35524);
nand U35952 (N_35952,N_35600,N_35647);
xor U35953 (N_35953,N_35684,N_35608);
xnor U35954 (N_35954,N_35743,N_35706);
nor U35955 (N_35955,N_35535,N_35613);
and U35956 (N_35956,N_35735,N_35585);
or U35957 (N_35957,N_35643,N_35545);
nor U35958 (N_35958,N_35523,N_35539);
and U35959 (N_35959,N_35663,N_35607);
nor U35960 (N_35960,N_35741,N_35576);
and U35961 (N_35961,N_35745,N_35567);
nand U35962 (N_35962,N_35588,N_35746);
nor U35963 (N_35963,N_35555,N_35688);
or U35964 (N_35964,N_35589,N_35646);
and U35965 (N_35965,N_35667,N_35581);
or U35966 (N_35966,N_35644,N_35549);
nor U35967 (N_35967,N_35741,N_35657);
nand U35968 (N_35968,N_35574,N_35516);
xnor U35969 (N_35969,N_35597,N_35539);
or U35970 (N_35970,N_35740,N_35678);
or U35971 (N_35971,N_35554,N_35594);
nor U35972 (N_35972,N_35676,N_35506);
nand U35973 (N_35973,N_35663,N_35503);
xnor U35974 (N_35974,N_35588,N_35744);
xnor U35975 (N_35975,N_35500,N_35671);
nor U35976 (N_35976,N_35520,N_35557);
xor U35977 (N_35977,N_35696,N_35552);
xor U35978 (N_35978,N_35538,N_35660);
and U35979 (N_35979,N_35545,N_35623);
xnor U35980 (N_35980,N_35588,N_35655);
and U35981 (N_35981,N_35553,N_35595);
xnor U35982 (N_35982,N_35746,N_35741);
nor U35983 (N_35983,N_35525,N_35724);
and U35984 (N_35984,N_35742,N_35697);
and U35985 (N_35985,N_35667,N_35547);
xor U35986 (N_35986,N_35700,N_35665);
nand U35987 (N_35987,N_35584,N_35563);
nor U35988 (N_35988,N_35681,N_35744);
nor U35989 (N_35989,N_35729,N_35714);
nor U35990 (N_35990,N_35538,N_35627);
and U35991 (N_35991,N_35571,N_35597);
nor U35992 (N_35992,N_35733,N_35511);
nand U35993 (N_35993,N_35545,N_35640);
nor U35994 (N_35994,N_35601,N_35538);
and U35995 (N_35995,N_35532,N_35696);
and U35996 (N_35996,N_35560,N_35734);
or U35997 (N_35997,N_35520,N_35532);
or U35998 (N_35998,N_35725,N_35633);
and U35999 (N_35999,N_35566,N_35516);
and U36000 (N_36000,N_35783,N_35890);
nand U36001 (N_36001,N_35996,N_35787);
nor U36002 (N_36002,N_35856,N_35779);
nor U36003 (N_36003,N_35894,N_35920);
xor U36004 (N_36004,N_35978,N_35767);
nor U36005 (N_36005,N_35919,N_35834);
and U36006 (N_36006,N_35992,N_35989);
and U36007 (N_36007,N_35949,N_35950);
and U36008 (N_36008,N_35980,N_35968);
or U36009 (N_36009,N_35991,N_35903);
or U36010 (N_36010,N_35922,N_35795);
nor U36011 (N_36011,N_35981,N_35803);
and U36012 (N_36012,N_35936,N_35877);
or U36013 (N_36013,N_35998,N_35824);
nand U36014 (N_36014,N_35826,N_35857);
nand U36015 (N_36015,N_35780,N_35768);
or U36016 (N_36016,N_35935,N_35751);
xnor U36017 (N_36017,N_35994,N_35771);
nor U36018 (N_36018,N_35808,N_35961);
nand U36019 (N_36019,N_35820,N_35909);
or U36020 (N_36020,N_35882,N_35831);
xnor U36021 (N_36021,N_35964,N_35871);
and U36022 (N_36022,N_35902,N_35911);
or U36023 (N_36023,N_35764,N_35847);
or U36024 (N_36024,N_35899,N_35900);
nor U36025 (N_36025,N_35770,N_35910);
xor U36026 (N_36026,N_35957,N_35931);
or U36027 (N_36027,N_35946,N_35889);
or U36028 (N_36028,N_35789,N_35801);
xor U36029 (N_36029,N_35757,N_35942);
and U36030 (N_36030,N_35867,N_35807);
nor U36031 (N_36031,N_35913,N_35796);
and U36032 (N_36032,N_35754,N_35761);
nand U36033 (N_36033,N_35921,N_35775);
and U36034 (N_36034,N_35883,N_35842);
nor U36035 (N_36035,N_35958,N_35849);
or U36036 (N_36036,N_35860,N_35925);
nor U36037 (N_36037,N_35893,N_35858);
xor U36038 (N_36038,N_35941,N_35865);
nand U36039 (N_36039,N_35854,N_35892);
nand U36040 (N_36040,N_35974,N_35818);
or U36041 (N_36041,N_35830,N_35792);
and U36042 (N_36042,N_35916,N_35896);
nor U36043 (N_36043,N_35859,N_35836);
and U36044 (N_36044,N_35945,N_35969);
nand U36045 (N_36045,N_35765,N_35844);
nand U36046 (N_36046,N_35986,N_35960);
and U36047 (N_36047,N_35993,N_35752);
nand U36048 (N_36048,N_35837,N_35846);
xor U36049 (N_36049,N_35982,N_35750);
nor U36050 (N_36050,N_35791,N_35979);
xor U36051 (N_36051,N_35813,N_35997);
or U36052 (N_36052,N_35891,N_35923);
and U36053 (N_36053,N_35901,N_35955);
xnor U36054 (N_36054,N_35845,N_35774);
and U36055 (N_36055,N_35804,N_35778);
xor U36056 (N_36056,N_35855,N_35797);
or U36057 (N_36057,N_35755,N_35758);
and U36058 (N_36058,N_35806,N_35759);
or U36059 (N_36059,N_35937,N_35832);
and U36060 (N_36060,N_35905,N_35835);
nor U36061 (N_36061,N_35785,N_35784);
xnor U36062 (N_36062,N_35888,N_35762);
nand U36063 (N_36063,N_35790,N_35753);
and U36064 (N_36064,N_35912,N_35776);
xnor U36065 (N_36065,N_35819,N_35948);
and U36066 (N_36066,N_35904,N_35929);
or U36067 (N_36067,N_35868,N_35821);
nor U36068 (N_36068,N_35988,N_35959);
and U36069 (N_36069,N_35930,N_35763);
and U36070 (N_36070,N_35866,N_35777);
and U36071 (N_36071,N_35947,N_35881);
nor U36072 (N_36072,N_35794,N_35863);
nor U36073 (N_36073,N_35862,N_35814);
or U36074 (N_36074,N_35873,N_35786);
nand U36075 (N_36075,N_35861,N_35875);
xnor U36076 (N_36076,N_35938,N_35906);
nor U36077 (N_36077,N_35869,N_35811);
nand U36078 (N_36078,N_35972,N_35932);
xnor U36079 (N_36079,N_35975,N_35876);
nor U36080 (N_36080,N_35766,N_35990);
or U36081 (N_36081,N_35833,N_35885);
xnor U36082 (N_36082,N_35943,N_35887);
nand U36083 (N_36083,N_35977,N_35933);
and U36084 (N_36084,N_35956,N_35984);
nor U36085 (N_36085,N_35828,N_35924);
and U36086 (N_36086,N_35850,N_35973);
nand U36087 (N_36087,N_35934,N_35843);
nand U36088 (N_36088,N_35822,N_35927);
xor U36089 (N_36089,N_35772,N_35962);
xnor U36090 (N_36090,N_35769,N_35798);
and U36091 (N_36091,N_35800,N_35878);
xnor U36092 (N_36092,N_35940,N_35983);
xor U36093 (N_36093,N_35985,N_35838);
and U36094 (N_36094,N_35952,N_35817);
or U36095 (N_36095,N_35886,N_35987);
nand U36096 (N_36096,N_35966,N_35965);
or U36097 (N_36097,N_35970,N_35884);
and U36098 (N_36098,N_35971,N_35812);
nand U36099 (N_36099,N_35852,N_35999);
or U36100 (N_36100,N_35823,N_35793);
nor U36101 (N_36101,N_35809,N_35756);
nand U36102 (N_36102,N_35760,N_35782);
xnor U36103 (N_36103,N_35781,N_35827);
or U36104 (N_36104,N_35895,N_35880);
nand U36105 (N_36105,N_35918,N_35951);
and U36106 (N_36106,N_35825,N_35907);
nor U36107 (N_36107,N_35815,N_35839);
xnor U36108 (N_36108,N_35976,N_35879);
and U36109 (N_36109,N_35851,N_35908);
or U36110 (N_36110,N_35953,N_35874);
nor U36111 (N_36111,N_35840,N_35788);
and U36112 (N_36112,N_35944,N_35954);
nand U36113 (N_36113,N_35995,N_35915);
and U36114 (N_36114,N_35914,N_35928);
nor U36115 (N_36115,N_35939,N_35897);
and U36116 (N_36116,N_35805,N_35967);
nand U36117 (N_36117,N_35917,N_35799);
nand U36118 (N_36118,N_35802,N_35872);
nand U36119 (N_36119,N_35853,N_35926);
nand U36120 (N_36120,N_35816,N_35870);
nor U36121 (N_36121,N_35841,N_35829);
or U36122 (N_36122,N_35898,N_35810);
nand U36123 (N_36123,N_35963,N_35864);
nor U36124 (N_36124,N_35773,N_35848);
or U36125 (N_36125,N_35829,N_35771);
nand U36126 (N_36126,N_35850,N_35949);
nor U36127 (N_36127,N_35892,N_35919);
and U36128 (N_36128,N_35838,N_35821);
or U36129 (N_36129,N_35918,N_35994);
nand U36130 (N_36130,N_35796,N_35819);
nor U36131 (N_36131,N_35852,N_35849);
xor U36132 (N_36132,N_35956,N_35851);
and U36133 (N_36133,N_35815,N_35843);
nor U36134 (N_36134,N_35943,N_35945);
and U36135 (N_36135,N_35989,N_35998);
xor U36136 (N_36136,N_35955,N_35908);
nor U36137 (N_36137,N_35949,N_35772);
nor U36138 (N_36138,N_35769,N_35860);
or U36139 (N_36139,N_35930,N_35990);
nand U36140 (N_36140,N_35780,N_35943);
or U36141 (N_36141,N_35888,N_35843);
nor U36142 (N_36142,N_35935,N_35970);
and U36143 (N_36143,N_35770,N_35832);
nand U36144 (N_36144,N_35819,N_35788);
nor U36145 (N_36145,N_35953,N_35890);
and U36146 (N_36146,N_35992,N_35786);
nor U36147 (N_36147,N_35973,N_35765);
or U36148 (N_36148,N_35792,N_35839);
xor U36149 (N_36149,N_35913,N_35818);
and U36150 (N_36150,N_35916,N_35820);
nand U36151 (N_36151,N_35846,N_35940);
or U36152 (N_36152,N_35917,N_35992);
nand U36153 (N_36153,N_35853,N_35934);
and U36154 (N_36154,N_35922,N_35821);
nand U36155 (N_36155,N_35933,N_35982);
or U36156 (N_36156,N_35810,N_35983);
and U36157 (N_36157,N_35900,N_35973);
nand U36158 (N_36158,N_35786,N_35902);
nand U36159 (N_36159,N_35926,N_35842);
nor U36160 (N_36160,N_35781,N_35939);
or U36161 (N_36161,N_35779,N_35959);
xor U36162 (N_36162,N_35997,N_35951);
or U36163 (N_36163,N_35769,N_35873);
or U36164 (N_36164,N_35886,N_35890);
xor U36165 (N_36165,N_35931,N_35853);
xor U36166 (N_36166,N_35772,N_35989);
nor U36167 (N_36167,N_35868,N_35785);
and U36168 (N_36168,N_35802,N_35853);
xnor U36169 (N_36169,N_35813,N_35815);
xor U36170 (N_36170,N_35853,N_35764);
xnor U36171 (N_36171,N_35938,N_35881);
xor U36172 (N_36172,N_35969,N_35938);
nand U36173 (N_36173,N_35757,N_35861);
xor U36174 (N_36174,N_35969,N_35792);
and U36175 (N_36175,N_35804,N_35982);
nand U36176 (N_36176,N_35910,N_35949);
and U36177 (N_36177,N_35806,N_35941);
xnor U36178 (N_36178,N_35867,N_35999);
and U36179 (N_36179,N_35851,N_35839);
or U36180 (N_36180,N_35997,N_35935);
nor U36181 (N_36181,N_35998,N_35758);
xor U36182 (N_36182,N_35867,N_35939);
and U36183 (N_36183,N_35807,N_35816);
or U36184 (N_36184,N_35811,N_35865);
or U36185 (N_36185,N_35935,N_35791);
or U36186 (N_36186,N_35780,N_35832);
or U36187 (N_36187,N_35809,N_35799);
nand U36188 (N_36188,N_35907,N_35783);
xnor U36189 (N_36189,N_35769,N_35790);
and U36190 (N_36190,N_35832,N_35783);
nand U36191 (N_36191,N_35982,N_35841);
nand U36192 (N_36192,N_35946,N_35844);
and U36193 (N_36193,N_35953,N_35948);
nand U36194 (N_36194,N_35974,N_35754);
nor U36195 (N_36195,N_35979,N_35963);
or U36196 (N_36196,N_35788,N_35757);
nand U36197 (N_36197,N_35874,N_35847);
or U36198 (N_36198,N_35960,N_35975);
nand U36199 (N_36199,N_35818,N_35875);
xnor U36200 (N_36200,N_35851,N_35762);
or U36201 (N_36201,N_35897,N_35962);
and U36202 (N_36202,N_35975,N_35973);
nor U36203 (N_36203,N_35857,N_35942);
or U36204 (N_36204,N_35835,N_35870);
xnor U36205 (N_36205,N_35765,N_35892);
nand U36206 (N_36206,N_35832,N_35912);
nand U36207 (N_36207,N_35754,N_35887);
or U36208 (N_36208,N_35860,N_35953);
or U36209 (N_36209,N_35774,N_35783);
nand U36210 (N_36210,N_35799,N_35800);
or U36211 (N_36211,N_35784,N_35845);
nand U36212 (N_36212,N_35982,N_35791);
and U36213 (N_36213,N_35959,N_35867);
and U36214 (N_36214,N_35911,N_35996);
nor U36215 (N_36215,N_35928,N_35845);
and U36216 (N_36216,N_35750,N_35915);
xnor U36217 (N_36217,N_35766,N_35826);
or U36218 (N_36218,N_35936,N_35906);
nand U36219 (N_36219,N_35801,N_35935);
nor U36220 (N_36220,N_35798,N_35977);
nand U36221 (N_36221,N_35916,N_35824);
and U36222 (N_36222,N_35892,N_35863);
nand U36223 (N_36223,N_35995,N_35848);
and U36224 (N_36224,N_35842,N_35829);
or U36225 (N_36225,N_35891,N_35765);
or U36226 (N_36226,N_35783,N_35775);
xor U36227 (N_36227,N_35938,N_35878);
nor U36228 (N_36228,N_35999,N_35807);
nor U36229 (N_36229,N_35790,N_35884);
or U36230 (N_36230,N_35929,N_35855);
or U36231 (N_36231,N_35853,N_35795);
nand U36232 (N_36232,N_35852,N_35794);
and U36233 (N_36233,N_35776,N_35780);
xnor U36234 (N_36234,N_35968,N_35977);
xor U36235 (N_36235,N_35771,N_35772);
and U36236 (N_36236,N_35894,N_35913);
and U36237 (N_36237,N_35996,N_35888);
or U36238 (N_36238,N_35844,N_35847);
and U36239 (N_36239,N_35986,N_35818);
nand U36240 (N_36240,N_35830,N_35821);
nand U36241 (N_36241,N_35801,N_35897);
nor U36242 (N_36242,N_35908,N_35972);
and U36243 (N_36243,N_35819,N_35966);
xor U36244 (N_36244,N_35947,N_35836);
nand U36245 (N_36245,N_35800,N_35782);
nor U36246 (N_36246,N_35966,N_35960);
or U36247 (N_36247,N_35956,N_35853);
or U36248 (N_36248,N_35762,N_35969);
or U36249 (N_36249,N_35889,N_35798);
and U36250 (N_36250,N_36020,N_36176);
xor U36251 (N_36251,N_36140,N_36246);
nor U36252 (N_36252,N_36214,N_36074);
or U36253 (N_36253,N_36056,N_36211);
or U36254 (N_36254,N_36148,N_36160);
nor U36255 (N_36255,N_36209,N_36234);
and U36256 (N_36256,N_36231,N_36072);
and U36257 (N_36257,N_36165,N_36185);
nand U36258 (N_36258,N_36193,N_36228);
nand U36259 (N_36259,N_36132,N_36046);
nor U36260 (N_36260,N_36057,N_36110);
or U36261 (N_36261,N_36180,N_36049);
xnor U36262 (N_36262,N_36221,N_36210);
and U36263 (N_36263,N_36219,N_36181);
nor U36264 (N_36264,N_36196,N_36096);
nand U36265 (N_36265,N_36038,N_36127);
or U36266 (N_36266,N_36146,N_36174);
and U36267 (N_36267,N_36183,N_36009);
nand U36268 (N_36268,N_36007,N_36075);
nand U36269 (N_36269,N_36120,N_36041);
nand U36270 (N_36270,N_36103,N_36017);
nor U36271 (N_36271,N_36188,N_36134);
xor U36272 (N_36272,N_36123,N_36192);
xor U36273 (N_36273,N_36131,N_36061);
nor U36274 (N_36274,N_36106,N_36147);
nor U36275 (N_36275,N_36073,N_36144);
xor U36276 (N_36276,N_36208,N_36244);
nand U36277 (N_36277,N_36059,N_36114);
and U36278 (N_36278,N_36032,N_36065);
nand U36279 (N_36279,N_36161,N_36085);
nand U36280 (N_36280,N_36170,N_36093);
and U36281 (N_36281,N_36014,N_36063);
or U36282 (N_36282,N_36159,N_36230);
or U36283 (N_36283,N_36145,N_36095);
nand U36284 (N_36284,N_36068,N_36249);
nand U36285 (N_36285,N_36101,N_36141);
nand U36286 (N_36286,N_36150,N_36153);
or U36287 (N_36287,N_36199,N_36067);
nor U36288 (N_36288,N_36179,N_36198);
xor U36289 (N_36289,N_36235,N_36109);
nor U36290 (N_36290,N_36055,N_36105);
nand U36291 (N_36291,N_36203,N_36173);
or U36292 (N_36292,N_36223,N_36117);
xor U36293 (N_36293,N_36248,N_36039);
or U36294 (N_36294,N_36078,N_36050);
nor U36295 (N_36295,N_36015,N_36030);
nor U36296 (N_36296,N_36058,N_36043);
or U36297 (N_36297,N_36004,N_36119);
or U36298 (N_36298,N_36034,N_36126);
or U36299 (N_36299,N_36191,N_36240);
nand U36300 (N_36300,N_36098,N_36182);
nand U36301 (N_36301,N_36197,N_36066);
and U36302 (N_36302,N_36129,N_36097);
xnor U36303 (N_36303,N_36115,N_36245);
nor U36304 (N_36304,N_36086,N_36128);
nand U36305 (N_36305,N_36216,N_36142);
xor U36306 (N_36306,N_36023,N_36028);
or U36307 (N_36307,N_36125,N_36006);
nand U36308 (N_36308,N_36155,N_36215);
or U36309 (N_36309,N_36163,N_36217);
nor U36310 (N_36310,N_36166,N_36042);
nand U36311 (N_36311,N_36062,N_36243);
or U36312 (N_36312,N_36229,N_36201);
xnor U36313 (N_36313,N_36001,N_36111);
nor U36314 (N_36314,N_36011,N_36033);
nor U36315 (N_36315,N_36175,N_36027);
or U36316 (N_36316,N_36239,N_36130);
and U36317 (N_36317,N_36118,N_36070);
nor U36318 (N_36318,N_36226,N_36082);
nor U36319 (N_36319,N_36051,N_36036);
xor U36320 (N_36320,N_36139,N_36158);
nor U36321 (N_36321,N_36025,N_36047);
and U36322 (N_36322,N_36241,N_36022);
or U36323 (N_36323,N_36026,N_36104);
nor U36324 (N_36324,N_36220,N_36054);
nand U36325 (N_36325,N_36008,N_36045);
nor U36326 (N_36326,N_36189,N_36064);
xnor U36327 (N_36327,N_36187,N_36247);
nand U36328 (N_36328,N_36060,N_36090);
and U36329 (N_36329,N_36152,N_36124);
or U36330 (N_36330,N_36031,N_36081);
nor U36331 (N_36331,N_36102,N_36016);
nand U36332 (N_36332,N_36167,N_36195);
nor U36333 (N_36333,N_36079,N_36169);
xnor U36334 (N_36334,N_36157,N_36136);
nor U36335 (N_36335,N_36164,N_36237);
xnor U36336 (N_36336,N_36162,N_36099);
and U36337 (N_36337,N_36108,N_36044);
nor U36338 (N_36338,N_36092,N_36003);
or U36339 (N_36339,N_36190,N_36071);
xnor U36340 (N_36340,N_36156,N_36048);
nor U36341 (N_36341,N_36083,N_36200);
or U36342 (N_36342,N_36087,N_36094);
xnor U36343 (N_36343,N_36122,N_36089);
nor U36344 (N_36344,N_36168,N_36113);
xor U36345 (N_36345,N_36178,N_36213);
or U36346 (N_36346,N_36035,N_36116);
nor U36347 (N_36347,N_36151,N_36010);
xnor U36348 (N_36348,N_36005,N_36232);
and U36349 (N_36349,N_36091,N_36225);
and U36350 (N_36350,N_36227,N_36002);
and U36351 (N_36351,N_36080,N_36121);
or U36352 (N_36352,N_36204,N_36242);
nor U36353 (N_36353,N_36040,N_36149);
and U36354 (N_36354,N_36236,N_36218);
or U36355 (N_36355,N_36212,N_36222);
xnor U36356 (N_36356,N_36186,N_36112);
nor U36357 (N_36357,N_36224,N_36177);
nor U36358 (N_36358,N_36143,N_36021);
nand U36359 (N_36359,N_36069,N_36024);
xor U36360 (N_36360,N_36100,N_36206);
nand U36361 (N_36361,N_36135,N_36171);
xor U36362 (N_36362,N_36238,N_36172);
or U36363 (N_36363,N_36019,N_36184);
xor U36364 (N_36364,N_36107,N_36154);
nand U36365 (N_36365,N_36013,N_36133);
nor U36366 (N_36366,N_36000,N_36018);
nand U36367 (N_36367,N_36012,N_36207);
and U36368 (N_36368,N_36202,N_36029);
nor U36369 (N_36369,N_36053,N_36088);
and U36370 (N_36370,N_36137,N_36077);
nand U36371 (N_36371,N_36194,N_36037);
or U36372 (N_36372,N_36076,N_36084);
or U36373 (N_36373,N_36205,N_36052);
nand U36374 (N_36374,N_36138,N_36233);
nand U36375 (N_36375,N_36039,N_36068);
and U36376 (N_36376,N_36169,N_36225);
xnor U36377 (N_36377,N_36070,N_36040);
and U36378 (N_36378,N_36050,N_36179);
and U36379 (N_36379,N_36247,N_36057);
nand U36380 (N_36380,N_36156,N_36084);
nand U36381 (N_36381,N_36079,N_36121);
nand U36382 (N_36382,N_36209,N_36141);
and U36383 (N_36383,N_36077,N_36148);
and U36384 (N_36384,N_36162,N_36176);
nand U36385 (N_36385,N_36083,N_36177);
xor U36386 (N_36386,N_36143,N_36249);
xor U36387 (N_36387,N_36000,N_36066);
nor U36388 (N_36388,N_36232,N_36172);
and U36389 (N_36389,N_36164,N_36222);
nor U36390 (N_36390,N_36156,N_36036);
or U36391 (N_36391,N_36236,N_36011);
or U36392 (N_36392,N_36133,N_36148);
and U36393 (N_36393,N_36015,N_36148);
and U36394 (N_36394,N_36227,N_36103);
or U36395 (N_36395,N_36067,N_36059);
and U36396 (N_36396,N_36182,N_36106);
nand U36397 (N_36397,N_36013,N_36101);
and U36398 (N_36398,N_36193,N_36103);
or U36399 (N_36399,N_36148,N_36014);
and U36400 (N_36400,N_36137,N_36219);
xor U36401 (N_36401,N_36065,N_36150);
nand U36402 (N_36402,N_36102,N_36172);
xnor U36403 (N_36403,N_36020,N_36072);
and U36404 (N_36404,N_36023,N_36063);
nand U36405 (N_36405,N_36217,N_36143);
or U36406 (N_36406,N_36042,N_36245);
xor U36407 (N_36407,N_36141,N_36016);
xnor U36408 (N_36408,N_36111,N_36165);
xor U36409 (N_36409,N_36240,N_36014);
nor U36410 (N_36410,N_36045,N_36081);
nand U36411 (N_36411,N_36242,N_36114);
nor U36412 (N_36412,N_36193,N_36210);
nand U36413 (N_36413,N_36230,N_36196);
or U36414 (N_36414,N_36029,N_36034);
and U36415 (N_36415,N_36105,N_36027);
nor U36416 (N_36416,N_36035,N_36037);
xor U36417 (N_36417,N_36233,N_36183);
xor U36418 (N_36418,N_36042,N_36225);
nand U36419 (N_36419,N_36211,N_36204);
nand U36420 (N_36420,N_36112,N_36226);
xor U36421 (N_36421,N_36006,N_36084);
xnor U36422 (N_36422,N_36117,N_36024);
xnor U36423 (N_36423,N_36017,N_36107);
nor U36424 (N_36424,N_36016,N_36171);
nor U36425 (N_36425,N_36193,N_36180);
or U36426 (N_36426,N_36060,N_36121);
nand U36427 (N_36427,N_36231,N_36058);
nand U36428 (N_36428,N_36190,N_36056);
and U36429 (N_36429,N_36185,N_36182);
or U36430 (N_36430,N_36098,N_36117);
nor U36431 (N_36431,N_36001,N_36158);
or U36432 (N_36432,N_36248,N_36213);
xnor U36433 (N_36433,N_36182,N_36227);
xnor U36434 (N_36434,N_36222,N_36189);
xor U36435 (N_36435,N_36119,N_36118);
xor U36436 (N_36436,N_36187,N_36022);
nand U36437 (N_36437,N_36109,N_36119);
or U36438 (N_36438,N_36031,N_36075);
nand U36439 (N_36439,N_36090,N_36144);
and U36440 (N_36440,N_36000,N_36170);
xor U36441 (N_36441,N_36165,N_36016);
nand U36442 (N_36442,N_36067,N_36107);
and U36443 (N_36443,N_36174,N_36226);
or U36444 (N_36444,N_36229,N_36163);
nand U36445 (N_36445,N_36028,N_36081);
and U36446 (N_36446,N_36148,N_36147);
nand U36447 (N_36447,N_36049,N_36046);
nand U36448 (N_36448,N_36097,N_36158);
and U36449 (N_36449,N_36111,N_36039);
nor U36450 (N_36450,N_36236,N_36104);
nor U36451 (N_36451,N_36193,N_36202);
nor U36452 (N_36452,N_36234,N_36118);
or U36453 (N_36453,N_36066,N_36201);
nor U36454 (N_36454,N_36213,N_36073);
xnor U36455 (N_36455,N_36133,N_36038);
nor U36456 (N_36456,N_36073,N_36179);
nand U36457 (N_36457,N_36041,N_36121);
or U36458 (N_36458,N_36114,N_36076);
xor U36459 (N_36459,N_36238,N_36033);
nor U36460 (N_36460,N_36247,N_36188);
xor U36461 (N_36461,N_36138,N_36248);
nor U36462 (N_36462,N_36156,N_36079);
and U36463 (N_36463,N_36057,N_36159);
and U36464 (N_36464,N_36173,N_36232);
nor U36465 (N_36465,N_36062,N_36089);
and U36466 (N_36466,N_36233,N_36008);
nand U36467 (N_36467,N_36088,N_36103);
nor U36468 (N_36468,N_36138,N_36040);
and U36469 (N_36469,N_36070,N_36137);
and U36470 (N_36470,N_36088,N_36117);
nor U36471 (N_36471,N_36101,N_36241);
nor U36472 (N_36472,N_36147,N_36186);
and U36473 (N_36473,N_36049,N_36000);
or U36474 (N_36474,N_36073,N_36074);
xnor U36475 (N_36475,N_36217,N_36140);
nand U36476 (N_36476,N_36049,N_36181);
nand U36477 (N_36477,N_36149,N_36175);
or U36478 (N_36478,N_36020,N_36159);
or U36479 (N_36479,N_36020,N_36076);
nand U36480 (N_36480,N_36200,N_36161);
or U36481 (N_36481,N_36181,N_36171);
and U36482 (N_36482,N_36209,N_36173);
or U36483 (N_36483,N_36090,N_36105);
or U36484 (N_36484,N_36221,N_36243);
or U36485 (N_36485,N_36019,N_36063);
nand U36486 (N_36486,N_36203,N_36064);
nand U36487 (N_36487,N_36003,N_36000);
and U36488 (N_36488,N_36140,N_36115);
and U36489 (N_36489,N_36074,N_36017);
nor U36490 (N_36490,N_36164,N_36190);
nor U36491 (N_36491,N_36091,N_36056);
nor U36492 (N_36492,N_36136,N_36044);
nor U36493 (N_36493,N_36061,N_36090);
and U36494 (N_36494,N_36006,N_36117);
or U36495 (N_36495,N_36055,N_36089);
and U36496 (N_36496,N_36019,N_36102);
nand U36497 (N_36497,N_36004,N_36140);
and U36498 (N_36498,N_36230,N_36064);
nand U36499 (N_36499,N_36118,N_36028);
and U36500 (N_36500,N_36427,N_36489);
xnor U36501 (N_36501,N_36292,N_36287);
and U36502 (N_36502,N_36379,N_36441);
nor U36503 (N_36503,N_36275,N_36337);
nor U36504 (N_36504,N_36381,N_36347);
or U36505 (N_36505,N_36250,N_36415);
or U36506 (N_36506,N_36321,N_36351);
nor U36507 (N_36507,N_36288,N_36326);
nand U36508 (N_36508,N_36327,N_36396);
or U36509 (N_36509,N_36466,N_36333);
xor U36510 (N_36510,N_36318,N_36284);
xnor U36511 (N_36511,N_36316,N_36463);
nor U36512 (N_36512,N_36276,N_36475);
and U36513 (N_36513,N_36440,N_36399);
xnor U36514 (N_36514,N_36290,N_36455);
and U36515 (N_36515,N_36467,N_36401);
nand U36516 (N_36516,N_36421,N_36361);
xor U36517 (N_36517,N_36389,N_36299);
nand U36518 (N_36518,N_36298,N_36331);
and U36519 (N_36519,N_36488,N_36386);
or U36520 (N_36520,N_36446,N_36358);
or U36521 (N_36521,N_36483,N_36498);
and U36522 (N_36522,N_36390,N_36492);
nand U36523 (N_36523,N_36408,N_36414);
nand U36524 (N_36524,N_36302,N_36285);
xor U36525 (N_36525,N_36269,N_36397);
nand U36526 (N_36526,N_36432,N_36480);
nor U36527 (N_36527,N_36260,N_36428);
nand U36528 (N_36528,N_36357,N_36422);
and U36529 (N_36529,N_36476,N_36359);
or U36530 (N_36530,N_36495,N_36309);
and U36531 (N_36531,N_36450,N_36374);
xnor U36532 (N_36532,N_36373,N_36270);
or U36533 (N_36533,N_36315,N_36452);
and U36534 (N_36534,N_36281,N_36457);
nor U36535 (N_36535,N_36312,N_36282);
nor U36536 (N_36536,N_36330,N_36332);
nand U36537 (N_36537,N_36261,N_36255);
nor U36538 (N_36538,N_36461,N_36491);
and U36539 (N_36539,N_36265,N_36295);
xor U36540 (N_36540,N_36482,N_36423);
xnor U36541 (N_36541,N_36437,N_36459);
nand U36542 (N_36542,N_36339,N_36375);
nand U36543 (N_36543,N_36385,N_36348);
or U36544 (N_36544,N_36494,N_36308);
or U36545 (N_36545,N_36490,N_36462);
nor U36546 (N_36546,N_36341,N_36259);
xnor U36547 (N_36547,N_36325,N_36363);
xnor U36548 (N_36548,N_36402,N_36484);
and U36549 (N_36549,N_36460,N_36251);
xor U36550 (N_36550,N_36346,N_36469);
or U36551 (N_36551,N_36294,N_36391);
nor U36552 (N_36552,N_36407,N_36439);
and U36553 (N_36553,N_36479,N_36378);
nand U36554 (N_36554,N_36413,N_36481);
nand U36555 (N_36555,N_36335,N_36384);
xnor U36556 (N_36556,N_36493,N_36354);
and U36557 (N_36557,N_36353,N_36279);
nand U36558 (N_36558,N_36257,N_36278);
xor U36559 (N_36559,N_36436,N_36387);
xnor U36560 (N_36560,N_36438,N_36485);
and U36561 (N_36561,N_36411,N_36487);
and U36562 (N_36562,N_36417,N_36253);
and U36563 (N_36563,N_36430,N_36264);
nor U36564 (N_36564,N_36273,N_36426);
nor U36565 (N_36565,N_36252,N_36256);
xor U36566 (N_36566,N_36405,N_36313);
xnor U36567 (N_36567,N_36317,N_36434);
and U36568 (N_36568,N_36355,N_36496);
or U36569 (N_36569,N_36478,N_36329);
and U36570 (N_36570,N_36274,N_36345);
nand U36571 (N_36571,N_36349,N_36497);
or U36572 (N_36572,N_36409,N_36304);
xnor U36573 (N_36573,N_36424,N_36473);
or U36574 (N_36574,N_36352,N_36388);
nor U36575 (N_36575,N_36293,N_36398);
xnor U36576 (N_36576,N_36362,N_36400);
or U36577 (N_36577,N_36334,N_36322);
or U36578 (N_36578,N_36443,N_36372);
nor U36579 (N_36579,N_36360,N_36271);
or U36580 (N_36580,N_36410,N_36307);
xor U36581 (N_36581,N_36403,N_36395);
or U36582 (N_36582,N_36314,N_36477);
nor U36583 (N_36583,N_36470,N_36420);
nand U36584 (N_36584,N_36419,N_36301);
and U36585 (N_36585,N_36263,N_36254);
xor U36586 (N_36586,N_36464,N_36291);
xor U36587 (N_36587,N_36444,N_36328);
xnor U36588 (N_36588,N_36499,N_36377);
xor U36589 (N_36589,N_36404,N_36297);
nor U36590 (N_36590,N_36350,N_36305);
nand U36591 (N_36591,N_36449,N_36343);
and U36592 (N_36592,N_36296,N_36280);
nor U36593 (N_36593,N_36268,N_36394);
nand U36594 (N_36594,N_36451,N_36453);
xnor U36595 (N_36595,N_36344,N_36340);
and U36596 (N_36596,N_36262,N_36283);
xor U36597 (N_36597,N_36286,N_36433);
or U36598 (N_36598,N_36320,N_36258);
or U36599 (N_36599,N_36310,N_36289);
or U36600 (N_36600,N_36370,N_36267);
nor U36601 (N_36601,N_36468,N_36338);
xor U36602 (N_36602,N_36447,N_36366);
nand U36603 (N_36603,N_36376,N_36323);
nand U36604 (N_36604,N_36474,N_36382);
nor U36605 (N_36605,N_36392,N_36448);
or U36606 (N_36606,N_36367,N_36277);
xor U36607 (N_36607,N_36342,N_36266);
nor U36608 (N_36608,N_36319,N_36458);
xor U36609 (N_36609,N_36435,N_36454);
xnor U36610 (N_36610,N_36486,N_36445);
xor U36611 (N_36611,N_36471,N_36300);
or U36612 (N_36612,N_36472,N_36416);
nor U36613 (N_36613,N_36380,N_36406);
nor U36614 (N_36614,N_36364,N_36365);
or U36615 (N_36615,N_36429,N_36465);
xor U36616 (N_36616,N_36456,N_36442);
or U36617 (N_36617,N_36306,N_36356);
nor U36618 (N_36618,N_36371,N_36412);
or U36619 (N_36619,N_36311,N_36383);
nor U36620 (N_36620,N_36431,N_36425);
or U36621 (N_36621,N_36303,N_36368);
nor U36622 (N_36622,N_36272,N_36418);
or U36623 (N_36623,N_36369,N_36336);
or U36624 (N_36624,N_36393,N_36324);
xor U36625 (N_36625,N_36309,N_36386);
nor U36626 (N_36626,N_36467,N_36279);
and U36627 (N_36627,N_36492,N_36255);
nand U36628 (N_36628,N_36256,N_36281);
and U36629 (N_36629,N_36341,N_36255);
nor U36630 (N_36630,N_36464,N_36328);
nand U36631 (N_36631,N_36418,N_36391);
xnor U36632 (N_36632,N_36497,N_36423);
nand U36633 (N_36633,N_36317,N_36429);
and U36634 (N_36634,N_36265,N_36330);
nand U36635 (N_36635,N_36295,N_36262);
xor U36636 (N_36636,N_36267,N_36409);
and U36637 (N_36637,N_36351,N_36415);
nand U36638 (N_36638,N_36463,N_36470);
or U36639 (N_36639,N_36417,N_36283);
and U36640 (N_36640,N_36392,N_36407);
nor U36641 (N_36641,N_36264,N_36461);
nand U36642 (N_36642,N_36318,N_36407);
nand U36643 (N_36643,N_36442,N_36367);
xnor U36644 (N_36644,N_36409,N_36438);
xor U36645 (N_36645,N_36411,N_36499);
xnor U36646 (N_36646,N_36496,N_36367);
nor U36647 (N_36647,N_36366,N_36348);
nor U36648 (N_36648,N_36330,N_36327);
nand U36649 (N_36649,N_36388,N_36265);
nand U36650 (N_36650,N_36488,N_36250);
nand U36651 (N_36651,N_36352,N_36387);
or U36652 (N_36652,N_36425,N_36293);
or U36653 (N_36653,N_36443,N_36286);
xor U36654 (N_36654,N_36320,N_36280);
or U36655 (N_36655,N_36408,N_36466);
or U36656 (N_36656,N_36357,N_36430);
nor U36657 (N_36657,N_36265,N_36352);
and U36658 (N_36658,N_36390,N_36376);
or U36659 (N_36659,N_36328,N_36353);
xnor U36660 (N_36660,N_36423,N_36463);
and U36661 (N_36661,N_36487,N_36325);
or U36662 (N_36662,N_36313,N_36412);
nor U36663 (N_36663,N_36423,N_36334);
xor U36664 (N_36664,N_36477,N_36320);
nand U36665 (N_36665,N_36265,N_36287);
nor U36666 (N_36666,N_36383,N_36436);
xor U36667 (N_36667,N_36322,N_36369);
nor U36668 (N_36668,N_36329,N_36260);
nor U36669 (N_36669,N_36274,N_36447);
xnor U36670 (N_36670,N_36272,N_36417);
and U36671 (N_36671,N_36265,N_36455);
nor U36672 (N_36672,N_36451,N_36309);
and U36673 (N_36673,N_36254,N_36497);
nand U36674 (N_36674,N_36297,N_36419);
and U36675 (N_36675,N_36462,N_36377);
nor U36676 (N_36676,N_36471,N_36423);
nor U36677 (N_36677,N_36492,N_36391);
nand U36678 (N_36678,N_36265,N_36379);
and U36679 (N_36679,N_36419,N_36455);
nand U36680 (N_36680,N_36255,N_36446);
nand U36681 (N_36681,N_36485,N_36495);
xnor U36682 (N_36682,N_36372,N_36360);
or U36683 (N_36683,N_36323,N_36415);
or U36684 (N_36684,N_36430,N_36436);
xor U36685 (N_36685,N_36462,N_36415);
xnor U36686 (N_36686,N_36443,N_36276);
nand U36687 (N_36687,N_36387,N_36371);
nand U36688 (N_36688,N_36478,N_36252);
or U36689 (N_36689,N_36492,N_36495);
nor U36690 (N_36690,N_36290,N_36399);
and U36691 (N_36691,N_36429,N_36435);
nor U36692 (N_36692,N_36281,N_36418);
xnor U36693 (N_36693,N_36445,N_36267);
nor U36694 (N_36694,N_36281,N_36368);
xnor U36695 (N_36695,N_36410,N_36321);
or U36696 (N_36696,N_36393,N_36390);
nor U36697 (N_36697,N_36252,N_36449);
or U36698 (N_36698,N_36297,N_36379);
nand U36699 (N_36699,N_36312,N_36455);
or U36700 (N_36700,N_36311,N_36350);
or U36701 (N_36701,N_36471,N_36395);
and U36702 (N_36702,N_36422,N_36268);
and U36703 (N_36703,N_36425,N_36463);
and U36704 (N_36704,N_36400,N_36321);
nor U36705 (N_36705,N_36291,N_36492);
xnor U36706 (N_36706,N_36262,N_36311);
nor U36707 (N_36707,N_36366,N_36308);
xor U36708 (N_36708,N_36263,N_36402);
or U36709 (N_36709,N_36348,N_36447);
or U36710 (N_36710,N_36459,N_36381);
nor U36711 (N_36711,N_36256,N_36349);
and U36712 (N_36712,N_36438,N_36408);
or U36713 (N_36713,N_36468,N_36267);
xnor U36714 (N_36714,N_36421,N_36283);
or U36715 (N_36715,N_36322,N_36272);
xor U36716 (N_36716,N_36469,N_36331);
nor U36717 (N_36717,N_36268,N_36376);
nor U36718 (N_36718,N_36343,N_36274);
nor U36719 (N_36719,N_36356,N_36487);
or U36720 (N_36720,N_36409,N_36309);
and U36721 (N_36721,N_36490,N_36280);
and U36722 (N_36722,N_36317,N_36406);
nor U36723 (N_36723,N_36411,N_36287);
and U36724 (N_36724,N_36448,N_36299);
nand U36725 (N_36725,N_36420,N_36285);
or U36726 (N_36726,N_36438,N_36294);
or U36727 (N_36727,N_36463,N_36472);
or U36728 (N_36728,N_36363,N_36366);
or U36729 (N_36729,N_36467,N_36345);
or U36730 (N_36730,N_36421,N_36327);
xor U36731 (N_36731,N_36266,N_36356);
and U36732 (N_36732,N_36294,N_36499);
nor U36733 (N_36733,N_36425,N_36464);
nor U36734 (N_36734,N_36490,N_36331);
nand U36735 (N_36735,N_36310,N_36443);
and U36736 (N_36736,N_36426,N_36423);
or U36737 (N_36737,N_36336,N_36429);
or U36738 (N_36738,N_36489,N_36418);
nand U36739 (N_36739,N_36497,N_36490);
and U36740 (N_36740,N_36293,N_36324);
nor U36741 (N_36741,N_36483,N_36362);
nand U36742 (N_36742,N_36462,N_36367);
nor U36743 (N_36743,N_36264,N_36463);
or U36744 (N_36744,N_36310,N_36354);
xor U36745 (N_36745,N_36337,N_36381);
and U36746 (N_36746,N_36313,N_36341);
nor U36747 (N_36747,N_36332,N_36270);
xor U36748 (N_36748,N_36296,N_36378);
xnor U36749 (N_36749,N_36309,N_36342);
and U36750 (N_36750,N_36680,N_36720);
or U36751 (N_36751,N_36658,N_36641);
and U36752 (N_36752,N_36667,N_36648);
or U36753 (N_36753,N_36608,N_36559);
or U36754 (N_36754,N_36504,N_36611);
or U36755 (N_36755,N_36689,N_36687);
xnor U36756 (N_36756,N_36676,N_36622);
xor U36757 (N_36757,N_36731,N_36515);
or U36758 (N_36758,N_36508,N_36690);
xor U36759 (N_36759,N_36519,N_36661);
and U36760 (N_36760,N_36694,N_36672);
nand U36761 (N_36761,N_36742,N_36710);
and U36762 (N_36762,N_36505,N_36696);
or U36763 (N_36763,N_36713,N_36637);
xor U36764 (N_36764,N_36551,N_36516);
xnor U36765 (N_36765,N_36591,N_36588);
xnor U36766 (N_36766,N_36502,N_36615);
nand U36767 (N_36767,N_36670,N_36617);
and U36768 (N_36768,N_36619,N_36522);
nand U36769 (N_36769,N_36703,N_36570);
and U36770 (N_36770,N_36527,N_36587);
or U36771 (N_36771,N_36717,N_36579);
xnor U36772 (N_36772,N_36701,N_36595);
nor U36773 (N_36773,N_36698,N_36653);
or U36774 (N_36774,N_36674,N_36733);
or U36775 (N_36775,N_36652,N_36517);
or U36776 (N_36776,N_36590,N_36691);
and U36777 (N_36777,N_36634,N_36639);
xnor U36778 (N_36778,N_36668,N_36663);
xnor U36779 (N_36779,N_36735,N_36620);
and U36780 (N_36780,N_36643,N_36649);
nor U36781 (N_36781,N_36707,N_36708);
and U36782 (N_36782,N_36521,N_36654);
or U36783 (N_36783,N_36700,N_36656);
or U36784 (N_36784,N_36610,N_36728);
or U36785 (N_36785,N_36638,N_36603);
or U36786 (N_36786,N_36518,N_36704);
xor U36787 (N_36787,N_36660,N_36623);
xor U36788 (N_36788,N_36514,N_36709);
and U36789 (N_36789,N_36600,N_36596);
and U36790 (N_36790,N_36627,N_36593);
or U36791 (N_36791,N_36509,N_36578);
or U36792 (N_36792,N_36726,N_36673);
nor U36793 (N_36793,N_36734,N_36534);
nand U36794 (N_36794,N_36659,N_36538);
and U36795 (N_36795,N_36662,N_36692);
and U36796 (N_36796,N_36568,N_36605);
and U36797 (N_36797,N_36586,N_36614);
or U36798 (N_36798,N_36724,N_36635);
or U36799 (N_36799,N_36729,N_36714);
and U36800 (N_36800,N_36565,N_36718);
or U36801 (N_36801,N_36618,N_36739);
and U36802 (N_36802,N_36530,N_36589);
and U36803 (N_36803,N_36548,N_36512);
or U36804 (N_36804,N_36598,N_36630);
and U36805 (N_36805,N_36582,N_36539);
nor U36806 (N_36806,N_36552,N_36669);
and U36807 (N_36807,N_36632,N_36543);
and U36808 (N_36808,N_36723,N_36646);
and U36809 (N_36809,N_36715,N_36712);
xor U36810 (N_36810,N_36686,N_36562);
or U36811 (N_36811,N_36592,N_36736);
or U36812 (N_36812,N_36609,N_36688);
xor U36813 (N_36813,N_36647,N_36563);
xnor U36814 (N_36814,N_36599,N_36666);
and U36815 (N_36815,N_36584,N_36681);
or U36816 (N_36816,N_36741,N_36711);
nand U36817 (N_36817,N_36645,N_36738);
or U36818 (N_36818,N_36746,N_36747);
nor U36819 (N_36819,N_36531,N_36601);
and U36820 (N_36820,N_36693,N_36544);
nor U36821 (N_36821,N_36640,N_36613);
xnor U36822 (N_36822,N_36557,N_36725);
or U36823 (N_36823,N_36561,N_36664);
nor U36824 (N_36824,N_36500,N_36555);
nor U36825 (N_36825,N_36625,N_36706);
or U36826 (N_36826,N_36684,N_36574);
nor U36827 (N_36827,N_36644,N_36526);
and U36828 (N_36828,N_36536,N_36671);
nand U36829 (N_36829,N_36567,N_36629);
nor U36830 (N_36830,N_36541,N_36730);
xnor U36831 (N_36831,N_36520,N_36604);
nand U36832 (N_36832,N_36727,N_36537);
xnor U36833 (N_36833,N_36507,N_36510);
or U36834 (N_36834,N_36597,N_36651);
or U36835 (N_36835,N_36683,N_36607);
and U36836 (N_36836,N_36553,N_36513);
and U36837 (N_36837,N_36554,N_36524);
or U36838 (N_36838,N_36564,N_36722);
nor U36839 (N_36839,N_36716,N_36525);
and U36840 (N_36840,N_36699,N_36523);
or U36841 (N_36841,N_36577,N_36575);
nor U36842 (N_36842,N_36558,N_36624);
xor U36843 (N_36843,N_36585,N_36685);
and U36844 (N_36844,N_36594,N_36581);
and U36845 (N_36845,N_36628,N_36719);
or U36846 (N_36846,N_36642,N_36556);
nor U36847 (N_36847,N_36540,N_36547);
nand U36848 (N_36848,N_36580,N_36612);
nor U36849 (N_36849,N_36573,N_36657);
xnor U36850 (N_36850,N_36721,N_36743);
and U36851 (N_36851,N_36576,N_36732);
nor U36852 (N_36852,N_36702,N_36675);
nor U36853 (N_36853,N_36569,N_36549);
or U36854 (N_36854,N_36744,N_36546);
and U36855 (N_36855,N_36737,N_36678);
xor U36856 (N_36856,N_36745,N_36633);
nand U36857 (N_36857,N_36572,N_36631);
nor U36858 (N_36858,N_36529,N_36535);
and U36859 (N_36859,N_36650,N_36655);
nor U36860 (N_36860,N_36542,N_36550);
nand U36861 (N_36861,N_36503,N_36583);
and U36862 (N_36862,N_36533,N_36566);
nor U36863 (N_36863,N_36705,N_36697);
xor U36864 (N_36864,N_36606,N_36626);
xnor U36865 (N_36865,N_36616,N_36528);
nor U36866 (N_36866,N_36602,N_36636);
nand U36867 (N_36867,N_36695,N_36506);
or U36868 (N_36868,N_36682,N_36560);
or U36869 (N_36869,N_36749,N_36511);
and U36870 (N_36870,N_36501,N_36621);
or U36871 (N_36871,N_36679,N_36740);
and U36872 (N_36872,N_36545,N_36748);
nand U36873 (N_36873,N_36532,N_36677);
nand U36874 (N_36874,N_36665,N_36571);
or U36875 (N_36875,N_36642,N_36623);
nor U36876 (N_36876,N_36604,N_36583);
nand U36877 (N_36877,N_36575,N_36623);
or U36878 (N_36878,N_36699,N_36708);
or U36879 (N_36879,N_36520,N_36712);
xnor U36880 (N_36880,N_36640,N_36558);
or U36881 (N_36881,N_36649,N_36701);
or U36882 (N_36882,N_36536,N_36656);
nor U36883 (N_36883,N_36556,N_36623);
or U36884 (N_36884,N_36665,N_36738);
nor U36885 (N_36885,N_36691,N_36535);
nor U36886 (N_36886,N_36599,N_36580);
and U36887 (N_36887,N_36573,N_36723);
xnor U36888 (N_36888,N_36712,N_36731);
xnor U36889 (N_36889,N_36570,N_36565);
nor U36890 (N_36890,N_36544,N_36568);
nand U36891 (N_36891,N_36661,N_36721);
nor U36892 (N_36892,N_36557,N_36736);
or U36893 (N_36893,N_36702,N_36523);
or U36894 (N_36894,N_36731,N_36645);
xnor U36895 (N_36895,N_36617,N_36735);
and U36896 (N_36896,N_36746,N_36625);
or U36897 (N_36897,N_36670,N_36509);
and U36898 (N_36898,N_36510,N_36691);
xnor U36899 (N_36899,N_36668,N_36505);
and U36900 (N_36900,N_36642,N_36530);
and U36901 (N_36901,N_36684,N_36674);
nor U36902 (N_36902,N_36586,N_36720);
and U36903 (N_36903,N_36601,N_36697);
or U36904 (N_36904,N_36651,N_36614);
nand U36905 (N_36905,N_36501,N_36719);
nand U36906 (N_36906,N_36632,N_36544);
or U36907 (N_36907,N_36566,N_36729);
and U36908 (N_36908,N_36624,N_36722);
nand U36909 (N_36909,N_36691,N_36679);
xnor U36910 (N_36910,N_36682,N_36665);
xnor U36911 (N_36911,N_36566,N_36605);
and U36912 (N_36912,N_36618,N_36541);
or U36913 (N_36913,N_36684,N_36503);
nand U36914 (N_36914,N_36618,N_36593);
and U36915 (N_36915,N_36600,N_36612);
and U36916 (N_36916,N_36725,N_36736);
nor U36917 (N_36917,N_36722,N_36590);
and U36918 (N_36918,N_36739,N_36571);
xnor U36919 (N_36919,N_36743,N_36603);
nor U36920 (N_36920,N_36685,N_36747);
xnor U36921 (N_36921,N_36720,N_36619);
nand U36922 (N_36922,N_36586,N_36525);
xnor U36923 (N_36923,N_36744,N_36739);
nand U36924 (N_36924,N_36514,N_36664);
xor U36925 (N_36925,N_36570,N_36630);
xnor U36926 (N_36926,N_36676,N_36500);
nor U36927 (N_36927,N_36553,N_36526);
and U36928 (N_36928,N_36669,N_36662);
nor U36929 (N_36929,N_36642,N_36678);
and U36930 (N_36930,N_36737,N_36562);
or U36931 (N_36931,N_36556,N_36610);
xor U36932 (N_36932,N_36584,N_36744);
and U36933 (N_36933,N_36519,N_36644);
or U36934 (N_36934,N_36734,N_36555);
or U36935 (N_36935,N_36666,N_36536);
and U36936 (N_36936,N_36623,N_36558);
or U36937 (N_36937,N_36530,N_36547);
or U36938 (N_36938,N_36719,N_36641);
and U36939 (N_36939,N_36560,N_36677);
nand U36940 (N_36940,N_36654,N_36541);
nor U36941 (N_36941,N_36670,N_36702);
or U36942 (N_36942,N_36599,N_36675);
and U36943 (N_36943,N_36509,N_36594);
nand U36944 (N_36944,N_36558,N_36653);
and U36945 (N_36945,N_36630,N_36731);
or U36946 (N_36946,N_36508,N_36573);
and U36947 (N_36947,N_36698,N_36661);
nand U36948 (N_36948,N_36731,N_36589);
xor U36949 (N_36949,N_36574,N_36739);
nor U36950 (N_36950,N_36744,N_36636);
nor U36951 (N_36951,N_36542,N_36604);
nor U36952 (N_36952,N_36534,N_36626);
or U36953 (N_36953,N_36703,N_36729);
nor U36954 (N_36954,N_36605,N_36509);
or U36955 (N_36955,N_36721,N_36517);
xor U36956 (N_36956,N_36709,N_36596);
xor U36957 (N_36957,N_36519,N_36673);
xnor U36958 (N_36958,N_36670,N_36535);
and U36959 (N_36959,N_36560,N_36559);
nand U36960 (N_36960,N_36665,N_36634);
or U36961 (N_36961,N_36726,N_36731);
nor U36962 (N_36962,N_36567,N_36649);
or U36963 (N_36963,N_36550,N_36635);
nand U36964 (N_36964,N_36581,N_36714);
or U36965 (N_36965,N_36710,N_36643);
and U36966 (N_36966,N_36534,N_36595);
nand U36967 (N_36967,N_36712,N_36608);
xnor U36968 (N_36968,N_36690,N_36522);
and U36969 (N_36969,N_36740,N_36518);
and U36970 (N_36970,N_36521,N_36733);
and U36971 (N_36971,N_36676,N_36526);
nor U36972 (N_36972,N_36577,N_36660);
xor U36973 (N_36973,N_36561,N_36699);
nand U36974 (N_36974,N_36563,N_36711);
or U36975 (N_36975,N_36660,N_36525);
nand U36976 (N_36976,N_36642,N_36541);
xnor U36977 (N_36977,N_36607,N_36567);
nand U36978 (N_36978,N_36738,N_36600);
nor U36979 (N_36979,N_36691,N_36530);
nor U36980 (N_36980,N_36675,N_36586);
or U36981 (N_36981,N_36520,N_36608);
or U36982 (N_36982,N_36649,N_36528);
nor U36983 (N_36983,N_36717,N_36674);
xor U36984 (N_36984,N_36725,N_36728);
nor U36985 (N_36985,N_36644,N_36735);
and U36986 (N_36986,N_36740,N_36588);
nand U36987 (N_36987,N_36582,N_36538);
xor U36988 (N_36988,N_36699,N_36603);
nand U36989 (N_36989,N_36615,N_36647);
xnor U36990 (N_36990,N_36550,N_36607);
nand U36991 (N_36991,N_36705,N_36652);
and U36992 (N_36992,N_36701,N_36689);
nor U36993 (N_36993,N_36664,N_36551);
nor U36994 (N_36994,N_36733,N_36640);
and U36995 (N_36995,N_36521,N_36544);
and U36996 (N_36996,N_36739,N_36690);
and U36997 (N_36997,N_36687,N_36749);
xor U36998 (N_36998,N_36596,N_36672);
nand U36999 (N_36999,N_36591,N_36648);
and U37000 (N_37000,N_36946,N_36870);
and U37001 (N_37001,N_36830,N_36767);
xnor U37002 (N_37002,N_36853,N_36852);
or U37003 (N_37003,N_36765,N_36943);
nand U37004 (N_37004,N_36976,N_36937);
xnor U37005 (N_37005,N_36820,N_36956);
and U37006 (N_37006,N_36944,N_36773);
and U37007 (N_37007,N_36993,N_36818);
and U37008 (N_37008,N_36903,N_36790);
and U37009 (N_37009,N_36823,N_36955);
and U37010 (N_37010,N_36966,N_36947);
nand U37011 (N_37011,N_36890,N_36856);
nor U37012 (N_37012,N_36928,N_36791);
or U37013 (N_37013,N_36807,N_36828);
or U37014 (N_37014,N_36922,N_36910);
and U37015 (N_37015,N_36926,N_36951);
or U37016 (N_37016,N_36838,N_36876);
nand U37017 (N_37017,N_36835,N_36898);
nor U37018 (N_37018,N_36771,N_36757);
or U37019 (N_37019,N_36932,N_36864);
and U37020 (N_37020,N_36836,N_36789);
nor U37021 (N_37021,N_36999,N_36760);
xnor U37022 (N_37022,N_36810,N_36840);
nor U37023 (N_37023,N_36822,N_36925);
xor U37024 (N_37024,N_36904,N_36848);
nand U37025 (N_37025,N_36874,N_36972);
or U37026 (N_37026,N_36968,N_36896);
and U37027 (N_37027,N_36970,N_36845);
nor U37028 (N_37028,N_36923,N_36986);
nor U37029 (N_37029,N_36973,N_36885);
nand U37030 (N_37030,N_36829,N_36819);
nand U37031 (N_37031,N_36984,N_36872);
xor U37032 (N_37032,N_36877,N_36935);
xor U37033 (N_37033,N_36803,N_36906);
nand U37034 (N_37034,N_36763,N_36770);
and U37035 (N_37035,N_36994,N_36891);
or U37036 (N_37036,N_36897,N_36957);
or U37037 (N_37037,N_36756,N_36806);
and U37038 (N_37038,N_36918,N_36815);
or U37039 (N_37039,N_36774,N_36964);
nand U37040 (N_37040,N_36905,N_36792);
xnor U37041 (N_37041,N_36758,N_36971);
xor U37042 (N_37042,N_36913,N_36768);
nand U37043 (N_37043,N_36772,N_36762);
nor U37044 (N_37044,N_36875,N_36814);
xnor U37045 (N_37045,N_36959,N_36952);
nor U37046 (N_37046,N_36826,N_36857);
or U37047 (N_37047,N_36858,N_36786);
xnor U37048 (N_37048,N_36886,N_36980);
nor U37049 (N_37049,N_36802,N_36839);
or U37050 (N_37050,N_36827,N_36778);
or U37051 (N_37051,N_36990,N_36843);
or U37052 (N_37052,N_36987,N_36793);
xnor U37053 (N_37053,N_36854,N_36974);
xnor U37054 (N_37054,N_36779,N_36794);
and U37055 (N_37055,N_36764,N_36834);
xor U37056 (N_37056,N_36961,N_36788);
or U37057 (N_37057,N_36983,N_36750);
or U37058 (N_37058,N_36900,N_36855);
xnor U37059 (N_37059,N_36908,N_36929);
nor U37060 (N_37060,N_36809,N_36945);
nand U37061 (N_37061,N_36780,N_36996);
nor U37062 (N_37062,N_36895,N_36920);
nor U37063 (N_37063,N_36958,N_36963);
xnor U37064 (N_37064,N_36909,N_36927);
xor U37065 (N_37065,N_36969,N_36901);
xor U37066 (N_37066,N_36784,N_36776);
and U37067 (N_37067,N_36954,N_36914);
or U37068 (N_37068,N_36883,N_36936);
or U37069 (N_37069,N_36881,N_36934);
xor U37070 (N_37070,N_36754,N_36907);
and U37071 (N_37071,N_36950,N_36953);
xnor U37072 (N_37072,N_36805,N_36862);
xor U37073 (N_37073,N_36981,N_36884);
or U37074 (N_37074,N_36832,N_36833);
and U37075 (N_37075,N_36782,N_36975);
and U37076 (N_37076,N_36992,N_36844);
or U37077 (N_37077,N_36893,N_36880);
nor U37078 (N_37078,N_36911,N_36785);
nand U37079 (N_37079,N_36948,N_36931);
and U37080 (N_37080,N_36861,N_36821);
xor U37081 (N_37081,N_36801,N_36985);
xor U37082 (N_37082,N_36982,N_36787);
and U37083 (N_37083,N_36869,N_36894);
xor U37084 (N_37084,N_36995,N_36977);
xnor U37085 (N_37085,N_36837,N_36991);
and U37086 (N_37086,N_36759,N_36997);
xnor U37087 (N_37087,N_36824,N_36939);
nor U37088 (N_37088,N_36808,N_36781);
xor U37089 (N_37089,N_36938,N_36878);
xnor U37090 (N_37090,N_36799,N_36860);
xor U37091 (N_37091,N_36859,N_36783);
xor U37092 (N_37092,N_36775,N_36879);
xor U37093 (N_37093,N_36912,N_36841);
and U37094 (N_37094,N_36755,N_36800);
nand U37095 (N_37095,N_36998,N_36921);
nand U37096 (N_37096,N_36919,N_36949);
and U37097 (N_37097,N_36777,N_36978);
or U37098 (N_37098,N_36989,N_36850);
or U37099 (N_37099,N_36941,N_36873);
nand U37100 (N_37100,N_36804,N_36915);
or U37101 (N_37101,N_36882,N_36863);
nor U37102 (N_37102,N_36962,N_36979);
or U37103 (N_37103,N_36796,N_36892);
nor U37104 (N_37104,N_36924,N_36889);
nand U37105 (N_37105,N_36988,N_36825);
nand U37106 (N_37106,N_36868,N_36798);
or U37107 (N_37107,N_36842,N_36887);
nand U37108 (N_37108,N_36813,N_36811);
nand U37109 (N_37109,N_36797,N_36866);
xnor U37110 (N_37110,N_36751,N_36930);
or U37111 (N_37111,N_36752,N_36960);
and U37112 (N_37112,N_36766,N_36761);
or U37113 (N_37113,N_36967,N_36849);
and U37114 (N_37114,N_36867,N_36899);
or U37115 (N_37115,N_36942,N_36795);
xnor U37116 (N_37116,N_36831,N_36816);
and U37117 (N_37117,N_36940,N_36865);
or U37118 (N_37118,N_36769,N_36871);
nor U37119 (N_37119,N_36933,N_36917);
nor U37120 (N_37120,N_36902,N_36851);
and U37121 (N_37121,N_36817,N_36812);
nor U37122 (N_37122,N_36888,N_36916);
and U37123 (N_37123,N_36965,N_36847);
xor U37124 (N_37124,N_36846,N_36753);
or U37125 (N_37125,N_36874,N_36940);
nand U37126 (N_37126,N_36826,N_36787);
and U37127 (N_37127,N_36820,N_36977);
or U37128 (N_37128,N_36948,N_36808);
or U37129 (N_37129,N_36890,N_36960);
nor U37130 (N_37130,N_36764,N_36780);
nor U37131 (N_37131,N_36968,N_36919);
nor U37132 (N_37132,N_36851,N_36998);
nand U37133 (N_37133,N_36785,N_36786);
or U37134 (N_37134,N_36992,N_36783);
or U37135 (N_37135,N_36851,N_36890);
nor U37136 (N_37136,N_36789,N_36903);
nand U37137 (N_37137,N_36811,N_36975);
xor U37138 (N_37138,N_36941,N_36901);
nand U37139 (N_37139,N_36858,N_36755);
and U37140 (N_37140,N_36969,N_36973);
nor U37141 (N_37141,N_36899,N_36920);
xnor U37142 (N_37142,N_36750,N_36803);
xor U37143 (N_37143,N_36867,N_36813);
and U37144 (N_37144,N_36977,N_36880);
nor U37145 (N_37145,N_36950,N_36993);
nand U37146 (N_37146,N_36915,N_36878);
and U37147 (N_37147,N_36946,N_36890);
nand U37148 (N_37148,N_36960,N_36759);
and U37149 (N_37149,N_36919,N_36887);
xnor U37150 (N_37150,N_36796,N_36994);
nor U37151 (N_37151,N_36757,N_36808);
or U37152 (N_37152,N_36995,N_36816);
nor U37153 (N_37153,N_36951,N_36886);
nand U37154 (N_37154,N_36898,N_36997);
nor U37155 (N_37155,N_36830,N_36843);
nand U37156 (N_37156,N_36818,N_36771);
xor U37157 (N_37157,N_36839,N_36960);
nor U37158 (N_37158,N_36801,N_36810);
or U37159 (N_37159,N_36824,N_36987);
xnor U37160 (N_37160,N_36852,N_36947);
and U37161 (N_37161,N_36827,N_36959);
xnor U37162 (N_37162,N_36951,N_36804);
nor U37163 (N_37163,N_36884,N_36816);
nand U37164 (N_37164,N_36868,N_36767);
xnor U37165 (N_37165,N_36842,N_36994);
or U37166 (N_37166,N_36784,N_36847);
nor U37167 (N_37167,N_36927,N_36963);
xnor U37168 (N_37168,N_36787,N_36773);
and U37169 (N_37169,N_36778,N_36782);
nand U37170 (N_37170,N_36799,N_36903);
xor U37171 (N_37171,N_36852,N_36938);
and U37172 (N_37172,N_36969,N_36941);
nand U37173 (N_37173,N_36936,N_36908);
nand U37174 (N_37174,N_36903,N_36807);
and U37175 (N_37175,N_36771,N_36908);
and U37176 (N_37176,N_36913,N_36890);
nor U37177 (N_37177,N_36902,N_36819);
and U37178 (N_37178,N_36995,N_36750);
and U37179 (N_37179,N_36885,N_36877);
xor U37180 (N_37180,N_36828,N_36905);
or U37181 (N_37181,N_36945,N_36791);
xnor U37182 (N_37182,N_36803,N_36933);
nor U37183 (N_37183,N_36993,N_36873);
nor U37184 (N_37184,N_36912,N_36788);
or U37185 (N_37185,N_36863,N_36784);
nand U37186 (N_37186,N_36786,N_36946);
xor U37187 (N_37187,N_36977,N_36756);
nand U37188 (N_37188,N_36974,N_36824);
nor U37189 (N_37189,N_36929,N_36803);
nand U37190 (N_37190,N_36756,N_36875);
or U37191 (N_37191,N_36902,N_36820);
nand U37192 (N_37192,N_36809,N_36803);
xor U37193 (N_37193,N_36791,N_36868);
xor U37194 (N_37194,N_36824,N_36935);
nand U37195 (N_37195,N_36921,N_36815);
and U37196 (N_37196,N_36799,N_36812);
or U37197 (N_37197,N_36759,N_36767);
nand U37198 (N_37198,N_36977,N_36825);
nor U37199 (N_37199,N_36828,N_36988);
and U37200 (N_37200,N_36845,N_36886);
xnor U37201 (N_37201,N_36777,N_36887);
or U37202 (N_37202,N_36988,N_36936);
xnor U37203 (N_37203,N_36859,N_36752);
nor U37204 (N_37204,N_36947,N_36940);
xor U37205 (N_37205,N_36773,N_36876);
or U37206 (N_37206,N_36901,N_36975);
and U37207 (N_37207,N_36825,N_36908);
nor U37208 (N_37208,N_36967,N_36925);
and U37209 (N_37209,N_36884,N_36905);
xnor U37210 (N_37210,N_36834,N_36762);
and U37211 (N_37211,N_36780,N_36959);
nor U37212 (N_37212,N_36772,N_36896);
xor U37213 (N_37213,N_36848,N_36887);
nand U37214 (N_37214,N_36859,N_36989);
nor U37215 (N_37215,N_36794,N_36776);
nor U37216 (N_37216,N_36837,N_36997);
or U37217 (N_37217,N_36842,N_36934);
or U37218 (N_37218,N_36844,N_36991);
or U37219 (N_37219,N_36756,N_36866);
nor U37220 (N_37220,N_36882,N_36858);
or U37221 (N_37221,N_36808,N_36840);
nor U37222 (N_37222,N_36973,N_36751);
and U37223 (N_37223,N_36961,N_36752);
nor U37224 (N_37224,N_36912,N_36992);
and U37225 (N_37225,N_36865,N_36936);
or U37226 (N_37226,N_36774,N_36958);
xnor U37227 (N_37227,N_36768,N_36977);
nor U37228 (N_37228,N_36853,N_36906);
xor U37229 (N_37229,N_36938,N_36756);
or U37230 (N_37230,N_36874,N_36980);
nand U37231 (N_37231,N_36757,N_36810);
and U37232 (N_37232,N_36751,N_36868);
xor U37233 (N_37233,N_36954,N_36934);
and U37234 (N_37234,N_36872,N_36783);
xnor U37235 (N_37235,N_36876,N_36769);
or U37236 (N_37236,N_36954,N_36871);
nand U37237 (N_37237,N_36825,N_36772);
and U37238 (N_37238,N_36785,N_36755);
or U37239 (N_37239,N_36843,N_36809);
or U37240 (N_37240,N_36995,N_36785);
or U37241 (N_37241,N_36894,N_36878);
nand U37242 (N_37242,N_36792,N_36914);
or U37243 (N_37243,N_36838,N_36881);
nor U37244 (N_37244,N_36916,N_36834);
nor U37245 (N_37245,N_36807,N_36951);
nand U37246 (N_37246,N_36897,N_36783);
nand U37247 (N_37247,N_36963,N_36921);
xor U37248 (N_37248,N_36826,N_36758);
and U37249 (N_37249,N_36845,N_36907);
and U37250 (N_37250,N_37059,N_37145);
nand U37251 (N_37251,N_37113,N_37052);
or U37252 (N_37252,N_37179,N_37181);
nor U37253 (N_37253,N_37075,N_37242);
nor U37254 (N_37254,N_37132,N_37177);
and U37255 (N_37255,N_37044,N_37225);
nand U37256 (N_37256,N_37019,N_37119);
nor U37257 (N_37257,N_37222,N_37175);
or U37258 (N_37258,N_37042,N_37227);
and U37259 (N_37259,N_37093,N_37095);
nand U37260 (N_37260,N_37065,N_37156);
or U37261 (N_37261,N_37055,N_37131);
xor U37262 (N_37262,N_37134,N_37069);
nand U37263 (N_37263,N_37161,N_37171);
nand U37264 (N_37264,N_37232,N_37192);
nand U37265 (N_37265,N_37207,N_37043);
nor U37266 (N_37266,N_37010,N_37153);
nand U37267 (N_37267,N_37048,N_37186);
and U37268 (N_37268,N_37117,N_37092);
nand U37269 (N_37269,N_37223,N_37024);
xnor U37270 (N_37270,N_37185,N_37082);
and U37271 (N_37271,N_37220,N_37146);
and U37272 (N_37272,N_37051,N_37032);
and U37273 (N_37273,N_37150,N_37229);
nand U37274 (N_37274,N_37204,N_37080);
nand U37275 (N_37275,N_37231,N_37169);
and U37276 (N_37276,N_37111,N_37138);
nor U37277 (N_37277,N_37187,N_37041);
and U37278 (N_37278,N_37123,N_37026);
nor U37279 (N_37279,N_37147,N_37205);
and U37280 (N_37280,N_37004,N_37139);
or U37281 (N_37281,N_37144,N_37040);
nand U37282 (N_37282,N_37249,N_37128);
nor U37283 (N_37283,N_37101,N_37083);
or U37284 (N_37284,N_37163,N_37200);
nor U37285 (N_37285,N_37039,N_37058);
nand U37286 (N_37286,N_37072,N_37151);
nand U37287 (N_37287,N_37049,N_37214);
nand U37288 (N_37288,N_37062,N_37014);
and U37289 (N_37289,N_37209,N_37215);
nor U37290 (N_37290,N_37003,N_37236);
or U37291 (N_37291,N_37164,N_37110);
nand U37292 (N_37292,N_37121,N_37140);
or U37293 (N_37293,N_37118,N_37074);
nor U37294 (N_37294,N_37099,N_37028);
or U37295 (N_37295,N_37071,N_37063);
and U37296 (N_37296,N_37212,N_37029);
xor U37297 (N_37297,N_37087,N_37016);
and U37298 (N_37298,N_37245,N_37105);
nor U37299 (N_37299,N_37114,N_37213);
or U37300 (N_37300,N_37085,N_37203);
nand U37301 (N_37301,N_37170,N_37217);
and U37302 (N_37302,N_37135,N_37188);
or U37303 (N_37303,N_37173,N_37027);
xor U37304 (N_37304,N_37006,N_37208);
xnor U37305 (N_37305,N_37096,N_37034);
xor U37306 (N_37306,N_37194,N_37184);
and U37307 (N_37307,N_37178,N_37104);
xor U37308 (N_37308,N_37002,N_37176);
and U37309 (N_37309,N_37077,N_37219);
and U37310 (N_37310,N_37155,N_37218);
and U37311 (N_37311,N_37073,N_37247);
and U37312 (N_37312,N_37122,N_37070);
nand U37313 (N_37313,N_37018,N_37091);
or U37314 (N_37314,N_37050,N_37120);
and U37315 (N_37315,N_37224,N_37168);
nand U37316 (N_37316,N_37025,N_37240);
nor U37317 (N_37317,N_37166,N_37127);
or U37318 (N_37318,N_37103,N_37180);
nand U37319 (N_37319,N_37015,N_37124);
or U37320 (N_37320,N_37081,N_37244);
and U37321 (N_37321,N_37159,N_37246);
xor U37322 (N_37322,N_37035,N_37202);
xnor U37323 (N_37323,N_37211,N_37013);
nor U37324 (N_37324,N_37076,N_37143);
nand U37325 (N_37325,N_37109,N_37154);
or U37326 (N_37326,N_37053,N_37061);
xnor U37327 (N_37327,N_37198,N_37129);
or U37328 (N_37328,N_37089,N_37102);
nand U37329 (N_37329,N_37001,N_37221);
or U37330 (N_37330,N_37116,N_37189);
nand U37331 (N_37331,N_37084,N_37088);
xor U37332 (N_37332,N_37125,N_37097);
nand U37333 (N_37333,N_37130,N_37158);
nand U37334 (N_37334,N_37115,N_37190);
nor U37335 (N_37335,N_37141,N_37210);
nor U37336 (N_37336,N_37165,N_37183);
xor U37337 (N_37337,N_37056,N_37031);
nand U37338 (N_37338,N_37136,N_37107);
or U37339 (N_37339,N_37191,N_37036);
and U37340 (N_37340,N_37008,N_37226);
nor U37341 (N_37341,N_37067,N_37248);
or U37342 (N_37342,N_37157,N_37167);
nor U37343 (N_37343,N_37235,N_37086);
or U37344 (N_37344,N_37182,N_37112);
nand U37345 (N_37345,N_37195,N_37007);
xnor U37346 (N_37346,N_37037,N_37137);
or U37347 (N_37347,N_37239,N_37094);
xor U37348 (N_37348,N_37106,N_37233);
nand U37349 (N_37349,N_37199,N_37142);
and U37350 (N_37350,N_37162,N_37047);
and U37351 (N_37351,N_37193,N_37100);
or U37352 (N_37352,N_37172,N_37149);
and U37353 (N_37353,N_37237,N_37160);
and U37354 (N_37354,N_37197,N_37064);
or U37355 (N_37355,N_37090,N_37020);
nor U37356 (N_37356,N_37012,N_37230);
nor U37357 (N_37357,N_37243,N_37078);
and U37358 (N_37358,N_37057,N_37079);
xor U37359 (N_37359,N_37201,N_37046);
nor U37360 (N_37360,N_37216,N_37148);
xor U37361 (N_37361,N_37030,N_37206);
nor U37362 (N_37362,N_37033,N_37021);
and U37363 (N_37363,N_37054,N_37060);
nand U37364 (N_37364,N_37066,N_37108);
xor U37365 (N_37365,N_37022,N_37017);
or U37366 (N_37366,N_37133,N_37152);
and U37367 (N_37367,N_37228,N_37011);
xnor U37368 (N_37368,N_37174,N_37009);
and U37369 (N_37369,N_37098,N_37005);
and U37370 (N_37370,N_37238,N_37234);
nor U37371 (N_37371,N_37196,N_37241);
nor U37372 (N_37372,N_37038,N_37068);
nand U37373 (N_37373,N_37045,N_37023);
xor U37374 (N_37374,N_37000,N_37126);
xor U37375 (N_37375,N_37076,N_37118);
and U37376 (N_37376,N_37068,N_37025);
nor U37377 (N_37377,N_37142,N_37182);
or U37378 (N_37378,N_37222,N_37240);
xnor U37379 (N_37379,N_37142,N_37209);
and U37380 (N_37380,N_37037,N_37122);
nor U37381 (N_37381,N_37085,N_37064);
nor U37382 (N_37382,N_37207,N_37211);
nand U37383 (N_37383,N_37217,N_37033);
nor U37384 (N_37384,N_37110,N_37210);
xnor U37385 (N_37385,N_37116,N_37215);
or U37386 (N_37386,N_37200,N_37092);
nand U37387 (N_37387,N_37191,N_37196);
xor U37388 (N_37388,N_37206,N_37061);
or U37389 (N_37389,N_37204,N_37203);
xnor U37390 (N_37390,N_37172,N_37098);
or U37391 (N_37391,N_37015,N_37067);
and U37392 (N_37392,N_37153,N_37096);
and U37393 (N_37393,N_37105,N_37198);
xnor U37394 (N_37394,N_37008,N_37055);
nor U37395 (N_37395,N_37113,N_37026);
or U37396 (N_37396,N_37240,N_37068);
or U37397 (N_37397,N_37093,N_37117);
nand U37398 (N_37398,N_37177,N_37192);
or U37399 (N_37399,N_37013,N_37087);
nor U37400 (N_37400,N_37153,N_37178);
or U37401 (N_37401,N_37224,N_37064);
or U37402 (N_37402,N_37028,N_37216);
and U37403 (N_37403,N_37207,N_37081);
xor U37404 (N_37404,N_37043,N_37121);
or U37405 (N_37405,N_37202,N_37100);
and U37406 (N_37406,N_37018,N_37059);
and U37407 (N_37407,N_37235,N_37058);
nor U37408 (N_37408,N_37178,N_37013);
xnor U37409 (N_37409,N_37111,N_37144);
xor U37410 (N_37410,N_37182,N_37029);
and U37411 (N_37411,N_37212,N_37064);
nor U37412 (N_37412,N_37125,N_37079);
and U37413 (N_37413,N_37010,N_37204);
xor U37414 (N_37414,N_37000,N_37165);
nor U37415 (N_37415,N_37026,N_37232);
nor U37416 (N_37416,N_37128,N_37140);
and U37417 (N_37417,N_37217,N_37226);
or U37418 (N_37418,N_37050,N_37097);
nand U37419 (N_37419,N_37109,N_37026);
xnor U37420 (N_37420,N_37103,N_37188);
nor U37421 (N_37421,N_37095,N_37182);
nor U37422 (N_37422,N_37021,N_37071);
nor U37423 (N_37423,N_37126,N_37025);
and U37424 (N_37424,N_37041,N_37248);
nor U37425 (N_37425,N_37212,N_37244);
or U37426 (N_37426,N_37214,N_37158);
and U37427 (N_37427,N_37025,N_37191);
nand U37428 (N_37428,N_37244,N_37192);
or U37429 (N_37429,N_37089,N_37202);
nor U37430 (N_37430,N_37169,N_37172);
xnor U37431 (N_37431,N_37002,N_37238);
and U37432 (N_37432,N_37184,N_37217);
xor U37433 (N_37433,N_37029,N_37067);
nor U37434 (N_37434,N_37124,N_37125);
and U37435 (N_37435,N_37193,N_37094);
and U37436 (N_37436,N_37099,N_37003);
or U37437 (N_37437,N_37096,N_37047);
xor U37438 (N_37438,N_37163,N_37239);
or U37439 (N_37439,N_37166,N_37064);
nand U37440 (N_37440,N_37123,N_37044);
or U37441 (N_37441,N_37165,N_37218);
xnor U37442 (N_37442,N_37175,N_37193);
or U37443 (N_37443,N_37087,N_37075);
xor U37444 (N_37444,N_37132,N_37039);
or U37445 (N_37445,N_37063,N_37185);
or U37446 (N_37446,N_37014,N_37010);
nand U37447 (N_37447,N_37007,N_37082);
nand U37448 (N_37448,N_37114,N_37094);
or U37449 (N_37449,N_37185,N_37062);
and U37450 (N_37450,N_37005,N_37170);
nand U37451 (N_37451,N_37074,N_37033);
xnor U37452 (N_37452,N_37031,N_37131);
nand U37453 (N_37453,N_37147,N_37045);
and U37454 (N_37454,N_37068,N_37210);
or U37455 (N_37455,N_37157,N_37187);
nand U37456 (N_37456,N_37145,N_37160);
nand U37457 (N_37457,N_37176,N_37066);
and U37458 (N_37458,N_37075,N_37120);
nor U37459 (N_37459,N_37117,N_37132);
nor U37460 (N_37460,N_37190,N_37169);
nor U37461 (N_37461,N_37122,N_37026);
xnor U37462 (N_37462,N_37195,N_37142);
nor U37463 (N_37463,N_37027,N_37153);
xnor U37464 (N_37464,N_37028,N_37080);
nor U37465 (N_37465,N_37114,N_37023);
and U37466 (N_37466,N_37054,N_37152);
or U37467 (N_37467,N_37156,N_37220);
and U37468 (N_37468,N_37225,N_37107);
nand U37469 (N_37469,N_37017,N_37034);
and U37470 (N_37470,N_37042,N_37150);
nand U37471 (N_37471,N_37102,N_37158);
or U37472 (N_37472,N_37193,N_37151);
and U37473 (N_37473,N_37215,N_37140);
and U37474 (N_37474,N_37078,N_37013);
or U37475 (N_37475,N_37013,N_37133);
or U37476 (N_37476,N_37126,N_37121);
nand U37477 (N_37477,N_37063,N_37204);
and U37478 (N_37478,N_37189,N_37095);
xnor U37479 (N_37479,N_37022,N_37143);
and U37480 (N_37480,N_37244,N_37189);
and U37481 (N_37481,N_37020,N_37164);
and U37482 (N_37482,N_37070,N_37228);
xor U37483 (N_37483,N_37132,N_37144);
and U37484 (N_37484,N_37142,N_37105);
nand U37485 (N_37485,N_37059,N_37031);
nand U37486 (N_37486,N_37075,N_37029);
xor U37487 (N_37487,N_37016,N_37212);
nor U37488 (N_37488,N_37168,N_37075);
xor U37489 (N_37489,N_37235,N_37001);
nor U37490 (N_37490,N_37208,N_37243);
xor U37491 (N_37491,N_37181,N_37207);
xnor U37492 (N_37492,N_37142,N_37205);
xnor U37493 (N_37493,N_37225,N_37033);
and U37494 (N_37494,N_37001,N_37128);
nor U37495 (N_37495,N_37167,N_37052);
and U37496 (N_37496,N_37211,N_37138);
and U37497 (N_37497,N_37209,N_37047);
nand U37498 (N_37498,N_37085,N_37213);
nor U37499 (N_37499,N_37071,N_37116);
xor U37500 (N_37500,N_37480,N_37327);
or U37501 (N_37501,N_37365,N_37318);
and U37502 (N_37502,N_37380,N_37460);
or U37503 (N_37503,N_37344,N_37278);
nand U37504 (N_37504,N_37343,N_37442);
xnor U37505 (N_37505,N_37309,N_37307);
xor U37506 (N_37506,N_37405,N_37349);
or U37507 (N_37507,N_37446,N_37410);
nor U37508 (N_37508,N_37464,N_37257);
and U37509 (N_37509,N_37323,N_37485);
or U37510 (N_37510,N_37375,N_37435);
nand U37511 (N_37511,N_37261,N_37373);
xnor U37512 (N_37512,N_37374,N_37302);
nor U37513 (N_37513,N_37385,N_37461);
nand U37514 (N_37514,N_37250,N_37481);
xor U37515 (N_37515,N_37407,N_37372);
xnor U37516 (N_37516,N_37390,N_37472);
nor U37517 (N_37517,N_37311,N_37259);
xor U37518 (N_37518,N_37449,N_37324);
nand U37519 (N_37519,N_37333,N_37388);
or U37520 (N_37520,N_37326,N_37383);
or U37521 (N_37521,N_37494,N_37419);
and U37522 (N_37522,N_37378,N_37384);
nand U37523 (N_37523,N_37470,N_37444);
and U37524 (N_37524,N_37267,N_37382);
nor U37525 (N_37525,N_37379,N_37412);
or U37526 (N_37526,N_37296,N_37499);
or U37527 (N_37527,N_37489,N_37463);
and U37528 (N_37528,N_37424,N_37299);
xor U37529 (N_37529,N_37254,N_37342);
nand U37530 (N_37530,N_37406,N_37255);
nor U37531 (N_37531,N_37290,N_37303);
xor U37532 (N_37532,N_37468,N_37427);
nor U37533 (N_37533,N_37260,N_37325);
xnor U37534 (N_37534,N_37253,N_37403);
nand U37535 (N_37535,N_37476,N_37386);
or U37536 (N_37536,N_37288,N_37440);
or U37537 (N_37537,N_37484,N_37462);
and U37538 (N_37538,N_37471,N_37488);
xor U37539 (N_37539,N_37477,N_37371);
nor U37540 (N_37540,N_37358,N_37399);
xor U37541 (N_37541,N_37493,N_37421);
or U37542 (N_37542,N_37338,N_37429);
xnor U37543 (N_37543,N_37401,N_37448);
xor U37544 (N_37544,N_37496,N_37474);
nor U37545 (N_37545,N_37355,N_37331);
and U37546 (N_37546,N_37391,N_37491);
xor U37547 (N_37547,N_37443,N_37498);
nand U37548 (N_37548,N_37368,N_37347);
nand U37549 (N_37549,N_37396,N_37350);
nand U37550 (N_37550,N_37293,N_37418);
or U37551 (N_37551,N_37420,N_37300);
nand U37552 (N_37552,N_37425,N_37269);
nor U37553 (N_37553,N_37433,N_37256);
nand U37554 (N_37554,N_37426,N_37436);
xor U37555 (N_37555,N_37363,N_37319);
nand U37556 (N_37556,N_37273,N_37428);
nor U37557 (N_37557,N_37459,N_37367);
xnor U37558 (N_37558,N_37357,N_37422);
xor U37559 (N_37559,N_37352,N_37346);
or U37560 (N_37560,N_37297,N_37451);
or U37561 (N_37561,N_37364,N_37279);
or U37562 (N_37562,N_37411,N_37432);
or U37563 (N_37563,N_37437,N_37285);
or U37564 (N_37564,N_37306,N_37397);
nor U37565 (N_37565,N_37392,N_37370);
nand U37566 (N_37566,N_37286,N_37294);
and U37567 (N_37567,N_37252,N_37337);
and U37568 (N_37568,N_37409,N_37295);
xor U37569 (N_37569,N_37291,N_37495);
or U37570 (N_37570,N_37402,N_37465);
or U37571 (N_37571,N_37359,N_37467);
or U37572 (N_37572,N_37339,N_37265);
nand U37573 (N_37573,N_37282,N_37457);
nand U37574 (N_37574,N_37366,N_37345);
nand U37575 (N_37575,N_37335,N_37354);
nand U37576 (N_37576,N_37492,N_37361);
or U37577 (N_37577,N_37473,N_37312);
nand U37578 (N_37578,N_37455,N_37362);
xor U37579 (N_37579,N_37415,N_37351);
nand U37580 (N_37580,N_37272,N_37431);
nor U37581 (N_37581,N_37490,N_37315);
nand U37582 (N_37582,N_37398,N_37453);
and U37583 (N_37583,N_37292,N_37456);
nand U37584 (N_37584,N_37356,N_37353);
or U37585 (N_37585,N_37439,N_37348);
nor U37586 (N_37586,N_37369,N_37332);
or U37587 (N_37587,N_37284,N_37447);
nand U37588 (N_37588,N_37454,N_37276);
nand U37589 (N_37589,N_37376,N_37263);
xor U37590 (N_37590,N_37387,N_37264);
nor U37591 (N_37591,N_37283,N_37281);
nand U37592 (N_37592,N_37336,N_37404);
nor U37593 (N_37593,N_37434,N_37430);
nand U37594 (N_37594,N_37258,N_37274);
or U37595 (N_37595,N_37417,N_37486);
or U37596 (N_37596,N_37450,N_37314);
nand U37597 (N_37597,N_37483,N_37340);
and U37598 (N_37598,N_37289,N_37423);
nor U37599 (N_37599,N_37308,N_37320);
nor U37600 (N_37600,N_37445,N_37416);
xnor U37601 (N_37601,N_37305,N_37377);
or U37602 (N_37602,N_37280,N_37381);
nand U37603 (N_37603,N_37393,N_37389);
nor U37604 (N_37604,N_37497,N_37408);
xor U37605 (N_37605,N_37329,N_37395);
or U37606 (N_37606,N_37270,N_37287);
xnor U37607 (N_37607,N_37266,N_37301);
and U37608 (N_37608,N_37317,N_37394);
nand U37609 (N_37609,N_37360,N_37271);
nand U37610 (N_37610,N_37322,N_37330);
and U37611 (N_37611,N_37341,N_37251);
or U37612 (N_37612,N_37304,N_37413);
or U37613 (N_37613,N_37321,N_37400);
nor U37614 (N_37614,N_37441,N_37469);
or U37615 (N_37615,N_37316,N_37268);
nand U37616 (N_37616,N_37298,N_37482);
nor U37617 (N_37617,N_37458,N_37466);
and U37618 (N_37618,N_37310,N_37313);
nand U37619 (N_37619,N_37487,N_37262);
and U37620 (N_37620,N_37438,N_37478);
or U37621 (N_37621,N_37275,N_37414);
and U37622 (N_37622,N_37475,N_37479);
and U37623 (N_37623,N_37334,N_37328);
or U37624 (N_37624,N_37452,N_37277);
xnor U37625 (N_37625,N_37287,N_37340);
nor U37626 (N_37626,N_37339,N_37393);
xnor U37627 (N_37627,N_37468,N_37312);
and U37628 (N_37628,N_37257,N_37400);
nand U37629 (N_37629,N_37351,N_37321);
or U37630 (N_37630,N_37291,N_37262);
and U37631 (N_37631,N_37447,N_37358);
xor U37632 (N_37632,N_37318,N_37483);
nand U37633 (N_37633,N_37337,N_37300);
nor U37634 (N_37634,N_37324,N_37307);
and U37635 (N_37635,N_37486,N_37476);
nand U37636 (N_37636,N_37457,N_37344);
xnor U37637 (N_37637,N_37338,N_37268);
or U37638 (N_37638,N_37309,N_37308);
and U37639 (N_37639,N_37312,N_37333);
nand U37640 (N_37640,N_37322,N_37454);
nor U37641 (N_37641,N_37404,N_37458);
and U37642 (N_37642,N_37343,N_37332);
and U37643 (N_37643,N_37399,N_37490);
nand U37644 (N_37644,N_37462,N_37290);
or U37645 (N_37645,N_37455,N_37499);
or U37646 (N_37646,N_37335,N_37381);
nor U37647 (N_37647,N_37353,N_37496);
and U37648 (N_37648,N_37388,N_37441);
nand U37649 (N_37649,N_37322,N_37326);
nand U37650 (N_37650,N_37351,N_37405);
and U37651 (N_37651,N_37423,N_37311);
nand U37652 (N_37652,N_37403,N_37472);
and U37653 (N_37653,N_37331,N_37295);
or U37654 (N_37654,N_37250,N_37267);
nand U37655 (N_37655,N_37419,N_37312);
nor U37656 (N_37656,N_37480,N_37389);
or U37657 (N_37657,N_37411,N_37391);
nor U37658 (N_37658,N_37309,N_37259);
nor U37659 (N_37659,N_37281,N_37254);
and U37660 (N_37660,N_37342,N_37409);
or U37661 (N_37661,N_37364,N_37486);
xnor U37662 (N_37662,N_37483,N_37251);
or U37663 (N_37663,N_37358,N_37258);
xor U37664 (N_37664,N_37483,N_37368);
nor U37665 (N_37665,N_37382,N_37322);
nand U37666 (N_37666,N_37497,N_37391);
xnor U37667 (N_37667,N_37316,N_37395);
xor U37668 (N_37668,N_37309,N_37470);
xor U37669 (N_37669,N_37452,N_37384);
and U37670 (N_37670,N_37345,N_37311);
nand U37671 (N_37671,N_37463,N_37258);
or U37672 (N_37672,N_37493,N_37471);
nor U37673 (N_37673,N_37282,N_37321);
nor U37674 (N_37674,N_37409,N_37412);
or U37675 (N_37675,N_37255,N_37279);
xor U37676 (N_37676,N_37496,N_37406);
nor U37677 (N_37677,N_37351,N_37402);
xnor U37678 (N_37678,N_37404,N_37471);
nand U37679 (N_37679,N_37466,N_37409);
xor U37680 (N_37680,N_37298,N_37318);
or U37681 (N_37681,N_37259,N_37399);
nand U37682 (N_37682,N_37398,N_37388);
and U37683 (N_37683,N_37265,N_37487);
and U37684 (N_37684,N_37288,N_37265);
nand U37685 (N_37685,N_37319,N_37263);
or U37686 (N_37686,N_37448,N_37420);
nand U37687 (N_37687,N_37414,N_37306);
or U37688 (N_37688,N_37465,N_37279);
or U37689 (N_37689,N_37260,N_37488);
and U37690 (N_37690,N_37314,N_37305);
nand U37691 (N_37691,N_37287,N_37300);
or U37692 (N_37692,N_37400,N_37334);
xor U37693 (N_37693,N_37282,N_37471);
and U37694 (N_37694,N_37427,N_37251);
nor U37695 (N_37695,N_37311,N_37286);
xor U37696 (N_37696,N_37418,N_37403);
nor U37697 (N_37697,N_37392,N_37361);
xor U37698 (N_37698,N_37396,N_37301);
nor U37699 (N_37699,N_37274,N_37486);
and U37700 (N_37700,N_37300,N_37259);
xor U37701 (N_37701,N_37353,N_37391);
nand U37702 (N_37702,N_37370,N_37484);
or U37703 (N_37703,N_37310,N_37424);
nor U37704 (N_37704,N_37409,N_37289);
or U37705 (N_37705,N_37264,N_37365);
or U37706 (N_37706,N_37345,N_37299);
nor U37707 (N_37707,N_37380,N_37424);
nor U37708 (N_37708,N_37371,N_37437);
and U37709 (N_37709,N_37400,N_37391);
nand U37710 (N_37710,N_37376,N_37424);
and U37711 (N_37711,N_37409,N_37290);
and U37712 (N_37712,N_37314,N_37494);
or U37713 (N_37713,N_37459,N_37489);
nand U37714 (N_37714,N_37337,N_37448);
nor U37715 (N_37715,N_37351,N_37288);
xor U37716 (N_37716,N_37296,N_37388);
and U37717 (N_37717,N_37423,N_37271);
or U37718 (N_37718,N_37428,N_37380);
or U37719 (N_37719,N_37446,N_37365);
nand U37720 (N_37720,N_37486,N_37392);
nand U37721 (N_37721,N_37495,N_37415);
nand U37722 (N_37722,N_37315,N_37359);
nand U37723 (N_37723,N_37250,N_37351);
or U37724 (N_37724,N_37410,N_37282);
nand U37725 (N_37725,N_37439,N_37311);
xnor U37726 (N_37726,N_37288,N_37403);
nor U37727 (N_37727,N_37333,N_37363);
and U37728 (N_37728,N_37335,N_37443);
nand U37729 (N_37729,N_37372,N_37340);
and U37730 (N_37730,N_37330,N_37406);
nand U37731 (N_37731,N_37286,N_37485);
or U37732 (N_37732,N_37330,N_37298);
xor U37733 (N_37733,N_37340,N_37478);
nor U37734 (N_37734,N_37341,N_37328);
and U37735 (N_37735,N_37305,N_37302);
or U37736 (N_37736,N_37280,N_37356);
and U37737 (N_37737,N_37376,N_37309);
and U37738 (N_37738,N_37482,N_37330);
and U37739 (N_37739,N_37418,N_37381);
nand U37740 (N_37740,N_37276,N_37407);
nand U37741 (N_37741,N_37295,N_37361);
xor U37742 (N_37742,N_37398,N_37319);
nand U37743 (N_37743,N_37377,N_37445);
and U37744 (N_37744,N_37347,N_37457);
xor U37745 (N_37745,N_37468,N_37307);
or U37746 (N_37746,N_37463,N_37290);
and U37747 (N_37747,N_37279,N_37433);
nor U37748 (N_37748,N_37353,N_37371);
nor U37749 (N_37749,N_37358,N_37468);
or U37750 (N_37750,N_37552,N_37582);
nor U37751 (N_37751,N_37671,N_37594);
or U37752 (N_37752,N_37507,N_37567);
nor U37753 (N_37753,N_37631,N_37731);
and U37754 (N_37754,N_37646,N_37626);
nand U37755 (N_37755,N_37571,N_37585);
nand U37756 (N_37756,N_37575,N_37559);
and U37757 (N_37757,N_37737,N_37636);
nor U37758 (N_37758,N_37612,N_37655);
nor U37759 (N_37759,N_37650,N_37639);
xnor U37760 (N_37760,N_37709,N_37659);
or U37761 (N_37761,N_37729,N_37697);
xnor U37762 (N_37762,N_37510,N_37668);
nand U37763 (N_37763,N_37657,N_37532);
nor U37764 (N_37764,N_37521,N_37537);
nand U37765 (N_37765,N_37747,N_37734);
or U37766 (N_37766,N_37564,N_37610);
nand U37767 (N_37767,N_37554,N_37678);
nand U37768 (N_37768,N_37540,N_37719);
nand U37769 (N_37769,N_37677,N_37550);
and U37770 (N_37770,N_37728,N_37568);
nor U37771 (N_37771,N_37539,N_37503);
nor U37772 (N_37772,N_37563,N_37581);
or U37773 (N_37773,N_37711,N_37613);
and U37774 (N_37774,N_37705,N_37529);
nand U37775 (N_37775,N_37538,N_37635);
xor U37776 (N_37776,N_37525,N_37608);
xor U37777 (N_37777,N_37722,N_37530);
nand U37778 (N_37778,N_37624,N_37666);
nand U37779 (N_37779,N_37716,N_37640);
nor U37780 (N_37780,N_37735,N_37604);
or U37781 (N_37781,N_37674,N_37620);
and U37782 (N_37782,N_37725,N_37528);
and U37783 (N_37783,N_37645,N_37717);
nand U37784 (N_37784,N_37694,N_37648);
and U37785 (N_37785,N_37616,N_37744);
or U37786 (N_37786,N_37553,N_37500);
xnor U37787 (N_37787,N_37549,N_37609);
xnor U37788 (N_37788,N_37685,N_37629);
and U37789 (N_37789,N_37634,N_37557);
xnor U37790 (N_37790,N_37593,N_37720);
and U37791 (N_37791,N_37733,N_37508);
and U37792 (N_37792,N_37504,N_37546);
xnor U37793 (N_37793,N_37543,N_37606);
xor U37794 (N_37794,N_37618,N_37672);
and U37795 (N_37795,N_37533,N_37623);
nand U37796 (N_37796,N_37627,N_37625);
nand U37797 (N_37797,N_37587,N_37562);
nand U37798 (N_37798,N_37732,N_37601);
or U37799 (N_37799,N_37520,N_37597);
xnor U37800 (N_37800,N_37617,N_37658);
nor U37801 (N_37801,N_37661,N_37622);
and U37802 (N_37802,N_37699,N_37580);
nor U37803 (N_37803,N_37673,N_37748);
and U37804 (N_37804,N_37715,N_37718);
and U37805 (N_37805,N_37565,N_37577);
nand U37806 (N_37806,N_37542,N_37545);
or U37807 (N_37807,N_37654,N_37664);
and U37808 (N_37808,N_37517,N_37534);
and U37809 (N_37809,N_37607,N_37667);
or U37810 (N_37810,N_37547,N_37619);
and U37811 (N_37811,N_37637,N_37535);
nor U37812 (N_37812,N_37665,N_37641);
nand U37813 (N_37813,N_37512,N_37633);
nor U37814 (N_37814,N_37741,N_37724);
nand U37815 (N_37815,N_37727,N_37700);
nor U37816 (N_37816,N_37643,N_37558);
xor U37817 (N_37817,N_37515,N_37586);
or U37818 (N_37818,N_37742,N_37516);
nand U37819 (N_37819,N_37522,N_37736);
nand U37820 (N_37820,N_37638,N_37614);
or U37821 (N_37821,N_37573,N_37588);
nor U37822 (N_37822,N_37745,N_37501);
and U37823 (N_37823,N_37688,N_37703);
or U37824 (N_37824,N_37739,N_37502);
nor U37825 (N_37825,N_37684,N_37642);
nand U37826 (N_37826,N_37570,N_37670);
nand U37827 (N_37827,N_37591,N_37698);
nand U37828 (N_37828,N_37656,N_37579);
nor U37829 (N_37829,N_37713,N_37696);
nand U37830 (N_37830,N_37721,N_37605);
and U37831 (N_37831,N_37511,N_37592);
and U37832 (N_37832,N_37598,N_37527);
xnor U37833 (N_37833,N_37544,N_37669);
nand U37834 (N_37834,N_37574,N_37560);
or U37835 (N_37835,N_37676,N_37555);
nand U37836 (N_37836,N_37682,N_37583);
and U37837 (N_37837,N_37509,N_37519);
nor U37838 (N_37838,N_37536,N_37590);
and U37839 (N_37839,N_37749,N_37706);
or U37840 (N_37840,N_37746,N_37589);
and U37841 (N_37841,N_37518,N_37686);
nor U37842 (N_37842,N_37691,N_37651);
nand U37843 (N_37843,N_37576,N_37695);
nor U37844 (N_37844,N_37514,N_37690);
or U37845 (N_37845,N_37660,N_37708);
nand U37846 (N_37846,N_37740,N_37714);
xnor U37847 (N_37847,N_37584,N_37566);
and U37848 (N_37848,N_37738,N_37743);
and U37849 (N_37849,N_37730,N_37702);
nand U37850 (N_37850,N_37523,N_37596);
xnor U37851 (N_37851,N_37541,N_37561);
nor U37852 (N_37852,N_37663,N_37611);
nor U37853 (N_37853,N_37707,N_37603);
xnor U37854 (N_37854,N_37578,N_37726);
and U37855 (N_37855,N_37595,N_37647);
nand U37856 (N_37856,N_37687,N_37615);
or U37857 (N_37857,N_37652,N_37569);
or U37858 (N_37858,N_37723,N_37679);
nand U37859 (N_37859,N_37710,N_37680);
or U37860 (N_37860,N_37505,N_37630);
nor U37861 (N_37861,N_37602,N_37681);
nand U37862 (N_37862,N_37556,N_37653);
or U37863 (N_37863,N_37693,N_37683);
and U37864 (N_37864,N_37551,N_37644);
nand U37865 (N_37865,N_37712,N_37513);
nand U37866 (N_37866,N_37621,N_37689);
or U37867 (N_37867,N_37599,N_37526);
nor U37868 (N_37868,N_37531,N_37628);
xor U37869 (N_37869,N_37572,N_37662);
or U37870 (N_37870,N_37548,N_37649);
or U37871 (N_37871,N_37701,N_37524);
xor U37872 (N_37872,N_37632,N_37675);
nand U37873 (N_37873,N_37600,N_37692);
nor U37874 (N_37874,N_37506,N_37704);
nor U37875 (N_37875,N_37590,N_37599);
xor U37876 (N_37876,N_37645,N_37546);
nor U37877 (N_37877,N_37741,N_37616);
xnor U37878 (N_37878,N_37596,N_37748);
nand U37879 (N_37879,N_37563,N_37621);
or U37880 (N_37880,N_37546,N_37563);
nor U37881 (N_37881,N_37589,N_37532);
or U37882 (N_37882,N_37542,N_37540);
nand U37883 (N_37883,N_37622,N_37692);
xnor U37884 (N_37884,N_37569,N_37613);
and U37885 (N_37885,N_37640,N_37555);
and U37886 (N_37886,N_37661,N_37718);
and U37887 (N_37887,N_37741,N_37565);
nand U37888 (N_37888,N_37559,N_37628);
nand U37889 (N_37889,N_37696,N_37607);
or U37890 (N_37890,N_37656,N_37545);
nor U37891 (N_37891,N_37657,N_37637);
or U37892 (N_37892,N_37549,N_37694);
nand U37893 (N_37893,N_37741,N_37593);
or U37894 (N_37894,N_37580,N_37589);
xnor U37895 (N_37895,N_37513,N_37700);
xor U37896 (N_37896,N_37571,N_37506);
and U37897 (N_37897,N_37712,N_37643);
nand U37898 (N_37898,N_37702,N_37663);
nor U37899 (N_37899,N_37622,N_37567);
and U37900 (N_37900,N_37529,N_37543);
nor U37901 (N_37901,N_37674,N_37561);
or U37902 (N_37902,N_37525,N_37721);
nand U37903 (N_37903,N_37580,N_37702);
nand U37904 (N_37904,N_37558,N_37624);
or U37905 (N_37905,N_37714,N_37546);
nand U37906 (N_37906,N_37542,N_37528);
nand U37907 (N_37907,N_37637,N_37641);
nand U37908 (N_37908,N_37739,N_37701);
and U37909 (N_37909,N_37726,N_37709);
xor U37910 (N_37910,N_37711,N_37516);
or U37911 (N_37911,N_37592,N_37596);
and U37912 (N_37912,N_37685,N_37545);
xnor U37913 (N_37913,N_37515,N_37694);
xor U37914 (N_37914,N_37557,N_37513);
xnor U37915 (N_37915,N_37667,N_37687);
xnor U37916 (N_37916,N_37569,N_37555);
nand U37917 (N_37917,N_37664,N_37617);
nand U37918 (N_37918,N_37695,N_37608);
or U37919 (N_37919,N_37536,N_37678);
xnor U37920 (N_37920,N_37560,N_37597);
xnor U37921 (N_37921,N_37634,N_37610);
nor U37922 (N_37922,N_37661,N_37613);
nor U37923 (N_37923,N_37589,N_37643);
or U37924 (N_37924,N_37537,N_37616);
nor U37925 (N_37925,N_37520,N_37595);
nor U37926 (N_37926,N_37507,N_37741);
nor U37927 (N_37927,N_37749,N_37536);
or U37928 (N_37928,N_37541,N_37646);
nand U37929 (N_37929,N_37654,N_37609);
nor U37930 (N_37930,N_37672,N_37500);
xor U37931 (N_37931,N_37677,N_37621);
or U37932 (N_37932,N_37744,N_37581);
xor U37933 (N_37933,N_37740,N_37564);
or U37934 (N_37934,N_37680,N_37737);
and U37935 (N_37935,N_37531,N_37605);
or U37936 (N_37936,N_37605,N_37517);
nand U37937 (N_37937,N_37524,N_37521);
nand U37938 (N_37938,N_37686,N_37509);
nand U37939 (N_37939,N_37505,N_37676);
or U37940 (N_37940,N_37586,N_37659);
xor U37941 (N_37941,N_37675,N_37542);
nand U37942 (N_37942,N_37630,N_37730);
xnor U37943 (N_37943,N_37733,N_37603);
or U37944 (N_37944,N_37540,N_37509);
or U37945 (N_37945,N_37740,N_37672);
nor U37946 (N_37946,N_37696,N_37566);
or U37947 (N_37947,N_37667,N_37673);
or U37948 (N_37948,N_37507,N_37564);
nor U37949 (N_37949,N_37517,N_37628);
nand U37950 (N_37950,N_37610,N_37557);
xnor U37951 (N_37951,N_37595,N_37744);
xor U37952 (N_37952,N_37676,N_37657);
nor U37953 (N_37953,N_37637,N_37561);
nor U37954 (N_37954,N_37724,N_37571);
nand U37955 (N_37955,N_37601,N_37508);
nand U37956 (N_37956,N_37599,N_37613);
and U37957 (N_37957,N_37567,N_37685);
xor U37958 (N_37958,N_37682,N_37704);
and U37959 (N_37959,N_37515,N_37619);
or U37960 (N_37960,N_37533,N_37543);
or U37961 (N_37961,N_37577,N_37515);
nand U37962 (N_37962,N_37736,N_37508);
and U37963 (N_37963,N_37696,N_37500);
nand U37964 (N_37964,N_37635,N_37681);
xor U37965 (N_37965,N_37666,N_37737);
xnor U37966 (N_37966,N_37527,N_37615);
and U37967 (N_37967,N_37561,N_37714);
nand U37968 (N_37968,N_37549,N_37666);
nor U37969 (N_37969,N_37566,N_37626);
nor U37970 (N_37970,N_37621,N_37505);
and U37971 (N_37971,N_37549,N_37641);
xnor U37972 (N_37972,N_37634,N_37613);
nand U37973 (N_37973,N_37575,N_37543);
nor U37974 (N_37974,N_37729,N_37500);
and U37975 (N_37975,N_37567,N_37602);
nor U37976 (N_37976,N_37650,N_37534);
xor U37977 (N_37977,N_37509,N_37634);
or U37978 (N_37978,N_37531,N_37670);
or U37979 (N_37979,N_37683,N_37502);
and U37980 (N_37980,N_37561,N_37746);
and U37981 (N_37981,N_37633,N_37570);
xnor U37982 (N_37982,N_37715,N_37689);
xor U37983 (N_37983,N_37529,N_37632);
nor U37984 (N_37984,N_37667,N_37612);
xor U37985 (N_37985,N_37698,N_37647);
xor U37986 (N_37986,N_37568,N_37502);
nor U37987 (N_37987,N_37648,N_37533);
and U37988 (N_37988,N_37636,N_37510);
nor U37989 (N_37989,N_37671,N_37614);
nor U37990 (N_37990,N_37600,N_37589);
and U37991 (N_37991,N_37666,N_37571);
xor U37992 (N_37992,N_37619,N_37720);
nand U37993 (N_37993,N_37741,N_37713);
or U37994 (N_37994,N_37560,N_37689);
xnor U37995 (N_37995,N_37570,N_37742);
nand U37996 (N_37996,N_37572,N_37728);
and U37997 (N_37997,N_37701,N_37546);
or U37998 (N_37998,N_37582,N_37620);
nor U37999 (N_37999,N_37617,N_37713);
nor U38000 (N_38000,N_37772,N_37803);
or U38001 (N_38001,N_37962,N_37814);
or U38002 (N_38002,N_37883,N_37931);
xnor U38003 (N_38003,N_37788,N_37840);
nand U38004 (N_38004,N_37880,N_37855);
nor U38005 (N_38005,N_37943,N_37783);
and U38006 (N_38006,N_37892,N_37971);
xnor U38007 (N_38007,N_37837,N_37887);
and U38008 (N_38008,N_37758,N_37928);
and U38009 (N_38009,N_37779,N_37789);
nand U38010 (N_38010,N_37947,N_37827);
xnor U38011 (N_38011,N_37897,N_37774);
xnor U38012 (N_38012,N_37974,N_37938);
xor U38013 (N_38013,N_37977,N_37912);
nand U38014 (N_38014,N_37843,N_37852);
nand U38015 (N_38015,N_37805,N_37961);
xnor U38016 (N_38016,N_37822,N_37982);
xnor U38017 (N_38017,N_37771,N_37754);
xor U38018 (N_38018,N_37750,N_37829);
or U38019 (N_38019,N_37957,N_37808);
xnor U38020 (N_38020,N_37800,N_37963);
nor U38021 (N_38021,N_37867,N_37879);
nand U38022 (N_38022,N_37874,N_37809);
xnor U38023 (N_38023,N_37911,N_37818);
or U38024 (N_38024,N_37775,N_37921);
and U38025 (N_38025,N_37770,N_37756);
nor U38026 (N_38026,N_37761,N_37993);
and U38027 (N_38027,N_37815,N_37953);
nor U38028 (N_38028,N_37752,N_37759);
or U38029 (N_38029,N_37807,N_37866);
or U38030 (N_38030,N_37776,N_37960);
or U38031 (N_38031,N_37755,N_37965);
and U38032 (N_38032,N_37834,N_37841);
nand U38033 (N_38033,N_37919,N_37766);
xnor U38034 (N_38034,N_37794,N_37985);
or U38035 (N_38035,N_37869,N_37828);
and U38036 (N_38036,N_37923,N_37877);
xnor U38037 (N_38037,N_37872,N_37966);
nor U38038 (N_38038,N_37915,N_37976);
nor U38039 (N_38039,N_37904,N_37973);
and U38040 (N_38040,N_37784,N_37933);
or U38041 (N_38041,N_37991,N_37995);
nor U38042 (N_38042,N_37764,N_37777);
nor U38043 (N_38043,N_37948,N_37790);
and U38044 (N_38044,N_37935,N_37835);
or U38045 (N_38045,N_37782,N_37964);
and U38046 (N_38046,N_37819,N_37916);
nor U38047 (N_38047,N_37884,N_37981);
and U38048 (N_38048,N_37988,N_37955);
nor U38049 (N_38049,N_37941,N_37786);
xnor U38050 (N_38050,N_37959,N_37894);
or U38051 (N_38051,N_37804,N_37831);
or U38052 (N_38052,N_37944,N_37860);
and U38053 (N_38053,N_37801,N_37856);
nand U38054 (N_38054,N_37757,N_37785);
or U38055 (N_38055,N_37773,N_37889);
nand U38056 (N_38056,N_37848,N_37929);
and U38057 (N_38057,N_37940,N_37954);
nor U38058 (N_38058,N_37845,N_37906);
nand U38059 (N_38059,N_37996,N_37997);
nor U38060 (N_38060,N_37876,N_37821);
nand U38061 (N_38061,N_37796,N_37909);
and U38062 (N_38062,N_37795,N_37968);
xnor U38063 (N_38063,N_37825,N_37908);
nor U38064 (N_38064,N_37989,N_37842);
nand U38065 (N_38065,N_37905,N_37768);
nand U38066 (N_38066,N_37868,N_37914);
nor U38067 (N_38067,N_37844,N_37990);
and U38068 (N_38068,N_37824,N_37763);
and U38069 (N_38069,N_37830,N_37760);
and U38070 (N_38070,N_37980,N_37924);
nand U38071 (N_38071,N_37813,N_37817);
nand U38072 (N_38072,N_37875,N_37994);
and U38073 (N_38073,N_37922,N_37970);
xor U38074 (N_38074,N_37802,N_37799);
and U38075 (N_38075,N_37946,N_37793);
and U38076 (N_38076,N_37992,N_37896);
or U38077 (N_38077,N_37901,N_37893);
nor U38078 (N_38078,N_37895,N_37833);
xor U38079 (N_38079,N_37853,N_37891);
or U38080 (N_38080,N_37811,N_37885);
nor U38081 (N_38081,N_37792,N_37797);
nor U38082 (N_38082,N_37969,N_37958);
and U38083 (N_38083,N_37987,N_37816);
or U38084 (N_38084,N_37956,N_37900);
nand U38085 (N_38085,N_37886,N_37798);
or U38086 (N_38086,N_37937,N_37863);
or U38087 (N_38087,N_37927,N_37975);
and U38088 (N_38088,N_37846,N_37820);
nor U38089 (N_38089,N_37949,N_37862);
and U38090 (N_38090,N_37890,N_37832);
and U38091 (N_38091,N_37918,N_37861);
nand U38092 (N_38092,N_37913,N_37945);
nand U38093 (N_38093,N_37870,N_37926);
or U38094 (N_38094,N_37787,N_37812);
and U38095 (N_38095,N_37823,N_37983);
nor U38096 (N_38096,N_37972,N_37942);
nand U38097 (N_38097,N_37850,N_37951);
nand U38098 (N_38098,N_37979,N_37780);
and U38099 (N_38099,N_37936,N_37838);
nor U38100 (N_38100,N_37903,N_37881);
xor U38101 (N_38101,N_37986,N_37920);
nand U38102 (N_38102,N_37847,N_37865);
nor U38103 (N_38103,N_37769,N_37902);
or U38104 (N_38104,N_37999,N_37934);
nor U38105 (N_38105,N_37854,N_37888);
xnor U38106 (N_38106,N_37778,N_37858);
or U38107 (N_38107,N_37864,N_37925);
or U38108 (N_38108,N_37873,N_37907);
and U38109 (N_38109,N_37836,N_37810);
and U38110 (N_38110,N_37984,N_37762);
nor U38111 (N_38111,N_37878,N_37917);
or U38112 (N_38112,N_37753,N_37978);
or U38113 (N_38113,N_37851,N_37882);
xnor U38114 (N_38114,N_37998,N_37899);
or U38115 (N_38115,N_37871,N_37898);
or U38116 (N_38116,N_37939,N_37791);
nand U38117 (N_38117,N_37967,N_37826);
and U38118 (N_38118,N_37806,N_37952);
and U38119 (N_38119,N_37910,N_37767);
nand U38120 (N_38120,N_37859,N_37849);
nor U38121 (N_38121,N_37930,N_37932);
and U38122 (N_38122,N_37751,N_37857);
nand U38123 (N_38123,N_37765,N_37950);
nor U38124 (N_38124,N_37839,N_37781);
and U38125 (N_38125,N_37893,N_37862);
or U38126 (N_38126,N_37882,N_37842);
and U38127 (N_38127,N_37908,N_37795);
or U38128 (N_38128,N_37989,N_37907);
nand U38129 (N_38129,N_37813,N_37785);
xnor U38130 (N_38130,N_37787,N_37990);
nor U38131 (N_38131,N_37941,N_37784);
nand U38132 (N_38132,N_37852,N_37957);
or U38133 (N_38133,N_37789,N_37772);
nand U38134 (N_38134,N_37781,N_37855);
nor U38135 (N_38135,N_37974,N_37896);
or U38136 (N_38136,N_37988,N_37818);
or U38137 (N_38137,N_37984,N_37864);
xnor U38138 (N_38138,N_37880,N_37753);
nand U38139 (N_38139,N_37762,N_37784);
xor U38140 (N_38140,N_37828,N_37884);
or U38141 (N_38141,N_37816,N_37894);
or U38142 (N_38142,N_37930,N_37927);
and U38143 (N_38143,N_37765,N_37956);
or U38144 (N_38144,N_37971,N_37958);
and U38145 (N_38145,N_37961,N_37787);
or U38146 (N_38146,N_37834,N_37886);
xnor U38147 (N_38147,N_37784,N_37884);
or U38148 (N_38148,N_37975,N_37907);
and U38149 (N_38149,N_37849,N_37895);
or U38150 (N_38150,N_37892,N_37940);
or U38151 (N_38151,N_37830,N_37794);
or U38152 (N_38152,N_37827,N_37901);
or U38153 (N_38153,N_37948,N_37848);
or U38154 (N_38154,N_37822,N_37783);
or U38155 (N_38155,N_37785,N_37756);
xnor U38156 (N_38156,N_37826,N_37753);
nand U38157 (N_38157,N_37981,N_37860);
nand U38158 (N_38158,N_37789,N_37780);
or U38159 (N_38159,N_37915,N_37926);
nand U38160 (N_38160,N_37961,N_37949);
or U38161 (N_38161,N_37857,N_37826);
nand U38162 (N_38162,N_37753,N_37988);
nand U38163 (N_38163,N_37837,N_37772);
xor U38164 (N_38164,N_37913,N_37778);
xnor U38165 (N_38165,N_37833,N_37828);
nand U38166 (N_38166,N_37980,N_37864);
or U38167 (N_38167,N_37884,N_37973);
xnor U38168 (N_38168,N_37798,N_37917);
nand U38169 (N_38169,N_37998,N_37852);
nor U38170 (N_38170,N_37806,N_37942);
xnor U38171 (N_38171,N_37775,N_37871);
xnor U38172 (N_38172,N_37969,N_37961);
xnor U38173 (N_38173,N_37987,N_37810);
nor U38174 (N_38174,N_37893,N_37944);
nor U38175 (N_38175,N_37756,N_37947);
nor U38176 (N_38176,N_37844,N_37941);
nor U38177 (N_38177,N_37916,N_37777);
nand U38178 (N_38178,N_37932,N_37880);
or U38179 (N_38179,N_37877,N_37938);
or U38180 (N_38180,N_37986,N_37907);
and U38181 (N_38181,N_37872,N_37916);
xnor U38182 (N_38182,N_37864,N_37983);
and U38183 (N_38183,N_37821,N_37967);
and U38184 (N_38184,N_37895,N_37904);
xor U38185 (N_38185,N_37750,N_37773);
nor U38186 (N_38186,N_37891,N_37914);
nand U38187 (N_38187,N_37876,N_37909);
xor U38188 (N_38188,N_37975,N_37991);
nor U38189 (N_38189,N_37922,N_37953);
and U38190 (N_38190,N_37834,N_37843);
or U38191 (N_38191,N_37912,N_37901);
nor U38192 (N_38192,N_37884,N_37999);
or U38193 (N_38193,N_37813,N_37951);
and U38194 (N_38194,N_37949,N_37795);
xor U38195 (N_38195,N_37964,N_37773);
or U38196 (N_38196,N_37984,N_37971);
and U38197 (N_38197,N_37982,N_37802);
and U38198 (N_38198,N_37997,N_37873);
and U38199 (N_38199,N_37929,N_37755);
nand U38200 (N_38200,N_37983,N_37965);
xnor U38201 (N_38201,N_37885,N_37877);
nor U38202 (N_38202,N_37879,N_37821);
nand U38203 (N_38203,N_37857,N_37911);
and U38204 (N_38204,N_37970,N_37981);
nor U38205 (N_38205,N_37783,N_37848);
and U38206 (N_38206,N_37985,N_37763);
nor U38207 (N_38207,N_37933,N_37845);
and U38208 (N_38208,N_37954,N_37962);
nand U38209 (N_38209,N_37794,N_37966);
nand U38210 (N_38210,N_37794,N_37817);
or U38211 (N_38211,N_37939,N_37920);
and U38212 (N_38212,N_37817,N_37833);
nand U38213 (N_38213,N_37785,N_37771);
nor U38214 (N_38214,N_37751,N_37971);
or U38215 (N_38215,N_37927,N_37761);
nor U38216 (N_38216,N_37986,N_37913);
nor U38217 (N_38217,N_37834,N_37952);
nand U38218 (N_38218,N_37954,N_37932);
nand U38219 (N_38219,N_37801,N_37811);
nor U38220 (N_38220,N_37941,N_37828);
nor U38221 (N_38221,N_37859,N_37831);
and U38222 (N_38222,N_37756,N_37944);
nand U38223 (N_38223,N_37928,N_37750);
or U38224 (N_38224,N_37973,N_37826);
and U38225 (N_38225,N_37928,N_37880);
or U38226 (N_38226,N_37850,N_37754);
and U38227 (N_38227,N_37940,N_37882);
or U38228 (N_38228,N_37918,N_37946);
nand U38229 (N_38229,N_37965,N_37920);
or U38230 (N_38230,N_37881,N_37816);
or U38231 (N_38231,N_37957,N_37989);
nand U38232 (N_38232,N_37989,N_37832);
and U38233 (N_38233,N_37946,N_37803);
and U38234 (N_38234,N_37844,N_37796);
nor U38235 (N_38235,N_37959,N_37801);
nor U38236 (N_38236,N_37837,N_37976);
nor U38237 (N_38237,N_37839,N_37984);
and U38238 (N_38238,N_37970,N_37881);
nor U38239 (N_38239,N_37926,N_37994);
nand U38240 (N_38240,N_37905,N_37779);
or U38241 (N_38241,N_37879,N_37974);
nand U38242 (N_38242,N_37893,N_37941);
and U38243 (N_38243,N_37844,N_37910);
or U38244 (N_38244,N_37932,N_37811);
nor U38245 (N_38245,N_37919,N_37763);
nor U38246 (N_38246,N_37944,N_37862);
nor U38247 (N_38247,N_37804,N_37888);
xnor U38248 (N_38248,N_37944,N_37802);
and U38249 (N_38249,N_37986,N_37881);
nand U38250 (N_38250,N_38076,N_38002);
nand U38251 (N_38251,N_38111,N_38227);
and U38252 (N_38252,N_38204,N_38032);
nor U38253 (N_38253,N_38126,N_38095);
nand U38254 (N_38254,N_38056,N_38011);
or U38255 (N_38255,N_38240,N_38192);
xnor U38256 (N_38256,N_38155,N_38021);
nor U38257 (N_38257,N_38096,N_38107);
xor U38258 (N_38258,N_38184,N_38067);
and U38259 (N_38259,N_38199,N_38113);
nor U38260 (N_38260,N_38087,N_38169);
nor U38261 (N_38261,N_38005,N_38085);
or U38262 (N_38262,N_38186,N_38228);
nand U38263 (N_38263,N_38180,N_38152);
nand U38264 (N_38264,N_38022,N_38048);
nor U38265 (N_38265,N_38216,N_38058);
or U38266 (N_38266,N_38018,N_38068);
or U38267 (N_38267,N_38112,N_38134);
xor U38268 (N_38268,N_38013,N_38144);
and U38269 (N_38269,N_38145,N_38066);
nor U38270 (N_38270,N_38024,N_38235);
or U38271 (N_38271,N_38000,N_38165);
xor U38272 (N_38272,N_38059,N_38229);
or U38273 (N_38273,N_38236,N_38221);
nor U38274 (N_38274,N_38247,N_38027);
nor U38275 (N_38275,N_38241,N_38166);
nor U38276 (N_38276,N_38043,N_38213);
or U38277 (N_38277,N_38123,N_38091);
and U38278 (N_38278,N_38161,N_38189);
and U38279 (N_38279,N_38139,N_38094);
nand U38280 (N_38280,N_38233,N_38162);
or U38281 (N_38281,N_38035,N_38119);
nor U38282 (N_38282,N_38146,N_38079);
xor U38283 (N_38283,N_38249,N_38200);
xor U38284 (N_38284,N_38223,N_38129);
xor U38285 (N_38285,N_38234,N_38072);
or U38286 (N_38286,N_38194,N_38177);
and U38287 (N_38287,N_38164,N_38178);
and U38288 (N_38288,N_38029,N_38054);
nand U38289 (N_38289,N_38090,N_38127);
nor U38290 (N_38290,N_38109,N_38246);
nor U38291 (N_38291,N_38010,N_38060);
xnor U38292 (N_38292,N_38201,N_38187);
nand U38293 (N_38293,N_38080,N_38209);
nor U38294 (N_38294,N_38081,N_38230);
nor U38295 (N_38295,N_38212,N_38210);
nand U38296 (N_38296,N_38219,N_38003);
or U38297 (N_38297,N_38158,N_38028);
nor U38298 (N_38298,N_38062,N_38114);
or U38299 (N_38299,N_38020,N_38041);
nor U38300 (N_38300,N_38104,N_38132);
xor U38301 (N_38301,N_38074,N_38055);
nand U38302 (N_38302,N_38245,N_38190);
nand U38303 (N_38303,N_38097,N_38049);
xnor U38304 (N_38304,N_38208,N_38140);
and U38305 (N_38305,N_38244,N_38135);
and U38306 (N_38306,N_38057,N_38042);
nand U38307 (N_38307,N_38016,N_38214);
and U38308 (N_38308,N_38007,N_38154);
nand U38309 (N_38309,N_38019,N_38105);
nor U38310 (N_38310,N_38218,N_38009);
nand U38311 (N_38311,N_38120,N_38149);
or U38312 (N_38312,N_38099,N_38093);
and U38313 (N_38313,N_38015,N_38141);
or U38314 (N_38314,N_38008,N_38038);
and U38315 (N_38315,N_38136,N_38116);
xor U38316 (N_38316,N_38086,N_38171);
nor U38317 (N_38317,N_38172,N_38051);
or U38318 (N_38318,N_38030,N_38224);
and U38319 (N_38319,N_38037,N_38121);
nand U38320 (N_38320,N_38157,N_38193);
nor U38321 (N_38321,N_38226,N_38122);
nand U38322 (N_38322,N_38118,N_38108);
and U38323 (N_38323,N_38198,N_38045);
nor U38324 (N_38324,N_38163,N_38065);
xor U38325 (N_38325,N_38168,N_38174);
or U38326 (N_38326,N_38175,N_38239);
and U38327 (N_38327,N_38222,N_38243);
xor U38328 (N_38328,N_38195,N_38117);
and U38329 (N_38329,N_38106,N_38033);
or U38330 (N_38330,N_38084,N_38064);
or U38331 (N_38331,N_38238,N_38047);
xnor U38332 (N_38332,N_38248,N_38089);
nand U38333 (N_38333,N_38046,N_38215);
nand U38334 (N_38334,N_38070,N_38205);
and U38335 (N_38335,N_38206,N_38138);
or U38336 (N_38336,N_38159,N_38156);
nor U38337 (N_38337,N_38176,N_38073);
nand U38338 (N_38338,N_38151,N_38004);
xnor U38339 (N_38339,N_38077,N_38237);
and U38340 (N_38340,N_38148,N_38052);
and U38341 (N_38341,N_38128,N_38071);
xor U38342 (N_38342,N_38207,N_38014);
and U38343 (N_38343,N_38031,N_38153);
nand U38344 (N_38344,N_38053,N_38217);
xnor U38345 (N_38345,N_38131,N_38173);
or U38346 (N_38346,N_38179,N_38088);
or U38347 (N_38347,N_38069,N_38197);
nand U38348 (N_38348,N_38098,N_38147);
nor U38349 (N_38349,N_38036,N_38050);
xor U38350 (N_38350,N_38110,N_38100);
nand U38351 (N_38351,N_38026,N_38231);
and U38352 (N_38352,N_38188,N_38040);
xor U38353 (N_38353,N_38034,N_38075);
nor U38354 (N_38354,N_38103,N_38017);
nor U38355 (N_38355,N_38130,N_38211);
nand U38356 (N_38356,N_38125,N_38167);
nand U38357 (N_38357,N_38133,N_38124);
nand U38358 (N_38358,N_38083,N_38092);
and U38359 (N_38359,N_38044,N_38061);
nand U38360 (N_38360,N_38082,N_38182);
or U38361 (N_38361,N_38220,N_38101);
and U38362 (N_38362,N_38078,N_38039);
nor U38363 (N_38363,N_38185,N_38025);
or U38364 (N_38364,N_38115,N_38006);
xnor U38365 (N_38365,N_38196,N_38170);
nor U38366 (N_38366,N_38143,N_38001);
or U38367 (N_38367,N_38202,N_38183);
or U38368 (N_38368,N_38012,N_38150);
nand U38369 (N_38369,N_38232,N_38142);
nand U38370 (N_38370,N_38063,N_38242);
xor U38371 (N_38371,N_38160,N_38191);
or U38372 (N_38372,N_38137,N_38023);
or U38373 (N_38373,N_38203,N_38181);
nor U38374 (N_38374,N_38102,N_38225);
or U38375 (N_38375,N_38080,N_38036);
and U38376 (N_38376,N_38213,N_38178);
nor U38377 (N_38377,N_38135,N_38133);
nand U38378 (N_38378,N_38233,N_38010);
nand U38379 (N_38379,N_38177,N_38220);
or U38380 (N_38380,N_38117,N_38183);
or U38381 (N_38381,N_38191,N_38017);
or U38382 (N_38382,N_38193,N_38109);
and U38383 (N_38383,N_38010,N_38011);
nor U38384 (N_38384,N_38143,N_38221);
or U38385 (N_38385,N_38070,N_38017);
or U38386 (N_38386,N_38019,N_38000);
nor U38387 (N_38387,N_38219,N_38094);
nand U38388 (N_38388,N_38192,N_38190);
and U38389 (N_38389,N_38014,N_38226);
and U38390 (N_38390,N_38068,N_38205);
xnor U38391 (N_38391,N_38083,N_38051);
nor U38392 (N_38392,N_38238,N_38249);
nor U38393 (N_38393,N_38167,N_38208);
nor U38394 (N_38394,N_38125,N_38113);
and U38395 (N_38395,N_38116,N_38076);
nor U38396 (N_38396,N_38007,N_38242);
nor U38397 (N_38397,N_38092,N_38024);
nand U38398 (N_38398,N_38020,N_38069);
and U38399 (N_38399,N_38081,N_38218);
nor U38400 (N_38400,N_38021,N_38148);
and U38401 (N_38401,N_38177,N_38225);
xor U38402 (N_38402,N_38172,N_38009);
nand U38403 (N_38403,N_38090,N_38241);
and U38404 (N_38404,N_38003,N_38026);
nor U38405 (N_38405,N_38125,N_38014);
nand U38406 (N_38406,N_38004,N_38102);
nand U38407 (N_38407,N_38039,N_38015);
and U38408 (N_38408,N_38170,N_38207);
nand U38409 (N_38409,N_38120,N_38103);
nand U38410 (N_38410,N_38191,N_38115);
nor U38411 (N_38411,N_38154,N_38180);
nand U38412 (N_38412,N_38184,N_38166);
and U38413 (N_38413,N_38158,N_38157);
and U38414 (N_38414,N_38073,N_38175);
or U38415 (N_38415,N_38242,N_38071);
nor U38416 (N_38416,N_38217,N_38223);
and U38417 (N_38417,N_38232,N_38147);
nor U38418 (N_38418,N_38154,N_38149);
xor U38419 (N_38419,N_38168,N_38214);
xnor U38420 (N_38420,N_38033,N_38074);
or U38421 (N_38421,N_38167,N_38229);
nand U38422 (N_38422,N_38119,N_38166);
or U38423 (N_38423,N_38231,N_38062);
and U38424 (N_38424,N_38126,N_38089);
nor U38425 (N_38425,N_38094,N_38171);
and U38426 (N_38426,N_38072,N_38162);
nand U38427 (N_38427,N_38047,N_38134);
or U38428 (N_38428,N_38116,N_38185);
nand U38429 (N_38429,N_38190,N_38193);
or U38430 (N_38430,N_38214,N_38155);
or U38431 (N_38431,N_38207,N_38236);
nor U38432 (N_38432,N_38240,N_38052);
nor U38433 (N_38433,N_38237,N_38068);
xor U38434 (N_38434,N_38231,N_38158);
nor U38435 (N_38435,N_38056,N_38041);
and U38436 (N_38436,N_38124,N_38128);
or U38437 (N_38437,N_38243,N_38092);
or U38438 (N_38438,N_38096,N_38053);
nand U38439 (N_38439,N_38018,N_38051);
nor U38440 (N_38440,N_38070,N_38120);
and U38441 (N_38441,N_38015,N_38153);
and U38442 (N_38442,N_38180,N_38189);
and U38443 (N_38443,N_38011,N_38177);
nor U38444 (N_38444,N_38067,N_38149);
xnor U38445 (N_38445,N_38172,N_38189);
and U38446 (N_38446,N_38020,N_38118);
or U38447 (N_38447,N_38240,N_38024);
xor U38448 (N_38448,N_38078,N_38209);
nand U38449 (N_38449,N_38093,N_38159);
xor U38450 (N_38450,N_38185,N_38245);
nand U38451 (N_38451,N_38109,N_38199);
or U38452 (N_38452,N_38025,N_38016);
xor U38453 (N_38453,N_38051,N_38187);
and U38454 (N_38454,N_38107,N_38142);
nand U38455 (N_38455,N_38128,N_38077);
and U38456 (N_38456,N_38236,N_38097);
xor U38457 (N_38457,N_38121,N_38066);
nand U38458 (N_38458,N_38158,N_38109);
nor U38459 (N_38459,N_38045,N_38112);
nor U38460 (N_38460,N_38208,N_38174);
nor U38461 (N_38461,N_38100,N_38157);
or U38462 (N_38462,N_38197,N_38070);
xnor U38463 (N_38463,N_38017,N_38129);
nand U38464 (N_38464,N_38010,N_38091);
xnor U38465 (N_38465,N_38112,N_38044);
nand U38466 (N_38466,N_38108,N_38082);
and U38467 (N_38467,N_38048,N_38185);
nor U38468 (N_38468,N_38013,N_38093);
and U38469 (N_38469,N_38219,N_38088);
nand U38470 (N_38470,N_38103,N_38104);
or U38471 (N_38471,N_38234,N_38102);
and U38472 (N_38472,N_38228,N_38009);
nor U38473 (N_38473,N_38130,N_38244);
and U38474 (N_38474,N_38080,N_38181);
xor U38475 (N_38475,N_38034,N_38008);
or U38476 (N_38476,N_38195,N_38190);
xor U38477 (N_38477,N_38218,N_38124);
nand U38478 (N_38478,N_38142,N_38044);
nor U38479 (N_38479,N_38074,N_38052);
nor U38480 (N_38480,N_38062,N_38144);
and U38481 (N_38481,N_38055,N_38183);
and U38482 (N_38482,N_38192,N_38079);
or U38483 (N_38483,N_38189,N_38156);
or U38484 (N_38484,N_38052,N_38036);
and U38485 (N_38485,N_38108,N_38192);
nor U38486 (N_38486,N_38237,N_38011);
xnor U38487 (N_38487,N_38199,N_38068);
nor U38488 (N_38488,N_38217,N_38026);
nor U38489 (N_38489,N_38077,N_38047);
and U38490 (N_38490,N_38007,N_38050);
nand U38491 (N_38491,N_38038,N_38178);
nand U38492 (N_38492,N_38018,N_38174);
nor U38493 (N_38493,N_38154,N_38163);
nor U38494 (N_38494,N_38130,N_38208);
nor U38495 (N_38495,N_38128,N_38114);
or U38496 (N_38496,N_38177,N_38059);
nor U38497 (N_38497,N_38147,N_38034);
or U38498 (N_38498,N_38210,N_38030);
nor U38499 (N_38499,N_38088,N_38178);
nor U38500 (N_38500,N_38491,N_38389);
and U38501 (N_38501,N_38306,N_38447);
and U38502 (N_38502,N_38258,N_38300);
and U38503 (N_38503,N_38251,N_38268);
xnor U38504 (N_38504,N_38302,N_38455);
nand U38505 (N_38505,N_38309,N_38462);
and U38506 (N_38506,N_38411,N_38367);
nor U38507 (N_38507,N_38274,N_38265);
xnor U38508 (N_38508,N_38341,N_38419);
and U38509 (N_38509,N_38312,N_38372);
nand U38510 (N_38510,N_38305,N_38392);
xor U38511 (N_38511,N_38488,N_38471);
or U38512 (N_38512,N_38402,N_38307);
and U38513 (N_38513,N_38476,N_38269);
and U38514 (N_38514,N_38267,N_38421);
nor U38515 (N_38515,N_38413,N_38313);
nor U38516 (N_38516,N_38428,N_38391);
xnor U38517 (N_38517,N_38423,N_38464);
or U38518 (N_38518,N_38325,N_38373);
or U38519 (N_38519,N_38452,N_38442);
or U38520 (N_38520,N_38328,N_38264);
or U38521 (N_38521,N_38396,N_38454);
xor U38522 (N_38522,N_38361,N_38427);
nand U38523 (N_38523,N_38398,N_38433);
xor U38524 (N_38524,N_38339,N_38381);
or U38525 (N_38525,N_38414,N_38422);
or U38526 (N_38526,N_38405,N_38388);
or U38527 (N_38527,N_38284,N_38352);
and U38528 (N_38528,N_38429,N_38438);
xnor U38529 (N_38529,N_38281,N_38408);
nor U38530 (N_38530,N_38382,N_38335);
nor U38531 (N_38531,N_38275,N_38271);
xor U38532 (N_38532,N_38395,N_38437);
nor U38533 (N_38533,N_38297,N_38263);
and U38534 (N_38534,N_38255,N_38420);
nor U38535 (N_38535,N_38358,N_38393);
or U38536 (N_38536,N_38278,N_38292);
xnor U38537 (N_38537,N_38282,N_38327);
nor U38538 (N_38538,N_38448,N_38470);
nand U38539 (N_38539,N_38404,N_38316);
nor U38540 (N_38540,N_38453,N_38291);
nand U38541 (N_38541,N_38477,N_38293);
or U38542 (N_38542,N_38461,N_38288);
nand U38543 (N_38543,N_38280,N_38479);
nor U38544 (N_38544,N_38322,N_38384);
nand U38545 (N_38545,N_38363,N_38348);
nor U38546 (N_38546,N_38369,N_38385);
and U38547 (N_38547,N_38468,N_38446);
and U38548 (N_38548,N_38425,N_38359);
nand U38549 (N_38549,N_38256,N_38276);
xnor U38550 (N_38550,N_38349,N_38380);
xnor U38551 (N_38551,N_38277,N_38368);
and U38552 (N_38552,N_38417,N_38336);
and U38553 (N_38553,N_38390,N_38334);
and U38554 (N_38554,N_38298,N_38406);
nand U38555 (N_38555,N_38301,N_38410);
nand U38556 (N_38556,N_38494,N_38270);
or U38557 (N_38557,N_38370,N_38492);
or U38558 (N_38558,N_38436,N_38400);
nor U38559 (N_38559,N_38387,N_38386);
nor U38560 (N_38560,N_38377,N_38456);
nand U38561 (N_38561,N_38344,N_38407);
nand U38562 (N_38562,N_38343,N_38329);
xnor U38563 (N_38563,N_38484,N_38303);
nand U38564 (N_38564,N_38469,N_38439);
nand U38565 (N_38565,N_38418,N_38371);
nand U38566 (N_38566,N_38355,N_38432);
xnor U38567 (N_38567,N_38289,N_38315);
or U38568 (N_38568,N_38250,N_38346);
nor U38569 (N_38569,N_38347,N_38486);
nor U38570 (N_38570,N_38356,N_38310);
or U38571 (N_38571,N_38330,N_38460);
and U38572 (N_38572,N_38262,N_38299);
and U38573 (N_38573,N_38483,N_38378);
nor U38574 (N_38574,N_38273,N_38357);
and U38575 (N_38575,N_38473,N_38286);
xnor U38576 (N_38576,N_38304,N_38498);
xnor U38577 (N_38577,N_38441,N_38383);
and U38578 (N_38578,N_38482,N_38365);
nor U38579 (N_38579,N_38458,N_38444);
nand U38580 (N_38580,N_38261,N_38440);
nor U38581 (N_38581,N_38253,N_38317);
and U38582 (N_38582,N_38332,N_38257);
nor U38583 (N_38583,N_38399,N_38495);
or U38584 (N_38584,N_38353,N_38333);
nor U38585 (N_38585,N_38457,N_38259);
and U38586 (N_38586,N_38287,N_38321);
and U38587 (N_38587,N_38485,N_38463);
nor U38588 (N_38588,N_38397,N_38415);
nor U38589 (N_38589,N_38449,N_38311);
nor U38590 (N_38590,N_38490,N_38295);
nand U38591 (N_38591,N_38478,N_38308);
or U38592 (N_38592,N_38416,N_38434);
xnor U38593 (N_38593,N_38472,N_38480);
or U38594 (N_38594,N_38338,N_38314);
nor U38595 (N_38595,N_38374,N_38360);
xnor U38596 (N_38596,N_38431,N_38323);
nand U38597 (N_38597,N_38324,N_38350);
or U38598 (N_38598,N_38403,N_38285);
xor U38599 (N_38599,N_38412,N_38424);
xnor U38600 (N_38600,N_38266,N_38260);
nand U38601 (N_38601,N_38451,N_38450);
nor U38602 (N_38602,N_38497,N_38354);
nand U38603 (N_38603,N_38364,N_38475);
xor U38604 (N_38604,N_38296,N_38426);
nand U38605 (N_38605,N_38319,N_38376);
and U38606 (N_38606,N_38379,N_38252);
and U38607 (N_38607,N_38342,N_38489);
nand U38608 (N_38608,N_38445,N_38394);
nand U38609 (N_38609,N_38279,N_38481);
or U38610 (N_38610,N_38326,N_38443);
nor U38611 (N_38611,N_38283,N_38487);
nor U38612 (N_38612,N_38340,N_38493);
nand U38613 (N_38613,N_38435,N_38409);
or U38614 (N_38614,N_38337,N_38430);
and U38615 (N_38615,N_38290,N_38320);
nor U38616 (N_38616,N_38366,N_38465);
or U38617 (N_38617,N_38254,N_38345);
or U38618 (N_38618,N_38467,N_38401);
nor U38619 (N_38619,N_38318,N_38294);
nand U38620 (N_38620,N_38459,N_38331);
and U38621 (N_38621,N_38351,N_38272);
nand U38622 (N_38622,N_38499,N_38466);
xor U38623 (N_38623,N_38474,N_38362);
xor U38624 (N_38624,N_38375,N_38496);
and U38625 (N_38625,N_38313,N_38484);
nand U38626 (N_38626,N_38329,N_38388);
and U38627 (N_38627,N_38261,N_38432);
or U38628 (N_38628,N_38307,N_38381);
xnor U38629 (N_38629,N_38488,N_38324);
or U38630 (N_38630,N_38268,N_38435);
and U38631 (N_38631,N_38475,N_38404);
or U38632 (N_38632,N_38292,N_38279);
or U38633 (N_38633,N_38250,N_38259);
nand U38634 (N_38634,N_38466,N_38319);
or U38635 (N_38635,N_38452,N_38344);
nand U38636 (N_38636,N_38373,N_38441);
xnor U38637 (N_38637,N_38361,N_38468);
nor U38638 (N_38638,N_38367,N_38310);
xnor U38639 (N_38639,N_38414,N_38388);
and U38640 (N_38640,N_38314,N_38428);
nor U38641 (N_38641,N_38274,N_38473);
or U38642 (N_38642,N_38283,N_38387);
nand U38643 (N_38643,N_38451,N_38414);
or U38644 (N_38644,N_38287,N_38306);
xor U38645 (N_38645,N_38423,N_38366);
nor U38646 (N_38646,N_38383,N_38440);
or U38647 (N_38647,N_38256,N_38415);
nor U38648 (N_38648,N_38382,N_38279);
xnor U38649 (N_38649,N_38292,N_38265);
nand U38650 (N_38650,N_38491,N_38256);
xor U38651 (N_38651,N_38401,N_38258);
nor U38652 (N_38652,N_38431,N_38268);
xnor U38653 (N_38653,N_38419,N_38442);
and U38654 (N_38654,N_38320,N_38380);
nor U38655 (N_38655,N_38467,N_38369);
nor U38656 (N_38656,N_38309,N_38476);
nand U38657 (N_38657,N_38311,N_38360);
or U38658 (N_38658,N_38428,N_38392);
nor U38659 (N_38659,N_38442,N_38368);
xor U38660 (N_38660,N_38352,N_38408);
and U38661 (N_38661,N_38264,N_38383);
xnor U38662 (N_38662,N_38366,N_38407);
nand U38663 (N_38663,N_38388,N_38347);
or U38664 (N_38664,N_38438,N_38287);
nor U38665 (N_38665,N_38337,N_38359);
and U38666 (N_38666,N_38403,N_38397);
or U38667 (N_38667,N_38307,N_38332);
and U38668 (N_38668,N_38295,N_38468);
nand U38669 (N_38669,N_38456,N_38275);
or U38670 (N_38670,N_38355,N_38379);
nand U38671 (N_38671,N_38256,N_38282);
or U38672 (N_38672,N_38330,N_38451);
and U38673 (N_38673,N_38386,N_38362);
or U38674 (N_38674,N_38483,N_38498);
nor U38675 (N_38675,N_38344,N_38493);
nor U38676 (N_38676,N_38451,N_38406);
and U38677 (N_38677,N_38421,N_38324);
nor U38678 (N_38678,N_38498,N_38434);
xnor U38679 (N_38679,N_38339,N_38430);
nor U38680 (N_38680,N_38475,N_38476);
nor U38681 (N_38681,N_38375,N_38459);
or U38682 (N_38682,N_38271,N_38314);
nor U38683 (N_38683,N_38358,N_38354);
and U38684 (N_38684,N_38427,N_38418);
xnor U38685 (N_38685,N_38394,N_38326);
nor U38686 (N_38686,N_38328,N_38434);
xor U38687 (N_38687,N_38326,N_38289);
or U38688 (N_38688,N_38310,N_38470);
or U38689 (N_38689,N_38408,N_38423);
nand U38690 (N_38690,N_38477,N_38499);
xnor U38691 (N_38691,N_38308,N_38452);
nor U38692 (N_38692,N_38403,N_38287);
and U38693 (N_38693,N_38344,N_38337);
xnor U38694 (N_38694,N_38498,N_38361);
nor U38695 (N_38695,N_38372,N_38396);
nor U38696 (N_38696,N_38342,N_38322);
nor U38697 (N_38697,N_38442,N_38285);
nand U38698 (N_38698,N_38320,N_38491);
and U38699 (N_38699,N_38329,N_38327);
xnor U38700 (N_38700,N_38322,N_38253);
nand U38701 (N_38701,N_38334,N_38335);
xnor U38702 (N_38702,N_38336,N_38379);
and U38703 (N_38703,N_38444,N_38398);
xnor U38704 (N_38704,N_38489,N_38494);
or U38705 (N_38705,N_38268,N_38494);
nand U38706 (N_38706,N_38438,N_38411);
and U38707 (N_38707,N_38398,N_38417);
xnor U38708 (N_38708,N_38287,N_38375);
xnor U38709 (N_38709,N_38295,N_38350);
nor U38710 (N_38710,N_38308,N_38402);
and U38711 (N_38711,N_38374,N_38333);
xnor U38712 (N_38712,N_38304,N_38495);
or U38713 (N_38713,N_38445,N_38304);
nor U38714 (N_38714,N_38329,N_38300);
and U38715 (N_38715,N_38395,N_38323);
xnor U38716 (N_38716,N_38462,N_38496);
nand U38717 (N_38717,N_38495,N_38453);
xor U38718 (N_38718,N_38385,N_38327);
nand U38719 (N_38719,N_38270,N_38422);
nor U38720 (N_38720,N_38308,N_38321);
and U38721 (N_38721,N_38432,N_38277);
or U38722 (N_38722,N_38485,N_38442);
and U38723 (N_38723,N_38487,N_38285);
or U38724 (N_38724,N_38404,N_38367);
and U38725 (N_38725,N_38370,N_38321);
and U38726 (N_38726,N_38274,N_38324);
or U38727 (N_38727,N_38379,N_38348);
or U38728 (N_38728,N_38434,N_38311);
nor U38729 (N_38729,N_38359,N_38393);
or U38730 (N_38730,N_38254,N_38495);
or U38731 (N_38731,N_38424,N_38263);
nor U38732 (N_38732,N_38307,N_38485);
xor U38733 (N_38733,N_38412,N_38445);
or U38734 (N_38734,N_38257,N_38325);
nor U38735 (N_38735,N_38420,N_38448);
and U38736 (N_38736,N_38475,N_38456);
or U38737 (N_38737,N_38444,N_38397);
or U38738 (N_38738,N_38293,N_38492);
xor U38739 (N_38739,N_38430,N_38462);
xor U38740 (N_38740,N_38286,N_38399);
xnor U38741 (N_38741,N_38267,N_38327);
nor U38742 (N_38742,N_38432,N_38325);
nor U38743 (N_38743,N_38490,N_38391);
and U38744 (N_38744,N_38405,N_38357);
or U38745 (N_38745,N_38331,N_38424);
and U38746 (N_38746,N_38490,N_38424);
and U38747 (N_38747,N_38406,N_38409);
and U38748 (N_38748,N_38363,N_38393);
and U38749 (N_38749,N_38324,N_38309);
and U38750 (N_38750,N_38684,N_38716);
or U38751 (N_38751,N_38546,N_38718);
nand U38752 (N_38752,N_38541,N_38674);
nand U38753 (N_38753,N_38722,N_38549);
xor U38754 (N_38754,N_38678,N_38730);
xor U38755 (N_38755,N_38696,N_38563);
and U38756 (N_38756,N_38590,N_38694);
or U38757 (N_38757,N_38559,N_38536);
nor U38758 (N_38758,N_38652,N_38721);
and U38759 (N_38759,N_38640,N_38616);
nand U38760 (N_38760,N_38569,N_38532);
xor U38761 (N_38761,N_38529,N_38713);
or U38762 (N_38762,N_38587,N_38598);
and U38763 (N_38763,N_38666,N_38676);
xor U38764 (N_38764,N_38518,N_38534);
and U38765 (N_38765,N_38523,N_38708);
xor U38766 (N_38766,N_38581,N_38601);
or U38767 (N_38767,N_38725,N_38733);
nor U38768 (N_38768,N_38702,N_38593);
and U38769 (N_38769,N_38649,N_38738);
nor U38770 (N_38770,N_38603,N_38726);
xnor U38771 (N_38771,N_38561,N_38527);
or U38772 (N_38772,N_38685,N_38739);
xnor U38773 (N_38773,N_38636,N_38508);
nor U38774 (N_38774,N_38642,N_38612);
and U38775 (N_38775,N_38717,N_38669);
xor U38776 (N_38776,N_38589,N_38629);
nor U38777 (N_38777,N_38633,N_38578);
nand U38778 (N_38778,N_38632,N_38740);
and U38779 (N_38779,N_38670,N_38553);
or U38780 (N_38780,N_38568,N_38657);
or U38781 (N_38781,N_38526,N_38661);
and U38782 (N_38782,N_38550,N_38552);
xor U38783 (N_38783,N_38648,N_38579);
or U38784 (N_38784,N_38659,N_38504);
nand U38785 (N_38785,N_38644,N_38606);
xnor U38786 (N_38786,N_38746,N_38608);
or U38787 (N_38787,N_38543,N_38690);
xnor U38788 (N_38788,N_38665,N_38528);
nor U38789 (N_38789,N_38591,N_38700);
and U38790 (N_38790,N_38575,N_38571);
nand U38791 (N_38791,N_38660,N_38683);
or U38792 (N_38792,N_38688,N_38663);
nand U38793 (N_38793,N_38530,N_38682);
nor U38794 (N_38794,N_38645,N_38545);
xnor U38795 (N_38795,N_38630,N_38723);
and U38796 (N_38796,N_38729,N_38654);
or U38797 (N_38797,N_38655,N_38680);
or U38798 (N_38798,N_38604,N_38662);
nor U38799 (N_38799,N_38505,N_38520);
and U38800 (N_38800,N_38677,N_38637);
nand U38801 (N_38801,N_38544,N_38748);
xor U38802 (N_38802,N_38566,N_38706);
nand U38803 (N_38803,N_38540,N_38620);
xor U38804 (N_38804,N_38744,N_38515);
xnor U38805 (N_38805,N_38679,N_38501);
nor U38806 (N_38806,N_38567,N_38576);
or U38807 (N_38807,N_38521,N_38516);
xnor U38808 (N_38808,N_38509,N_38502);
and U38809 (N_38809,N_38582,N_38638);
nand U38810 (N_38810,N_38735,N_38599);
and U38811 (N_38811,N_38562,N_38600);
nor U38812 (N_38812,N_38622,N_38728);
nor U38813 (N_38813,N_38699,N_38675);
nor U38814 (N_38814,N_38743,N_38539);
xnor U38815 (N_38815,N_38535,N_38556);
xor U38816 (N_38816,N_38709,N_38547);
or U38817 (N_38817,N_38513,N_38584);
nor U38818 (N_38818,N_38609,N_38564);
xor U38819 (N_38819,N_38719,N_38512);
nand U38820 (N_38820,N_38626,N_38511);
and U38821 (N_38821,N_38623,N_38731);
and U38822 (N_38822,N_38749,N_38691);
and U38823 (N_38823,N_38689,N_38624);
nor U38824 (N_38824,N_38586,N_38614);
or U38825 (N_38825,N_38607,N_38588);
xnor U38826 (N_38826,N_38500,N_38647);
xor U38827 (N_38827,N_38697,N_38574);
or U38828 (N_38828,N_38613,N_38577);
nor U38829 (N_38829,N_38560,N_38596);
xor U38830 (N_38830,N_38594,N_38573);
and U38831 (N_38831,N_38742,N_38707);
xor U38832 (N_38832,N_38695,N_38724);
xor U38833 (N_38833,N_38635,N_38538);
or U38834 (N_38834,N_38650,N_38595);
or U38835 (N_38835,N_38686,N_38570);
or U38836 (N_38836,N_38737,N_38610);
and U38837 (N_38837,N_38704,N_38667);
and U38838 (N_38838,N_38745,N_38664);
nand U38839 (N_38839,N_38734,N_38698);
nor U38840 (N_38840,N_38651,N_38551);
or U38841 (N_38841,N_38687,N_38557);
and U38842 (N_38842,N_38703,N_38618);
and U38843 (N_38843,N_38533,N_38542);
or U38844 (N_38844,N_38673,N_38639);
nor U38845 (N_38845,N_38517,N_38537);
and U38846 (N_38846,N_38631,N_38506);
nand U38847 (N_38847,N_38705,N_38554);
nand U38848 (N_38848,N_38592,N_38597);
xor U38849 (N_38849,N_38711,N_38732);
and U38850 (N_38850,N_38617,N_38681);
and U38851 (N_38851,N_38585,N_38628);
xnor U38852 (N_38852,N_38580,N_38611);
xor U38853 (N_38853,N_38701,N_38715);
nand U38854 (N_38854,N_38615,N_38653);
or U38855 (N_38855,N_38619,N_38602);
nand U38856 (N_38856,N_38627,N_38641);
xor U38857 (N_38857,N_38710,N_38658);
or U38858 (N_38858,N_38736,N_38741);
nor U38859 (N_38859,N_38572,N_38714);
nor U38860 (N_38860,N_38671,N_38503);
nor U38861 (N_38861,N_38747,N_38525);
nor U38862 (N_38862,N_38558,N_38672);
nor U38863 (N_38863,N_38634,N_38720);
xnor U38864 (N_38864,N_38548,N_38668);
and U38865 (N_38865,N_38522,N_38519);
nor U38866 (N_38866,N_38531,N_38621);
nand U38867 (N_38867,N_38625,N_38565);
nor U38868 (N_38868,N_38514,N_38692);
or U38869 (N_38869,N_38555,N_38712);
or U38870 (N_38870,N_38646,N_38524);
or U38871 (N_38871,N_38727,N_38643);
nand U38872 (N_38872,N_38605,N_38507);
nor U38873 (N_38873,N_38583,N_38510);
nand U38874 (N_38874,N_38656,N_38693);
and U38875 (N_38875,N_38548,N_38563);
xor U38876 (N_38876,N_38725,N_38604);
and U38877 (N_38877,N_38712,N_38516);
xor U38878 (N_38878,N_38543,N_38638);
and U38879 (N_38879,N_38553,N_38700);
and U38880 (N_38880,N_38520,N_38616);
nand U38881 (N_38881,N_38571,N_38693);
nor U38882 (N_38882,N_38544,N_38728);
xor U38883 (N_38883,N_38565,N_38544);
and U38884 (N_38884,N_38667,N_38539);
xnor U38885 (N_38885,N_38525,N_38746);
xnor U38886 (N_38886,N_38502,N_38536);
nor U38887 (N_38887,N_38665,N_38503);
or U38888 (N_38888,N_38728,N_38624);
nor U38889 (N_38889,N_38567,N_38579);
and U38890 (N_38890,N_38665,N_38535);
or U38891 (N_38891,N_38517,N_38657);
nand U38892 (N_38892,N_38522,N_38720);
or U38893 (N_38893,N_38642,N_38574);
and U38894 (N_38894,N_38737,N_38547);
xor U38895 (N_38895,N_38632,N_38589);
nand U38896 (N_38896,N_38602,N_38747);
xor U38897 (N_38897,N_38681,N_38636);
or U38898 (N_38898,N_38702,N_38560);
nor U38899 (N_38899,N_38656,N_38636);
and U38900 (N_38900,N_38590,N_38502);
xnor U38901 (N_38901,N_38744,N_38676);
and U38902 (N_38902,N_38638,N_38724);
nand U38903 (N_38903,N_38533,N_38646);
xnor U38904 (N_38904,N_38602,N_38517);
nor U38905 (N_38905,N_38544,N_38595);
xnor U38906 (N_38906,N_38725,N_38636);
nor U38907 (N_38907,N_38578,N_38694);
nand U38908 (N_38908,N_38683,N_38669);
xor U38909 (N_38909,N_38657,N_38569);
nor U38910 (N_38910,N_38557,N_38745);
nand U38911 (N_38911,N_38550,N_38555);
and U38912 (N_38912,N_38546,N_38531);
nor U38913 (N_38913,N_38618,N_38568);
xnor U38914 (N_38914,N_38661,N_38701);
xnor U38915 (N_38915,N_38643,N_38677);
xor U38916 (N_38916,N_38709,N_38665);
nand U38917 (N_38917,N_38692,N_38560);
nor U38918 (N_38918,N_38679,N_38552);
or U38919 (N_38919,N_38600,N_38715);
or U38920 (N_38920,N_38698,N_38637);
nand U38921 (N_38921,N_38517,N_38728);
nor U38922 (N_38922,N_38724,N_38636);
nand U38923 (N_38923,N_38566,N_38714);
nor U38924 (N_38924,N_38576,N_38731);
nand U38925 (N_38925,N_38547,N_38607);
nor U38926 (N_38926,N_38709,N_38570);
or U38927 (N_38927,N_38644,N_38641);
nand U38928 (N_38928,N_38520,N_38601);
or U38929 (N_38929,N_38646,N_38715);
nor U38930 (N_38930,N_38507,N_38588);
xor U38931 (N_38931,N_38700,N_38520);
or U38932 (N_38932,N_38686,N_38671);
or U38933 (N_38933,N_38686,N_38608);
nand U38934 (N_38934,N_38509,N_38592);
and U38935 (N_38935,N_38596,N_38605);
nand U38936 (N_38936,N_38574,N_38556);
nor U38937 (N_38937,N_38645,N_38735);
nand U38938 (N_38938,N_38565,N_38596);
nor U38939 (N_38939,N_38607,N_38738);
nor U38940 (N_38940,N_38632,N_38549);
nor U38941 (N_38941,N_38708,N_38623);
and U38942 (N_38942,N_38602,N_38608);
or U38943 (N_38943,N_38688,N_38735);
and U38944 (N_38944,N_38579,N_38707);
or U38945 (N_38945,N_38558,N_38702);
nor U38946 (N_38946,N_38629,N_38523);
and U38947 (N_38947,N_38539,N_38607);
xnor U38948 (N_38948,N_38560,N_38601);
nand U38949 (N_38949,N_38582,N_38597);
xor U38950 (N_38950,N_38599,N_38682);
nor U38951 (N_38951,N_38591,N_38529);
nor U38952 (N_38952,N_38680,N_38645);
nand U38953 (N_38953,N_38571,N_38611);
nor U38954 (N_38954,N_38717,N_38526);
and U38955 (N_38955,N_38602,N_38709);
and U38956 (N_38956,N_38558,N_38509);
or U38957 (N_38957,N_38651,N_38747);
xnor U38958 (N_38958,N_38749,N_38700);
xor U38959 (N_38959,N_38671,N_38585);
xor U38960 (N_38960,N_38670,N_38564);
xnor U38961 (N_38961,N_38504,N_38641);
xnor U38962 (N_38962,N_38531,N_38573);
and U38963 (N_38963,N_38505,N_38688);
nand U38964 (N_38964,N_38598,N_38707);
nand U38965 (N_38965,N_38704,N_38559);
xor U38966 (N_38966,N_38706,N_38572);
nor U38967 (N_38967,N_38666,N_38655);
and U38968 (N_38968,N_38737,N_38623);
nor U38969 (N_38969,N_38722,N_38570);
or U38970 (N_38970,N_38675,N_38583);
and U38971 (N_38971,N_38564,N_38575);
nor U38972 (N_38972,N_38609,N_38597);
nand U38973 (N_38973,N_38565,N_38664);
xnor U38974 (N_38974,N_38705,N_38642);
or U38975 (N_38975,N_38531,N_38714);
and U38976 (N_38976,N_38578,N_38550);
or U38977 (N_38977,N_38534,N_38553);
nor U38978 (N_38978,N_38722,N_38522);
or U38979 (N_38979,N_38684,N_38741);
xnor U38980 (N_38980,N_38511,N_38606);
or U38981 (N_38981,N_38589,N_38512);
nor U38982 (N_38982,N_38556,N_38724);
nor U38983 (N_38983,N_38605,N_38525);
nand U38984 (N_38984,N_38539,N_38666);
and U38985 (N_38985,N_38670,N_38658);
or U38986 (N_38986,N_38734,N_38511);
or U38987 (N_38987,N_38673,N_38602);
and U38988 (N_38988,N_38518,N_38574);
nand U38989 (N_38989,N_38640,N_38667);
xor U38990 (N_38990,N_38563,N_38555);
xor U38991 (N_38991,N_38704,N_38538);
nor U38992 (N_38992,N_38690,N_38563);
or U38993 (N_38993,N_38500,N_38640);
xnor U38994 (N_38994,N_38617,N_38724);
and U38995 (N_38995,N_38654,N_38570);
xnor U38996 (N_38996,N_38501,N_38743);
nor U38997 (N_38997,N_38667,N_38611);
nor U38998 (N_38998,N_38625,N_38748);
or U38999 (N_38999,N_38669,N_38624);
nor U39000 (N_39000,N_38786,N_38925);
xor U39001 (N_39001,N_38976,N_38836);
and U39002 (N_39002,N_38927,N_38900);
and U39003 (N_39003,N_38938,N_38959);
nor U39004 (N_39004,N_38989,N_38957);
nand U39005 (N_39005,N_38899,N_38823);
or U39006 (N_39006,N_38847,N_38956);
xnor U39007 (N_39007,N_38793,N_38854);
or U39008 (N_39008,N_38750,N_38965);
or U39009 (N_39009,N_38843,N_38851);
nor U39010 (N_39010,N_38771,N_38935);
nor U39011 (N_39011,N_38894,N_38831);
nor U39012 (N_39012,N_38890,N_38926);
nand U39013 (N_39013,N_38797,N_38895);
nand U39014 (N_39014,N_38961,N_38997);
xnor U39015 (N_39015,N_38783,N_38969);
nand U39016 (N_39016,N_38909,N_38811);
or U39017 (N_39017,N_38818,N_38868);
or U39018 (N_39018,N_38758,N_38940);
or U39019 (N_39019,N_38878,N_38782);
and U39020 (N_39020,N_38856,N_38880);
nor U39021 (N_39021,N_38807,N_38883);
or U39022 (N_39022,N_38799,N_38873);
nor U39023 (N_39023,N_38974,N_38780);
nor U39024 (N_39024,N_38845,N_38817);
nor U39025 (N_39025,N_38892,N_38784);
xor U39026 (N_39026,N_38844,N_38917);
xnor U39027 (N_39027,N_38765,N_38766);
or U39028 (N_39028,N_38752,N_38977);
xnor U39029 (N_39029,N_38955,N_38903);
xnor U39030 (N_39030,N_38970,N_38803);
or U39031 (N_39031,N_38779,N_38920);
nand U39032 (N_39032,N_38981,N_38882);
xor U39033 (N_39033,N_38833,N_38952);
nand U39034 (N_39034,N_38821,N_38924);
xnor U39035 (N_39035,N_38830,N_38958);
or U39036 (N_39036,N_38754,N_38846);
xor U39037 (N_39037,N_38824,N_38874);
xor U39038 (N_39038,N_38891,N_38808);
and U39039 (N_39039,N_38852,N_38798);
nor U39040 (N_39040,N_38893,N_38810);
and U39041 (N_39041,N_38948,N_38767);
and U39042 (N_39042,N_38763,N_38901);
and U39043 (N_39043,N_38879,N_38937);
and U39044 (N_39044,N_38964,N_38790);
and U39045 (N_39045,N_38944,N_38776);
and U39046 (N_39046,N_38864,N_38967);
nor U39047 (N_39047,N_38933,N_38910);
xor U39048 (N_39048,N_38960,N_38777);
nor U39049 (N_39049,N_38902,N_38773);
or U39050 (N_39050,N_38753,N_38772);
nand U39051 (N_39051,N_38820,N_38794);
and U39052 (N_39052,N_38966,N_38858);
or U39053 (N_39053,N_38813,N_38908);
nor U39054 (N_39054,N_38814,N_38946);
nand U39055 (N_39055,N_38881,N_38825);
and U39056 (N_39056,N_38999,N_38778);
xnor U39057 (N_39057,N_38986,N_38875);
xnor U39058 (N_39058,N_38988,N_38934);
nor U39059 (N_39059,N_38923,N_38888);
nand U39060 (N_39060,N_38889,N_38993);
and U39061 (N_39061,N_38816,N_38978);
or U39062 (N_39062,N_38787,N_38990);
or U39063 (N_39063,N_38828,N_38885);
xnor U39064 (N_39064,N_38947,N_38984);
nand U39065 (N_39065,N_38953,N_38916);
nor U39066 (N_39066,N_38857,N_38853);
and U39067 (N_39067,N_38918,N_38928);
xnor U39068 (N_39068,N_38987,N_38855);
xor U39069 (N_39069,N_38796,N_38760);
nor U39070 (N_39070,N_38781,N_38768);
xor U39071 (N_39071,N_38822,N_38809);
or U39072 (N_39072,N_38789,N_38975);
and U39073 (N_39073,N_38804,N_38982);
xor U39074 (N_39074,N_38896,N_38911);
and U39075 (N_39075,N_38842,N_38762);
nor U39076 (N_39076,N_38755,N_38905);
or U39077 (N_39077,N_38827,N_38839);
or U39078 (N_39078,N_38826,N_38764);
and U39079 (N_39079,N_38815,N_38904);
or U39080 (N_39080,N_38971,N_38862);
nand U39081 (N_39081,N_38812,N_38871);
xor U39082 (N_39082,N_38985,N_38801);
and U39083 (N_39083,N_38898,N_38921);
or U39084 (N_39084,N_38943,N_38848);
and U39085 (N_39085,N_38968,N_38941);
xnor U39086 (N_39086,N_38865,N_38991);
nor U39087 (N_39087,N_38929,N_38860);
nand U39088 (N_39088,N_38834,N_38887);
and U39089 (N_39089,N_38806,N_38867);
or U39090 (N_39090,N_38995,N_38913);
and U39091 (N_39091,N_38761,N_38876);
xor U39092 (N_39092,N_38819,N_38973);
nor U39093 (N_39093,N_38835,N_38866);
or U39094 (N_39094,N_38950,N_38954);
xor U39095 (N_39095,N_38907,N_38906);
nor U39096 (N_39096,N_38838,N_38980);
nand U39097 (N_39097,N_38930,N_38870);
nor U39098 (N_39098,N_38829,N_38942);
nand U39099 (N_39099,N_38791,N_38756);
xnor U39100 (N_39100,N_38832,N_38872);
or U39101 (N_39101,N_38962,N_38994);
or U39102 (N_39102,N_38915,N_38769);
or U39103 (N_39103,N_38996,N_38919);
nand U39104 (N_39104,N_38963,N_38785);
or U39105 (N_39105,N_38850,N_38863);
nand U39106 (N_39106,N_38945,N_38792);
xnor U39107 (N_39107,N_38979,N_38770);
xnor U39108 (N_39108,N_38869,N_38897);
or U39109 (N_39109,N_38983,N_38932);
nand U39110 (N_39110,N_38849,N_38949);
xnor U39111 (N_39111,N_38802,N_38998);
nor U39112 (N_39112,N_38884,N_38914);
or U39113 (N_39113,N_38951,N_38877);
and U39114 (N_39114,N_38775,N_38922);
and U39115 (N_39115,N_38931,N_38912);
nand U39116 (N_39116,N_38795,N_38800);
xnor U39117 (N_39117,N_38972,N_38774);
xnor U39118 (N_39118,N_38886,N_38837);
nor U39119 (N_39119,N_38939,N_38859);
and U39120 (N_39120,N_38992,N_38788);
nor U39121 (N_39121,N_38751,N_38841);
nand U39122 (N_39122,N_38936,N_38759);
nand U39123 (N_39123,N_38805,N_38861);
and U39124 (N_39124,N_38757,N_38840);
nand U39125 (N_39125,N_38814,N_38873);
and U39126 (N_39126,N_38903,N_38815);
nand U39127 (N_39127,N_38854,N_38873);
or U39128 (N_39128,N_38996,N_38865);
nor U39129 (N_39129,N_38875,N_38993);
and U39130 (N_39130,N_38918,N_38966);
nand U39131 (N_39131,N_38789,N_38911);
and U39132 (N_39132,N_38938,N_38953);
nor U39133 (N_39133,N_38949,N_38923);
xnor U39134 (N_39134,N_38784,N_38891);
nor U39135 (N_39135,N_38881,N_38810);
or U39136 (N_39136,N_38977,N_38800);
and U39137 (N_39137,N_38845,N_38875);
or U39138 (N_39138,N_38976,N_38775);
xor U39139 (N_39139,N_38784,N_38755);
nor U39140 (N_39140,N_38754,N_38885);
nor U39141 (N_39141,N_38901,N_38955);
nand U39142 (N_39142,N_38767,N_38967);
xnor U39143 (N_39143,N_38975,N_38838);
nor U39144 (N_39144,N_38941,N_38865);
or U39145 (N_39145,N_38898,N_38805);
and U39146 (N_39146,N_38782,N_38803);
and U39147 (N_39147,N_38852,N_38766);
and U39148 (N_39148,N_38868,N_38776);
or U39149 (N_39149,N_38797,N_38771);
or U39150 (N_39150,N_38807,N_38767);
nor U39151 (N_39151,N_38932,N_38844);
xor U39152 (N_39152,N_38792,N_38954);
xor U39153 (N_39153,N_38935,N_38872);
nor U39154 (N_39154,N_38986,N_38892);
nor U39155 (N_39155,N_38916,N_38854);
nand U39156 (N_39156,N_38904,N_38858);
or U39157 (N_39157,N_38998,N_38881);
nand U39158 (N_39158,N_38829,N_38793);
nand U39159 (N_39159,N_38799,N_38782);
nor U39160 (N_39160,N_38960,N_38803);
or U39161 (N_39161,N_38775,N_38764);
or U39162 (N_39162,N_38863,N_38769);
or U39163 (N_39163,N_38875,N_38987);
nor U39164 (N_39164,N_38928,N_38830);
xor U39165 (N_39165,N_38872,N_38799);
nor U39166 (N_39166,N_38784,N_38774);
and U39167 (N_39167,N_38855,N_38991);
and U39168 (N_39168,N_38823,N_38976);
and U39169 (N_39169,N_38985,N_38786);
xnor U39170 (N_39170,N_38943,N_38849);
nor U39171 (N_39171,N_38915,N_38856);
nor U39172 (N_39172,N_38909,N_38870);
nand U39173 (N_39173,N_38905,N_38819);
and U39174 (N_39174,N_38811,N_38988);
nand U39175 (N_39175,N_38892,N_38959);
nor U39176 (N_39176,N_38964,N_38994);
nand U39177 (N_39177,N_38761,N_38943);
and U39178 (N_39178,N_38894,N_38947);
nand U39179 (N_39179,N_38961,N_38772);
nand U39180 (N_39180,N_38978,N_38870);
xor U39181 (N_39181,N_38884,N_38886);
xnor U39182 (N_39182,N_38762,N_38935);
and U39183 (N_39183,N_38817,N_38996);
and U39184 (N_39184,N_38759,N_38832);
xnor U39185 (N_39185,N_38915,N_38820);
and U39186 (N_39186,N_38969,N_38825);
nor U39187 (N_39187,N_38982,N_38955);
xor U39188 (N_39188,N_38858,N_38926);
or U39189 (N_39189,N_38920,N_38994);
or U39190 (N_39190,N_38938,N_38928);
nand U39191 (N_39191,N_38815,N_38936);
xnor U39192 (N_39192,N_38803,N_38786);
nor U39193 (N_39193,N_38798,N_38841);
and U39194 (N_39194,N_38982,N_38939);
nor U39195 (N_39195,N_38901,N_38888);
nor U39196 (N_39196,N_38975,N_38825);
nor U39197 (N_39197,N_38970,N_38805);
and U39198 (N_39198,N_38933,N_38808);
nand U39199 (N_39199,N_38752,N_38907);
nor U39200 (N_39200,N_38767,N_38947);
nand U39201 (N_39201,N_38995,N_38974);
nand U39202 (N_39202,N_38756,N_38842);
or U39203 (N_39203,N_38779,N_38828);
nor U39204 (N_39204,N_38895,N_38969);
nor U39205 (N_39205,N_38774,N_38971);
or U39206 (N_39206,N_38799,N_38961);
nor U39207 (N_39207,N_38868,N_38848);
nor U39208 (N_39208,N_38985,N_38858);
nor U39209 (N_39209,N_38756,N_38755);
nor U39210 (N_39210,N_38995,N_38756);
or U39211 (N_39211,N_38894,N_38800);
and U39212 (N_39212,N_38992,N_38983);
or U39213 (N_39213,N_38886,N_38785);
and U39214 (N_39214,N_38855,N_38864);
or U39215 (N_39215,N_38857,N_38974);
or U39216 (N_39216,N_38885,N_38917);
nand U39217 (N_39217,N_38949,N_38809);
nor U39218 (N_39218,N_38823,N_38794);
nand U39219 (N_39219,N_38949,N_38881);
nor U39220 (N_39220,N_38984,N_38763);
and U39221 (N_39221,N_38776,N_38991);
and U39222 (N_39222,N_38963,N_38998);
nand U39223 (N_39223,N_38799,N_38779);
nor U39224 (N_39224,N_38845,N_38771);
or U39225 (N_39225,N_38907,N_38918);
nor U39226 (N_39226,N_38954,N_38895);
and U39227 (N_39227,N_38778,N_38794);
xor U39228 (N_39228,N_38837,N_38958);
or U39229 (N_39229,N_38918,N_38838);
xor U39230 (N_39230,N_38966,N_38947);
and U39231 (N_39231,N_38843,N_38789);
and U39232 (N_39232,N_38853,N_38997);
nand U39233 (N_39233,N_38792,N_38833);
nand U39234 (N_39234,N_38884,N_38764);
xor U39235 (N_39235,N_38874,N_38897);
and U39236 (N_39236,N_38990,N_38993);
xnor U39237 (N_39237,N_38772,N_38782);
nand U39238 (N_39238,N_38768,N_38878);
or U39239 (N_39239,N_38775,N_38865);
xnor U39240 (N_39240,N_38812,N_38757);
xor U39241 (N_39241,N_38828,N_38769);
nor U39242 (N_39242,N_38832,N_38914);
nand U39243 (N_39243,N_38751,N_38853);
or U39244 (N_39244,N_38812,N_38944);
nor U39245 (N_39245,N_38769,N_38895);
xnor U39246 (N_39246,N_38963,N_38822);
or U39247 (N_39247,N_38772,N_38886);
and U39248 (N_39248,N_38830,N_38862);
nand U39249 (N_39249,N_38827,N_38837);
nor U39250 (N_39250,N_39072,N_39036);
nor U39251 (N_39251,N_39200,N_39016);
and U39252 (N_39252,N_39037,N_39025);
xnor U39253 (N_39253,N_39160,N_39121);
nand U39254 (N_39254,N_39223,N_39229);
nand U39255 (N_39255,N_39218,N_39056);
nor U39256 (N_39256,N_39248,N_39064);
nand U39257 (N_39257,N_39051,N_39130);
nor U39258 (N_39258,N_39166,N_39133);
or U39259 (N_39259,N_39182,N_39199);
nor U39260 (N_39260,N_39006,N_39127);
or U39261 (N_39261,N_39076,N_39090);
xnor U39262 (N_39262,N_39108,N_39134);
nor U39263 (N_39263,N_39209,N_39228);
nand U39264 (N_39264,N_39118,N_39171);
and U39265 (N_39265,N_39015,N_39139);
nand U39266 (N_39266,N_39247,N_39012);
nand U39267 (N_39267,N_39152,N_39031);
xor U39268 (N_39268,N_39236,N_39120);
nand U39269 (N_39269,N_39097,N_39086);
or U39270 (N_39270,N_39143,N_39009);
and U39271 (N_39271,N_39119,N_39125);
or U39272 (N_39272,N_39181,N_39138);
or U39273 (N_39273,N_39000,N_39093);
nand U39274 (N_39274,N_39211,N_39220);
nor U39275 (N_39275,N_39089,N_39017);
or U39276 (N_39276,N_39245,N_39205);
nor U39277 (N_39277,N_39188,N_39044);
and U39278 (N_39278,N_39179,N_39193);
nand U39279 (N_39279,N_39194,N_39170);
or U39280 (N_39280,N_39176,N_39109);
nand U39281 (N_39281,N_39233,N_39238);
or U39282 (N_39282,N_39158,N_39062);
nand U39283 (N_39283,N_39135,N_39183);
and U39284 (N_39284,N_39032,N_39189);
or U39285 (N_39285,N_39007,N_39243);
nor U39286 (N_39286,N_39103,N_39107);
xor U39287 (N_39287,N_39178,N_39180);
nand U39288 (N_39288,N_39094,N_39219);
or U39289 (N_39289,N_39029,N_39234);
nor U39290 (N_39290,N_39046,N_39136);
and U39291 (N_39291,N_39147,N_39175);
nand U39292 (N_39292,N_39095,N_39048);
nor U39293 (N_39293,N_39227,N_39246);
xnor U39294 (N_39294,N_39002,N_39073);
xor U39295 (N_39295,N_39106,N_39074);
or U39296 (N_39296,N_39132,N_39244);
or U39297 (N_39297,N_39004,N_39061);
and U39298 (N_39298,N_39001,N_39126);
and U39299 (N_39299,N_39240,N_39070);
and U39300 (N_39300,N_39249,N_39225);
xnor U39301 (N_39301,N_39242,N_39163);
and U39302 (N_39302,N_39042,N_39195);
xor U39303 (N_39303,N_39156,N_39174);
or U39304 (N_39304,N_39039,N_39150);
nor U39305 (N_39305,N_39068,N_39018);
or U39306 (N_39306,N_39045,N_39060);
nand U39307 (N_39307,N_39075,N_39155);
nor U39308 (N_39308,N_39235,N_39028);
nor U39309 (N_39309,N_39112,N_39040);
or U39310 (N_39310,N_39067,N_39214);
or U39311 (N_39311,N_39208,N_39116);
nand U39312 (N_39312,N_39058,N_39052);
xor U39313 (N_39313,N_39148,N_39035);
nor U39314 (N_39314,N_39212,N_39080);
nor U39315 (N_39315,N_39047,N_39237);
nand U39316 (N_39316,N_39079,N_39085);
nor U39317 (N_39317,N_39226,N_39034);
or U39318 (N_39318,N_39167,N_39197);
xor U39319 (N_39319,N_39063,N_39038);
xor U39320 (N_39320,N_39165,N_39131);
nand U39321 (N_39321,N_39124,N_39146);
nand U39322 (N_39322,N_39099,N_39157);
nor U39323 (N_39323,N_39071,N_39210);
or U39324 (N_39324,N_39066,N_39030);
or U39325 (N_39325,N_39213,N_39154);
nor U39326 (N_39326,N_39078,N_39113);
nand U39327 (N_39327,N_39230,N_39096);
nor U39328 (N_39328,N_39123,N_39177);
or U39329 (N_39329,N_39203,N_39169);
or U39330 (N_39330,N_39008,N_39129);
nand U39331 (N_39331,N_39221,N_39151);
nor U39332 (N_39332,N_39083,N_39027);
xnor U39333 (N_39333,N_39145,N_39105);
nor U39334 (N_39334,N_39162,N_39172);
and U39335 (N_39335,N_39023,N_39010);
xor U39336 (N_39336,N_39102,N_39100);
nand U39337 (N_39337,N_39164,N_39059);
and U39338 (N_39338,N_39050,N_39114);
nor U39339 (N_39339,N_39173,N_39011);
nor U39340 (N_39340,N_39231,N_39041);
and U39341 (N_39341,N_39077,N_39019);
and U39342 (N_39342,N_39087,N_39115);
nand U39343 (N_39343,N_39239,N_39149);
xnor U39344 (N_39344,N_39224,N_39190);
and U39345 (N_39345,N_39186,N_39153);
xor U39346 (N_39346,N_39021,N_39159);
and U39347 (N_39347,N_39122,N_39003);
and U39348 (N_39348,N_39082,N_39055);
nor U39349 (N_39349,N_39207,N_39081);
xnor U39350 (N_39350,N_39092,N_39014);
nor U39351 (N_39351,N_39128,N_39191);
and U39352 (N_39352,N_39141,N_39185);
and U39353 (N_39353,N_39091,N_39140);
xor U39354 (N_39354,N_39168,N_39192);
nand U39355 (N_39355,N_39098,N_39187);
nor U39356 (N_39356,N_39144,N_39204);
nand U39357 (N_39357,N_39024,N_39215);
and U39358 (N_39358,N_39222,N_39206);
xnor U39359 (N_39359,N_39216,N_39022);
nor U39360 (N_39360,N_39057,N_39117);
nor U39361 (N_39361,N_39110,N_39184);
nor U39362 (N_39362,N_39013,N_39196);
or U39363 (N_39363,N_39033,N_39053);
or U39364 (N_39364,N_39202,N_39137);
xnor U39365 (N_39365,N_39142,N_39065);
nand U39366 (N_39366,N_39217,N_39084);
xor U39367 (N_39367,N_39198,N_39005);
nand U39368 (N_39368,N_39161,N_39104);
nand U39369 (N_39369,N_39020,N_39111);
nand U39370 (N_39370,N_39026,N_39088);
xor U39371 (N_39371,N_39069,N_39101);
xnor U39372 (N_39372,N_39201,N_39241);
xor U39373 (N_39373,N_39049,N_39232);
xor U39374 (N_39374,N_39054,N_39043);
nand U39375 (N_39375,N_39131,N_39088);
xnor U39376 (N_39376,N_39109,N_39112);
xor U39377 (N_39377,N_39082,N_39008);
xor U39378 (N_39378,N_39019,N_39149);
or U39379 (N_39379,N_39071,N_39245);
nand U39380 (N_39380,N_39167,N_39033);
and U39381 (N_39381,N_39053,N_39076);
nor U39382 (N_39382,N_39182,N_39039);
xor U39383 (N_39383,N_39073,N_39233);
nor U39384 (N_39384,N_39149,N_39117);
xor U39385 (N_39385,N_39026,N_39027);
or U39386 (N_39386,N_39101,N_39104);
xor U39387 (N_39387,N_39049,N_39140);
nand U39388 (N_39388,N_39248,N_39058);
and U39389 (N_39389,N_39069,N_39173);
and U39390 (N_39390,N_39193,N_39028);
and U39391 (N_39391,N_39217,N_39181);
and U39392 (N_39392,N_39074,N_39003);
xnor U39393 (N_39393,N_39017,N_39056);
xnor U39394 (N_39394,N_39162,N_39147);
and U39395 (N_39395,N_39124,N_39165);
nand U39396 (N_39396,N_39198,N_39218);
and U39397 (N_39397,N_39247,N_39204);
xor U39398 (N_39398,N_39102,N_39209);
xnor U39399 (N_39399,N_39183,N_39170);
nand U39400 (N_39400,N_39076,N_39110);
and U39401 (N_39401,N_39078,N_39007);
nand U39402 (N_39402,N_39149,N_39130);
and U39403 (N_39403,N_39074,N_39015);
nor U39404 (N_39404,N_39022,N_39209);
and U39405 (N_39405,N_39246,N_39057);
and U39406 (N_39406,N_39214,N_39123);
or U39407 (N_39407,N_39238,N_39093);
xnor U39408 (N_39408,N_39169,N_39095);
xnor U39409 (N_39409,N_39227,N_39138);
or U39410 (N_39410,N_39100,N_39042);
xnor U39411 (N_39411,N_39229,N_39076);
nor U39412 (N_39412,N_39103,N_39055);
or U39413 (N_39413,N_39084,N_39095);
nand U39414 (N_39414,N_39122,N_39180);
nand U39415 (N_39415,N_39077,N_39111);
and U39416 (N_39416,N_39240,N_39146);
nor U39417 (N_39417,N_39036,N_39184);
nand U39418 (N_39418,N_39099,N_39040);
or U39419 (N_39419,N_39052,N_39094);
or U39420 (N_39420,N_39072,N_39218);
or U39421 (N_39421,N_39087,N_39044);
or U39422 (N_39422,N_39008,N_39184);
nand U39423 (N_39423,N_39055,N_39156);
or U39424 (N_39424,N_39044,N_39216);
or U39425 (N_39425,N_39041,N_39006);
nand U39426 (N_39426,N_39115,N_39099);
nor U39427 (N_39427,N_39082,N_39113);
or U39428 (N_39428,N_39057,N_39027);
and U39429 (N_39429,N_39193,N_39065);
nor U39430 (N_39430,N_39219,N_39016);
nor U39431 (N_39431,N_39056,N_39196);
nor U39432 (N_39432,N_39238,N_39146);
or U39433 (N_39433,N_39000,N_39137);
and U39434 (N_39434,N_39050,N_39203);
nor U39435 (N_39435,N_39090,N_39159);
and U39436 (N_39436,N_39221,N_39020);
or U39437 (N_39437,N_39137,N_39243);
nor U39438 (N_39438,N_39086,N_39013);
or U39439 (N_39439,N_39063,N_39144);
and U39440 (N_39440,N_39139,N_39244);
nor U39441 (N_39441,N_39225,N_39011);
and U39442 (N_39442,N_39179,N_39165);
and U39443 (N_39443,N_39221,N_39239);
and U39444 (N_39444,N_39100,N_39226);
and U39445 (N_39445,N_39229,N_39165);
and U39446 (N_39446,N_39085,N_39063);
nand U39447 (N_39447,N_39122,N_39067);
nor U39448 (N_39448,N_39193,N_39228);
xnor U39449 (N_39449,N_39018,N_39103);
nor U39450 (N_39450,N_39100,N_39216);
nand U39451 (N_39451,N_39098,N_39245);
and U39452 (N_39452,N_39238,N_39199);
xor U39453 (N_39453,N_39203,N_39076);
and U39454 (N_39454,N_39052,N_39141);
nor U39455 (N_39455,N_39195,N_39166);
xnor U39456 (N_39456,N_39154,N_39145);
nor U39457 (N_39457,N_39046,N_39019);
nor U39458 (N_39458,N_39207,N_39224);
and U39459 (N_39459,N_39161,N_39231);
nand U39460 (N_39460,N_39043,N_39225);
nand U39461 (N_39461,N_39157,N_39001);
xnor U39462 (N_39462,N_39090,N_39197);
or U39463 (N_39463,N_39019,N_39028);
and U39464 (N_39464,N_39206,N_39136);
nand U39465 (N_39465,N_39206,N_39135);
nand U39466 (N_39466,N_39097,N_39114);
nand U39467 (N_39467,N_39209,N_39067);
nor U39468 (N_39468,N_39006,N_39208);
nor U39469 (N_39469,N_39097,N_39106);
nor U39470 (N_39470,N_39081,N_39147);
xor U39471 (N_39471,N_39113,N_39159);
or U39472 (N_39472,N_39015,N_39178);
or U39473 (N_39473,N_39070,N_39103);
and U39474 (N_39474,N_39069,N_39142);
nand U39475 (N_39475,N_39200,N_39001);
or U39476 (N_39476,N_39156,N_39124);
and U39477 (N_39477,N_39159,N_39135);
xnor U39478 (N_39478,N_39034,N_39000);
nor U39479 (N_39479,N_39000,N_39191);
or U39480 (N_39480,N_39059,N_39202);
and U39481 (N_39481,N_39090,N_39222);
nor U39482 (N_39482,N_39066,N_39112);
and U39483 (N_39483,N_39070,N_39040);
nor U39484 (N_39484,N_39215,N_39061);
and U39485 (N_39485,N_39242,N_39077);
or U39486 (N_39486,N_39200,N_39147);
and U39487 (N_39487,N_39220,N_39209);
nor U39488 (N_39488,N_39052,N_39145);
and U39489 (N_39489,N_39194,N_39067);
nand U39490 (N_39490,N_39225,N_39012);
nor U39491 (N_39491,N_39086,N_39159);
and U39492 (N_39492,N_39205,N_39149);
nor U39493 (N_39493,N_39028,N_39156);
or U39494 (N_39494,N_39186,N_39074);
xnor U39495 (N_39495,N_39013,N_39131);
xnor U39496 (N_39496,N_39107,N_39161);
nor U39497 (N_39497,N_39034,N_39216);
xor U39498 (N_39498,N_39180,N_39019);
xor U39499 (N_39499,N_39073,N_39232);
xor U39500 (N_39500,N_39402,N_39282);
or U39501 (N_39501,N_39256,N_39393);
xor U39502 (N_39502,N_39499,N_39262);
nor U39503 (N_39503,N_39404,N_39492);
nand U39504 (N_39504,N_39355,N_39412);
xor U39505 (N_39505,N_39275,N_39306);
and U39506 (N_39506,N_39297,N_39364);
nor U39507 (N_39507,N_39263,N_39455);
or U39508 (N_39508,N_39386,N_39448);
nor U39509 (N_39509,N_39477,N_39330);
or U39510 (N_39510,N_39435,N_39493);
and U39511 (N_39511,N_39349,N_39445);
or U39512 (N_39512,N_39385,N_39365);
xnor U39513 (N_39513,N_39315,N_39298);
xnor U39514 (N_39514,N_39254,N_39406);
nor U39515 (N_39515,N_39328,N_39481);
nand U39516 (N_39516,N_39257,N_39361);
nand U39517 (N_39517,N_39373,N_39292);
nor U39518 (N_39518,N_39442,N_39483);
nand U39519 (N_39519,N_39416,N_39486);
or U39520 (N_39520,N_39490,N_39382);
nor U39521 (N_39521,N_39434,N_39265);
and U39522 (N_39522,N_39398,N_39400);
and U39523 (N_39523,N_39429,N_39459);
or U39524 (N_39524,N_39321,N_39437);
nor U39525 (N_39525,N_39342,N_39424);
or U39526 (N_39526,N_39320,N_39383);
xnor U39527 (N_39527,N_39409,N_39329);
or U39528 (N_39528,N_39339,N_39475);
and U39529 (N_39529,N_39472,N_39418);
nor U39530 (N_39530,N_39381,N_39305);
or U39531 (N_39531,N_39301,N_39428);
xnor U39532 (N_39532,N_39359,N_39423);
nor U39533 (N_39533,N_39266,N_39425);
nor U39534 (N_39534,N_39344,N_39449);
and U39535 (N_39535,N_39443,N_39452);
or U39536 (N_39536,N_39388,N_39269);
and U39537 (N_39537,N_39303,N_39470);
nand U39538 (N_39538,N_39347,N_39458);
and U39539 (N_39539,N_39464,N_39274);
and U39540 (N_39540,N_39446,N_39277);
xor U39541 (N_39541,N_39422,N_39270);
nand U39542 (N_39542,N_39340,N_39285);
or U39543 (N_39543,N_39426,N_39496);
xor U39544 (N_39544,N_39444,N_39272);
nor U39545 (N_39545,N_39408,N_39467);
nor U39546 (N_39546,N_39494,N_39334);
nand U39547 (N_39547,N_39264,N_39350);
nor U39548 (N_39548,N_39296,N_39387);
nand U39549 (N_39549,N_39420,N_39440);
or U39550 (N_39550,N_39432,N_39430);
nand U39551 (N_39551,N_39433,N_39326);
xnor U39552 (N_39552,N_39271,N_39267);
nor U39553 (N_39553,N_39352,N_39497);
xnor U39554 (N_39554,N_39345,N_39336);
xnor U39555 (N_39555,N_39293,N_39307);
nor U39556 (N_39556,N_39371,N_39366);
xnor U39557 (N_39557,N_39313,N_39380);
or U39558 (N_39558,N_39337,N_39353);
xor U39559 (N_39559,N_39447,N_39357);
or U39560 (N_39560,N_39253,N_39362);
nor U39561 (N_39561,N_39289,N_39394);
and U39562 (N_39562,N_39333,N_39436);
nor U39563 (N_39563,N_39367,N_39405);
nand U39564 (N_39564,N_39300,N_39255);
or U39565 (N_39565,N_39392,N_39407);
nand U39566 (N_39566,N_39335,N_39251);
or U39567 (N_39567,N_39346,N_39395);
or U39568 (N_39568,N_39411,N_39397);
nand U39569 (N_39569,N_39323,N_39290);
and U39570 (N_39570,N_39327,N_39419);
nand U39571 (N_39571,N_39466,N_39439);
xor U39572 (N_39572,N_39304,N_39311);
and U39573 (N_39573,N_39341,N_39431);
xnor U39574 (N_39574,N_39378,N_39417);
or U39575 (N_39575,N_39403,N_39457);
and U39576 (N_39576,N_39302,N_39491);
nand U39577 (N_39577,N_39338,N_39363);
nor U39578 (N_39578,N_39377,N_39332);
nand U39579 (N_39579,N_39498,N_39317);
and U39580 (N_39580,N_39453,N_39358);
or U39581 (N_39581,N_39391,N_39482);
or U39582 (N_39582,N_39250,N_39469);
xor U39583 (N_39583,N_39260,N_39463);
xnor U39584 (N_39584,N_39476,N_39356);
nand U39585 (N_39585,N_39268,N_39488);
or U39586 (N_39586,N_39276,N_39325);
xnor U39587 (N_39587,N_39368,N_39376);
or U39588 (N_39588,N_39360,N_39281);
nand U39589 (N_39589,N_39273,N_39421);
xor U39590 (N_39590,N_39294,N_39413);
nor U39591 (N_39591,N_39414,N_39489);
xor U39592 (N_39592,N_39318,N_39369);
or U39593 (N_39593,N_39309,N_39354);
xnor U39594 (N_39594,N_39372,N_39441);
nand U39595 (N_39595,N_39460,N_39480);
or U39596 (N_39596,N_39379,N_39478);
xnor U39597 (N_39597,N_39258,N_39370);
nor U39598 (N_39598,N_39389,N_39286);
xnor U39599 (N_39599,N_39485,N_39374);
or U39600 (N_39600,N_39316,N_39259);
nand U39601 (N_39601,N_39319,N_39283);
and U39602 (N_39602,N_39384,N_39351);
nor U39603 (N_39603,N_39456,N_39280);
xnor U39604 (N_39604,N_39343,N_39474);
nor U39605 (N_39605,N_39299,N_39322);
nor U39606 (N_39606,N_39324,N_39399);
and U39607 (N_39607,N_39287,N_39390);
nand U39608 (N_39608,N_39278,N_39375);
and U39609 (N_39609,N_39465,N_39314);
xor U39610 (N_39610,N_39495,N_39252);
or U39611 (N_39611,N_39261,N_39295);
xnor U39612 (N_39612,N_39310,N_39487);
nand U39613 (N_39613,N_39348,N_39401);
and U39614 (N_39614,N_39331,N_39288);
nor U39615 (N_39615,N_39484,N_39473);
xnor U39616 (N_39616,N_39462,N_39396);
nand U39617 (N_39617,N_39279,N_39291);
nand U39618 (N_39618,N_39308,N_39438);
nor U39619 (N_39619,N_39479,N_39284);
xnor U39620 (N_39620,N_39312,N_39415);
xnor U39621 (N_39621,N_39471,N_39410);
xnor U39622 (N_39622,N_39461,N_39451);
and U39623 (N_39623,N_39454,N_39427);
and U39624 (N_39624,N_39468,N_39450);
and U39625 (N_39625,N_39380,N_39310);
or U39626 (N_39626,N_39266,N_39443);
nor U39627 (N_39627,N_39426,N_39347);
nand U39628 (N_39628,N_39254,N_39291);
or U39629 (N_39629,N_39384,N_39293);
nand U39630 (N_39630,N_39266,N_39471);
nor U39631 (N_39631,N_39348,N_39404);
nand U39632 (N_39632,N_39400,N_39420);
or U39633 (N_39633,N_39277,N_39310);
or U39634 (N_39634,N_39301,N_39471);
xor U39635 (N_39635,N_39259,N_39315);
nand U39636 (N_39636,N_39393,N_39277);
nand U39637 (N_39637,N_39258,N_39329);
nor U39638 (N_39638,N_39283,N_39299);
nor U39639 (N_39639,N_39428,N_39370);
xnor U39640 (N_39640,N_39416,N_39383);
and U39641 (N_39641,N_39417,N_39360);
nand U39642 (N_39642,N_39404,N_39421);
and U39643 (N_39643,N_39325,N_39320);
or U39644 (N_39644,N_39466,N_39288);
nor U39645 (N_39645,N_39396,N_39328);
or U39646 (N_39646,N_39263,N_39357);
xor U39647 (N_39647,N_39429,N_39385);
xnor U39648 (N_39648,N_39328,N_39310);
xor U39649 (N_39649,N_39458,N_39489);
xnor U39650 (N_39650,N_39281,N_39321);
nand U39651 (N_39651,N_39338,N_39284);
nor U39652 (N_39652,N_39417,N_39369);
xor U39653 (N_39653,N_39374,N_39401);
xor U39654 (N_39654,N_39433,N_39297);
nand U39655 (N_39655,N_39278,N_39460);
nand U39656 (N_39656,N_39484,N_39270);
and U39657 (N_39657,N_39418,N_39456);
nand U39658 (N_39658,N_39270,N_39291);
and U39659 (N_39659,N_39488,N_39435);
and U39660 (N_39660,N_39373,N_39338);
or U39661 (N_39661,N_39435,N_39312);
xnor U39662 (N_39662,N_39442,N_39457);
nor U39663 (N_39663,N_39318,N_39404);
nor U39664 (N_39664,N_39347,N_39259);
xor U39665 (N_39665,N_39374,N_39346);
nor U39666 (N_39666,N_39346,N_39454);
and U39667 (N_39667,N_39428,N_39405);
and U39668 (N_39668,N_39312,N_39444);
nor U39669 (N_39669,N_39354,N_39414);
or U39670 (N_39670,N_39473,N_39318);
xnor U39671 (N_39671,N_39487,N_39277);
and U39672 (N_39672,N_39356,N_39355);
nand U39673 (N_39673,N_39262,N_39392);
and U39674 (N_39674,N_39494,N_39465);
xnor U39675 (N_39675,N_39285,N_39323);
nand U39676 (N_39676,N_39481,N_39405);
or U39677 (N_39677,N_39424,N_39314);
nor U39678 (N_39678,N_39407,N_39349);
nand U39679 (N_39679,N_39261,N_39312);
nand U39680 (N_39680,N_39339,N_39353);
nand U39681 (N_39681,N_39366,N_39487);
nor U39682 (N_39682,N_39443,N_39407);
nor U39683 (N_39683,N_39371,N_39278);
and U39684 (N_39684,N_39258,N_39423);
or U39685 (N_39685,N_39426,N_39285);
or U39686 (N_39686,N_39289,N_39398);
nand U39687 (N_39687,N_39325,N_39340);
xor U39688 (N_39688,N_39278,N_39327);
nor U39689 (N_39689,N_39357,N_39438);
and U39690 (N_39690,N_39385,N_39407);
or U39691 (N_39691,N_39384,N_39485);
or U39692 (N_39692,N_39280,N_39356);
or U39693 (N_39693,N_39421,N_39401);
or U39694 (N_39694,N_39435,N_39367);
and U39695 (N_39695,N_39398,N_39366);
xnor U39696 (N_39696,N_39359,N_39314);
xnor U39697 (N_39697,N_39463,N_39406);
nand U39698 (N_39698,N_39487,N_39307);
nor U39699 (N_39699,N_39302,N_39382);
nor U39700 (N_39700,N_39329,N_39394);
xor U39701 (N_39701,N_39281,N_39301);
nand U39702 (N_39702,N_39307,N_39467);
nor U39703 (N_39703,N_39361,N_39434);
xor U39704 (N_39704,N_39339,N_39487);
nor U39705 (N_39705,N_39358,N_39450);
and U39706 (N_39706,N_39291,N_39259);
or U39707 (N_39707,N_39440,N_39466);
or U39708 (N_39708,N_39295,N_39490);
nor U39709 (N_39709,N_39269,N_39306);
and U39710 (N_39710,N_39441,N_39318);
nand U39711 (N_39711,N_39252,N_39417);
nor U39712 (N_39712,N_39452,N_39361);
nand U39713 (N_39713,N_39458,N_39490);
xor U39714 (N_39714,N_39343,N_39321);
and U39715 (N_39715,N_39314,N_39394);
nor U39716 (N_39716,N_39332,N_39462);
xnor U39717 (N_39717,N_39368,N_39322);
nor U39718 (N_39718,N_39320,N_39426);
and U39719 (N_39719,N_39408,N_39444);
nor U39720 (N_39720,N_39479,N_39458);
nor U39721 (N_39721,N_39265,N_39475);
nand U39722 (N_39722,N_39397,N_39352);
xor U39723 (N_39723,N_39316,N_39358);
and U39724 (N_39724,N_39470,N_39298);
xnor U39725 (N_39725,N_39314,N_39428);
xor U39726 (N_39726,N_39489,N_39433);
xor U39727 (N_39727,N_39371,N_39497);
or U39728 (N_39728,N_39331,N_39345);
or U39729 (N_39729,N_39309,N_39366);
or U39730 (N_39730,N_39449,N_39378);
xor U39731 (N_39731,N_39302,N_39281);
or U39732 (N_39732,N_39497,N_39416);
and U39733 (N_39733,N_39367,N_39408);
nand U39734 (N_39734,N_39287,N_39319);
or U39735 (N_39735,N_39324,N_39471);
and U39736 (N_39736,N_39419,N_39478);
nor U39737 (N_39737,N_39388,N_39477);
nor U39738 (N_39738,N_39375,N_39402);
or U39739 (N_39739,N_39488,N_39257);
or U39740 (N_39740,N_39310,N_39302);
nor U39741 (N_39741,N_39253,N_39310);
nand U39742 (N_39742,N_39385,N_39489);
and U39743 (N_39743,N_39357,N_39456);
nand U39744 (N_39744,N_39393,N_39490);
and U39745 (N_39745,N_39305,N_39452);
and U39746 (N_39746,N_39462,N_39428);
nor U39747 (N_39747,N_39280,N_39427);
and U39748 (N_39748,N_39414,N_39433);
nand U39749 (N_39749,N_39481,N_39459);
nor U39750 (N_39750,N_39658,N_39526);
xor U39751 (N_39751,N_39509,N_39726);
nor U39752 (N_39752,N_39689,N_39605);
and U39753 (N_39753,N_39550,N_39534);
or U39754 (N_39754,N_39731,N_39717);
nand U39755 (N_39755,N_39553,N_39743);
or U39756 (N_39756,N_39657,N_39711);
or U39757 (N_39757,N_39632,N_39571);
or U39758 (N_39758,N_39662,N_39660);
or U39759 (N_39759,N_39502,N_39646);
nor U39760 (N_39760,N_39670,N_39671);
and U39761 (N_39761,N_39531,N_39722);
and U39762 (N_39762,N_39615,N_39674);
and U39763 (N_39763,N_39572,N_39709);
or U39764 (N_39764,N_39513,N_39608);
or U39765 (N_39765,N_39563,N_39593);
and U39766 (N_39766,N_39595,N_39638);
nand U39767 (N_39767,N_39611,N_39721);
xnor U39768 (N_39768,N_39644,N_39610);
xor U39769 (N_39769,N_39654,N_39697);
and U39770 (N_39770,N_39533,N_39728);
or U39771 (N_39771,N_39516,N_39524);
or U39772 (N_39772,N_39588,N_39740);
or U39773 (N_39773,N_39624,N_39590);
nand U39774 (N_39774,N_39681,N_39505);
xor U39775 (N_39775,N_39555,N_39659);
and U39776 (N_39776,N_39639,N_39506);
nor U39777 (N_39777,N_39562,N_39637);
or U39778 (N_39778,N_39700,N_39733);
and U39779 (N_39779,N_39621,N_39735);
nor U39780 (N_39780,N_39596,N_39656);
nand U39781 (N_39781,N_39585,N_39742);
xnor U39782 (N_39782,N_39633,N_39650);
or U39783 (N_39783,N_39529,N_39609);
nand U39784 (N_39784,N_39518,N_39686);
nor U39785 (N_39785,N_39747,N_39629);
or U39786 (N_39786,N_39554,N_39668);
xor U39787 (N_39787,N_39661,N_39545);
nand U39788 (N_39788,N_39580,N_39577);
xor U39789 (N_39789,N_39582,N_39692);
or U39790 (N_39790,N_39647,N_39521);
nand U39791 (N_39791,N_39579,N_39586);
or U39792 (N_39792,N_39578,N_39520);
nand U39793 (N_39793,N_39535,N_39548);
and U39794 (N_39794,N_39745,N_39527);
xnor U39795 (N_39795,N_39699,N_39549);
nor U39796 (N_39796,N_39667,N_39669);
nor U39797 (N_39797,N_39634,N_39616);
nand U39798 (N_39798,N_39687,N_39641);
or U39799 (N_39799,N_39591,N_39623);
nor U39800 (N_39800,N_39741,N_39613);
and U39801 (N_39801,N_39603,N_39501);
xnor U39802 (N_39802,N_39685,N_39708);
nand U39803 (N_39803,N_39503,N_39748);
xor U39804 (N_39804,N_39515,N_39665);
xnor U39805 (N_39805,N_39507,N_39604);
nor U39806 (N_39806,N_39607,N_39569);
xor U39807 (N_39807,N_39560,N_39636);
nand U39808 (N_39808,N_39725,N_39703);
and U39809 (N_39809,N_39683,N_39532);
nand U39810 (N_39810,N_39508,N_39598);
nor U39811 (N_39811,N_39587,N_39592);
or U39812 (N_39812,N_39602,N_39525);
xnor U39813 (N_39813,N_39694,N_39583);
xor U39814 (N_39814,N_39576,N_39677);
nand U39815 (N_39815,N_39626,N_39652);
xor U39816 (N_39816,N_39619,N_39540);
or U39817 (N_39817,N_39566,N_39600);
nand U39818 (N_39818,N_39723,N_39691);
nand U39819 (N_39819,N_39589,N_39517);
nand U39820 (N_39820,N_39710,N_39736);
and U39821 (N_39821,N_39749,N_39599);
nand U39822 (N_39822,N_39706,N_39564);
and U39823 (N_39823,N_39541,N_39746);
nand U39824 (N_39824,N_39631,N_39559);
and U39825 (N_39825,N_39575,N_39614);
nand U39826 (N_39826,N_39538,N_39622);
nor U39827 (N_39827,N_39567,N_39594);
and U39828 (N_39828,N_39556,N_39730);
xor U39829 (N_39829,N_39537,N_39546);
and U39830 (N_39830,N_39744,N_39584);
nor U39831 (N_39831,N_39542,N_39682);
and U39832 (N_39832,N_39678,N_39568);
nand U39833 (N_39833,N_39719,N_39701);
nor U39834 (N_39834,N_39734,N_39528);
nor U39835 (N_39835,N_39617,N_39739);
xor U39836 (N_39836,N_39544,N_39536);
or U39837 (N_39837,N_39597,N_39601);
or U39838 (N_39838,N_39547,N_39581);
or U39839 (N_39839,N_39514,N_39565);
and U39840 (N_39840,N_39630,N_39684);
nand U39841 (N_39841,N_39504,N_39695);
nand U39842 (N_39842,N_39557,N_39643);
nand U39843 (N_39843,N_39673,N_39651);
nand U39844 (N_39844,N_39628,N_39642);
or U39845 (N_39845,N_39672,N_39698);
xnor U39846 (N_39846,N_39663,N_39618);
and U39847 (N_39847,N_39655,N_39612);
or U39848 (N_39848,N_39606,N_39570);
nor U39849 (N_39849,N_39724,N_39511);
nand U39850 (N_39850,N_39649,N_39648);
nor U39851 (N_39851,N_39737,N_39705);
nor U39852 (N_39852,N_39552,N_39558);
nor U39853 (N_39853,N_39551,N_39543);
and U39854 (N_39854,N_39696,N_39519);
nor U39855 (N_39855,N_39512,N_39635);
nand U39856 (N_39856,N_39653,N_39688);
and U39857 (N_39857,N_39713,N_39707);
or U39858 (N_39858,N_39625,N_39573);
or U39859 (N_39859,N_39738,N_39727);
nand U39860 (N_39860,N_39732,N_39693);
nor U39861 (N_39861,N_39714,N_39680);
nor U39862 (N_39862,N_39574,N_39712);
xnor U39863 (N_39863,N_39500,N_39666);
and U39864 (N_39864,N_39716,N_39522);
nand U39865 (N_39865,N_39561,N_39729);
and U39866 (N_39866,N_39690,N_39720);
and U39867 (N_39867,N_39704,N_39676);
and U39868 (N_39868,N_39627,N_39523);
xor U39869 (N_39869,N_39718,N_39645);
or U39870 (N_39870,N_39675,N_39530);
nand U39871 (N_39871,N_39702,N_39620);
nand U39872 (N_39872,N_39715,N_39539);
xnor U39873 (N_39873,N_39510,N_39679);
and U39874 (N_39874,N_39640,N_39664);
nor U39875 (N_39875,N_39655,N_39718);
and U39876 (N_39876,N_39730,N_39582);
nand U39877 (N_39877,N_39587,N_39729);
xnor U39878 (N_39878,N_39617,N_39737);
or U39879 (N_39879,N_39748,N_39550);
or U39880 (N_39880,N_39653,N_39690);
nand U39881 (N_39881,N_39748,N_39731);
xnor U39882 (N_39882,N_39707,N_39606);
nand U39883 (N_39883,N_39551,N_39701);
nor U39884 (N_39884,N_39555,N_39576);
or U39885 (N_39885,N_39621,N_39581);
and U39886 (N_39886,N_39667,N_39537);
nand U39887 (N_39887,N_39585,N_39661);
or U39888 (N_39888,N_39683,N_39641);
and U39889 (N_39889,N_39516,N_39543);
nand U39890 (N_39890,N_39740,N_39744);
nand U39891 (N_39891,N_39532,N_39743);
and U39892 (N_39892,N_39698,N_39624);
nor U39893 (N_39893,N_39554,N_39660);
xnor U39894 (N_39894,N_39503,N_39674);
and U39895 (N_39895,N_39521,N_39630);
or U39896 (N_39896,N_39641,N_39734);
nor U39897 (N_39897,N_39734,N_39507);
nor U39898 (N_39898,N_39676,N_39728);
and U39899 (N_39899,N_39582,N_39689);
nor U39900 (N_39900,N_39593,N_39623);
nor U39901 (N_39901,N_39720,N_39727);
or U39902 (N_39902,N_39642,N_39661);
nor U39903 (N_39903,N_39715,N_39555);
nor U39904 (N_39904,N_39666,N_39589);
xnor U39905 (N_39905,N_39582,N_39607);
nand U39906 (N_39906,N_39559,N_39546);
nand U39907 (N_39907,N_39574,N_39694);
xnor U39908 (N_39908,N_39741,N_39746);
or U39909 (N_39909,N_39539,N_39536);
and U39910 (N_39910,N_39596,N_39558);
or U39911 (N_39911,N_39634,N_39507);
xor U39912 (N_39912,N_39639,N_39698);
or U39913 (N_39913,N_39540,N_39593);
and U39914 (N_39914,N_39510,N_39656);
and U39915 (N_39915,N_39719,N_39728);
nand U39916 (N_39916,N_39555,N_39738);
and U39917 (N_39917,N_39736,N_39601);
nor U39918 (N_39918,N_39677,N_39613);
nand U39919 (N_39919,N_39713,N_39617);
nor U39920 (N_39920,N_39746,N_39561);
or U39921 (N_39921,N_39598,N_39709);
and U39922 (N_39922,N_39538,N_39712);
or U39923 (N_39923,N_39739,N_39565);
nor U39924 (N_39924,N_39699,N_39671);
or U39925 (N_39925,N_39718,N_39631);
xnor U39926 (N_39926,N_39725,N_39563);
xnor U39927 (N_39927,N_39581,N_39573);
and U39928 (N_39928,N_39537,N_39615);
and U39929 (N_39929,N_39501,N_39593);
and U39930 (N_39930,N_39595,N_39531);
or U39931 (N_39931,N_39713,N_39748);
nand U39932 (N_39932,N_39512,N_39662);
nor U39933 (N_39933,N_39741,N_39531);
nor U39934 (N_39934,N_39706,N_39557);
or U39935 (N_39935,N_39731,N_39594);
or U39936 (N_39936,N_39675,N_39682);
or U39937 (N_39937,N_39576,N_39675);
nor U39938 (N_39938,N_39553,N_39746);
xor U39939 (N_39939,N_39519,N_39511);
and U39940 (N_39940,N_39631,N_39545);
nand U39941 (N_39941,N_39715,N_39617);
nand U39942 (N_39942,N_39697,N_39681);
nand U39943 (N_39943,N_39656,N_39644);
xor U39944 (N_39944,N_39624,N_39593);
or U39945 (N_39945,N_39565,N_39702);
and U39946 (N_39946,N_39566,N_39693);
and U39947 (N_39947,N_39586,N_39738);
nand U39948 (N_39948,N_39599,N_39546);
nand U39949 (N_39949,N_39592,N_39516);
or U39950 (N_39950,N_39743,N_39513);
or U39951 (N_39951,N_39510,N_39519);
and U39952 (N_39952,N_39543,N_39624);
or U39953 (N_39953,N_39724,N_39732);
nand U39954 (N_39954,N_39612,N_39509);
or U39955 (N_39955,N_39670,N_39689);
or U39956 (N_39956,N_39721,N_39693);
nand U39957 (N_39957,N_39669,N_39508);
and U39958 (N_39958,N_39710,N_39732);
or U39959 (N_39959,N_39560,N_39577);
and U39960 (N_39960,N_39585,N_39517);
and U39961 (N_39961,N_39703,N_39600);
xor U39962 (N_39962,N_39708,N_39748);
xor U39963 (N_39963,N_39692,N_39684);
or U39964 (N_39964,N_39718,N_39600);
nor U39965 (N_39965,N_39649,N_39736);
or U39966 (N_39966,N_39537,N_39530);
or U39967 (N_39967,N_39602,N_39556);
nand U39968 (N_39968,N_39704,N_39505);
nor U39969 (N_39969,N_39682,N_39690);
and U39970 (N_39970,N_39626,N_39631);
xnor U39971 (N_39971,N_39568,N_39732);
xnor U39972 (N_39972,N_39622,N_39566);
or U39973 (N_39973,N_39667,N_39503);
and U39974 (N_39974,N_39573,N_39602);
or U39975 (N_39975,N_39709,N_39675);
nand U39976 (N_39976,N_39730,N_39609);
xor U39977 (N_39977,N_39617,N_39596);
or U39978 (N_39978,N_39745,N_39581);
nand U39979 (N_39979,N_39666,N_39509);
or U39980 (N_39980,N_39678,N_39585);
or U39981 (N_39981,N_39509,N_39650);
nand U39982 (N_39982,N_39532,N_39682);
nor U39983 (N_39983,N_39673,N_39534);
nand U39984 (N_39984,N_39589,N_39656);
or U39985 (N_39985,N_39568,N_39513);
and U39986 (N_39986,N_39685,N_39508);
or U39987 (N_39987,N_39621,N_39542);
nor U39988 (N_39988,N_39518,N_39558);
and U39989 (N_39989,N_39526,N_39587);
and U39990 (N_39990,N_39711,N_39655);
nand U39991 (N_39991,N_39664,N_39724);
nand U39992 (N_39992,N_39523,N_39737);
or U39993 (N_39993,N_39744,N_39633);
or U39994 (N_39994,N_39560,N_39714);
or U39995 (N_39995,N_39515,N_39626);
nand U39996 (N_39996,N_39565,N_39721);
or U39997 (N_39997,N_39736,N_39528);
xor U39998 (N_39998,N_39680,N_39603);
nor U39999 (N_39999,N_39716,N_39642);
nand U40000 (N_40000,N_39823,N_39842);
xor U40001 (N_40001,N_39762,N_39989);
nor U40002 (N_40002,N_39759,N_39908);
and U40003 (N_40003,N_39856,N_39904);
nand U40004 (N_40004,N_39943,N_39988);
and U40005 (N_40005,N_39792,N_39852);
nor U40006 (N_40006,N_39986,N_39814);
and U40007 (N_40007,N_39952,N_39895);
nand U40008 (N_40008,N_39974,N_39880);
or U40009 (N_40009,N_39956,N_39836);
nor U40010 (N_40010,N_39793,N_39821);
or U40011 (N_40011,N_39907,N_39915);
xor U40012 (N_40012,N_39857,N_39991);
or U40013 (N_40013,N_39910,N_39838);
xnor U40014 (N_40014,N_39903,N_39841);
xor U40015 (N_40015,N_39861,N_39794);
nand U40016 (N_40016,N_39833,N_39977);
or U40017 (N_40017,N_39869,N_39960);
nor U40018 (N_40018,N_39967,N_39978);
nand U40019 (N_40019,N_39775,N_39800);
nand U40020 (N_40020,N_39834,N_39958);
or U40021 (N_40021,N_39892,N_39939);
nor U40022 (N_40022,N_39803,N_39786);
or U40023 (N_40023,N_39763,N_39783);
nand U40024 (N_40024,N_39914,N_39755);
and U40025 (N_40025,N_39980,N_39864);
xnor U40026 (N_40026,N_39931,N_39828);
or U40027 (N_40027,N_39971,N_39934);
nor U40028 (N_40028,N_39900,N_39999);
xor U40029 (N_40029,N_39951,N_39965);
xnor U40030 (N_40030,N_39940,N_39901);
nand U40031 (N_40031,N_39799,N_39805);
and U40032 (N_40032,N_39837,N_39987);
nand U40033 (N_40033,N_39964,N_39947);
nor U40034 (N_40034,N_39764,N_39825);
xor U40035 (N_40035,N_39995,N_39822);
nand U40036 (N_40036,N_39813,N_39916);
and U40037 (N_40037,N_39998,N_39984);
and U40038 (N_40038,N_39871,N_39779);
nor U40039 (N_40039,N_39877,N_39961);
or U40040 (N_40040,N_39906,N_39854);
xor U40041 (N_40041,N_39752,N_39750);
nor U40042 (N_40042,N_39795,N_39777);
nand U40043 (N_40043,N_39885,N_39992);
or U40044 (N_40044,N_39846,N_39886);
xor U40045 (N_40045,N_39982,N_39948);
nand U40046 (N_40046,N_39928,N_39776);
nor U40047 (N_40047,N_39949,N_39754);
xnor U40048 (N_40048,N_39831,N_39913);
nor U40049 (N_40049,N_39756,N_39769);
nand U40050 (N_40050,N_39780,N_39839);
and U40051 (N_40051,N_39757,N_39894);
nor U40052 (N_40052,N_39772,N_39898);
nor U40053 (N_40053,N_39774,N_39850);
and U40054 (N_40054,N_39881,N_39860);
xnor U40055 (N_40055,N_39851,N_39816);
and U40056 (N_40056,N_39879,N_39981);
xor U40057 (N_40057,N_39890,N_39758);
xnor U40058 (N_40058,N_39897,N_39902);
or U40059 (N_40059,N_39870,N_39953);
nand U40060 (N_40060,N_39873,N_39760);
nor U40061 (N_40061,N_39927,N_39941);
xnor U40062 (N_40062,N_39801,N_39920);
nor U40063 (N_40063,N_39933,N_39843);
and U40064 (N_40064,N_39863,N_39945);
nor U40065 (N_40065,N_39924,N_39918);
xor U40066 (N_40066,N_39993,N_39950);
or U40067 (N_40067,N_39787,N_39847);
xnor U40068 (N_40068,N_39808,N_39824);
or U40069 (N_40069,N_39909,N_39936);
and U40070 (N_40070,N_39942,N_39938);
and U40071 (N_40071,N_39753,N_39922);
xor U40072 (N_40072,N_39855,N_39973);
or U40073 (N_40073,N_39815,N_39806);
nand U40074 (N_40074,N_39893,N_39859);
and U40075 (N_40075,N_39807,N_39921);
nand U40076 (N_40076,N_39853,N_39882);
nand U40077 (N_40077,N_39896,N_39874);
xnor U40078 (N_40078,N_39925,N_39875);
nor U40079 (N_40079,N_39791,N_39996);
nor U40080 (N_40080,N_39970,N_39862);
and U40081 (N_40081,N_39983,N_39751);
nand U40082 (N_40082,N_39818,N_39866);
xor U40083 (N_40083,N_39935,N_39826);
nor U40084 (N_40084,N_39923,N_39972);
nand U40085 (N_40085,N_39832,N_39761);
nor U40086 (N_40086,N_39946,N_39809);
or U40087 (N_40087,N_39932,N_39883);
xor U40088 (N_40088,N_39835,N_39830);
nand U40089 (N_40089,N_39990,N_39849);
nor U40090 (N_40090,N_39976,N_39929);
nor U40091 (N_40091,N_39785,N_39868);
or U40092 (N_40092,N_39802,N_39781);
nor U40093 (N_40093,N_39889,N_39899);
or U40094 (N_40094,N_39926,N_39966);
nand U40095 (N_40095,N_39789,N_39810);
and U40096 (N_40096,N_39829,N_39905);
xor U40097 (N_40097,N_39765,N_39876);
or U40098 (N_40098,N_39937,N_39930);
nand U40099 (N_40099,N_39975,N_39827);
and U40100 (N_40100,N_39865,N_39817);
nor U40101 (N_40101,N_39944,N_39848);
or U40102 (N_40102,N_39954,N_39878);
and U40103 (N_40103,N_39917,N_39812);
and U40104 (N_40104,N_39985,N_39912);
and U40105 (N_40105,N_39955,N_39969);
or U40106 (N_40106,N_39820,N_39957);
xor U40107 (N_40107,N_39784,N_39804);
and U40108 (N_40108,N_39819,N_39962);
and U40109 (N_40109,N_39811,N_39767);
nor U40110 (N_40110,N_39773,N_39845);
nand U40111 (N_40111,N_39959,N_39782);
nand U40112 (N_40112,N_39884,N_39778);
nor U40113 (N_40113,N_39844,N_39979);
xor U40114 (N_40114,N_39858,N_39798);
xor U40115 (N_40115,N_39888,N_39768);
nor U40116 (N_40116,N_39796,N_39919);
and U40117 (N_40117,N_39770,N_39994);
and U40118 (N_40118,N_39766,N_39891);
xor U40119 (N_40119,N_39797,N_39790);
nor U40120 (N_40120,N_39963,N_39911);
xor U40121 (N_40121,N_39872,N_39968);
or U40122 (N_40122,N_39997,N_39840);
nand U40123 (N_40123,N_39771,N_39867);
nand U40124 (N_40124,N_39788,N_39887);
nor U40125 (N_40125,N_39811,N_39786);
xor U40126 (N_40126,N_39854,N_39828);
or U40127 (N_40127,N_39823,N_39784);
xor U40128 (N_40128,N_39762,N_39876);
or U40129 (N_40129,N_39892,N_39823);
and U40130 (N_40130,N_39885,N_39855);
and U40131 (N_40131,N_39903,N_39788);
nor U40132 (N_40132,N_39923,N_39779);
xnor U40133 (N_40133,N_39784,N_39886);
xor U40134 (N_40134,N_39773,N_39889);
xor U40135 (N_40135,N_39901,N_39758);
nor U40136 (N_40136,N_39787,N_39867);
nor U40137 (N_40137,N_39884,N_39787);
or U40138 (N_40138,N_39898,N_39838);
or U40139 (N_40139,N_39764,N_39947);
or U40140 (N_40140,N_39796,N_39857);
or U40141 (N_40141,N_39807,N_39810);
and U40142 (N_40142,N_39784,N_39830);
nand U40143 (N_40143,N_39897,N_39777);
and U40144 (N_40144,N_39909,N_39952);
xnor U40145 (N_40145,N_39853,N_39931);
nor U40146 (N_40146,N_39810,N_39774);
and U40147 (N_40147,N_39753,N_39771);
xnor U40148 (N_40148,N_39998,N_39959);
nor U40149 (N_40149,N_39767,N_39940);
nor U40150 (N_40150,N_39851,N_39994);
or U40151 (N_40151,N_39903,N_39810);
or U40152 (N_40152,N_39764,N_39768);
xnor U40153 (N_40153,N_39751,N_39928);
nand U40154 (N_40154,N_39938,N_39774);
xnor U40155 (N_40155,N_39810,N_39866);
or U40156 (N_40156,N_39928,N_39768);
xnor U40157 (N_40157,N_39878,N_39862);
nand U40158 (N_40158,N_39957,N_39909);
and U40159 (N_40159,N_39902,N_39914);
xor U40160 (N_40160,N_39765,N_39860);
nor U40161 (N_40161,N_39800,N_39905);
nand U40162 (N_40162,N_39945,N_39758);
or U40163 (N_40163,N_39776,N_39940);
xnor U40164 (N_40164,N_39791,N_39790);
or U40165 (N_40165,N_39992,N_39912);
xor U40166 (N_40166,N_39750,N_39819);
nand U40167 (N_40167,N_39941,N_39957);
xor U40168 (N_40168,N_39799,N_39854);
xnor U40169 (N_40169,N_39919,N_39865);
or U40170 (N_40170,N_39923,N_39810);
or U40171 (N_40171,N_39770,N_39880);
xor U40172 (N_40172,N_39914,N_39786);
xnor U40173 (N_40173,N_39754,N_39791);
or U40174 (N_40174,N_39926,N_39984);
nand U40175 (N_40175,N_39938,N_39921);
nor U40176 (N_40176,N_39921,N_39802);
xor U40177 (N_40177,N_39822,N_39998);
nor U40178 (N_40178,N_39959,N_39836);
and U40179 (N_40179,N_39774,N_39936);
nor U40180 (N_40180,N_39906,N_39982);
and U40181 (N_40181,N_39993,N_39825);
or U40182 (N_40182,N_39772,N_39863);
xnor U40183 (N_40183,N_39763,N_39815);
xor U40184 (N_40184,N_39805,N_39858);
or U40185 (N_40185,N_39789,N_39814);
and U40186 (N_40186,N_39913,N_39797);
nor U40187 (N_40187,N_39961,N_39808);
nor U40188 (N_40188,N_39977,N_39750);
xor U40189 (N_40189,N_39883,N_39979);
and U40190 (N_40190,N_39771,N_39878);
xnor U40191 (N_40191,N_39852,N_39970);
nor U40192 (N_40192,N_39780,N_39812);
xnor U40193 (N_40193,N_39872,N_39995);
xnor U40194 (N_40194,N_39996,N_39770);
or U40195 (N_40195,N_39902,N_39975);
or U40196 (N_40196,N_39973,N_39829);
xnor U40197 (N_40197,N_39917,N_39839);
and U40198 (N_40198,N_39985,N_39904);
nor U40199 (N_40199,N_39963,N_39992);
nor U40200 (N_40200,N_39894,N_39798);
or U40201 (N_40201,N_39773,N_39765);
xor U40202 (N_40202,N_39985,N_39896);
or U40203 (N_40203,N_39759,N_39814);
and U40204 (N_40204,N_39883,N_39753);
nor U40205 (N_40205,N_39772,N_39855);
xnor U40206 (N_40206,N_39909,N_39889);
xor U40207 (N_40207,N_39810,N_39863);
nand U40208 (N_40208,N_39846,N_39902);
xor U40209 (N_40209,N_39758,N_39775);
and U40210 (N_40210,N_39750,N_39764);
or U40211 (N_40211,N_39869,N_39881);
or U40212 (N_40212,N_39815,N_39906);
xnor U40213 (N_40213,N_39820,N_39786);
and U40214 (N_40214,N_39777,N_39959);
or U40215 (N_40215,N_39804,N_39963);
or U40216 (N_40216,N_39792,N_39768);
nor U40217 (N_40217,N_39754,N_39830);
nor U40218 (N_40218,N_39915,N_39908);
nand U40219 (N_40219,N_39817,N_39921);
and U40220 (N_40220,N_39773,N_39877);
nor U40221 (N_40221,N_39903,N_39784);
and U40222 (N_40222,N_39979,N_39982);
xor U40223 (N_40223,N_39853,N_39875);
nand U40224 (N_40224,N_39806,N_39886);
or U40225 (N_40225,N_39985,N_39909);
nor U40226 (N_40226,N_39978,N_39841);
and U40227 (N_40227,N_39937,N_39906);
nor U40228 (N_40228,N_39869,N_39985);
nand U40229 (N_40229,N_39946,N_39863);
or U40230 (N_40230,N_39900,N_39842);
or U40231 (N_40231,N_39765,N_39958);
nand U40232 (N_40232,N_39868,N_39775);
xnor U40233 (N_40233,N_39758,N_39825);
xnor U40234 (N_40234,N_39829,N_39985);
nor U40235 (N_40235,N_39762,N_39786);
nor U40236 (N_40236,N_39832,N_39967);
xnor U40237 (N_40237,N_39771,N_39963);
xor U40238 (N_40238,N_39755,N_39809);
or U40239 (N_40239,N_39921,N_39844);
nand U40240 (N_40240,N_39784,N_39911);
and U40241 (N_40241,N_39862,N_39884);
nor U40242 (N_40242,N_39842,N_39847);
xnor U40243 (N_40243,N_39905,N_39818);
xnor U40244 (N_40244,N_39953,N_39949);
xor U40245 (N_40245,N_39824,N_39977);
and U40246 (N_40246,N_39933,N_39768);
nor U40247 (N_40247,N_39914,N_39941);
xnor U40248 (N_40248,N_39772,N_39814);
nor U40249 (N_40249,N_39962,N_39914);
and U40250 (N_40250,N_40049,N_40230);
nand U40251 (N_40251,N_40108,N_40127);
xnor U40252 (N_40252,N_40027,N_40074);
or U40253 (N_40253,N_40103,N_40234);
and U40254 (N_40254,N_40000,N_40132);
or U40255 (N_40255,N_40231,N_40058);
and U40256 (N_40256,N_40240,N_40140);
and U40257 (N_40257,N_40122,N_40023);
nor U40258 (N_40258,N_40118,N_40065);
nor U40259 (N_40259,N_40172,N_40150);
xnor U40260 (N_40260,N_40025,N_40204);
xor U40261 (N_40261,N_40142,N_40081);
nor U40262 (N_40262,N_40021,N_40246);
nor U40263 (N_40263,N_40163,N_40038);
xor U40264 (N_40264,N_40003,N_40046);
xor U40265 (N_40265,N_40193,N_40123);
xor U40266 (N_40266,N_40220,N_40181);
nand U40267 (N_40267,N_40121,N_40094);
nor U40268 (N_40268,N_40047,N_40226);
nor U40269 (N_40269,N_40107,N_40198);
and U40270 (N_40270,N_40171,N_40066);
nor U40271 (N_40271,N_40174,N_40165);
or U40272 (N_40272,N_40008,N_40239);
nand U40273 (N_40273,N_40153,N_40031);
nand U40274 (N_40274,N_40005,N_40120);
nor U40275 (N_40275,N_40125,N_40068);
nand U40276 (N_40276,N_40102,N_40004);
or U40277 (N_40277,N_40117,N_40087);
nor U40278 (N_40278,N_40183,N_40148);
xnor U40279 (N_40279,N_40137,N_40196);
nor U40280 (N_40280,N_40055,N_40219);
xor U40281 (N_40281,N_40166,N_40061);
nand U40282 (N_40282,N_40216,N_40072);
nand U40283 (N_40283,N_40029,N_40156);
nor U40284 (N_40284,N_40147,N_40212);
and U40285 (N_40285,N_40160,N_40069);
or U40286 (N_40286,N_40217,N_40113);
xor U40287 (N_40287,N_40187,N_40151);
or U40288 (N_40288,N_40135,N_40085);
nor U40289 (N_40289,N_40026,N_40152);
xnor U40290 (N_40290,N_40018,N_40001);
and U40291 (N_40291,N_40073,N_40225);
nand U40292 (N_40292,N_40042,N_40243);
nand U40293 (N_40293,N_40017,N_40173);
nor U40294 (N_40294,N_40112,N_40009);
nand U40295 (N_40295,N_40157,N_40095);
or U40296 (N_40296,N_40247,N_40090);
nand U40297 (N_40297,N_40197,N_40161);
nor U40298 (N_40298,N_40075,N_40249);
and U40299 (N_40299,N_40080,N_40209);
or U40300 (N_40300,N_40201,N_40126);
nor U40301 (N_40301,N_40109,N_40050);
nor U40302 (N_40302,N_40099,N_40010);
xnor U40303 (N_40303,N_40052,N_40070);
nand U40304 (N_40304,N_40175,N_40245);
nor U40305 (N_40305,N_40097,N_40028);
or U40306 (N_40306,N_40054,N_40096);
and U40307 (N_40307,N_40228,N_40200);
xor U40308 (N_40308,N_40242,N_40144);
xnor U40309 (N_40309,N_40128,N_40088);
nand U40310 (N_40310,N_40168,N_40015);
nor U40311 (N_40311,N_40215,N_40138);
and U40312 (N_40312,N_40213,N_40040);
nor U40313 (N_40313,N_40111,N_40169);
or U40314 (N_40314,N_40011,N_40104);
xor U40315 (N_40315,N_40149,N_40227);
nand U40316 (N_40316,N_40019,N_40034);
nor U40317 (N_40317,N_40022,N_40244);
nor U40318 (N_40318,N_40179,N_40237);
nand U40319 (N_40319,N_40032,N_40098);
xor U40320 (N_40320,N_40083,N_40006);
xnor U40321 (N_40321,N_40170,N_40101);
xor U40322 (N_40322,N_40207,N_40091);
xor U40323 (N_40323,N_40202,N_40235);
xor U40324 (N_40324,N_40192,N_40191);
and U40325 (N_40325,N_40116,N_40036);
nor U40326 (N_40326,N_40189,N_40063);
or U40327 (N_40327,N_40092,N_40035);
xor U40328 (N_40328,N_40139,N_40110);
and U40329 (N_40329,N_40182,N_40007);
xnor U40330 (N_40330,N_40030,N_40154);
xnor U40331 (N_40331,N_40248,N_40199);
and U40332 (N_40332,N_40190,N_40041);
or U40333 (N_40333,N_40186,N_40057);
nand U40334 (N_40334,N_40155,N_40124);
and U40335 (N_40335,N_40079,N_40229);
and U40336 (N_40336,N_40134,N_40059);
or U40337 (N_40337,N_40013,N_40039);
nand U40338 (N_40338,N_40131,N_40067);
nand U40339 (N_40339,N_40176,N_40221);
or U40340 (N_40340,N_40214,N_40222);
and U40341 (N_40341,N_40082,N_40146);
xnor U40342 (N_40342,N_40053,N_40188);
nand U40343 (N_40343,N_40205,N_40002);
or U40344 (N_40344,N_40224,N_40100);
or U40345 (N_40345,N_40012,N_40093);
xor U40346 (N_40346,N_40185,N_40143);
nand U40347 (N_40347,N_40145,N_40133);
or U40348 (N_40348,N_40194,N_40195);
xnor U40349 (N_40349,N_40130,N_40203);
nor U40350 (N_40350,N_40105,N_40033);
nor U40351 (N_40351,N_40180,N_40115);
or U40352 (N_40352,N_40086,N_40020);
nor U40353 (N_40353,N_40223,N_40084);
nand U40354 (N_40354,N_40159,N_40236);
xnor U40355 (N_40355,N_40208,N_40106);
xnor U40356 (N_40356,N_40044,N_40119);
or U40357 (N_40357,N_40051,N_40211);
and U40358 (N_40358,N_40162,N_40136);
xor U40359 (N_40359,N_40232,N_40177);
and U40360 (N_40360,N_40071,N_40178);
nor U40361 (N_40361,N_40210,N_40241);
nor U40362 (N_40362,N_40238,N_40060);
and U40363 (N_40363,N_40233,N_40218);
and U40364 (N_40364,N_40114,N_40158);
nor U40365 (N_40365,N_40141,N_40076);
xnor U40366 (N_40366,N_40045,N_40024);
xor U40367 (N_40367,N_40089,N_40129);
nor U40368 (N_40368,N_40014,N_40184);
and U40369 (N_40369,N_40206,N_40167);
and U40370 (N_40370,N_40164,N_40064);
or U40371 (N_40371,N_40077,N_40078);
nor U40372 (N_40372,N_40062,N_40048);
or U40373 (N_40373,N_40043,N_40037);
nand U40374 (N_40374,N_40056,N_40016);
and U40375 (N_40375,N_40179,N_40086);
nand U40376 (N_40376,N_40057,N_40056);
nor U40377 (N_40377,N_40043,N_40227);
nor U40378 (N_40378,N_40182,N_40148);
nand U40379 (N_40379,N_40014,N_40130);
nand U40380 (N_40380,N_40174,N_40087);
xor U40381 (N_40381,N_40160,N_40116);
nand U40382 (N_40382,N_40224,N_40229);
or U40383 (N_40383,N_40192,N_40116);
nor U40384 (N_40384,N_40095,N_40206);
and U40385 (N_40385,N_40010,N_40209);
nand U40386 (N_40386,N_40089,N_40205);
nor U40387 (N_40387,N_40088,N_40157);
nand U40388 (N_40388,N_40082,N_40171);
and U40389 (N_40389,N_40241,N_40086);
xnor U40390 (N_40390,N_40008,N_40048);
and U40391 (N_40391,N_40006,N_40189);
and U40392 (N_40392,N_40169,N_40057);
nand U40393 (N_40393,N_40063,N_40231);
or U40394 (N_40394,N_40052,N_40150);
and U40395 (N_40395,N_40096,N_40052);
xnor U40396 (N_40396,N_40119,N_40139);
xor U40397 (N_40397,N_40047,N_40021);
and U40398 (N_40398,N_40207,N_40224);
or U40399 (N_40399,N_40068,N_40135);
nand U40400 (N_40400,N_40094,N_40213);
or U40401 (N_40401,N_40075,N_40042);
nand U40402 (N_40402,N_40233,N_40157);
or U40403 (N_40403,N_40236,N_40083);
and U40404 (N_40404,N_40222,N_40026);
xor U40405 (N_40405,N_40171,N_40137);
or U40406 (N_40406,N_40089,N_40196);
nor U40407 (N_40407,N_40179,N_40188);
or U40408 (N_40408,N_40000,N_40074);
and U40409 (N_40409,N_40243,N_40183);
or U40410 (N_40410,N_40211,N_40048);
nor U40411 (N_40411,N_40171,N_40236);
or U40412 (N_40412,N_40037,N_40157);
nor U40413 (N_40413,N_40177,N_40079);
and U40414 (N_40414,N_40132,N_40227);
nor U40415 (N_40415,N_40055,N_40184);
nand U40416 (N_40416,N_40235,N_40037);
nor U40417 (N_40417,N_40245,N_40017);
nor U40418 (N_40418,N_40116,N_40062);
nor U40419 (N_40419,N_40042,N_40148);
xor U40420 (N_40420,N_40233,N_40014);
or U40421 (N_40421,N_40140,N_40122);
nand U40422 (N_40422,N_40193,N_40121);
nand U40423 (N_40423,N_40238,N_40205);
nand U40424 (N_40424,N_40152,N_40221);
and U40425 (N_40425,N_40174,N_40004);
nor U40426 (N_40426,N_40122,N_40225);
or U40427 (N_40427,N_40205,N_40230);
and U40428 (N_40428,N_40166,N_40117);
or U40429 (N_40429,N_40204,N_40238);
xor U40430 (N_40430,N_40043,N_40158);
and U40431 (N_40431,N_40030,N_40047);
nor U40432 (N_40432,N_40212,N_40185);
and U40433 (N_40433,N_40111,N_40207);
and U40434 (N_40434,N_40057,N_40085);
nor U40435 (N_40435,N_40183,N_40246);
or U40436 (N_40436,N_40038,N_40066);
nor U40437 (N_40437,N_40182,N_40064);
nor U40438 (N_40438,N_40052,N_40188);
nand U40439 (N_40439,N_40222,N_40190);
or U40440 (N_40440,N_40062,N_40225);
or U40441 (N_40441,N_40097,N_40146);
and U40442 (N_40442,N_40219,N_40121);
nand U40443 (N_40443,N_40129,N_40046);
and U40444 (N_40444,N_40103,N_40111);
xor U40445 (N_40445,N_40163,N_40008);
nand U40446 (N_40446,N_40042,N_40072);
nand U40447 (N_40447,N_40182,N_40013);
nand U40448 (N_40448,N_40126,N_40249);
nand U40449 (N_40449,N_40192,N_40068);
xor U40450 (N_40450,N_40044,N_40003);
xor U40451 (N_40451,N_40069,N_40232);
xnor U40452 (N_40452,N_40048,N_40156);
nor U40453 (N_40453,N_40193,N_40076);
xnor U40454 (N_40454,N_40240,N_40138);
or U40455 (N_40455,N_40234,N_40166);
nor U40456 (N_40456,N_40056,N_40180);
nor U40457 (N_40457,N_40155,N_40091);
or U40458 (N_40458,N_40237,N_40050);
or U40459 (N_40459,N_40150,N_40227);
xnor U40460 (N_40460,N_40193,N_40084);
nand U40461 (N_40461,N_40133,N_40100);
or U40462 (N_40462,N_40242,N_40200);
or U40463 (N_40463,N_40134,N_40126);
and U40464 (N_40464,N_40076,N_40065);
xnor U40465 (N_40465,N_40231,N_40050);
or U40466 (N_40466,N_40023,N_40224);
nor U40467 (N_40467,N_40152,N_40149);
xor U40468 (N_40468,N_40246,N_40154);
xnor U40469 (N_40469,N_40051,N_40074);
nor U40470 (N_40470,N_40243,N_40234);
and U40471 (N_40471,N_40067,N_40126);
nand U40472 (N_40472,N_40124,N_40035);
xnor U40473 (N_40473,N_40036,N_40143);
or U40474 (N_40474,N_40244,N_40065);
or U40475 (N_40475,N_40055,N_40179);
xnor U40476 (N_40476,N_40050,N_40022);
or U40477 (N_40477,N_40220,N_40161);
or U40478 (N_40478,N_40041,N_40096);
nand U40479 (N_40479,N_40038,N_40069);
nand U40480 (N_40480,N_40142,N_40145);
or U40481 (N_40481,N_40151,N_40168);
and U40482 (N_40482,N_40199,N_40160);
nand U40483 (N_40483,N_40090,N_40068);
xor U40484 (N_40484,N_40036,N_40061);
xnor U40485 (N_40485,N_40190,N_40206);
and U40486 (N_40486,N_40063,N_40225);
nor U40487 (N_40487,N_40040,N_40115);
and U40488 (N_40488,N_40077,N_40248);
or U40489 (N_40489,N_40249,N_40196);
and U40490 (N_40490,N_40175,N_40001);
and U40491 (N_40491,N_40078,N_40052);
and U40492 (N_40492,N_40207,N_40007);
or U40493 (N_40493,N_40052,N_40223);
and U40494 (N_40494,N_40212,N_40135);
nand U40495 (N_40495,N_40071,N_40028);
xor U40496 (N_40496,N_40046,N_40016);
nor U40497 (N_40497,N_40225,N_40045);
nand U40498 (N_40498,N_40071,N_40216);
nor U40499 (N_40499,N_40173,N_40171);
nor U40500 (N_40500,N_40394,N_40293);
nor U40501 (N_40501,N_40262,N_40473);
nor U40502 (N_40502,N_40375,N_40315);
and U40503 (N_40503,N_40359,N_40435);
and U40504 (N_40504,N_40344,N_40499);
nor U40505 (N_40505,N_40379,N_40498);
or U40506 (N_40506,N_40430,N_40322);
or U40507 (N_40507,N_40309,N_40376);
and U40508 (N_40508,N_40405,N_40366);
xor U40509 (N_40509,N_40440,N_40288);
xnor U40510 (N_40510,N_40373,N_40357);
and U40511 (N_40511,N_40341,N_40462);
and U40512 (N_40512,N_40392,N_40444);
and U40513 (N_40513,N_40459,N_40370);
nand U40514 (N_40514,N_40419,N_40424);
and U40515 (N_40515,N_40338,N_40453);
and U40516 (N_40516,N_40330,N_40377);
and U40517 (N_40517,N_40305,N_40445);
or U40518 (N_40518,N_40490,N_40294);
xnor U40519 (N_40519,N_40439,N_40464);
and U40520 (N_40520,N_40275,N_40354);
or U40521 (N_40521,N_40396,N_40329);
and U40522 (N_40522,N_40280,N_40421);
and U40523 (N_40523,N_40401,N_40496);
and U40524 (N_40524,N_40428,N_40446);
or U40525 (N_40525,N_40284,N_40467);
xor U40526 (N_40526,N_40449,N_40402);
or U40527 (N_40527,N_40420,N_40255);
nor U40528 (N_40528,N_40272,N_40455);
nand U40529 (N_40529,N_40450,N_40398);
nor U40530 (N_40530,N_40438,N_40426);
xor U40531 (N_40531,N_40381,N_40476);
xnor U40532 (N_40532,N_40451,N_40372);
nand U40533 (N_40533,N_40253,N_40340);
nand U40534 (N_40534,N_40346,N_40486);
nor U40535 (N_40535,N_40335,N_40468);
nor U40536 (N_40536,N_40312,N_40395);
and U40537 (N_40537,N_40321,N_40427);
or U40538 (N_40538,N_40286,N_40478);
and U40539 (N_40539,N_40360,N_40256);
xnor U40540 (N_40540,N_40480,N_40349);
and U40541 (N_40541,N_40304,N_40334);
nand U40542 (N_40542,N_40443,N_40271);
xor U40543 (N_40543,N_40448,N_40399);
xor U40544 (N_40544,N_40415,N_40432);
xor U40545 (N_40545,N_40265,N_40434);
or U40546 (N_40546,N_40386,N_40342);
nand U40547 (N_40547,N_40447,N_40289);
nand U40548 (N_40548,N_40492,N_40316);
and U40549 (N_40549,N_40318,N_40298);
or U40550 (N_40550,N_40482,N_40264);
nand U40551 (N_40551,N_40308,N_40484);
or U40552 (N_40552,N_40303,N_40472);
nand U40553 (N_40553,N_40385,N_40259);
xor U40554 (N_40554,N_40413,N_40317);
or U40555 (N_40555,N_40358,N_40350);
and U40556 (N_40556,N_40274,N_40367);
nor U40557 (N_40557,N_40362,N_40347);
nand U40558 (N_40558,N_40311,N_40404);
nand U40559 (N_40559,N_40493,N_40485);
and U40560 (N_40560,N_40387,N_40260);
nand U40561 (N_40561,N_40418,N_40417);
xnor U40562 (N_40562,N_40261,N_40465);
and U40563 (N_40563,N_40361,N_40300);
or U40564 (N_40564,N_40380,N_40412);
nand U40565 (N_40565,N_40277,N_40252);
or U40566 (N_40566,N_40287,N_40295);
or U40567 (N_40567,N_40283,N_40273);
xnor U40568 (N_40568,N_40251,N_40461);
or U40569 (N_40569,N_40296,N_40364);
nor U40570 (N_40570,N_40269,N_40302);
xnor U40571 (N_40571,N_40469,N_40353);
and U40572 (N_40572,N_40371,N_40278);
nor U40573 (N_40573,N_40352,N_40475);
nand U40574 (N_40574,N_40481,N_40429);
nand U40575 (N_40575,N_40285,N_40281);
nor U40576 (N_40576,N_40355,N_40414);
nor U40577 (N_40577,N_40423,N_40437);
xor U40578 (N_40578,N_40491,N_40407);
nand U40579 (N_40579,N_40483,N_40254);
nor U40580 (N_40580,N_40365,N_40479);
nor U40581 (N_40581,N_40408,N_40487);
or U40582 (N_40582,N_40291,N_40314);
and U40583 (N_40583,N_40337,N_40416);
or U40584 (N_40584,N_40452,N_40471);
xor U40585 (N_40585,N_40257,N_40441);
and U40586 (N_40586,N_40494,N_40400);
and U40587 (N_40587,N_40422,N_40489);
xor U40588 (N_40588,N_40292,N_40333);
nor U40589 (N_40589,N_40299,N_40301);
xor U40590 (N_40590,N_40266,N_40282);
nor U40591 (N_40591,N_40495,N_40327);
and U40592 (N_40592,N_40369,N_40290);
nand U40593 (N_40593,N_40391,N_40258);
and U40594 (N_40594,N_40457,N_40409);
nand U40595 (N_40595,N_40463,N_40356);
nor U40596 (N_40596,N_40276,N_40307);
nor U40597 (N_40597,N_40332,N_40488);
or U40598 (N_40598,N_40384,N_40390);
nor U40599 (N_40599,N_40319,N_40368);
xor U40600 (N_40600,N_40324,N_40363);
or U40601 (N_40601,N_40406,N_40460);
and U40602 (N_40602,N_40425,N_40397);
nand U40603 (N_40603,N_40310,N_40383);
or U40604 (N_40604,N_40326,N_40466);
nor U40605 (N_40605,N_40306,N_40270);
nand U40606 (N_40606,N_40339,N_40343);
or U40607 (N_40607,N_40313,N_40470);
nor U40608 (N_40608,N_40403,N_40456);
and U40609 (N_40609,N_40268,N_40477);
xor U40610 (N_40610,N_40411,N_40279);
nand U40611 (N_40611,N_40454,N_40378);
and U40612 (N_40612,N_40267,N_40436);
nand U40613 (N_40613,N_40431,N_40393);
xnor U40614 (N_40614,N_40250,N_40345);
and U40615 (N_40615,N_40297,N_40328);
nand U40616 (N_40616,N_40410,N_40389);
xnor U40617 (N_40617,N_40325,N_40331);
nand U40618 (N_40618,N_40336,N_40458);
nor U40619 (N_40619,N_40323,N_40320);
and U40620 (N_40620,N_40442,N_40348);
nand U40621 (N_40621,N_40382,N_40433);
or U40622 (N_40622,N_40388,N_40497);
and U40623 (N_40623,N_40374,N_40263);
xor U40624 (N_40624,N_40474,N_40351);
or U40625 (N_40625,N_40442,N_40445);
or U40626 (N_40626,N_40473,N_40389);
nand U40627 (N_40627,N_40420,N_40262);
xnor U40628 (N_40628,N_40339,N_40261);
nor U40629 (N_40629,N_40324,N_40307);
nand U40630 (N_40630,N_40333,N_40434);
nor U40631 (N_40631,N_40293,N_40285);
or U40632 (N_40632,N_40459,N_40471);
or U40633 (N_40633,N_40270,N_40455);
nor U40634 (N_40634,N_40404,N_40474);
nand U40635 (N_40635,N_40306,N_40445);
nor U40636 (N_40636,N_40334,N_40467);
or U40637 (N_40637,N_40434,N_40352);
nand U40638 (N_40638,N_40408,N_40370);
nor U40639 (N_40639,N_40468,N_40457);
or U40640 (N_40640,N_40327,N_40440);
and U40641 (N_40641,N_40407,N_40433);
nand U40642 (N_40642,N_40493,N_40318);
and U40643 (N_40643,N_40418,N_40295);
or U40644 (N_40644,N_40346,N_40493);
xor U40645 (N_40645,N_40352,N_40292);
nand U40646 (N_40646,N_40389,N_40427);
or U40647 (N_40647,N_40256,N_40422);
and U40648 (N_40648,N_40319,N_40350);
nor U40649 (N_40649,N_40268,N_40462);
nor U40650 (N_40650,N_40329,N_40258);
nand U40651 (N_40651,N_40392,N_40484);
or U40652 (N_40652,N_40267,N_40331);
nand U40653 (N_40653,N_40366,N_40323);
or U40654 (N_40654,N_40452,N_40316);
nand U40655 (N_40655,N_40287,N_40489);
nand U40656 (N_40656,N_40341,N_40286);
xnor U40657 (N_40657,N_40405,N_40302);
nor U40658 (N_40658,N_40487,N_40429);
or U40659 (N_40659,N_40443,N_40401);
and U40660 (N_40660,N_40309,N_40367);
nor U40661 (N_40661,N_40303,N_40478);
nor U40662 (N_40662,N_40305,N_40392);
xor U40663 (N_40663,N_40462,N_40458);
xnor U40664 (N_40664,N_40383,N_40453);
and U40665 (N_40665,N_40258,N_40268);
nor U40666 (N_40666,N_40436,N_40272);
nor U40667 (N_40667,N_40360,N_40432);
xnor U40668 (N_40668,N_40484,N_40334);
nor U40669 (N_40669,N_40489,N_40391);
nand U40670 (N_40670,N_40257,N_40390);
nor U40671 (N_40671,N_40490,N_40418);
and U40672 (N_40672,N_40251,N_40291);
xnor U40673 (N_40673,N_40464,N_40385);
or U40674 (N_40674,N_40287,N_40305);
and U40675 (N_40675,N_40432,N_40451);
xnor U40676 (N_40676,N_40385,N_40374);
xnor U40677 (N_40677,N_40393,N_40324);
nand U40678 (N_40678,N_40285,N_40387);
xor U40679 (N_40679,N_40279,N_40278);
and U40680 (N_40680,N_40352,N_40317);
nand U40681 (N_40681,N_40279,N_40448);
and U40682 (N_40682,N_40481,N_40427);
and U40683 (N_40683,N_40403,N_40484);
xnor U40684 (N_40684,N_40330,N_40392);
xor U40685 (N_40685,N_40456,N_40291);
xnor U40686 (N_40686,N_40484,N_40349);
or U40687 (N_40687,N_40419,N_40267);
xnor U40688 (N_40688,N_40258,N_40322);
nor U40689 (N_40689,N_40317,N_40452);
and U40690 (N_40690,N_40386,N_40318);
xor U40691 (N_40691,N_40480,N_40292);
nor U40692 (N_40692,N_40271,N_40417);
or U40693 (N_40693,N_40464,N_40353);
nand U40694 (N_40694,N_40362,N_40497);
and U40695 (N_40695,N_40379,N_40360);
and U40696 (N_40696,N_40296,N_40286);
nor U40697 (N_40697,N_40423,N_40492);
nand U40698 (N_40698,N_40474,N_40370);
or U40699 (N_40699,N_40360,N_40437);
and U40700 (N_40700,N_40466,N_40484);
xnor U40701 (N_40701,N_40255,N_40326);
and U40702 (N_40702,N_40496,N_40260);
or U40703 (N_40703,N_40456,N_40343);
xnor U40704 (N_40704,N_40448,N_40447);
or U40705 (N_40705,N_40373,N_40317);
nor U40706 (N_40706,N_40271,N_40390);
nor U40707 (N_40707,N_40404,N_40459);
nand U40708 (N_40708,N_40285,N_40272);
xor U40709 (N_40709,N_40406,N_40285);
nand U40710 (N_40710,N_40498,N_40352);
nor U40711 (N_40711,N_40419,N_40371);
or U40712 (N_40712,N_40413,N_40340);
nand U40713 (N_40713,N_40261,N_40266);
nor U40714 (N_40714,N_40358,N_40433);
or U40715 (N_40715,N_40490,N_40272);
nand U40716 (N_40716,N_40288,N_40308);
and U40717 (N_40717,N_40361,N_40260);
xnor U40718 (N_40718,N_40297,N_40261);
nand U40719 (N_40719,N_40268,N_40473);
xor U40720 (N_40720,N_40296,N_40362);
and U40721 (N_40721,N_40289,N_40450);
nand U40722 (N_40722,N_40395,N_40409);
or U40723 (N_40723,N_40313,N_40432);
nor U40724 (N_40724,N_40250,N_40445);
xor U40725 (N_40725,N_40390,N_40400);
or U40726 (N_40726,N_40302,N_40448);
nor U40727 (N_40727,N_40254,N_40402);
nand U40728 (N_40728,N_40256,N_40355);
xor U40729 (N_40729,N_40460,N_40483);
nor U40730 (N_40730,N_40478,N_40360);
or U40731 (N_40731,N_40461,N_40456);
and U40732 (N_40732,N_40320,N_40416);
nor U40733 (N_40733,N_40455,N_40462);
and U40734 (N_40734,N_40367,N_40324);
or U40735 (N_40735,N_40454,N_40483);
nor U40736 (N_40736,N_40383,N_40324);
and U40737 (N_40737,N_40257,N_40450);
and U40738 (N_40738,N_40337,N_40492);
and U40739 (N_40739,N_40302,N_40281);
nand U40740 (N_40740,N_40278,N_40467);
or U40741 (N_40741,N_40463,N_40454);
xor U40742 (N_40742,N_40388,N_40337);
or U40743 (N_40743,N_40345,N_40390);
nand U40744 (N_40744,N_40282,N_40255);
and U40745 (N_40745,N_40341,N_40459);
nand U40746 (N_40746,N_40430,N_40425);
nand U40747 (N_40747,N_40402,N_40454);
nand U40748 (N_40748,N_40295,N_40428);
xnor U40749 (N_40749,N_40278,N_40475);
nand U40750 (N_40750,N_40687,N_40560);
and U40751 (N_40751,N_40514,N_40575);
xnor U40752 (N_40752,N_40617,N_40643);
nand U40753 (N_40753,N_40573,N_40658);
nor U40754 (N_40754,N_40539,N_40608);
xnor U40755 (N_40755,N_40686,N_40599);
nand U40756 (N_40756,N_40728,N_40741);
nor U40757 (N_40757,N_40579,N_40586);
and U40758 (N_40758,N_40559,N_40601);
nor U40759 (N_40759,N_40562,N_40600);
nand U40760 (N_40760,N_40564,N_40739);
xnor U40761 (N_40761,N_40665,N_40696);
xnor U40762 (N_40762,N_40533,N_40558);
xor U40763 (N_40763,N_40590,N_40509);
xnor U40764 (N_40764,N_40522,N_40611);
or U40765 (N_40765,N_40729,N_40667);
or U40766 (N_40766,N_40519,N_40688);
nand U40767 (N_40767,N_40661,N_40527);
nand U40768 (N_40768,N_40660,N_40505);
nand U40769 (N_40769,N_40636,N_40653);
and U40770 (N_40770,N_40715,N_40528);
or U40771 (N_40771,N_40689,N_40535);
nand U40772 (N_40772,N_40543,N_40627);
and U40773 (N_40773,N_40690,N_40638);
and U40774 (N_40774,N_40708,N_40721);
nor U40775 (N_40775,N_40656,N_40662);
nand U40776 (N_40776,N_40628,N_40532);
and U40777 (N_40777,N_40531,N_40645);
and U40778 (N_40778,N_40518,N_40577);
nor U40779 (N_40779,N_40582,N_40706);
nor U40780 (N_40780,N_40571,N_40530);
or U40781 (N_40781,N_40591,N_40675);
xnor U40782 (N_40782,N_40712,N_40583);
or U40783 (N_40783,N_40644,N_40730);
or U40784 (N_40784,N_40733,N_40674);
xnor U40785 (N_40785,N_40517,N_40609);
xor U40786 (N_40786,N_40618,N_40742);
xor U40787 (N_40787,N_40673,N_40516);
and U40788 (N_40788,N_40620,N_40719);
nand U40789 (N_40789,N_40574,N_40705);
and U40790 (N_40790,N_40631,N_40717);
nand U40791 (N_40791,N_40698,N_40589);
xnor U40792 (N_40792,N_40671,N_40624);
and U40793 (N_40793,N_40576,N_40666);
nor U40794 (N_40794,N_40536,N_40614);
or U40795 (N_40795,N_40670,N_40637);
or U40796 (N_40796,N_40580,N_40693);
nor U40797 (N_40797,N_40735,N_40707);
nor U40798 (N_40798,N_40743,N_40585);
nor U40799 (N_40799,N_40548,N_40597);
nor U40800 (N_40800,N_40625,N_40529);
nand U40801 (N_40801,N_40727,N_40551);
and U40802 (N_40802,N_40557,N_40545);
nor U40803 (N_40803,N_40595,N_40596);
nand U40804 (N_40804,N_40642,N_40737);
nor U40805 (N_40805,N_40736,N_40732);
and U40806 (N_40806,N_40738,N_40731);
and U40807 (N_40807,N_40744,N_40605);
xnor U40808 (N_40808,N_40646,N_40503);
nand U40809 (N_40809,N_40534,N_40629);
nor U40810 (N_40810,N_40507,N_40649);
nor U40811 (N_40811,N_40659,N_40568);
and U40812 (N_40812,N_40578,N_40635);
nor U40813 (N_40813,N_40526,N_40648);
nor U40814 (N_40814,N_40594,N_40672);
nand U40815 (N_40815,N_40722,N_40504);
xnor U40816 (N_40816,N_40512,N_40550);
nand U40817 (N_40817,N_40544,N_40734);
or U40818 (N_40818,N_40540,N_40565);
and U40819 (N_40819,N_40684,N_40513);
nand U40820 (N_40820,N_40547,N_40682);
nand U40821 (N_40821,N_40640,N_40555);
nor U40822 (N_40822,N_40634,N_40570);
and U40823 (N_40823,N_40724,N_40593);
xor U40824 (N_40824,N_40606,N_40701);
nand U40825 (N_40825,N_40678,N_40553);
and U40826 (N_40826,N_40740,N_40704);
or U40827 (N_40827,N_40702,N_40521);
and U40828 (N_40828,N_40537,N_40679);
xor U40829 (N_40829,N_40616,N_40726);
nand U40830 (N_40830,N_40581,N_40538);
nand U40831 (N_40831,N_40541,N_40748);
nor U40832 (N_40832,N_40663,N_40619);
or U40833 (N_40833,N_40510,N_40716);
nand U40834 (N_40834,N_40718,N_40676);
xor U40835 (N_40835,N_40587,N_40652);
or U40836 (N_40836,N_40703,N_40699);
and U40837 (N_40837,N_40598,N_40655);
nor U40838 (N_40838,N_40694,N_40723);
nand U40839 (N_40839,N_40561,N_40592);
nand U40840 (N_40840,N_40588,N_40552);
nor U40841 (N_40841,N_40668,N_40691);
xnor U40842 (N_40842,N_40502,N_40714);
xnor U40843 (N_40843,N_40612,N_40622);
nand U40844 (N_40844,N_40711,N_40523);
and U40845 (N_40845,N_40626,N_40685);
nor U40846 (N_40846,N_40566,N_40603);
nand U40847 (N_40847,N_40615,N_40669);
or U40848 (N_40848,N_40695,N_40713);
nor U40849 (N_40849,N_40633,N_40680);
and U40850 (N_40850,N_40610,N_40650);
xnor U40851 (N_40851,N_40524,N_40654);
nand U40852 (N_40852,N_40623,N_40720);
xnor U40853 (N_40853,N_40709,N_40584);
and U40854 (N_40854,N_40500,N_40692);
or U40855 (N_40855,N_40613,N_40563);
nand U40856 (N_40856,N_40664,N_40697);
and U40857 (N_40857,N_40681,N_40630);
and U40858 (N_40858,N_40700,N_40639);
and U40859 (N_40859,N_40657,N_40683);
nand U40860 (N_40860,N_40525,N_40569);
nor U40861 (N_40861,N_40542,N_40506);
nand U40862 (N_40862,N_40501,N_40572);
nand U40863 (N_40863,N_40632,N_40677);
or U40864 (N_40864,N_40604,N_40567);
nor U40865 (N_40865,N_40508,N_40641);
nor U40866 (N_40866,N_40515,N_40511);
xnor U40867 (N_40867,N_40520,N_40549);
or U40868 (N_40868,N_40647,N_40747);
or U40869 (N_40869,N_40546,N_40651);
nand U40870 (N_40870,N_40607,N_40602);
and U40871 (N_40871,N_40725,N_40556);
nand U40872 (N_40872,N_40554,N_40749);
nor U40873 (N_40873,N_40710,N_40621);
nand U40874 (N_40874,N_40746,N_40745);
nor U40875 (N_40875,N_40666,N_40749);
and U40876 (N_40876,N_40714,N_40516);
or U40877 (N_40877,N_40746,N_40702);
xor U40878 (N_40878,N_40502,N_40677);
xnor U40879 (N_40879,N_40673,N_40628);
xnor U40880 (N_40880,N_40692,N_40602);
and U40881 (N_40881,N_40575,N_40707);
and U40882 (N_40882,N_40520,N_40544);
xor U40883 (N_40883,N_40588,N_40613);
and U40884 (N_40884,N_40581,N_40596);
xnor U40885 (N_40885,N_40575,N_40704);
or U40886 (N_40886,N_40618,N_40738);
nor U40887 (N_40887,N_40574,N_40728);
or U40888 (N_40888,N_40632,N_40523);
or U40889 (N_40889,N_40583,N_40723);
and U40890 (N_40890,N_40748,N_40699);
xnor U40891 (N_40891,N_40738,N_40643);
nand U40892 (N_40892,N_40725,N_40718);
xnor U40893 (N_40893,N_40575,N_40661);
nand U40894 (N_40894,N_40665,N_40670);
nor U40895 (N_40895,N_40503,N_40608);
xor U40896 (N_40896,N_40606,N_40555);
xor U40897 (N_40897,N_40640,N_40713);
and U40898 (N_40898,N_40698,N_40627);
and U40899 (N_40899,N_40634,N_40571);
or U40900 (N_40900,N_40603,N_40682);
nor U40901 (N_40901,N_40667,N_40575);
and U40902 (N_40902,N_40748,N_40508);
xor U40903 (N_40903,N_40571,N_40616);
or U40904 (N_40904,N_40654,N_40606);
or U40905 (N_40905,N_40532,N_40549);
nor U40906 (N_40906,N_40643,N_40718);
or U40907 (N_40907,N_40538,N_40532);
nor U40908 (N_40908,N_40730,N_40647);
or U40909 (N_40909,N_40517,N_40693);
and U40910 (N_40910,N_40673,N_40534);
nor U40911 (N_40911,N_40725,N_40668);
nor U40912 (N_40912,N_40701,N_40609);
xor U40913 (N_40913,N_40608,N_40693);
xnor U40914 (N_40914,N_40559,N_40678);
nand U40915 (N_40915,N_40704,N_40727);
nand U40916 (N_40916,N_40516,N_40615);
nand U40917 (N_40917,N_40658,N_40523);
xnor U40918 (N_40918,N_40726,N_40579);
xnor U40919 (N_40919,N_40505,N_40533);
xnor U40920 (N_40920,N_40583,N_40599);
xnor U40921 (N_40921,N_40552,N_40529);
xor U40922 (N_40922,N_40702,N_40651);
nor U40923 (N_40923,N_40512,N_40634);
nand U40924 (N_40924,N_40603,N_40673);
xor U40925 (N_40925,N_40679,N_40517);
xnor U40926 (N_40926,N_40643,N_40727);
nor U40927 (N_40927,N_40521,N_40689);
nor U40928 (N_40928,N_40502,N_40621);
nor U40929 (N_40929,N_40560,N_40637);
xnor U40930 (N_40930,N_40712,N_40720);
and U40931 (N_40931,N_40601,N_40608);
nand U40932 (N_40932,N_40500,N_40510);
nand U40933 (N_40933,N_40731,N_40613);
nor U40934 (N_40934,N_40579,N_40544);
and U40935 (N_40935,N_40698,N_40643);
and U40936 (N_40936,N_40688,N_40542);
nor U40937 (N_40937,N_40670,N_40721);
nor U40938 (N_40938,N_40716,N_40500);
and U40939 (N_40939,N_40561,N_40720);
or U40940 (N_40940,N_40569,N_40614);
and U40941 (N_40941,N_40622,N_40557);
nand U40942 (N_40942,N_40597,N_40559);
or U40943 (N_40943,N_40646,N_40732);
xnor U40944 (N_40944,N_40560,N_40672);
nand U40945 (N_40945,N_40501,N_40510);
or U40946 (N_40946,N_40580,N_40717);
nand U40947 (N_40947,N_40591,N_40575);
or U40948 (N_40948,N_40546,N_40681);
or U40949 (N_40949,N_40616,N_40522);
or U40950 (N_40950,N_40661,N_40706);
or U40951 (N_40951,N_40598,N_40582);
xnor U40952 (N_40952,N_40639,N_40674);
or U40953 (N_40953,N_40631,N_40527);
nor U40954 (N_40954,N_40589,N_40681);
xnor U40955 (N_40955,N_40701,N_40677);
xor U40956 (N_40956,N_40543,N_40595);
nor U40957 (N_40957,N_40531,N_40686);
nand U40958 (N_40958,N_40500,N_40515);
or U40959 (N_40959,N_40554,N_40669);
nor U40960 (N_40960,N_40548,N_40585);
and U40961 (N_40961,N_40714,N_40639);
nand U40962 (N_40962,N_40662,N_40727);
or U40963 (N_40963,N_40741,N_40628);
nand U40964 (N_40964,N_40608,N_40535);
and U40965 (N_40965,N_40593,N_40565);
xor U40966 (N_40966,N_40669,N_40520);
nor U40967 (N_40967,N_40592,N_40674);
nor U40968 (N_40968,N_40620,N_40669);
and U40969 (N_40969,N_40693,N_40653);
xnor U40970 (N_40970,N_40610,N_40627);
nor U40971 (N_40971,N_40607,N_40676);
nor U40972 (N_40972,N_40582,N_40609);
nor U40973 (N_40973,N_40627,N_40535);
nand U40974 (N_40974,N_40531,N_40507);
and U40975 (N_40975,N_40564,N_40727);
nand U40976 (N_40976,N_40608,N_40521);
and U40977 (N_40977,N_40577,N_40676);
nand U40978 (N_40978,N_40651,N_40689);
and U40979 (N_40979,N_40514,N_40620);
xor U40980 (N_40980,N_40584,N_40599);
nor U40981 (N_40981,N_40624,N_40743);
xor U40982 (N_40982,N_40715,N_40682);
and U40983 (N_40983,N_40517,N_40539);
and U40984 (N_40984,N_40650,N_40729);
nand U40985 (N_40985,N_40528,N_40601);
xor U40986 (N_40986,N_40578,N_40551);
nor U40987 (N_40987,N_40704,N_40633);
nor U40988 (N_40988,N_40664,N_40720);
nor U40989 (N_40989,N_40594,N_40603);
nor U40990 (N_40990,N_40555,N_40530);
or U40991 (N_40991,N_40744,N_40541);
or U40992 (N_40992,N_40579,N_40694);
nand U40993 (N_40993,N_40604,N_40574);
nand U40994 (N_40994,N_40707,N_40669);
and U40995 (N_40995,N_40528,N_40724);
xnor U40996 (N_40996,N_40683,N_40505);
or U40997 (N_40997,N_40594,N_40747);
xnor U40998 (N_40998,N_40592,N_40582);
xnor U40999 (N_40999,N_40703,N_40578);
and U41000 (N_41000,N_40984,N_40940);
nand U41001 (N_41001,N_40957,N_40985);
and U41002 (N_41002,N_40762,N_40885);
and U41003 (N_41003,N_40859,N_40939);
xor U41004 (N_41004,N_40979,N_40818);
nand U41005 (N_41005,N_40944,N_40848);
and U41006 (N_41006,N_40910,N_40993);
and U41007 (N_41007,N_40888,N_40887);
xnor U41008 (N_41008,N_40803,N_40788);
and U41009 (N_41009,N_40778,N_40856);
xor U41010 (N_41010,N_40750,N_40982);
and U41011 (N_41011,N_40849,N_40896);
or U41012 (N_41012,N_40908,N_40805);
xor U41013 (N_41013,N_40995,N_40783);
nor U41014 (N_41014,N_40964,N_40757);
or U41015 (N_41015,N_40784,N_40855);
or U41016 (N_41016,N_40980,N_40947);
or U41017 (N_41017,N_40821,N_40771);
and U41018 (N_41018,N_40862,N_40827);
nor U41019 (N_41019,N_40925,N_40937);
xnor U41020 (N_41020,N_40852,N_40988);
nor U41021 (N_41021,N_40917,N_40945);
or U41022 (N_41022,N_40973,N_40869);
xor U41023 (N_41023,N_40822,N_40971);
or U41024 (N_41024,N_40898,N_40765);
nand U41025 (N_41025,N_40758,N_40899);
and U41026 (N_41026,N_40930,N_40923);
or U41027 (N_41027,N_40968,N_40934);
or U41028 (N_41028,N_40851,N_40867);
xor U41029 (N_41029,N_40812,N_40839);
or U41030 (N_41030,N_40897,N_40967);
and U41031 (N_41031,N_40933,N_40768);
nand U41032 (N_41032,N_40808,N_40965);
and U41033 (N_41033,N_40951,N_40953);
or U41034 (N_41034,N_40799,N_40832);
or U41035 (N_41035,N_40916,N_40882);
nor U41036 (N_41036,N_40789,N_40817);
xnor U41037 (N_41037,N_40935,N_40936);
nor U41038 (N_41038,N_40753,N_40785);
xnor U41039 (N_41039,N_40797,N_40959);
nor U41040 (N_41040,N_40977,N_40807);
or U41041 (N_41041,N_40786,N_40919);
xor U41042 (N_41042,N_40902,N_40779);
nand U41043 (N_41043,N_40870,N_40764);
and U41044 (N_41044,N_40837,N_40858);
nand U41045 (N_41045,N_40826,N_40836);
nand U41046 (N_41046,N_40920,N_40997);
and U41047 (N_41047,N_40850,N_40834);
xnor U41048 (N_41048,N_40815,N_40884);
and U41049 (N_41049,N_40912,N_40877);
xnor U41050 (N_41050,N_40796,N_40791);
nor U41051 (N_41051,N_40811,N_40905);
and U41052 (N_41052,N_40751,N_40806);
nor U41053 (N_41053,N_40857,N_40861);
xnor U41054 (N_41054,N_40831,N_40976);
and U41055 (N_41055,N_40886,N_40820);
nor U41056 (N_41056,N_40915,N_40865);
xnor U41057 (N_41057,N_40775,N_40893);
nor U41058 (N_41058,N_40838,N_40798);
nand U41059 (N_41059,N_40847,N_40983);
and U41060 (N_41060,N_40754,N_40890);
nand U41061 (N_41061,N_40879,N_40792);
nor U41062 (N_41062,N_40814,N_40880);
or U41063 (N_41063,N_40780,N_40952);
xor U41064 (N_41064,N_40904,N_40990);
or U41065 (N_41065,N_40795,N_40755);
and U41066 (N_41066,N_40813,N_40840);
nor U41067 (N_41067,N_40883,N_40843);
nand U41068 (N_41068,N_40906,N_40978);
xor U41069 (N_41069,N_40801,N_40863);
xor U41070 (N_41070,N_40829,N_40866);
and U41071 (N_41071,N_40874,N_40854);
and U41072 (N_41072,N_40963,N_40891);
nor U41073 (N_41073,N_40860,N_40956);
and U41074 (N_41074,N_40961,N_40932);
nand U41075 (N_41075,N_40986,N_40761);
or U41076 (N_41076,N_40844,N_40769);
nor U41077 (N_41077,N_40872,N_40931);
xnor U41078 (N_41078,N_40966,N_40846);
or U41079 (N_41079,N_40929,N_40770);
and U41080 (N_41080,N_40752,N_40763);
xor U41081 (N_41081,N_40835,N_40955);
and U41082 (N_41082,N_40772,N_40974);
and U41083 (N_41083,N_40777,N_40790);
or U41084 (N_41084,N_40950,N_40819);
nand U41085 (N_41085,N_40800,N_40946);
or U41086 (N_41086,N_40913,N_40901);
xnor U41087 (N_41087,N_40830,N_40900);
or U41088 (N_41088,N_40810,N_40975);
nor U41089 (N_41089,N_40903,N_40926);
nor U41090 (N_41090,N_40895,N_40760);
nor U41091 (N_41091,N_40873,N_40864);
or U41092 (N_41092,N_40845,N_40991);
or U41093 (N_41093,N_40938,N_40962);
or U41094 (N_41094,N_40868,N_40871);
xor U41095 (N_41095,N_40999,N_40960);
xnor U41096 (N_41096,N_40894,N_40766);
and U41097 (N_41097,N_40881,N_40756);
or U41098 (N_41098,N_40972,N_40948);
nand U41099 (N_41099,N_40781,N_40809);
nand U41100 (N_41100,N_40774,N_40816);
nand U41101 (N_41101,N_40878,N_40928);
or U41102 (N_41102,N_40841,N_40892);
or U41103 (N_41103,N_40992,N_40927);
and U41104 (N_41104,N_40958,N_40994);
or U41105 (N_41105,N_40828,N_40793);
nor U41106 (N_41106,N_40907,N_40876);
xor U41107 (N_41107,N_40833,N_40987);
nor U41108 (N_41108,N_40941,N_40918);
xor U41109 (N_41109,N_40773,N_40759);
xor U41110 (N_41110,N_40942,N_40823);
nor U41111 (N_41111,N_40922,N_40970);
and U41112 (N_41112,N_40981,N_40875);
nor U41113 (N_41113,N_40889,N_40911);
nand U41114 (N_41114,N_40842,N_40782);
nor U41115 (N_41115,N_40996,N_40954);
and U41116 (N_41116,N_40776,N_40998);
or U41117 (N_41117,N_40921,N_40804);
and U41118 (N_41118,N_40914,N_40853);
nor U41119 (N_41119,N_40909,N_40943);
xnor U41120 (N_41120,N_40787,N_40802);
nor U41121 (N_41121,N_40989,N_40824);
and U41122 (N_41122,N_40825,N_40949);
nor U41123 (N_41123,N_40767,N_40794);
nor U41124 (N_41124,N_40924,N_40969);
xor U41125 (N_41125,N_40795,N_40879);
nor U41126 (N_41126,N_40938,N_40869);
nand U41127 (N_41127,N_40933,N_40897);
or U41128 (N_41128,N_40761,N_40759);
nand U41129 (N_41129,N_40790,N_40808);
nand U41130 (N_41130,N_40896,N_40783);
nand U41131 (N_41131,N_40763,N_40841);
nand U41132 (N_41132,N_40993,N_40812);
and U41133 (N_41133,N_40891,N_40807);
xor U41134 (N_41134,N_40892,N_40815);
or U41135 (N_41135,N_40777,N_40889);
xor U41136 (N_41136,N_40999,N_40835);
nand U41137 (N_41137,N_40831,N_40826);
and U41138 (N_41138,N_40980,N_40776);
xnor U41139 (N_41139,N_40847,N_40890);
nor U41140 (N_41140,N_40992,N_40792);
or U41141 (N_41141,N_40756,N_40754);
nand U41142 (N_41142,N_40857,N_40845);
or U41143 (N_41143,N_40830,N_40852);
xor U41144 (N_41144,N_40767,N_40896);
nand U41145 (N_41145,N_40756,N_40942);
xor U41146 (N_41146,N_40854,N_40910);
xor U41147 (N_41147,N_40993,N_40901);
or U41148 (N_41148,N_40823,N_40902);
xor U41149 (N_41149,N_40850,N_40802);
nand U41150 (N_41150,N_40838,N_40875);
nor U41151 (N_41151,N_40897,N_40966);
and U41152 (N_41152,N_40891,N_40832);
and U41153 (N_41153,N_40923,N_40960);
nand U41154 (N_41154,N_40793,N_40995);
nor U41155 (N_41155,N_40951,N_40752);
and U41156 (N_41156,N_40909,N_40753);
nand U41157 (N_41157,N_40815,N_40836);
xnor U41158 (N_41158,N_40826,N_40837);
and U41159 (N_41159,N_40851,N_40904);
and U41160 (N_41160,N_40805,N_40838);
xor U41161 (N_41161,N_40928,N_40788);
and U41162 (N_41162,N_40866,N_40898);
nand U41163 (N_41163,N_40891,N_40775);
nor U41164 (N_41164,N_40841,N_40935);
xnor U41165 (N_41165,N_40964,N_40817);
nor U41166 (N_41166,N_40796,N_40931);
xor U41167 (N_41167,N_40752,N_40809);
or U41168 (N_41168,N_40844,N_40755);
nand U41169 (N_41169,N_40756,N_40770);
xnor U41170 (N_41170,N_40920,N_40790);
or U41171 (N_41171,N_40766,N_40797);
xnor U41172 (N_41172,N_40934,N_40905);
or U41173 (N_41173,N_40874,N_40948);
xor U41174 (N_41174,N_40860,N_40755);
or U41175 (N_41175,N_40885,N_40939);
nor U41176 (N_41176,N_40860,N_40927);
or U41177 (N_41177,N_40942,N_40761);
or U41178 (N_41178,N_40810,N_40781);
or U41179 (N_41179,N_40850,N_40894);
nor U41180 (N_41180,N_40957,N_40893);
and U41181 (N_41181,N_40876,N_40766);
nor U41182 (N_41182,N_40901,N_40857);
xor U41183 (N_41183,N_40888,N_40819);
nor U41184 (N_41184,N_40821,N_40895);
nor U41185 (N_41185,N_40943,N_40753);
or U41186 (N_41186,N_40800,N_40982);
or U41187 (N_41187,N_40895,N_40993);
or U41188 (N_41188,N_40824,N_40976);
or U41189 (N_41189,N_40839,N_40758);
nor U41190 (N_41190,N_40990,N_40913);
or U41191 (N_41191,N_40828,N_40895);
and U41192 (N_41192,N_40753,N_40903);
nand U41193 (N_41193,N_40909,N_40986);
nand U41194 (N_41194,N_40938,N_40987);
xnor U41195 (N_41195,N_40944,N_40995);
xnor U41196 (N_41196,N_40940,N_40764);
and U41197 (N_41197,N_40927,N_40772);
or U41198 (N_41198,N_40766,N_40752);
or U41199 (N_41199,N_40916,N_40796);
and U41200 (N_41200,N_40779,N_40982);
nor U41201 (N_41201,N_40800,N_40973);
or U41202 (N_41202,N_40965,N_40964);
nor U41203 (N_41203,N_40808,N_40897);
and U41204 (N_41204,N_40960,N_40805);
nand U41205 (N_41205,N_40948,N_40890);
and U41206 (N_41206,N_40799,N_40827);
or U41207 (N_41207,N_40888,N_40866);
or U41208 (N_41208,N_40790,N_40874);
nand U41209 (N_41209,N_40784,N_40826);
nor U41210 (N_41210,N_40948,N_40843);
or U41211 (N_41211,N_40985,N_40922);
and U41212 (N_41212,N_40976,N_40858);
or U41213 (N_41213,N_40756,N_40786);
xnor U41214 (N_41214,N_40875,N_40969);
xor U41215 (N_41215,N_40870,N_40928);
xnor U41216 (N_41216,N_40784,N_40865);
xor U41217 (N_41217,N_40769,N_40800);
or U41218 (N_41218,N_40798,N_40808);
xnor U41219 (N_41219,N_40891,N_40758);
or U41220 (N_41220,N_40998,N_40951);
xor U41221 (N_41221,N_40815,N_40754);
xor U41222 (N_41222,N_40976,N_40896);
nand U41223 (N_41223,N_40772,N_40936);
nand U41224 (N_41224,N_40806,N_40936);
and U41225 (N_41225,N_40790,N_40998);
xnor U41226 (N_41226,N_40993,N_40941);
nor U41227 (N_41227,N_40966,N_40972);
nand U41228 (N_41228,N_40999,N_40785);
and U41229 (N_41229,N_40953,N_40968);
or U41230 (N_41230,N_40882,N_40949);
and U41231 (N_41231,N_40792,N_40997);
and U41232 (N_41232,N_40817,N_40830);
xnor U41233 (N_41233,N_40795,N_40914);
nor U41234 (N_41234,N_40959,N_40879);
nand U41235 (N_41235,N_40849,N_40758);
nor U41236 (N_41236,N_40795,N_40875);
and U41237 (N_41237,N_40977,N_40937);
or U41238 (N_41238,N_40918,N_40953);
and U41239 (N_41239,N_40881,N_40797);
xnor U41240 (N_41240,N_40769,N_40801);
xnor U41241 (N_41241,N_40848,N_40832);
and U41242 (N_41242,N_40787,N_40927);
nand U41243 (N_41243,N_40934,N_40857);
xor U41244 (N_41244,N_40820,N_40958);
nand U41245 (N_41245,N_40930,N_40842);
and U41246 (N_41246,N_40766,N_40926);
nand U41247 (N_41247,N_40833,N_40878);
and U41248 (N_41248,N_40790,N_40812);
and U41249 (N_41249,N_40876,N_40934);
nor U41250 (N_41250,N_41069,N_41101);
and U41251 (N_41251,N_41054,N_41236);
or U41252 (N_41252,N_41064,N_41086);
and U41253 (N_41253,N_41026,N_41149);
and U41254 (N_41254,N_41225,N_41235);
nand U41255 (N_41255,N_41098,N_41056);
nand U41256 (N_41256,N_41172,N_41090);
nor U41257 (N_41257,N_41070,N_41078);
and U41258 (N_41258,N_41115,N_41221);
xor U41259 (N_41259,N_41004,N_41219);
and U41260 (N_41260,N_41139,N_41216);
and U41261 (N_41261,N_41034,N_41093);
xor U41262 (N_41262,N_41043,N_41220);
and U41263 (N_41263,N_41127,N_41059);
nor U41264 (N_41264,N_41077,N_41052);
and U41265 (N_41265,N_41017,N_41045);
or U41266 (N_41266,N_41143,N_41103);
or U41267 (N_41267,N_41016,N_41163);
or U41268 (N_41268,N_41232,N_41071);
xnor U41269 (N_41269,N_41111,N_41075);
and U41270 (N_41270,N_41186,N_41227);
and U41271 (N_41271,N_41030,N_41014);
xnor U41272 (N_41272,N_41193,N_41205);
and U41273 (N_41273,N_41131,N_41245);
nor U41274 (N_41274,N_41124,N_41224);
and U41275 (N_41275,N_41191,N_41140);
xnor U41276 (N_41276,N_41249,N_41035);
nand U41277 (N_41277,N_41173,N_41006);
or U41278 (N_41278,N_41242,N_41113);
nor U41279 (N_41279,N_41047,N_41095);
nor U41280 (N_41280,N_41157,N_41123);
nor U41281 (N_41281,N_41137,N_41226);
xnor U41282 (N_41282,N_41151,N_41000);
and U41283 (N_41283,N_41114,N_41066);
and U41284 (N_41284,N_41058,N_41023);
or U41285 (N_41285,N_41020,N_41207);
xnor U41286 (N_41286,N_41110,N_41190);
nor U41287 (N_41287,N_41087,N_41015);
xnor U41288 (N_41288,N_41196,N_41187);
or U41289 (N_41289,N_41042,N_41146);
or U41290 (N_41290,N_41018,N_41108);
nor U41291 (N_41291,N_41073,N_41182);
xor U41292 (N_41292,N_41008,N_41141);
xnor U41293 (N_41293,N_41119,N_41233);
nor U41294 (N_41294,N_41177,N_41032);
or U41295 (N_41295,N_41229,N_41048);
or U41296 (N_41296,N_41097,N_41144);
xor U41297 (N_41297,N_41105,N_41046);
nand U41298 (N_41298,N_41028,N_41003);
xor U41299 (N_41299,N_41228,N_41145);
nor U41300 (N_41300,N_41125,N_41230);
and U41301 (N_41301,N_41150,N_41060);
nand U41302 (N_41302,N_41171,N_41112);
nand U41303 (N_41303,N_41199,N_41092);
nand U41304 (N_41304,N_41244,N_41062);
xnor U41305 (N_41305,N_41036,N_41197);
or U41306 (N_41306,N_41162,N_41084);
or U41307 (N_41307,N_41021,N_41174);
nand U41308 (N_41308,N_41049,N_41051);
and U41309 (N_41309,N_41188,N_41179);
nand U41310 (N_41310,N_41134,N_41159);
xor U41311 (N_41311,N_41041,N_41002);
or U41312 (N_41312,N_41169,N_41027);
and U41313 (N_41313,N_41135,N_41012);
xnor U41314 (N_41314,N_41133,N_41176);
xnor U41315 (N_41315,N_41106,N_41185);
and U41316 (N_41316,N_41234,N_41198);
nand U41317 (N_41317,N_41120,N_41104);
nor U41318 (N_41318,N_41237,N_41096);
or U41319 (N_41319,N_41248,N_41136);
or U41320 (N_41320,N_41116,N_41132);
nor U41321 (N_41321,N_41240,N_41184);
and U41322 (N_41322,N_41033,N_41167);
and U41323 (N_41323,N_41223,N_41118);
or U41324 (N_41324,N_41091,N_41154);
and U41325 (N_41325,N_41168,N_41181);
nand U41326 (N_41326,N_41094,N_41222);
or U41327 (N_41327,N_41231,N_41215);
nor U41328 (N_41328,N_41038,N_41044);
xor U41329 (N_41329,N_41107,N_41192);
xnor U41330 (N_41330,N_41130,N_41153);
or U41331 (N_41331,N_41005,N_41164);
and U41332 (N_41332,N_41156,N_41210);
nand U41333 (N_41333,N_41109,N_41039);
or U41334 (N_41334,N_41009,N_41001);
or U41335 (N_41335,N_41218,N_41074);
nor U41336 (N_41336,N_41081,N_41129);
and U41337 (N_41337,N_41161,N_41195);
nand U41338 (N_41338,N_41065,N_41209);
or U41339 (N_41339,N_41063,N_41175);
or U41340 (N_41340,N_41126,N_41155);
nand U41341 (N_41341,N_41100,N_41089);
or U41342 (N_41342,N_41055,N_41147);
nor U41343 (N_41343,N_41079,N_41010);
or U41344 (N_41344,N_41099,N_41057);
and U41345 (N_41345,N_41067,N_41025);
nand U41346 (N_41346,N_41022,N_41142);
xnor U41347 (N_41347,N_41165,N_41208);
or U41348 (N_41348,N_41031,N_41178);
nand U41349 (N_41349,N_41200,N_41061);
nor U41350 (N_41350,N_41053,N_41138);
and U41351 (N_41351,N_41206,N_41019);
nor U41352 (N_41352,N_41243,N_41068);
and U41353 (N_41353,N_41050,N_41217);
xnor U41354 (N_41354,N_41239,N_41029);
nand U41355 (N_41355,N_41076,N_41024);
or U41356 (N_41356,N_41080,N_41211);
nand U41357 (N_41357,N_41088,N_41247);
nand U41358 (N_41358,N_41121,N_41083);
and U41359 (N_41359,N_41213,N_41166);
nand U41360 (N_41360,N_41160,N_41040);
and U41361 (N_41361,N_41204,N_41180);
nand U41362 (N_41362,N_41152,N_41102);
nor U41363 (N_41363,N_41011,N_41203);
and U41364 (N_41364,N_41007,N_41183);
xor U41365 (N_41365,N_41013,N_41037);
nor U41366 (N_41366,N_41212,N_41128);
nor U41367 (N_41367,N_41082,N_41122);
or U41368 (N_41368,N_41072,N_41241);
nand U41369 (N_41369,N_41117,N_41201);
xor U41370 (N_41370,N_41246,N_41170);
nor U41371 (N_41371,N_41148,N_41194);
and U41372 (N_41372,N_41214,N_41202);
nand U41373 (N_41373,N_41238,N_41189);
or U41374 (N_41374,N_41158,N_41085);
nor U41375 (N_41375,N_41124,N_41029);
or U41376 (N_41376,N_41214,N_41028);
and U41377 (N_41377,N_41184,N_41145);
xor U41378 (N_41378,N_41207,N_41236);
or U41379 (N_41379,N_41239,N_41152);
or U41380 (N_41380,N_41051,N_41112);
or U41381 (N_41381,N_41133,N_41233);
xnor U41382 (N_41382,N_41048,N_41206);
nand U41383 (N_41383,N_41183,N_41069);
or U41384 (N_41384,N_41173,N_41142);
nor U41385 (N_41385,N_41182,N_41117);
nand U41386 (N_41386,N_41200,N_41208);
xor U41387 (N_41387,N_41110,N_41154);
or U41388 (N_41388,N_41121,N_41079);
xor U41389 (N_41389,N_41062,N_41229);
nand U41390 (N_41390,N_41082,N_41016);
and U41391 (N_41391,N_41179,N_41023);
xnor U41392 (N_41392,N_41105,N_41192);
nor U41393 (N_41393,N_41002,N_41079);
xnor U41394 (N_41394,N_41069,N_41143);
xnor U41395 (N_41395,N_41075,N_41175);
and U41396 (N_41396,N_41184,N_41177);
xor U41397 (N_41397,N_41065,N_41072);
nor U41398 (N_41398,N_41231,N_41103);
nor U41399 (N_41399,N_41210,N_41057);
or U41400 (N_41400,N_41062,N_41034);
nand U41401 (N_41401,N_41145,N_41113);
nor U41402 (N_41402,N_41233,N_41228);
or U41403 (N_41403,N_41051,N_41108);
nand U41404 (N_41404,N_41053,N_41004);
xor U41405 (N_41405,N_41007,N_41043);
xor U41406 (N_41406,N_41119,N_41132);
or U41407 (N_41407,N_41100,N_41068);
nor U41408 (N_41408,N_41194,N_41179);
nand U41409 (N_41409,N_41120,N_41045);
nand U41410 (N_41410,N_41075,N_41123);
nand U41411 (N_41411,N_41142,N_41240);
xnor U41412 (N_41412,N_41142,N_41016);
and U41413 (N_41413,N_41231,N_41236);
xor U41414 (N_41414,N_41236,N_41171);
xor U41415 (N_41415,N_41090,N_41143);
or U41416 (N_41416,N_41163,N_41049);
nor U41417 (N_41417,N_41085,N_41127);
xor U41418 (N_41418,N_41188,N_41165);
or U41419 (N_41419,N_41041,N_41024);
nand U41420 (N_41420,N_41153,N_41029);
or U41421 (N_41421,N_41149,N_41170);
or U41422 (N_41422,N_41003,N_41061);
nand U41423 (N_41423,N_41147,N_41053);
xnor U41424 (N_41424,N_41010,N_41177);
or U41425 (N_41425,N_41174,N_41034);
xor U41426 (N_41426,N_41161,N_41035);
xor U41427 (N_41427,N_41172,N_41147);
nor U41428 (N_41428,N_41089,N_41122);
or U41429 (N_41429,N_41001,N_41183);
nor U41430 (N_41430,N_41080,N_41062);
nor U41431 (N_41431,N_41120,N_41210);
or U41432 (N_41432,N_41206,N_41002);
nand U41433 (N_41433,N_41180,N_41038);
nand U41434 (N_41434,N_41003,N_41224);
xnor U41435 (N_41435,N_41221,N_41070);
and U41436 (N_41436,N_41044,N_41238);
nor U41437 (N_41437,N_41181,N_41056);
nor U41438 (N_41438,N_41204,N_41151);
and U41439 (N_41439,N_41193,N_41218);
nand U41440 (N_41440,N_41131,N_41041);
nand U41441 (N_41441,N_41080,N_41035);
xnor U41442 (N_41442,N_41031,N_41208);
nand U41443 (N_41443,N_41090,N_41112);
nor U41444 (N_41444,N_41043,N_41030);
nor U41445 (N_41445,N_41132,N_41071);
and U41446 (N_41446,N_41219,N_41056);
nor U41447 (N_41447,N_41085,N_41072);
and U41448 (N_41448,N_41048,N_41158);
and U41449 (N_41449,N_41043,N_41037);
or U41450 (N_41450,N_41245,N_41180);
nand U41451 (N_41451,N_41209,N_41100);
nand U41452 (N_41452,N_41207,N_41105);
nand U41453 (N_41453,N_41071,N_41081);
or U41454 (N_41454,N_41131,N_41219);
nand U41455 (N_41455,N_41229,N_41021);
nor U41456 (N_41456,N_41013,N_41025);
xnor U41457 (N_41457,N_41197,N_41180);
and U41458 (N_41458,N_41103,N_41025);
xor U41459 (N_41459,N_41170,N_41242);
xor U41460 (N_41460,N_41185,N_41169);
or U41461 (N_41461,N_41223,N_41187);
and U41462 (N_41462,N_41015,N_41029);
nor U41463 (N_41463,N_41084,N_41049);
and U41464 (N_41464,N_41178,N_41146);
and U41465 (N_41465,N_41182,N_41173);
xnor U41466 (N_41466,N_41182,N_41151);
or U41467 (N_41467,N_41097,N_41000);
or U41468 (N_41468,N_41172,N_41058);
nand U41469 (N_41469,N_41033,N_41052);
and U41470 (N_41470,N_41205,N_41048);
nand U41471 (N_41471,N_41236,N_41005);
or U41472 (N_41472,N_41247,N_41055);
xor U41473 (N_41473,N_41244,N_41125);
and U41474 (N_41474,N_41240,N_41008);
and U41475 (N_41475,N_41220,N_41074);
or U41476 (N_41476,N_41236,N_41138);
nor U41477 (N_41477,N_41085,N_41075);
xor U41478 (N_41478,N_41073,N_41148);
or U41479 (N_41479,N_41146,N_41161);
xnor U41480 (N_41480,N_41229,N_41241);
nand U41481 (N_41481,N_41227,N_41079);
xnor U41482 (N_41482,N_41067,N_41103);
nand U41483 (N_41483,N_41008,N_41202);
xor U41484 (N_41484,N_41230,N_41100);
nand U41485 (N_41485,N_41239,N_41044);
xnor U41486 (N_41486,N_41235,N_41019);
xor U41487 (N_41487,N_41062,N_41046);
nor U41488 (N_41488,N_41220,N_41194);
nor U41489 (N_41489,N_41130,N_41192);
nor U41490 (N_41490,N_41208,N_41003);
xor U41491 (N_41491,N_41000,N_41057);
or U41492 (N_41492,N_41144,N_41006);
nor U41493 (N_41493,N_41008,N_41067);
nand U41494 (N_41494,N_41227,N_41065);
nor U41495 (N_41495,N_41107,N_41052);
and U41496 (N_41496,N_41111,N_41057);
nand U41497 (N_41497,N_41181,N_41186);
xnor U41498 (N_41498,N_41200,N_41195);
nor U41499 (N_41499,N_41189,N_41129);
or U41500 (N_41500,N_41310,N_41463);
nor U41501 (N_41501,N_41419,N_41482);
nand U41502 (N_41502,N_41481,N_41483);
nand U41503 (N_41503,N_41465,N_41315);
nand U41504 (N_41504,N_41458,N_41496);
or U41505 (N_41505,N_41308,N_41394);
xnor U41506 (N_41506,N_41401,N_41352);
nand U41507 (N_41507,N_41464,N_41274);
and U41508 (N_41508,N_41428,N_41385);
nand U41509 (N_41509,N_41413,N_41408);
xnor U41510 (N_41510,N_41280,N_41422);
or U41511 (N_41511,N_41372,N_41314);
and U41512 (N_41512,N_41326,N_41291);
nor U41513 (N_41513,N_41384,N_41305);
nor U41514 (N_41514,N_41477,N_41474);
nor U41515 (N_41515,N_41479,N_41415);
nand U41516 (N_41516,N_41388,N_41398);
nand U41517 (N_41517,N_41375,N_41432);
or U41518 (N_41518,N_41475,N_41368);
or U41519 (N_41519,N_41282,N_41383);
xor U41520 (N_41520,N_41396,N_41302);
xnor U41521 (N_41521,N_41351,N_41251);
or U41522 (N_41522,N_41370,N_41341);
xnor U41523 (N_41523,N_41473,N_41488);
or U41524 (N_41524,N_41381,N_41279);
nor U41525 (N_41525,N_41424,N_41467);
and U41526 (N_41526,N_41292,N_41268);
nor U41527 (N_41527,N_41412,N_41471);
nor U41528 (N_41528,N_41491,N_41250);
and U41529 (N_41529,N_41363,N_41276);
xor U41530 (N_41530,N_41318,N_41367);
nand U41531 (N_41531,N_41322,N_41329);
and U41532 (N_41532,N_41454,N_41346);
xnor U41533 (N_41533,N_41373,N_41300);
or U41534 (N_41534,N_41357,N_41301);
xor U41535 (N_41535,N_41369,N_41362);
or U41536 (N_41536,N_41466,N_41309);
nand U41537 (N_41537,N_41321,N_41429);
xnor U41538 (N_41538,N_41495,N_41445);
xor U41539 (N_41539,N_41418,N_41349);
nand U41540 (N_41540,N_41253,N_41452);
nor U41541 (N_41541,N_41453,N_41441);
nor U41542 (N_41542,N_41430,N_41260);
and U41543 (N_41543,N_41283,N_41399);
xnor U41544 (N_41544,N_41252,N_41431);
and U41545 (N_41545,N_41350,N_41438);
and U41546 (N_41546,N_41320,N_41258);
xnor U41547 (N_41547,N_41306,N_41400);
xnor U41548 (N_41548,N_41275,N_41284);
or U41549 (N_41549,N_41286,N_41333);
nor U41550 (N_41550,N_41358,N_41397);
nor U41551 (N_41551,N_41393,N_41450);
or U41552 (N_41552,N_41311,N_41457);
nor U41553 (N_41553,N_41371,N_41435);
nor U41554 (N_41554,N_41290,N_41489);
nand U41555 (N_41555,N_41355,N_41295);
nor U41556 (N_41556,N_41386,N_41492);
or U41557 (N_41557,N_41426,N_41469);
xnor U41558 (N_41558,N_41478,N_41271);
nor U41559 (N_41559,N_41376,N_41497);
xor U41560 (N_41560,N_41294,N_41296);
xnor U41561 (N_41561,N_41262,N_41377);
or U41562 (N_41562,N_41379,N_41344);
nor U41563 (N_41563,N_41328,N_41267);
nand U41564 (N_41564,N_41392,N_41403);
and U41565 (N_41565,N_41347,N_41406);
or U41566 (N_41566,N_41484,N_41323);
xor U41567 (N_41567,N_41345,N_41331);
nand U41568 (N_41568,N_41325,N_41493);
or U41569 (N_41569,N_41263,N_41330);
nand U41570 (N_41570,N_41427,N_41281);
nor U41571 (N_41571,N_41340,N_41324);
and U41572 (N_41572,N_41269,N_41356);
and U41573 (N_41573,N_41449,N_41382);
or U41574 (N_41574,N_41451,N_41289);
xor U41575 (N_41575,N_41462,N_41421);
or U41576 (N_41576,N_41444,N_41256);
or U41577 (N_41577,N_41440,N_41277);
xor U41578 (N_41578,N_41299,N_41338);
or U41579 (N_41579,N_41380,N_41316);
nor U41580 (N_41580,N_41442,N_41312);
and U41581 (N_41581,N_41342,N_41332);
or U41582 (N_41582,N_41288,N_41254);
and U41583 (N_41583,N_41434,N_41270);
and U41584 (N_41584,N_41339,N_41410);
nand U41585 (N_41585,N_41287,N_41468);
nor U41586 (N_41586,N_41334,N_41272);
or U41587 (N_41587,N_41361,N_41387);
nand U41588 (N_41588,N_41461,N_41335);
or U41589 (N_41589,N_41494,N_41264);
xnor U41590 (N_41590,N_41317,N_41404);
and U41591 (N_41591,N_41266,N_41259);
xor U41592 (N_41592,N_41336,N_41354);
xor U41593 (N_41593,N_41261,N_41439);
or U41594 (N_41594,N_41364,N_41498);
xnor U41595 (N_41595,N_41472,N_41447);
or U41596 (N_41596,N_41389,N_41391);
nand U41597 (N_41597,N_41298,N_41307);
xor U41598 (N_41598,N_41409,N_41353);
xnor U41599 (N_41599,N_41499,N_41297);
or U41600 (N_41600,N_41348,N_41304);
xor U41601 (N_41601,N_41486,N_41337);
nor U41602 (N_41602,N_41278,N_41480);
xnor U41603 (N_41603,N_41285,N_41374);
nand U41604 (N_41604,N_41402,N_41257);
nor U41605 (N_41605,N_41265,N_41414);
and U41606 (N_41606,N_41425,N_41319);
nand U41607 (N_41607,N_41443,N_41390);
or U41608 (N_41608,N_41417,N_41420);
nand U41609 (N_41609,N_41327,N_41366);
nand U41610 (N_41610,N_41365,N_41487);
xnor U41611 (N_41611,N_41359,N_41416);
nand U41612 (N_41612,N_41448,N_41470);
or U41613 (N_41613,N_41395,N_41456);
or U41614 (N_41614,N_41455,N_41303);
or U41615 (N_41615,N_41378,N_41446);
nand U41616 (N_41616,N_41437,N_41407);
nand U41617 (N_41617,N_41490,N_41460);
nor U41618 (N_41618,N_41459,N_41485);
or U41619 (N_41619,N_41360,N_41436);
nor U41620 (N_41620,N_41343,N_41411);
nor U41621 (N_41621,N_41313,N_41293);
nand U41622 (N_41622,N_41476,N_41255);
and U41623 (N_41623,N_41433,N_41273);
or U41624 (N_41624,N_41423,N_41405);
nand U41625 (N_41625,N_41476,N_41467);
xor U41626 (N_41626,N_41409,N_41434);
xor U41627 (N_41627,N_41402,N_41273);
or U41628 (N_41628,N_41337,N_41253);
xor U41629 (N_41629,N_41379,N_41434);
xnor U41630 (N_41630,N_41297,N_41430);
xor U41631 (N_41631,N_41469,N_41460);
or U41632 (N_41632,N_41412,N_41335);
and U41633 (N_41633,N_41387,N_41303);
xnor U41634 (N_41634,N_41464,N_41289);
xnor U41635 (N_41635,N_41291,N_41432);
nor U41636 (N_41636,N_41444,N_41474);
xnor U41637 (N_41637,N_41283,N_41409);
and U41638 (N_41638,N_41254,N_41372);
and U41639 (N_41639,N_41475,N_41388);
or U41640 (N_41640,N_41429,N_41316);
nand U41641 (N_41641,N_41402,N_41464);
nor U41642 (N_41642,N_41367,N_41299);
xor U41643 (N_41643,N_41480,N_41360);
and U41644 (N_41644,N_41435,N_41338);
and U41645 (N_41645,N_41344,N_41293);
or U41646 (N_41646,N_41491,N_41359);
nor U41647 (N_41647,N_41260,N_41490);
nand U41648 (N_41648,N_41348,N_41281);
or U41649 (N_41649,N_41261,N_41283);
nand U41650 (N_41650,N_41300,N_41442);
nand U41651 (N_41651,N_41320,N_41353);
nand U41652 (N_41652,N_41289,N_41443);
and U41653 (N_41653,N_41260,N_41458);
and U41654 (N_41654,N_41269,N_41416);
and U41655 (N_41655,N_41271,N_41267);
and U41656 (N_41656,N_41338,N_41380);
xor U41657 (N_41657,N_41451,N_41422);
xnor U41658 (N_41658,N_41339,N_41432);
nor U41659 (N_41659,N_41423,N_41307);
nand U41660 (N_41660,N_41401,N_41479);
and U41661 (N_41661,N_41328,N_41461);
nor U41662 (N_41662,N_41250,N_41275);
nor U41663 (N_41663,N_41272,N_41347);
or U41664 (N_41664,N_41288,N_41444);
and U41665 (N_41665,N_41403,N_41405);
nor U41666 (N_41666,N_41372,N_41279);
and U41667 (N_41667,N_41365,N_41364);
and U41668 (N_41668,N_41282,N_41347);
nor U41669 (N_41669,N_41300,N_41342);
and U41670 (N_41670,N_41498,N_41470);
nor U41671 (N_41671,N_41273,N_41286);
nand U41672 (N_41672,N_41317,N_41491);
nor U41673 (N_41673,N_41287,N_41251);
and U41674 (N_41674,N_41462,N_41370);
nor U41675 (N_41675,N_41414,N_41392);
nand U41676 (N_41676,N_41471,N_41375);
xnor U41677 (N_41677,N_41482,N_41372);
nand U41678 (N_41678,N_41439,N_41417);
nand U41679 (N_41679,N_41477,N_41266);
xnor U41680 (N_41680,N_41332,N_41268);
xnor U41681 (N_41681,N_41260,N_41395);
xnor U41682 (N_41682,N_41465,N_41311);
nor U41683 (N_41683,N_41467,N_41359);
nand U41684 (N_41684,N_41389,N_41416);
nor U41685 (N_41685,N_41321,N_41327);
or U41686 (N_41686,N_41351,N_41453);
and U41687 (N_41687,N_41355,N_41387);
nand U41688 (N_41688,N_41323,N_41406);
or U41689 (N_41689,N_41463,N_41427);
nand U41690 (N_41690,N_41480,N_41390);
and U41691 (N_41691,N_41432,N_41342);
and U41692 (N_41692,N_41490,N_41345);
and U41693 (N_41693,N_41305,N_41488);
xnor U41694 (N_41694,N_41400,N_41499);
and U41695 (N_41695,N_41426,N_41398);
or U41696 (N_41696,N_41388,N_41430);
nand U41697 (N_41697,N_41353,N_41307);
nor U41698 (N_41698,N_41386,N_41497);
nand U41699 (N_41699,N_41418,N_41314);
nor U41700 (N_41700,N_41288,N_41317);
xnor U41701 (N_41701,N_41273,N_41431);
xnor U41702 (N_41702,N_41464,N_41465);
nand U41703 (N_41703,N_41402,N_41433);
nor U41704 (N_41704,N_41492,N_41446);
nor U41705 (N_41705,N_41407,N_41326);
nor U41706 (N_41706,N_41458,N_41447);
xnor U41707 (N_41707,N_41278,N_41252);
nand U41708 (N_41708,N_41279,N_41311);
and U41709 (N_41709,N_41257,N_41286);
and U41710 (N_41710,N_41388,N_41330);
or U41711 (N_41711,N_41294,N_41356);
nor U41712 (N_41712,N_41397,N_41252);
nor U41713 (N_41713,N_41271,N_41259);
nor U41714 (N_41714,N_41287,N_41351);
nor U41715 (N_41715,N_41459,N_41332);
and U41716 (N_41716,N_41474,N_41487);
xor U41717 (N_41717,N_41318,N_41410);
or U41718 (N_41718,N_41364,N_41308);
xor U41719 (N_41719,N_41278,N_41327);
xor U41720 (N_41720,N_41273,N_41487);
nand U41721 (N_41721,N_41309,N_41264);
or U41722 (N_41722,N_41253,N_41374);
nor U41723 (N_41723,N_41348,N_41421);
nand U41724 (N_41724,N_41452,N_41368);
nor U41725 (N_41725,N_41471,N_41483);
or U41726 (N_41726,N_41366,N_41477);
nand U41727 (N_41727,N_41409,N_41262);
and U41728 (N_41728,N_41373,N_41327);
or U41729 (N_41729,N_41499,N_41489);
or U41730 (N_41730,N_41294,N_41476);
nor U41731 (N_41731,N_41368,N_41365);
and U41732 (N_41732,N_41357,N_41334);
xor U41733 (N_41733,N_41341,N_41304);
and U41734 (N_41734,N_41448,N_41414);
nor U41735 (N_41735,N_41371,N_41444);
xnor U41736 (N_41736,N_41397,N_41425);
xnor U41737 (N_41737,N_41320,N_41302);
or U41738 (N_41738,N_41323,N_41269);
xnor U41739 (N_41739,N_41283,N_41431);
or U41740 (N_41740,N_41488,N_41264);
nand U41741 (N_41741,N_41384,N_41269);
or U41742 (N_41742,N_41447,N_41325);
or U41743 (N_41743,N_41407,N_41290);
xnor U41744 (N_41744,N_41296,N_41458);
or U41745 (N_41745,N_41323,N_41452);
nand U41746 (N_41746,N_41359,N_41342);
or U41747 (N_41747,N_41494,N_41411);
xnor U41748 (N_41748,N_41270,N_41326);
nor U41749 (N_41749,N_41395,N_41329);
or U41750 (N_41750,N_41643,N_41700);
or U41751 (N_41751,N_41648,N_41600);
and U41752 (N_41752,N_41689,N_41738);
or U41753 (N_41753,N_41595,N_41554);
nor U41754 (N_41754,N_41535,N_41638);
nor U41755 (N_41755,N_41647,N_41641);
nor U41756 (N_41756,N_41705,N_41518);
or U41757 (N_41757,N_41618,N_41704);
xor U41758 (N_41758,N_41530,N_41695);
xnor U41759 (N_41759,N_41670,N_41517);
nand U41760 (N_41760,N_41718,N_41708);
xnor U41761 (N_41761,N_41559,N_41692);
xor U41762 (N_41762,N_41674,N_41748);
or U41763 (N_41763,N_41657,N_41693);
or U41764 (N_41764,N_41685,N_41587);
and U41765 (N_41765,N_41745,N_41697);
nand U41766 (N_41766,N_41666,N_41548);
nand U41767 (N_41767,N_41734,N_41654);
and U41768 (N_41768,N_41507,N_41709);
xnor U41769 (N_41769,N_41653,N_41529);
xnor U41770 (N_41770,N_41582,N_41525);
xor U41771 (N_41771,N_41570,N_41551);
and U41772 (N_41772,N_41545,N_41658);
or U41773 (N_41773,N_41546,N_41651);
nor U41774 (N_41774,N_41702,N_41564);
nand U41775 (N_41775,N_41568,N_41544);
and U41776 (N_41776,N_41522,N_41690);
nand U41777 (N_41777,N_41605,N_41668);
or U41778 (N_41778,N_41642,N_41632);
or U41779 (N_41779,N_41677,N_41727);
and U41780 (N_41780,N_41593,N_41678);
nand U41781 (N_41781,N_41550,N_41541);
and U41782 (N_41782,N_41608,N_41649);
and U41783 (N_41783,N_41749,N_41601);
xor U41784 (N_41784,N_41591,N_41631);
nand U41785 (N_41785,N_41565,N_41664);
or U41786 (N_41786,N_41520,N_41661);
or U41787 (N_41787,N_41725,N_41562);
or U41788 (N_41788,N_41533,N_41699);
or U41789 (N_41789,N_41662,N_41573);
or U41790 (N_41790,N_41509,N_41719);
and U41791 (N_41791,N_41731,N_41592);
and U41792 (N_41792,N_41603,N_41583);
nand U41793 (N_41793,N_41706,N_41558);
or U41794 (N_41794,N_41621,N_41504);
xor U41795 (N_41795,N_41625,N_41640);
nor U41796 (N_41796,N_41694,N_41531);
xor U41797 (N_41797,N_41577,N_41511);
or U41798 (N_41798,N_41627,N_41710);
or U41799 (N_41799,N_41566,N_41644);
xor U41800 (N_41800,N_41684,N_41519);
or U41801 (N_41801,N_41510,N_41736);
xor U41802 (N_41802,N_41629,N_41744);
xnor U41803 (N_41803,N_41691,N_41610);
nand U41804 (N_41804,N_41597,N_41740);
xor U41805 (N_41805,N_41672,N_41660);
or U41806 (N_41806,N_41619,N_41534);
or U41807 (N_41807,N_41688,N_41675);
and U41808 (N_41808,N_41584,N_41626);
nor U41809 (N_41809,N_41630,N_41729);
and U41810 (N_41810,N_41521,N_41622);
nand U41811 (N_41811,N_41588,N_41623);
nor U41812 (N_41812,N_41624,N_41613);
nand U41813 (N_41813,N_41604,N_41538);
and U41814 (N_41814,N_41542,N_41527);
nand U41815 (N_41815,N_41569,N_41502);
nor U41816 (N_41816,N_41615,N_41720);
or U41817 (N_41817,N_41506,N_41737);
xnor U41818 (N_41818,N_41724,N_41614);
nand U41819 (N_41819,N_41743,N_41717);
or U41820 (N_41820,N_41579,N_41572);
and U41821 (N_41821,N_41594,N_41571);
xnor U41822 (N_41822,N_41655,N_41707);
xnor U41823 (N_41823,N_41682,N_41528);
and U41824 (N_41824,N_41721,N_41512);
xor U41825 (N_41825,N_41501,N_41611);
nand U41826 (N_41826,N_41513,N_41500);
nand U41827 (N_41827,N_41616,N_41747);
nor U41828 (N_41828,N_41516,N_41650);
xor U41829 (N_41829,N_41563,N_41671);
nand U41830 (N_41830,N_41742,N_41578);
and U41831 (N_41831,N_41679,N_41557);
nand U41832 (N_41832,N_41540,N_41634);
nand U41833 (N_41833,N_41508,N_41609);
nand U41834 (N_41834,N_41686,N_41552);
nor U41835 (N_41835,N_41585,N_41561);
nor U41836 (N_41836,N_41680,N_41711);
and U41837 (N_41837,N_41556,N_41543);
or U41838 (N_41838,N_41732,N_41726);
or U41839 (N_41839,N_41712,N_41505);
or U41840 (N_41840,N_41620,N_41515);
and U41841 (N_41841,N_41607,N_41722);
and U41842 (N_41842,N_41628,N_41602);
or U41843 (N_41843,N_41537,N_41555);
nor U41844 (N_41844,N_41547,N_41524);
nand U41845 (N_41845,N_41636,N_41696);
nand U41846 (N_41846,N_41576,N_41652);
or U41847 (N_41847,N_41635,N_41598);
xnor U41848 (N_41848,N_41687,N_41669);
and U41849 (N_41849,N_41667,N_41575);
nor U41850 (N_41850,N_41746,N_41560);
and U41851 (N_41851,N_41665,N_41739);
nand U41852 (N_41852,N_41713,N_41733);
xor U41853 (N_41853,N_41567,N_41599);
nand U41854 (N_41854,N_41580,N_41735);
nand U41855 (N_41855,N_41741,N_41703);
or U41856 (N_41856,N_41646,N_41617);
nand U41857 (N_41857,N_41659,N_41523);
nor U41858 (N_41858,N_41728,N_41681);
nand U41859 (N_41859,N_41676,N_41596);
or U41860 (N_41860,N_41549,N_41639);
nor U41861 (N_41861,N_41698,N_41701);
and U41862 (N_41862,N_41683,N_41723);
and U41863 (N_41863,N_41574,N_41656);
or U41864 (N_41864,N_41553,N_41633);
or U41865 (N_41865,N_41581,N_41645);
and U41866 (N_41866,N_41503,N_41514);
nor U41867 (N_41867,N_41716,N_41590);
or U41868 (N_41868,N_41637,N_41673);
nor U41869 (N_41869,N_41536,N_41714);
nand U41870 (N_41870,N_41526,N_41532);
nand U41871 (N_41871,N_41539,N_41606);
nand U41872 (N_41872,N_41589,N_41586);
nand U41873 (N_41873,N_41612,N_41715);
and U41874 (N_41874,N_41663,N_41730);
or U41875 (N_41875,N_41677,N_41608);
or U41876 (N_41876,N_41551,N_41554);
xor U41877 (N_41877,N_41596,N_41615);
nor U41878 (N_41878,N_41598,N_41532);
xnor U41879 (N_41879,N_41695,N_41557);
xor U41880 (N_41880,N_41737,N_41520);
or U41881 (N_41881,N_41609,N_41688);
nand U41882 (N_41882,N_41675,N_41552);
xnor U41883 (N_41883,N_41587,N_41598);
xnor U41884 (N_41884,N_41677,N_41573);
xor U41885 (N_41885,N_41705,N_41654);
xor U41886 (N_41886,N_41614,N_41563);
and U41887 (N_41887,N_41608,N_41506);
nand U41888 (N_41888,N_41515,N_41514);
nand U41889 (N_41889,N_41683,N_41677);
nor U41890 (N_41890,N_41697,N_41728);
xnor U41891 (N_41891,N_41548,N_41647);
xnor U41892 (N_41892,N_41740,N_41578);
or U41893 (N_41893,N_41748,N_41703);
or U41894 (N_41894,N_41601,N_41689);
or U41895 (N_41895,N_41516,N_41661);
nand U41896 (N_41896,N_41557,N_41678);
and U41897 (N_41897,N_41546,N_41718);
nand U41898 (N_41898,N_41544,N_41712);
nand U41899 (N_41899,N_41573,N_41578);
or U41900 (N_41900,N_41646,N_41717);
and U41901 (N_41901,N_41588,N_41738);
nor U41902 (N_41902,N_41688,N_41717);
nand U41903 (N_41903,N_41653,N_41614);
and U41904 (N_41904,N_41521,N_41535);
nand U41905 (N_41905,N_41698,N_41680);
xor U41906 (N_41906,N_41598,N_41564);
nor U41907 (N_41907,N_41520,N_41508);
nor U41908 (N_41908,N_41702,N_41533);
and U41909 (N_41909,N_41589,N_41605);
or U41910 (N_41910,N_41724,N_41705);
nor U41911 (N_41911,N_41737,N_41707);
nor U41912 (N_41912,N_41702,N_41662);
nand U41913 (N_41913,N_41527,N_41723);
and U41914 (N_41914,N_41525,N_41560);
and U41915 (N_41915,N_41513,N_41655);
xor U41916 (N_41916,N_41637,N_41624);
nand U41917 (N_41917,N_41585,N_41677);
nor U41918 (N_41918,N_41501,N_41732);
and U41919 (N_41919,N_41729,N_41673);
or U41920 (N_41920,N_41590,N_41578);
and U41921 (N_41921,N_41747,N_41501);
and U41922 (N_41922,N_41573,N_41598);
and U41923 (N_41923,N_41742,N_41554);
and U41924 (N_41924,N_41687,N_41514);
xor U41925 (N_41925,N_41591,N_41656);
nor U41926 (N_41926,N_41509,N_41720);
xnor U41927 (N_41927,N_41676,N_41561);
nand U41928 (N_41928,N_41715,N_41584);
xor U41929 (N_41929,N_41515,N_41533);
and U41930 (N_41930,N_41617,N_41518);
xor U41931 (N_41931,N_41608,N_41597);
xnor U41932 (N_41932,N_41530,N_41625);
xnor U41933 (N_41933,N_41749,N_41591);
nand U41934 (N_41934,N_41670,N_41593);
nand U41935 (N_41935,N_41721,N_41675);
xnor U41936 (N_41936,N_41727,N_41649);
nand U41937 (N_41937,N_41514,N_41624);
and U41938 (N_41938,N_41643,N_41611);
nand U41939 (N_41939,N_41533,N_41527);
nand U41940 (N_41940,N_41639,N_41714);
or U41941 (N_41941,N_41598,N_41667);
xor U41942 (N_41942,N_41530,N_41612);
nand U41943 (N_41943,N_41653,N_41654);
xnor U41944 (N_41944,N_41644,N_41684);
nand U41945 (N_41945,N_41666,N_41628);
nand U41946 (N_41946,N_41712,N_41736);
and U41947 (N_41947,N_41690,N_41654);
nand U41948 (N_41948,N_41612,N_41503);
and U41949 (N_41949,N_41620,N_41683);
nor U41950 (N_41950,N_41640,N_41638);
nor U41951 (N_41951,N_41655,N_41521);
or U41952 (N_41952,N_41651,N_41533);
nor U41953 (N_41953,N_41651,N_41606);
nand U41954 (N_41954,N_41519,N_41708);
nand U41955 (N_41955,N_41567,N_41710);
nor U41956 (N_41956,N_41692,N_41579);
and U41957 (N_41957,N_41553,N_41701);
and U41958 (N_41958,N_41692,N_41700);
and U41959 (N_41959,N_41515,N_41695);
xor U41960 (N_41960,N_41683,N_41664);
nand U41961 (N_41961,N_41624,N_41516);
nor U41962 (N_41962,N_41716,N_41749);
nor U41963 (N_41963,N_41521,N_41684);
nor U41964 (N_41964,N_41692,N_41747);
nor U41965 (N_41965,N_41659,N_41728);
nand U41966 (N_41966,N_41530,N_41701);
or U41967 (N_41967,N_41646,N_41504);
nor U41968 (N_41968,N_41664,N_41661);
xnor U41969 (N_41969,N_41624,N_41589);
nand U41970 (N_41970,N_41677,N_41631);
or U41971 (N_41971,N_41652,N_41606);
and U41972 (N_41972,N_41507,N_41505);
nor U41973 (N_41973,N_41519,N_41556);
nor U41974 (N_41974,N_41627,N_41729);
and U41975 (N_41975,N_41590,N_41546);
or U41976 (N_41976,N_41724,N_41526);
nor U41977 (N_41977,N_41509,N_41663);
nand U41978 (N_41978,N_41732,N_41637);
or U41979 (N_41979,N_41725,N_41697);
or U41980 (N_41980,N_41688,N_41629);
nor U41981 (N_41981,N_41626,N_41710);
nand U41982 (N_41982,N_41703,N_41658);
and U41983 (N_41983,N_41530,N_41596);
nand U41984 (N_41984,N_41631,N_41707);
nand U41985 (N_41985,N_41716,N_41736);
xor U41986 (N_41986,N_41682,N_41553);
or U41987 (N_41987,N_41703,N_41660);
or U41988 (N_41988,N_41511,N_41547);
xnor U41989 (N_41989,N_41730,N_41654);
nand U41990 (N_41990,N_41658,N_41526);
and U41991 (N_41991,N_41566,N_41702);
xnor U41992 (N_41992,N_41566,N_41529);
nand U41993 (N_41993,N_41718,N_41608);
nor U41994 (N_41994,N_41664,N_41668);
nand U41995 (N_41995,N_41701,N_41625);
nor U41996 (N_41996,N_41667,N_41694);
or U41997 (N_41997,N_41662,N_41513);
nand U41998 (N_41998,N_41577,N_41539);
nor U41999 (N_41999,N_41686,N_41558);
nor U42000 (N_42000,N_41922,N_41960);
nor U42001 (N_42001,N_41984,N_41900);
and U42002 (N_42002,N_41821,N_41959);
xnor U42003 (N_42003,N_41961,N_41957);
and U42004 (N_42004,N_41983,N_41840);
or U42005 (N_42005,N_41844,N_41928);
nor U42006 (N_42006,N_41810,N_41942);
or U42007 (N_42007,N_41758,N_41848);
nand U42008 (N_42008,N_41986,N_41854);
nor U42009 (N_42009,N_41949,N_41884);
or U42010 (N_42010,N_41988,N_41858);
or U42011 (N_42011,N_41901,N_41765);
and U42012 (N_42012,N_41896,N_41750);
nor U42013 (N_42013,N_41895,N_41773);
nor U42014 (N_42014,N_41891,N_41991);
and U42015 (N_42015,N_41793,N_41938);
nand U42016 (N_42016,N_41831,N_41910);
nor U42017 (N_42017,N_41812,N_41846);
nand U42018 (N_42018,N_41973,N_41985);
and U42019 (N_42019,N_41827,N_41813);
nor U42020 (N_42020,N_41953,N_41766);
and U42021 (N_42021,N_41764,N_41935);
nor U42022 (N_42022,N_41877,N_41994);
and U42023 (N_42023,N_41950,N_41776);
nor U42024 (N_42024,N_41852,N_41930);
or U42025 (N_42025,N_41948,N_41876);
and U42026 (N_42026,N_41923,N_41753);
xnor U42027 (N_42027,N_41967,N_41759);
nand U42028 (N_42028,N_41804,N_41795);
nor U42029 (N_42029,N_41826,N_41979);
nor U42030 (N_42030,N_41894,N_41865);
and U42031 (N_42031,N_41995,N_41871);
and U42032 (N_42032,N_41860,N_41911);
or U42033 (N_42033,N_41952,N_41853);
or U42034 (N_42034,N_41816,N_41751);
and U42035 (N_42035,N_41838,N_41880);
nand U42036 (N_42036,N_41921,N_41996);
xnor U42037 (N_42037,N_41917,N_41885);
nor U42038 (N_42038,N_41752,N_41822);
or U42039 (N_42039,N_41770,N_41968);
nand U42040 (N_42040,N_41886,N_41847);
nand U42041 (N_42041,N_41760,N_41805);
and U42042 (N_42042,N_41835,N_41802);
xnor U42043 (N_42043,N_41883,N_41807);
and U42044 (N_42044,N_41974,N_41989);
nand U42045 (N_42045,N_41788,N_41966);
nor U42046 (N_42046,N_41888,N_41964);
or U42047 (N_42047,N_41898,N_41841);
nand U42048 (N_42048,N_41999,N_41825);
xor U42049 (N_42049,N_41947,N_41990);
xnor U42050 (N_42050,N_41951,N_41814);
nor U42051 (N_42051,N_41798,N_41833);
xnor U42052 (N_42052,N_41828,N_41820);
and U42053 (N_42053,N_41944,N_41780);
or U42054 (N_42054,N_41934,N_41762);
or U42055 (N_42055,N_41796,N_41954);
nand U42056 (N_42056,N_41763,N_41940);
or U42057 (N_42057,N_41851,N_41893);
xor U42058 (N_42058,N_41799,N_41927);
and U42059 (N_42059,N_41970,N_41897);
and U42060 (N_42060,N_41916,N_41800);
and U42061 (N_42061,N_41830,N_41756);
nand U42062 (N_42062,N_41987,N_41857);
or U42063 (N_42063,N_41855,N_41913);
nor U42064 (N_42064,N_41811,N_41992);
and U42065 (N_42065,N_41783,N_41842);
xor U42066 (N_42066,N_41905,N_41754);
or U42067 (N_42067,N_41834,N_41778);
xor U42068 (N_42068,N_41843,N_41904);
xor U42069 (N_42069,N_41978,N_41787);
and U42070 (N_42070,N_41774,N_41909);
nor U42071 (N_42071,N_41870,N_41920);
and U42072 (N_42072,N_41823,N_41829);
nor U42073 (N_42073,N_41878,N_41769);
or U42074 (N_42074,N_41824,N_41839);
and U42075 (N_42075,N_41908,N_41859);
xnor U42076 (N_42076,N_41963,N_41863);
and U42077 (N_42077,N_41803,N_41771);
nand U42078 (N_42078,N_41819,N_41789);
and U42079 (N_42079,N_41919,N_41757);
xor U42080 (N_42080,N_41969,N_41815);
and U42081 (N_42081,N_41941,N_41955);
and U42082 (N_42082,N_41932,N_41777);
or U42083 (N_42083,N_41775,N_41976);
nand U42084 (N_42084,N_41936,N_41903);
nor U42085 (N_42085,N_41912,N_41925);
and U42086 (N_42086,N_41933,N_41926);
nand U42087 (N_42087,N_41975,N_41761);
nor U42088 (N_42088,N_41977,N_41982);
or U42089 (N_42089,N_41806,N_41768);
or U42090 (N_42090,N_41907,N_41882);
nand U42091 (N_42091,N_41862,N_41937);
xor U42092 (N_42092,N_41931,N_41869);
and U42093 (N_42093,N_41887,N_41971);
or U42094 (N_42094,N_41914,N_41866);
xor U42095 (N_42095,N_41998,N_41875);
and U42096 (N_42096,N_41958,N_41779);
and U42097 (N_42097,N_41889,N_41790);
nand U42098 (N_42098,N_41856,N_41906);
and U42099 (N_42099,N_41962,N_41818);
nor U42100 (N_42100,N_41801,N_41956);
or U42101 (N_42101,N_41832,N_41879);
and U42102 (N_42102,N_41972,N_41980);
xnor U42103 (N_42103,N_41808,N_41872);
and U42104 (N_42104,N_41915,N_41784);
nor U42105 (N_42105,N_41792,N_41868);
xor U42106 (N_42106,N_41772,N_41767);
or U42107 (N_42107,N_41929,N_41755);
nand U42108 (N_42108,N_41791,N_41946);
nand U42109 (N_42109,N_41836,N_41849);
xor U42110 (N_42110,N_41845,N_41993);
xnor U42111 (N_42111,N_41924,N_41965);
or U42112 (N_42112,N_41997,N_41943);
xor U42113 (N_42113,N_41786,N_41945);
nand U42114 (N_42114,N_41794,N_41797);
or U42115 (N_42115,N_41785,N_41782);
nor U42116 (N_42116,N_41781,N_41902);
and U42117 (N_42117,N_41867,N_41939);
and U42118 (N_42118,N_41881,N_41873);
and U42119 (N_42119,N_41874,N_41864);
nand U42120 (N_42120,N_41890,N_41837);
nor U42121 (N_42121,N_41809,N_41817);
or U42122 (N_42122,N_41981,N_41861);
nor U42123 (N_42123,N_41899,N_41918);
nor U42124 (N_42124,N_41892,N_41850);
xor U42125 (N_42125,N_41840,N_41923);
or U42126 (N_42126,N_41785,N_41780);
or U42127 (N_42127,N_41961,N_41826);
nand U42128 (N_42128,N_41909,N_41763);
and U42129 (N_42129,N_41780,N_41995);
nor U42130 (N_42130,N_41768,N_41919);
or U42131 (N_42131,N_41946,N_41955);
nor U42132 (N_42132,N_41805,N_41975);
or U42133 (N_42133,N_41833,N_41945);
or U42134 (N_42134,N_41775,N_41830);
xnor U42135 (N_42135,N_41878,N_41922);
or U42136 (N_42136,N_41841,N_41886);
nor U42137 (N_42137,N_41931,N_41857);
nand U42138 (N_42138,N_41828,N_41850);
and U42139 (N_42139,N_41959,N_41754);
nor U42140 (N_42140,N_41927,N_41896);
or U42141 (N_42141,N_41813,N_41840);
nand U42142 (N_42142,N_41941,N_41965);
nand U42143 (N_42143,N_41946,N_41867);
and U42144 (N_42144,N_41790,N_41970);
xor U42145 (N_42145,N_41971,N_41948);
xor U42146 (N_42146,N_41960,N_41861);
and U42147 (N_42147,N_41863,N_41908);
nor U42148 (N_42148,N_41799,N_41965);
and U42149 (N_42149,N_41864,N_41974);
nand U42150 (N_42150,N_41859,N_41782);
and U42151 (N_42151,N_41847,N_41822);
nor U42152 (N_42152,N_41798,N_41784);
and U42153 (N_42153,N_41792,N_41828);
xor U42154 (N_42154,N_41890,N_41989);
nor U42155 (N_42155,N_41787,N_41921);
or U42156 (N_42156,N_41928,N_41782);
and U42157 (N_42157,N_41979,N_41805);
xor U42158 (N_42158,N_41968,N_41937);
xnor U42159 (N_42159,N_41876,N_41795);
and U42160 (N_42160,N_41919,N_41960);
nor U42161 (N_42161,N_41785,N_41949);
nor U42162 (N_42162,N_41838,N_41825);
or U42163 (N_42163,N_41866,N_41756);
nand U42164 (N_42164,N_41943,N_41841);
or U42165 (N_42165,N_41894,N_41919);
or U42166 (N_42166,N_41925,N_41883);
nor U42167 (N_42167,N_41915,N_41801);
and U42168 (N_42168,N_41753,N_41963);
nor U42169 (N_42169,N_41894,N_41792);
nand U42170 (N_42170,N_41952,N_41897);
or U42171 (N_42171,N_41850,N_41794);
nand U42172 (N_42172,N_41862,N_41986);
xnor U42173 (N_42173,N_41896,N_41910);
xor U42174 (N_42174,N_41999,N_41780);
nor U42175 (N_42175,N_41973,N_41853);
or U42176 (N_42176,N_41760,N_41902);
xnor U42177 (N_42177,N_41948,N_41861);
and U42178 (N_42178,N_41761,N_41995);
or U42179 (N_42179,N_41795,N_41987);
nor U42180 (N_42180,N_41911,N_41834);
or U42181 (N_42181,N_41770,N_41852);
xor U42182 (N_42182,N_41935,N_41787);
nor U42183 (N_42183,N_41851,N_41750);
or U42184 (N_42184,N_41895,N_41970);
or U42185 (N_42185,N_41812,N_41870);
and U42186 (N_42186,N_41779,N_41979);
nand U42187 (N_42187,N_41797,N_41863);
nand U42188 (N_42188,N_41988,N_41811);
nand U42189 (N_42189,N_41878,N_41792);
and U42190 (N_42190,N_41978,N_41811);
nand U42191 (N_42191,N_41990,N_41888);
xnor U42192 (N_42192,N_41988,N_41752);
and U42193 (N_42193,N_41752,N_41985);
nand U42194 (N_42194,N_41789,N_41970);
or U42195 (N_42195,N_41996,N_41885);
nor U42196 (N_42196,N_41977,N_41809);
or U42197 (N_42197,N_41801,N_41881);
nor U42198 (N_42198,N_41936,N_41921);
xnor U42199 (N_42199,N_41864,N_41882);
and U42200 (N_42200,N_41850,N_41827);
nand U42201 (N_42201,N_41751,N_41829);
and U42202 (N_42202,N_41949,N_41771);
nand U42203 (N_42203,N_41913,N_41774);
nand U42204 (N_42204,N_41901,N_41895);
nor U42205 (N_42205,N_41857,N_41958);
nand U42206 (N_42206,N_41760,N_41764);
xnor U42207 (N_42207,N_41752,N_41865);
nor U42208 (N_42208,N_41907,N_41883);
xor U42209 (N_42209,N_41936,N_41802);
xnor U42210 (N_42210,N_41924,N_41952);
xor U42211 (N_42211,N_41819,N_41965);
and U42212 (N_42212,N_41759,N_41941);
nand U42213 (N_42213,N_41966,N_41957);
nand U42214 (N_42214,N_41987,N_41796);
or U42215 (N_42215,N_41993,N_41899);
or U42216 (N_42216,N_41770,N_41787);
nand U42217 (N_42217,N_41981,N_41904);
nand U42218 (N_42218,N_41947,N_41842);
and U42219 (N_42219,N_41937,N_41967);
or U42220 (N_42220,N_41972,N_41950);
xnor U42221 (N_42221,N_41761,N_41754);
and U42222 (N_42222,N_41766,N_41984);
nand U42223 (N_42223,N_41870,N_41916);
and U42224 (N_42224,N_41858,N_41992);
or U42225 (N_42225,N_41928,N_41941);
nor U42226 (N_42226,N_41895,N_41790);
or U42227 (N_42227,N_41999,N_41947);
or U42228 (N_42228,N_41962,N_41751);
nor U42229 (N_42229,N_41940,N_41867);
nor U42230 (N_42230,N_41952,N_41859);
and U42231 (N_42231,N_41906,N_41874);
and U42232 (N_42232,N_41876,N_41789);
xor U42233 (N_42233,N_41841,N_41984);
nor U42234 (N_42234,N_41880,N_41766);
or U42235 (N_42235,N_41798,N_41786);
xnor U42236 (N_42236,N_41816,N_41802);
nand U42237 (N_42237,N_41868,N_41964);
and U42238 (N_42238,N_41812,N_41788);
and U42239 (N_42239,N_41830,N_41893);
or U42240 (N_42240,N_41784,N_41883);
nor U42241 (N_42241,N_41851,N_41913);
xnor U42242 (N_42242,N_41774,N_41796);
nand U42243 (N_42243,N_41812,N_41768);
nand U42244 (N_42244,N_41794,N_41867);
and U42245 (N_42245,N_41795,N_41854);
xnor U42246 (N_42246,N_41752,N_41900);
and U42247 (N_42247,N_41759,N_41840);
or U42248 (N_42248,N_41981,N_41795);
and U42249 (N_42249,N_41910,N_41805);
nor U42250 (N_42250,N_42021,N_42150);
and U42251 (N_42251,N_42030,N_42061);
nand U42252 (N_42252,N_42207,N_42128);
nor U42253 (N_42253,N_42186,N_42182);
or U42254 (N_42254,N_42176,N_42071);
nand U42255 (N_42255,N_42104,N_42116);
and U42256 (N_42256,N_42154,N_42157);
or U42257 (N_42257,N_42245,N_42189);
nand U42258 (N_42258,N_42006,N_42008);
nand U42259 (N_42259,N_42249,N_42046);
nand U42260 (N_42260,N_42023,N_42027);
and U42261 (N_42261,N_42109,N_42138);
or U42262 (N_42262,N_42166,N_42136);
nand U42263 (N_42263,N_42124,N_42226);
nand U42264 (N_42264,N_42025,N_42221);
or U42265 (N_42265,N_42078,N_42044);
nor U42266 (N_42266,N_42019,N_42196);
xor U42267 (N_42267,N_42090,N_42220);
or U42268 (N_42268,N_42243,N_42033);
or U42269 (N_42269,N_42206,N_42232);
nand U42270 (N_42270,N_42056,N_42062);
nand U42271 (N_42271,N_42001,N_42171);
nor U42272 (N_42272,N_42175,N_42098);
xnor U42273 (N_42273,N_42014,N_42054);
nor U42274 (N_42274,N_42106,N_42123);
xnor U42275 (N_42275,N_42065,N_42013);
nor U42276 (N_42276,N_42092,N_42086);
nor U42277 (N_42277,N_42051,N_42228);
nor U42278 (N_42278,N_42000,N_42110);
or U42279 (N_42279,N_42129,N_42026);
and U42280 (N_42280,N_42087,N_42066);
nor U42281 (N_42281,N_42088,N_42190);
xnor U42282 (N_42282,N_42007,N_42035);
and U42283 (N_42283,N_42241,N_42057);
xnor U42284 (N_42284,N_42134,N_42219);
nor U42285 (N_42285,N_42130,N_42053);
or U42286 (N_42286,N_42178,N_42185);
nand U42287 (N_42287,N_42084,N_42063);
or U42288 (N_42288,N_42045,N_42198);
xor U42289 (N_42289,N_42173,N_42024);
and U42290 (N_42290,N_42139,N_42179);
nor U42291 (N_42291,N_42003,N_42094);
nor U42292 (N_42292,N_42216,N_42225);
nor U42293 (N_42293,N_42127,N_42015);
or U42294 (N_42294,N_42097,N_42239);
or U42295 (N_42295,N_42140,N_42042);
nor U42296 (N_42296,N_42017,N_42167);
nor U42297 (N_42297,N_42122,N_42093);
xnor U42298 (N_42298,N_42005,N_42002);
nor U42299 (N_42299,N_42037,N_42102);
and U42300 (N_42300,N_42016,N_42010);
and U42301 (N_42301,N_42163,N_42230);
nand U42302 (N_42302,N_42187,N_42073);
nor U42303 (N_42303,N_42064,N_42208);
xor U42304 (N_42304,N_42169,N_42161);
and U42305 (N_42305,N_42031,N_42246);
xor U42306 (N_42306,N_42145,N_42012);
nor U42307 (N_42307,N_42091,N_42131);
or U42308 (N_42308,N_42162,N_42222);
xor U42309 (N_42309,N_42022,N_42055);
nor U42310 (N_42310,N_42137,N_42101);
and U42311 (N_42311,N_42107,N_42205);
xor U42312 (N_42312,N_42223,N_42237);
or U42313 (N_42313,N_42089,N_42174);
nand U42314 (N_42314,N_42172,N_42077);
or U42315 (N_42315,N_42149,N_42234);
and U42316 (N_42316,N_42200,N_42195);
xor U42317 (N_42317,N_42212,N_42100);
nor U42318 (N_42318,N_42142,N_42047);
xnor U42319 (N_42319,N_42075,N_42158);
nand U42320 (N_42320,N_42121,N_42240);
nor U42321 (N_42321,N_42184,N_42183);
and U42322 (N_42322,N_42068,N_42119);
nand U42323 (N_42323,N_42112,N_42074);
nand U42324 (N_42324,N_42160,N_42080);
and U42325 (N_42325,N_42020,N_42235);
and U42326 (N_42326,N_42199,N_42151);
xnor U42327 (N_42327,N_42096,N_42108);
nor U42328 (N_42328,N_42118,N_42141);
nor U42329 (N_42329,N_42059,N_42194);
or U42330 (N_42330,N_42060,N_42132);
xor U42331 (N_42331,N_42038,N_42192);
or U42332 (N_42332,N_42011,N_42113);
or U42333 (N_42333,N_42028,N_42236);
or U42334 (N_42334,N_42204,N_42153);
nor U42335 (N_42335,N_42156,N_42120);
nand U42336 (N_42336,N_42018,N_42165);
nand U42337 (N_42337,N_42242,N_42180);
xnor U42338 (N_42338,N_42050,N_42111);
nand U42339 (N_42339,N_42164,N_42126);
nand U42340 (N_42340,N_42233,N_42004);
nor U42341 (N_42341,N_42177,N_42032);
and U42342 (N_42342,N_42070,N_42040);
and U42343 (N_42343,N_42103,N_42224);
xor U42344 (N_42344,N_42135,N_42069);
nor U42345 (N_42345,N_42193,N_42076);
nand U42346 (N_42346,N_42152,N_42247);
xor U42347 (N_42347,N_42188,N_42036);
xor U42348 (N_42348,N_42105,N_42048);
and U42349 (N_42349,N_42041,N_42067);
xor U42350 (N_42350,N_42202,N_42034);
nand U42351 (N_42351,N_42218,N_42082);
or U42352 (N_42352,N_42168,N_42201);
and U42353 (N_42353,N_42058,N_42229);
and U42354 (N_42354,N_42049,N_42039);
or U42355 (N_42355,N_42115,N_42244);
and U42356 (N_42356,N_42052,N_42125);
and U42357 (N_42357,N_42114,N_42210);
nor U42358 (N_42358,N_42211,N_42072);
nor U42359 (N_42359,N_42209,N_42231);
nor U42360 (N_42360,N_42099,N_42181);
nor U42361 (N_42361,N_42159,N_42081);
or U42362 (N_42362,N_42248,N_42214);
nor U42363 (N_42363,N_42227,N_42217);
nand U42364 (N_42364,N_42213,N_42143);
or U42365 (N_42365,N_42170,N_42147);
nor U42366 (N_42366,N_42144,N_42029);
nand U42367 (N_42367,N_42009,N_42238);
and U42368 (N_42368,N_42079,N_42148);
or U42369 (N_42369,N_42146,N_42083);
and U42370 (N_42370,N_42155,N_42197);
and U42371 (N_42371,N_42191,N_42203);
and U42372 (N_42372,N_42133,N_42085);
and U42373 (N_42373,N_42095,N_42043);
xor U42374 (N_42374,N_42117,N_42215);
nand U42375 (N_42375,N_42147,N_42032);
or U42376 (N_42376,N_42004,N_42158);
or U42377 (N_42377,N_42101,N_42037);
nor U42378 (N_42378,N_42138,N_42153);
nor U42379 (N_42379,N_42101,N_42107);
and U42380 (N_42380,N_42027,N_42043);
and U42381 (N_42381,N_42113,N_42204);
nand U42382 (N_42382,N_42151,N_42090);
and U42383 (N_42383,N_42187,N_42026);
nor U42384 (N_42384,N_42023,N_42243);
or U42385 (N_42385,N_42107,N_42141);
nand U42386 (N_42386,N_42070,N_42033);
or U42387 (N_42387,N_42210,N_42090);
nor U42388 (N_42388,N_42046,N_42045);
or U42389 (N_42389,N_42182,N_42137);
nor U42390 (N_42390,N_42097,N_42095);
and U42391 (N_42391,N_42017,N_42037);
xnor U42392 (N_42392,N_42243,N_42142);
or U42393 (N_42393,N_42155,N_42044);
and U42394 (N_42394,N_42094,N_42098);
xor U42395 (N_42395,N_42017,N_42201);
or U42396 (N_42396,N_42140,N_42241);
xor U42397 (N_42397,N_42070,N_42220);
nand U42398 (N_42398,N_42073,N_42230);
xnor U42399 (N_42399,N_42057,N_42013);
or U42400 (N_42400,N_42222,N_42227);
nor U42401 (N_42401,N_42016,N_42101);
nand U42402 (N_42402,N_42146,N_42118);
nand U42403 (N_42403,N_42247,N_42187);
or U42404 (N_42404,N_42184,N_42188);
nand U42405 (N_42405,N_42003,N_42127);
and U42406 (N_42406,N_42029,N_42074);
nand U42407 (N_42407,N_42215,N_42229);
nand U42408 (N_42408,N_42137,N_42162);
nor U42409 (N_42409,N_42042,N_42216);
nand U42410 (N_42410,N_42138,N_42005);
nor U42411 (N_42411,N_42096,N_42151);
or U42412 (N_42412,N_42170,N_42094);
nand U42413 (N_42413,N_42035,N_42186);
nand U42414 (N_42414,N_42237,N_42203);
nor U42415 (N_42415,N_42134,N_42027);
and U42416 (N_42416,N_42218,N_42134);
or U42417 (N_42417,N_42147,N_42076);
nand U42418 (N_42418,N_42157,N_42080);
and U42419 (N_42419,N_42038,N_42243);
and U42420 (N_42420,N_42113,N_42024);
nor U42421 (N_42421,N_42084,N_42191);
and U42422 (N_42422,N_42085,N_42230);
nor U42423 (N_42423,N_42234,N_42227);
nor U42424 (N_42424,N_42232,N_42067);
nor U42425 (N_42425,N_42062,N_42154);
or U42426 (N_42426,N_42152,N_42024);
nand U42427 (N_42427,N_42074,N_42161);
nand U42428 (N_42428,N_42232,N_42001);
or U42429 (N_42429,N_42013,N_42221);
xor U42430 (N_42430,N_42093,N_42220);
nand U42431 (N_42431,N_42022,N_42182);
nor U42432 (N_42432,N_42044,N_42144);
and U42433 (N_42433,N_42202,N_42056);
or U42434 (N_42434,N_42118,N_42133);
or U42435 (N_42435,N_42093,N_42118);
nor U42436 (N_42436,N_42171,N_42084);
and U42437 (N_42437,N_42073,N_42034);
and U42438 (N_42438,N_42172,N_42167);
nand U42439 (N_42439,N_42092,N_42169);
or U42440 (N_42440,N_42176,N_42049);
nand U42441 (N_42441,N_42147,N_42249);
and U42442 (N_42442,N_42240,N_42213);
and U42443 (N_42443,N_42004,N_42212);
or U42444 (N_42444,N_42162,N_42023);
xor U42445 (N_42445,N_42175,N_42157);
and U42446 (N_42446,N_42249,N_42157);
nor U42447 (N_42447,N_42099,N_42090);
xor U42448 (N_42448,N_42101,N_42068);
xnor U42449 (N_42449,N_42158,N_42028);
nand U42450 (N_42450,N_42233,N_42104);
or U42451 (N_42451,N_42054,N_42078);
nor U42452 (N_42452,N_42136,N_42214);
nor U42453 (N_42453,N_42006,N_42094);
and U42454 (N_42454,N_42122,N_42240);
nor U42455 (N_42455,N_42099,N_42146);
xor U42456 (N_42456,N_42032,N_42208);
nor U42457 (N_42457,N_42242,N_42192);
nor U42458 (N_42458,N_42105,N_42199);
and U42459 (N_42459,N_42232,N_42175);
xor U42460 (N_42460,N_42047,N_42115);
nand U42461 (N_42461,N_42034,N_42100);
xnor U42462 (N_42462,N_42177,N_42042);
and U42463 (N_42463,N_42186,N_42092);
nand U42464 (N_42464,N_42021,N_42174);
xor U42465 (N_42465,N_42140,N_42118);
nand U42466 (N_42466,N_42144,N_42037);
nor U42467 (N_42467,N_42160,N_42241);
xor U42468 (N_42468,N_42237,N_42023);
nand U42469 (N_42469,N_42138,N_42189);
xnor U42470 (N_42470,N_42209,N_42023);
nor U42471 (N_42471,N_42166,N_42001);
xor U42472 (N_42472,N_42043,N_42052);
nor U42473 (N_42473,N_42035,N_42173);
nor U42474 (N_42474,N_42243,N_42165);
or U42475 (N_42475,N_42020,N_42114);
xnor U42476 (N_42476,N_42046,N_42162);
and U42477 (N_42477,N_42007,N_42193);
nand U42478 (N_42478,N_42104,N_42067);
and U42479 (N_42479,N_42098,N_42191);
or U42480 (N_42480,N_42154,N_42156);
and U42481 (N_42481,N_42248,N_42242);
nor U42482 (N_42482,N_42108,N_42104);
nand U42483 (N_42483,N_42091,N_42190);
xor U42484 (N_42484,N_42039,N_42073);
nand U42485 (N_42485,N_42040,N_42194);
nor U42486 (N_42486,N_42228,N_42200);
nor U42487 (N_42487,N_42150,N_42142);
xnor U42488 (N_42488,N_42172,N_42232);
nor U42489 (N_42489,N_42035,N_42195);
and U42490 (N_42490,N_42153,N_42043);
and U42491 (N_42491,N_42044,N_42100);
or U42492 (N_42492,N_42069,N_42218);
xor U42493 (N_42493,N_42227,N_42130);
and U42494 (N_42494,N_42141,N_42061);
and U42495 (N_42495,N_42114,N_42198);
or U42496 (N_42496,N_42023,N_42015);
and U42497 (N_42497,N_42018,N_42177);
xor U42498 (N_42498,N_42143,N_42078);
nand U42499 (N_42499,N_42213,N_42090);
and U42500 (N_42500,N_42406,N_42388);
nor U42501 (N_42501,N_42254,N_42417);
or U42502 (N_42502,N_42376,N_42362);
nand U42503 (N_42503,N_42328,N_42432);
nor U42504 (N_42504,N_42356,N_42401);
xor U42505 (N_42505,N_42322,N_42379);
or U42506 (N_42506,N_42424,N_42421);
or U42507 (N_42507,N_42305,N_42291);
and U42508 (N_42508,N_42350,N_42450);
or U42509 (N_42509,N_42403,N_42412);
and U42510 (N_42510,N_42426,N_42252);
nand U42511 (N_42511,N_42273,N_42290);
nand U42512 (N_42512,N_42404,N_42452);
nand U42513 (N_42513,N_42486,N_42324);
or U42514 (N_42514,N_42344,N_42387);
nand U42515 (N_42515,N_42367,N_42438);
nor U42516 (N_42516,N_42439,N_42365);
nor U42517 (N_42517,N_42495,N_42283);
nor U42518 (N_42518,N_42327,N_42487);
and U42519 (N_42519,N_42384,N_42451);
and U42520 (N_42520,N_42316,N_42378);
nor U42521 (N_42521,N_42371,N_42416);
or U42522 (N_42522,N_42334,N_42383);
and U42523 (N_42523,N_42278,N_42289);
and U42524 (N_42524,N_42440,N_42483);
or U42525 (N_42525,N_42477,N_42405);
nand U42526 (N_42526,N_42366,N_42390);
and U42527 (N_42527,N_42332,N_42335);
xor U42528 (N_42528,N_42263,N_42266);
nand U42529 (N_42529,N_42295,N_42418);
nor U42530 (N_42530,N_42315,N_42275);
or U42531 (N_42531,N_42399,N_42294);
nand U42532 (N_42532,N_42341,N_42260);
or U42533 (N_42533,N_42314,N_42349);
nand U42534 (N_42534,N_42425,N_42496);
nand U42535 (N_42535,N_42377,N_42274);
nand U42536 (N_42536,N_42287,N_42470);
and U42537 (N_42537,N_42436,N_42479);
nand U42538 (N_42538,N_42343,N_42299);
xor U42539 (N_42539,N_42462,N_42296);
xnor U42540 (N_42540,N_42265,N_42397);
and U42541 (N_42541,N_42369,N_42389);
or U42542 (N_42542,N_42372,N_42256);
nand U42543 (N_42543,N_42308,N_42381);
or U42544 (N_42544,N_42474,N_42339);
and U42545 (N_42545,N_42455,N_42374);
xor U42546 (N_42546,N_42392,N_42330);
nand U42547 (N_42547,N_42300,N_42422);
nand U42548 (N_42548,N_42472,N_42414);
nand U42549 (N_42549,N_42352,N_42429);
nor U42550 (N_42550,N_42297,N_42396);
xor U42551 (N_42551,N_42269,N_42494);
or U42552 (N_42552,N_42493,N_42358);
or U42553 (N_42553,N_42435,N_42491);
xnor U42554 (N_42554,N_42329,N_42268);
or U42555 (N_42555,N_42468,N_42354);
and U42556 (N_42556,N_42411,N_42480);
nor U42557 (N_42557,N_42489,N_42364);
and U42558 (N_42558,N_42326,N_42484);
or U42559 (N_42559,N_42442,N_42340);
nor U42560 (N_42560,N_42293,N_42463);
nand U42561 (N_42561,N_42361,N_42443);
and U42562 (N_42562,N_42351,N_42393);
nand U42563 (N_42563,N_42321,N_42261);
nand U42564 (N_42564,N_42313,N_42258);
nand U42565 (N_42565,N_42395,N_42370);
and U42566 (N_42566,N_42368,N_42469);
nor U42567 (N_42567,N_42382,N_42280);
nor U42568 (N_42568,N_42445,N_42460);
nor U42569 (N_42569,N_42423,N_42453);
xor U42570 (N_42570,N_42380,N_42267);
nor U42571 (N_42571,N_42394,N_42410);
or U42572 (N_42572,N_42427,N_42375);
or U42573 (N_42573,N_42386,N_42409);
nor U42574 (N_42574,N_42400,N_42449);
or U42575 (N_42575,N_42457,N_42288);
and U42576 (N_42576,N_42492,N_42407);
nand U42577 (N_42577,N_42402,N_42465);
and U42578 (N_42578,N_42347,N_42342);
or U42579 (N_42579,N_42359,N_42337);
and U42580 (N_42580,N_42331,N_42441);
nand U42581 (N_42581,N_42257,N_42363);
nand U42582 (N_42582,N_42498,N_42385);
nor U42583 (N_42583,N_42320,N_42433);
xor U42584 (N_42584,N_42467,N_42262);
xor U42585 (N_42585,N_42454,N_42431);
xor U42586 (N_42586,N_42357,N_42490);
nand U42587 (N_42587,N_42360,N_42353);
nand U42588 (N_42588,N_42419,N_42338);
nor U42589 (N_42589,N_42475,N_42281);
nor U42590 (N_42590,N_42304,N_42481);
nand U42591 (N_42591,N_42285,N_42310);
or U42592 (N_42592,N_42250,N_42336);
nand U42593 (N_42593,N_42319,N_42437);
nand U42594 (N_42594,N_42499,N_42270);
nand U42595 (N_42595,N_42408,N_42253);
nand U42596 (N_42596,N_42413,N_42471);
xor U42597 (N_42597,N_42473,N_42346);
and U42598 (N_42598,N_42430,N_42434);
and U42599 (N_42599,N_42264,N_42282);
nor U42600 (N_42600,N_42311,N_42272);
xor U42601 (N_42601,N_42271,N_42318);
nand U42602 (N_42602,N_42415,N_42345);
nand U42603 (N_42603,N_42292,N_42276);
or U42604 (N_42604,N_42464,N_42482);
and U42605 (N_42605,N_42391,N_42323);
or U42606 (N_42606,N_42446,N_42312);
or U42607 (N_42607,N_42373,N_42348);
xnor U42608 (N_42608,N_42398,N_42476);
nand U42609 (N_42609,N_42298,N_42456);
xnor U42610 (N_42610,N_42488,N_42309);
and U42611 (N_42611,N_42428,N_42255);
nand U42612 (N_42612,N_42303,N_42466);
or U42613 (N_42613,N_42420,N_42444);
or U42614 (N_42614,N_42333,N_42317);
xor U42615 (N_42615,N_42279,N_42286);
or U42616 (N_42616,N_42459,N_42251);
nand U42617 (N_42617,N_42478,N_42259);
nor U42618 (N_42618,N_42302,N_42301);
nor U42619 (N_42619,N_42497,N_42284);
and U42620 (N_42620,N_42277,N_42325);
nand U42621 (N_42621,N_42355,N_42485);
xor U42622 (N_42622,N_42447,N_42307);
nor U42623 (N_42623,N_42306,N_42461);
nor U42624 (N_42624,N_42458,N_42448);
xnor U42625 (N_42625,N_42441,N_42292);
nand U42626 (N_42626,N_42382,N_42370);
or U42627 (N_42627,N_42365,N_42481);
nor U42628 (N_42628,N_42277,N_42379);
xnor U42629 (N_42629,N_42319,N_42375);
and U42630 (N_42630,N_42314,N_42446);
xor U42631 (N_42631,N_42372,N_42471);
nand U42632 (N_42632,N_42464,N_42367);
nor U42633 (N_42633,N_42271,N_42262);
nor U42634 (N_42634,N_42499,N_42372);
and U42635 (N_42635,N_42413,N_42293);
or U42636 (N_42636,N_42313,N_42251);
xor U42637 (N_42637,N_42399,N_42482);
or U42638 (N_42638,N_42332,N_42426);
and U42639 (N_42639,N_42318,N_42288);
xor U42640 (N_42640,N_42376,N_42346);
nand U42641 (N_42641,N_42296,N_42459);
nand U42642 (N_42642,N_42394,N_42461);
xnor U42643 (N_42643,N_42467,N_42314);
xor U42644 (N_42644,N_42314,N_42280);
or U42645 (N_42645,N_42250,N_42304);
nor U42646 (N_42646,N_42461,N_42329);
xor U42647 (N_42647,N_42317,N_42302);
or U42648 (N_42648,N_42364,N_42442);
xor U42649 (N_42649,N_42369,N_42424);
and U42650 (N_42650,N_42407,N_42475);
xor U42651 (N_42651,N_42267,N_42460);
or U42652 (N_42652,N_42328,N_42309);
nor U42653 (N_42653,N_42346,N_42411);
xnor U42654 (N_42654,N_42443,N_42463);
nor U42655 (N_42655,N_42416,N_42358);
or U42656 (N_42656,N_42382,N_42276);
xnor U42657 (N_42657,N_42446,N_42250);
and U42658 (N_42658,N_42391,N_42395);
and U42659 (N_42659,N_42360,N_42408);
nand U42660 (N_42660,N_42299,N_42476);
xor U42661 (N_42661,N_42477,N_42460);
xor U42662 (N_42662,N_42444,N_42282);
xor U42663 (N_42663,N_42496,N_42317);
and U42664 (N_42664,N_42256,N_42334);
nand U42665 (N_42665,N_42394,N_42388);
xor U42666 (N_42666,N_42376,N_42470);
xnor U42667 (N_42667,N_42365,N_42488);
and U42668 (N_42668,N_42313,N_42284);
and U42669 (N_42669,N_42466,N_42409);
or U42670 (N_42670,N_42257,N_42386);
xnor U42671 (N_42671,N_42469,N_42358);
xor U42672 (N_42672,N_42490,N_42462);
and U42673 (N_42673,N_42270,N_42432);
or U42674 (N_42674,N_42336,N_42496);
and U42675 (N_42675,N_42497,N_42263);
and U42676 (N_42676,N_42445,N_42347);
or U42677 (N_42677,N_42491,N_42416);
xnor U42678 (N_42678,N_42391,N_42294);
and U42679 (N_42679,N_42271,N_42311);
and U42680 (N_42680,N_42336,N_42401);
or U42681 (N_42681,N_42449,N_42444);
xnor U42682 (N_42682,N_42310,N_42298);
or U42683 (N_42683,N_42343,N_42304);
nand U42684 (N_42684,N_42475,N_42289);
or U42685 (N_42685,N_42427,N_42259);
and U42686 (N_42686,N_42329,N_42365);
nor U42687 (N_42687,N_42382,N_42250);
and U42688 (N_42688,N_42472,N_42491);
nand U42689 (N_42689,N_42458,N_42479);
nand U42690 (N_42690,N_42369,N_42254);
xor U42691 (N_42691,N_42301,N_42492);
nor U42692 (N_42692,N_42388,N_42335);
or U42693 (N_42693,N_42300,N_42490);
xnor U42694 (N_42694,N_42383,N_42268);
and U42695 (N_42695,N_42359,N_42310);
nand U42696 (N_42696,N_42364,N_42413);
nand U42697 (N_42697,N_42338,N_42470);
or U42698 (N_42698,N_42362,N_42287);
nor U42699 (N_42699,N_42360,N_42430);
and U42700 (N_42700,N_42489,N_42251);
nor U42701 (N_42701,N_42434,N_42433);
and U42702 (N_42702,N_42347,N_42426);
nand U42703 (N_42703,N_42474,N_42404);
nor U42704 (N_42704,N_42253,N_42356);
or U42705 (N_42705,N_42370,N_42313);
nand U42706 (N_42706,N_42336,N_42300);
or U42707 (N_42707,N_42432,N_42483);
or U42708 (N_42708,N_42278,N_42365);
xor U42709 (N_42709,N_42395,N_42313);
and U42710 (N_42710,N_42360,N_42426);
nor U42711 (N_42711,N_42333,N_42380);
and U42712 (N_42712,N_42339,N_42388);
nor U42713 (N_42713,N_42398,N_42266);
nand U42714 (N_42714,N_42285,N_42319);
or U42715 (N_42715,N_42273,N_42383);
or U42716 (N_42716,N_42374,N_42296);
xor U42717 (N_42717,N_42294,N_42258);
nor U42718 (N_42718,N_42415,N_42485);
nor U42719 (N_42719,N_42496,N_42441);
nor U42720 (N_42720,N_42323,N_42334);
nor U42721 (N_42721,N_42272,N_42281);
or U42722 (N_42722,N_42355,N_42343);
and U42723 (N_42723,N_42290,N_42388);
nor U42724 (N_42724,N_42466,N_42465);
xor U42725 (N_42725,N_42365,N_42473);
nand U42726 (N_42726,N_42282,N_42337);
and U42727 (N_42727,N_42398,N_42474);
nor U42728 (N_42728,N_42436,N_42459);
xor U42729 (N_42729,N_42460,N_42462);
or U42730 (N_42730,N_42262,N_42483);
nor U42731 (N_42731,N_42278,N_42326);
xor U42732 (N_42732,N_42435,N_42330);
and U42733 (N_42733,N_42264,N_42397);
nand U42734 (N_42734,N_42372,N_42354);
xnor U42735 (N_42735,N_42311,N_42327);
xor U42736 (N_42736,N_42259,N_42285);
xor U42737 (N_42737,N_42430,N_42306);
nand U42738 (N_42738,N_42456,N_42395);
nor U42739 (N_42739,N_42443,N_42319);
xnor U42740 (N_42740,N_42322,N_42427);
nor U42741 (N_42741,N_42341,N_42477);
and U42742 (N_42742,N_42447,N_42382);
xor U42743 (N_42743,N_42345,N_42337);
nand U42744 (N_42744,N_42410,N_42433);
nand U42745 (N_42745,N_42407,N_42338);
nand U42746 (N_42746,N_42415,N_42270);
nor U42747 (N_42747,N_42421,N_42353);
and U42748 (N_42748,N_42348,N_42428);
and U42749 (N_42749,N_42356,N_42448);
nand U42750 (N_42750,N_42663,N_42515);
and U42751 (N_42751,N_42573,N_42659);
and U42752 (N_42752,N_42534,N_42550);
xor U42753 (N_42753,N_42586,N_42649);
nor U42754 (N_42754,N_42640,N_42653);
nor U42755 (N_42755,N_42570,N_42611);
xor U42756 (N_42756,N_42609,N_42603);
nor U42757 (N_42757,N_42569,N_42744);
nand U42758 (N_42758,N_42678,N_42544);
or U42759 (N_42759,N_42541,N_42566);
nand U42760 (N_42760,N_42644,N_42561);
xnor U42761 (N_42761,N_42574,N_42720);
nand U42762 (N_42762,N_42519,N_42583);
xor U42763 (N_42763,N_42664,N_42710);
nand U42764 (N_42764,N_42636,N_42707);
nor U42765 (N_42765,N_42668,N_42715);
and U42766 (N_42766,N_42672,N_42627);
nand U42767 (N_42767,N_42656,N_42542);
and U42768 (N_42768,N_42528,N_42702);
or U42769 (N_42769,N_42575,N_42645);
nor U42770 (N_42770,N_42568,N_42598);
and U42771 (N_42771,N_42556,N_42719);
or U42772 (N_42772,N_42706,N_42741);
nor U42773 (N_42773,N_42726,N_42631);
or U42774 (N_42774,N_42617,N_42745);
nand U42775 (N_42775,N_42648,N_42504);
nor U42776 (N_42776,N_42547,N_42584);
xor U42777 (N_42777,N_42728,N_42554);
nand U42778 (N_42778,N_42622,N_42508);
and U42779 (N_42779,N_42589,N_42642);
and U42780 (N_42780,N_42703,N_42552);
and U42781 (N_42781,N_42701,N_42697);
xor U42782 (N_42782,N_42717,N_42602);
and U42783 (N_42783,N_42695,N_42647);
and U42784 (N_42784,N_42654,N_42746);
xor U42785 (N_42785,N_42633,N_42551);
nor U42786 (N_42786,N_42709,N_42527);
nor U42787 (N_42787,N_42608,N_42662);
or U42788 (N_42788,N_42543,N_42621);
xnor U42789 (N_42789,N_42600,N_42607);
nor U42790 (N_42790,N_42503,N_42591);
nor U42791 (N_42791,N_42588,N_42723);
xnor U42792 (N_42792,N_42630,N_42595);
nand U42793 (N_42793,N_42628,N_42674);
or U42794 (N_42794,N_42730,N_42536);
xnor U42795 (N_42795,N_42538,N_42634);
xor U42796 (N_42796,N_42576,N_42637);
and U42797 (N_42797,N_42587,N_42712);
xnor U42798 (N_42798,N_42567,N_42673);
nor U42799 (N_42799,N_42572,N_42713);
or U42800 (N_42800,N_42683,N_42671);
or U42801 (N_42801,N_42629,N_42520);
or U42802 (N_42802,N_42732,N_42511);
nand U42803 (N_42803,N_42688,N_42632);
nor U42804 (N_42804,N_42526,N_42523);
and U42805 (N_42805,N_42599,N_42548);
nor U42806 (N_42806,N_42646,N_42545);
xnor U42807 (N_42807,N_42650,N_42563);
nor U42808 (N_42808,N_42616,N_42643);
or U42809 (N_42809,N_42742,N_42537);
and U42810 (N_42810,N_42665,N_42601);
nor U42811 (N_42811,N_42693,N_42509);
and U42812 (N_42812,N_42675,N_42593);
or U42813 (N_42813,N_42546,N_42577);
nor U42814 (N_42814,N_42718,N_42510);
or U42815 (N_42815,N_42539,N_42558);
nand U42816 (N_42816,N_42549,N_42516);
and U42817 (N_42817,N_42560,N_42735);
nand U42818 (N_42818,N_42506,N_42734);
xor U42819 (N_42819,N_42618,N_42553);
nor U42820 (N_42820,N_42500,N_42530);
and U42821 (N_42821,N_42651,N_42738);
or U42822 (N_42822,N_42747,N_42605);
nor U42823 (N_42823,N_42559,N_42721);
xor U42824 (N_42824,N_42667,N_42580);
or U42825 (N_42825,N_42729,N_42540);
nand U42826 (N_42826,N_42613,N_42639);
and U42827 (N_42827,N_42660,N_42532);
or U42828 (N_42828,N_42597,N_42562);
nand U42829 (N_42829,N_42623,N_42733);
or U42830 (N_42830,N_42739,N_42705);
and U42831 (N_42831,N_42661,N_42596);
and U42832 (N_42832,N_42529,N_42652);
xnor U42833 (N_42833,N_42690,N_42679);
nor U42834 (N_42834,N_42525,N_42522);
nor U42835 (N_42835,N_42518,N_42686);
or U42836 (N_42836,N_42581,N_42676);
or U42837 (N_42837,N_42700,N_42711);
or U42838 (N_42838,N_42521,N_42578);
nand U42839 (N_42839,N_42749,N_42689);
xor U42840 (N_42840,N_42743,N_42725);
nor U42841 (N_42841,N_42505,N_42612);
xnor U42842 (N_42842,N_42513,N_42517);
nor U42843 (N_42843,N_42655,N_42716);
or U42844 (N_42844,N_42502,N_42692);
xnor U42845 (N_42845,N_42696,N_42687);
and U42846 (N_42846,N_42564,N_42714);
xnor U42847 (N_42847,N_42582,N_42606);
or U42848 (N_42848,N_42698,N_42699);
xor U42849 (N_42849,N_42594,N_42694);
nor U42850 (N_42850,N_42691,N_42748);
xor U42851 (N_42851,N_42579,N_42535);
and U42852 (N_42852,N_42670,N_42737);
xnor U42853 (N_42853,N_42708,N_42681);
nand U42854 (N_42854,N_42727,N_42531);
or U42855 (N_42855,N_42657,N_42624);
nor U42856 (N_42856,N_42658,N_42724);
nand U42857 (N_42857,N_42590,N_42736);
or U42858 (N_42858,N_42571,N_42680);
nor U42859 (N_42859,N_42610,N_42684);
and U42860 (N_42860,N_42533,N_42565);
or U42861 (N_42861,N_42625,N_42669);
xnor U42862 (N_42862,N_42615,N_42682);
nand U42863 (N_42863,N_42512,N_42514);
nor U42864 (N_42864,N_42666,N_42619);
or U42865 (N_42865,N_42626,N_42501);
or U42866 (N_42866,N_42524,N_42638);
or U42867 (N_42867,N_42592,N_42555);
nor U42868 (N_42868,N_42604,N_42635);
xnor U42869 (N_42869,N_42585,N_42614);
or U42870 (N_42870,N_42740,N_42620);
nand U42871 (N_42871,N_42722,N_42507);
nand U42872 (N_42872,N_42557,N_42677);
nand U42873 (N_42873,N_42731,N_42704);
nand U42874 (N_42874,N_42641,N_42685);
or U42875 (N_42875,N_42679,N_42743);
nor U42876 (N_42876,N_42661,N_42700);
or U42877 (N_42877,N_42740,N_42508);
xor U42878 (N_42878,N_42590,N_42580);
or U42879 (N_42879,N_42662,N_42584);
nor U42880 (N_42880,N_42547,N_42713);
nor U42881 (N_42881,N_42705,N_42623);
nand U42882 (N_42882,N_42635,N_42585);
and U42883 (N_42883,N_42718,N_42542);
and U42884 (N_42884,N_42720,N_42700);
xnor U42885 (N_42885,N_42555,N_42710);
xor U42886 (N_42886,N_42596,N_42589);
or U42887 (N_42887,N_42688,N_42664);
and U42888 (N_42888,N_42653,N_42710);
nor U42889 (N_42889,N_42682,N_42596);
nand U42890 (N_42890,N_42697,N_42648);
nand U42891 (N_42891,N_42683,N_42646);
xnor U42892 (N_42892,N_42515,N_42622);
nand U42893 (N_42893,N_42555,N_42526);
and U42894 (N_42894,N_42681,N_42583);
nor U42895 (N_42895,N_42563,N_42720);
xnor U42896 (N_42896,N_42610,N_42549);
xor U42897 (N_42897,N_42740,N_42699);
and U42898 (N_42898,N_42509,N_42530);
nand U42899 (N_42899,N_42655,N_42725);
or U42900 (N_42900,N_42650,N_42747);
or U42901 (N_42901,N_42574,N_42738);
nor U42902 (N_42902,N_42606,N_42714);
or U42903 (N_42903,N_42566,N_42684);
nand U42904 (N_42904,N_42590,N_42701);
or U42905 (N_42905,N_42746,N_42690);
nand U42906 (N_42906,N_42654,N_42743);
nor U42907 (N_42907,N_42689,N_42609);
nor U42908 (N_42908,N_42507,N_42713);
and U42909 (N_42909,N_42673,N_42506);
or U42910 (N_42910,N_42595,N_42547);
or U42911 (N_42911,N_42520,N_42639);
or U42912 (N_42912,N_42539,N_42703);
nor U42913 (N_42913,N_42600,N_42680);
nor U42914 (N_42914,N_42616,N_42737);
nand U42915 (N_42915,N_42734,N_42707);
nand U42916 (N_42916,N_42706,N_42707);
xnor U42917 (N_42917,N_42678,N_42728);
or U42918 (N_42918,N_42591,N_42530);
or U42919 (N_42919,N_42748,N_42716);
and U42920 (N_42920,N_42538,N_42505);
nand U42921 (N_42921,N_42534,N_42700);
or U42922 (N_42922,N_42734,N_42719);
xnor U42923 (N_42923,N_42632,N_42626);
nand U42924 (N_42924,N_42736,N_42739);
and U42925 (N_42925,N_42722,N_42626);
and U42926 (N_42926,N_42644,N_42543);
or U42927 (N_42927,N_42523,N_42534);
nand U42928 (N_42928,N_42612,N_42542);
nor U42929 (N_42929,N_42558,N_42694);
xnor U42930 (N_42930,N_42717,N_42582);
and U42931 (N_42931,N_42678,N_42745);
nand U42932 (N_42932,N_42683,N_42635);
nor U42933 (N_42933,N_42629,N_42559);
nor U42934 (N_42934,N_42576,N_42560);
nor U42935 (N_42935,N_42658,N_42527);
nor U42936 (N_42936,N_42631,N_42611);
and U42937 (N_42937,N_42594,N_42658);
nand U42938 (N_42938,N_42728,N_42570);
xnor U42939 (N_42939,N_42653,N_42709);
or U42940 (N_42940,N_42730,N_42671);
nor U42941 (N_42941,N_42748,N_42516);
nand U42942 (N_42942,N_42723,N_42694);
or U42943 (N_42943,N_42612,N_42650);
xnor U42944 (N_42944,N_42681,N_42690);
nand U42945 (N_42945,N_42649,N_42715);
nand U42946 (N_42946,N_42745,N_42622);
xnor U42947 (N_42947,N_42734,N_42597);
and U42948 (N_42948,N_42638,N_42520);
nand U42949 (N_42949,N_42695,N_42727);
nor U42950 (N_42950,N_42610,N_42632);
and U42951 (N_42951,N_42707,N_42644);
nand U42952 (N_42952,N_42699,N_42541);
or U42953 (N_42953,N_42616,N_42647);
nand U42954 (N_42954,N_42528,N_42740);
xnor U42955 (N_42955,N_42594,N_42512);
xor U42956 (N_42956,N_42523,N_42551);
xor U42957 (N_42957,N_42646,N_42501);
xnor U42958 (N_42958,N_42692,N_42712);
or U42959 (N_42959,N_42605,N_42571);
and U42960 (N_42960,N_42739,N_42523);
nand U42961 (N_42961,N_42714,N_42589);
or U42962 (N_42962,N_42600,N_42670);
xor U42963 (N_42963,N_42504,N_42727);
xor U42964 (N_42964,N_42607,N_42735);
or U42965 (N_42965,N_42611,N_42550);
nor U42966 (N_42966,N_42718,N_42613);
or U42967 (N_42967,N_42722,N_42745);
nand U42968 (N_42968,N_42582,N_42545);
nand U42969 (N_42969,N_42748,N_42617);
nor U42970 (N_42970,N_42725,N_42501);
or U42971 (N_42971,N_42536,N_42578);
or U42972 (N_42972,N_42519,N_42605);
nor U42973 (N_42973,N_42581,N_42737);
and U42974 (N_42974,N_42738,N_42533);
or U42975 (N_42975,N_42675,N_42703);
xor U42976 (N_42976,N_42696,N_42501);
xnor U42977 (N_42977,N_42559,N_42617);
or U42978 (N_42978,N_42555,N_42512);
or U42979 (N_42979,N_42660,N_42696);
xnor U42980 (N_42980,N_42686,N_42558);
nand U42981 (N_42981,N_42700,N_42684);
nand U42982 (N_42982,N_42703,N_42702);
xnor U42983 (N_42983,N_42526,N_42702);
and U42984 (N_42984,N_42616,N_42710);
or U42985 (N_42985,N_42652,N_42628);
or U42986 (N_42986,N_42586,N_42530);
nand U42987 (N_42987,N_42649,N_42711);
xnor U42988 (N_42988,N_42560,N_42542);
and U42989 (N_42989,N_42545,N_42623);
xor U42990 (N_42990,N_42650,N_42541);
and U42991 (N_42991,N_42687,N_42647);
nand U42992 (N_42992,N_42730,N_42594);
and U42993 (N_42993,N_42744,N_42602);
and U42994 (N_42994,N_42583,N_42588);
xnor U42995 (N_42995,N_42623,N_42633);
or U42996 (N_42996,N_42527,N_42632);
nand U42997 (N_42997,N_42591,N_42576);
xnor U42998 (N_42998,N_42687,N_42568);
and U42999 (N_42999,N_42550,N_42712);
and U43000 (N_43000,N_42886,N_42924);
xnor U43001 (N_43001,N_42843,N_42885);
xnor U43002 (N_43002,N_42805,N_42896);
nor U43003 (N_43003,N_42840,N_42905);
nor U43004 (N_43004,N_42862,N_42775);
and U43005 (N_43005,N_42999,N_42920);
xor U43006 (N_43006,N_42816,N_42892);
and U43007 (N_43007,N_42903,N_42763);
and U43008 (N_43008,N_42877,N_42904);
or U43009 (N_43009,N_42778,N_42867);
nor U43010 (N_43010,N_42811,N_42956);
and U43011 (N_43011,N_42829,N_42753);
and U43012 (N_43012,N_42972,N_42837);
xor U43013 (N_43013,N_42767,N_42947);
and U43014 (N_43014,N_42758,N_42939);
and U43015 (N_43015,N_42860,N_42828);
xnor U43016 (N_43016,N_42825,N_42801);
nor U43017 (N_43017,N_42998,N_42965);
nand U43018 (N_43018,N_42781,N_42821);
xor U43019 (N_43019,N_42823,N_42990);
or U43020 (N_43020,N_42911,N_42808);
xor U43021 (N_43021,N_42938,N_42832);
nand U43022 (N_43022,N_42919,N_42916);
or U43023 (N_43023,N_42987,N_42968);
xor U43024 (N_43024,N_42909,N_42879);
xnor U43025 (N_43025,N_42834,N_42777);
nand U43026 (N_43026,N_42766,N_42934);
nand U43027 (N_43027,N_42769,N_42959);
and U43028 (N_43028,N_42914,N_42951);
nand U43029 (N_43029,N_42944,N_42923);
nor U43030 (N_43030,N_42983,N_42776);
xor U43031 (N_43031,N_42949,N_42865);
xnor U43032 (N_43032,N_42815,N_42803);
xor U43033 (N_43033,N_42858,N_42994);
or U43034 (N_43034,N_42806,N_42946);
or U43035 (N_43035,N_42910,N_42785);
and U43036 (N_43036,N_42849,N_42940);
xnor U43037 (N_43037,N_42935,N_42883);
nor U43038 (N_43038,N_42848,N_42982);
xnor U43039 (N_43039,N_42888,N_42985);
and U43040 (N_43040,N_42899,N_42774);
and U43041 (N_43041,N_42966,N_42793);
or U43042 (N_43042,N_42979,N_42817);
nor U43043 (N_43043,N_42812,N_42851);
nand U43044 (N_43044,N_42901,N_42798);
xor U43045 (N_43045,N_42827,N_42988);
nand U43046 (N_43046,N_42783,N_42974);
and U43047 (N_43047,N_42772,N_42876);
or U43048 (N_43048,N_42895,N_42894);
nor U43049 (N_43049,N_42820,N_42809);
or U43050 (N_43050,N_42818,N_42853);
or U43051 (N_43051,N_42804,N_42857);
xnor U43052 (N_43052,N_42967,N_42932);
and U43053 (N_43053,N_42937,N_42992);
nand U43054 (N_43054,N_42917,N_42796);
nand U43055 (N_43055,N_42977,N_42866);
xor U43056 (N_43056,N_42969,N_42770);
nand U43057 (N_43057,N_42915,N_42791);
nor U43058 (N_43058,N_42764,N_42841);
and U43059 (N_43059,N_42995,N_42978);
nand U43060 (N_43060,N_42838,N_42850);
nand U43061 (N_43061,N_42782,N_42800);
nor U43062 (N_43062,N_42964,N_42819);
and U43063 (N_43063,N_42861,N_42868);
and U43064 (N_43064,N_42976,N_42873);
nor U43065 (N_43065,N_42790,N_42771);
and U43066 (N_43066,N_42844,N_42779);
xor U43067 (N_43067,N_42891,N_42822);
xnor U43068 (N_43068,N_42890,N_42797);
and U43069 (N_43069,N_42952,N_42773);
or U43070 (N_43070,N_42845,N_42854);
or U43071 (N_43071,N_42997,N_42786);
or U43072 (N_43072,N_42871,N_42863);
xor U43073 (N_43073,N_42780,N_42870);
nand U43074 (N_43074,N_42925,N_42882);
and U43075 (N_43075,N_42856,N_42839);
nor U43076 (N_43076,N_42931,N_42913);
and U43077 (N_43077,N_42807,N_42926);
nand U43078 (N_43078,N_42788,N_42954);
nor U43079 (N_43079,N_42933,N_42963);
and U43080 (N_43080,N_42927,N_42922);
nor U43081 (N_43081,N_42765,N_42880);
and U43082 (N_43082,N_42761,N_42887);
nand U43083 (N_43083,N_42955,N_42826);
and U43084 (N_43084,N_42852,N_42756);
nor U43085 (N_43085,N_42874,N_42941);
nor U43086 (N_43086,N_42893,N_42921);
or U43087 (N_43087,N_42872,N_42833);
nor U43088 (N_43088,N_42961,N_42962);
nor U43089 (N_43089,N_42864,N_42799);
xor U43090 (N_43090,N_42902,N_42875);
nor U43091 (N_43091,N_42918,N_42810);
or U43092 (N_43092,N_42950,N_42842);
nor U43093 (N_43093,N_42980,N_42760);
nand U43094 (N_43094,N_42953,N_42898);
xnor U43095 (N_43095,N_42906,N_42831);
and U43096 (N_43096,N_42907,N_42762);
and U43097 (N_43097,N_42957,N_42846);
and U43098 (N_43098,N_42869,N_42794);
nand U43099 (N_43099,N_42757,N_42802);
and U43100 (N_43100,N_42975,N_42936);
xor U43101 (N_43101,N_42908,N_42795);
xnor U43102 (N_43102,N_42847,N_42792);
and U43103 (N_43103,N_42750,N_42897);
nand U43104 (N_43104,N_42930,N_42993);
xor U43105 (N_43105,N_42768,N_42996);
or U43106 (N_43106,N_42973,N_42836);
and U43107 (N_43107,N_42958,N_42787);
nand U43108 (N_43108,N_42989,N_42881);
or U43109 (N_43109,N_42928,N_42889);
or U43110 (N_43110,N_42859,N_42878);
nor U43111 (N_43111,N_42981,N_42754);
nand U43112 (N_43112,N_42912,N_42900);
xnor U43113 (N_43113,N_42824,N_42784);
nand U43114 (N_43114,N_42986,N_42814);
xor U43115 (N_43115,N_42835,N_42789);
nand U43116 (N_43116,N_42948,N_42943);
nor U43117 (N_43117,N_42971,N_42970);
nand U43118 (N_43118,N_42755,N_42929);
nand U43119 (N_43119,N_42751,N_42759);
nor U43120 (N_43120,N_42960,N_42991);
nor U43121 (N_43121,N_42942,N_42855);
or U43122 (N_43122,N_42984,N_42884);
xor U43123 (N_43123,N_42830,N_42945);
xnor U43124 (N_43124,N_42813,N_42752);
nand U43125 (N_43125,N_42778,N_42900);
and U43126 (N_43126,N_42883,N_42761);
or U43127 (N_43127,N_42914,N_42787);
or U43128 (N_43128,N_42936,N_42999);
nand U43129 (N_43129,N_42864,N_42861);
nor U43130 (N_43130,N_42885,N_42944);
nor U43131 (N_43131,N_42922,N_42924);
and U43132 (N_43132,N_42789,N_42859);
and U43133 (N_43133,N_42958,N_42968);
or U43134 (N_43134,N_42803,N_42949);
xor U43135 (N_43135,N_42996,N_42751);
and U43136 (N_43136,N_42759,N_42787);
nor U43137 (N_43137,N_42992,N_42880);
nand U43138 (N_43138,N_42834,N_42771);
and U43139 (N_43139,N_42910,N_42812);
nor U43140 (N_43140,N_42894,N_42792);
and U43141 (N_43141,N_42750,N_42822);
nor U43142 (N_43142,N_42813,N_42946);
or U43143 (N_43143,N_42835,N_42909);
xor U43144 (N_43144,N_42896,N_42969);
or U43145 (N_43145,N_42837,N_42864);
nand U43146 (N_43146,N_42918,N_42966);
and U43147 (N_43147,N_42987,N_42768);
xnor U43148 (N_43148,N_42805,N_42942);
and U43149 (N_43149,N_42972,N_42862);
or U43150 (N_43150,N_42941,N_42759);
nand U43151 (N_43151,N_42766,N_42998);
and U43152 (N_43152,N_42817,N_42791);
nor U43153 (N_43153,N_42799,N_42869);
nand U43154 (N_43154,N_42858,N_42816);
nor U43155 (N_43155,N_42813,N_42785);
xor U43156 (N_43156,N_42991,N_42911);
xor U43157 (N_43157,N_42881,N_42771);
xnor U43158 (N_43158,N_42765,N_42757);
or U43159 (N_43159,N_42825,N_42989);
and U43160 (N_43160,N_42998,N_42840);
nor U43161 (N_43161,N_42994,N_42823);
nand U43162 (N_43162,N_42970,N_42992);
or U43163 (N_43163,N_42892,N_42813);
or U43164 (N_43164,N_42860,N_42939);
nand U43165 (N_43165,N_42966,N_42901);
nand U43166 (N_43166,N_42963,N_42866);
and U43167 (N_43167,N_42988,N_42765);
xor U43168 (N_43168,N_42768,N_42992);
nor U43169 (N_43169,N_42997,N_42951);
nand U43170 (N_43170,N_42755,N_42836);
or U43171 (N_43171,N_42998,N_42812);
xnor U43172 (N_43172,N_42900,N_42938);
xnor U43173 (N_43173,N_42782,N_42854);
nor U43174 (N_43174,N_42854,N_42950);
and U43175 (N_43175,N_42992,N_42831);
nand U43176 (N_43176,N_42850,N_42813);
or U43177 (N_43177,N_42875,N_42952);
nor U43178 (N_43178,N_42965,N_42942);
nor U43179 (N_43179,N_42945,N_42961);
nand U43180 (N_43180,N_42886,N_42751);
nand U43181 (N_43181,N_42808,N_42762);
nor U43182 (N_43182,N_42824,N_42864);
or U43183 (N_43183,N_42853,N_42761);
nor U43184 (N_43184,N_42810,N_42843);
xnor U43185 (N_43185,N_42826,N_42993);
nand U43186 (N_43186,N_42803,N_42971);
nand U43187 (N_43187,N_42859,N_42819);
or U43188 (N_43188,N_42917,N_42994);
nor U43189 (N_43189,N_42805,N_42842);
nand U43190 (N_43190,N_42780,N_42922);
and U43191 (N_43191,N_42753,N_42913);
or U43192 (N_43192,N_42842,N_42922);
nand U43193 (N_43193,N_42764,N_42868);
xnor U43194 (N_43194,N_42831,N_42822);
xnor U43195 (N_43195,N_42869,N_42879);
nor U43196 (N_43196,N_42953,N_42841);
and U43197 (N_43197,N_42941,N_42796);
nand U43198 (N_43198,N_42829,N_42778);
nand U43199 (N_43199,N_42961,N_42788);
nand U43200 (N_43200,N_42883,N_42998);
nor U43201 (N_43201,N_42817,N_42859);
nor U43202 (N_43202,N_42858,N_42974);
or U43203 (N_43203,N_42894,N_42837);
nand U43204 (N_43204,N_42787,N_42951);
or U43205 (N_43205,N_42793,N_42999);
nand U43206 (N_43206,N_42817,N_42795);
or U43207 (N_43207,N_42927,N_42764);
or U43208 (N_43208,N_42807,N_42790);
xnor U43209 (N_43209,N_42774,N_42888);
nand U43210 (N_43210,N_42809,N_42934);
or U43211 (N_43211,N_42768,N_42836);
or U43212 (N_43212,N_42813,N_42753);
and U43213 (N_43213,N_42855,N_42758);
and U43214 (N_43214,N_42936,N_42985);
or U43215 (N_43215,N_42849,N_42805);
or U43216 (N_43216,N_42814,N_42884);
nor U43217 (N_43217,N_42773,N_42764);
or U43218 (N_43218,N_42882,N_42824);
xnor U43219 (N_43219,N_42888,N_42787);
nor U43220 (N_43220,N_42930,N_42992);
xnor U43221 (N_43221,N_42965,N_42772);
or U43222 (N_43222,N_42849,N_42885);
xor U43223 (N_43223,N_42785,N_42881);
and U43224 (N_43224,N_42819,N_42760);
xor U43225 (N_43225,N_42944,N_42880);
and U43226 (N_43226,N_42997,N_42803);
and U43227 (N_43227,N_42780,N_42797);
xor U43228 (N_43228,N_42874,N_42955);
xnor U43229 (N_43229,N_42939,N_42794);
nor U43230 (N_43230,N_42750,N_42962);
nor U43231 (N_43231,N_42866,N_42909);
nor U43232 (N_43232,N_42953,N_42938);
and U43233 (N_43233,N_42811,N_42759);
xor U43234 (N_43234,N_42752,N_42887);
and U43235 (N_43235,N_42920,N_42986);
xor U43236 (N_43236,N_42945,N_42814);
and U43237 (N_43237,N_42976,N_42874);
nor U43238 (N_43238,N_42974,N_42980);
xnor U43239 (N_43239,N_42903,N_42971);
or U43240 (N_43240,N_42866,N_42783);
nor U43241 (N_43241,N_42889,N_42978);
xnor U43242 (N_43242,N_42804,N_42811);
and U43243 (N_43243,N_42953,N_42879);
nor U43244 (N_43244,N_42797,N_42785);
or U43245 (N_43245,N_42944,N_42886);
and U43246 (N_43246,N_42763,N_42875);
nor U43247 (N_43247,N_42921,N_42975);
or U43248 (N_43248,N_42793,N_42816);
nor U43249 (N_43249,N_42948,N_42982);
or U43250 (N_43250,N_43222,N_43180);
nand U43251 (N_43251,N_43164,N_43132);
and U43252 (N_43252,N_43120,N_43189);
xor U43253 (N_43253,N_43213,N_43092);
nand U43254 (N_43254,N_43068,N_43020);
nor U43255 (N_43255,N_43097,N_43188);
nor U43256 (N_43256,N_43015,N_43245);
or U43257 (N_43257,N_43077,N_43002);
xnor U43258 (N_43258,N_43172,N_43244);
and U43259 (N_43259,N_43158,N_43035);
nand U43260 (N_43260,N_43218,N_43049);
and U43261 (N_43261,N_43181,N_43126);
nor U43262 (N_43262,N_43215,N_43051);
nor U43263 (N_43263,N_43050,N_43118);
nand U43264 (N_43264,N_43059,N_43010);
nor U43265 (N_43265,N_43073,N_43144);
xor U43266 (N_43266,N_43153,N_43226);
or U43267 (N_43267,N_43219,N_43155);
and U43268 (N_43268,N_43101,N_43127);
xor U43269 (N_43269,N_43028,N_43193);
and U43270 (N_43270,N_43006,N_43106);
or U43271 (N_43271,N_43100,N_43096);
or U43272 (N_43272,N_43129,N_43034);
and U43273 (N_43273,N_43242,N_43210);
nor U43274 (N_43274,N_43037,N_43030);
nand U43275 (N_43275,N_43113,N_43044);
xor U43276 (N_43276,N_43115,N_43178);
and U43277 (N_43277,N_43093,N_43225);
or U43278 (N_43278,N_43067,N_43249);
xor U43279 (N_43279,N_43124,N_43098);
and U43280 (N_43280,N_43200,N_43208);
and U43281 (N_43281,N_43065,N_43169);
and U43282 (N_43282,N_43198,N_43243);
or U43283 (N_43283,N_43196,N_43229);
nand U43284 (N_43284,N_43151,N_43133);
xor U43285 (N_43285,N_43248,N_43081);
or U43286 (N_43286,N_43103,N_43109);
nor U43287 (N_43287,N_43139,N_43056);
and U43288 (N_43288,N_43197,N_43005);
nand U43289 (N_43289,N_43023,N_43060);
or U43290 (N_43290,N_43041,N_43165);
and U43291 (N_43291,N_43122,N_43230);
nor U43292 (N_43292,N_43177,N_43183);
or U43293 (N_43293,N_43085,N_43227);
xor U43294 (N_43294,N_43013,N_43039);
and U43295 (N_43295,N_43221,N_43021);
nand U43296 (N_43296,N_43147,N_43209);
xor U43297 (N_43297,N_43094,N_43022);
or U43298 (N_43298,N_43228,N_43232);
or U43299 (N_43299,N_43205,N_43176);
xnor U43300 (N_43300,N_43102,N_43187);
or U43301 (N_43301,N_43182,N_43104);
nand U43302 (N_43302,N_43003,N_43086);
nor U43303 (N_43303,N_43114,N_43237);
xnor U43304 (N_43304,N_43138,N_43069);
nand U43305 (N_43305,N_43112,N_43224);
nand U43306 (N_43306,N_43131,N_43149);
nor U43307 (N_43307,N_43231,N_43072);
or U43308 (N_43308,N_43157,N_43123);
xor U43309 (N_43309,N_43091,N_43110);
xor U43310 (N_43310,N_43089,N_43247);
nor U43311 (N_43311,N_43004,N_43170);
and U43312 (N_43312,N_43134,N_43001);
or U43313 (N_43313,N_43084,N_43063);
nand U43314 (N_43314,N_43007,N_43162);
xor U43315 (N_43315,N_43026,N_43166);
nor U43316 (N_43316,N_43038,N_43057);
or U43317 (N_43317,N_43075,N_43199);
and U43318 (N_43318,N_43024,N_43239);
xor U43319 (N_43319,N_43079,N_43192);
nand U43320 (N_43320,N_43058,N_43223);
nand U43321 (N_43321,N_43053,N_43117);
and U43322 (N_43322,N_43195,N_43047);
nand U43323 (N_43323,N_43148,N_43240);
or U43324 (N_43324,N_43066,N_43083);
nor U43325 (N_43325,N_43236,N_43052);
or U43326 (N_43326,N_43207,N_43027);
or U43327 (N_43327,N_43216,N_43241);
xnor U43328 (N_43328,N_43043,N_43150);
xor U43329 (N_43329,N_43042,N_43186);
and U43330 (N_43330,N_43204,N_43019);
or U43331 (N_43331,N_43212,N_43202);
nor U43332 (N_43332,N_43174,N_43136);
nor U43333 (N_43333,N_43175,N_43111);
xnor U43334 (N_43334,N_43029,N_43143);
and U43335 (N_43335,N_43099,N_43008);
or U43336 (N_43336,N_43190,N_43154);
or U43337 (N_43337,N_43036,N_43088);
and U43338 (N_43338,N_43234,N_43128);
nor U43339 (N_43339,N_43090,N_43233);
nor U43340 (N_43340,N_43211,N_43017);
and U43341 (N_43341,N_43009,N_43082);
nor U43342 (N_43342,N_43137,N_43238);
or U43343 (N_43343,N_43119,N_43214);
nand U43344 (N_43344,N_43142,N_43140);
nand U43345 (N_43345,N_43171,N_43217);
nor U43346 (N_43346,N_43033,N_43016);
xor U43347 (N_43347,N_43203,N_43025);
and U43348 (N_43348,N_43116,N_43107);
xnor U43349 (N_43349,N_43235,N_43161);
nor U43350 (N_43350,N_43054,N_43080);
nand U43351 (N_43351,N_43173,N_43000);
xnor U43352 (N_43352,N_43105,N_43064);
xnor U43353 (N_43353,N_43145,N_43156);
or U43354 (N_43354,N_43220,N_43168);
or U43355 (N_43355,N_43071,N_43206);
nand U43356 (N_43356,N_43130,N_43135);
and U43357 (N_43357,N_43163,N_43055);
nor U43358 (N_43358,N_43141,N_43031);
xnor U43359 (N_43359,N_43062,N_43012);
xor U43360 (N_43360,N_43179,N_43167);
nand U43361 (N_43361,N_43087,N_43191);
and U43362 (N_43362,N_43108,N_43194);
xor U43363 (N_43363,N_43046,N_43018);
nor U43364 (N_43364,N_43014,N_43048);
nor U43365 (N_43365,N_43076,N_43061);
xor U43366 (N_43366,N_43201,N_43152);
or U43367 (N_43367,N_43125,N_43246);
nand U43368 (N_43368,N_43045,N_43146);
and U43369 (N_43369,N_43185,N_43095);
nor U43370 (N_43370,N_43160,N_43040);
nand U43371 (N_43371,N_43184,N_43159);
nor U43372 (N_43372,N_43074,N_43011);
nand U43373 (N_43373,N_43032,N_43121);
xnor U43374 (N_43374,N_43078,N_43070);
nand U43375 (N_43375,N_43081,N_43030);
nand U43376 (N_43376,N_43022,N_43062);
nand U43377 (N_43377,N_43140,N_43188);
nand U43378 (N_43378,N_43081,N_43111);
or U43379 (N_43379,N_43156,N_43158);
xnor U43380 (N_43380,N_43097,N_43152);
or U43381 (N_43381,N_43163,N_43017);
nor U43382 (N_43382,N_43150,N_43195);
or U43383 (N_43383,N_43045,N_43204);
and U43384 (N_43384,N_43076,N_43227);
and U43385 (N_43385,N_43015,N_43044);
and U43386 (N_43386,N_43012,N_43009);
or U43387 (N_43387,N_43055,N_43034);
or U43388 (N_43388,N_43236,N_43244);
and U43389 (N_43389,N_43247,N_43093);
or U43390 (N_43390,N_43029,N_43216);
and U43391 (N_43391,N_43015,N_43071);
or U43392 (N_43392,N_43088,N_43152);
xnor U43393 (N_43393,N_43003,N_43007);
nor U43394 (N_43394,N_43096,N_43195);
and U43395 (N_43395,N_43177,N_43004);
or U43396 (N_43396,N_43043,N_43239);
nor U43397 (N_43397,N_43201,N_43190);
nor U43398 (N_43398,N_43229,N_43159);
nor U43399 (N_43399,N_43059,N_43079);
nor U43400 (N_43400,N_43056,N_43042);
and U43401 (N_43401,N_43066,N_43188);
and U43402 (N_43402,N_43055,N_43017);
xnor U43403 (N_43403,N_43064,N_43187);
nor U43404 (N_43404,N_43103,N_43211);
and U43405 (N_43405,N_43225,N_43014);
nand U43406 (N_43406,N_43140,N_43045);
xnor U43407 (N_43407,N_43054,N_43149);
xor U43408 (N_43408,N_43129,N_43170);
and U43409 (N_43409,N_43141,N_43177);
or U43410 (N_43410,N_43077,N_43146);
and U43411 (N_43411,N_43134,N_43061);
nor U43412 (N_43412,N_43096,N_43002);
nand U43413 (N_43413,N_43136,N_43166);
xnor U43414 (N_43414,N_43135,N_43207);
and U43415 (N_43415,N_43034,N_43109);
or U43416 (N_43416,N_43030,N_43046);
nor U43417 (N_43417,N_43046,N_43093);
and U43418 (N_43418,N_43053,N_43044);
or U43419 (N_43419,N_43081,N_43007);
and U43420 (N_43420,N_43030,N_43178);
or U43421 (N_43421,N_43167,N_43019);
nor U43422 (N_43422,N_43072,N_43154);
and U43423 (N_43423,N_43162,N_43046);
xnor U43424 (N_43424,N_43001,N_43233);
nand U43425 (N_43425,N_43017,N_43142);
nor U43426 (N_43426,N_43030,N_43158);
nor U43427 (N_43427,N_43074,N_43221);
nand U43428 (N_43428,N_43142,N_43082);
or U43429 (N_43429,N_43156,N_43207);
or U43430 (N_43430,N_43129,N_43230);
and U43431 (N_43431,N_43226,N_43195);
nor U43432 (N_43432,N_43108,N_43206);
xnor U43433 (N_43433,N_43070,N_43032);
nand U43434 (N_43434,N_43163,N_43068);
nand U43435 (N_43435,N_43193,N_43185);
nand U43436 (N_43436,N_43234,N_43211);
nor U43437 (N_43437,N_43096,N_43011);
nor U43438 (N_43438,N_43117,N_43150);
or U43439 (N_43439,N_43088,N_43084);
and U43440 (N_43440,N_43016,N_43062);
nor U43441 (N_43441,N_43014,N_43036);
or U43442 (N_43442,N_43206,N_43186);
and U43443 (N_43443,N_43165,N_43247);
nor U43444 (N_43444,N_43012,N_43248);
or U43445 (N_43445,N_43031,N_43155);
xor U43446 (N_43446,N_43231,N_43105);
xor U43447 (N_43447,N_43061,N_43092);
and U43448 (N_43448,N_43142,N_43102);
nor U43449 (N_43449,N_43073,N_43246);
nor U43450 (N_43450,N_43216,N_43032);
nand U43451 (N_43451,N_43051,N_43045);
and U43452 (N_43452,N_43119,N_43205);
nand U43453 (N_43453,N_43199,N_43238);
or U43454 (N_43454,N_43086,N_43036);
and U43455 (N_43455,N_43110,N_43199);
nand U43456 (N_43456,N_43099,N_43223);
and U43457 (N_43457,N_43182,N_43139);
or U43458 (N_43458,N_43233,N_43234);
nand U43459 (N_43459,N_43108,N_43144);
nor U43460 (N_43460,N_43150,N_43249);
or U43461 (N_43461,N_43007,N_43054);
and U43462 (N_43462,N_43033,N_43064);
and U43463 (N_43463,N_43152,N_43102);
or U43464 (N_43464,N_43157,N_43016);
xnor U43465 (N_43465,N_43195,N_43022);
xnor U43466 (N_43466,N_43062,N_43235);
and U43467 (N_43467,N_43097,N_43128);
xor U43468 (N_43468,N_43196,N_43026);
or U43469 (N_43469,N_43154,N_43015);
xor U43470 (N_43470,N_43143,N_43078);
nand U43471 (N_43471,N_43017,N_43081);
and U43472 (N_43472,N_43237,N_43159);
xnor U43473 (N_43473,N_43159,N_43056);
and U43474 (N_43474,N_43247,N_43154);
or U43475 (N_43475,N_43236,N_43101);
nor U43476 (N_43476,N_43164,N_43229);
and U43477 (N_43477,N_43090,N_43018);
and U43478 (N_43478,N_43179,N_43116);
or U43479 (N_43479,N_43100,N_43028);
xor U43480 (N_43480,N_43169,N_43002);
nor U43481 (N_43481,N_43146,N_43175);
nand U43482 (N_43482,N_43091,N_43060);
nor U43483 (N_43483,N_43226,N_43066);
and U43484 (N_43484,N_43074,N_43089);
xor U43485 (N_43485,N_43181,N_43207);
and U43486 (N_43486,N_43110,N_43089);
nor U43487 (N_43487,N_43034,N_43176);
and U43488 (N_43488,N_43119,N_43032);
nor U43489 (N_43489,N_43064,N_43221);
nor U43490 (N_43490,N_43044,N_43091);
nand U43491 (N_43491,N_43153,N_43181);
nand U43492 (N_43492,N_43130,N_43037);
nand U43493 (N_43493,N_43178,N_43079);
or U43494 (N_43494,N_43131,N_43158);
or U43495 (N_43495,N_43127,N_43138);
and U43496 (N_43496,N_43127,N_43117);
nand U43497 (N_43497,N_43071,N_43060);
xnor U43498 (N_43498,N_43066,N_43208);
nor U43499 (N_43499,N_43234,N_43195);
nor U43500 (N_43500,N_43424,N_43313);
nand U43501 (N_43501,N_43344,N_43371);
nand U43502 (N_43502,N_43347,N_43289);
xor U43503 (N_43503,N_43298,N_43314);
or U43504 (N_43504,N_43497,N_43479);
nand U43505 (N_43505,N_43340,N_43267);
and U43506 (N_43506,N_43356,N_43331);
nand U43507 (N_43507,N_43264,N_43462);
or U43508 (N_43508,N_43461,N_43450);
xnor U43509 (N_43509,N_43297,N_43433);
nor U43510 (N_43510,N_43402,N_43287);
or U43511 (N_43511,N_43251,N_43386);
or U43512 (N_43512,N_43390,N_43373);
xor U43513 (N_43513,N_43327,N_43421);
and U43514 (N_43514,N_43438,N_43397);
xnor U43515 (N_43515,N_43477,N_43376);
nand U43516 (N_43516,N_43447,N_43367);
and U43517 (N_43517,N_43322,N_43423);
xnor U43518 (N_43518,N_43355,N_43398);
or U43519 (N_43519,N_43266,N_43427);
xnor U43520 (N_43520,N_43299,N_43359);
nor U43521 (N_43521,N_43329,N_43354);
or U43522 (N_43522,N_43481,N_43303);
xor U43523 (N_43523,N_43432,N_43494);
xnor U43524 (N_43524,N_43403,N_43417);
nor U43525 (N_43525,N_43429,N_43368);
and U43526 (N_43526,N_43414,N_43441);
nor U43527 (N_43527,N_43280,N_43288);
xor U43528 (N_43528,N_43319,N_43454);
and U43529 (N_43529,N_43286,N_43457);
nand U43530 (N_43530,N_43250,N_43338);
xor U43531 (N_43531,N_43446,N_43475);
xor U43532 (N_43532,N_43255,N_43361);
xnor U43533 (N_43533,N_43408,N_43436);
or U43534 (N_43534,N_43422,N_43320);
xnor U43535 (N_43535,N_43310,N_43404);
nand U43536 (N_43536,N_43326,N_43366);
nor U43537 (N_43537,N_43258,N_43316);
or U43538 (N_43538,N_43295,N_43315);
or U43539 (N_43539,N_43352,N_43259);
nor U43540 (N_43540,N_43453,N_43296);
nor U43541 (N_43541,N_43499,N_43269);
nand U43542 (N_43542,N_43407,N_43469);
nor U43543 (N_43543,N_43253,N_43484);
nand U43544 (N_43544,N_43437,N_43379);
xnor U43545 (N_43545,N_43349,N_43276);
nand U43546 (N_43546,N_43318,N_43274);
and U43547 (N_43547,N_43463,N_43485);
nor U43548 (N_43548,N_43419,N_43409);
and U43549 (N_43549,N_43363,N_43336);
nor U43550 (N_43550,N_43442,N_43337);
and U43551 (N_43551,N_43440,N_43439);
and U43552 (N_43552,N_43343,N_43473);
and U43553 (N_43553,N_43489,N_43305);
nand U43554 (N_43554,N_43333,N_43448);
or U43555 (N_43555,N_43396,N_43444);
xor U43556 (N_43556,N_43480,N_43478);
xnor U43557 (N_43557,N_43418,N_43411);
nor U43558 (N_43558,N_43293,N_43341);
nor U43559 (N_43559,N_43375,N_43393);
xor U43560 (N_43560,N_43456,N_43377);
nor U43561 (N_43561,N_43474,N_43487);
or U43562 (N_43562,N_43496,N_43372);
or U43563 (N_43563,N_43370,N_43323);
and U43564 (N_43564,N_43385,N_43278);
nand U43565 (N_43565,N_43490,N_43256);
or U43566 (N_43566,N_43459,N_43304);
nand U43567 (N_43567,N_43300,N_43260);
nor U43568 (N_43568,N_43428,N_43348);
and U43569 (N_43569,N_43262,N_43351);
nand U43570 (N_43570,N_43282,N_43283);
and U43571 (N_43571,N_43415,N_43334);
and U43572 (N_43572,N_43395,N_43291);
xnor U43573 (N_43573,N_43321,N_43335);
nor U43574 (N_43574,N_43412,N_43272);
and U43575 (N_43575,N_43380,N_43382);
and U43576 (N_43576,N_43277,N_43261);
or U43577 (N_43577,N_43265,N_43330);
nor U43578 (N_43578,N_43400,N_43471);
nor U43579 (N_43579,N_43464,N_43468);
xnor U43580 (N_43580,N_43275,N_43342);
or U43581 (N_43581,N_43425,N_43362);
nand U43582 (N_43582,N_43345,N_43290);
or U43583 (N_43583,N_43460,N_43394);
xnor U43584 (N_43584,N_43328,N_43399);
nand U43585 (N_43585,N_43324,N_43353);
xnor U43586 (N_43586,N_43452,N_43284);
xor U43587 (N_43587,N_43498,N_43426);
and U43588 (N_43588,N_43431,N_43346);
nand U43589 (N_43589,N_43410,N_43451);
nor U43590 (N_43590,N_43443,N_43430);
nand U43591 (N_43591,N_43306,N_43383);
xnor U43592 (N_43592,N_43369,N_43389);
or U43593 (N_43593,N_43401,N_43413);
or U43594 (N_43594,N_43378,N_43263);
nand U43595 (N_43595,N_43332,N_43492);
xor U43596 (N_43596,N_43360,N_43466);
xnor U43597 (N_43597,N_43406,N_43252);
or U43598 (N_43598,N_43365,N_43488);
or U43599 (N_43599,N_43388,N_43495);
xor U43600 (N_43600,N_43455,N_43358);
nand U43601 (N_43601,N_43301,N_43482);
and U43602 (N_43602,N_43364,N_43387);
nand U43603 (N_43603,N_43281,N_43350);
xnor U43604 (N_43604,N_43465,N_43302);
and U43605 (N_43605,N_43405,N_43486);
nand U43606 (N_43606,N_43420,N_43493);
nor U43607 (N_43607,N_43308,N_43476);
xnor U43608 (N_43608,N_43445,N_43470);
and U43609 (N_43609,N_43458,N_43311);
xor U43610 (N_43610,N_43294,N_43491);
nand U43611 (N_43611,N_43416,N_43312);
or U43612 (N_43612,N_43307,N_43392);
nand U43613 (N_43613,N_43271,N_43391);
nor U43614 (N_43614,N_43339,N_43435);
and U43615 (N_43615,N_43309,N_43285);
and U43616 (N_43616,N_43381,N_43279);
xor U43617 (N_43617,N_43317,N_43254);
nand U43618 (N_43618,N_43325,N_43257);
xor U43619 (N_43619,N_43467,N_43357);
and U43620 (N_43620,N_43384,N_43472);
nand U43621 (N_43621,N_43374,N_43434);
nand U43622 (N_43622,N_43273,N_43268);
or U43623 (N_43623,N_43270,N_43449);
nor U43624 (N_43624,N_43483,N_43292);
and U43625 (N_43625,N_43342,N_43358);
nand U43626 (N_43626,N_43256,N_43460);
xor U43627 (N_43627,N_43401,N_43409);
nand U43628 (N_43628,N_43269,N_43436);
nor U43629 (N_43629,N_43347,N_43252);
nor U43630 (N_43630,N_43341,N_43471);
nor U43631 (N_43631,N_43391,N_43450);
and U43632 (N_43632,N_43364,N_43330);
and U43633 (N_43633,N_43418,N_43279);
nand U43634 (N_43634,N_43424,N_43380);
xnor U43635 (N_43635,N_43314,N_43342);
nor U43636 (N_43636,N_43395,N_43352);
xnor U43637 (N_43637,N_43339,N_43373);
nand U43638 (N_43638,N_43492,N_43411);
or U43639 (N_43639,N_43295,N_43457);
xor U43640 (N_43640,N_43431,N_43295);
or U43641 (N_43641,N_43329,N_43456);
xor U43642 (N_43642,N_43409,N_43317);
or U43643 (N_43643,N_43453,N_43263);
xnor U43644 (N_43644,N_43465,N_43269);
xor U43645 (N_43645,N_43258,N_43437);
and U43646 (N_43646,N_43360,N_43424);
nand U43647 (N_43647,N_43401,N_43334);
nand U43648 (N_43648,N_43368,N_43357);
or U43649 (N_43649,N_43453,N_43430);
xnor U43650 (N_43650,N_43411,N_43450);
and U43651 (N_43651,N_43488,N_43482);
xor U43652 (N_43652,N_43464,N_43429);
xnor U43653 (N_43653,N_43426,N_43285);
and U43654 (N_43654,N_43457,N_43287);
nand U43655 (N_43655,N_43399,N_43495);
nand U43656 (N_43656,N_43367,N_43354);
nand U43657 (N_43657,N_43460,N_43277);
or U43658 (N_43658,N_43334,N_43475);
nor U43659 (N_43659,N_43470,N_43262);
xor U43660 (N_43660,N_43260,N_43370);
or U43661 (N_43661,N_43286,N_43351);
or U43662 (N_43662,N_43265,N_43329);
and U43663 (N_43663,N_43358,N_43357);
nor U43664 (N_43664,N_43286,N_43495);
nor U43665 (N_43665,N_43475,N_43384);
or U43666 (N_43666,N_43288,N_43258);
and U43667 (N_43667,N_43355,N_43362);
nand U43668 (N_43668,N_43370,N_43359);
nand U43669 (N_43669,N_43447,N_43432);
nor U43670 (N_43670,N_43478,N_43367);
or U43671 (N_43671,N_43292,N_43256);
nor U43672 (N_43672,N_43490,N_43428);
nor U43673 (N_43673,N_43427,N_43482);
xnor U43674 (N_43674,N_43357,N_43430);
or U43675 (N_43675,N_43276,N_43439);
xor U43676 (N_43676,N_43485,N_43401);
and U43677 (N_43677,N_43338,N_43341);
nand U43678 (N_43678,N_43292,N_43382);
nand U43679 (N_43679,N_43282,N_43348);
xor U43680 (N_43680,N_43302,N_43488);
nor U43681 (N_43681,N_43449,N_43345);
nor U43682 (N_43682,N_43489,N_43422);
xnor U43683 (N_43683,N_43269,N_43491);
nand U43684 (N_43684,N_43302,N_43431);
xnor U43685 (N_43685,N_43353,N_43262);
nor U43686 (N_43686,N_43485,N_43311);
and U43687 (N_43687,N_43435,N_43345);
nand U43688 (N_43688,N_43348,N_43328);
xor U43689 (N_43689,N_43361,N_43346);
nor U43690 (N_43690,N_43360,N_43491);
and U43691 (N_43691,N_43463,N_43460);
and U43692 (N_43692,N_43255,N_43401);
nand U43693 (N_43693,N_43340,N_43370);
xnor U43694 (N_43694,N_43341,N_43420);
or U43695 (N_43695,N_43446,N_43477);
nor U43696 (N_43696,N_43329,N_43416);
or U43697 (N_43697,N_43483,N_43301);
or U43698 (N_43698,N_43429,N_43451);
and U43699 (N_43699,N_43321,N_43349);
xor U43700 (N_43700,N_43384,N_43441);
nand U43701 (N_43701,N_43302,N_43412);
or U43702 (N_43702,N_43298,N_43359);
or U43703 (N_43703,N_43434,N_43483);
xnor U43704 (N_43704,N_43355,N_43271);
xor U43705 (N_43705,N_43302,N_43296);
nor U43706 (N_43706,N_43319,N_43352);
xnor U43707 (N_43707,N_43428,N_43340);
or U43708 (N_43708,N_43363,N_43258);
or U43709 (N_43709,N_43350,N_43479);
and U43710 (N_43710,N_43414,N_43443);
and U43711 (N_43711,N_43392,N_43385);
and U43712 (N_43712,N_43278,N_43383);
xnor U43713 (N_43713,N_43391,N_43301);
nor U43714 (N_43714,N_43468,N_43386);
nor U43715 (N_43715,N_43293,N_43361);
xnor U43716 (N_43716,N_43373,N_43272);
nand U43717 (N_43717,N_43325,N_43309);
nand U43718 (N_43718,N_43300,N_43396);
and U43719 (N_43719,N_43415,N_43333);
or U43720 (N_43720,N_43276,N_43409);
and U43721 (N_43721,N_43359,N_43430);
and U43722 (N_43722,N_43451,N_43400);
nor U43723 (N_43723,N_43328,N_43403);
nor U43724 (N_43724,N_43299,N_43349);
nand U43725 (N_43725,N_43425,N_43405);
and U43726 (N_43726,N_43275,N_43296);
or U43727 (N_43727,N_43401,N_43412);
nand U43728 (N_43728,N_43367,N_43262);
or U43729 (N_43729,N_43486,N_43465);
nand U43730 (N_43730,N_43262,N_43364);
nor U43731 (N_43731,N_43445,N_43480);
nand U43732 (N_43732,N_43417,N_43454);
nor U43733 (N_43733,N_43420,N_43372);
and U43734 (N_43734,N_43454,N_43415);
nor U43735 (N_43735,N_43362,N_43383);
nor U43736 (N_43736,N_43342,N_43302);
xor U43737 (N_43737,N_43468,N_43423);
nor U43738 (N_43738,N_43485,N_43304);
and U43739 (N_43739,N_43495,N_43342);
nor U43740 (N_43740,N_43310,N_43339);
nor U43741 (N_43741,N_43359,N_43301);
nor U43742 (N_43742,N_43391,N_43492);
xnor U43743 (N_43743,N_43310,N_43323);
or U43744 (N_43744,N_43404,N_43304);
or U43745 (N_43745,N_43307,N_43443);
and U43746 (N_43746,N_43414,N_43438);
and U43747 (N_43747,N_43497,N_43354);
xnor U43748 (N_43748,N_43475,N_43448);
or U43749 (N_43749,N_43354,N_43405);
xnor U43750 (N_43750,N_43673,N_43588);
or U43751 (N_43751,N_43713,N_43674);
or U43752 (N_43752,N_43648,N_43709);
nor U43753 (N_43753,N_43604,N_43638);
nand U43754 (N_43754,N_43660,N_43542);
xor U43755 (N_43755,N_43639,N_43567);
nor U43756 (N_43756,N_43520,N_43685);
nand U43757 (N_43757,N_43668,N_43507);
or U43758 (N_43758,N_43579,N_43562);
nor U43759 (N_43759,N_43557,N_43624);
or U43760 (N_43760,N_43595,N_43530);
and U43761 (N_43761,N_43597,N_43587);
nand U43762 (N_43762,N_43523,N_43565);
and U43763 (N_43763,N_43656,N_43695);
nand U43764 (N_43764,N_43657,N_43744);
and U43765 (N_43765,N_43611,N_43641);
or U43766 (N_43766,N_43566,N_43593);
nor U43767 (N_43767,N_43727,N_43719);
nor U43768 (N_43768,N_43549,N_43669);
or U43769 (N_43769,N_43678,N_43741);
and U43770 (N_43770,N_43723,N_43555);
xnor U43771 (N_43771,N_43516,N_43578);
and U43772 (N_43772,N_43540,N_43580);
xnor U43773 (N_43773,N_43650,N_43728);
nor U43774 (N_43774,N_43550,N_43636);
or U43775 (N_43775,N_43538,N_43531);
nor U43776 (N_43776,N_43712,N_43513);
nor U43777 (N_43777,N_43598,N_43568);
or U43778 (N_43778,N_43574,N_43738);
xor U43779 (N_43779,N_43602,N_43576);
or U43780 (N_43780,N_43642,N_43635);
nor U43781 (N_43781,N_43586,N_43739);
or U43782 (N_43782,N_43608,N_43687);
xnor U43783 (N_43783,N_43688,N_43706);
xor U43784 (N_43784,N_43570,N_43690);
or U43785 (N_43785,N_43572,N_43553);
nor U43786 (N_43786,N_43505,N_43509);
nor U43787 (N_43787,N_43526,N_43670);
and U43788 (N_43788,N_43692,N_43546);
and U43789 (N_43789,N_43698,N_43734);
and U43790 (N_43790,N_43644,N_43623);
xor U43791 (N_43791,N_43679,N_43658);
or U43792 (N_43792,N_43665,N_43697);
nor U43793 (N_43793,N_43708,N_43672);
xnor U43794 (N_43794,N_43681,N_43518);
nand U43795 (N_43795,N_43514,N_43655);
xor U43796 (N_43796,N_43683,N_43680);
nor U43797 (N_43797,N_43544,N_43700);
xor U43798 (N_43798,N_43522,N_43731);
xor U43799 (N_43799,N_43605,N_43631);
nor U43800 (N_43800,N_43561,N_43637);
nand U43801 (N_43801,N_43525,N_43705);
nand U43802 (N_43802,N_43745,N_43564);
nor U43803 (N_43803,N_43533,N_43691);
nor U43804 (N_43804,N_43537,N_43626);
nand U43805 (N_43805,N_43618,N_43545);
or U43806 (N_43806,N_43515,N_43600);
and U43807 (N_43807,N_43554,N_43527);
and U43808 (N_43808,N_43502,N_43603);
nand U43809 (N_43809,N_43675,N_43649);
nand U43810 (N_43810,N_43652,N_43699);
xnor U43811 (N_43811,N_43558,N_43634);
nand U43812 (N_43812,N_43551,N_43591);
xor U43813 (N_43813,N_43590,N_43743);
xnor U43814 (N_43814,N_43614,N_43733);
and U43815 (N_43815,N_43548,N_43736);
and U43816 (N_43816,N_43726,N_43646);
xnor U43817 (N_43817,N_43569,N_43559);
xnor U43818 (N_43818,N_43735,N_43556);
or U43819 (N_43819,N_43651,N_43577);
nand U43820 (N_43820,N_43594,N_43715);
or U43821 (N_43821,N_43504,N_43500);
and U43822 (N_43822,N_43711,N_43632);
nand U43823 (N_43823,N_43647,N_43552);
nor U43824 (N_43824,N_43610,N_43663);
nand U43825 (N_43825,N_43599,N_43671);
nand U43826 (N_43826,N_43629,N_43585);
and U43827 (N_43827,N_43682,N_43529);
or U43828 (N_43828,N_43740,N_43701);
xnor U43829 (N_43829,N_43716,N_43584);
nand U43830 (N_43830,N_43640,N_43619);
and U43831 (N_43831,N_43666,N_43510);
or U43832 (N_43832,N_43547,N_43714);
and U43833 (N_43833,N_43613,N_43737);
and U43834 (N_43834,N_43702,N_43732);
xnor U43835 (N_43835,N_43645,N_43696);
nand U43836 (N_43836,N_43575,N_43524);
xor U43837 (N_43837,N_43630,N_43601);
xor U43838 (N_43838,N_43606,N_43729);
xnor U43839 (N_43839,N_43528,N_43694);
and U43840 (N_43840,N_43749,N_43703);
xnor U43841 (N_43841,N_43541,N_43581);
nor U43842 (N_43842,N_43722,N_43625);
xor U43843 (N_43843,N_43746,N_43617);
nor U43844 (N_43844,N_43654,N_43620);
xnor U43845 (N_43845,N_43536,N_43511);
nor U43846 (N_43846,N_43508,N_43539);
xor U43847 (N_43847,N_43573,N_43534);
nor U43848 (N_43848,N_43633,N_43686);
or U43849 (N_43849,N_43721,N_43506);
or U43850 (N_43850,N_43532,N_43707);
and U43851 (N_43851,N_43560,N_43677);
or U43852 (N_43852,N_43662,N_43717);
or U43853 (N_43853,N_43653,N_43503);
xor U43854 (N_43854,N_43724,N_43748);
xor U43855 (N_43855,N_43659,N_43667);
xor U43856 (N_43856,N_43718,N_43607);
nand U43857 (N_43857,N_43676,N_43612);
or U43858 (N_43858,N_43589,N_43582);
or U43859 (N_43859,N_43583,N_43571);
or U43860 (N_43860,N_43628,N_43704);
nor U43861 (N_43861,N_43720,N_43563);
xnor U43862 (N_43862,N_43622,N_43730);
nor U43863 (N_43863,N_43725,N_43664);
xnor U43864 (N_43864,N_43661,N_43742);
and U43865 (N_43865,N_43689,N_43521);
or U43866 (N_43866,N_43747,N_43643);
or U43867 (N_43867,N_43627,N_43684);
and U43868 (N_43868,N_43693,N_43535);
nand U43869 (N_43869,N_43710,N_43621);
and U43870 (N_43870,N_43512,N_43517);
nand U43871 (N_43871,N_43519,N_43501);
or U43872 (N_43872,N_43616,N_43609);
nand U43873 (N_43873,N_43592,N_43596);
nand U43874 (N_43874,N_43615,N_43543);
nand U43875 (N_43875,N_43523,N_43506);
and U43876 (N_43876,N_43502,N_43527);
and U43877 (N_43877,N_43714,N_43653);
and U43878 (N_43878,N_43630,N_43738);
xnor U43879 (N_43879,N_43573,N_43597);
and U43880 (N_43880,N_43539,N_43560);
and U43881 (N_43881,N_43533,N_43710);
and U43882 (N_43882,N_43706,N_43748);
and U43883 (N_43883,N_43666,N_43635);
nor U43884 (N_43884,N_43614,N_43540);
nand U43885 (N_43885,N_43614,N_43626);
nand U43886 (N_43886,N_43548,N_43553);
nor U43887 (N_43887,N_43680,N_43717);
xor U43888 (N_43888,N_43600,N_43716);
nand U43889 (N_43889,N_43585,N_43672);
xnor U43890 (N_43890,N_43544,N_43734);
and U43891 (N_43891,N_43707,N_43604);
or U43892 (N_43892,N_43662,N_43683);
xor U43893 (N_43893,N_43651,N_43516);
nor U43894 (N_43894,N_43544,N_43672);
and U43895 (N_43895,N_43569,N_43566);
nor U43896 (N_43896,N_43678,N_43588);
nor U43897 (N_43897,N_43689,N_43704);
xnor U43898 (N_43898,N_43523,N_43583);
xor U43899 (N_43899,N_43604,N_43699);
or U43900 (N_43900,N_43652,N_43612);
and U43901 (N_43901,N_43625,N_43718);
nand U43902 (N_43902,N_43717,N_43603);
or U43903 (N_43903,N_43617,N_43689);
nor U43904 (N_43904,N_43504,N_43553);
nor U43905 (N_43905,N_43615,N_43684);
nand U43906 (N_43906,N_43501,N_43668);
nand U43907 (N_43907,N_43520,N_43629);
nor U43908 (N_43908,N_43617,N_43729);
nor U43909 (N_43909,N_43558,N_43665);
xor U43910 (N_43910,N_43559,N_43679);
or U43911 (N_43911,N_43633,N_43727);
xnor U43912 (N_43912,N_43554,N_43731);
xor U43913 (N_43913,N_43573,N_43717);
nand U43914 (N_43914,N_43530,N_43543);
and U43915 (N_43915,N_43547,N_43600);
nand U43916 (N_43916,N_43736,N_43677);
nand U43917 (N_43917,N_43607,N_43522);
and U43918 (N_43918,N_43687,N_43639);
nor U43919 (N_43919,N_43592,N_43712);
or U43920 (N_43920,N_43516,N_43735);
and U43921 (N_43921,N_43745,N_43557);
xor U43922 (N_43922,N_43579,N_43686);
or U43923 (N_43923,N_43568,N_43700);
xor U43924 (N_43924,N_43556,N_43654);
nand U43925 (N_43925,N_43610,N_43517);
nand U43926 (N_43926,N_43732,N_43711);
and U43927 (N_43927,N_43570,N_43658);
nand U43928 (N_43928,N_43690,N_43741);
or U43929 (N_43929,N_43500,N_43645);
nand U43930 (N_43930,N_43696,N_43578);
xor U43931 (N_43931,N_43739,N_43729);
or U43932 (N_43932,N_43625,N_43542);
and U43933 (N_43933,N_43680,N_43657);
xor U43934 (N_43934,N_43540,N_43571);
or U43935 (N_43935,N_43522,N_43749);
nor U43936 (N_43936,N_43680,N_43685);
and U43937 (N_43937,N_43636,N_43613);
nor U43938 (N_43938,N_43691,N_43618);
xnor U43939 (N_43939,N_43539,N_43694);
xnor U43940 (N_43940,N_43508,N_43521);
nor U43941 (N_43941,N_43533,N_43651);
nor U43942 (N_43942,N_43580,N_43532);
or U43943 (N_43943,N_43573,N_43655);
xnor U43944 (N_43944,N_43711,N_43597);
or U43945 (N_43945,N_43713,N_43519);
or U43946 (N_43946,N_43618,N_43547);
or U43947 (N_43947,N_43731,N_43629);
nand U43948 (N_43948,N_43697,N_43630);
nor U43949 (N_43949,N_43573,N_43613);
nor U43950 (N_43950,N_43657,N_43512);
and U43951 (N_43951,N_43500,N_43624);
or U43952 (N_43952,N_43723,N_43676);
nand U43953 (N_43953,N_43578,N_43632);
nand U43954 (N_43954,N_43580,N_43616);
nand U43955 (N_43955,N_43674,N_43678);
nor U43956 (N_43956,N_43710,N_43639);
nand U43957 (N_43957,N_43733,N_43597);
nand U43958 (N_43958,N_43693,N_43602);
or U43959 (N_43959,N_43520,N_43540);
xor U43960 (N_43960,N_43640,N_43507);
and U43961 (N_43961,N_43716,N_43575);
nor U43962 (N_43962,N_43587,N_43555);
and U43963 (N_43963,N_43718,N_43723);
nor U43964 (N_43964,N_43581,N_43692);
xnor U43965 (N_43965,N_43627,N_43630);
or U43966 (N_43966,N_43713,N_43691);
xnor U43967 (N_43967,N_43565,N_43559);
nor U43968 (N_43968,N_43598,N_43629);
nor U43969 (N_43969,N_43572,N_43674);
or U43970 (N_43970,N_43637,N_43624);
xor U43971 (N_43971,N_43546,N_43686);
nor U43972 (N_43972,N_43698,N_43680);
nand U43973 (N_43973,N_43525,N_43588);
xor U43974 (N_43974,N_43619,N_43749);
nand U43975 (N_43975,N_43652,N_43558);
and U43976 (N_43976,N_43632,N_43526);
xnor U43977 (N_43977,N_43563,N_43692);
or U43978 (N_43978,N_43587,N_43739);
or U43979 (N_43979,N_43631,N_43711);
nand U43980 (N_43980,N_43583,N_43703);
nand U43981 (N_43981,N_43649,N_43619);
nand U43982 (N_43982,N_43672,N_43582);
nand U43983 (N_43983,N_43642,N_43617);
nor U43984 (N_43984,N_43742,N_43682);
or U43985 (N_43985,N_43659,N_43694);
xnor U43986 (N_43986,N_43516,N_43670);
or U43987 (N_43987,N_43544,N_43588);
xor U43988 (N_43988,N_43659,N_43679);
nor U43989 (N_43989,N_43589,N_43620);
nand U43990 (N_43990,N_43588,N_43710);
and U43991 (N_43991,N_43609,N_43581);
nor U43992 (N_43992,N_43663,N_43678);
nor U43993 (N_43993,N_43534,N_43543);
nor U43994 (N_43994,N_43659,N_43729);
xor U43995 (N_43995,N_43674,N_43607);
nand U43996 (N_43996,N_43577,N_43634);
nor U43997 (N_43997,N_43556,N_43604);
and U43998 (N_43998,N_43594,N_43657);
nand U43999 (N_43999,N_43553,N_43679);
xnor U44000 (N_44000,N_43797,N_43946);
nand U44001 (N_44001,N_43939,N_43770);
nor U44002 (N_44002,N_43938,N_43844);
xnor U44003 (N_44003,N_43789,N_43869);
nor U44004 (N_44004,N_43846,N_43786);
or U44005 (N_44005,N_43929,N_43751);
xor U44006 (N_44006,N_43949,N_43787);
nand U44007 (N_44007,N_43874,N_43912);
nand U44008 (N_44008,N_43792,N_43788);
or U44009 (N_44009,N_43858,N_43877);
or U44010 (N_44010,N_43754,N_43913);
or U44011 (N_44011,N_43785,N_43993);
nor U44012 (N_44012,N_43943,N_43979);
and U44013 (N_44013,N_43981,N_43879);
nor U44014 (N_44014,N_43933,N_43815);
or U44015 (N_44015,N_43819,N_43902);
and U44016 (N_44016,N_43821,N_43894);
nand U44017 (N_44017,N_43823,N_43764);
nand U44018 (N_44018,N_43982,N_43865);
and U44019 (N_44019,N_43759,N_43908);
nand U44020 (N_44020,N_43983,N_43899);
or U44021 (N_44021,N_43779,N_43904);
nor U44022 (N_44022,N_43996,N_43762);
xor U44023 (N_44023,N_43852,N_43833);
xor U44024 (N_44024,N_43773,N_43911);
nand U44025 (N_44025,N_43969,N_43950);
nand U44026 (N_44026,N_43980,N_43976);
or U44027 (N_44027,N_43906,N_43934);
and U44028 (N_44028,N_43897,N_43804);
nand U44029 (N_44029,N_43924,N_43992);
nand U44030 (N_44030,N_43951,N_43809);
or U44031 (N_44031,N_43935,N_43853);
xor U44032 (N_44032,N_43861,N_43842);
xnor U44033 (N_44033,N_43963,N_43891);
and U44034 (N_44034,N_43932,N_43817);
xnor U44035 (N_44035,N_43851,N_43760);
and U44036 (N_44036,N_43970,N_43953);
and U44037 (N_44037,N_43888,N_43954);
xnor U44038 (N_44038,N_43813,N_43780);
nor U44039 (N_44039,N_43881,N_43826);
xnor U44040 (N_44040,N_43837,N_43753);
or U44041 (N_44041,N_43926,N_43995);
or U44042 (N_44042,N_43986,N_43956);
and U44043 (N_44043,N_43974,N_43977);
and U44044 (N_44044,N_43893,N_43914);
nor U44045 (N_44045,N_43783,N_43776);
nor U44046 (N_44046,N_43758,N_43985);
or U44047 (N_44047,N_43838,N_43818);
nand U44048 (N_44048,N_43918,N_43820);
and U44049 (N_44049,N_43790,N_43755);
and U44050 (N_44050,N_43812,N_43972);
or U44051 (N_44051,N_43828,N_43964);
xnor U44052 (N_44052,N_43984,N_43878);
and U44053 (N_44053,N_43973,N_43855);
or U44054 (N_44054,N_43774,N_43859);
or U44055 (N_44055,N_43756,N_43798);
xor U44056 (N_44056,N_43942,N_43795);
xnor U44057 (N_44057,N_43998,N_43917);
nand U44058 (N_44058,N_43771,N_43763);
xnor U44059 (N_44059,N_43937,N_43960);
nand U44060 (N_44060,N_43827,N_43948);
nand U44061 (N_44061,N_43752,N_43957);
or U44062 (N_44062,N_43947,N_43940);
xor U44063 (N_44063,N_43840,N_43885);
or U44064 (N_44064,N_43890,N_43799);
nor U44065 (N_44065,N_43843,N_43968);
xnor U44066 (N_44066,N_43873,N_43801);
or U44067 (N_44067,N_43903,N_43772);
nor U44068 (N_44068,N_43868,N_43781);
xnor U44069 (N_44069,N_43931,N_43794);
and U44070 (N_44070,N_43830,N_43769);
or U44071 (N_44071,N_43850,N_43866);
or U44072 (N_44072,N_43997,N_43848);
and U44073 (N_44073,N_43909,N_43936);
and U44074 (N_44074,N_43962,N_43777);
xnor U44075 (N_44075,N_43845,N_43990);
xnor U44076 (N_44076,N_43775,N_43849);
or U44077 (N_44077,N_43805,N_43889);
nor U44078 (N_44078,N_43808,N_43925);
nand U44079 (N_44079,N_43967,N_43999);
or U44080 (N_44080,N_43806,N_43831);
nor U44081 (N_44081,N_43988,N_43778);
nand U44082 (N_44082,N_43887,N_43901);
nor U44083 (N_44083,N_43895,N_43807);
and U44084 (N_44084,N_43860,N_43814);
nand U44085 (N_44085,N_43768,N_43898);
nand U44086 (N_44086,N_43919,N_43886);
or U44087 (N_44087,N_43765,N_43870);
nor U44088 (N_44088,N_43875,N_43978);
or U44089 (N_44089,N_43791,N_43923);
or U44090 (N_44090,N_43958,N_43989);
nor U44091 (N_44091,N_43862,N_43796);
nor U44092 (N_44092,N_43952,N_43835);
xnor U44093 (N_44093,N_43959,N_43782);
or U44094 (N_44094,N_43955,N_43994);
nand U44095 (N_44095,N_43905,N_43965);
nor U44096 (N_44096,N_43834,N_43971);
nand U44097 (N_44097,N_43810,N_43857);
nand U44098 (N_44098,N_43927,N_43761);
and U44099 (N_44099,N_43841,N_43863);
xnor U44100 (N_44100,N_43871,N_43847);
and U44101 (N_44101,N_43944,N_43802);
or U44102 (N_44102,N_43872,N_43816);
xor U44103 (N_44103,N_43928,N_43856);
xnor U44104 (N_44104,N_43800,N_43945);
nor U44105 (N_44105,N_43864,N_43824);
nand U44106 (N_44106,N_43896,N_43915);
nand U44107 (N_44107,N_43922,N_43910);
nand U44108 (N_44108,N_43811,N_43975);
nor U44109 (N_44109,N_43991,N_43907);
xnor U44110 (N_44110,N_43766,N_43803);
nor U44111 (N_44111,N_43793,N_43750);
or U44112 (N_44112,N_43941,N_43839);
and U44113 (N_44113,N_43825,N_43987);
and U44114 (N_44114,N_43876,N_43884);
nor U44115 (N_44115,N_43829,N_43892);
and U44116 (N_44116,N_43822,N_43867);
xnor U44117 (N_44117,N_43757,N_43854);
nor U44118 (N_44118,N_43836,N_43920);
nor U44119 (N_44119,N_43921,N_43784);
nand U44120 (N_44120,N_43767,N_43880);
or U44121 (N_44121,N_43961,N_43930);
or U44122 (N_44122,N_43832,N_43900);
or U44123 (N_44123,N_43916,N_43882);
and U44124 (N_44124,N_43883,N_43966);
and U44125 (N_44125,N_43772,N_43913);
or U44126 (N_44126,N_43840,N_43878);
and U44127 (N_44127,N_43959,N_43947);
or U44128 (N_44128,N_43876,N_43798);
and U44129 (N_44129,N_43803,N_43779);
xnor U44130 (N_44130,N_43876,N_43988);
xor U44131 (N_44131,N_43873,N_43957);
nor U44132 (N_44132,N_43837,N_43798);
xor U44133 (N_44133,N_43941,N_43787);
and U44134 (N_44134,N_43947,N_43784);
xnor U44135 (N_44135,N_43892,N_43868);
xnor U44136 (N_44136,N_43891,N_43836);
xnor U44137 (N_44137,N_43973,N_43927);
and U44138 (N_44138,N_43996,N_43985);
nor U44139 (N_44139,N_43899,N_43809);
and U44140 (N_44140,N_43805,N_43769);
nor U44141 (N_44141,N_43763,N_43851);
xor U44142 (N_44142,N_43895,N_43862);
or U44143 (N_44143,N_43805,N_43753);
nand U44144 (N_44144,N_43915,N_43824);
nand U44145 (N_44145,N_43792,N_43963);
nor U44146 (N_44146,N_43895,N_43898);
xor U44147 (N_44147,N_43795,N_43963);
or U44148 (N_44148,N_43914,N_43775);
and U44149 (N_44149,N_43856,N_43943);
xnor U44150 (N_44150,N_43965,N_43994);
and U44151 (N_44151,N_43776,N_43831);
and U44152 (N_44152,N_43911,N_43961);
or U44153 (N_44153,N_43850,N_43891);
nand U44154 (N_44154,N_43877,N_43989);
xnor U44155 (N_44155,N_43949,N_43777);
and U44156 (N_44156,N_43859,N_43954);
xor U44157 (N_44157,N_43867,N_43943);
nor U44158 (N_44158,N_43765,N_43773);
xnor U44159 (N_44159,N_43861,N_43953);
nand U44160 (N_44160,N_43831,N_43889);
xor U44161 (N_44161,N_43997,N_43870);
or U44162 (N_44162,N_43798,N_43975);
xor U44163 (N_44163,N_43829,N_43822);
or U44164 (N_44164,N_43983,N_43796);
xor U44165 (N_44165,N_43785,N_43944);
or U44166 (N_44166,N_43869,N_43944);
nand U44167 (N_44167,N_43824,N_43793);
or U44168 (N_44168,N_43918,N_43751);
or U44169 (N_44169,N_43821,N_43811);
nand U44170 (N_44170,N_43959,N_43955);
and U44171 (N_44171,N_43926,N_43754);
nand U44172 (N_44172,N_43944,N_43988);
and U44173 (N_44173,N_43927,N_43948);
nand U44174 (N_44174,N_43752,N_43760);
xor U44175 (N_44175,N_43784,N_43995);
xnor U44176 (N_44176,N_43887,N_43953);
and U44177 (N_44177,N_43816,N_43949);
nor U44178 (N_44178,N_43893,N_43787);
and U44179 (N_44179,N_43803,N_43791);
nand U44180 (N_44180,N_43979,N_43843);
xor U44181 (N_44181,N_43906,N_43975);
nand U44182 (N_44182,N_43778,N_43925);
and U44183 (N_44183,N_43819,N_43973);
nand U44184 (N_44184,N_43774,N_43758);
xnor U44185 (N_44185,N_43775,N_43772);
xnor U44186 (N_44186,N_43899,N_43798);
xor U44187 (N_44187,N_43813,N_43938);
or U44188 (N_44188,N_43833,N_43909);
nand U44189 (N_44189,N_43946,N_43823);
or U44190 (N_44190,N_43922,N_43999);
or U44191 (N_44191,N_43956,N_43761);
xnor U44192 (N_44192,N_43923,N_43982);
or U44193 (N_44193,N_43847,N_43981);
nand U44194 (N_44194,N_43787,N_43907);
xnor U44195 (N_44195,N_43943,N_43934);
nor U44196 (N_44196,N_43772,N_43992);
and U44197 (N_44197,N_43953,N_43932);
and U44198 (N_44198,N_43945,N_43892);
nor U44199 (N_44199,N_43965,N_43937);
xor U44200 (N_44200,N_43938,N_43980);
xor U44201 (N_44201,N_43899,N_43857);
nand U44202 (N_44202,N_43988,N_43952);
xnor U44203 (N_44203,N_43833,N_43904);
xor U44204 (N_44204,N_43962,N_43931);
nand U44205 (N_44205,N_43902,N_43945);
xor U44206 (N_44206,N_43908,N_43829);
nand U44207 (N_44207,N_43867,N_43801);
nor U44208 (N_44208,N_43788,N_43995);
nand U44209 (N_44209,N_43932,N_43956);
xnor U44210 (N_44210,N_43901,N_43763);
and U44211 (N_44211,N_43781,N_43940);
and U44212 (N_44212,N_43941,N_43892);
and U44213 (N_44213,N_43921,N_43873);
nand U44214 (N_44214,N_43832,N_43914);
or U44215 (N_44215,N_43877,N_43772);
nand U44216 (N_44216,N_43829,N_43992);
or U44217 (N_44217,N_43813,N_43858);
xnor U44218 (N_44218,N_43783,N_43828);
or U44219 (N_44219,N_43880,N_43758);
xnor U44220 (N_44220,N_43923,N_43929);
nor U44221 (N_44221,N_43828,N_43959);
nor U44222 (N_44222,N_43817,N_43973);
or U44223 (N_44223,N_43839,N_43825);
nor U44224 (N_44224,N_43856,N_43766);
nor U44225 (N_44225,N_43933,N_43777);
and U44226 (N_44226,N_43996,N_43828);
nor U44227 (N_44227,N_43876,N_43768);
and U44228 (N_44228,N_43944,N_43859);
nand U44229 (N_44229,N_43982,N_43830);
nand U44230 (N_44230,N_43957,N_43882);
nand U44231 (N_44231,N_43822,N_43795);
and U44232 (N_44232,N_43941,N_43960);
nor U44233 (N_44233,N_43998,N_43808);
or U44234 (N_44234,N_43979,N_43855);
and U44235 (N_44235,N_43949,N_43940);
nor U44236 (N_44236,N_43918,N_43826);
and U44237 (N_44237,N_43785,N_43820);
or U44238 (N_44238,N_43850,N_43843);
or U44239 (N_44239,N_43979,N_43879);
nand U44240 (N_44240,N_43854,N_43957);
xnor U44241 (N_44241,N_43774,N_43876);
nor U44242 (N_44242,N_43977,N_43812);
nor U44243 (N_44243,N_43791,N_43785);
nand U44244 (N_44244,N_43987,N_43960);
and U44245 (N_44245,N_43825,N_43809);
nor U44246 (N_44246,N_43957,N_43999);
xnor U44247 (N_44247,N_43999,N_43803);
nor U44248 (N_44248,N_43924,N_43905);
or U44249 (N_44249,N_43890,N_43860);
or U44250 (N_44250,N_44094,N_44037);
xnor U44251 (N_44251,N_44022,N_44114);
nand U44252 (N_44252,N_44243,N_44183);
and U44253 (N_44253,N_44069,N_44159);
nor U44254 (N_44254,N_44075,N_44098);
nor U44255 (N_44255,N_44084,N_44121);
and U44256 (N_44256,N_44210,N_44126);
xor U44257 (N_44257,N_44051,N_44237);
xor U44258 (N_44258,N_44004,N_44007);
nand U44259 (N_44259,N_44165,N_44133);
xor U44260 (N_44260,N_44209,N_44081);
and U44261 (N_44261,N_44052,N_44003);
or U44262 (N_44262,N_44247,N_44025);
or U44263 (N_44263,N_44021,N_44205);
nor U44264 (N_44264,N_44031,N_44236);
nand U44265 (N_44265,N_44002,N_44218);
xnor U44266 (N_44266,N_44189,N_44244);
nand U44267 (N_44267,N_44093,N_44203);
nand U44268 (N_44268,N_44235,N_44169);
or U44269 (N_44269,N_44234,N_44162);
or U44270 (N_44270,N_44113,N_44194);
and U44271 (N_44271,N_44129,N_44134);
or U44272 (N_44272,N_44005,N_44196);
and U44273 (N_44273,N_44061,N_44174);
and U44274 (N_44274,N_44228,N_44156);
xnor U44275 (N_44275,N_44208,N_44153);
and U44276 (N_44276,N_44248,N_44230);
xnor U44277 (N_44277,N_44180,N_44015);
xor U44278 (N_44278,N_44170,N_44006);
nand U44279 (N_44279,N_44016,N_44112);
nor U44280 (N_44280,N_44138,N_44017);
xnor U44281 (N_44281,N_44225,N_44188);
nor U44282 (N_44282,N_44168,N_44144);
nor U44283 (N_44283,N_44122,N_44148);
or U44284 (N_44284,N_44000,N_44186);
and U44285 (N_44285,N_44009,N_44106);
nand U44286 (N_44286,N_44166,N_44101);
nand U44287 (N_44287,N_44105,N_44115);
and U44288 (N_44288,N_44027,N_44139);
nor U44289 (N_44289,N_44146,N_44095);
or U44290 (N_44290,N_44001,N_44010);
and U44291 (N_44291,N_44085,N_44012);
nand U44292 (N_44292,N_44019,N_44103);
nand U44293 (N_44293,N_44145,N_44076);
or U44294 (N_44294,N_44249,N_44163);
nand U44295 (N_44295,N_44053,N_44035);
xor U44296 (N_44296,N_44033,N_44050);
nor U44297 (N_44297,N_44111,N_44072);
nor U44298 (N_44298,N_44063,N_44044);
nand U44299 (N_44299,N_44046,N_44147);
xor U44300 (N_44300,N_44107,N_44078);
xnor U44301 (N_44301,N_44200,N_44212);
nor U44302 (N_44302,N_44067,N_44181);
nor U44303 (N_44303,N_44023,N_44074);
or U44304 (N_44304,N_44219,N_44008);
nand U44305 (N_44305,N_44223,N_44086);
xnor U44306 (N_44306,N_44216,N_44062);
or U44307 (N_44307,N_44018,N_44043);
nor U44308 (N_44308,N_44201,N_44057);
xor U44309 (N_44309,N_44211,N_44049);
and U44310 (N_44310,N_44020,N_44193);
xnor U44311 (N_44311,N_44179,N_44150);
xor U44312 (N_44312,N_44065,N_44124);
xor U44313 (N_44313,N_44042,N_44140);
nor U44314 (N_44314,N_44048,N_44118);
and U44315 (N_44315,N_44036,N_44161);
and U44316 (N_44316,N_44026,N_44071);
nand U44317 (N_44317,N_44120,N_44029);
nand U44318 (N_44318,N_44088,N_44152);
and U44319 (N_44319,N_44242,N_44055);
xor U44320 (N_44320,N_44030,N_44059);
or U44321 (N_44321,N_44039,N_44083);
xnor U44322 (N_44322,N_44233,N_44082);
and U44323 (N_44323,N_44038,N_44239);
and U44324 (N_44324,N_44176,N_44227);
nand U44325 (N_44325,N_44117,N_44232);
or U44326 (N_44326,N_44104,N_44079);
and U44327 (N_44327,N_44056,N_44131);
xor U44328 (N_44328,N_44155,N_44217);
and U44329 (N_44329,N_44190,N_44167);
nand U44330 (N_44330,N_44191,N_44206);
or U44331 (N_44331,N_44178,N_44199);
and U44332 (N_44332,N_44245,N_44041);
nor U44333 (N_44333,N_44097,N_44198);
and U44334 (N_44334,N_44102,N_44185);
or U44335 (N_44335,N_44207,N_44142);
or U44336 (N_44336,N_44215,N_44011);
nand U44337 (N_44337,N_44034,N_44220);
and U44338 (N_44338,N_44164,N_44116);
nand U44339 (N_44339,N_44032,N_44092);
or U44340 (N_44340,N_44157,N_44123);
or U44341 (N_44341,N_44132,N_44202);
or U44342 (N_44342,N_44240,N_44060);
and U44343 (N_44343,N_44231,N_44171);
xnor U44344 (N_44344,N_44089,N_44028);
and U44345 (N_44345,N_44110,N_44058);
or U44346 (N_44346,N_44136,N_44172);
nor U44347 (N_44347,N_44125,N_44135);
xnor U44348 (N_44348,N_44214,N_44246);
nand U44349 (N_44349,N_44158,N_44100);
nor U44350 (N_44350,N_44226,N_44087);
nor U44351 (N_44351,N_44229,N_44222);
and U44352 (N_44352,N_44127,N_44221);
nand U44353 (N_44353,N_44177,N_44160);
nor U44354 (N_44354,N_44192,N_44197);
nand U44355 (N_44355,N_44224,N_44213);
and U44356 (N_44356,N_44014,N_44064);
nor U44357 (N_44357,N_44070,N_44195);
xor U44358 (N_44358,N_44149,N_44040);
and U44359 (N_44359,N_44241,N_44068);
or U44360 (N_44360,N_44154,N_44045);
and U44361 (N_44361,N_44099,N_44108);
and U44362 (N_44362,N_44238,N_44184);
or U44363 (N_44363,N_44054,N_44119);
nor U44364 (N_44364,N_44024,N_44073);
and U44365 (N_44365,N_44047,N_44187);
or U44366 (N_44366,N_44091,N_44143);
or U44367 (N_44367,N_44173,N_44066);
nand U44368 (N_44368,N_44077,N_44175);
nand U44369 (N_44369,N_44141,N_44137);
and U44370 (N_44370,N_44109,N_44151);
xor U44371 (N_44371,N_44090,N_44130);
and U44372 (N_44372,N_44204,N_44013);
xnor U44373 (N_44373,N_44182,N_44128);
nor U44374 (N_44374,N_44080,N_44096);
or U44375 (N_44375,N_44218,N_44230);
nor U44376 (N_44376,N_44078,N_44024);
or U44377 (N_44377,N_44143,N_44193);
and U44378 (N_44378,N_44191,N_44232);
or U44379 (N_44379,N_44212,N_44224);
and U44380 (N_44380,N_44240,N_44001);
xor U44381 (N_44381,N_44126,N_44177);
or U44382 (N_44382,N_44141,N_44076);
nand U44383 (N_44383,N_44072,N_44095);
nor U44384 (N_44384,N_44059,N_44069);
and U44385 (N_44385,N_44159,N_44017);
and U44386 (N_44386,N_44063,N_44222);
or U44387 (N_44387,N_44133,N_44136);
or U44388 (N_44388,N_44045,N_44023);
and U44389 (N_44389,N_44229,N_44146);
or U44390 (N_44390,N_44154,N_44249);
or U44391 (N_44391,N_44245,N_44113);
nand U44392 (N_44392,N_44094,N_44181);
nand U44393 (N_44393,N_44037,N_44135);
and U44394 (N_44394,N_44003,N_44134);
xor U44395 (N_44395,N_44111,N_44211);
nor U44396 (N_44396,N_44033,N_44219);
and U44397 (N_44397,N_44007,N_44129);
or U44398 (N_44398,N_44225,N_44029);
nand U44399 (N_44399,N_44024,N_44217);
xor U44400 (N_44400,N_44114,N_44246);
nor U44401 (N_44401,N_44200,N_44211);
nor U44402 (N_44402,N_44022,N_44156);
and U44403 (N_44403,N_44211,N_44217);
xor U44404 (N_44404,N_44071,N_44054);
or U44405 (N_44405,N_44207,N_44094);
or U44406 (N_44406,N_44045,N_44060);
and U44407 (N_44407,N_44205,N_44114);
xnor U44408 (N_44408,N_44019,N_44147);
and U44409 (N_44409,N_44117,N_44156);
nor U44410 (N_44410,N_44028,N_44231);
xor U44411 (N_44411,N_44108,N_44242);
and U44412 (N_44412,N_44078,N_44068);
and U44413 (N_44413,N_44015,N_44172);
or U44414 (N_44414,N_44029,N_44047);
and U44415 (N_44415,N_44065,N_44218);
nand U44416 (N_44416,N_44232,N_44129);
or U44417 (N_44417,N_44117,N_44186);
nor U44418 (N_44418,N_44063,N_44248);
or U44419 (N_44419,N_44101,N_44120);
nand U44420 (N_44420,N_44003,N_44160);
nor U44421 (N_44421,N_44195,N_44007);
xor U44422 (N_44422,N_44155,N_44235);
xnor U44423 (N_44423,N_44125,N_44233);
xnor U44424 (N_44424,N_44047,N_44107);
nand U44425 (N_44425,N_44111,N_44034);
nor U44426 (N_44426,N_44000,N_44240);
and U44427 (N_44427,N_44035,N_44156);
or U44428 (N_44428,N_44173,N_44020);
xnor U44429 (N_44429,N_44126,N_44230);
xnor U44430 (N_44430,N_44223,N_44180);
or U44431 (N_44431,N_44199,N_44050);
and U44432 (N_44432,N_44128,N_44246);
nor U44433 (N_44433,N_44217,N_44019);
nand U44434 (N_44434,N_44127,N_44249);
xor U44435 (N_44435,N_44066,N_44074);
and U44436 (N_44436,N_44218,N_44016);
and U44437 (N_44437,N_44050,N_44109);
or U44438 (N_44438,N_44077,N_44127);
nand U44439 (N_44439,N_44083,N_44073);
or U44440 (N_44440,N_44128,N_44179);
nand U44441 (N_44441,N_44139,N_44053);
or U44442 (N_44442,N_44051,N_44094);
or U44443 (N_44443,N_44135,N_44038);
nand U44444 (N_44444,N_44015,N_44092);
or U44445 (N_44445,N_44021,N_44022);
xnor U44446 (N_44446,N_44234,N_44021);
nor U44447 (N_44447,N_44117,N_44075);
nand U44448 (N_44448,N_44166,N_44095);
or U44449 (N_44449,N_44213,N_44074);
xnor U44450 (N_44450,N_44181,N_44026);
nand U44451 (N_44451,N_44155,N_44056);
or U44452 (N_44452,N_44158,N_44081);
or U44453 (N_44453,N_44080,N_44177);
nor U44454 (N_44454,N_44235,N_44070);
nor U44455 (N_44455,N_44142,N_44137);
or U44456 (N_44456,N_44240,N_44002);
and U44457 (N_44457,N_44038,N_44014);
nor U44458 (N_44458,N_44164,N_44087);
nor U44459 (N_44459,N_44046,N_44048);
nand U44460 (N_44460,N_44174,N_44130);
nand U44461 (N_44461,N_44203,N_44022);
xnor U44462 (N_44462,N_44163,N_44105);
nand U44463 (N_44463,N_44057,N_44082);
nand U44464 (N_44464,N_44109,N_44090);
and U44465 (N_44465,N_44248,N_44188);
nor U44466 (N_44466,N_44127,N_44218);
xor U44467 (N_44467,N_44214,N_44045);
or U44468 (N_44468,N_44102,N_44078);
nor U44469 (N_44469,N_44223,N_44036);
and U44470 (N_44470,N_44036,N_44160);
nor U44471 (N_44471,N_44196,N_44204);
or U44472 (N_44472,N_44063,N_44052);
or U44473 (N_44473,N_44191,N_44133);
nor U44474 (N_44474,N_44214,N_44096);
nand U44475 (N_44475,N_44230,N_44054);
and U44476 (N_44476,N_44208,N_44004);
or U44477 (N_44477,N_44002,N_44145);
and U44478 (N_44478,N_44140,N_44019);
nor U44479 (N_44479,N_44001,N_44025);
and U44480 (N_44480,N_44218,N_44200);
and U44481 (N_44481,N_44197,N_44011);
or U44482 (N_44482,N_44060,N_44036);
xnor U44483 (N_44483,N_44004,N_44220);
nand U44484 (N_44484,N_44072,N_44114);
nor U44485 (N_44485,N_44013,N_44115);
xor U44486 (N_44486,N_44019,N_44242);
nand U44487 (N_44487,N_44210,N_44092);
xor U44488 (N_44488,N_44048,N_44133);
xnor U44489 (N_44489,N_44176,N_44043);
nand U44490 (N_44490,N_44218,N_44051);
xnor U44491 (N_44491,N_44241,N_44092);
nor U44492 (N_44492,N_44131,N_44080);
nand U44493 (N_44493,N_44095,N_44057);
nand U44494 (N_44494,N_44005,N_44161);
or U44495 (N_44495,N_44184,N_44065);
or U44496 (N_44496,N_44088,N_44179);
xnor U44497 (N_44497,N_44120,N_44113);
or U44498 (N_44498,N_44035,N_44199);
xor U44499 (N_44499,N_44070,N_44162);
nand U44500 (N_44500,N_44272,N_44421);
and U44501 (N_44501,N_44422,N_44328);
nand U44502 (N_44502,N_44382,N_44292);
xor U44503 (N_44503,N_44322,N_44418);
xor U44504 (N_44504,N_44323,N_44487);
xnor U44505 (N_44505,N_44486,N_44398);
nor U44506 (N_44506,N_44330,N_44415);
or U44507 (N_44507,N_44493,N_44408);
xnor U44508 (N_44508,N_44263,N_44468);
nor U44509 (N_44509,N_44474,N_44400);
nor U44510 (N_44510,N_44276,N_44416);
nand U44511 (N_44511,N_44495,N_44399);
nor U44512 (N_44512,N_44463,N_44369);
and U44513 (N_44513,N_44279,N_44342);
and U44514 (N_44514,N_44489,N_44447);
or U44515 (N_44515,N_44407,N_44364);
nor U44516 (N_44516,N_44443,N_44310);
and U44517 (N_44517,N_44444,N_44333);
and U44518 (N_44518,N_44395,N_44308);
nor U44519 (N_44519,N_44290,N_44402);
or U44520 (N_44520,N_44485,N_44451);
or U44521 (N_44521,N_44484,N_44355);
nor U44522 (N_44522,N_44258,N_44339);
nand U44523 (N_44523,N_44315,N_44265);
xnor U44524 (N_44524,N_44331,N_44388);
and U44525 (N_44525,N_44394,N_44427);
xnor U44526 (N_44526,N_44282,N_44285);
nor U44527 (N_44527,N_44304,N_44450);
xor U44528 (N_44528,N_44481,N_44251);
xor U44529 (N_44529,N_44419,N_44326);
xnor U44530 (N_44530,N_44437,N_44253);
and U44531 (N_44531,N_44381,N_44476);
and U44532 (N_44532,N_44329,N_44383);
nand U44533 (N_44533,N_44306,N_44371);
or U44534 (N_44534,N_44291,N_44464);
nor U44535 (N_44535,N_44467,N_44337);
nor U44536 (N_44536,N_44363,N_44286);
xnor U44537 (N_44537,N_44365,N_44469);
or U44538 (N_44538,N_44472,N_44344);
nand U44539 (N_44539,N_44411,N_44455);
and U44540 (N_44540,N_44403,N_44492);
or U44541 (N_44541,N_44275,N_44338);
nor U44542 (N_44542,N_44378,N_44314);
nor U44543 (N_44543,N_44499,N_44352);
nor U44544 (N_44544,N_44312,N_44264);
or U44545 (N_44545,N_44423,N_44387);
nor U44546 (N_44546,N_44336,N_44321);
nand U44547 (N_44547,N_44431,N_44268);
xor U44548 (N_44548,N_44300,N_44262);
or U44549 (N_44549,N_44483,N_44307);
nand U44550 (N_44550,N_44457,N_44305);
and U44551 (N_44551,N_44488,N_44494);
and U44552 (N_44552,N_44479,N_44462);
xnor U44553 (N_44553,N_44277,N_44346);
or U44554 (N_44554,N_44368,N_44362);
xnor U44555 (N_44555,N_44319,N_44347);
and U44556 (N_44556,N_44317,N_44295);
nand U44557 (N_44557,N_44456,N_44458);
nor U44558 (N_44558,N_44377,N_44391);
or U44559 (N_44559,N_44303,N_44257);
or U44560 (N_44560,N_44281,N_44446);
nand U44561 (N_44561,N_44430,N_44298);
and U44562 (N_44562,N_44490,N_44414);
or U44563 (N_44563,N_44397,N_44366);
nand U44564 (N_44564,N_44357,N_44280);
nand U44565 (N_44565,N_44287,N_44324);
or U44566 (N_44566,N_44360,N_44250);
xnor U44567 (N_44567,N_44367,N_44433);
or U44568 (N_44568,N_44466,N_44471);
nand U44569 (N_44569,N_44335,N_44309);
and U44570 (N_44570,N_44445,N_44440);
and U44571 (N_44571,N_44498,N_44348);
xor U44572 (N_44572,N_44351,N_44278);
nand U44573 (N_44573,N_44293,N_44420);
xnor U44574 (N_44574,N_44296,N_44254);
xnor U44575 (N_44575,N_44404,N_44406);
xnor U44576 (N_44576,N_44273,N_44332);
and U44577 (N_44577,N_44269,N_44271);
nor U44578 (N_44578,N_44390,N_44497);
nand U44579 (N_44579,N_44361,N_44294);
or U44580 (N_44580,N_44349,N_44441);
or U44581 (N_44581,N_44380,N_44259);
or U44582 (N_44582,N_44318,N_44393);
xor U44583 (N_44583,N_44384,N_44410);
nor U44584 (N_44584,N_44311,N_44299);
or U44585 (N_44585,N_44386,N_44370);
or U44586 (N_44586,N_44316,N_44432);
or U44587 (N_44587,N_44412,N_44350);
or U44588 (N_44588,N_44392,N_44274);
nor U44589 (N_44589,N_44442,N_44482);
xnor U44590 (N_44590,N_44327,N_44435);
nor U44591 (N_44591,N_44425,N_44270);
or U44592 (N_44592,N_44373,N_44454);
and U44593 (N_44593,N_44256,N_44448);
or U44594 (N_44594,N_44459,N_44429);
or U44595 (N_44595,N_44473,N_44266);
xnor U44596 (N_44596,N_44372,N_44358);
or U44597 (N_44597,N_44436,N_44353);
nand U44598 (N_44598,N_44405,N_44428);
xor U44599 (N_44599,N_44284,N_44267);
or U44600 (N_44600,N_44374,N_44460);
xnor U44601 (N_44601,N_44341,N_44434);
nor U44602 (N_44602,N_44452,N_44356);
and U44603 (N_44603,N_44465,N_44261);
nand U44604 (N_44604,N_44480,N_44354);
nor U44605 (N_44605,N_44320,N_44334);
or U44606 (N_44606,N_44413,N_44375);
or U44607 (N_44607,N_44477,N_44289);
nor U44608 (N_44608,N_44345,N_44453);
nor U44609 (N_44609,N_44343,N_44470);
xnor U44610 (N_44610,N_44396,N_44385);
nand U44611 (N_44611,N_44301,N_44288);
nand U44612 (N_44612,N_44496,N_44449);
xnor U44613 (N_44613,N_44283,N_44426);
xor U44614 (N_44614,N_44376,N_44389);
xor U44615 (N_44615,N_44252,N_44461);
or U44616 (N_44616,N_44359,N_44439);
or U44617 (N_44617,N_44438,N_44302);
nor U44618 (N_44618,N_44491,N_44379);
nand U44619 (N_44619,N_44325,N_44313);
nor U44620 (N_44620,N_44475,N_44417);
or U44621 (N_44621,N_44260,N_44401);
or U44622 (N_44622,N_44340,N_44255);
and U44623 (N_44623,N_44409,N_44424);
and U44624 (N_44624,N_44297,N_44478);
and U44625 (N_44625,N_44485,N_44378);
and U44626 (N_44626,N_44478,N_44341);
nand U44627 (N_44627,N_44320,N_44479);
or U44628 (N_44628,N_44308,N_44349);
nand U44629 (N_44629,N_44360,N_44304);
nor U44630 (N_44630,N_44487,N_44419);
nor U44631 (N_44631,N_44498,N_44259);
xnor U44632 (N_44632,N_44461,N_44380);
xor U44633 (N_44633,N_44294,N_44321);
and U44634 (N_44634,N_44488,N_44256);
nand U44635 (N_44635,N_44264,N_44377);
nand U44636 (N_44636,N_44334,N_44376);
and U44637 (N_44637,N_44373,N_44332);
xnor U44638 (N_44638,N_44489,N_44459);
or U44639 (N_44639,N_44394,N_44495);
nand U44640 (N_44640,N_44477,N_44424);
or U44641 (N_44641,N_44433,N_44380);
xnor U44642 (N_44642,N_44359,N_44444);
nand U44643 (N_44643,N_44479,N_44307);
nor U44644 (N_44644,N_44421,N_44382);
or U44645 (N_44645,N_44287,N_44319);
nand U44646 (N_44646,N_44453,N_44404);
xnor U44647 (N_44647,N_44430,N_44446);
nor U44648 (N_44648,N_44422,N_44463);
nand U44649 (N_44649,N_44412,N_44390);
or U44650 (N_44650,N_44389,N_44266);
nor U44651 (N_44651,N_44449,N_44453);
and U44652 (N_44652,N_44375,N_44465);
and U44653 (N_44653,N_44254,N_44308);
nor U44654 (N_44654,N_44409,N_44418);
nor U44655 (N_44655,N_44339,N_44489);
nand U44656 (N_44656,N_44280,N_44498);
and U44657 (N_44657,N_44264,N_44417);
or U44658 (N_44658,N_44314,N_44418);
xor U44659 (N_44659,N_44448,N_44309);
nor U44660 (N_44660,N_44477,N_44333);
xor U44661 (N_44661,N_44295,N_44259);
xor U44662 (N_44662,N_44368,N_44387);
or U44663 (N_44663,N_44349,N_44297);
nand U44664 (N_44664,N_44327,N_44270);
and U44665 (N_44665,N_44393,N_44323);
nand U44666 (N_44666,N_44382,N_44443);
and U44667 (N_44667,N_44348,N_44399);
xnor U44668 (N_44668,N_44411,N_44424);
xor U44669 (N_44669,N_44310,N_44315);
nor U44670 (N_44670,N_44494,N_44468);
xor U44671 (N_44671,N_44334,N_44327);
nand U44672 (N_44672,N_44434,N_44327);
nor U44673 (N_44673,N_44308,N_44321);
and U44674 (N_44674,N_44395,N_44445);
xor U44675 (N_44675,N_44418,N_44292);
nor U44676 (N_44676,N_44368,N_44396);
nand U44677 (N_44677,N_44296,N_44499);
xor U44678 (N_44678,N_44288,N_44322);
xor U44679 (N_44679,N_44428,N_44363);
or U44680 (N_44680,N_44268,N_44375);
nor U44681 (N_44681,N_44390,N_44264);
and U44682 (N_44682,N_44482,N_44343);
nor U44683 (N_44683,N_44311,N_44499);
xor U44684 (N_44684,N_44482,N_44372);
and U44685 (N_44685,N_44376,N_44312);
xnor U44686 (N_44686,N_44417,N_44322);
and U44687 (N_44687,N_44484,N_44311);
nand U44688 (N_44688,N_44367,N_44476);
or U44689 (N_44689,N_44366,N_44370);
nand U44690 (N_44690,N_44281,N_44408);
or U44691 (N_44691,N_44397,N_44346);
nand U44692 (N_44692,N_44490,N_44416);
and U44693 (N_44693,N_44332,N_44384);
nand U44694 (N_44694,N_44294,N_44329);
xor U44695 (N_44695,N_44372,N_44348);
xnor U44696 (N_44696,N_44262,N_44367);
nand U44697 (N_44697,N_44479,N_44422);
and U44698 (N_44698,N_44461,N_44399);
xor U44699 (N_44699,N_44358,N_44407);
and U44700 (N_44700,N_44283,N_44284);
and U44701 (N_44701,N_44262,N_44286);
or U44702 (N_44702,N_44446,N_44404);
nor U44703 (N_44703,N_44480,N_44470);
or U44704 (N_44704,N_44399,N_44409);
and U44705 (N_44705,N_44337,N_44297);
nand U44706 (N_44706,N_44426,N_44425);
xor U44707 (N_44707,N_44308,N_44397);
and U44708 (N_44708,N_44475,N_44303);
and U44709 (N_44709,N_44301,N_44473);
xor U44710 (N_44710,N_44324,N_44470);
or U44711 (N_44711,N_44263,N_44273);
nor U44712 (N_44712,N_44334,N_44452);
nor U44713 (N_44713,N_44261,N_44298);
and U44714 (N_44714,N_44363,N_44453);
nor U44715 (N_44715,N_44418,N_44284);
nand U44716 (N_44716,N_44373,N_44430);
nand U44717 (N_44717,N_44459,N_44471);
xnor U44718 (N_44718,N_44471,N_44456);
nor U44719 (N_44719,N_44263,N_44274);
nand U44720 (N_44720,N_44337,N_44437);
nor U44721 (N_44721,N_44343,N_44374);
or U44722 (N_44722,N_44389,N_44283);
xnor U44723 (N_44723,N_44370,N_44414);
or U44724 (N_44724,N_44370,N_44354);
nand U44725 (N_44725,N_44388,N_44461);
xnor U44726 (N_44726,N_44427,N_44461);
and U44727 (N_44727,N_44295,N_44366);
or U44728 (N_44728,N_44329,N_44261);
or U44729 (N_44729,N_44465,N_44251);
xnor U44730 (N_44730,N_44303,N_44355);
or U44731 (N_44731,N_44459,N_44411);
and U44732 (N_44732,N_44375,N_44372);
xor U44733 (N_44733,N_44349,N_44253);
xor U44734 (N_44734,N_44352,N_44397);
nand U44735 (N_44735,N_44323,N_44267);
or U44736 (N_44736,N_44265,N_44305);
nor U44737 (N_44737,N_44330,N_44361);
or U44738 (N_44738,N_44253,N_44270);
nand U44739 (N_44739,N_44318,N_44333);
nand U44740 (N_44740,N_44364,N_44319);
nand U44741 (N_44741,N_44396,N_44379);
nor U44742 (N_44742,N_44445,N_44435);
or U44743 (N_44743,N_44435,N_44499);
or U44744 (N_44744,N_44436,N_44333);
nor U44745 (N_44745,N_44388,N_44476);
nand U44746 (N_44746,N_44431,N_44399);
nor U44747 (N_44747,N_44266,N_44405);
nand U44748 (N_44748,N_44302,N_44336);
nand U44749 (N_44749,N_44342,N_44294);
and U44750 (N_44750,N_44618,N_44675);
nor U44751 (N_44751,N_44652,N_44678);
and U44752 (N_44752,N_44672,N_44621);
nand U44753 (N_44753,N_44550,N_44548);
xnor U44754 (N_44754,N_44643,N_44627);
xor U44755 (N_44755,N_44715,N_44654);
and U44756 (N_44756,N_44684,N_44582);
xor U44757 (N_44757,N_44543,N_44593);
and U44758 (N_44758,N_44502,N_44739);
xnor U44759 (N_44759,N_44703,N_44699);
nor U44760 (N_44760,N_44668,N_44686);
or U44761 (N_44761,N_44730,N_44748);
and U44762 (N_44762,N_44610,N_44720);
nor U44763 (N_44763,N_44580,N_44705);
or U44764 (N_44764,N_44646,N_44524);
nor U44765 (N_44765,N_44536,N_44556);
or U44766 (N_44766,N_44530,N_44619);
or U44767 (N_44767,N_44608,N_44625);
xnor U44768 (N_44768,N_44728,N_44590);
nand U44769 (N_44769,N_44641,N_44565);
nor U44770 (N_44770,N_44508,N_44596);
xor U44771 (N_44771,N_44574,N_44673);
and U44772 (N_44772,N_44642,N_44500);
nand U44773 (N_44773,N_44659,N_44712);
nand U44774 (N_44774,N_44601,N_44681);
nor U44775 (N_44775,N_44592,N_44503);
and U44776 (N_44776,N_44692,N_44611);
or U44777 (N_44777,N_44628,N_44585);
or U44778 (N_44778,N_44538,N_44507);
and U44779 (N_44779,N_44744,N_44648);
nand U44780 (N_44780,N_44521,N_44571);
nand U44781 (N_44781,N_44589,N_44525);
and U44782 (N_44782,N_44519,N_44575);
or U44783 (N_44783,N_44622,N_44526);
and U44784 (N_44784,N_44598,N_44632);
or U44785 (N_44785,N_44722,N_44616);
xnor U44786 (N_44786,N_44595,N_44513);
xor U44787 (N_44787,N_44661,N_44636);
xnor U44788 (N_44788,N_44662,N_44564);
nor U44789 (N_44789,N_44742,N_44649);
or U44790 (N_44790,N_44558,N_44572);
or U44791 (N_44791,N_44510,N_44653);
nor U44792 (N_44792,N_44749,N_44562);
or U44793 (N_44793,N_44685,N_44644);
or U44794 (N_44794,N_44604,N_44549);
nand U44795 (N_44795,N_44542,N_44617);
nand U44796 (N_44796,N_44613,N_44734);
or U44797 (N_44797,N_44566,N_44696);
xnor U44798 (N_44798,N_44591,N_44745);
nand U44799 (N_44799,N_44506,N_44724);
nor U44800 (N_44800,N_44537,N_44573);
nor U44801 (N_44801,N_44509,N_44717);
or U44802 (N_44802,N_44697,N_44732);
or U44803 (N_44803,N_44553,N_44588);
and U44804 (N_44804,N_44682,N_44624);
nor U44805 (N_44805,N_44719,N_44711);
xor U44806 (N_44806,N_44505,N_44532);
nand U44807 (N_44807,N_44586,N_44743);
nand U44808 (N_44808,N_44637,N_44679);
nand U44809 (N_44809,N_44576,N_44747);
xor U44810 (N_44810,N_44688,N_44516);
or U44811 (N_44811,N_44638,N_44523);
and U44812 (N_44812,N_44714,N_44657);
and U44813 (N_44813,N_44706,N_44623);
xor U44814 (N_44814,N_44708,N_44647);
or U44815 (N_44815,N_44725,N_44680);
or U44816 (N_44816,N_44658,N_44735);
xnor U44817 (N_44817,N_44701,N_44540);
or U44818 (N_44818,N_44667,N_44609);
xor U44819 (N_44819,N_44693,N_44671);
nor U44820 (N_44820,N_44517,N_44736);
xor U44821 (N_44821,N_44718,N_44674);
or U44822 (N_44822,N_44529,N_44710);
or U44823 (N_44823,N_44547,N_44666);
nor U44824 (N_44824,N_44731,N_44607);
xnor U44825 (N_44825,N_44512,N_44631);
and U44826 (N_44826,N_44534,N_44716);
nor U44827 (N_44827,N_44560,N_44511);
nand U44828 (N_44828,N_44713,N_44727);
nand U44829 (N_44829,N_44614,N_44528);
and U44830 (N_44830,N_44602,N_44501);
or U44831 (N_44831,N_44737,N_44746);
nand U44832 (N_44832,N_44570,N_44545);
xor U44833 (N_44833,N_44522,N_44635);
xor U44834 (N_44834,N_44723,N_44660);
nand U44835 (N_44835,N_44704,N_44656);
xor U44836 (N_44836,N_44615,N_44640);
nand U44837 (N_44837,N_44541,N_44535);
nor U44838 (N_44838,N_44683,N_44733);
or U44839 (N_44839,N_44605,N_44515);
or U44840 (N_44840,N_44630,N_44677);
and U44841 (N_44841,N_44729,N_44544);
nand U44842 (N_44842,N_44639,N_44633);
and U44843 (N_44843,N_44578,N_44561);
nor U44844 (N_44844,N_44554,N_44691);
nor U44845 (N_44845,N_44670,N_44650);
or U44846 (N_44846,N_44709,N_44669);
nand U44847 (N_44847,N_44567,N_44520);
and U44848 (N_44848,N_44555,N_44655);
and U44849 (N_44849,N_44698,N_44563);
xnor U44850 (N_44850,N_44645,N_44726);
xnor U44851 (N_44851,N_44531,N_44676);
nor U44852 (N_44852,N_44620,N_44702);
nand U44853 (N_44853,N_44599,N_44629);
nor U44854 (N_44854,N_44606,N_44741);
or U44855 (N_44855,N_44651,N_44527);
nor U44856 (N_44856,N_44569,N_44603);
xnor U44857 (N_44857,N_44568,N_44551);
or U44858 (N_44858,N_44612,N_44707);
nor U44859 (N_44859,N_44581,N_44694);
xnor U44860 (N_44860,N_44539,N_44533);
and U44861 (N_44861,N_44738,N_44600);
nand U44862 (N_44862,N_44689,N_44579);
or U44863 (N_44863,N_44587,N_44626);
nand U44864 (N_44864,N_44700,N_44546);
or U44865 (N_44865,N_44559,N_44514);
and U44866 (N_44866,N_44665,N_44577);
nor U44867 (N_44867,N_44557,N_44740);
nor U44868 (N_44868,N_44664,N_44690);
nor U44869 (N_44869,N_44663,N_44552);
and U44870 (N_44870,N_44687,N_44504);
and U44871 (N_44871,N_44721,N_44634);
and U44872 (N_44872,N_44518,N_44583);
xor U44873 (N_44873,N_44695,N_44597);
nand U44874 (N_44874,N_44594,N_44584);
nand U44875 (N_44875,N_44647,N_44710);
nor U44876 (N_44876,N_44511,N_44543);
nand U44877 (N_44877,N_44605,N_44607);
or U44878 (N_44878,N_44589,N_44514);
or U44879 (N_44879,N_44501,N_44576);
or U44880 (N_44880,N_44600,N_44661);
or U44881 (N_44881,N_44729,N_44684);
or U44882 (N_44882,N_44503,N_44621);
xor U44883 (N_44883,N_44571,N_44523);
and U44884 (N_44884,N_44718,N_44609);
xor U44885 (N_44885,N_44614,N_44603);
nand U44886 (N_44886,N_44509,N_44515);
nand U44887 (N_44887,N_44600,N_44613);
xnor U44888 (N_44888,N_44738,N_44667);
nor U44889 (N_44889,N_44586,N_44730);
and U44890 (N_44890,N_44577,N_44534);
and U44891 (N_44891,N_44638,N_44739);
or U44892 (N_44892,N_44661,N_44694);
nand U44893 (N_44893,N_44605,N_44529);
xor U44894 (N_44894,N_44679,N_44694);
nand U44895 (N_44895,N_44661,N_44604);
xnor U44896 (N_44896,N_44522,N_44545);
and U44897 (N_44897,N_44675,N_44611);
xnor U44898 (N_44898,N_44531,N_44596);
xor U44899 (N_44899,N_44599,N_44740);
nand U44900 (N_44900,N_44695,N_44696);
nor U44901 (N_44901,N_44665,N_44707);
nor U44902 (N_44902,N_44666,N_44533);
or U44903 (N_44903,N_44726,N_44521);
or U44904 (N_44904,N_44592,N_44562);
or U44905 (N_44905,N_44635,N_44680);
xor U44906 (N_44906,N_44649,N_44602);
nor U44907 (N_44907,N_44628,N_44528);
nand U44908 (N_44908,N_44598,N_44745);
nor U44909 (N_44909,N_44537,N_44686);
nor U44910 (N_44910,N_44665,N_44746);
or U44911 (N_44911,N_44571,N_44703);
nand U44912 (N_44912,N_44516,N_44626);
nand U44913 (N_44913,N_44690,N_44589);
or U44914 (N_44914,N_44595,N_44528);
or U44915 (N_44915,N_44722,N_44577);
nor U44916 (N_44916,N_44638,N_44543);
and U44917 (N_44917,N_44574,N_44593);
xor U44918 (N_44918,N_44708,N_44656);
xnor U44919 (N_44919,N_44570,N_44553);
xor U44920 (N_44920,N_44668,N_44522);
nand U44921 (N_44921,N_44629,N_44643);
and U44922 (N_44922,N_44593,N_44689);
or U44923 (N_44923,N_44691,N_44709);
xor U44924 (N_44924,N_44556,N_44686);
and U44925 (N_44925,N_44581,N_44678);
xor U44926 (N_44926,N_44556,N_44731);
nor U44927 (N_44927,N_44563,N_44539);
and U44928 (N_44928,N_44563,N_44676);
nor U44929 (N_44929,N_44668,N_44735);
and U44930 (N_44930,N_44526,N_44711);
or U44931 (N_44931,N_44713,N_44648);
or U44932 (N_44932,N_44573,N_44694);
xnor U44933 (N_44933,N_44525,N_44733);
xor U44934 (N_44934,N_44640,N_44715);
or U44935 (N_44935,N_44572,N_44717);
and U44936 (N_44936,N_44562,N_44746);
nor U44937 (N_44937,N_44660,N_44562);
and U44938 (N_44938,N_44595,N_44681);
xnor U44939 (N_44939,N_44740,N_44683);
or U44940 (N_44940,N_44710,N_44722);
nor U44941 (N_44941,N_44631,N_44608);
xor U44942 (N_44942,N_44595,N_44698);
nand U44943 (N_44943,N_44597,N_44642);
nand U44944 (N_44944,N_44623,N_44636);
nor U44945 (N_44945,N_44665,N_44675);
xnor U44946 (N_44946,N_44638,N_44700);
and U44947 (N_44947,N_44508,N_44651);
nor U44948 (N_44948,N_44663,N_44507);
nand U44949 (N_44949,N_44724,N_44545);
or U44950 (N_44950,N_44650,N_44599);
or U44951 (N_44951,N_44559,N_44645);
or U44952 (N_44952,N_44503,N_44595);
nor U44953 (N_44953,N_44650,N_44672);
or U44954 (N_44954,N_44534,N_44579);
nor U44955 (N_44955,N_44663,N_44642);
nor U44956 (N_44956,N_44683,N_44602);
and U44957 (N_44957,N_44650,N_44723);
or U44958 (N_44958,N_44541,N_44703);
xor U44959 (N_44959,N_44629,N_44546);
and U44960 (N_44960,N_44556,N_44636);
and U44961 (N_44961,N_44653,N_44694);
and U44962 (N_44962,N_44707,N_44577);
xor U44963 (N_44963,N_44657,N_44652);
or U44964 (N_44964,N_44513,N_44535);
and U44965 (N_44965,N_44704,N_44509);
nor U44966 (N_44966,N_44616,N_44732);
or U44967 (N_44967,N_44729,N_44504);
and U44968 (N_44968,N_44584,N_44531);
nand U44969 (N_44969,N_44621,N_44530);
nor U44970 (N_44970,N_44564,N_44588);
nand U44971 (N_44971,N_44676,N_44547);
xnor U44972 (N_44972,N_44730,N_44724);
and U44973 (N_44973,N_44717,N_44738);
nor U44974 (N_44974,N_44526,N_44713);
nand U44975 (N_44975,N_44524,N_44602);
nand U44976 (N_44976,N_44659,N_44726);
nor U44977 (N_44977,N_44723,N_44523);
or U44978 (N_44978,N_44748,N_44649);
or U44979 (N_44979,N_44515,N_44584);
or U44980 (N_44980,N_44645,N_44695);
nor U44981 (N_44981,N_44554,N_44740);
nor U44982 (N_44982,N_44657,N_44532);
xnor U44983 (N_44983,N_44587,N_44701);
or U44984 (N_44984,N_44528,N_44700);
nand U44985 (N_44985,N_44726,N_44564);
and U44986 (N_44986,N_44624,N_44518);
xor U44987 (N_44987,N_44531,N_44551);
or U44988 (N_44988,N_44523,N_44632);
or U44989 (N_44989,N_44526,N_44580);
or U44990 (N_44990,N_44608,N_44713);
xor U44991 (N_44991,N_44698,N_44745);
or U44992 (N_44992,N_44724,N_44664);
and U44993 (N_44993,N_44575,N_44718);
and U44994 (N_44994,N_44680,N_44528);
nand U44995 (N_44995,N_44641,N_44636);
and U44996 (N_44996,N_44741,N_44597);
xnor U44997 (N_44997,N_44733,N_44678);
nor U44998 (N_44998,N_44692,N_44632);
xnor U44999 (N_44999,N_44659,N_44500);
nor U45000 (N_45000,N_44960,N_44766);
and U45001 (N_45001,N_44968,N_44793);
xnor U45002 (N_45002,N_44771,N_44761);
and U45003 (N_45003,N_44873,N_44966);
xor U45004 (N_45004,N_44946,N_44949);
nor U45005 (N_45005,N_44980,N_44767);
or U45006 (N_45006,N_44947,N_44986);
or U45007 (N_45007,N_44774,N_44833);
xor U45008 (N_45008,N_44804,N_44851);
and U45009 (N_45009,N_44842,N_44890);
nor U45010 (N_45010,N_44918,N_44958);
nor U45011 (N_45011,N_44930,N_44756);
nand U45012 (N_45012,N_44956,N_44907);
nand U45013 (N_45013,N_44803,N_44805);
xnor U45014 (N_45014,N_44780,N_44938);
nand U45015 (N_45015,N_44885,N_44855);
xor U45016 (N_45016,N_44863,N_44777);
and U45017 (N_45017,N_44820,N_44818);
or U45018 (N_45018,N_44853,N_44982);
or U45019 (N_45019,N_44868,N_44898);
and U45020 (N_45020,N_44825,N_44891);
xor U45021 (N_45021,N_44915,N_44900);
nor U45022 (N_45022,N_44840,N_44936);
and U45023 (N_45023,N_44867,N_44995);
or U45024 (N_45024,N_44763,N_44954);
or U45025 (N_45025,N_44928,N_44810);
xnor U45026 (N_45026,N_44832,N_44990);
nand U45027 (N_45027,N_44878,N_44903);
and U45028 (N_45028,N_44939,N_44912);
nor U45029 (N_45029,N_44830,N_44758);
nand U45030 (N_45030,N_44797,N_44865);
xnor U45031 (N_45031,N_44970,N_44913);
xnor U45032 (N_45032,N_44933,N_44857);
and U45033 (N_45033,N_44893,N_44998);
or U45034 (N_45034,N_44925,N_44974);
and U45035 (N_45035,N_44942,N_44792);
and U45036 (N_45036,N_44874,N_44881);
nor U45037 (N_45037,N_44789,N_44940);
nand U45038 (N_45038,N_44862,N_44821);
nor U45039 (N_45039,N_44879,N_44997);
nand U45040 (N_45040,N_44914,N_44876);
xnor U45041 (N_45041,N_44852,N_44899);
nand U45042 (N_45042,N_44957,N_44790);
xnor U45043 (N_45043,N_44837,N_44843);
nand U45044 (N_45044,N_44993,N_44989);
xnor U45045 (N_45045,N_44769,N_44884);
and U45046 (N_45046,N_44943,N_44858);
nand U45047 (N_45047,N_44935,N_44757);
or U45048 (N_45048,N_44963,N_44779);
or U45049 (N_45049,N_44760,N_44854);
or U45050 (N_45050,N_44800,N_44969);
or U45051 (N_45051,N_44812,N_44984);
or U45052 (N_45052,N_44838,N_44870);
nand U45053 (N_45053,N_44831,N_44904);
and U45054 (N_45054,N_44847,N_44828);
and U45055 (N_45055,N_44994,N_44937);
xnor U45056 (N_45056,N_44752,N_44869);
nor U45057 (N_45057,N_44962,N_44866);
or U45058 (N_45058,N_44848,N_44905);
xnor U45059 (N_45059,N_44952,N_44791);
nand U45060 (N_45060,N_44944,N_44826);
and U45061 (N_45061,N_44861,N_44909);
or U45062 (N_45062,N_44950,N_44765);
nor U45063 (N_45063,N_44754,N_44886);
nand U45064 (N_45064,N_44911,N_44927);
or U45065 (N_45065,N_44973,N_44850);
or U45066 (N_45066,N_44948,N_44753);
and U45067 (N_45067,N_44750,N_44934);
or U45068 (N_45068,N_44896,N_44906);
and U45069 (N_45069,N_44809,N_44965);
and U45070 (N_45070,N_44815,N_44795);
xnor U45071 (N_45071,N_44964,N_44841);
nor U45072 (N_45072,N_44961,N_44931);
or U45073 (N_45073,N_44786,N_44953);
nand U45074 (N_45074,N_44834,N_44971);
nand U45075 (N_45075,N_44976,N_44979);
xor U45076 (N_45076,N_44856,N_44883);
and U45077 (N_45077,N_44864,N_44817);
nand U45078 (N_45078,N_44807,N_44875);
xor U45079 (N_45079,N_44887,N_44916);
or U45080 (N_45080,N_44992,N_44902);
or U45081 (N_45081,N_44827,N_44813);
or U45082 (N_45082,N_44770,N_44859);
or U45083 (N_45083,N_44996,N_44768);
xor U45084 (N_45084,N_44816,N_44806);
or U45085 (N_45085,N_44991,N_44849);
and U45086 (N_45086,N_44764,N_44917);
or U45087 (N_45087,N_44889,N_44778);
or U45088 (N_45088,N_44932,N_44784);
nor U45089 (N_45089,N_44823,N_44781);
xor U45090 (N_45090,N_44888,N_44796);
xnor U45091 (N_45091,N_44776,N_44999);
xor U45092 (N_45092,N_44895,N_44983);
nand U45093 (N_45093,N_44798,N_44773);
xor U45094 (N_45094,N_44908,N_44801);
and U45095 (N_45095,N_44819,N_44762);
and U45096 (N_45096,N_44787,N_44967);
or U45097 (N_45097,N_44985,N_44951);
or U45098 (N_45098,N_44802,N_44839);
and U45099 (N_45099,N_44959,N_44844);
or U45100 (N_45100,N_44783,N_44882);
nor U45101 (N_45101,N_44835,N_44782);
nor U45102 (N_45102,N_44845,N_44794);
or U45103 (N_45103,N_44788,N_44978);
or U45104 (N_45104,N_44901,N_44775);
nand U45105 (N_45105,N_44836,N_44846);
nand U45106 (N_45106,N_44799,N_44877);
xor U45107 (N_45107,N_44785,N_44759);
xnor U45108 (N_45108,N_44872,N_44972);
nor U45109 (N_45109,N_44977,N_44920);
nor U45110 (N_45110,N_44814,N_44880);
and U45111 (N_45111,N_44919,N_44860);
or U45112 (N_45112,N_44924,N_44987);
xor U45113 (N_45113,N_44922,N_44955);
nor U45114 (N_45114,N_44897,N_44811);
xor U45115 (N_45115,N_44929,N_44988);
or U45116 (N_45116,N_44824,N_44808);
nand U45117 (N_45117,N_44926,N_44945);
nor U45118 (N_45118,N_44921,N_44751);
nand U45119 (N_45119,N_44871,N_44941);
and U45120 (N_45120,N_44892,N_44981);
xor U45121 (N_45121,N_44910,N_44894);
and U45122 (N_45122,N_44755,N_44975);
nand U45123 (N_45123,N_44822,N_44772);
and U45124 (N_45124,N_44829,N_44923);
or U45125 (N_45125,N_44787,N_44813);
nand U45126 (N_45126,N_44985,N_44816);
or U45127 (N_45127,N_44752,N_44790);
or U45128 (N_45128,N_44890,N_44858);
or U45129 (N_45129,N_44918,N_44885);
nor U45130 (N_45130,N_44784,N_44860);
nor U45131 (N_45131,N_44900,N_44990);
nand U45132 (N_45132,N_44967,N_44932);
or U45133 (N_45133,N_44852,N_44955);
nor U45134 (N_45134,N_44772,N_44910);
nand U45135 (N_45135,N_44971,N_44811);
nand U45136 (N_45136,N_44857,N_44846);
nand U45137 (N_45137,N_44984,N_44883);
or U45138 (N_45138,N_44801,N_44837);
and U45139 (N_45139,N_44983,N_44783);
or U45140 (N_45140,N_44944,N_44899);
nand U45141 (N_45141,N_44753,N_44831);
xnor U45142 (N_45142,N_44892,N_44795);
or U45143 (N_45143,N_44853,N_44900);
nor U45144 (N_45144,N_44754,N_44955);
xor U45145 (N_45145,N_44975,N_44943);
or U45146 (N_45146,N_44752,N_44883);
xor U45147 (N_45147,N_44785,N_44767);
nand U45148 (N_45148,N_44814,N_44863);
nor U45149 (N_45149,N_44971,N_44900);
nor U45150 (N_45150,N_44770,N_44918);
or U45151 (N_45151,N_44941,N_44861);
nor U45152 (N_45152,N_44823,N_44907);
and U45153 (N_45153,N_44802,N_44906);
xnor U45154 (N_45154,N_44849,N_44777);
nand U45155 (N_45155,N_44797,N_44885);
and U45156 (N_45156,N_44766,N_44898);
or U45157 (N_45157,N_44802,N_44996);
or U45158 (N_45158,N_44970,N_44750);
or U45159 (N_45159,N_44820,N_44784);
and U45160 (N_45160,N_44977,N_44891);
xnor U45161 (N_45161,N_44924,N_44991);
xor U45162 (N_45162,N_44876,N_44893);
and U45163 (N_45163,N_44984,N_44822);
or U45164 (N_45164,N_44902,N_44873);
or U45165 (N_45165,N_44757,N_44862);
nor U45166 (N_45166,N_44801,N_44796);
and U45167 (N_45167,N_44770,N_44853);
or U45168 (N_45168,N_44996,N_44783);
xor U45169 (N_45169,N_44882,N_44951);
and U45170 (N_45170,N_44962,N_44827);
xnor U45171 (N_45171,N_44859,N_44994);
and U45172 (N_45172,N_44770,N_44940);
nand U45173 (N_45173,N_44750,N_44759);
and U45174 (N_45174,N_44818,N_44970);
nand U45175 (N_45175,N_44897,N_44885);
nor U45176 (N_45176,N_44883,N_44964);
xor U45177 (N_45177,N_44898,N_44758);
xor U45178 (N_45178,N_44968,N_44848);
nor U45179 (N_45179,N_44775,N_44839);
nor U45180 (N_45180,N_44904,N_44787);
or U45181 (N_45181,N_44972,N_44930);
nand U45182 (N_45182,N_44842,N_44968);
nand U45183 (N_45183,N_44751,N_44926);
or U45184 (N_45184,N_44793,N_44902);
nand U45185 (N_45185,N_44956,N_44766);
nor U45186 (N_45186,N_44984,N_44814);
nor U45187 (N_45187,N_44847,N_44999);
or U45188 (N_45188,N_44866,N_44892);
and U45189 (N_45189,N_44916,N_44820);
nor U45190 (N_45190,N_44836,N_44792);
and U45191 (N_45191,N_44904,N_44947);
or U45192 (N_45192,N_44953,N_44836);
xor U45193 (N_45193,N_44864,N_44917);
and U45194 (N_45194,N_44921,N_44998);
nand U45195 (N_45195,N_44766,N_44887);
or U45196 (N_45196,N_44967,N_44759);
xor U45197 (N_45197,N_44842,N_44780);
xnor U45198 (N_45198,N_44767,N_44779);
xor U45199 (N_45199,N_44755,N_44951);
nor U45200 (N_45200,N_44963,N_44786);
nor U45201 (N_45201,N_44998,N_44990);
xor U45202 (N_45202,N_44905,N_44755);
and U45203 (N_45203,N_44839,N_44754);
xnor U45204 (N_45204,N_44798,N_44878);
xnor U45205 (N_45205,N_44963,N_44875);
nand U45206 (N_45206,N_44970,N_44923);
or U45207 (N_45207,N_44909,N_44817);
nor U45208 (N_45208,N_44913,N_44888);
nand U45209 (N_45209,N_44931,N_44977);
or U45210 (N_45210,N_44813,N_44814);
nand U45211 (N_45211,N_44951,N_44922);
nand U45212 (N_45212,N_44995,N_44818);
or U45213 (N_45213,N_44904,N_44807);
or U45214 (N_45214,N_44936,N_44778);
or U45215 (N_45215,N_44919,N_44912);
or U45216 (N_45216,N_44867,N_44851);
and U45217 (N_45217,N_44933,N_44990);
nand U45218 (N_45218,N_44917,N_44992);
and U45219 (N_45219,N_44943,N_44863);
and U45220 (N_45220,N_44969,N_44772);
nor U45221 (N_45221,N_44793,N_44885);
or U45222 (N_45222,N_44797,N_44913);
or U45223 (N_45223,N_44876,N_44856);
xor U45224 (N_45224,N_44899,N_44980);
xor U45225 (N_45225,N_44885,N_44770);
xor U45226 (N_45226,N_44826,N_44951);
and U45227 (N_45227,N_44752,N_44936);
xor U45228 (N_45228,N_44890,N_44869);
nor U45229 (N_45229,N_44916,N_44902);
and U45230 (N_45230,N_44882,N_44869);
or U45231 (N_45231,N_44947,N_44834);
or U45232 (N_45232,N_44789,N_44945);
xor U45233 (N_45233,N_44875,N_44818);
nand U45234 (N_45234,N_44942,N_44794);
and U45235 (N_45235,N_44833,N_44864);
and U45236 (N_45236,N_44829,N_44881);
nand U45237 (N_45237,N_44884,N_44828);
xor U45238 (N_45238,N_44768,N_44884);
and U45239 (N_45239,N_44787,N_44968);
or U45240 (N_45240,N_44827,N_44829);
xnor U45241 (N_45241,N_44770,N_44780);
nor U45242 (N_45242,N_44926,N_44812);
nand U45243 (N_45243,N_44920,N_44814);
nand U45244 (N_45244,N_44910,N_44848);
and U45245 (N_45245,N_44963,N_44759);
nand U45246 (N_45246,N_44771,N_44946);
or U45247 (N_45247,N_44991,N_44750);
xnor U45248 (N_45248,N_44793,N_44847);
nor U45249 (N_45249,N_44908,N_44984);
or U45250 (N_45250,N_45101,N_45155);
nor U45251 (N_45251,N_45024,N_45233);
or U45252 (N_45252,N_45234,N_45049);
xnor U45253 (N_45253,N_45135,N_45042);
nor U45254 (N_45254,N_45227,N_45225);
nand U45255 (N_45255,N_45221,N_45050);
xnor U45256 (N_45256,N_45170,N_45109);
xnor U45257 (N_45257,N_45040,N_45048);
xnor U45258 (N_45258,N_45194,N_45028);
nand U45259 (N_45259,N_45191,N_45235);
xor U45260 (N_45260,N_45016,N_45237);
nand U45261 (N_45261,N_45153,N_45126);
or U45262 (N_45262,N_45168,N_45177);
and U45263 (N_45263,N_45120,N_45007);
nand U45264 (N_45264,N_45154,N_45211);
or U45265 (N_45265,N_45148,N_45215);
xor U45266 (N_45266,N_45118,N_45231);
nor U45267 (N_45267,N_45236,N_45151);
xnor U45268 (N_45268,N_45038,N_45008);
or U45269 (N_45269,N_45208,N_45037);
nand U45270 (N_45270,N_45137,N_45136);
nand U45271 (N_45271,N_45183,N_45093);
and U45272 (N_45272,N_45054,N_45242);
nand U45273 (N_45273,N_45067,N_45036);
xnor U45274 (N_45274,N_45196,N_45140);
nor U45275 (N_45275,N_45011,N_45133);
nand U45276 (N_45276,N_45088,N_45080);
nand U45277 (N_45277,N_45238,N_45083);
nor U45278 (N_45278,N_45057,N_45125);
or U45279 (N_45279,N_45230,N_45239);
nand U45280 (N_45280,N_45245,N_45045);
nand U45281 (N_45281,N_45090,N_45097);
or U45282 (N_45282,N_45022,N_45127);
nor U45283 (N_45283,N_45030,N_45199);
or U45284 (N_45284,N_45094,N_45033);
nand U45285 (N_45285,N_45174,N_45069);
nor U45286 (N_45286,N_45032,N_45071);
and U45287 (N_45287,N_45066,N_45213);
and U45288 (N_45288,N_45147,N_45072);
nor U45289 (N_45289,N_45190,N_45006);
xor U45290 (N_45290,N_45128,N_45124);
and U45291 (N_45291,N_45226,N_45058);
xor U45292 (N_45292,N_45070,N_45223);
xnor U45293 (N_45293,N_45089,N_45092);
and U45294 (N_45294,N_45001,N_45025);
and U45295 (N_45295,N_45130,N_45084);
xnor U45296 (N_45296,N_45074,N_45144);
and U45297 (N_45297,N_45000,N_45107);
xnor U45298 (N_45298,N_45059,N_45162);
xnor U45299 (N_45299,N_45210,N_45027);
and U45300 (N_45300,N_45053,N_45102);
and U45301 (N_45301,N_45014,N_45158);
nand U45302 (N_45302,N_45115,N_45246);
or U45303 (N_45303,N_45005,N_45171);
and U45304 (N_45304,N_45141,N_45184);
nor U45305 (N_45305,N_45222,N_45198);
nor U45306 (N_45306,N_45039,N_45220);
nor U45307 (N_45307,N_45013,N_45076);
nor U45308 (N_45308,N_45248,N_45023);
or U45309 (N_45309,N_45123,N_45240);
nor U45310 (N_45310,N_45161,N_45003);
nand U45311 (N_45311,N_45145,N_45085);
nand U45312 (N_45312,N_45002,N_45150);
xnor U45313 (N_45313,N_45219,N_45182);
or U45314 (N_45314,N_45202,N_45157);
nor U45315 (N_45315,N_45019,N_45209);
nand U45316 (N_45316,N_45010,N_45026);
nor U45317 (N_45317,N_45009,N_45114);
nand U45318 (N_45318,N_45173,N_45212);
xor U45319 (N_45319,N_45216,N_45186);
nor U45320 (N_45320,N_45160,N_45091);
nor U45321 (N_45321,N_45193,N_45041);
and U45322 (N_45322,N_45105,N_45146);
nor U45323 (N_45323,N_45138,N_45063);
or U45324 (N_45324,N_45121,N_45176);
nand U45325 (N_45325,N_45081,N_45247);
xnor U45326 (N_45326,N_45078,N_45132);
nor U45327 (N_45327,N_45178,N_45077);
nand U45328 (N_45328,N_45020,N_45205);
xnor U45329 (N_45329,N_45229,N_45104);
or U45330 (N_45330,N_45043,N_45111);
and U45331 (N_45331,N_45086,N_45131);
nor U45332 (N_45332,N_45163,N_45197);
xor U45333 (N_45333,N_45156,N_45015);
nor U45334 (N_45334,N_45228,N_45051);
or U45335 (N_45335,N_45029,N_45164);
xnor U45336 (N_45336,N_45249,N_45004);
or U45337 (N_45337,N_45224,N_45232);
or U45338 (N_45338,N_45187,N_45087);
or U45339 (N_45339,N_45201,N_45166);
nand U45340 (N_45340,N_45064,N_45047);
and U45341 (N_45341,N_45167,N_45044);
and U45342 (N_45342,N_45110,N_45034);
nor U45343 (N_45343,N_45099,N_45244);
and U45344 (N_45344,N_45181,N_45206);
xor U45345 (N_45345,N_45062,N_45103);
and U45346 (N_45346,N_45134,N_45195);
or U45347 (N_45347,N_45055,N_45204);
and U45348 (N_45348,N_45152,N_45189);
nor U45349 (N_45349,N_45073,N_45035);
nor U45350 (N_45350,N_45169,N_45119);
and U45351 (N_45351,N_45056,N_45192);
nor U45352 (N_45352,N_45052,N_45203);
nand U45353 (N_45353,N_45082,N_45112);
xor U45354 (N_45354,N_45061,N_45165);
and U45355 (N_45355,N_45217,N_45200);
or U45356 (N_45356,N_45241,N_45108);
or U45357 (N_45357,N_45117,N_45185);
and U45358 (N_45358,N_45243,N_45031);
or U45359 (N_45359,N_45106,N_45175);
nor U45360 (N_45360,N_45018,N_45095);
nand U45361 (N_45361,N_45098,N_45113);
nand U45362 (N_45362,N_45075,N_45149);
or U45363 (N_45363,N_45180,N_45060);
nor U45364 (N_45364,N_45143,N_45046);
or U45365 (N_45365,N_45207,N_45116);
nand U45366 (N_45366,N_45068,N_45096);
xor U45367 (N_45367,N_45021,N_45172);
nand U45368 (N_45368,N_45179,N_45139);
and U45369 (N_45369,N_45129,N_45214);
or U45370 (N_45370,N_45017,N_45065);
nand U45371 (N_45371,N_45012,N_45218);
xor U45372 (N_45372,N_45079,N_45142);
nor U45373 (N_45373,N_45188,N_45122);
xnor U45374 (N_45374,N_45100,N_45159);
nor U45375 (N_45375,N_45005,N_45111);
and U45376 (N_45376,N_45032,N_45161);
xnor U45377 (N_45377,N_45043,N_45115);
nand U45378 (N_45378,N_45246,N_45102);
nand U45379 (N_45379,N_45248,N_45091);
xnor U45380 (N_45380,N_45048,N_45078);
xnor U45381 (N_45381,N_45220,N_45221);
or U45382 (N_45382,N_45227,N_45088);
or U45383 (N_45383,N_45138,N_45176);
xor U45384 (N_45384,N_45102,N_45177);
or U45385 (N_45385,N_45050,N_45016);
or U45386 (N_45386,N_45220,N_45235);
xnor U45387 (N_45387,N_45061,N_45065);
nand U45388 (N_45388,N_45069,N_45207);
nor U45389 (N_45389,N_45154,N_45021);
and U45390 (N_45390,N_45098,N_45009);
or U45391 (N_45391,N_45188,N_45183);
xor U45392 (N_45392,N_45244,N_45064);
and U45393 (N_45393,N_45103,N_45160);
nor U45394 (N_45394,N_45188,N_45044);
nor U45395 (N_45395,N_45047,N_45155);
and U45396 (N_45396,N_45120,N_45239);
or U45397 (N_45397,N_45198,N_45157);
nor U45398 (N_45398,N_45030,N_45232);
or U45399 (N_45399,N_45180,N_45069);
nor U45400 (N_45400,N_45123,N_45170);
and U45401 (N_45401,N_45121,N_45040);
nand U45402 (N_45402,N_45247,N_45168);
and U45403 (N_45403,N_45054,N_45018);
nand U45404 (N_45404,N_45183,N_45117);
nor U45405 (N_45405,N_45132,N_45158);
and U45406 (N_45406,N_45227,N_45137);
or U45407 (N_45407,N_45241,N_45245);
nor U45408 (N_45408,N_45004,N_45240);
xor U45409 (N_45409,N_45191,N_45150);
xnor U45410 (N_45410,N_45127,N_45244);
or U45411 (N_45411,N_45045,N_45234);
or U45412 (N_45412,N_45189,N_45080);
xor U45413 (N_45413,N_45128,N_45146);
nand U45414 (N_45414,N_45104,N_45124);
and U45415 (N_45415,N_45017,N_45169);
nand U45416 (N_45416,N_45196,N_45199);
or U45417 (N_45417,N_45062,N_45064);
nor U45418 (N_45418,N_45192,N_45030);
nor U45419 (N_45419,N_45082,N_45057);
and U45420 (N_45420,N_45103,N_45204);
nand U45421 (N_45421,N_45134,N_45219);
nand U45422 (N_45422,N_45139,N_45239);
or U45423 (N_45423,N_45120,N_45029);
and U45424 (N_45424,N_45033,N_45081);
and U45425 (N_45425,N_45158,N_45186);
or U45426 (N_45426,N_45219,N_45112);
nor U45427 (N_45427,N_45027,N_45058);
or U45428 (N_45428,N_45021,N_45217);
nor U45429 (N_45429,N_45110,N_45228);
nand U45430 (N_45430,N_45100,N_45235);
nor U45431 (N_45431,N_45201,N_45115);
nand U45432 (N_45432,N_45226,N_45057);
or U45433 (N_45433,N_45023,N_45077);
nor U45434 (N_45434,N_45153,N_45079);
xor U45435 (N_45435,N_45016,N_45176);
nor U45436 (N_45436,N_45060,N_45118);
nor U45437 (N_45437,N_45042,N_45113);
nor U45438 (N_45438,N_45232,N_45047);
nor U45439 (N_45439,N_45201,N_45151);
nor U45440 (N_45440,N_45015,N_45231);
nor U45441 (N_45441,N_45099,N_45124);
and U45442 (N_45442,N_45031,N_45220);
nand U45443 (N_45443,N_45149,N_45207);
or U45444 (N_45444,N_45130,N_45164);
or U45445 (N_45445,N_45035,N_45083);
nand U45446 (N_45446,N_45097,N_45197);
xor U45447 (N_45447,N_45095,N_45092);
and U45448 (N_45448,N_45178,N_45112);
xnor U45449 (N_45449,N_45070,N_45100);
nand U45450 (N_45450,N_45238,N_45033);
and U45451 (N_45451,N_45104,N_45151);
or U45452 (N_45452,N_45202,N_45249);
or U45453 (N_45453,N_45247,N_45117);
and U45454 (N_45454,N_45246,N_45016);
and U45455 (N_45455,N_45110,N_45002);
xor U45456 (N_45456,N_45072,N_45103);
nand U45457 (N_45457,N_45105,N_45119);
nand U45458 (N_45458,N_45231,N_45216);
nand U45459 (N_45459,N_45083,N_45220);
nor U45460 (N_45460,N_45199,N_45041);
or U45461 (N_45461,N_45061,N_45041);
or U45462 (N_45462,N_45112,N_45003);
nand U45463 (N_45463,N_45225,N_45103);
and U45464 (N_45464,N_45163,N_45104);
and U45465 (N_45465,N_45125,N_45097);
nand U45466 (N_45466,N_45092,N_45038);
and U45467 (N_45467,N_45222,N_45212);
nand U45468 (N_45468,N_45048,N_45012);
and U45469 (N_45469,N_45054,N_45158);
or U45470 (N_45470,N_45074,N_45190);
xor U45471 (N_45471,N_45053,N_45069);
and U45472 (N_45472,N_45175,N_45228);
or U45473 (N_45473,N_45030,N_45126);
xnor U45474 (N_45474,N_45078,N_45184);
or U45475 (N_45475,N_45036,N_45110);
or U45476 (N_45476,N_45033,N_45154);
or U45477 (N_45477,N_45214,N_45072);
nor U45478 (N_45478,N_45182,N_45194);
and U45479 (N_45479,N_45153,N_45021);
xor U45480 (N_45480,N_45065,N_45220);
xnor U45481 (N_45481,N_45111,N_45023);
xnor U45482 (N_45482,N_45124,N_45002);
nor U45483 (N_45483,N_45161,N_45128);
or U45484 (N_45484,N_45232,N_45037);
or U45485 (N_45485,N_45081,N_45108);
nor U45486 (N_45486,N_45011,N_45015);
xnor U45487 (N_45487,N_45177,N_45022);
nand U45488 (N_45488,N_45078,N_45101);
and U45489 (N_45489,N_45124,N_45027);
and U45490 (N_45490,N_45102,N_45196);
xnor U45491 (N_45491,N_45035,N_45090);
or U45492 (N_45492,N_45144,N_45158);
nor U45493 (N_45493,N_45067,N_45136);
nand U45494 (N_45494,N_45227,N_45079);
nor U45495 (N_45495,N_45158,N_45234);
and U45496 (N_45496,N_45030,N_45035);
or U45497 (N_45497,N_45185,N_45164);
nand U45498 (N_45498,N_45063,N_45004);
nand U45499 (N_45499,N_45026,N_45052);
nand U45500 (N_45500,N_45355,N_45344);
nand U45501 (N_45501,N_45378,N_45380);
nand U45502 (N_45502,N_45415,N_45438);
xor U45503 (N_45503,N_45354,N_45454);
nor U45504 (N_45504,N_45467,N_45381);
and U45505 (N_45505,N_45262,N_45338);
nand U45506 (N_45506,N_45429,N_45409);
and U45507 (N_45507,N_45495,N_45283);
or U45508 (N_45508,N_45319,N_45316);
xnor U45509 (N_45509,N_45308,N_45386);
nand U45510 (N_45510,N_45395,N_45443);
xnor U45511 (N_45511,N_45497,N_45309);
xor U45512 (N_45512,N_45461,N_45496);
xnor U45513 (N_45513,N_45321,N_45337);
or U45514 (N_45514,N_45423,N_45484);
xnor U45515 (N_45515,N_45404,N_45469);
and U45516 (N_45516,N_45250,N_45372);
nand U45517 (N_45517,N_45313,N_45434);
nor U45518 (N_45518,N_45435,N_45340);
xnor U45519 (N_45519,N_45458,N_45470);
and U45520 (N_45520,N_45418,N_45272);
xor U45521 (N_45521,N_45267,N_45274);
or U45522 (N_45522,N_45329,N_45492);
nand U45523 (N_45523,N_45396,N_45485);
xnor U45524 (N_45524,N_45424,N_45252);
or U45525 (N_45525,N_45268,N_45482);
xnor U45526 (N_45526,N_45433,N_45315);
nor U45527 (N_45527,N_45260,N_45298);
nor U45528 (N_45528,N_45493,N_45285);
and U45529 (N_45529,N_45310,N_45306);
and U45530 (N_45530,N_45450,N_45343);
and U45531 (N_45531,N_45400,N_45393);
nor U45532 (N_45532,N_45322,N_45473);
nor U45533 (N_45533,N_45451,N_45312);
and U45534 (N_45534,N_45453,N_45323);
or U45535 (N_45535,N_45420,N_45333);
or U45536 (N_45536,N_45363,N_45463);
xor U45537 (N_45537,N_45281,N_45431);
nor U45538 (N_45538,N_45276,N_45320);
nand U45539 (N_45539,N_45425,N_45266);
xor U45540 (N_45540,N_45279,N_45362);
and U45541 (N_45541,N_45401,N_45376);
or U45542 (N_45542,N_45264,N_45271);
or U45543 (N_45543,N_45472,N_45325);
or U45544 (N_45544,N_45368,N_45498);
nand U45545 (N_45545,N_45375,N_45477);
and U45546 (N_45546,N_45374,N_45334);
xor U45547 (N_45547,N_45416,N_45361);
or U45548 (N_45548,N_45476,N_45326);
nand U45549 (N_45549,N_45455,N_45366);
nor U45550 (N_45550,N_45304,N_45452);
nand U45551 (N_45551,N_45410,N_45307);
nand U45552 (N_45552,N_45373,N_45462);
nor U45553 (N_45553,N_45351,N_45341);
nor U45554 (N_45554,N_45254,N_45448);
nor U45555 (N_45555,N_45287,N_45446);
xor U45556 (N_45556,N_45350,N_45311);
and U45557 (N_45557,N_45426,N_45499);
or U45558 (N_45558,N_45392,N_45474);
nor U45559 (N_45559,N_45399,N_45494);
and U45560 (N_45560,N_45295,N_45336);
nor U45561 (N_45561,N_45391,N_45457);
nor U45562 (N_45562,N_45468,N_45317);
xnor U45563 (N_45563,N_45471,N_45352);
and U45564 (N_45564,N_45327,N_45456);
and U45565 (N_45565,N_45278,N_45365);
or U45566 (N_45566,N_45277,N_45465);
xor U45567 (N_45567,N_45275,N_45379);
nand U45568 (N_45568,N_45360,N_45488);
xor U45569 (N_45569,N_45258,N_45293);
and U45570 (N_45570,N_45367,N_45257);
and U45571 (N_45571,N_45357,N_45412);
nor U45572 (N_45572,N_45270,N_45314);
nor U45573 (N_45573,N_45407,N_45292);
nand U45574 (N_45574,N_45263,N_45251);
nor U45575 (N_45575,N_45486,N_45324);
xor U45576 (N_45576,N_45436,N_45331);
nor U45577 (N_45577,N_45347,N_45441);
nor U45578 (N_45578,N_45345,N_45405);
nor U45579 (N_45579,N_45300,N_45478);
or U45580 (N_45580,N_45358,N_45356);
nor U45581 (N_45581,N_45273,N_45377);
or U45582 (N_45582,N_45284,N_45294);
nand U45583 (N_45583,N_45387,N_45353);
or U45584 (N_45584,N_45346,N_45385);
nand U45585 (N_45585,N_45475,N_45390);
xnor U45586 (N_45586,N_45389,N_45259);
nand U45587 (N_45587,N_45437,N_45447);
or U45588 (N_45588,N_45466,N_45288);
or U45589 (N_45589,N_45349,N_45439);
xor U45590 (N_45590,N_45370,N_45442);
and U45591 (N_45591,N_45342,N_45369);
or U45592 (N_45592,N_45280,N_45318);
or U45593 (N_45593,N_45428,N_45296);
or U45594 (N_45594,N_45480,N_45291);
nand U45595 (N_45595,N_45297,N_45388);
nor U45596 (N_45596,N_45282,N_45332);
xnor U45597 (N_45597,N_45427,N_45299);
xnor U45598 (N_45598,N_45491,N_45255);
nor U45599 (N_45599,N_45359,N_45490);
xor U45600 (N_45600,N_45440,N_45397);
and U45601 (N_45601,N_45411,N_45286);
and U45602 (N_45602,N_45335,N_45289);
nand U45603 (N_45603,N_45348,N_45464);
nor U45604 (N_45604,N_45290,N_45445);
xor U45605 (N_45605,N_45269,N_45487);
xor U45606 (N_45606,N_45417,N_45394);
nand U45607 (N_45607,N_45489,N_45305);
and U45608 (N_45608,N_45384,N_45414);
nand U45609 (N_45609,N_45256,N_45339);
or U45610 (N_45610,N_45444,N_45383);
xnor U45611 (N_45611,N_45432,N_45413);
xor U45612 (N_45612,N_45382,N_45330);
xnor U45613 (N_45613,N_45265,N_45302);
nand U45614 (N_45614,N_45364,N_45419);
nand U45615 (N_45615,N_45421,N_45303);
or U45616 (N_45616,N_45403,N_45301);
nand U45617 (N_45617,N_45430,N_45253);
and U45618 (N_45618,N_45398,N_45261);
and U45619 (N_45619,N_45479,N_45483);
and U45620 (N_45620,N_45459,N_45328);
nand U45621 (N_45621,N_45371,N_45408);
or U45622 (N_45622,N_45406,N_45449);
xnor U45623 (N_45623,N_45481,N_45402);
nor U45624 (N_45624,N_45422,N_45460);
and U45625 (N_45625,N_45281,N_45306);
xnor U45626 (N_45626,N_45496,N_45270);
or U45627 (N_45627,N_45401,N_45402);
nand U45628 (N_45628,N_45498,N_45316);
and U45629 (N_45629,N_45438,N_45345);
xnor U45630 (N_45630,N_45270,N_45266);
nor U45631 (N_45631,N_45359,N_45398);
xnor U45632 (N_45632,N_45353,N_45412);
nor U45633 (N_45633,N_45341,N_45339);
and U45634 (N_45634,N_45417,N_45266);
xnor U45635 (N_45635,N_45410,N_45282);
xor U45636 (N_45636,N_45336,N_45454);
nor U45637 (N_45637,N_45402,N_45459);
nand U45638 (N_45638,N_45496,N_45381);
nand U45639 (N_45639,N_45414,N_45342);
nand U45640 (N_45640,N_45427,N_45311);
and U45641 (N_45641,N_45395,N_45348);
nand U45642 (N_45642,N_45396,N_45496);
or U45643 (N_45643,N_45306,N_45348);
or U45644 (N_45644,N_45271,N_45392);
xnor U45645 (N_45645,N_45283,N_45278);
and U45646 (N_45646,N_45472,N_45273);
and U45647 (N_45647,N_45315,N_45289);
and U45648 (N_45648,N_45485,N_45284);
and U45649 (N_45649,N_45318,N_45391);
nor U45650 (N_45650,N_45465,N_45431);
nand U45651 (N_45651,N_45269,N_45312);
or U45652 (N_45652,N_45347,N_45339);
nand U45653 (N_45653,N_45259,N_45360);
or U45654 (N_45654,N_45394,N_45393);
xnor U45655 (N_45655,N_45252,N_45300);
nor U45656 (N_45656,N_45447,N_45305);
nor U45657 (N_45657,N_45261,N_45397);
nor U45658 (N_45658,N_45424,N_45265);
or U45659 (N_45659,N_45499,N_45260);
nor U45660 (N_45660,N_45298,N_45366);
xnor U45661 (N_45661,N_45496,N_45417);
or U45662 (N_45662,N_45347,N_45269);
and U45663 (N_45663,N_45357,N_45445);
nand U45664 (N_45664,N_45482,N_45467);
or U45665 (N_45665,N_45264,N_45316);
nor U45666 (N_45666,N_45263,N_45336);
or U45667 (N_45667,N_45329,N_45341);
xor U45668 (N_45668,N_45365,N_45262);
nand U45669 (N_45669,N_45307,N_45421);
or U45670 (N_45670,N_45291,N_45372);
nand U45671 (N_45671,N_45430,N_45462);
or U45672 (N_45672,N_45496,N_45283);
xnor U45673 (N_45673,N_45429,N_45320);
and U45674 (N_45674,N_45339,N_45328);
and U45675 (N_45675,N_45291,N_45350);
and U45676 (N_45676,N_45375,N_45254);
nand U45677 (N_45677,N_45408,N_45309);
nor U45678 (N_45678,N_45357,N_45428);
xnor U45679 (N_45679,N_45413,N_45386);
or U45680 (N_45680,N_45271,N_45254);
nor U45681 (N_45681,N_45497,N_45387);
or U45682 (N_45682,N_45407,N_45390);
xor U45683 (N_45683,N_45306,N_45340);
or U45684 (N_45684,N_45312,N_45301);
nor U45685 (N_45685,N_45465,N_45495);
nor U45686 (N_45686,N_45389,N_45381);
nor U45687 (N_45687,N_45381,N_45400);
and U45688 (N_45688,N_45289,N_45344);
and U45689 (N_45689,N_45267,N_45409);
nor U45690 (N_45690,N_45452,N_45293);
or U45691 (N_45691,N_45446,N_45406);
nor U45692 (N_45692,N_45269,N_45459);
xor U45693 (N_45693,N_45307,N_45460);
nor U45694 (N_45694,N_45481,N_45397);
xor U45695 (N_45695,N_45364,N_45294);
nand U45696 (N_45696,N_45306,N_45382);
xor U45697 (N_45697,N_45265,N_45489);
and U45698 (N_45698,N_45394,N_45346);
or U45699 (N_45699,N_45338,N_45344);
nand U45700 (N_45700,N_45256,N_45467);
and U45701 (N_45701,N_45433,N_45451);
or U45702 (N_45702,N_45298,N_45365);
nor U45703 (N_45703,N_45302,N_45492);
xor U45704 (N_45704,N_45254,N_45425);
nand U45705 (N_45705,N_45285,N_45365);
or U45706 (N_45706,N_45380,N_45286);
nand U45707 (N_45707,N_45433,N_45420);
or U45708 (N_45708,N_45444,N_45287);
and U45709 (N_45709,N_45371,N_45268);
nor U45710 (N_45710,N_45419,N_45380);
xor U45711 (N_45711,N_45282,N_45446);
nand U45712 (N_45712,N_45351,N_45278);
xnor U45713 (N_45713,N_45430,N_45353);
or U45714 (N_45714,N_45346,N_45494);
nand U45715 (N_45715,N_45335,N_45443);
or U45716 (N_45716,N_45459,N_45418);
and U45717 (N_45717,N_45303,N_45442);
and U45718 (N_45718,N_45283,N_45402);
xor U45719 (N_45719,N_45319,N_45367);
nor U45720 (N_45720,N_45437,N_45320);
nor U45721 (N_45721,N_45470,N_45372);
nor U45722 (N_45722,N_45445,N_45480);
and U45723 (N_45723,N_45342,N_45257);
xnor U45724 (N_45724,N_45359,N_45280);
xor U45725 (N_45725,N_45299,N_45382);
and U45726 (N_45726,N_45299,N_45339);
xor U45727 (N_45727,N_45280,N_45373);
and U45728 (N_45728,N_45445,N_45354);
xnor U45729 (N_45729,N_45357,N_45323);
or U45730 (N_45730,N_45417,N_45407);
nand U45731 (N_45731,N_45462,N_45272);
nand U45732 (N_45732,N_45318,N_45381);
nor U45733 (N_45733,N_45322,N_45454);
nor U45734 (N_45734,N_45318,N_45373);
and U45735 (N_45735,N_45448,N_45291);
xnor U45736 (N_45736,N_45325,N_45301);
and U45737 (N_45737,N_45384,N_45335);
nand U45738 (N_45738,N_45250,N_45257);
or U45739 (N_45739,N_45295,N_45312);
nand U45740 (N_45740,N_45488,N_45480);
or U45741 (N_45741,N_45402,N_45369);
nand U45742 (N_45742,N_45273,N_45255);
and U45743 (N_45743,N_45444,N_45284);
nand U45744 (N_45744,N_45329,N_45306);
or U45745 (N_45745,N_45366,N_45267);
and U45746 (N_45746,N_45363,N_45409);
nor U45747 (N_45747,N_45360,N_45485);
and U45748 (N_45748,N_45293,N_45263);
xor U45749 (N_45749,N_45358,N_45349);
nor U45750 (N_45750,N_45736,N_45669);
nor U45751 (N_45751,N_45711,N_45663);
nand U45752 (N_45752,N_45512,N_45652);
xnor U45753 (N_45753,N_45680,N_45577);
or U45754 (N_45754,N_45614,N_45662);
and U45755 (N_45755,N_45588,N_45698);
nor U45756 (N_45756,N_45547,N_45697);
or U45757 (N_45757,N_45673,N_45715);
nand U45758 (N_45758,N_45548,N_45608);
and U45759 (N_45759,N_45668,N_45705);
nand U45760 (N_45760,N_45585,N_45621);
and U45761 (N_45761,N_45619,N_45545);
nor U45762 (N_45762,N_45661,N_45598);
nand U45763 (N_45763,N_45583,N_45687);
or U45764 (N_45764,N_45591,N_45510);
nor U45765 (N_45765,N_45695,N_45513);
nand U45766 (N_45766,N_45678,N_45523);
and U45767 (N_45767,N_45683,N_45543);
nor U45768 (N_45768,N_45519,N_45601);
and U45769 (N_45769,N_45604,N_45534);
or U45770 (N_45770,N_45655,N_45639);
or U45771 (N_45771,N_45551,N_45657);
xnor U45772 (N_45772,N_45617,N_45546);
and U45773 (N_45773,N_45729,N_45738);
xor U45774 (N_45774,N_45539,N_45560);
xor U45775 (N_45775,N_45643,N_45740);
or U45776 (N_45776,N_45568,N_45647);
nand U45777 (N_45777,N_45508,N_45730);
or U45778 (N_45778,N_45709,N_45501);
nor U45779 (N_45779,N_45563,N_45593);
xnor U45780 (N_45780,N_45587,N_45739);
and U45781 (N_45781,N_45575,N_45618);
or U45782 (N_45782,N_45612,N_45620);
nand U45783 (N_45783,N_45693,N_45542);
xnor U45784 (N_45784,N_45670,N_45688);
or U45785 (N_45785,N_45700,N_45732);
nand U45786 (N_45786,N_45746,N_45712);
nor U45787 (N_45787,N_45727,N_45742);
nor U45788 (N_45788,N_45525,N_45672);
nor U45789 (N_45789,N_45656,N_45564);
xor U45790 (N_45790,N_45648,N_45566);
and U45791 (N_45791,N_45558,N_45611);
nand U45792 (N_45792,N_45685,N_45692);
nor U45793 (N_45793,N_45505,N_45616);
and U45794 (N_45794,N_45518,N_45701);
and U45795 (N_45795,N_45702,N_45671);
and U45796 (N_45796,N_45649,N_45703);
or U45797 (N_45797,N_45531,N_45667);
and U45798 (N_45798,N_45694,N_45615);
xor U45799 (N_45799,N_45626,N_45666);
nand U45800 (N_45800,N_45704,N_45520);
nor U45801 (N_45801,N_45550,N_45676);
nor U45802 (N_45802,N_45610,N_45691);
nor U45803 (N_45803,N_45743,N_45516);
nor U45804 (N_45804,N_45530,N_45607);
and U45805 (N_45805,N_45589,N_45748);
xor U45806 (N_45806,N_45600,N_45749);
xnor U45807 (N_45807,N_45674,N_45572);
nor U45808 (N_45808,N_45716,N_45719);
and U45809 (N_45809,N_45646,N_45664);
nor U45810 (N_45810,N_45713,N_45675);
xor U45811 (N_45811,N_45651,N_45557);
or U45812 (N_45812,N_45609,N_45707);
and U45813 (N_45813,N_45684,N_45689);
and U45814 (N_45814,N_45561,N_45517);
nor U45815 (N_45815,N_45638,N_45659);
and U45816 (N_45816,N_45570,N_45574);
and U45817 (N_45817,N_45696,N_45559);
xor U45818 (N_45818,N_45628,N_45722);
nor U45819 (N_45819,N_45708,N_45690);
nor U45820 (N_45820,N_45595,N_45580);
xnor U45821 (N_45821,N_45506,N_45650);
xnor U45822 (N_45822,N_45503,N_45735);
nand U45823 (N_45823,N_45532,N_45734);
nor U45824 (N_45824,N_45665,N_45509);
nor U45825 (N_45825,N_45654,N_45624);
and U45826 (N_45826,N_45747,N_45586);
xor U45827 (N_45827,N_45515,N_45502);
nor U45828 (N_45828,N_45511,N_45535);
or U45829 (N_45829,N_45699,N_45504);
or U45830 (N_45830,N_45605,N_45592);
xor U45831 (N_45831,N_45526,N_45625);
xor U45832 (N_45832,N_45541,N_45640);
xnor U45833 (N_45833,N_45725,N_45507);
xor U45834 (N_45834,N_45569,N_45636);
nor U45835 (N_45835,N_45645,N_45660);
nand U45836 (N_45836,N_45641,N_45629);
xnor U45837 (N_45837,N_45522,N_45644);
nand U45838 (N_45838,N_45528,N_45533);
nor U45839 (N_45839,N_45536,N_45552);
xor U45840 (N_45840,N_45737,N_45581);
nor U45841 (N_45841,N_45733,N_45642);
and U45842 (N_45842,N_45529,N_45579);
and U45843 (N_45843,N_45717,N_45627);
and U45844 (N_45844,N_45630,N_45631);
xnor U45845 (N_45845,N_45524,N_45623);
and U45846 (N_45846,N_45603,N_45632);
nand U45847 (N_45847,N_45635,N_45681);
or U45848 (N_45848,N_45744,N_45538);
or U45849 (N_45849,N_45527,N_45537);
nand U45850 (N_45850,N_45634,N_45555);
nand U45851 (N_45851,N_45554,N_45706);
xnor U45852 (N_45852,N_45726,N_45596);
and U45853 (N_45853,N_45584,N_45724);
nor U45854 (N_45854,N_45633,N_45599);
nand U45855 (N_45855,N_45567,N_45565);
nand U45856 (N_45856,N_45745,N_45576);
and U45857 (N_45857,N_45594,N_45553);
nand U45858 (N_45858,N_45514,N_45679);
xor U45859 (N_45859,N_45500,N_45582);
nor U45860 (N_45860,N_45544,N_45571);
nand U45861 (N_45861,N_45741,N_45613);
or U45862 (N_45862,N_45653,N_45714);
xnor U45863 (N_45863,N_45720,N_45578);
or U45864 (N_45864,N_45573,N_45540);
or U45865 (N_45865,N_45718,N_45590);
or U45866 (N_45866,N_45606,N_45556);
or U45867 (N_45867,N_45658,N_45562);
or U45868 (N_45868,N_45682,N_45728);
xnor U45869 (N_45869,N_45521,N_45723);
xor U45870 (N_45870,N_45731,N_45602);
nor U45871 (N_45871,N_45637,N_45597);
xnor U45872 (N_45872,N_45721,N_45622);
nor U45873 (N_45873,N_45677,N_45549);
nand U45874 (N_45874,N_45686,N_45710);
and U45875 (N_45875,N_45581,N_45509);
and U45876 (N_45876,N_45549,N_45535);
nand U45877 (N_45877,N_45737,N_45675);
or U45878 (N_45878,N_45652,N_45615);
nor U45879 (N_45879,N_45605,N_45675);
and U45880 (N_45880,N_45712,N_45671);
or U45881 (N_45881,N_45651,N_45730);
and U45882 (N_45882,N_45662,N_45739);
and U45883 (N_45883,N_45671,N_45689);
and U45884 (N_45884,N_45694,N_45605);
nand U45885 (N_45885,N_45504,N_45587);
nand U45886 (N_45886,N_45728,N_45696);
nor U45887 (N_45887,N_45515,N_45679);
and U45888 (N_45888,N_45585,N_45671);
nor U45889 (N_45889,N_45683,N_45605);
nor U45890 (N_45890,N_45701,N_45552);
nand U45891 (N_45891,N_45671,N_45641);
nand U45892 (N_45892,N_45518,N_45570);
xnor U45893 (N_45893,N_45617,N_45533);
and U45894 (N_45894,N_45735,N_45643);
and U45895 (N_45895,N_45635,N_45685);
and U45896 (N_45896,N_45536,N_45601);
or U45897 (N_45897,N_45500,N_45722);
or U45898 (N_45898,N_45650,N_45586);
xnor U45899 (N_45899,N_45595,N_45591);
nor U45900 (N_45900,N_45688,N_45641);
or U45901 (N_45901,N_45518,N_45616);
and U45902 (N_45902,N_45721,N_45597);
nor U45903 (N_45903,N_45722,N_45526);
and U45904 (N_45904,N_45560,N_45515);
or U45905 (N_45905,N_45685,N_45655);
and U45906 (N_45906,N_45537,N_45686);
and U45907 (N_45907,N_45693,N_45621);
or U45908 (N_45908,N_45575,N_45504);
nor U45909 (N_45909,N_45749,N_45726);
xnor U45910 (N_45910,N_45511,N_45521);
nor U45911 (N_45911,N_45592,N_45721);
xnor U45912 (N_45912,N_45716,N_45533);
nor U45913 (N_45913,N_45607,N_45553);
nor U45914 (N_45914,N_45731,N_45639);
and U45915 (N_45915,N_45730,N_45583);
or U45916 (N_45916,N_45617,N_45628);
xnor U45917 (N_45917,N_45599,N_45720);
nand U45918 (N_45918,N_45568,N_45559);
xor U45919 (N_45919,N_45550,N_45717);
or U45920 (N_45920,N_45727,N_45512);
nand U45921 (N_45921,N_45670,N_45573);
nand U45922 (N_45922,N_45516,N_45675);
and U45923 (N_45923,N_45543,N_45610);
xnor U45924 (N_45924,N_45725,N_45709);
or U45925 (N_45925,N_45622,N_45710);
and U45926 (N_45926,N_45692,N_45611);
or U45927 (N_45927,N_45738,N_45659);
nand U45928 (N_45928,N_45710,N_45581);
or U45929 (N_45929,N_45657,N_45625);
or U45930 (N_45930,N_45535,N_45512);
xor U45931 (N_45931,N_45696,N_45718);
xnor U45932 (N_45932,N_45542,N_45700);
and U45933 (N_45933,N_45568,N_45684);
nor U45934 (N_45934,N_45691,N_45671);
xor U45935 (N_45935,N_45526,N_45525);
or U45936 (N_45936,N_45548,N_45556);
nand U45937 (N_45937,N_45673,N_45660);
nand U45938 (N_45938,N_45504,N_45640);
and U45939 (N_45939,N_45655,N_45739);
xnor U45940 (N_45940,N_45513,N_45587);
xnor U45941 (N_45941,N_45586,N_45572);
xor U45942 (N_45942,N_45519,N_45565);
xnor U45943 (N_45943,N_45596,N_45534);
nor U45944 (N_45944,N_45652,N_45674);
or U45945 (N_45945,N_45539,N_45708);
nor U45946 (N_45946,N_45701,N_45665);
or U45947 (N_45947,N_45748,N_45503);
nand U45948 (N_45948,N_45609,N_45702);
nand U45949 (N_45949,N_45596,N_45629);
and U45950 (N_45950,N_45513,N_45606);
nor U45951 (N_45951,N_45534,N_45532);
nor U45952 (N_45952,N_45541,N_45568);
nand U45953 (N_45953,N_45530,N_45639);
nor U45954 (N_45954,N_45613,N_45668);
nand U45955 (N_45955,N_45595,N_45500);
nand U45956 (N_45956,N_45594,N_45664);
or U45957 (N_45957,N_45593,N_45722);
nor U45958 (N_45958,N_45595,N_45511);
nand U45959 (N_45959,N_45555,N_45729);
or U45960 (N_45960,N_45721,N_45639);
nor U45961 (N_45961,N_45574,N_45655);
or U45962 (N_45962,N_45587,N_45590);
nor U45963 (N_45963,N_45664,N_45732);
nor U45964 (N_45964,N_45728,N_45566);
nand U45965 (N_45965,N_45724,N_45534);
nor U45966 (N_45966,N_45706,N_45636);
or U45967 (N_45967,N_45600,N_45696);
xnor U45968 (N_45968,N_45671,N_45528);
nor U45969 (N_45969,N_45719,N_45607);
xor U45970 (N_45970,N_45616,N_45669);
and U45971 (N_45971,N_45657,N_45574);
or U45972 (N_45972,N_45558,N_45560);
nand U45973 (N_45973,N_45520,N_45749);
nor U45974 (N_45974,N_45532,N_45593);
nand U45975 (N_45975,N_45669,N_45510);
or U45976 (N_45976,N_45606,N_45575);
nand U45977 (N_45977,N_45714,N_45624);
nor U45978 (N_45978,N_45504,N_45706);
and U45979 (N_45979,N_45536,N_45560);
nand U45980 (N_45980,N_45528,N_45552);
nand U45981 (N_45981,N_45695,N_45586);
or U45982 (N_45982,N_45542,N_45574);
xor U45983 (N_45983,N_45690,N_45673);
xnor U45984 (N_45984,N_45726,N_45617);
and U45985 (N_45985,N_45538,N_45578);
and U45986 (N_45986,N_45704,N_45644);
or U45987 (N_45987,N_45622,N_45749);
and U45988 (N_45988,N_45600,N_45630);
and U45989 (N_45989,N_45501,N_45641);
and U45990 (N_45990,N_45673,N_45637);
and U45991 (N_45991,N_45585,N_45704);
nand U45992 (N_45992,N_45642,N_45589);
or U45993 (N_45993,N_45666,N_45683);
nand U45994 (N_45994,N_45603,N_45638);
or U45995 (N_45995,N_45569,N_45645);
xnor U45996 (N_45996,N_45597,N_45714);
nand U45997 (N_45997,N_45545,N_45634);
and U45998 (N_45998,N_45606,N_45677);
nor U45999 (N_45999,N_45612,N_45653);
xor U46000 (N_46000,N_45987,N_45994);
nand U46001 (N_46001,N_45916,N_45982);
or U46002 (N_46002,N_45860,N_45838);
and U46003 (N_46003,N_45938,N_45822);
and U46004 (N_46004,N_45990,N_45984);
and U46005 (N_46005,N_45887,N_45973);
or U46006 (N_46006,N_45773,N_45915);
and U46007 (N_46007,N_45955,N_45934);
and U46008 (N_46008,N_45926,N_45911);
or U46009 (N_46009,N_45872,N_45886);
nor U46010 (N_46010,N_45992,N_45841);
nor U46011 (N_46011,N_45948,N_45906);
or U46012 (N_46012,N_45802,N_45880);
or U46013 (N_46013,N_45929,N_45801);
nor U46014 (N_46014,N_45753,N_45898);
xor U46015 (N_46015,N_45965,N_45989);
and U46016 (N_46016,N_45780,N_45888);
and U46017 (N_46017,N_45851,N_45751);
nor U46018 (N_46018,N_45769,N_45980);
xor U46019 (N_46019,N_45787,N_45789);
and U46020 (N_46020,N_45956,N_45759);
and U46021 (N_46021,N_45823,N_45931);
nand U46022 (N_46022,N_45762,N_45899);
or U46023 (N_46023,N_45756,N_45968);
or U46024 (N_46024,N_45870,N_45917);
nor U46025 (N_46025,N_45991,N_45834);
or U46026 (N_46026,N_45806,N_45998);
and U46027 (N_46027,N_45889,N_45848);
xnor U46028 (N_46028,N_45814,N_45988);
xor U46029 (N_46029,N_45975,N_45912);
and U46030 (N_46030,N_45840,N_45797);
or U46031 (N_46031,N_45776,N_45824);
or U46032 (N_46032,N_45967,N_45809);
nor U46033 (N_46033,N_45947,N_45777);
xnor U46034 (N_46034,N_45845,N_45795);
xor U46035 (N_46035,N_45937,N_45862);
nor U46036 (N_46036,N_45864,N_45770);
or U46037 (N_46037,N_45974,N_45942);
nor U46038 (N_46038,N_45933,N_45859);
and U46039 (N_46039,N_45874,N_45794);
nor U46040 (N_46040,N_45995,N_45936);
nor U46041 (N_46041,N_45784,N_45952);
or U46042 (N_46042,N_45964,N_45861);
or U46043 (N_46043,N_45798,N_45771);
and U46044 (N_46044,N_45999,N_45878);
or U46045 (N_46045,N_45791,N_45792);
or U46046 (N_46046,N_45966,N_45796);
nor U46047 (N_46047,N_45951,N_45807);
nand U46048 (N_46048,N_45993,N_45953);
or U46049 (N_46049,N_45909,N_45954);
nor U46050 (N_46050,N_45818,N_45904);
nor U46051 (N_46051,N_45907,N_45812);
and U46052 (N_46052,N_45986,N_45891);
nor U46053 (N_46053,N_45856,N_45875);
and U46054 (N_46054,N_45981,N_45945);
and U46055 (N_46055,N_45785,N_45997);
or U46056 (N_46056,N_45808,N_45913);
xor U46057 (N_46057,N_45963,N_45835);
and U46058 (N_46058,N_45847,N_45853);
xor U46059 (N_46059,N_45817,N_45884);
nand U46060 (N_46060,N_45788,N_45935);
nor U46061 (N_46061,N_45896,N_45786);
xnor U46062 (N_46062,N_45978,N_45831);
nor U46063 (N_46063,N_45869,N_45800);
nor U46064 (N_46064,N_45849,N_45815);
and U46065 (N_46065,N_45781,N_45763);
and U46066 (N_46066,N_45754,N_45846);
xor U46067 (N_46067,N_45901,N_45971);
and U46068 (N_46068,N_45821,N_45895);
or U46069 (N_46069,N_45819,N_45779);
nand U46070 (N_46070,N_45905,N_45943);
and U46071 (N_46071,N_45890,N_45939);
nand U46072 (N_46072,N_45922,N_45959);
and U46073 (N_46073,N_45930,N_45946);
nor U46074 (N_46074,N_45919,N_45876);
xor U46075 (N_46075,N_45866,N_45783);
or U46076 (N_46076,N_45764,N_45857);
or U46077 (N_46077,N_45816,N_45805);
nand U46078 (N_46078,N_45902,N_45826);
nor U46079 (N_46079,N_45761,N_45871);
or U46080 (N_46080,N_45829,N_45828);
nor U46081 (N_46081,N_45897,N_45882);
nand U46082 (N_46082,N_45827,N_45920);
nor U46083 (N_46083,N_45837,N_45910);
xnor U46084 (N_46084,N_45969,N_45977);
or U46085 (N_46085,N_45765,N_45842);
and U46086 (N_46086,N_45775,N_45832);
nor U46087 (N_46087,N_45892,N_45768);
nor U46088 (N_46088,N_45918,N_45903);
xnor U46089 (N_46089,N_45758,N_45774);
and U46090 (N_46090,N_45972,N_45925);
or U46091 (N_46091,N_45760,N_45811);
xor U46092 (N_46092,N_45900,N_45790);
nand U46093 (N_46093,N_45820,N_45858);
nor U46094 (N_46094,N_45894,N_45877);
nor U46095 (N_46095,N_45873,N_45962);
and U46096 (N_46096,N_45782,N_45865);
and U46097 (N_46097,N_45970,N_45844);
or U46098 (N_46098,N_45810,N_45881);
nor U46099 (N_46099,N_45950,N_45932);
nand U46100 (N_46100,N_45914,N_45893);
and U46101 (N_46101,N_45996,N_45804);
and U46102 (N_46102,N_45960,N_45855);
nand U46103 (N_46103,N_45813,N_45767);
or U46104 (N_46104,N_45961,N_45803);
nor U46105 (N_46105,N_45836,N_45799);
nand U46106 (N_46106,N_45883,N_45985);
nor U46107 (N_46107,N_45927,N_45944);
and U46108 (N_46108,N_45833,N_45885);
nand U46109 (N_46109,N_45949,N_45752);
or U46110 (N_46110,N_45979,N_45854);
and U46111 (N_46111,N_45983,N_45793);
and U46112 (N_46112,N_45850,N_45958);
xor U46113 (N_46113,N_45924,N_45863);
or U46114 (N_46114,N_45755,N_45941);
and U46115 (N_46115,N_45839,N_45852);
nor U46116 (N_46116,N_45766,N_45957);
nor U46117 (N_46117,N_45867,N_45750);
nor U46118 (N_46118,N_45923,N_45778);
or U46119 (N_46119,N_45825,N_45830);
and U46120 (N_46120,N_45908,N_45928);
and U46121 (N_46121,N_45843,N_45868);
and U46122 (N_46122,N_45757,N_45879);
or U46123 (N_46123,N_45921,N_45976);
nor U46124 (N_46124,N_45940,N_45772);
xnor U46125 (N_46125,N_45917,N_45830);
or U46126 (N_46126,N_45787,N_45752);
nor U46127 (N_46127,N_45824,N_45989);
or U46128 (N_46128,N_45985,N_45893);
xor U46129 (N_46129,N_45980,N_45796);
nand U46130 (N_46130,N_45927,N_45833);
xnor U46131 (N_46131,N_45839,N_45840);
or U46132 (N_46132,N_45992,N_45812);
nor U46133 (N_46133,N_45981,N_45948);
or U46134 (N_46134,N_45894,N_45804);
nor U46135 (N_46135,N_45977,N_45790);
nand U46136 (N_46136,N_45890,N_45766);
or U46137 (N_46137,N_45980,N_45976);
nor U46138 (N_46138,N_45897,N_45866);
nand U46139 (N_46139,N_45907,N_45850);
or U46140 (N_46140,N_45984,N_45782);
and U46141 (N_46141,N_45993,N_45870);
nor U46142 (N_46142,N_45962,N_45875);
nor U46143 (N_46143,N_45750,N_45785);
and U46144 (N_46144,N_45763,N_45921);
or U46145 (N_46145,N_45982,N_45884);
nor U46146 (N_46146,N_45923,N_45908);
and U46147 (N_46147,N_45927,N_45777);
nor U46148 (N_46148,N_45895,N_45948);
nand U46149 (N_46149,N_45751,N_45932);
nand U46150 (N_46150,N_45814,N_45997);
nor U46151 (N_46151,N_45883,N_45923);
nand U46152 (N_46152,N_45904,N_45850);
or U46153 (N_46153,N_45967,N_45842);
or U46154 (N_46154,N_45866,N_45777);
and U46155 (N_46155,N_45750,N_45758);
xnor U46156 (N_46156,N_45776,N_45860);
or U46157 (N_46157,N_45906,N_45839);
nand U46158 (N_46158,N_45929,N_45790);
nor U46159 (N_46159,N_45885,N_45853);
nor U46160 (N_46160,N_45792,N_45816);
and U46161 (N_46161,N_45813,N_45891);
and U46162 (N_46162,N_45816,N_45933);
and U46163 (N_46163,N_45955,N_45976);
nand U46164 (N_46164,N_45850,N_45849);
nor U46165 (N_46165,N_45993,N_45805);
nor U46166 (N_46166,N_45952,N_45856);
xor U46167 (N_46167,N_45939,N_45774);
nand U46168 (N_46168,N_45972,N_45993);
nand U46169 (N_46169,N_45909,N_45778);
or U46170 (N_46170,N_45889,N_45828);
nor U46171 (N_46171,N_45990,N_45881);
or U46172 (N_46172,N_45789,N_45915);
nor U46173 (N_46173,N_45833,N_45882);
nor U46174 (N_46174,N_45924,N_45889);
xor U46175 (N_46175,N_45918,N_45830);
or U46176 (N_46176,N_45869,N_45788);
nor U46177 (N_46177,N_45767,N_45988);
nor U46178 (N_46178,N_45871,N_45951);
xnor U46179 (N_46179,N_45785,N_45788);
or U46180 (N_46180,N_45846,N_45859);
and U46181 (N_46181,N_45773,N_45885);
xor U46182 (N_46182,N_45869,N_45976);
and U46183 (N_46183,N_45960,N_45958);
nor U46184 (N_46184,N_45974,N_45763);
xnor U46185 (N_46185,N_45763,N_45849);
or U46186 (N_46186,N_45804,N_45946);
nand U46187 (N_46187,N_45832,N_45843);
or U46188 (N_46188,N_45972,N_45856);
or U46189 (N_46189,N_45946,N_45829);
nor U46190 (N_46190,N_45809,N_45753);
xor U46191 (N_46191,N_45761,N_45875);
nand U46192 (N_46192,N_45906,N_45921);
nand U46193 (N_46193,N_45819,N_45802);
xor U46194 (N_46194,N_45851,N_45932);
or U46195 (N_46195,N_45771,N_45937);
nor U46196 (N_46196,N_45761,N_45786);
and U46197 (N_46197,N_45774,N_45851);
nor U46198 (N_46198,N_45874,N_45885);
nand U46199 (N_46199,N_45853,N_45930);
xnor U46200 (N_46200,N_45969,N_45884);
or U46201 (N_46201,N_45786,N_45907);
nor U46202 (N_46202,N_45763,N_45851);
or U46203 (N_46203,N_45964,N_45852);
or U46204 (N_46204,N_45912,N_45773);
or U46205 (N_46205,N_45895,N_45836);
xnor U46206 (N_46206,N_45761,N_45973);
and U46207 (N_46207,N_45993,N_45966);
nor U46208 (N_46208,N_45852,N_45832);
nor U46209 (N_46209,N_45860,N_45896);
nor U46210 (N_46210,N_45989,N_45926);
nand U46211 (N_46211,N_45930,N_45840);
nand U46212 (N_46212,N_45783,N_45971);
nor U46213 (N_46213,N_45889,N_45774);
nor U46214 (N_46214,N_45990,N_45963);
xor U46215 (N_46215,N_45944,N_45788);
and U46216 (N_46216,N_45800,N_45906);
and U46217 (N_46217,N_45903,N_45755);
and U46218 (N_46218,N_45823,N_45930);
or U46219 (N_46219,N_45779,N_45916);
nand U46220 (N_46220,N_45934,N_45915);
nor U46221 (N_46221,N_45834,N_45912);
xnor U46222 (N_46222,N_45788,N_45876);
nand U46223 (N_46223,N_45813,N_45971);
and U46224 (N_46224,N_45844,N_45931);
nor U46225 (N_46225,N_45910,N_45886);
and U46226 (N_46226,N_45775,N_45818);
and U46227 (N_46227,N_45779,N_45918);
nor U46228 (N_46228,N_45823,N_45810);
xor U46229 (N_46229,N_45948,N_45982);
nor U46230 (N_46230,N_45951,N_45966);
xor U46231 (N_46231,N_45949,N_45850);
nor U46232 (N_46232,N_45801,N_45928);
and U46233 (N_46233,N_45929,N_45871);
and U46234 (N_46234,N_45861,N_45907);
nor U46235 (N_46235,N_45861,N_45984);
nand U46236 (N_46236,N_45932,N_45900);
and U46237 (N_46237,N_45825,N_45984);
nor U46238 (N_46238,N_45958,N_45785);
nand U46239 (N_46239,N_45801,N_45981);
nor U46240 (N_46240,N_45853,N_45867);
and U46241 (N_46241,N_45767,N_45925);
or U46242 (N_46242,N_45787,N_45841);
and U46243 (N_46243,N_45859,N_45947);
or U46244 (N_46244,N_45902,N_45953);
or U46245 (N_46245,N_45903,N_45952);
and U46246 (N_46246,N_45778,N_45929);
and U46247 (N_46247,N_45958,N_45770);
xnor U46248 (N_46248,N_45979,N_45830);
nor U46249 (N_46249,N_45895,N_45880);
or U46250 (N_46250,N_46047,N_46036);
or U46251 (N_46251,N_46238,N_46041);
and U46252 (N_46252,N_46189,N_46114);
or U46253 (N_46253,N_46219,N_46098);
xnor U46254 (N_46254,N_46110,N_46016);
nand U46255 (N_46255,N_46152,N_46058);
nand U46256 (N_46256,N_46153,N_46086);
and U46257 (N_46257,N_46128,N_46132);
nand U46258 (N_46258,N_46097,N_46164);
xnor U46259 (N_46259,N_46112,N_46147);
xor U46260 (N_46260,N_46077,N_46148);
and U46261 (N_46261,N_46229,N_46082);
nand U46262 (N_46262,N_46145,N_46165);
nor U46263 (N_46263,N_46103,N_46043);
or U46264 (N_46264,N_46139,N_46040);
xnor U46265 (N_46265,N_46166,N_46208);
nand U46266 (N_46266,N_46083,N_46154);
nor U46267 (N_46267,N_46236,N_46020);
nor U46268 (N_46268,N_46242,N_46220);
nor U46269 (N_46269,N_46234,N_46031);
or U46270 (N_46270,N_46158,N_46009);
xnor U46271 (N_46271,N_46194,N_46249);
xnor U46272 (N_46272,N_46201,N_46237);
nor U46273 (N_46273,N_46187,N_46143);
xnor U46274 (N_46274,N_46207,N_46046);
nor U46275 (N_46275,N_46169,N_46095);
nand U46276 (N_46276,N_46063,N_46021);
and U46277 (N_46277,N_46186,N_46074);
nor U46278 (N_46278,N_46006,N_46030);
or U46279 (N_46279,N_46174,N_46087);
nor U46280 (N_46280,N_46068,N_46150);
nand U46281 (N_46281,N_46204,N_46127);
or U46282 (N_46282,N_46039,N_46073);
nand U46283 (N_46283,N_46146,N_46056);
nor U46284 (N_46284,N_46213,N_46115);
or U46285 (N_46285,N_46178,N_46037);
xor U46286 (N_46286,N_46179,N_46203);
and U46287 (N_46287,N_46245,N_46050);
or U46288 (N_46288,N_46069,N_46120);
or U46289 (N_46289,N_46188,N_46010);
or U46290 (N_46290,N_46241,N_46217);
xnor U46291 (N_46291,N_46211,N_46195);
xor U46292 (N_46292,N_46210,N_46027);
xnor U46293 (N_46293,N_46130,N_46025);
and U46294 (N_46294,N_46197,N_46244);
nand U46295 (N_46295,N_46137,N_46038);
or U46296 (N_46296,N_46227,N_46138);
nor U46297 (N_46297,N_46105,N_46026);
or U46298 (N_46298,N_46005,N_46096);
xor U46299 (N_46299,N_46181,N_46091);
xnor U46300 (N_46300,N_46018,N_46045);
xor U46301 (N_46301,N_46042,N_46060);
or U46302 (N_46302,N_46185,N_46012);
nand U46303 (N_46303,N_46136,N_46017);
and U46304 (N_46304,N_46221,N_46001);
or U46305 (N_46305,N_46228,N_46144);
nor U46306 (N_46306,N_46079,N_46084);
nand U46307 (N_46307,N_46033,N_46107);
nor U46308 (N_46308,N_46162,N_46160);
or U46309 (N_46309,N_46072,N_46224);
and U46310 (N_46310,N_46134,N_46081);
nand U46311 (N_46311,N_46131,N_46151);
or U46312 (N_46312,N_46196,N_46167);
and U46313 (N_46313,N_46190,N_46171);
and U46314 (N_46314,N_46226,N_46064);
or U46315 (N_46315,N_46066,N_46168);
and U46316 (N_46316,N_46182,N_46177);
and U46317 (N_46317,N_46109,N_46240);
nor U46318 (N_46318,N_46003,N_46014);
and U46319 (N_46319,N_46004,N_46231);
and U46320 (N_46320,N_46090,N_46156);
nor U46321 (N_46321,N_46239,N_46106);
and U46322 (N_46322,N_46141,N_46123);
xor U46323 (N_46323,N_46053,N_46243);
and U46324 (N_46324,N_46122,N_46117);
xor U46325 (N_46325,N_46089,N_46199);
nand U46326 (N_46326,N_46246,N_46118);
nand U46327 (N_46327,N_46111,N_46214);
or U46328 (N_46328,N_46235,N_46232);
nand U46329 (N_46329,N_46057,N_46008);
nor U46330 (N_46330,N_46015,N_46104);
nand U46331 (N_46331,N_46215,N_46124);
xnor U46332 (N_46332,N_46205,N_46116);
xor U46333 (N_46333,N_46013,N_46065);
and U46334 (N_46334,N_46088,N_46155);
or U46335 (N_46335,N_46175,N_46024);
xor U46336 (N_46336,N_46176,N_46163);
nand U46337 (N_46337,N_46129,N_46075);
or U46338 (N_46338,N_46121,N_46135);
and U46339 (N_46339,N_46035,N_46192);
or U46340 (N_46340,N_46070,N_46059);
nand U46341 (N_46341,N_46200,N_46173);
nand U46342 (N_46342,N_46184,N_46078);
xnor U46343 (N_46343,N_46198,N_46085);
and U46344 (N_46344,N_46092,N_46206);
nor U46345 (N_46345,N_46022,N_46161);
and U46346 (N_46346,N_46071,N_46142);
nor U46347 (N_46347,N_46032,N_46034);
and U46348 (N_46348,N_46108,N_46044);
or U46349 (N_46349,N_46093,N_46202);
xor U46350 (N_46350,N_46140,N_46212);
or U46351 (N_46351,N_46051,N_46218);
xor U46352 (N_46352,N_46172,N_46080);
xnor U46353 (N_46353,N_46223,N_46100);
xnor U46354 (N_46354,N_46052,N_46061);
and U46355 (N_46355,N_46076,N_46054);
or U46356 (N_46356,N_46157,N_46193);
xnor U46357 (N_46357,N_46099,N_46170);
nor U46358 (N_46358,N_46191,N_46247);
and U46359 (N_46359,N_46007,N_46233);
nor U46360 (N_46360,N_46113,N_46230);
nor U46361 (N_46361,N_46216,N_46029);
or U46362 (N_46362,N_46002,N_46149);
and U46363 (N_46363,N_46225,N_46222);
or U46364 (N_46364,N_46101,N_46011);
xor U46365 (N_46365,N_46094,N_46049);
nor U46366 (N_46366,N_46183,N_46126);
nand U46367 (N_46367,N_46180,N_46159);
xnor U46368 (N_46368,N_46209,N_46102);
nand U46369 (N_46369,N_46055,N_46125);
and U46370 (N_46370,N_46133,N_46023);
xnor U46371 (N_46371,N_46119,N_46028);
nand U46372 (N_46372,N_46067,N_46019);
nor U46373 (N_46373,N_46048,N_46248);
or U46374 (N_46374,N_46000,N_46062);
and U46375 (N_46375,N_46005,N_46004);
xnor U46376 (N_46376,N_46221,N_46147);
nor U46377 (N_46377,N_46092,N_46154);
nor U46378 (N_46378,N_46088,N_46106);
and U46379 (N_46379,N_46073,N_46062);
xor U46380 (N_46380,N_46062,N_46190);
and U46381 (N_46381,N_46187,N_46063);
and U46382 (N_46382,N_46073,N_46146);
and U46383 (N_46383,N_46061,N_46164);
or U46384 (N_46384,N_46177,N_46249);
and U46385 (N_46385,N_46222,N_46228);
and U46386 (N_46386,N_46143,N_46107);
xor U46387 (N_46387,N_46124,N_46197);
nor U46388 (N_46388,N_46163,N_46220);
xnor U46389 (N_46389,N_46057,N_46177);
nand U46390 (N_46390,N_46214,N_46123);
xnor U46391 (N_46391,N_46054,N_46022);
or U46392 (N_46392,N_46019,N_46003);
or U46393 (N_46393,N_46020,N_46045);
nor U46394 (N_46394,N_46199,N_46101);
or U46395 (N_46395,N_46236,N_46235);
xor U46396 (N_46396,N_46174,N_46128);
nor U46397 (N_46397,N_46137,N_46028);
nor U46398 (N_46398,N_46075,N_46191);
nor U46399 (N_46399,N_46218,N_46229);
nand U46400 (N_46400,N_46083,N_46048);
nand U46401 (N_46401,N_46219,N_46026);
or U46402 (N_46402,N_46187,N_46140);
nor U46403 (N_46403,N_46134,N_46038);
xnor U46404 (N_46404,N_46059,N_46046);
nor U46405 (N_46405,N_46208,N_46087);
or U46406 (N_46406,N_46089,N_46178);
or U46407 (N_46407,N_46104,N_46054);
nor U46408 (N_46408,N_46199,N_46190);
and U46409 (N_46409,N_46144,N_46052);
xor U46410 (N_46410,N_46245,N_46073);
nand U46411 (N_46411,N_46072,N_46001);
nor U46412 (N_46412,N_46040,N_46245);
and U46413 (N_46413,N_46012,N_46035);
nand U46414 (N_46414,N_46089,N_46053);
nor U46415 (N_46415,N_46113,N_46162);
nor U46416 (N_46416,N_46065,N_46218);
and U46417 (N_46417,N_46128,N_46218);
xor U46418 (N_46418,N_46045,N_46107);
or U46419 (N_46419,N_46239,N_46078);
nor U46420 (N_46420,N_46042,N_46030);
and U46421 (N_46421,N_46081,N_46208);
nand U46422 (N_46422,N_46023,N_46244);
and U46423 (N_46423,N_46131,N_46229);
xor U46424 (N_46424,N_46156,N_46016);
or U46425 (N_46425,N_46107,N_46007);
and U46426 (N_46426,N_46245,N_46200);
or U46427 (N_46427,N_46031,N_46140);
nand U46428 (N_46428,N_46167,N_46107);
xor U46429 (N_46429,N_46029,N_46086);
nand U46430 (N_46430,N_46053,N_46068);
and U46431 (N_46431,N_46190,N_46098);
xor U46432 (N_46432,N_46068,N_46100);
nor U46433 (N_46433,N_46224,N_46060);
or U46434 (N_46434,N_46178,N_46202);
nor U46435 (N_46435,N_46081,N_46195);
xnor U46436 (N_46436,N_46035,N_46062);
or U46437 (N_46437,N_46058,N_46053);
or U46438 (N_46438,N_46241,N_46123);
nand U46439 (N_46439,N_46186,N_46155);
or U46440 (N_46440,N_46015,N_46101);
nand U46441 (N_46441,N_46208,N_46004);
nand U46442 (N_46442,N_46045,N_46207);
nand U46443 (N_46443,N_46157,N_46247);
or U46444 (N_46444,N_46199,N_46024);
and U46445 (N_46445,N_46094,N_46096);
nand U46446 (N_46446,N_46166,N_46093);
nor U46447 (N_46447,N_46214,N_46072);
xor U46448 (N_46448,N_46058,N_46002);
and U46449 (N_46449,N_46185,N_46183);
nand U46450 (N_46450,N_46008,N_46211);
nor U46451 (N_46451,N_46017,N_46107);
or U46452 (N_46452,N_46152,N_46165);
xor U46453 (N_46453,N_46060,N_46222);
and U46454 (N_46454,N_46171,N_46191);
xor U46455 (N_46455,N_46044,N_46234);
xnor U46456 (N_46456,N_46178,N_46029);
xnor U46457 (N_46457,N_46003,N_46236);
nand U46458 (N_46458,N_46015,N_46237);
xor U46459 (N_46459,N_46155,N_46045);
or U46460 (N_46460,N_46107,N_46058);
or U46461 (N_46461,N_46121,N_46143);
nor U46462 (N_46462,N_46060,N_46163);
nand U46463 (N_46463,N_46187,N_46112);
or U46464 (N_46464,N_46188,N_46151);
nand U46465 (N_46465,N_46034,N_46157);
xor U46466 (N_46466,N_46234,N_46023);
nand U46467 (N_46467,N_46167,N_46248);
or U46468 (N_46468,N_46157,N_46050);
xnor U46469 (N_46469,N_46065,N_46027);
or U46470 (N_46470,N_46019,N_46161);
nor U46471 (N_46471,N_46057,N_46190);
xor U46472 (N_46472,N_46204,N_46153);
nand U46473 (N_46473,N_46008,N_46230);
and U46474 (N_46474,N_46121,N_46111);
nor U46475 (N_46475,N_46197,N_46032);
and U46476 (N_46476,N_46161,N_46222);
xnor U46477 (N_46477,N_46154,N_46169);
nor U46478 (N_46478,N_46178,N_46105);
or U46479 (N_46479,N_46038,N_46022);
nand U46480 (N_46480,N_46248,N_46086);
xor U46481 (N_46481,N_46219,N_46198);
nor U46482 (N_46482,N_46137,N_46057);
and U46483 (N_46483,N_46089,N_46103);
nor U46484 (N_46484,N_46081,N_46115);
nor U46485 (N_46485,N_46202,N_46160);
or U46486 (N_46486,N_46067,N_46060);
nand U46487 (N_46487,N_46138,N_46194);
and U46488 (N_46488,N_46184,N_46027);
and U46489 (N_46489,N_46140,N_46008);
xnor U46490 (N_46490,N_46108,N_46101);
or U46491 (N_46491,N_46127,N_46209);
nor U46492 (N_46492,N_46039,N_46162);
nor U46493 (N_46493,N_46030,N_46016);
xnor U46494 (N_46494,N_46115,N_46002);
or U46495 (N_46495,N_46087,N_46017);
and U46496 (N_46496,N_46182,N_46205);
nor U46497 (N_46497,N_46197,N_46058);
and U46498 (N_46498,N_46016,N_46229);
nor U46499 (N_46499,N_46096,N_46015);
nor U46500 (N_46500,N_46276,N_46439);
nor U46501 (N_46501,N_46264,N_46433);
and U46502 (N_46502,N_46283,N_46446);
nor U46503 (N_46503,N_46391,N_46437);
xor U46504 (N_46504,N_46357,N_46275);
nand U46505 (N_46505,N_46288,N_46420);
xnor U46506 (N_46506,N_46473,N_46431);
nor U46507 (N_46507,N_46432,N_46422);
nor U46508 (N_46508,N_46396,N_46408);
nor U46509 (N_46509,N_46333,N_46454);
and U46510 (N_46510,N_46321,N_46470);
nor U46511 (N_46511,N_46499,N_46462);
xor U46512 (N_46512,N_46477,N_46471);
xor U46513 (N_46513,N_46443,N_46486);
or U46514 (N_46514,N_46378,N_46384);
xor U46515 (N_46515,N_46330,N_46488);
nor U46516 (N_46516,N_46303,N_46375);
xor U46517 (N_46517,N_46365,N_46340);
nand U46518 (N_46518,N_46417,N_46299);
or U46519 (N_46519,N_46329,N_46402);
nand U46520 (N_46520,N_46398,N_46259);
or U46521 (N_46521,N_46412,N_46325);
or U46522 (N_46522,N_46387,N_46388);
nand U46523 (N_46523,N_46421,N_46348);
and U46524 (N_46524,N_46338,N_46260);
nor U46525 (N_46525,N_46465,N_46363);
and U46526 (N_46526,N_46304,N_46290);
and U46527 (N_46527,N_46377,N_46278);
or U46528 (N_46528,N_46293,N_46425);
nand U46529 (N_46529,N_46460,N_46267);
nor U46530 (N_46530,N_46487,N_46492);
or U46531 (N_46531,N_46282,N_46406);
or U46532 (N_46532,N_46478,N_46281);
nor U46533 (N_46533,N_46482,N_46258);
nor U46534 (N_46534,N_46450,N_46494);
nand U46535 (N_46535,N_46400,N_46265);
nand U46536 (N_46536,N_46262,N_46289);
nor U46537 (N_46537,N_46453,N_46409);
nand U46538 (N_46538,N_46383,N_46356);
nand U46539 (N_46539,N_46498,N_46419);
nand U46540 (N_46540,N_46274,N_46269);
xnor U46541 (N_46541,N_46305,N_46351);
or U46542 (N_46542,N_46287,N_46292);
xnor U46543 (N_46543,N_46393,N_46251);
xnor U46544 (N_46544,N_46364,N_46355);
xnor U46545 (N_46545,N_46342,N_46445);
nor U46546 (N_46546,N_46277,N_46261);
nand U46547 (N_46547,N_46253,N_46327);
and U46548 (N_46548,N_46279,N_46373);
nand U46549 (N_46549,N_46440,N_46472);
nor U46550 (N_46550,N_46266,N_46497);
or U46551 (N_46551,N_46339,N_46313);
xor U46552 (N_46552,N_46294,N_46345);
nand U46553 (N_46553,N_46270,N_46395);
xnor U46554 (N_46554,N_46370,N_46320);
xnor U46555 (N_46555,N_46254,N_46436);
nor U46556 (N_46556,N_46314,N_46343);
nor U46557 (N_46557,N_46347,N_46427);
or U46558 (N_46558,N_46268,N_46297);
or U46559 (N_46559,N_46369,N_46332);
xor U46560 (N_46560,N_46256,N_46317);
nor U46561 (N_46561,N_46481,N_46309);
or U46562 (N_46562,N_46374,N_46456);
nor U46563 (N_46563,N_46405,N_46380);
or U46564 (N_46564,N_46467,N_46263);
nand U46565 (N_46565,N_46415,N_46366);
and U46566 (N_46566,N_46397,N_46344);
xor U46567 (N_46567,N_46490,N_46455);
nor U46568 (N_46568,N_46407,N_46452);
nand U46569 (N_46569,N_46441,N_46449);
xnor U46570 (N_46570,N_46352,N_46485);
nor U46571 (N_46571,N_46484,N_46381);
nand U46572 (N_46572,N_46362,N_46444);
or U46573 (N_46573,N_46479,N_46495);
nand U46574 (N_46574,N_46295,N_46350);
or U46575 (N_46575,N_46346,N_46358);
nor U46576 (N_46576,N_46489,N_46447);
xor U46577 (N_46577,N_46410,N_46442);
xor U46578 (N_46578,N_46308,N_46475);
or U46579 (N_46579,N_46315,N_46458);
or U46580 (N_46580,N_46414,N_46413);
xor U46581 (N_46581,N_46483,N_46349);
nand U46582 (N_46582,N_46326,N_46335);
or U46583 (N_46583,N_46418,N_46311);
or U46584 (N_46584,N_46493,N_46361);
and U46585 (N_46585,N_46469,N_46360);
and U46586 (N_46586,N_46296,N_46322);
xnor U46587 (N_46587,N_46371,N_46491);
and U46588 (N_46588,N_46429,N_46323);
and U46589 (N_46589,N_46411,N_46389);
xnor U46590 (N_46590,N_46298,N_46312);
nand U46591 (N_46591,N_46310,N_46319);
nand U46592 (N_46592,N_46376,N_46341);
or U46593 (N_46593,N_46336,N_46461);
and U46594 (N_46594,N_46424,N_46318);
or U46595 (N_46595,N_46480,N_46307);
nor U46596 (N_46596,N_46291,N_46386);
and U46597 (N_46597,N_46337,N_46331);
and U46598 (N_46598,N_46434,N_46401);
nand U46599 (N_46599,N_46379,N_46328);
xnor U46600 (N_46600,N_46451,N_46468);
or U46601 (N_46601,N_46316,N_46250);
nor U46602 (N_46602,N_46416,N_46367);
nor U46603 (N_46603,N_46476,N_46435);
and U46604 (N_46604,N_46272,N_46403);
xnor U46605 (N_46605,N_46428,N_46334);
and U46606 (N_46606,N_46423,N_46385);
or U46607 (N_46607,N_46463,N_46457);
nand U46608 (N_46608,N_46255,N_46252);
and U46609 (N_46609,N_46286,N_46448);
nand U46610 (N_46610,N_46399,N_46301);
nor U46611 (N_46611,N_46392,N_46474);
nor U46612 (N_46612,N_46271,N_46353);
nand U46613 (N_46613,N_46324,N_46430);
nor U46614 (N_46614,N_46372,N_46285);
or U46615 (N_46615,N_46426,N_46280);
xor U46616 (N_46616,N_46306,N_46464);
or U46617 (N_46617,N_46390,N_46300);
xor U46618 (N_46618,N_46354,N_46368);
or U46619 (N_46619,N_46257,N_46459);
xnor U46620 (N_46620,N_46273,N_46466);
and U46621 (N_46621,N_46359,N_46496);
or U46622 (N_46622,N_46394,N_46284);
nand U46623 (N_46623,N_46382,N_46438);
nor U46624 (N_46624,N_46302,N_46404);
nor U46625 (N_46625,N_46270,N_46311);
nor U46626 (N_46626,N_46480,N_46456);
xnor U46627 (N_46627,N_46424,N_46438);
nor U46628 (N_46628,N_46311,N_46261);
nand U46629 (N_46629,N_46339,N_46453);
and U46630 (N_46630,N_46415,N_46347);
and U46631 (N_46631,N_46331,N_46313);
nor U46632 (N_46632,N_46263,N_46290);
nand U46633 (N_46633,N_46384,N_46336);
and U46634 (N_46634,N_46459,N_46406);
nor U46635 (N_46635,N_46496,N_46267);
nand U46636 (N_46636,N_46400,N_46441);
or U46637 (N_46637,N_46455,N_46393);
nand U46638 (N_46638,N_46285,N_46470);
xor U46639 (N_46639,N_46355,N_46287);
nor U46640 (N_46640,N_46252,N_46462);
nand U46641 (N_46641,N_46451,N_46310);
or U46642 (N_46642,N_46384,N_46444);
xor U46643 (N_46643,N_46316,N_46342);
or U46644 (N_46644,N_46336,N_46450);
xor U46645 (N_46645,N_46272,N_46260);
xor U46646 (N_46646,N_46264,N_46324);
or U46647 (N_46647,N_46329,N_46264);
or U46648 (N_46648,N_46302,N_46496);
and U46649 (N_46649,N_46391,N_46287);
nor U46650 (N_46650,N_46372,N_46250);
nand U46651 (N_46651,N_46382,N_46371);
xnor U46652 (N_46652,N_46310,N_46450);
nand U46653 (N_46653,N_46316,N_46493);
nand U46654 (N_46654,N_46428,N_46289);
and U46655 (N_46655,N_46258,N_46296);
and U46656 (N_46656,N_46434,N_46363);
nor U46657 (N_46657,N_46440,N_46346);
nor U46658 (N_46658,N_46329,N_46314);
xnor U46659 (N_46659,N_46400,N_46449);
or U46660 (N_46660,N_46458,N_46378);
or U46661 (N_46661,N_46359,N_46397);
nand U46662 (N_46662,N_46447,N_46456);
nor U46663 (N_46663,N_46261,N_46460);
nand U46664 (N_46664,N_46259,N_46276);
nor U46665 (N_46665,N_46491,N_46303);
or U46666 (N_46666,N_46369,N_46446);
and U46667 (N_46667,N_46438,N_46465);
and U46668 (N_46668,N_46312,N_46416);
nand U46669 (N_46669,N_46271,N_46459);
nor U46670 (N_46670,N_46327,N_46318);
and U46671 (N_46671,N_46477,N_46459);
xnor U46672 (N_46672,N_46362,N_46419);
nand U46673 (N_46673,N_46398,N_46490);
xor U46674 (N_46674,N_46371,N_46414);
and U46675 (N_46675,N_46475,N_46369);
xor U46676 (N_46676,N_46374,N_46306);
xor U46677 (N_46677,N_46282,N_46469);
xnor U46678 (N_46678,N_46465,N_46376);
nand U46679 (N_46679,N_46371,N_46489);
nor U46680 (N_46680,N_46265,N_46483);
nand U46681 (N_46681,N_46342,N_46464);
nor U46682 (N_46682,N_46455,N_46425);
nand U46683 (N_46683,N_46281,N_46398);
xnor U46684 (N_46684,N_46436,N_46392);
nor U46685 (N_46685,N_46482,N_46377);
nand U46686 (N_46686,N_46404,N_46458);
and U46687 (N_46687,N_46301,N_46417);
nor U46688 (N_46688,N_46403,N_46362);
and U46689 (N_46689,N_46358,N_46496);
or U46690 (N_46690,N_46348,N_46320);
xor U46691 (N_46691,N_46480,N_46299);
or U46692 (N_46692,N_46487,N_46369);
nand U46693 (N_46693,N_46399,N_46319);
and U46694 (N_46694,N_46261,N_46387);
nor U46695 (N_46695,N_46494,N_46439);
or U46696 (N_46696,N_46435,N_46364);
or U46697 (N_46697,N_46269,N_46420);
or U46698 (N_46698,N_46438,N_46377);
or U46699 (N_46699,N_46288,N_46257);
nand U46700 (N_46700,N_46316,N_46465);
xor U46701 (N_46701,N_46387,N_46424);
xor U46702 (N_46702,N_46458,N_46471);
xor U46703 (N_46703,N_46460,N_46327);
or U46704 (N_46704,N_46328,N_46494);
nand U46705 (N_46705,N_46323,N_46484);
or U46706 (N_46706,N_46328,N_46440);
nand U46707 (N_46707,N_46250,N_46297);
or U46708 (N_46708,N_46294,N_46300);
nand U46709 (N_46709,N_46289,N_46336);
and U46710 (N_46710,N_46308,N_46343);
or U46711 (N_46711,N_46409,N_46286);
nand U46712 (N_46712,N_46469,N_46417);
and U46713 (N_46713,N_46438,N_46470);
nand U46714 (N_46714,N_46437,N_46392);
nand U46715 (N_46715,N_46456,N_46277);
nor U46716 (N_46716,N_46472,N_46303);
nand U46717 (N_46717,N_46496,N_46466);
nand U46718 (N_46718,N_46435,N_46382);
nor U46719 (N_46719,N_46451,N_46406);
and U46720 (N_46720,N_46482,N_46397);
or U46721 (N_46721,N_46387,N_46484);
and U46722 (N_46722,N_46394,N_46256);
or U46723 (N_46723,N_46327,N_46478);
and U46724 (N_46724,N_46325,N_46338);
xor U46725 (N_46725,N_46460,N_46474);
or U46726 (N_46726,N_46319,N_46445);
xnor U46727 (N_46727,N_46417,N_46323);
or U46728 (N_46728,N_46306,N_46302);
or U46729 (N_46729,N_46425,N_46430);
xor U46730 (N_46730,N_46447,N_46337);
nor U46731 (N_46731,N_46269,N_46334);
and U46732 (N_46732,N_46363,N_46460);
nor U46733 (N_46733,N_46491,N_46337);
and U46734 (N_46734,N_46491,N_46498);
and U46735 (N_46735,N_46396,N_46415);
nand U46736 (N_46736,N_46384,N_46439);
and U46737 (N_46737,N_46457,N_46492);
xnor U46738 (N_46738,N_46316,N_46478);
xor U46739 (N_46739,N_46365,N_46416);
and U46740 (N_46740,N_46481,N_46466);
or U46741 (N_46741,N_46481,N_46311);
and U46742 (N_46742,N_46439,N_46416);
nor U46743 (N_46743,N_46348,N_46331);
and U46744 (N_46744,N_46254,N_46449);
xor U46745 (N_46745,N_46379,N_46320);
xor U46746 (N_46746,N_46344,N_46262);
or U46747 (N_46747,N_46418,N_46499);
and U46748 (N_46748,N_46439,N_46356);
and U46749 (N_46749,N_46441,N_46261);
and U46750 (N_46750,N_46569,N_46736);
and U46751 (N_46751,N_46657,N_46525);
nor U46752 (N_46752,N_46587,N_46722);
xor U46753 (N_46753,N_46519,N_46524);
nor U46754 (N_46754,N_46595,N_46656);
xnor U46755 (N_46755,N_46568,N_46682);
nor U46756 (N_46756,N_46522,N_46585);
or U46757 (N_46757,N_46741,N_46548);
or U46758 (N_46758,N_46734,N_46534);
nand U46759 (N_46759,N_46581,N_46579);
nor U46760 (N_46760,N_46537,N_46635);
nand U46761 (N_46761,N_46527,N_46673);
xnor U46762 (N_46762,N_46624,N_46670);
or U46763 (N_46763,N_46705,N_46714);
nor U46764 (N_46764,N_46557,N_46598);
xor U46765 (N_46765,N_46500,N_46570);
nand U46766 (N_46766,N_46743,N_46501);
nor U46767 (N_46767,N_46550,N_46720);
nand U46768 (N_46768,N_46749,N_46707);
and U46769 (N_46769,N_46612,N_46697);
xnor U46770 (N_46770,N_46647,N_46592);
xnor U46771 (N_46771,N_46577,N_46559);
xor U46772 (N_46772,N_46605,N_46502);
xnor U46773 (N_46773,N_46694,N_46740);
or U46774 (N_46774,N_46589,N_46591);
and U46775 (N_46775,N_46718,N_46688);
nand U46776 (N_46776,N_46563,N_46703);
nor U46777 (N_46777,N_46683,N_46737);
nor U46778 (N_46778,N_46690,N_46669);
and U46779 (N_46779,N_46629,N_46662);
nand U46780 (N_46780,N_46611,N_46599);
xnor U46781 (N_46781,N_46632,N_46729);
nand U46782 (N_46782,N_46544,N_46521);
nand U46783 (N_46783,N_46681,N_46618);
and U46784 (N_46784,N_46564,N_46721);
nand U46785 (N_46785,N_46584,N_46560);
and U46786 (N_46786,N_46710,N_46551);
xnor U46787 (N_46787,N_46706,N_46529);
nand U46788 (N_46788,N_46555,N_46696);
and U46789 (N_46789,N_46651,N_46704);
nand U46790 (N_46790,N_46746,N_46613);
nand U46791 (N_46791,N_46539,N_46649);
nor U46792 (N_46792,N_46660,N_46672);
xnor U46793 (N_46793,N_46634,N_46620);
and U46794 (N_46794,N_46713,N_46742);
or U46795 (N_46795,N_46685,N_46687);
xnor U46796 (N_46796,N_46523,N_46546);
or U46797 (N_46797,N_46668,N_46545);
nand U46798 (N_46798,N_46726,N_46671);
or U46799 (N_46799,N_46650,N_46695);
or U46800 (N_46800,N_46715,N_46562);
and U46801 (N_46801,N_46666,N_46526);
or U46802 (N_46802,N_46588,N_46616);
xor U46803 (N_46803,N_46607,N_46640);
nand U46804 (N_46804,N_46590,N_46693);
nand U46805 (N_46805,N_46549,N_46573);
and U46806 (N_46806,N_46745,N_46617);
xnor U46807 (N_46807,N_46597,N_46503);
or U46808 (N_46808,N_46692,N_46552);
xnor U46809 (N_46809,N_46645,N_46731);
and U46810 (N_46810,N_46725,N_46514);
and U46811 (N_46811,N_46504,N_46700);
or U46812 (N_46812,N_46637,N_46636);
nor U46813 (N_46813,N_46604,N_46702);
or U46814 (N_46814,N_46512,N_46728);
and U46815 (N_46815,N_46648,N_46578);
xor U46816 (N_46816,N_46628,N_46665);
and U46817 (N_46817,N_46533,N_46679);
or U46818 (N_46818,N_46606,N_46517);
and U46819 (N_46819,N_46621,N_46507);
and U46820 (N_46820,N_46542,N_46506);
nor U46821 (N_46821,N_46653,N_46732);
nand U46822 (N_46822,N_46646,N_46639);
nor U46823 (N_46823,N_46593,N_46615);
or U46824 (N_46824,N_46691,N_46667);
nand U46825 (N_46825,N_46554,N_46642);
and U46826 (N_46826,N_46735,N_46717);
and U46827 (N_46827,N_46515,N_46747);
and U46828 (N_46828,N_46509,N_46608);
and U46829 (N_46829,N_46596,N_46716);
nand U46830 (N_46830,N_46709,N_46586);
nor U46831 (N_46831,N_46603,N_46520);
or U46832 (N_46832,N_46719,N_46582);
nand U46833 (N_46833,N_46677,N_46583);
xor U46834 (N_46834,N_46712,N_46518);
and U46835 (N_46835,N_46727,N_46575);
or U46836 (N_46836,N_46609,N_46508);
and U46837 (N_46837,N_46571,N_46708);
nor U46838 (N_46838,N_46625,N_46567);
nor U46839 (N_46839,N_46580,N_46678);
xnor U46840 (N_46840,N_46619,N_46684);
xor U46841 (N_46841,N_46652,N_46744);
xnor U46842 (N_46842,N_46531,N_46516);
and U46843 (N_46843,N_46643,N_46664);
xnor U46844 (N_46844,N_46574,N_46676);
nor U46845 (N_46845,N_46535,N_46638);
xnor U46846 (N_46846,N_46663,N_46543);
or U46847 (N_46847,N_46623,N_46556);
nor U46848 (N_46848,N_46601,N_46627);
or U46849 (N_46849,N_46622,N_46644);
nand U46850 (N_46850,N_46655,N_46633);
or U46851 (N_46851,N_46699,N_46654);
nor U46852 (N_46852,N_46738,N_46674);
xor U46853 (N_46853,N_46566,N_46602);
xor U46854 (N_46854,N_46675,N_46547);
and U46855 (N_46855,N_46733,N_46594);
nand U46856 (N_46856,N_46530,N_46610);
nand U46857 (N_46857,N_46661,N_46614);
nor U46858 (N_46858,N_46565,N_46630);
xor U46859 (N_46859,N_46626,N_46553);
nor U46860 (N_46860,N_46558,N_46711);
nand U46861 (N_46861,N_46748,N_46528);
nor U46862 (N_46862,N_46730,N_46561);
or U46863 (N_46863,N_46698,N_46689);
or U46864 (N_46864,N_46641,N_46540);
or U46865 (N_46865,N_46505,N_46572);
nor U46866 (N_46866,N_46576,N_46541);
nor U46867 (N_46867,N_46600,N_46536);
nand U46868 (N_46868,N_46739,N_46538);
nor U46869 (N_46869,N_46532,N_46659);
nor U46870 (N_46870,N_46510,N_46680);
nand U46871 (N_46871,N_46658,N_46723);
and U46872 (N_46872,N_46513,N_46724);
xnor U46873 (N_46873,N_46701,N_46686);
and U46874 (N_46874,N_46631,N_46511);
nor U46875 (N_46875,N_46737,N_46623);
and U46876 (N_46876,N_46632,N_46744);
or U46877 (N_46877,N_46673,N_46622);
or U46878 (N_46878,N_46551,N_46556);
nand U46879 (N_46879,N_46588,N_46501);
xor U46880 (N_46880,N_46544,N_46747);
and U46881 (N_46881,N_46700,N_46652);
nand U46882 (N_46882,N_46582,N_46633);
nand U46883 (N_46883,N_46694,N_46742);
and U46884 (N_46884,N_46629,N_46569);
and U46885 (N_46885,N_46660,N_46738);
nor U46886 (N_46886,N_46714,N_46748);
or U46887 (N_46887,N_46690,N_46609);
nor U46888 (N_46888,N_46706,N_46620);
or U46889 (N_46889,N_46719,N_46609);
xnor U46890 (N_46890,N_46660,N_46718);
or U46891 (N_46891,N_46691,N_46579);
nor U46892 (N_46892,N_46544,N_46647);
nand U46893 (N_46893,N_46557,N_46558);
and U46894 (N_46894,N_46660,N_46588);
nor U46895 (N_46895,N_46720,N_46702);
and U46896 (N_46896,N_46538,N_46712);
nand U46897 (N_46897,N_46620,N_46692);
nor U46898 (N_46898,N_46626,N_46558);
or U46899 (N_46899,N_46551,N_46570);
xor U46900 (N_46900,N_46521,N_46567);
nor U46901 (N_46901,N_46520,N_46680);
nand U46902 (N_46902,N_46657,N_46630);
and U46903 (N_46903,N_46541,N_46554);
or U46904 (N_46904,N_46699,N_46749);
xnor U46905 (N_46905,N_46586,N_46726);
or U46906 (N_46906,N_46716,N_46538);
and U46907 (N_46907,N_46618,N_46540);
nand U46908 (N_46908,N_46576,N_46702);
nor U46909 (N_46909,N_46627,N_46611);
xor U46910 (N_46910,N_46663,N_46599);
xor U46911 (N_46911,N_46514,N_46577);
nor U46912 (N_46912,N_46611,N_46647);
nor U46913 (N_46913,N_46662,N_46581);
nand U46914 (N_46914,N_46523,N_46718);
nor U46915 (N_46915,N_46555,N_46543);
xnor U46916 (N_46916,N_46644,N_46519);
nand U46917 (N_46917,N_46646,N_46597);
and U46918 (N_46918,N_46639,N_46553);
xor U46919 (N_46919,N_46524,N_46699);
and U46920 (N_46920,N_46586,N_46649);
xor U46921 (N_46921,N_46721,N_46725);
nor U46922 (N_46922,N_46576,N_46711);
xor U46923 (N_46923,N_46587,N_46565);
nand U46924 (N_46924,N_46655,N_46578);
nor U46925 (N_46925,N_46631,N_46603);
nand U46926 (N_46926,N_46558,N_46538);
and U46927 (N_46927,N_46696,N_46600);
nor U46928 (N_46928,N_46575,N_46506);
and U46929 (N_46929,N_46529,N_46542);
or U46930 (N_46930,N_46544,N_46523);
or U46931 (N_46931,N_46600,N_46511);
nor U46932 (N_46932,N_46517,N_46505);
and U46933 (N_46933,N_46619,N_46519);
xor U46934 (N_46934,N_46633,N_46537);
nor U46935 (N_46935,N_46508,N_46526);
nand U46936 (N_46936,N_46643,N_46539);
or U46937 (N_46937,N_46591,N_46642);
or U46938 (N_46938,N_46625,N_46713);
or U46939 (N_46939,N_46524,N_46624);
nand U46940 (N_46940,N_46538,N_46599);
nor U46941 (N_46941,N_46676,N_46601);
nand U46942 (N_46942,N_46689,N_46675);
nand U46943 (N_46943,N_46687,N_46743);
or U46944 (N_46944,N_46571,N_46634);
xor U46945 (N_46945,N_46625,N_46614);
nand U46946 (N_46946,N_46536,N_46679);
xor U46947 (N_46947,N_46604,N_46520);
and U46948 (N_46948,N_46500,N_46732);
nor U46949 (N_46949,N_46590,N_46583);
nor U46950 (N_46950,N_46543,N_46622);
and U46951 (N_46951,N_46705,N_46709);
or U46952 (N_46952,N_46518,N_46746);
xor U46953 (N_46953,N_46645,N_46633);
and U46954 (N_46954,N_46561,N_46582);
nand U46955 (N_46955,N_46627,N_46641);
or U46956 (N_46956,N_46621,N_46652);
and U46957 (N_46957,N_46646,N_46616);
nor U46958 (N_46958,N_46532,N_46578);
and U46959 (N_46959,N_46526,N_46523);
nor U46960 (N_46960,N_46730,N_46674);
and U46961 (N_46961,N_46523,N_46663);
nand U46962 (N_46962,N_46580,N_46633);
nand U46963 (N_46963,N_46622,N_46558);
xnor U46964 (N_46964,N_46748,N_46561);
and U46965 (N_46965,N_46541,N_46625);
xnor U46966 (N_46966,N_46528,N_46563);
nor U46967 (N_46967,N_46518,N_46724);
xnor U46968 (N_46968,N_46567,N_46618);
or U46969 (N_46969,N_46704,N_46707);
nand U46970 (N_46970,N_46529,N_46659);
xor U46971 (N_46971,N_46609,N_46701);
nand U46972 (N_46972,N_46502,N_46657);
nand U46973 (N_46973,N_46709,N_46523);
xnor U46974 (N_46974,N_46516,N_46662);
and U46975 (N_46975,N_46647,N_46512);
and U46976 (N_46976,N_46649,N_46565);
nor U46977 (N_46977,N_46531,N_46654);
xor U46978 (N_46978,N_46572,N_46678);
nor U46979 (N_46979,N_46689,N_46593);
nor U46980 (N_46980,N_46541,N_46686);
and U46981 (N_46981,N_46634,N_46530);
or U46982 (N_46982,N_46661,N_46514);
nand U46983 (N_46983,N_46691,N_46562);
or U46984 (N_46984,N_46509,N_46662);
xor U46985 (N_46985,N_46577,N_46699);
xnor U46986 (N_46986,N_46606,N_46663);
or U46987 (N_46987,N_46694,N_46621);
or U46988 (N_46988,N_46570,N_46613);
nor U46989 (N_46989,N_46571,N_46525);
xor U46990 (N_46990,N_46508,N_46727);
or U46991 (N_46991,N_46635,N_46615);
and U46992 (N_46992,N_46633,N_46678);
and U46993 (N_46993,N_46648,N_46715);
or U46994 (N_46994,N_46674,N_46532);
xor U46995 (N_46995,N_46591,N_46513);
nand U46996 (N_46996,N_46567,N_46747);
xnor U46997 (N_46997,N_46645,N_46631);
and U46998 (N_46998,N_46507,N_46619);
xnor U46999 (N_46999,N_46685,N_46654);
or U47000 (N_47000,N_46972,N_46961);
and U47001 (N_47001,N_46832,N_46788);
or U47002 (N_47002,N_46858,N_46865);
xor U47003 (N_47003,N_46946,N_46848);
and U47004 (N_47004,N_46779,N_46979);
xor U47005 (N_47005,N_46884,N_46840);
and U47006 (N_47006,N_46758,N_46815);
xnor U47007 (N_47007,N_46837,N_46846);
or U47008 (N_47008,N_46803,N_46906);
nand U47009 (N_47009,N_46992,N_46915);
xnor U47010 (N_47010,N_46921,N_46863);
xnor U47011 (N_47011,N_46957,N_46860);
nand U47012 (N_47012,N_46785,N_46952);
or U47013 (N_47013,N_46804,N_46967);
and U47014 (N_47014,N_46930,N_46867);
xor U47015 (N_47015,N_46920,N_46782);
xor U47016 (N_47016,N_46950,N_46931);
xnor U47017 (N_47017,N_46987,N_46770);
or U47018 (N_47018,N_46787,N_46869);
or U47019 (N_47019,N_46943,N_46900);
nand U47020 (N_47020,N_46813,N_46773);
and U47021 (N_47021,N_46754,N_46861);
nand U47022 (N_47022,N_46995,N_46970);
xor U47023 (N_47023,N_46802,N_46766);
or U47024 (N_47024,N_46775,N_46821);
or U47025 (N_47025,N_46897,N_46866);
or U47026 (N_47026,N_46889,N_46940);
xor U47027 (N_47027,N_46907,N_46912);
nand U47028 (N_47028,N_46896,N_46820);
and U47029 (N_47029,N_46951,N_46971);
or U47030 (N_47030,N_46856,N_46903);
or U47031 (N_47031,N_46895,N_46978);
xor U47032 (N_47032,N_46893,N_46885);
xor U47033 (N_47033,N_46894,N_46990);
or U47034 (N_47034,N_46963,N_46964);
and U47035 (N_47035,N_46752,N_46826);
and U47036 (N_47036,N_46795,N_46917);
or U47037 (N_47037,N_46793,N_46960);
nor U47038 (N_47038,N_46852,N_46844);
xor U47039 (N_47039,N_46945,N_46872);
or U47040 (N_47040,N_46776,N_46827);
or U47041 (N_47041,N_46916,N_46955);
and U47042 (N_47042,N_46924,N_46809);
or U47043 (N_47043,N_46927,N_46847);
nand U47044 (N_47044,N_46834,N_46784);
or U47045 (N_47045,N_46814,N_46973);
or U47046 (N_47046,N_46999,N_46936);
nand U47047 (N_47047,N_46983,N_46807);
nand U47048 (N_47048,N_46911,N_46939);
or U47049 (N_47049,N_46756,N_46871);
nand U47050 (N_47050,N_46958,N_46812);
and U47051 (N_47051,N_46887,N_46969);
nor U47052 (N_47052,N_46989,N_46956);
nor U47053 (N_47053,N_46901,N_46792);
nor U47054 (N_47054,N_46959,N_46801);
nand U47055 (N_47055,N_46942,N_46842);
nand U47056 (N_47056,N_46774,N_46908);
nand U47057 (N_47057,N_46874,N_46965);
and U47058 (N_47058,N_46800,N_46928);
or U47059 (N_47059,N_46751,N_46875);
nor U47060 (N_47060,N_46993,N_46949);
nor U47061 (N_47061,N_46891,N_46822);
and U47062 (N_47062,N_46910,N_46877);
or U47063 (N_47063,N_46994,N_46750);
or U47064 (N_47064,N_46948,N_46818);
nand U47065 (N_47065,N_46777,N_46868);
xnor U47066 (N_47066,N_46833,N_46878);
nor U47067 (N_47067,N_46797,N_46980);
and U47068 (N_47068,N_46918,N_46888);
nor U47069 (N_47069,N_46783,N_46781);
or U47070 (N_47070,N_46919,N_46892);
nand U47071 (N_47071,N_46925,N_46853);
and U47072 (N_47072,N_46986,N_46976);
or U47073 (N_47073,N_46904,N_46926);
xnor U47074 (N_47074,N_46922,N_46762);
and U47075 (N_47075,N_46977,N_46870);
and U47076 (N_47076,N_46838,N_46786);
nand U47077 (N_47077,N_46765,N_46941);
nor U47078 (N_47078,N_46836,N_46879);
nor U47079 (N_47079,N_46882,N_46851);
or U47080 (N_47080,N_46794,N_46760);
and U47081 (N_47081,N_46769,N_46996);
nor U47082 (N_47082,N_46857,N_46876);
or U47083 (N_47083,N_46899,N_46823);
and U47084 (N_47084,N_46953,N_46975);
and U47085 (N_47085,N_46808,N_46934);
nand U47086 (N_47086,N_46859,N_46831);
or U47087 (N_47087,N_46862,N_46839);
xnor U47088 (N_47088,N_46811,N_46772);
nand U47089 (N_47089,N_46914,N_46841);
xnor U47090 (N_47090,N_46761,N_46880);
nor U47091 (N_47091,N_46944,N_46974);
or U47092 (N_47092,N_46845,N_46824);
and U47093 (N_47093,N_46791,N_46984);
nand U47094 (N_47094,N_46938,N_46817);
nand U47095 (N_47095,N_46757,N_46806);
xor U47096 (N_47096,N_46883,N_46805);
nand U47097 (N_47097,N_46830,N_46819);
xor U47098 (N_47098,N_46864,N_46843);
and U47099 (N_47099,N_46825,N_46828);
xnor U47100 (N_47100,N_46835,N_46855);
nor U47101 (N_47101,N_46850,N_46768);
xor U47102 (N_47102,N_46981,N_46798);
nand U47103 (N_47103,N_46816,N_46796);
xor U47104 (N_47104,N_46962,N_46829);
and U47105 (N_47105,N_46933,N_46898);
and U47106 (N_47106,N_46873,N_46810);
or U47107 (N_47107,N_46771,N_46966);
or U47108 (N_47108,N_46998,N_46905);
and U47109 (N_47109,N_46759,N_46755);
nand U47110 (N_47110,N_46923,N_46790);
and U47111 (N_47111,N_46935,N_46954);
nand U47112 (N_47112,N_46913,N_46854);
and U47113 (N_47113,N_46937,N_46982);
nand U47114 (N_47114,N_46789,N_46764);
nor U47115 (N_47115,N_46997,N_46881);
and U47116 (N_47116,N_46753,N_46778);
nor U47117 (N_47117,N_46947,N_46991);
and U47118 (N_47118,N_46886,N_46909);
and U47119 (N_47119,N_46929,N_46890);
nand U47120 (N_47120,N_46985,N_46932);
and U47121 (N_47121,N_46968,N_46767);
and U47122 (N_47122,N_46763,N_46799);
or U47123 (N_47123,N_46902,N_46988);
nor U47124 (N_47124,N_46849,N_46780);
nand U47125 (N_47125,N_46922,N_46825);
or U47126 (N_47126,N_46881,N_46834);
nor U47127 (N_47127,N_46962,N_46890);
nor U47128 (N_47128,N_46872,N_46818);
nor U47129 (N_47129,N_46751,N_46913);
nor U47130 (N_47130,N_46851,N_46850);
and U47131 (N_47131,N_46960,N_46988);
xnor U47132 (N_47132,N_46994,N_46907);
and U47133 (N_47133,N_46857,N_46985);
nand U47134 (N_47134,N_46981,N_46915);
xor U47135 (N_47135,N_46804,N_46984);
and U47136 (N_47136,N_46866,N_46851);
nand U47137 (N_47137,N_46959,N_46910);
nor U47138 (N_47138,N_46854,N_46967);
and U47139 (N_47139,N_46948,N_46827);
nand U47140 (N_47140,N_46778,N_46829);
or U47141 (N_47141,N_46880,N_46788);
or U47142 (N_47142,N_46812,N_46905);
or U47143 (N_47143,N_46908,N_46922);
and U47144 (N_47144,N_46918,N_46895);
or U47145 (N_47145,N_46964,N_46887);
xor U47146 (N_47146,N_46969,N_46960);
nor U47147 (N_47147,N_46984,N_46839);
nor U47148 (N_47148,N_46961,N_46875);
nand U47149 (N_47149,N_46812,N_46781);
nand U47150 (N_47150,N_46986,N_46812);
nand U47151 (N_47151,N_46838,N_46845);
and U47152 (N_47152,N_46870,N_46826);
xor U47153 (N_47153,N_46856,N_46886);
xnor U47154 (N_47154,N_46964,N_46941);
nand U47155 (N_47155,N_46820,N_46756);
nand U47156 (N_47156,N_46979,N_46918);
nand U47157 (N_47157,N_46963,N_46935);
or U47158 (N_47158,N_46776,N_46811);
and U47159 (N_47159,N_46755,N_46951);
or U47160 (N_47160,N_46836,N_46782);
and U47161 (N_47161,N_46877,N_46890);
and U47162 (N_47162,N_46774,N_46967);
nor U47163 (N_47163,N_46976,N_46929);
and U47164 (N_47164,N_46877,N_46757);
xor U47165 (N_47165,N_46938,N_46795);
or U47166 (N_47166,N_46837,N_46911);
and U47167 (N_47167,N_46963,N_46842);
nand U47168 (N_47168,N_46797,N_46868);
or U47169 (N_47169,N_46835,N_46772);
or U47170 (N_47170,N_46905,N_46860);
nand U47171 (N_47171,N_46835,N_46839);
nand U47172 (N_47172,N_46930,N_46804);
xnor U47173 (N_47173,N_46860,N_46835);
xor U47174 (N_47174,N_46831,N_46801);
xnor U47175 (N_47175,N_46814,N_46981);
and U47176 (N_47176,N_46972,N_46821);
and U47177 (N_47177,N_46776,N_46952);
or U47178 (N_47178,N_46999,N_46903);
and U47179 (N_47179,N_46851,N_46890);
nand U47180 (N_47180,N_46967,N_46880);
or U47181 (N_47181,N_46846,N_46866);
or U47182 (N_47182,N_46900,N_46847);
nor U47183 (N_47183,N_46929,N_46785);
or U47184 (N_47184,N_46779,N_46951);
xor U47185 (N_47185,N_46800,N_46959);
nand U47186 (N_47186,N_46885,N_46917);
xor U47187 (N_47187,N_46770,N_46810);
or U47188 (N_47188,N_46990,N_46947);
nand U47189 (N_47189,N_46818,N_46947);
and U47190 (N_47190,N_46884,N_46780);
nor U47191 (N_47191,N_46887,N_46833);
and U47192 (N_47192,N_46985,N_46950);
and U47193 (N_47193,N_46796,N_46930);
or U47194 (N_47194,N_46972,N_46959);
xnor U47195 (N_47195,N_46830,N_46886);
nor U47196 (N_47196,N_46966,N_46820);
or U47197 (N_47197,N_46941,N_46875);
xor U47198 (N_47198,N_46770,N_46890);
xnor U47199 (N_47199,N_46957,N_46780);
nor U47200 (N_47200,N_46884,N_46799);
or U47201 (N_47201,N_46863,N_46918);
and U47202 (N_47202,N_46994,N_46911);
and U47203 (N_47203,N_46762,N_46880);
and U47204 (N_47204,N_46922,N_46917);
or U47205 (N_47205,N_46752,N_46961);
and U47206 (N_47206,N_46915,N_46956);
nor U47207 (N_47207,N_46779,N_46760);
nand U47208 (N_47208,N_46846,N_46892);
and U47209 (N_47209,N_46850,N_46991);
nand U47210 (N_47210,N_46786,N_46951);
nor U47211 (N_47211,N_46775,N_46866);
nand U47212 (N_47212,N_46803,N_46865);
and U47213 (N_47213,N_46799,N_46860);
and U47214 (N_47214,N_46925,N_46818);
xor U47215 (N_47215,N_46826,N_46921);
nand U47216 (N_47216,N_46818,N_46929);
xor U47217 (N_47217,N_46908,N_46814);
and U47218 (N_47218,N_46755,N_46989);
xnor U47219 (N_47219,N_46869,N_46863);
nand U47220 (N_47220,N_46941,N_46851);
nand U47221 (N_47221,N_46920,N_46750);
nor U47222 (N_47222,N_46823,N_46760);
xnor U47223 (N_47223,N_46791,N_46998);
xnor U47224 (N_47224,N_46973,N_46819);
and U47225 (N_47225,N_46873,N_46921);
or U47226 (N_47226,N_46884,N_46938);
nand U47227 (N_47227,N_46831,N_46993);
nand U47228 (N_47228,N_46754,N_46891);
and U47229 (N_47229,N_46929,N_46874);
nand U47230 (N_47230,N_46961,N_46777);
nor U47231 (N_47231,N_46779,N_46918);
and U47232 (N_47232,N_46915,N_46752);
nand U47233 (N_47233,N_46781,N_46989);
nor U47234 (N_47234,N_46881,N_46827);
nand U47235 (N_47235,N_46908,N_46800);
nand U47236 (N_47236,N_46765,N_46810);
or U47237 (N_47237,N_46958,N_46848);
or U47238 (N_47238,N_46939,N_46791);
and U47239 (N_47239,N_46909,N_46882);
or U47240 (N_47240,N_46996,N_46883);
and U47241 (N_47241,N_46798,N_46873);
or U47242 (N_47242,N_46891,N_46968);
or U47243 (N_47243,N_46923,N_46816);
and U47244 (N_47244,N_46964,N_46839);
and U47245 (N_47245,N_46905,N_46818);
or U47246 (N_47246,N_46877,N_46762);
nor U47247 (N_47247,N_46858,N_46902);
nand U47248 (N_47248,N_46824,N_46792);
nand U47249 (N_47249,N_46877,N_46838);
nand U47250 (N_47250,N_47158,N_47114);
xnor U47251 (N_47251,N_47004,N_47239);
nand U47252 (N_47252,N_47091,N_47058);
xor U47253 (N_47253,N_47174,N_47123);
nand U47254 (N_47254,N_47019,N_47104);
xnor U47255 (N_47255,N_47038,N_47115);
or U47256 (N_47256,N_47163,N_47106);
xor U47257 (N_47257,N_47110,N_47111);
nand U47258 (N_47258,N_47067,N_47092);
nor U47259 (N_47259,N_47017,N_47228);
xor U47260 (N_47260,N_47050,N_47015);
and U47261 (N_47261,N_47082,N_47087);
nand U47262 (N_47262,N_47006,N_47003);
xor U47263 (N_47263,N_47037,N_47047);
or U47264 (N_47264,N_47055,N_47241);
and U47265 (N_47265,N_47020,N_47211);
nand U47266 (N_47266,N_47154,N_47014);
nor U47267 (N_47267,N_47045,N_47200);
or U47268 (N_47268,N_47249,N_47031);
xor U47269 (N_47269,N_47233,N_47235);
and U47270 (N_47270,N_47005,N_47044);
and U47271 (N_47271,N_47032,N_47046);
nand U47272 (N_47272,N_47073,N_47121);
and U47273 (N_47273,N_47220,N_47053);
nand U47274 (N_47274,N_47130,N_47107);
and U47275 (N_47275,N_47160,N_47009);
xor U47276 (N_47276,N_47124,N_47223);
and U47277 (N_47277,N_47023,N_47170);
nand U47278 (N_47278,N_47247,N_47069);
nand U47279 (N_47279,N_47025,N_47093);
nor U47280 (N_47280,N_47139,N_47024);
nor U47281 (N_47281,N_47205,N_47065);
or U47282 (N_47282,N_47068,N_47159);
or U47283 (N_47283,N_47149,N_47076);
or U47284 (N_47284,N_47095,N_47101);
and U47285 (N_47285,N_47195,N_47216);
and U47286 (N_47286,N_47048,N_47193);
xnor U47287 (N_47287,N_47141,N_47077);
and U47288 (N_47288,N_47016,N_47248);
and U47289 (N_47289,N_47071,N_47183);
or U47290 (N_47290,N_47012,N_47081);
or U47291 (N_47291,N_47208,N_47140);
and U47292 (N_47292,N_47083,N_47178);
xnor U47293 (N_47293,N_47222,N_47175);
nor U47294 (N_47294,N_47052,N_47054);
xnor U47295 (N_47295,N_47134,N_47212);
and U47296 (N_47296,N_47144,N_47018);
nand U47297 (N_47297,N_47243,N_47180);
xnor U47298 (N_47298,N_47162,N_47242);
or U47299 (N_47299,N_47138,N_47225);
xor U47300 (N_47300,N_47105,N_47129);
or U47301 (N_47301,N_47039,N_47177);
xnor U47302 (N_47302,N_47244,N_47173);
or U47303 (N_47303,N_47030,N_47007);
nor U47304 (N_47304,N_47097,N_47185);
or U47305 (N_47305,N_47064,N_47150);
nand U47306 (N_47306,N_47066,N_47148);
or U47307 (N_47307,N_47232,N_47230);
nand U47308 (N_47308,N_47245,N_47062);
and U47309 (N_47309,N_47089,N_47119);
or U47310 (N_47310,N_47221,N_47181);
xnor U47311 (N_47311,N_47001,N_47215);
or U47312 (N_47312,N_47188,N_47164);
nor U47313 (N_47313,N_47147,N_47078);
nand U47314 (N_47314,N_47033,N_47204);
or U47315 (N_47315,N_47051,N_47132);
xnor U47316 (N_47316,N_47086,N_47227);
nand U47317 (N_47317,N_47098,N_47207);
nor U47318 (N_47318,N_47172,N_47197);
and U47319 (N_47319,N_47206,N_47157);
and U47320 (N_47320,N_47234,N_47099);
xnor U47321 (N_47321,N_47125,N_47190);
and U47322 (N_47322,N_47008,N_47063);
or U47323 (N_47323,N_47217,N_47152);
xor U47324 (N_47324,N_47128,N_47194);
nand U47325 (N_47325,N_47102,N_47126);
nand U47326 (N_47326,N_47237,N_47029);
nand U47327 (N_47327,N_47153,N_47040);
and U47328 (N_47328,N_47060,N_47100);
or U47329 (N_47329,N_47231,N_47010);
or U47330 (N_47330,N_47084,N_47072);
nand U47331 (N_47331,N_47198,N_47120);
or U47332 (N_47332,N_47219,N_47146);
and U47333 (N_47333,N_47187,N_47176);
xor U47334 (N_47334,N_47210,N_47041);
or U47335 (N_47335,N_47085,N_47182);
and U47336 (N_47336,N_47151,N_47034);
and U47337 (N_47337,N_47201,N_47203);
nand U47338 (N_47338,N_47113,N_47059);
or U47339 (N_47339,N_47116,N_47088);
nor U47340 (N_47340,N_47209,N_47061);
or U47341 (N_47341,N_47127,N_47156);
and U47342 (N_47342,N_47057,N_47202);
or U47343 (N_47343,N_47229,N_47192);
or U47344 (N_47344,N_47196,N_47168);
xnor U47345 (N_47345,N_47090,N_47191);
and U47346 (N_47346,N_47000,N_47079);
or U47347 (N_47347,N_47167,N_47117);
nor U47348 (N_47348,N_47075,N_47224);
xnor U47349 (N_47349,N_47145,N_47136);
nor U47350 (N_47350,N_47137,N_47246);
nor U47351 (N_47351,N_47035,N_47218);
and U47352 (N_47352,N_47142,N_47213);
nand U47353 (N_47353,N_47011,N_47056);
and U47354 (N_47354,N_47074,N_47143);
nor U47355 (N_47355,N_47043,N_47184);
nand U47356 (N_47356,N_47171,N_47042);
nor U47357 (N_47357,N_47021,N_47238);
nand U47358 (N_47358,N_47028,N_47135);
xor U47359 (N_47359,N_47013,N_47161);
nand U47360 (N_47360,N_47226,N_47049);
and U47361 (N_47361,N_47169,N_47179);
xnor U47362 (N_47362,N_47080,N_47103);
and U47363 (N_47363,N_47165,N_47036);
and U47364 (N_47364,N_47199,N_47002);
and U47365 (N_47365,N_47236,N_47109);
or U47366 (N_47366,N_47214,N_47027);
xnor U47367 (N_47367,N_47131,N_47133);
nor U47368 (N_47368,N_47186,N_47108);
nor U47369 (N_47369,N_47094,N_47240);
or U47370 (N_47370,N_47166,N_47118);
xnor U47371 (N_47371,N_47189,N_47122);
xnor U47372 (N_47372,N_47022,N_47096);
nor U47373 (N_47373,N_47026,N_47070);
or U47374 (N_47374,N_47155,N_47112);
xor U47375 (N_47375,N_47062,N_47137);
xor U47376 (N_47376,N_47063,N_47086);
and U47377 (N_47377,N_47240,N_47163);
xor U47378 (N_47378,N_47109,N_47124);
and U47379 (N_47379,N_47132,N_47168);
xnor U47380 (N_47380,N_47214,N_47129);
xnor U47381 (N_47381,N_47163,N_47227);
or U47382 (N_47382,N_47035,N_47107);
nand U47383 (N_47383,N_47115,N_47117);
nand U47384 (N_47384,N_47122,N_47214);
xor U47385 (N_47385,N_47085,N_47148);
and U47386 (N_47386,N_47067,N_47220);
or U47387 (N_47387,N_47218,N_47127);
xnor U47388 (N_47388,N_47066,N_47073);
xor U47389 (N_47389,N_47015,N_47144);
nand U47390 (N_47390,N_47139,N_47147);
and U47391 (N_47391,N_47012,N_47247);
nand U47392 (N_47392,N_47181,N_47131);
xnor U47393 (N_47393,N_47220,N_47011);
nor U47394 (N_47394,N_47077,N_47027);
nor U47395 (N_47395,N_47000,N_47083);
nand U47396 (N_47396,N_47179,N_47144);
nor U47397 (N_47397,N_47099,N_47018);
nor U47398 (N_47398,N_47178,N_47102);
nand U47399 (N_47399,N_47034,N_47006);
nor U47400 (N_47400,N_47014,N_47007);
or U47401 (N_47401,N_47151,N_47026);
xor U47402 (N_47402,N_47127,N_47144);
nor U47403 (N_47403,N_47234,N_47081);
and U47404 (N_47404,N_47033,N_47227);
xnor U47405 (N_47405,N_47177,N_47249);
and U47406 (N_47406,N_47092,N_47125);
and U47407 (N_47407,N_47087,N_47237);
nor U47408 (N_47408,N_47023,N_47059);
nand U47409 (N_47409,N_47185,N_47002);
and U47410 (N_47410,N_47177,N_47024);
and U47411 (N_47411,N_47013,N_47154);
and U47412 (N_47412,N_47061,N_47225);
and U47413 (N_47413,N_47142,N_47216);
or U47414 (N_47414,N_47020,N_47066);
or U47415 (N_47415,N_47246,N_47168);
and U47416 (N_47416,N_47060,N_47049);
or U47417 (N_47417,N_47000,N_47032);
nor U47418 (N_47418,N_47048,N_47203);
or U47419 (N_47419,N_47079,N_47173);
and U47420 (N_47420,N_47147,N_47035);
and U47421 (N_47421,N_47122,N_47156);
nand U47422 (N_47422,N_47071,N_47236);
and U47423 (N_47423,N_47111,N_47034);
nor U47424 (N_47424,N_47238,N_47239);
or U47425 (N_47425,N_47067,N_47098);
xnor U47426 (N_47426,N_47025,N_47148);
and U47427 (N_47427,N_47188,N_47111);
and U47428 (N_47428,N_47123,N_47204);
xnor U47429 (N_47429,N_47007,N_47156);
nor U47430 (N_47430,N_47026,N_47073);
nand U47431 (N_47431,N_47243,N_47069);
nand U47432 (N_47432,N_47092,N_47152);
or U47433 (N_47433,N_47078,N_47196);
or U47434 (N_47434,N_47245,N_47037);
nand U47435 (N_47435,N_47173,N_47069);
nand U47436 (N_47436,N_47076,N_47197);
and U47437 (N_47437,N_47119,N_47128);
nand U47438 (N_47438,N_47155,N_47197);
or U47439 (N_47439,N_47107,N_47125);
or U47440 (N_47440,N_47218,N_47040);
xnor U47441 (N_47441,N_47125,N_47071);
xnor U47442 (N_47442,N_47048,N_47162);
nor U47443 (N_47443,N_47043,N_47034);
nand U47444 (N_47444,N_47059,N_47095);
nor U47445 (N_47445,N_47173,N_47141);
nor U47446 (N_47446,N_47059,N_47186);
or U47447 (N_47447,N_47055,N_47116);
nand U47448 (N_47448,N_47092,N_47186);
or U47449 (N_47449,N_47246,N_47227);
nand U47450 (N_47450,N_47002,N_47009);
or U47451 (N_47451,N_47133,N_47053);
nor U47452 (N_47452,N_47131,N_47149);
nand U47453 (N_47453,N_47013,N_47228);
nor U47454 (N_47454,N_47001,N_47074);
nand U47455 (N_47455,N_47138,N_47183);
nand U47456 (N_47456,N_47088,N_47205);
or U47457 (N_47457,N_47105,N_47113);
nand U47458 (N_47458,N_47010,N_47088);
or U47459 (N_47459,N_47018,N_47200);
nand U47460 (N_47460,N_47027,N_47024);
nand U47461 (N_47461,N_47080,N_47097);
or U47462 (N_47462,N_47205,N_47011);
and U47463 (N_47463,N_47160,N_47249);
or U47464 (N_47464,N_47179,N_47167);
xor U47465 (N_47465,N_47112,N_47177);
or U47466 (N_47466,N_47128,N_47070);
nand U47467 (N_47467,N_47039,N_47020);
nand U47468 (N_47468,N_47208,N_47088);
nand U47469 (N_47469,N_47242,N_47249);
xnor U47470 (N_47470,N_47176,N_47241);
xor U47471 (N_47471,N_47013,N_47084);
and U47472 (N_47472,N_47210,N_47156);
nor U47473 (N_47473,N_47036,N_47135);
nand U47474 (N_47474,N_47246,N_47108);
xnor U47475 (N_47475,N_47062,N_47215);
and U47476 (N_47476,N_47160,N_47193);
nor U47477 (N_47477,N_47004,N_47097);
xnor U47478 (N_47478,N_47060,N_47235);
nand U47479 (N_47479,N_47157,N_47093);
nand U47480 (N_47480,N_47185,N_47071);
nor U47481 (N_47481,N_47144,N_47055);
or U47482 (N_47482,N_47217,N_47179);
xnor U47483 (N_47483,N_47016,N_47120);
nand U47484 (N_47484,N_47003,N_47068);
and U47485 (N_47485,N_47202,N_47006);
or U47486 (N_47486,N_47223,N_47181);
nand U47487 (N_47487,N_47183,N_47217);
nor U47488 (N_47488,N_47057,N_47109);
nor U47489 (N_47489,N_47107,N_47044);
xnor U47490 (N_47490,N_47074,N_47168);
nand U47491 (N_47491,N_47154,N_47038);
nand U47492 (N_47492,N_47166,N_47143);
nand U47493 (N_47493,N_47164,N_47224);
nor U47494 (N_47494,N_47051,N_47243);
and U47495 (N_47495,N_47148,N_47110);
xor U47496 (N_47496,N_47074,N_47157);
or U47497 (N_47497,N_47157,N_47048);
and U47498 (N_47498,N_47058,N_47046);
nand U47499 (N_47499,N_47240,N_47246);
nor U47500 (N_47500,N_47288,N_47280);
xnor U47501 (N_47501,N_47393,N_47366);
nor U47502 (N_47502,N_47303,N_47416);
or U47503 (N_47503,N_47267,N_47474);
and U47504 (N_47504,N_47478,N_47386);
or U47505 (N_47505,N_47256,N_47375);
xnor U47506 (N_47506,N_47401,N_47379);
xnor U47507 (N_47507,N_47335,N_47314);
and U47508 (N_47508,N_47261,N_47396);
and U47509 (N_47509,N_47454,N_47458);
and U47510 (N_47510,N_47345,N_47272);
and U47511 (N_47511,N_47462,N_47355);
nand U47512 (N_47512,N_47490,N_47499);
nor U47513 (N_47513,N_47285,N_47425);
nand U47514 (N_47514,N_47481,N_47340);
or U47515 (N_47515,N_47449,N_47299);
or U47516 (N_47516,N_47262,N_47313);
and U47517 (N_47517,N_47381,N_47459);
nand U47518 (N_47518,N_47463,N_47252);
xnor U47519 (N_47519,N_47258,N_47259);
nand U47520 (N_47520,N_47287,N_47333);
or U47521 (N_47521,N_47435,N_47403);
and U47522 (N_47522,N_47266,N_47385);
nor U47523 (N_47523,N_47325,N_47376);
and U47524 (N_47524,N_47482,N_47358);
xor U47525 (N_47525,N_47440,N_47384);
xor U47526 (N_47526,N_47337,N_47297);
nor U47527 (N_47527,N_47467,N_47476);
and U47528 (N_47528,N_47405,N_47457);
xnor U47529 (N_47529,N_47455,N_47432);
xor U47530 (N_47530,N_47319,N_47364);
nand U47531 (N_47531,N_47307,N_47309);
nor U47532 (N_47532,N_47293,N_47341);
nor U47533 (N_47533,N_47485,N_47330);
xnor U47534 (N_47534,N_47468,N_47360);
and U47535 (N_47535,N_47268,N_47399);
nor U47536 (N_47536,N_47343,N_47278);
nand U47537 (N_47537,N_47413,N_47354);
or U47538 (N_47538,N_47269,N_47357);
and U47539 (N_47539,N_47332,N_47370);
xnor U47540 (N_47540,N_47257,N_47483);
and U47541 (N_47541,N_47250,N_47441);
xnor U47542 (N_47542,N_47423,N_47368);
xnor U47543 (N_47543,N_47361,N_47327);
or U47544 (N_47544,N_47494,N_47447);
nand U47545 (N_47545,N_47450,N_47390);
nand U47546 (N_47546,N_47469,N_47484);
nand U47547 (N_47547,N_47373,N_47424);
or U47548 (N_47548,N_47452,N_47426);
nand U47549 (N_47549,N_47349,N_47437);
and U47550 (N_47550,N_47328,N_47398);
and U47551 (N_47551,N_47265,N_47400);
nor U47552 (N_47552,N_47419,N_47260);
or U47553 (N_47553,N_47312,N_47318);
nor U47554 (N_47554,N_47428,N_47316);
nand U47555 (N_47555,N_47417,N_47442);
and U47556 (N_47556,N_47279,N_47443);
xnor U47557 (N_47557,N_47298,N_47470);
nor U47558 (N_47558,N_47274,N_47444);
nand U47559 (N_47559,N_47394,N_47404);
nand U47560 (N_47560,N_47479,N_47277);
and U47561 (N_47561,N_47276,N_47480);
xnor U47562 (N_47562,N_47290,N_47430);
and U47563 (N_47563,N_47323,N_47451);
and U47564 (N_47564,N_47387,N_47397);
xnor U47565 (N_47565,N_47477,N_47475);
xnor U47566 (N_47566,N_47353,N_47270);
xor U47567 (N_47567,N_47295,N_47466);
or U47568 (N_47568,N_47310,N_47365);
nand U47569 (N_47569,N_47411,N_47326);
xnor U47570 (N_47570,N_47383,N_47292);
nand U47571 (N_47571,N_47306,N_47301);
xnor U47572 (N_47572,N_47329,N_47492);
nor U47573 (N_47573,N_47334,N_47429);
or U47574 (N_47574,N_47291,N_47495);
nand U47575 (N_47575,N_47286,N_47308);
nand U47576 (N_47576,N_47346,N_47374);
or U47577 (N_47577,N_47251,N_47324);
nand U47578 (N_47578,N_47351,N_47336);
or U47579 (N_47579,N_47471,N_47254);
nand U47580 (N_47580,N_47439,N_47322);
or U47581 (N_47581,N_47282,N_47320);
and U47582 (N_47582,N_47497,N_47392);
nor U47583 (N_47583,N_47431,N_47421);
nor U47584 (N_47584,N_47407,N_47275);
and U47585 (N_47585,N_47377,N_47409);
xnor U47586 (N_47586,N_47253,N_47294);
and U47587 (N_47587,N_47255,N_47460);
xnor U47588 (N_47588,N_47498,N_47342);
xnor U47589 (N_47589,N_47388,N_47412);
xnor U47590 (N_47590,N_47402,N_47296);
nor U47591 (N_47591,N_47491,N_47311);
nor U47592 (N_47592,N_47264,N_47473);
nand U47593 (N_47593,N_47415,N_47453);
nor U47594 (N_47594,N_47446,N_47422);
or U47595 (N_47595,N_47317,N_47359);
xor U47596 (N_47596,N_47378,N_47367);
nor U47597 (N_47597,N_47356,N_47363);
and U47598 (N_47598,N_47281,N_47461);
nor U47599 (N_47599,N_47371,N_47321);
nand U47600 (N_47600,N_47420,N_47486);
nor U47601 (N_47601,N_47300,N_47283);
nand U47602 (N_47602,N_47418,N_47408);
or U47603 (N_47603,N_47284,N_47464);
xnor U47604 (N_47604,N_47339,N_47391);
xor U47605 (N_47605,N_47434,N_47348);
and U47606 (N_47606,N_47489,N_47271);
and U47607 (N_47607,N_47315,N_47433);
and U47608 (N_47608,N_47338,N_47436);
xnor U47609 (N_47609,N_47302,N_47472);
nor U47610 (N_47610,N_47427,N_47488);
xnor U47611 (N_47611,N_47350,N_47493);
xnor U47612 (N_47612,N_47331,N_47362);
nor U47613 (N_47613,N_47352,N_47263);
nor U47614 (N_47614,N_47406,N_47305);
xor U47615 (N_47615,N_47465,N_47344);
or U47616 (N_47616,N_47410,N_47414);
nand U47617 (N_47617,N_47389,N_47289);
or U47618 (N_47618,N_47438,N_47456);
nor U47619 (N_47619,N_47347,N_47496);
or U47620 (N_47620,N_47487,N_47445);
nor U47621 (N_47621,N_47395,N_47372);
and U47622 (N_47622,N_47382,N_47448);
and U47623 (N_47623,N_47304,N_47273);
xnor U47624 (N_47624,N_47380,N_47369);
or U47625 (N_47625,N_47398,N_47442);
and U47626 (N_47626,N_47428,N_47487);
xnor U47627 (N_47627,N_47263,N_47422);
or U47628 (N_47628,N_47323,N_47380);
and U47629 (N_47629,N_47276,N_47302);
and U47630 (N_47630,N_47368,N_47303);
xor U47631 (N_47631,N_47422,N_47498);
xnor U47632 (N_47632,N_47418,N_47417);
nand U47633 (N_47633,N_47447,N_47361);
or U47634 (N_47634,N_47305,N_47345);
nor U47635 (N_47635,N_47356,N_47492);
xor U47636 (N_47636,N_47373,N_47264);
or U47637 (N_47637,N_47462,N_47409);
nor U47638 (N_47638,N_47448,N_47336);
xnor U47639 (N_47639,N_47432,N_47482);
and U47640 (N_47640,N_47488,N_47298);
or U47641 (N_47641,N_47302,N_47327);
nand U47642 (N_47642,N_47372,N_47362);
nor U47643 (N_47643,N_47478,N_47318);
nor U47644 (N_47644,N_47352,N_47265);
nand U47645 (N_47645,N_47373,N_47451);
nand U47646 (N_47646,N_47369,N_47274);
xor U47647 (N_47647,N_47377,N_47359);
xnor U47648 (N_47648,N_47481,N_47372);
and U47649 (N_47649,N_47289,N_47326);
nor U47650 (N_47650,N_47268,N_47458);
nor U47651 (N_47651,N_47326,N_47256);
xnor U47652 (N_47652,N_47309,N_47485);
or U47653 (N_47653,N_47371,N_47473);
nand U47654 (N_47654,N_47426,N_47472);
nand U47655 (N_47655,N_47395,N_47488);
or U47656 (N_47656,N_47440,N_47368);
or U47657 (N_47657,N_47424,N_47415);
or U47658 (N_47658,N_47435,N_47485);
nand U47659 (N_47659,N_47406,N_47328);
xnor U47660 (N_47660,N_47307,N_47384);
nand U47661 (N_47661,N_47493,N_47272);
or U47662 (N_47662,N_47442,N_47499);
xor U47663 (N_47663,N_47357,N_47453);
xor U47664 (N_47664,N_47280,N_47390);
and U47665 (N_47665,N_47361,N_47330);
nor U47666 (N_47666,N_47430,N_47295);
nor U47667 (N_47667,N_47386,N_47438);
nand U47668 (N_47668,N_47434,N_47324);
xor U47669 (N_47669,N_47451,N_47474);
xnor U47670 (N_47670,N_47484,N_47411);
or U47671 (N_47671,N_47425,N_47461);
or U47672 (N_47672,N_47498,N_47282);
or U47673 (N_47673,N_47442,N_47377);
or U47674 (N_47674,N_47357,N_47420);
nor U47675 (N_47675,N_47432,N_47291);
nor U47676 (N_47676,N_47411,N_47364);
or U47677 (N_47677,N_47301,N_47361);
and U47678 (N_47678,N_47489,N_47474);
nand U47679 (N_47679,N_47443,N_47252);
or U47680 (N_47680,N_47353,N_47482);
or U47681 (N_47681,N_47305,N_47485);
and U47682 (N_47682,N_47330,N_47411);
or U47683 (N_47683,N_47472,N_47263);
nor U47684 (N_47684,N_47385,N_47435);
and U47685 (N_47685,N_47347,N_47257);
xor U47686 (N_47686,N_47419,N_47472);
nor U47687 (N_47687,N_47458,N_47411);
xnor U47688 (N_47688,N_47402,N_47450);
and U47689 (N_47689,N_47263,N_47446);
and U47690 (N_47690,N_47441,N_47431);
nand U47691 (N_47691,N_47478,N_47371);
or U47692 (N_47692,N_47443,N_47259);
and U47693 (N_47693,N_47325,N_47420);
or U47694 (N_47694,N_47420,N_47467);
and U47695 (N_47695,N_47324,N_47301);
nor U47696 (N_47696,N_47463,N_47374);
and U47697 (N_47697,N_47257,N_47302);
and U47698 (N_47698,N_47399,N_47323);
and U47699 (N_47699,N_47252,N_47308);
and U47700 (N_47700,N_47476,N_47340);
nand U47701 (N_47701,N_47482,N_47294);
or U47702 (N_47702,N_47314,N_47358);
nor U47703 (N_47703,N_47390,N_47330);
xnor U47704 (N_47704,N_47264,N_47319);
nor U47705 (N_47705,N_47464,N_47339);
nor U47706 (N_47706,N_47383,N_47486);
or U47707 (N_47707,N_47371,N_47320);
and U47708 (N_47708,N_47250,N_47340);
xor U47709 (N_47709,N_47454,N_47361);
xnor U47710 (N_47710,N_47364,N_47437);
xor U47711 (N_47711,N_47418,N_47290);
nand U47712 (N_47712,N_47451,N_47362);
nor U47713 (N_47713,N_47425,N_47256);
and U47714 (N_47714,N_47417,N_47289);
or U47715 (N_47715,N_47277,N_47385);
xnor U47716 (N_47716,N_47311,N_47383);
nor U47717 (N_47717,N_47375,N_47462);
and U47718 (N_47718,N_47441,N_47493);
xor U47719 (N_47719,N_47340,N_47338);
and U47720 (N_47720,N_47321,N_47398);
and U47721 (N_47721,N_47424,N_47402);
nor U47722 (N_47722,N_47380,N_47435);
nand U47723 (N_47723,N_47338,N_47269);
or U47724 (N_47724,N_47496,N_47251);
and U47725 (N_47725,N_47356,N_47413);
xor U47726 (N_47726,N_47410,N_47473);
or U47727 (N_47727,N_47463,N_47262);
nand U47728 (N_47728,N_47473,N_47317);
or U47729 (N_47729,N_47328,N_47494);
or U47730 (N_47730,N_47392,N_47371);
and U47731 (N_47731,N_47495,N_47316);
xnor U47732 (N_47732,N_47353,N_47379);
nand U47733 (N_47733,N_47325,N_47453);
nor U47734 (N_47734,N_47310,N_47374);
xor U47735 (N_47735,N_47433,N_47399);
or U47736 (N_47736,N_47432,N_47386);
nand U47737 (N_47737,N_47479,N_47493);
or U47738 (N_47738,N_47308,N_47362);
xor U47739 (N_47739,N_47318,N_47316);
nand U47740 (N_47740,N_47287,N_47274);
or U47741 (N_47741,N_47328,N_47471);
nand U47742 (N_47742,N_47444,N_47496);
and U47743 (N_47743,N_47262,N_47267);
xnor U47744 (N_47744,N_47260,N_47302);
nor U47745 (N_47745,N_47278,N_47432);
or U47746 (N_47746,N_47475,N_47350);
nand U47747 (N_47747,N_47295,N_47391);
nor U47748 (N_47748,N_47479,N_47386);
xnor U47749 (N_47749,N_47265,N_47393);
xor U47750 (N_47750,N_47686,N_47671);
nand U47751 (N_47751,N_47589,N_47599);
xor U47752 (N_47752,N_47684,N_47534);
and U47753 (N_47753,N_47695,N_47632);
or U47754 (N_47754,N_47722,N_47731);
xor U47755 (N_47755,N_47736,N_47724);
nor U47756 (N_47756,N_47652,N_47634);
xnor U47757 (N_47757,N_47604,N_47714);
and U47758 (N_47758,N_47537,N_47526);
nor U47759 (N_47759,N_47542,N_47651);
xor U47760 (N_47760,N_47590,N_47616);
nand U47761 (N_47761,N_47546,N_47533);
nand U47762 (N_47762,N_47527,N_47554);
xor U47763 (N_47763,N_47568,N_47726);
nor U47764 (N_47764,N_47563,N_47561);
nor U47765 (N_47765,N_47524,N_47569);
nand U47766 (N_47766,N_47596,N_47612);
or U47767 (N_47767,N_47518,N_47566);
xnor U47768 (N_47768,N_47531,N_47707);
xnor U47769 (N_47769,N_47580,N_47683);
and U47770 (N_47770,N_47633,N_47739);
or U47771 (N_47771,N_47532,N_47575);
or U47772 (N_47772,N_47510,N_47548);
and U47773 (N_47773,N_47625,N_47549);
or U47774 (N_47774,N_47574,N_47509);
nand U47775 (N_47775,N_47647,N_47728);
nand U47776 (N_47776,N_47661,N_47617);
nor U47777 (N_47777,N_47703,N_47620);
nor U47778 (N_47778,N_47700,N_47582);
nand U47779 (N_47779,N_47595,N_47658);
or U47780 (N_47780,N_47730,N_47729);
xnor U47781 (N_47781,N_47501,N_47545);
and U47782 (N_47782,N_47565,N_47511);
and U47783 (N_47783,N_47734,N_47667);
or U47784 (N_47784,N_47522,N_47613);
or U47785 (N_47785,N_47649,N_47610);
or U47786 (N_47786,N_47637,N_47701);
or U47787 (N_47787,N_47740,N_47699);
xor U47788 (N_47788,N_47540,N_47747);
xnor U47789 (N_47789,N_47648,N_47529);
nor U47790 (N_47790,N_47578,N_47696);
or U47791 (N_47791,N_47626,N_47675);
nand U47792 (N_47792,N_47680,N_47682);
and U47793 (N_47793,N_47668,N_47502);
and U47794 (N_47794,N_47678,N_47743);
nor U47795 (N_47795,N_47603,N_47664);
or U47796 (N_47796,N_47636,N_47641);
or U47797 (N_47797,N_47601,N_47706);
and U47798 (N_47798,N_47660,N_47716);
nand U47799 (N_47799,N_47521,N_47689);
or U47800 (N_47800,N_47583,N_47516);
and U47801 (N_47801,N_47619,N_47577);
xnor U47802 (N_47802,N_47640,N_47579);
nor U47803 (N_47803,N_47674,N_47515);
xnor U47804 (N_47804,N_47666,N_47588);
or U47805 (N_47805,N_47639,N_47506);
nand U47806 (N_47806,N_47523,N_47607);
nand U47807 (N_47807,N_47500,N_47547);
nor U47808 (N_47808,N_47744,N_47525);
or U47809 (N_47809,N_47646,N_47720);
xor U47810 (N_47810,N_47705,N_47552);
xnor U47811 (N_47811,N_47503,N_47642);
nand U47812 (N_47812,N_47713,N_47572);
and U47813 (N_47813,N_47517,N_47587);
nor U47814 (N_47814,N_47550,N_47662);
nand U47815 (N_47815,N_47687,N_47621);
xor U47816 (N_47816,N_47741,N_47555);
nand U47817 (N_47817,N_47514,N_47638);
or U47818 (N_47818,N_47654,N_47738);
xor U47819 (N_47819,N_47602,N_47544);
and U47820 (N_47820,N_47663,N_47535);
and U47821 (N_47821,N_47645,N_47742);
nand U47822 (N_47822,N_47560,N_47657);
and U47823 (N_47823,N_47543,N_47553);
xnor U47824 (N_47824,N_47507,N_47672);
nand U47825 (N_47825,N_47623,N_47598);
nor U47826 (N_47826,N_47593,N_47712);
nand U47827 (N_47827,N_47592,N_47624);
nand U47828 (N_47828,N_47591,N_47581);
nor U47829 (N_47829,N_47690,N_47570);
nand U47830 (N_47830,N_47618,N_47615);
nand U47831 (N_47831,N_47673,N_47732);
nor U47832 (N_47832,N_47677,N_47528);
and U47833 (N_47833,N_47656,N_47622);
xor U47834 (N_47834,N_47562,N_47559);
or U47835 (N_47835,N_47557,N_47611);
and U47836 (N_47836,N_47505,N_47571);
or U47837 (N_47837,N_47586,N_47608);
nor U47838 (N_47838,N_47558,N_47693);
or U47839 (N_47839,N_47504,N_47573);
nand U47840 (N_47840,N_47606,N_47691);
and U47841 (N_47841,N_47512,N_47698);
and U47842 (N_47842,N_47685,N_47745);
nor U47843 (N_47843,N_47669,N_47508);
and U47844 (N_47844,N_47564,N_47541);
xor U47845 (N_47845,N_47718,N_47717);
or U47846 (N_47846,N_47727,N_47635);
xnor U47847 (N_47847,N_47600,N_47688);
xor U47848 (N_47848,N_47629,N_47567);
nand U47849 (N_47849,N_47530,N_47708);
and U47850 (N_47850,N_47721,N_47536);
nand U47851 (N_47851,N_47735,N_47584);
and U47852 (N_47852,N_47692,N_47715);
or U47853 (N_47853,N_47733,N_47679);
nand U47854 (N_47854,N_47538,N_47520);
or U47855 (N_47855,N_47709,N_47594);
and U47856 (N_47856,N_47676,N_47631);
xor U47857 (N_47857,N_47723,N_47704);
nor U47858 (N_47858,N_47609,N_47653);
and U47859 (N_47859,N_47585,N_47539);
or U47860 (N_47860,N_47519,N_47725);
or U47861 (N_47861,N_47710,N_47737);
nor U47862 (N_47862,N_47628,N_47665);
and U47863 (N_47863,N_47670,N_47597);
and U47864 (N_47864,N_47719,N_47749);
nor U47865 (N_47865,N_47643,N_47650);
nand U47866 (N_47866,N_47644,N_47614);
and U47867 (N_47867,N_47627,N_47697);
nand U47868 (N_47868,N_47556,N_47655);
nor U47869 (N_47869,N_47694,N_47605);
or U47870 (N_47870,N_47746,N_47576);
and U47871 (N_47871,N_47711,N_47702);
or U47872 (N_47872,N_47513,N_47748);
and U47873 (N_47873,N_47551,N_47681);
or U47874 (N_47874,N_47630,N_47659);
nand U47875 (N_47875,N_47679,N_47595);
nand U47876 (N_47876,N_47724,N_47502);
xor U47877 (N_47877,N_47711,N_47696);
nand U47878 (N_47878,N_47505,N_47738);
nor U47879 (N_47879,N_47531,N_47516);
or U47880 (N_47880,N_47527,N_47524);
or U47881 (N_47881,N_47739,N_47695);
and U47882 (N_47882,N_47749,N_47627);
xor U47883 (N_47883,N_47562,N_47557);
or U47884 (N_47884,N_47626,N_47733);
nor U47885 (N_47885,N_47711,N_47568);
and U47886 (N_47886,N_47677,N_47712);
nand U47887 (N_47887,N_47639,N_47547);
nor U47888 (N_47888,N_47697,N_47669);
nand U47889 (N_47889,N_47680,N_47541);
or U47890 (N_47890,N_47528,N_47711);
and U47891 (N_47891,N_47539,N_47596);
nand U47892 (N_47892,N_47517,N_47582);
nand U47893 (N_47893,N_47701,N_47521);
and U47894 (N_47894,N_47599,N_47702);
and U47895 (N_47895,N_47675,N_47594);
nor U47896 (N_47896,N_47542,N_47599);
nand U47897 (N_47897,N_47586,N_47518);
nand U47898 (N_47898,N_47723,N_47677);
and U47899 (N_47899,N_47590,N_47660);
and U47900 (N_47900,N_47660,N_47546);
nand U47901 (N_47901,N_47510,N_47691);
or U47902 (N_47902,N_47590,N_47567);
xor U47903 (N_47903,N_47738,N_47658);
and U47904 (N_47904,N_47594,N_47723);
and U47905 (N_47905,N_47546,N_47707);
xnor U47906 (N_47906,N_47573,N_47732);
and U47907 (N_47907,N_47594,N_47603);
or U47908 (N_47908,N_47698,N_47619);
xor U47909 (N_47909,N_47598,N_47505);
nor U47910 (N_47910,N_47571,N_47590);
nor U47911 (N_47911,N_47692,N_47675);
and U47912 (N_47912,N_47628,N_47500);
nand U47913 (N_47913,N_47529,N_47571);
nor U47914 (N_47914,N_47542,N_47634);
xor U47915 (N_47915,N_47594,N_47543);
and U47916 (N_47916,N_47593,N_47541);
nor U47917 (N_47917,N_47728,N_47729);
or U47918 (N_47918,N_47639,N_47576);
or U47919 (N_47919,N_47586,N_47723);
or U47920 (N_47920,N_47538,N_47726);
or U47921 (N_47921,N_47681,N_47748);
and U47922 (N_47922,N_47533,N_47720);
nor U47923 (N_47923,N_47704,N_47603);
and U47924 (N_47924,N_47601,N_47737);
nand U47925 (N_47925,N_47705,N_47513);
or U47926 (N_47926,N_47618,N_47671);
nor U47927 (N_47927,N_47680,N_47589);
nor U47928 (N_47928,N_47712,N_47610);
nand U47929 (N_47929,N_47631,N_47501);
xor U47930 (N_47930,N_47502,N_47660);
xnor U47931 (N_47931,N_47638,N_47694);
xnor U47932 (N_47932,N_47740,N_47640);
or U47933 (N_47933,N_47687,N_47724);
or U47934 (N_47934,N_47590,N_47545);
nor U47935 (N_47935,N_47679,N_47635);
nand U47936 (N_47936,N_47620,N_47727);
nor U47937 (N_47937,N_47720,N_47555);
or U47938 (N_47938,N_47631,N_47664);
and U47939 (N_47939,N_47658,N_47741);
nor U47940 (N_47940,N_47740,N_47513);
and U47941 (N_47941,N_47675,N_47558);
nand U47942 (N_47942,N_47528,N_47661);
nor U47943 (N_47943,N_47737,N_47529);
and U47944 (N_47944,N_47519,N_47718);
xnor U47945 (N_47945,N_47610,N_47605);
xnor U47946 (N_47946,N_47520,N_47544);
nor U47947 (N_47947,N_47699,N_47688);
nor U47948 (N_47948,N_47651,N_47635);
xor U47949 (N_47949,N_47725,N_47711);
nand U47950 (N_47950,N_47636,N_47612);
nor U47951 (N_47951,N_47573,N_47634);
xor U47952 (N_47952,N_47601,N_47594);
xnor U47953 (N_47953,N_47581,N_47675);
xor U47954 (N_47954,N_47652,N_47661);
nor U47955 (N_47955,N_47526,N_47538);
xor U47956 (N_47956,N_47544,N_47578);
xnor U47957 (N_47957,N_47530,N_47532);
xor U47958 (N_47958,N_47724,N_47526);
xnor U47959 (N_47959,N_47651,N_47636);
and U47960 (N_47960,N_47624,N_47746);
xnor U47961 (N_47961,N_47561,N_47552);
xor U47962 (N_47962,N_47527,N_47513);
nor U47963 (N_47963,N_47700,N_47529);
and U47964 (N_47964,N_47508,N_47623);
or U47965 (N_47965,N_47721,N_47632);
or U47966 (N_47966,N_47573,N_47737);
nand U47967 (N_47967,N_47631,N_47738);
and U47968 (N_47968,N_47633,N_47563);
and U47969 (N_47969,N_47691,N_47592);
nor U47970 (N_47970,N_47601,N_47739);
xnor U47971 (N_47971,N_47742,N_47587);
and U47972 (N_47972,N_47654,N_47741);
or U47973 (N_47973,N_47735,N_47616);
nor U47974 (N_47974,N_47639,N_47525);
or U47975 (N_47975,N_47625,N_47621);
and U47976 (N_47976,N_47698,N_47517);
nand U47977 (N_47977,N_47527,N_47548);
or U47978 (N_47978,N_47564,N_47619);
nor U47979 (N_47979,N_47524,N_47639);
nor U47980 (N_47980,N_47593,N_47642);
xor U47981 (N_47981,N_47745,N_47582);
xnor U47982 (N_47982,N_47686,N_47745);
or U47983 (N_47983,N_47672,N_47630);
nand U47984 (N_47984,N_47523,N_47717);
nor U47985 (N_47985,N_47660,N_47558);
or U47986 (N_47986,N_47549,N_47622);
or U47987 (N_47987,N_47749,N_47610);
and U47988 (N_47988,N_47724,N_47537);
nand U47989 (N_47989,N_47539,N_47623);
xor U47990 (N_47990,N_47681,N_47626);
xnor U47991 (N_47991,N_47536,N_47742);
and U47992 (N_47992,N_47687,N_47727);
xnor U47993 (N_47993,N_47609,N_47606);
nand U47994 (N_47994,N_47581,N_47654);
nand U47995 (N_47995,N_47528,N_47607);
nor U47996 (N_47996,N_47705,N_47627);
nor U47997 (N_47997,N_47547,N_47652);
and U47998 (N_47998,N_47524,N_47588);
nand U47999 (N_47999,N_47725,N_47721);
and U48000 (N_48000,N_47885,N_47963);
nand U48001 (N_48001,N_47896,N_47916);
nor U48002 (N_48002,N_47899,N_47952);
and U48003 (N_48003,N_47793,N_47783);
and U48004 (N_48004,N_47986,N_47787);
nand U48005 (N_48005,N_47819,N_47951);
nand U48006 (N_48006,N_47877,N_47922);
xor U48007 (N_48007,N_47869,N_47908);
or U48008 (N_48008,N_47932,N_47829);
and U48009 (N_48009,N_47798,N_47790);
nor U48010 (N_48010,N_47821,N_47863);
or U48011 (N_48011,N_47902,N_47981);
or U48012 (N_48012,N_47892,N_47800);
xor U48013 (N_48013,N_47751,N_47797);
xnor U48014 (N_48014,N_47815,N_47855);
or U48015 (N_48015,N_47913,N_47903);
nor U48016 (N_48016,N_47977,N_47866);
xor U48017 (N_48017,N_47972,N_47928);
xor U48018 (N_48018,N_47988,N_47976);
or U48019 (N_48019,N_47758,N_47867);
and U48020 (N_48020,N_47954,N_47956);
xnor U48021 (N_48021,N_47875,N_47985);
nand U48022 (N_48022,N_47817,N_47763);
nor U48023 (N_48023,N_47964,N_47918);
xnor U48024 (N_48024,N_47890,N_47872);
xor U48025 (N_48025,N_47959,N_47961);
or U48026 (N_48026,N_47827,N_47774);
and U48027 (N_48027,N_47836,N_47923);
or U48028 (N_48028,N_47935,N_47936);
nand U48029 (N_48029,N_47870,N_47931);
or U48030 (N_48030,N_47934,N_47860);
and U48031 (N_48031,N_47808,N_47907);
nor U48032 (N_48032,N_47761,N_47888);
nor U48033 (N_48033,N_47843,N_47937);
nor U48034 (N_48034,N_47856,N_47853);
nor U48035 (N_48035,N_47926,N_47830);
or U48036 (N_48036,N_47984,N_47753);
nand U48037 (N_48037,N_47912,N_47945);
nor U48038 (N_48038,N_47778,N_47982);
nor U48039 (N_48039,N_47909,N_47939);
nand U48040 (N_48040,N_47772,N_47764);
nand U48041 (N_48041,N_47770,N_47920);
and U48042 (N_48042,N_47884,N_47823);
xor U48043 (N_48043,N_47777,N_47814);
nand U48044 (N_48044,N_47850,N_47983);
nor U48045 (N_48045,N_47837,N_47980);
and U48046 (N_48046,N_47801,N_47788);
nor U48047 (N_48047,N_47786,N_47759);
and U48048 (N_48048,N_47993,N_47938);
nand U48049 (N_48049,N_47832,N_47905);
xor U48050 (N_48050,N_47999,N_47991);
xnor U48051 (N_48051,N_47795,N_47887);
and U48052 (N_48052,N_47775,N_47768);
and U48053 (N_48053,N_47873,N_47810);
nand U48054 (N_48054,N_47944,N_47833);
nand U48055 (N_48055,N_47941,N_47886);
or U48056 (N_48056,N_47820,N_47978);
and U48057 (N_48057,N_47998,N_47969);
and U48058 (N_48058,N_47754,N_47766);
xnor U48059 (N_48059,N_47960,N_47940);
nor U48060 (N_48060,N_47958,N_47792);
nor U48061 (N_48061,N_47974,N_47990);
nor U48062 (N_48062,N_47765,N_47965);
xor U48063 (N_48063,N_47862,N_47894);
xnor U48064 (N_48064,N_47874,N_47813);
or U48065 (N_48065,N_47857,N_47762);
xor U48066 (N_48066,N_47780,N_47947);
nand U48067 (N_48067,N_47975,N_47844);
or U48068 (N_48068,N_47858,N_47910);
or U48069 (N_48069,N_47919,N_47996);
nor U48070 (N_48070,N_47897,N_47811);
xnor U48071 (N_48071,N_47950,N_47955);
nand U48072 (N_48072,N_47864,N_47848);
xor U48073 (N_48073,N_47971,N_47911);
nor U48074 (N_48074,N_47900,N_47839);
nand U48075 (N_48075,N_47824,N_47760);
and U48076 (N_48076,N_47915,N_47838);
nor U48077 (N_48077,N_47769,N_47962);
nor U48078 (N_48078,N_47791,N_47806);
and U48079 (N_48079,N_47828,N_47946);
nor U48080 (N_48080,N_47782,N_47826);
nor U48081 (N_48081,N_47841,N_47876);
xnor U48082 (N_48082,N_47898,N_47943);
nor U48083 (N_48083,N_47997,N_47776);
or U48084 (N_48084,N_47861,N_47871);
nor U48085 (N_48085,N_47812,N_47883);
and U48086 (N_48086,N_47849,N_47948);
nor U48087 (N_48087,N_47979,N_47847);
or U48088 (N_48088,N_47881,N_47895);
nand U48089 (N_48089,N_47973,N_47921);
nor U48090 (N_48090,N_47789,N_47822);
and U48091 (N_48091,N_47840,N_47796);
and U48092 (N_48092,N_47781,N_47906);
nor U48093 (N_48093,N_47925,N_47805);
xor U48094 (N_48094,N_47757,N_47924);
nor U48095 (N_48095,N_47859,N_47970);
or U48096 (N_48096,N_47803,N_47929);
xnor U48097 (N_48097,N_47893,N_47807);
or U48098 (N_48098,N_47794,N_47784);
or U48099 (N_48099,N_47865,N_47995);
xnor U48100 (N_48100,N_47878,N_47880);
nand U48101 (N_48101,N_47779,N_47755);
nand U48102 (N_48102,N_47804,N_47879);
or U48103 (N_48103,N_47831,N_47852);
and U48104 (N_48104,N_47771,N_47802);
xnor U48105 (N_48105,N_47835,N_47992);
nor U48106 (N_48106,N_47750,N_47942);
and U48107 (N_48107,N_47889,N_47868);
and U48108 (N_48108,N_47901,N_47809);
nor U48109 (N_48109,N_47927,N_47854);
or U48110 (N_48110,N_47933,N_47953);
nand U48111 (N_48111,N_47930,N_47914);
nor U48112 (N_48112,N_47752,N_47842);
or U48113 (N_48113,N_47846,N_47816);
nor U48114 (N_48114,N_47987,N_47967);
nor U48115 (N_48115,N_47966,N_47957);
nand U48116 (N_48116,N_47917,N_47851);
or U48117 (N_48117,N_47818,N_47904);
nand U48118 (N_48118,N_47825,N_47756);
xor U48119 (N_48119,N_47994,N_47785);
or U48120 (N_48120,N_47845,N_47989);
or U48121 (N_48121,N_47767,N_47834);
or U48122 (N_48122,N_47882,N_47773);
or U48123 (N_48123,N_47949,N_47968);
or U48124 (N_48124,N_47891,N_47799);
xor U48125 (N_48125,N_47988,N_47906);
and U48126 (N_48126,N_47842,N_47903);
nand U48127 (N_48127,N_47782,N_47769);
xnor U48128 (N_48128,N_47797,N_47827);
or U48129 (N_48129,N_47973,N_47936);
xor U48130 (N_48130,N_47876,N_47923);
or U48131 (N_48131,N_47969,N_47763);
nand U48132 (N_48132,N_47860,N_47810);
xor U48133 (N_48133,N_47954,N_47780);
xnor U48134 (N_48134,N_47851,N_47785);
or U48135 (N_48135,N_47817,N_47767);
xor U48136 (N_48136,N_47902,N_47927);
xnor U48137 (N_48137,N_47961,N_47955);
or U48138 (N_48138,N_47997,N_47871);
nand U48139 (N_48139,N_47862,N_47877);
xnor U48140 (N_48140,N_47832,N_47953);
nor U48141 (N_48141,N_47760,N_47889);
and U48142 (N_48142,N_47852,N_47959);
nor U48143 (N_48143,N_47907,N_47782);
and U48144 (N_48144,N_47840,N_47786);
xor U48145 (N_48145,N_47997,N_47876);
nand U48146 (N_48146,N_47894,N_47791);
and U48147 (N_48147,N_47768,N_47866);
nor U48148 (N_48148,N_47885,N_47993);
nor U48149 (N_48149,N_47872,N_47782);
nor U48150 (N_48150,N_47799,N_47918);
nand U48151 (N_48151,N_47931,N_47950);
nand U48152 (N_48152,N_47908,N_47880);
and U48153 (N_48153,N_47992,N_47986);
and U48154 (N_48154,N_47804,N_47838);
nand U48155 (N_48155,N_47751,N_47755);
nor U48156 (N_48156,N_47979,N_47830);
xor U48157 (N_48157,N_47932,N_47761);
or U48158 (N_48158,N_47915,N_47822);
or U48159 (N_48159,N_47911,N_47981);
xor U48160 (N_48160,N_47855,N_47879);
and U48161 (N_48161,N_47765,N_47875);
nand U48162 (N_48162,N_47871,N_47922);
nor U48163 (N_48163,N_47754,N_47836);
nand U48164 (N_48164,N_47914,N_47997);
nor U48165 (N_48165,N_47942,N_47913);
nand U48166 (N_48166,N_47970,N_47752);
and U48167 (N_48167,N_47821,N_47760);
or U48168 (N_48168,N_47786,N_47888);
nand U48169 (N_48169,N_47914,N_47911);
xor U48170 (N_48170,N_47948,N_47763);
nor U48171 (N_48171,N_47999,N_47838);
xor U48172 (N_48172,N_47906,N_47902);
or U48173 (N_48173,N_47825,N_47914);
and U48174 (N_48174,N_47923,N_47879);
nor U48175 (N_48175,N_47986,N_47937);
xor U48176 (N_48176,N_47931,N_47995);
nand U48177 (N_48177,N_47879,N_47927);
nand U48178 (N_48178,N_47815,N_47756);
nand U48179 (N_48179,N_47895,N_47828);
nand U48180 (N_48180,N_47887,N_47873);
or U48181 (N_48181,N_47940,N_47963);
or U48182 (N_48182,N_47824,N_47861);
nand U48183 (N_48183,N_47931,N_47929);
nor U48184 (N_48184,N_47947,N_47863);
xnor U48185 (N_48185,N_47850,N_47880);
and U48186 (N_48186,N_47875,N_47835);
nor U48187 (N_48187,N_47932,N_47976);
or U48188 (N_48188,N_47906,N_47764);
nand U48189 (N_48189,N_47785,N_47980);
xnor U48190 (N_48190,N_47798,N_47926);
nand U48191 (N_48191,N_47959,N_47752);
or U48192 (N_48192,N_47937,N_47830);
nor U48193 (N_48193,N_47802,N_47776);
nor U48194 (N_48194,N_47916,N_47802);
or U48195 (N_48195,N_47885,N_47776);
and U48196 (N_48196,N_47892,N_47884);
xor U48197 (N_48197,N_47953,N_47994);
nor U48198 (N_48198,N_47938,N_47818);
xor U48199 (N_48199,N_47779,N_47959);
nor U48200 (N_48200,N_47967,N_47975);
and U48201 (N_48201,N_47811,N_47815);
nor U48202 (N_48202,N_47860,N_47834);
and U48203 (N_48203,N_47784,N_47779);
nand U48204 (N_48204,N_47911,N_47856);
nor U48205 (N_48205,N_47758,N_47936);
nand U48206 (N_48206,N_47888,N_47849);
and U48207 (N_48207,N_47792,N_47770);
or U48208 (N_48208,N_47807,N_47766);
or U48209 (N_48209,N_47792,N_47982);
or U48210 (N_48210,N_47784,N_47774);
nor U48211 (N_48211,N_47777,N_47937);
xnor U48212 (N_48212,N_47808,N_47936);
xor U48213 (N_48213,N_47760,N_47959);
and U48214 (N_48214,N_47796,N_47850);
nand U48215 (N_48215,N_47858,N_47786);
nor U48216 (N_48216,N_47943,N_47825);
xor U48217 (N_48217,N_47897,N_47889);
nand U48218 (N_48218,N_47828,N_47845);
xnor U48219 (N_48219,N_47914,N_47836);
nor U48220 (N_48220,N_47914,N_47920);
nand U48221 (N_48221,N_47777,N_47927);
nor U48222 (N_48222,N_47903,N_47866);
and U48223 (N_48223,N_47881,N_47804);
or U48224 (N_48224,N_47975,N_47964);
xnor U48225 (N_48225,N_47796,N_47858);
nor U48226 (N_48226,N_47869,N_47939);
and U48227 (N_48227,N_47815,N_47913);
or U48228 (N_48228,N_47842,N_47807);
nor U48229 (N_48229,N_47835,N_47851);
and U48230 (N_48230,N_47820,N_47894);
xor U48231 (N_48231,N_47774,N_47913);
or U48232 (N_48232,N_47922,N_47750);
and U48233 (N_48233,N_47931,N_47985);
xor U48234 (N_48234,N_47768,N_47777);
or U48235 (N_48235,N_47879,N_47903);
nor U48236 (N_48236,N_47766,N_47992);
and U48237 (N_48237,N_47996,N_47900);
or U48238 (N_48238,N_47919,N_47978);
nand U48239 (N_48239,N_47957,N_47998);
and U48240 (N_48240,N_47864,N_47939);
and U48241 (N_48241,N_47974,N_47849);
and U48242 (N_48242,N_47879,N_47840);
xnor U48243 (N_48243,N_47795,N_47986);
nand U48244 (N_48244,N_47783,N_47858);
xnor U48245 (N_48245,N_47799,N_47892);
nand U48246 (N_48246,N_47781,N_47891);
nor U48247 (N_48247,N_47947,N_47890);
nor U48248 (N_48248,N_47831,N_47980);
and U48249 (N_48249,N_47791,N_47945);
or U48250 (N_48250,N_48163,N_48182);
xor U48251 (N_48251,N_48188,N_48121);
nor U48252 (N_48252,N_48213,N_48210);
nand U48253 (N_48253,N_48212,N_48098);
nor U48254 (N_48254,N_48181,N_48144);
nand U48255 (N_48255,N_48146,N_48239);
nand U48256 (N_48256,N_48183,N_48109);
nor U48257 (N_48257,N_48000,N_48081);
or U48258 (N_48258,N_48127,N_48236);
nand U48259 (N_48259,N_48067,N_48241);
nor U48260 (N_48260,N_48060,N_48131);
xnor U48261 (N_48261,N_48009,N_48080);
and U48262 (N_48262,N_48072,N_48045);
nor U48263 (N_48263,N_48101,N_48216);
xor U48264 (N_48264,N_48222,N_48008);
nand U48265 (N_48265,N_48186,N_48028);
or U48266 (N_48266,N_48026,N_48024);
nor U48267 (N_48267,N_48108,N_48065);
xor U48268 (N_48268,N_48090,N_48056);
nand U48269 (N_48269,N_48164,N_48202);
nand U48270 (N_48270,N_48134,N_48225);
xor U48271 (N_48271,N_48159,N_48016);
and U48272 (N_48272,N_48244,N_48166);
xor U48273 (N_48273,N_48150,N_48227);
and U48274 (N_48274,N_48054,N_48038);
xnor U48275 (N_48275,N_48177,N_48013);
or U48276 (N_48276,N_48092,N_48019);
nor U48277 (N_48277,N_48169,N_48125);
xnor U48278 (N_48278,N_48189,N_48178);
xor U48279 (N_48279,N_48033,N_48003);
nand U48280 (N_48280,N_48208,N_48145);
nor U48281 (N_48281,N_48075,N_48099);
nor U48282 (N_48282,N_48161,N_48014);
xor U48283 (N_48283,N_48199,N_48233);
xnor U48284 (N_48284,N_48057,N_48138);
and U48285 (N_48285,N_48192,N_48004);
nand U48286 (N_48286,N_48153,N_48195);
and U48287 (N_48287,N_48228,N_48018);
nand U48288 (N_48288,N_48068,N_48168);
nor U48289 (N_48289,N_48155,N_48066);
nor U48290 (N_48290,N_48105,N_48132);
nand U48291 (N_48291,N_48096,N_48086);
and U48292 (N_48292,N_48017,N_48115);
xor U48293 (N_48293,N_48139,N_48046);
nor U48294 (N_48294,N_48082,N_48128);
nand U48295 (N_48295,N_48051,N_48207);
xor U48296 (N_48296,N_48123,N_48135);
xnor U48297 (N_48297,N_48077,N_48093);
xor U48298 (N_48298,N_48247,N_48088);
nand U48299 (N_48299,N_48200,N_48073);
and U48300 (N_48300,N_48047,N_48036);
nor U48301 (N_48301,N_48196,N_48172);
and U48302 (N_48302,N_48006,N_48160);
xnor U48303 (N_48303,N_48104,N_48230);
and U48304 (N_48304,N_48107,N_48059);
nor U48305 (N_48305,N_48242,N_48097);
xnor U48306 (N_48306,N_48120,N_48193);
or U48307 (N_48307,N_48112,N_48091);
xor U48308 (N_48308,N_48012,N_48063);
or U48309 (N_48309,N_48126,N_48224);
or U48310 (N_48310,N_48151,N_48114);
nand U48311 (N_48311,N_48111,N_48234);
or U48312 (N_48312,N_48030,N_48007);
and U48313 (N_48313,N_48173,N_48174);
nor U48314 (N_48314,N_48218,N_48170);
or U48315 (N_48315,N_48142,N_48203);
xnor U48316 (N_48316,N_48235,N_48130);
xor U48317 (N_48317,N_48025,N_48175);
xnor U48318 (N_48318,N_48215,N_48084);
xor U48319 (N_48319,N_48023,N_48143);
nor U48320 (N_48320,N_48221,N_48156);
xor U48321 (N_48321,N_48122,N_48103);
or U48322 (N_48322,N_48152,N_48076);
nand U48323 (N_48323,N_48100,N_48240);
and U48324 (N_48324,N_48187,N_48083);
nor U48325 (N_48325,N_48042,N_48117);
nand U48326 (N_48326,N_48029,N_48087);
nand U48327 (N_48327,N_48157,N_48041);
nor U48328 (N_48328,N_48078,N_48079);
nand U48329 (N_48329,N_48113,N_48198);
and U48330 (N_48330,N_48053,N_48062);
nand U48331 (N_48331,N_48022,N_48197);
and U48332 (N_48332,N_48185,N_48043);
nand U48333 (N_48333,N_48070,N_48220);
or U48334 (N_48334,N_48167,N_48061);
nor U48335 (N_48335,N_48039,N_48205);
and U48336 (N_48336,N_48136,N_48020);
xnor U48337 (N_48337,N_48095,N_48141);
and U48338 (N_48338,N_48052,N_48124);
or U48339 (N_48339,N_48214,N_48001);
nand U48340 (N_48340,N_48037,N_48094);
or U48341 (N_48341,N_48217,N_48147);
xnor U48342 (N_48342,N_48162,N_48223);
nor U48343 (N_48343,N_48055,N_48226);
nor U48344 (N_48344,N_48201,N_48048);
xor U48345 (N_48345,N_48089,N_48191);
nor U48346 (N_48346,N_48040,N_48232);
or U48347 (N_48347,N_48118,N_48035);
nand U48348 (N_48348,N_48044,N_48204);
nor U48349 (N_48349,N_48248,N_48106);
or U48350 (N_48350,N_48165,N_48050);
and U48351 (N_48351,N_48219,N_48209);
and U48352 (N_48352,N_48137,N_48074);
nand U48353 (N_48353,N_48179,N_48231);
xnor U48354 (N_48354,N_48211,N_48110);
xor U48355 (N_48355,N_48049,N_48245);
xor U48356 (N_48356,N_48246,N_48027);
nand U48357 (N_48357,N_48085,N_48021);
xnor U48358 (N_48358,N_48206,N_48069);
or U48359 (N_48359,N_48176,N_48015);
nand U48360 (N_48360,N_48133,N_48229);
or U48361 (N_48361,N_48058,N_48190);
xor U48362 (N_48362,N_48184,N_48116);
or U48363 (N_48363,N_48149,N_48071);
xor U48364 (N_48364,N_48002,N_48243);
nand U48365 (N_48365,N_48032,N_48011);
nand U48366 (N_48366,N_48031,N_48249);
or U48367 (N_48367,N_48102,N_48034);
and U48368 (N_48368,N_48194,N_48238);
and U48369 (N_48369,N_48129,N_48148);
nor U48370 (N_48370,N_48005,N_48171);
and U48371 (N_48371,N_48119,N_48158);
or U48372 (N_48372,N_48010,N_48154);
and U48373 (N_48373,N_48140,N_48237);
or U48374 (N_48374,N_48064,N_48180);
xor U48375 (N_48375,N_48066,N_48210);
or U48376 (N_48376,N_48110,N_48100);
nand U48377 (N_48377,N_48179,N_48024);
nor U48378 (N_48378,N_48055,N_48231);
nand U48379 (N_48379,N_48082,N_48115);
nor U48380 (N_48380,N_48191,N_48160);
nor U48381 (N_48381,N_48185,N_48095);
xnor U48382 (N_48382,N_48175,N_48089);
and U48383 (N_48383,N_48052,N_48075);
nor U48384 (N_48384,N_48209,N_48187);
or U48385 (N_48385,N_48227,N_48044);
nor U48386 (N_48386,N_48025,N_48091);
or U48387 (N_48387,N_48072,N_48022);
and U48388 (N_48388,N_48144,N_48146);
and U48389 (N_48389,N_48209,N_48228);
and U48390 (N_48390,N_48125,N_48188);
and U48391 (N_48391,N_48082,N_48136);
nor U48392 (N_48392,N_48190,N_48236);
xor U48393 (N_48393,N_48172,N_48229);
or U48394 (N_48394,N_48202,N_48113);
or U48395 (N_48395,N_48185,N_48076);
nor U48396 (N_48396,N_48137,N_48231);
and U48397 (N_48397,N_48013,N_48121);
and U48398 (N_48398,N_48173,N_48014);
xor U48399 (N_48399,N_48143,N_48105);
xnor U48400 (N_48400,N_48126,N_48110);
and U48401 (N_48401,N_48007,N_48135);
and U48402 (N_48402,N_48038,N_48173);
xnor U48403 (N_48403,N_48226,N_48218);
nor U48404 (N_48404,N_48242,N_48187);
nor U48405 (N_48405,N_48242,N_48068);
xnor U48406 (N_48406,N_48143,N_48067);
nor U48407 (N_48407,N_48016,N_48110);
and U48408 (N_48408,N_48065,N_48055);
or U48409 (N_48409,N_48142,N_48062);
and U48410 (N_48410,N_48212,N_48190);
and U48411 (N_48411,N_48038,N_48003);
or U48412 (N_48412,N_48193,N_48184);
nand U48413 (N_48413,N_48168,N_48244);
and U48414 (N_48414,N_48082,N_48161);
xor U48415 (N_48415,N_48185,N_48093);
or U48416 (N_48416,N_48138,N_48135);
xor U48417 (N_48417,N_48063,N_48136);
and U48418 (N_48418,N_48072,N_48245);
and U48419 (N_48419,N_48210,N_48184);
xor U48420 (N_48420,N_48032,N_48020);
nand U48421 (N_48421,N_48060,N_48221);
nand U48422 (N_48422,N_48187,N_48212);
and U48423 (N_48423,N_48235,N_48159);
xor U48424 (N_48424,N_48215,N_48101);
or U48425 (N_48425,N_48049,N_48127);
or U48426 (N_48426,N_48036,N_48074);
nor U48427 (N_48427,N_48077,N_48106);
or U48428 (N_48428,N_48242,N_48229);
nand U48429 (N_48429,N_48120,N_48161);
or U48430 (N_48430,N_48153,N_48009);
and U48431 (N_48431,N_48133,N_48076);
nand U48432 (N_48432,N_48140,N_48192);
or U48433 (N_48433,N_48235,N_48201);
and U48434 (N_48434,N_48045,N_48035);
nand U48435 (N_48435,N_48192,N_48016);
xnor U48436 (N_48436,N_48006,N_48099);
or U48437 (N_48437,N_48225,N_48224);
nor U48438 (N_48438,N_48241,N_48191);
nand U48439 (N_48439,N_48196,N_48022);
xnor U48440 (N_48440,N_48028,N_48140);
or U48441 (N_48441,N_48073,N_48225);
or U48442 (N_48442,N_48076,N_48141);
nand U48443 (N_48443,N_48098,N_48153);
or U48444 (N_48444,N_48034,N_48110);
xnor U48445 (N_48445,N_48199,N_48167);
and U48446 (N_48446,N_48107,N_48019);
or U48447 (N_48447,N_48170,N_48158);
nand U48448 (N_48448,N_48013,N_48026);
nor U48449 (N_48449,N_48073,N_48210);
and U48450 (N_48450,N_48229,N_48017);
nor U48451 (N_48451,N_48009,N_48007);
and U48452 (N_48452,N_48007,N_48006);
nand U48453 (N_48453,N_48001,N_48172);
or U48454 (N_48454,N_48026,N_48226);
nor U48455 (N_48455,N_48014,N_48053);
or U48456 (N_48456,N_48064,N_48089);
and U48457 (N_48457,N_48107,N_48202);
xor U48458 (N_48458,N_48213,N_48207);
or U48459 (N_48459,N_48132,N_48137);
nand U48460 (N_48460,N_48171,N_48130);
and U48461 (N_48461,N_48097,N_48107);
xnor U48462 (N_48462,N_48139,N_48034);
nor U48463 (N_48463,N_48051,N_48213);
and U48464 (N_48464,N_48023,N_48088);
nor U48465 (N_48465,N_48084,N_48244);
xnor U48466 (N_48466,N_48116,N_48178);
and U48467 (N_48467,N_48180,N_48004);
or U48468 (N_48468,N_48088,N_48015);
nor U48469 (N_48469,N_48051,N_48216);
nand U48470 (N_48470,N_48163,N_48245);
nor U48471 (N_48471,N_48228,N_48039);
nand U48472 (N_48472,N_48220,N_48146);
nor U48473 (N_48473,N_48171,N_48121);
nor U48474 (N_48474,N_48229,N_48248);
xor U48475 (N_48475,N_48145,N_48036);
nand U48476 (N_48476,N_48194,N_48147);
nor U48477 (N_48477,N_48212,N_48245);
and U48478 (N_48478,N_48163,N_48117);
or U48479 (N_48479,N_48160,N_48059);
and U48480 (N_48480,N_48082,N_48189);
and U48481 (N_48481,N_48028,N_48051);
and U48482 (N_48482,N_48092,N_48187);
and U48483 (N_48483,N_48123,N_48034);
nor U48484 (N_48484,N_48099,N_48212);
nand U48485 (N_48485,N_48076,N_48171);
xor U48486 (N_48486,N_48144,N_48248);
nor U48487 (N_48487,N_48008,N_48173);
and U48488 (N_48488,N_48023,N_48135);
or U48489 (N_48489,N_48236,N_48134);
nor U48490 (N_48490,N_48112,N_48204);
nor U48491 (N_48491,N_48068,N_48101);
xnor U48492 (N_48492,N_48241,N_48059);
or U48493 (N_48493,N_48111,N_48169);
and U48494 (N_48494,N_48230,N_48213);
and U48495 (N_48495,N_48097,N_48179);
nand U48496 (N_48496,N_48053,N_48095);
nand U48497 (N_48497,N_48004,N_48153);
xnor U48498 (N_48498,N_48101,N_48035);
nor U48499 (N_48499,N_48227,N_48225);
or U48500 (N_48500,N_48335,N_48389);
nor U48501 (N_48501,N_48433,N_48370);
and U48502 (N_48502,N_48392,N_48378);
or U48503 (N_48503,N_48406,N_48405);
nor U48504 (N_48504,N_48302,N_48288);
or U48505 (N_48505,N_48330,N_48496);
nor U48506 (N_48506,N_48390,N_48256);
nand U48507 (N_48507,N_48254,N_48316);
or U48508 (N_48508,N_48482,N_48385);
and U48509 (N_48509,N_48439,N_48473);
xor U48510 (N_48510,N_48437,N_48391);
nand U48511 (N_48511,N_48467,N_48322);
nand U48512 (N_48512,N_48279,N_48325);
or U48513 (N_48513,N_48435,N_48308);
nand U48514 (N_48514,N_48402,N_48468);
xor U48515 (N_48515,N_48273,N_48347);
and U48516 (N_48516,N_48491,N_48451);
nand U48517 (N_48517,N_48266,N_48376);
and U48518 (N_48518,N_48354,N_48463);
or U48519 (N_48519,N_48494,N_48315);
nor U48520 (N_48520,N_48282,N_48331);
xor U48521 (N_48521,N_48295,N_48409);
and U48522 (N_48522,N_48386,N_48440);
xnor U48523 (N_48523,N_48480,N_48351);
xnor U48524 (N_48524,N_48303,N_48344);
xor U48525 (N_48525,N_48411,N_48292);
or U48526 (N_48526,N_48277,N_48445);
or U48527 (N_48527,N_48479,N_48380);
xor U48528 (N_48528,N_48349,N_48407);
and U48529 (N_48529,N_48498,N_48353);
xor U48530 (N_48530,N_48458,N_48436);
and U48531 (N_48531,N_48362,N_48269);
xnor U48532 (N_48532,N_48404,N_48311);
or U48533 (N_48533,N_48313,N_48306);
nor U48534 (N_48534,N_48395,N_48324);
nor U48535 (N_48535,N_48429,N_48477);
nor U48536 (N_48536,N_48336,N_48393);
nand U48537 (N_48537,N_48488,N_48490);
nand U48538 (N_48538,N_48487,N_48280);
or U48539 (N_48539,N_48450,N_48276);
nor U48540 (N_48540,N_48412,N_48421);
xor U48541 (N_48541,N_48352,N_48260);
or U48542 (N_48542,N_48371,N_48470);
or U48543 (N_48543,N_48413,N_48307);
nand U48544 (N_48544,N_48368,N_48340);
nor U48545 (N_48545,N_48384,N_48387);
nor U48546 (N_48546,N_48483,N_48305);
xnor U48547 (N_48547,N_48449,N_48418);
or U48548 (N_48548,N_48275,N_48334);
and U48549 (N_48549,N_48396,N_48442);
nand U48550 (N_48550,N_48297,N_48318);
nor U48551 (N_48551,N_48461,N_48294);
nor U48552 (N_48552,N_48299,N_48360);
nor U48553 (N_48553,N_48300,N_48264);
xnor U48554 (N_48554,N_48377,N_48323);
xnor U48555 (N_48555,N_48489,N_48348);
nor U48556 (N_48556,N_48492,N_48281);
and U48557 (N_48557,N_48253,N_48417);
and U48558 (N_48558,N_48382,N_48251);
xor U48559 (N_48559,N_48444,N_48363);
or U48560 (N_48560,N_48366,N_48422);
nor U48561 (N_48561,N_48394,N_48367);
or U48562 (N_48562,N_48454,N_48272);
nand U48563 (N_48563,N_48459,N_48296);
nand U48564 (N_48564,N_48481,N_48472);
xnor U48565 (N_48565,N_48321,N_48414);
nor U48566 (N_48566,N_48438,N_48257);
or U48567 (N_48567,N_48310,N_48457);
nand U48568 (N_48568,N_48443,N_48298);
nand U48569 (N_48569,N_48416,N_48493);
and U48570 (N_48570,N_48259,N_48304);
and U48571 (N_48571,N_48397,N_48486);
or U48572 (N_48572,N_48283,N_48466);
nor U48573 (N_48573,N_48268,N_48428);
nor U48574 (N_48574,N_48369,N_48420);
xnor U48575 (N_48575,N_48293,N_48441);
and U48576 (N_48576,N_48426,N_48497);
xnor U48577 (N_48577,N_48359,N_48339);
xor U48578 (N_48578,N_48398,N_48401);
xnor U48579 (N_48579,N_48333,N_48427);
nor U48580 (N_48580,N_48356,N_48383);
and U48581 (N_48581,N_48460,N_48285);
and U48582 (N_48582,N_48345,N_48456);
or U48583 (N_48583,N_48263,N_48290);
and U48584 (N_48584,N_48261,N_48291);
nand U48585 (N_48585,N_48319,N_48364);
and U48586 (N_48586,N_48250,N_48431);
nor U48587 (N_48587,N_48410,N_48289);
and U48588 (N_48588,N_48309,N_48374);
and U48589 (N_48589,N_48284,N_48271);
xnor U48590 (N_48590,N_48400,N_48312);
nor U48591 (N_48591,N_48286,N_48357);
and U48592 (N_48592,N_48341,N_48419);
xor U48593 (N_48593,N_48448,N_48373);
xnor U48594 (N_48594,N_48471,N_48258);
nor U48595 (N_48595,N_48314,N_48262);
nor U48596 (N_48596,N_48484,N_48446);
and U48597 (N_48597,N_48464,N_48469);
or U48598 (N_48598,N_48270,N_48432);
or U48599 (N_48599,N_48423,N_48434);
or U48600 (N_48600,N_48447,N_48452);
and U48601 (N_48601,N_48320,N_48328);
nor U48602 (N_48602,N_48267,N_48278);
or U48603 (N_48603,N_48252,N_48476);
nand U48604 (N_48604,N_48478,N_48465);
and U48605 (N_48605,N_48274,N_48301);
and U48606 (N_48606,N_48355,N_48372);
nor U48607 (N_48607,N_48408,N_48317);
nand U48608 (N_48608,N_48346,N_48329);
nand U48609 (N_48609,N_48337,N_48255);
nor U48610 (N_48610,N_48327,N_48326);
and U48611 (N_48611,N_48375,N_48388);
xor U48612 (N_48612,N_48430,N_48415);
and U48613 (N_48613,N_48462,N_48379);
nand U48614 (N_48614,N_48358,N_48265);
nor U48615 (N_48615,N_48365,N_48474);
nand U48616 (N_48616,N_48403,N_48499);
xor U48617 (N_48617,N_48424,N_48381);
nor U48618 (N_48618,N_48425,N_48342);
nor U48619 (N_48619,N_48361,N_48350);
nor U48620 (N_48620,N_48455,N_48495);
or U48621 (N_48621,N_48475,N_48453);
nor U48622 (N_48622,N_48332,N_48343);
nand U48623 (N_48623,N_48485,N_48287);
nand U48624 (N_48624,N_48338,N_48399);
and U48625 (N_48625,N_48443,N_48485);
nor U48626 (N_48626,N_48347,N_48380);
nand U48627 (N_48627,N_48477,N_48270);
nand U48628 (N_48628,N_48313,N_48393);
xnor U48629 (N_48629,N_48448,N_48403);
nor U48630 (N_48630,N_48392,N_48259);
nor U48631 (N_48631,N_48281,N_48333);
or U48632 (N_48632,N_48418,N_48304);
nand U48633 (N_48633,N_48346,N_48389);
or U48634 (N_48634,N_48497,N_48393);
and U48635 (N_48635,N_48441,N_48291);
and U48636 (N_48636,N_48420,N_48398);
xnor U48637 (N_48637,N_48411,N_48274);
and U48638 (N_48638,N_48260,N_48395);
and U48639 (N_48639,N_48400,N_48288);
or U48640 (N_48640,N_48339,N_48276);
nand U48641 (N_48641,N_48470,N_48289);
and U48642 (N_48642,N_48257,N_48484);
nor U48643 (N_48643,N_48281,N_48468);
xnor U48644 (N_48644,N_48279,N_48329);
nor U48645 (N_48645,N_48284,N_48483);
nor U48646 (N_48646,N_48332,N_48342);
nor U48647 (N_48647,N_48481,N_48438);
xnor U48648 (N_48648,N_48270,N_48284);
nor U48649 (N_48649,N_48310,N_48280);
nand U48650 (N_48650,N_48348,N_48491);
nand U48651 (N_48651,N_48470,N_48273);
or U48652 (N_48652,N_48453,N_48326);
and U48653 (N_48653,N_48494,N_48432);
or U48654 (N_48654,N_48346,N_48268);
xnor U48655 (N_48655,N_48383,N_48388);
or U48656 (N_48656,N_48420,N_48427);
xor U48657 (N_48657,N_48389,N_48315);
and U48658 (N_48658,N_48344,N_48382);
or U48659 (N_48659,N_48307,N_48294);
nand U48660 (N_48660,N_48308,N_48392);
and U48661 (N_48661,N_48288,N_48323);
and U48662 (N_48662,N_48401,N_48281);
nor U48663 (N_48663,N_48463,N_48286);
and U48664 (N_48664,N_48457,N_48387);
or U48665 (N_48665,N_48383,N_48440);
nor U48666 (N_48666,N_48480,N_48343);
xnor U48667 (N_48667,N_48431,N_48269);
nor U48668 (N_48668,N_48281,N_48427);
xor U48669 (N_48669,N_48353,N_48384);
nand U48670 (N_48670,N_48348,N_48486);
and U48671 (N_48671,N_48291,N_48447);
and U48672 (N_48672,N_48396,N_48403);
xor U48673 (N_48673,N_48409,N_48309);
or U48674 (N_48674,N_48336,N_48327);
nand U48675 (N_48675,N_48304,N_48332);
xnor U48676 (N_48676,N_48266,N_48262);
nand U48677 (N_48677,N_48304,N_48285);
nor U48678 (N_48678,N_48271,N_48437);
nand U48679 (N_48679,N_48350,N_48446);
nand U48680 (N_48680,N_48395,N_48429);
xor U48681 (N_48681,N_48263,N_48317);
or U48682 (N_48682,N_48426,N_48482);
or U48683 (N_48683,N_48330,N_48423);
xnor U48684 (N_48684,N_48291,N_48365);
and U48685 (N_48685,N_48375,N_48392);
nand U48686 (N_48686,N_48316,N_48310);
and U48687 (N_48687,N_48427,N_48271);
nand U48688 (N_48688,N_48460,N_48453);
and U48689 (N_48689,N_48379,N_48367);
and U48690 (N_48690,N_48483,N_48316);
and U48691 (N_48691,N_48460,N_48261);
nor U48692 (N_48692,N_48422,N_48455);
nor U48693 (N_48693,N_48321,N_48491);
nor U48694 (N_48694,N_48362,N_48416);
xnor U48695 (N_48695,N_48444,N_48495);
xor U48696 (N_48696,N_48467,N_48359);
nand U48697 (N_48697,N_48323,N_48387);
or U48698 (N_48698,N_48471,N_48287);
nor U48699 (N_48699,N_48326,N_48417);
and U48700 (N_48700,N_48382,N_48383);
nand U48701 (N_48701,N_48414,N_48488);
or U48702 (N_48702,N_48362,N_48294);
nor U48703 (N_48703,N_48273,N_48299);
xnor U48704 (N_48704,N_48321,N_48477);
and U48705 (N_48705,N_48331,N_48266);
nand U48706 (N_48706,N_48424,N_48408);
nand U48707 (N_48707,N_48406,N_48326);
xor U48708 (N_48708,N_48321,N_48291);
nand U48709 (N_48709,N_48451,N_48261);
and U48710 (N_48710,N_48293,N_48323);
and U48711 (N_48711,N_48384,N_48440);
nand U48712 (N_48712,N_48382,N_48305);
nand U48713 (N_48713,N_48427,N_48274);
nand U48714 (N_48714,N_48293,N_48334);
or U48715 (N_48715,N_48494,N_48319);
and U48716 (N_48716,N_48347,N_48439);
xor U48717 (N_48717,N_48351,N_48380);
xor U48718 (N_48718,N_48332,N_48266);
or U48719 (N_48719,N_48486,N_48490);
nand U48720 (N_48720,N_48339,N_48266);
nor U48721 (N_48721,N_48390,N_48322);
or U48722 (N_48722,N_48469,N_48372);
and U48723 (N_48723,N_48346,N_48383);
or U48724 (N_48724,N_48347,N_48336);
xnor U48725 (N_48725,N_48397,N_48328);
and U48726 (N_48726,N_48362,N_48393);
xor U48727 (N_48727,N_48434,N_48259);
and U48728 (N_48728,N_48308,N_48475);
or U48729 (N_48729,N_48387,N_48490);
xor U48730 (N_48730,N_48409,N_48499);
and U48731 (N_48731,N_48293,N_48444);
nand U48732 (N_48732,N_48483,N_48343);
and U48733 (N_48733,N_48469,N_48274);
xnor U48734 (N_48734,N_48497,N_48312);
nand U48735 (N_48735,N_48273,N_48490);
nand U48736 (N_48736,N_48276,N_48373);
and U48737 (N_48737,N_48375,N_48472);
nand U48738 (N_48738,N_48458,N_48341);
or U48739 (N_48739,N_48470,N_48403);
nand U48740 (N_48740,N_48298,N_48270);
xor U48741 (N_48741,N_48454,N_48298);
nand U48742 (N_48742,N_48455,N_48470);
or U48743 (N_48743,N_48300,N_48414);
nor U48744 (N_48744,N_48290,N_48277);
xor U48745 (N_48745,N_48328,N_48451);
xor U48746 (N_48746,N_48458,N_48250);
nor U48747 (N_48747,N_48265,N_48484);
nand U48748 (N_48748,N_48381,N_48269);
xor U48749 (N_48749,N_48424,N_48364);
xnor U48750 (N_48750,N_48523,N_48520);
and U48751 (N_48751,N_48598,N_48573);
xnor U48752 (N_48752,N_48544,N_48532);
xnor U48753 (N_48753,N_48697,N_48537);
or U48754 (N_48754,N_48600,N_48654);
or U48755 (N_48755,N_48622,N_48500);
nand U48756 (N_48756,N_48538,N_48620);
and U48757 (N_48757,N_48530,N_48578);
xnor U48758 (N_48758,N_48547,N_48664);
or U48759 (N_48759,N_48658,N_48713);
or U48760 (N_48760,N_48735,N_48648);
xnor U48761 (N_48761,N_48553,N_48683);
nand U48762 (N_48762,N_48638,N_48728);
xnor U48763 (N_48763,N_48724,N_48727);
xor U48764 (N_48764,N_48597,N_48723);
xor U48765 (N_48765,N_48639,N_48700);
nor U48766 (N_48766,N_48703,N_48725);
nand U48767 (N_48767,N_48514,N_48702);
or U48768 (N_48768,N_48696,N_48592);
and U48769 (N_48769,N_48693,N_48593);
nand U48770 (N_48770,N_48528,N_48706);
or U48771 (N_48771,N_48733,N_48572);
xnor U48772 (N_48772,N_48541,N_48681);
nand U48773 (N_48773,N_48741,N_48591);
xnor U48774 (N_48774,N_48555,N_48628);
or U48775 (N_48775,N_48565,N_48534);
nor U48776 (N_48776,N_48743,N_48580);
nor U48777 (N_48777,N_48617,N_48692);
nor U48778 (N_48778,N_48709,N_48655);
nor U48779 (N_48779,N_48698,N_48557);
nor U48780 (N_48780,N_48601,N_48686);
or U48781 (N_48781,N_48732,N_48720);
and U48782 (N_48782,N_48531,N_48548);
nand U48783 (N_48783,N_48662,N_48614);
nand U48784 (N_48784,N_48651,N_48734);
nor U48785 (N_48785,N_48582,N_48521);
nand U48786 (N_48786,N_48558,N_48586);
xor U48787 (N_48787,N_48623,N_48695);
and U48788 (N_48788,N_48667,N_48561);
xnor U48789 (N_48789,N_48744,N_48563);
nor U48790 (N_48790,N_48571,N_48513);
and U48791 (N_48791,N_48745,N_48650);
nand U48792 (N_48792,N_48653,N_48504);
nor U48793 (N_48793,N_48595,N_48596);
and U48794 (N_48794,N_48642,N_48705);
xor U48795 (N_48795,N_48568,N_48740);
xor U48796 (N_48796,N_48673,N_48640);
nand U48797 (N_48797,N_48619,N_48739);
and U48798 (N_48798,N_48549,N_48682);
nor U48799 (N_48799,N_48659,N_48570);
and U48800 (N_48800,N_48577,N_48699);
nor U48801 (N_48801,N_48503,N_48737);
and U48802 (N_48802,N_48707,N_48540);
nand U48803 (N_48803,N_48714,N_48581);
and U48804 (N_48804,N_48590,N_48661);
nand U48805 (N_48805,N_48506,N_48527);
or U48806 (N_48806,N_48731,N_48677);
xor U48807 (N_48807,N_48660,N_48637);
xor U48808 (N_48808,N_48625,N_48652);
nor U48809 (N_48809,N_48704,N_48501);
nand U48810 (N_48810,N_48621,N_48564);
xnor U48811 (N_48811,N_48644,N_48626);
and U48812 (N_48812,N_48738,N_48689);
or U48813 (N_48813,N_48566,N_48574);
xnor U48814 (N_48814,N_48605,N_48630);
or U48815 (N_48815,N_48618,N_48516);
or U48816 (N_48816,N_48672,N_48676);
nand U48817 (N_48817,N_48730,N_48663);
or U48818 (N_48818,N_48665,N_48610);
or U48819 (N_48819,N_48701,N_48583);
and U48820 (N_48820,N_48721,N_48694);
nand U48821 (N_48821,N_48656,N_48559);
and U48822 (N_48822,N_48515,N_48669);
xor U48823 (N_48823,N_48602,N_48518);
or U48824 (N_48824,N_48729,N_48576);
or U48825 (N_48825,N_48675,N_48685);
xor U48826 (N_48826,N_48641,N_48613);
or U48827 (N_48827,N_48616,N_48509);
nand U48828 (N_48828,N_48569,N_48615);
xnor U48829 (N_48829,N_48552,N_48687);
and U48830 (N_48830,N_48624,N_48711);
nor U48831 (N_48831,N_48708,N_48585);
nor U48832 (N_48832,N_48512,N_48594);
and U48833 (N_48833,N_48668,N_48562);
and U48834 (N_48834,N_48631,N_48643);
and U48835 (N_48835,N_48554,N_48535);
or U48836 (N_48836,N_48636,N_48533);
nor U48837 (N_48837,N_48680,N_48678);
and U48838 (N_48838,N_48584,N_48670);
nand U48839 (N_48839,N_48715,N_48684);
nor U48840 (N_48840,N_48525,N_48609);
or U48841 (N_48841,N_48567,N_48632);
and U48842 (N_48842,N_48719,N_48666);
nand U48843 (N_48843,N_48749,N_48671);
nor U48844 (N_48844,N_48606,N_48629);
and U48845 (N_48845,N_48551,N_48603);
nor U48846 (N_48846,N_48647,N_48505);
nand U48847 (N_48847,N_48635,N_48545);
xnor U48848 (N_48848,N_48608,N_48679);
and U48849 (N_48849,N_48646,N_48717);
and U48850 (N_48850,N_48550,N_48604);
xor U48851 (N_48851,N_48587,N_48726);
xnor U48852 (N_48852,N_48560,N_48526);
or U48853 (N_48853,N_48722,N_48688);
and U48854 (N_48854,N_48502,N_48657);
nor U48855 (N_48855,N_48607,N_48718);
xnor U48856 (N_48856,N_48599,N_48556);
nor U48857 (N_48857,N_48519,N_48690);
nand U48858 (N_48858,N_48611,N_48710);
and U48859 (N_48859,N_48539,N_48508);
or U48860 (N_48860,N_48529,N_48746);
nand U48861 (N_48861,N_48536,N_48511);
or U48862 (N_48862,N_48627,N_48712);
nor U48863 (N_48863,N_48612,N_48510);
nor U48864 (N_48864,N_48579,N_48748);
xnor U48865 (N_48865,N_48517,N_48507);
nor U48866 (N_48866,N_48588,N_48634);
nand U48867 (N_48867,N_48543,N_48522);
and U48868 (N_48868,N_48716,N_48633);
or U48869 (N_48869,N_48691,N_48589);
nand U48870 (N_48870,N_48742,N_48575);
nand U48871 (N_48871,N_48649,N_48546);
xor U48872 (N_48872,N_48645,N_48747);
nor U48873 (N_48873,N_48736,N_48674);
or U48874 (N_48874,N_48524,N_48542);
nand U48875 (N_48875,N_48598,N_48582);
or U48876 (N_48876,N_48566,N_48533);
nand U48877 (N_48877,N_48690,N_48646);
and U48878 (N_48878,N_48670,N_48535);
nor U48879 (N_48879,N_48707,N_48727);
nor U48880 (N_48880,N_48602,N_48545);
and U48881 (N_48881,N_48536,N_48628);
and U48882 (N_48882,N_48594,N_48707);
and U48883 (N_48883,N_48669,N_48548);
or U48884 (N_48884,N_48540,N_48582);
nand U48885 (N_48885,N_48513,N_48706);
or U48886 (N_48886,N_48644,N_48506);
nand U48887 (N_48887,N_48664,N_48732);
and U48888 (N_48888,N_48642,N_48728);
xor U48889 (N_48889,N_48730,N_48731);
nor U48890 (N_48890,N_48594,N_48504);
xnor U48891 (N_48891,N_48551,N_48555);
or U48892 (N_48892,N_48711,N_48671);
or U48893 (N_48893,N_48665,N_48675);
and U48894 (N_48894,N_48614,N_48549);
nor U48895 (N_48895,N_48532,N_48626);
nor U48896 (N_48896,N_48541,N_48522);
nor U48897 (N_48897,N_48503,N_48746);
xnor U48898 (N_48898,N_48658,N_48631);
and U48899 (N_48899,N_48583,N_48673);
nor U48900 (N_48900,N_48702,N_48614);
nor U48901 (N_48901,N_48570,N_48645);
and U48902 (N_48902,N_48610,N_48583);
and U48903 (N_48903,N_48645,N_48687);
xnor U48904 (N_48904,N_48651,N_48714);
xnor U48905 (N_48905,N_48647,N_48681);
or U48906 (N_48906,N_48660,N_48631);
or U48907 (N_48907,N_48596,N_48630);
xor U48908 (N_48908,N_48588,N_48508);
and U48909 (N_48909,N_48633,N_48555);
and U48910 (N_48910,N_48687,N_48675);
and U48911 (N_48911,N_48726,N_48563);
and U48912 (N_48912,N_48714,N_48621);
and U48913 (N_48913,N_48701,N_48717);
and U48914 (N_48914,N_48725,N_48665);
xor U48915 (N_48915,N_48576,N_48722);
nand U48916 (N_48916,N_48690,N_48711);
and U48917 (N_48917,N_48633,N_48526);
nand U48918 (N_48918,N_48513,N_48545);
and U48919 (N_48919,N_48607,N_48572);
and U48920 (N_48920,N_48699,N_48501);
nor U48921 (N_48921,N_48657,N_48745);
nand U48922 (N_48922,N_48686,N_48733);
and U48923 (N_48923,N_48621,N_48602);
or U48924 (N_48924,N_48515,N_48574);
nor U48925 (N_48925,N_48507,N_48739);
and U48926 (N_48926,N_48693,N_48628);
nand U48927 (N_48927,N_48672,N_48649);
nand U48928 (N_48928,N_48745,N_48513);
nand U48929 (N_48929,N_48514,N_48736);
or U48930 (N_48930,N_48633,N_48597);
nand U48931 (N_48931,N_48549,N_48716);
nand U48932 (N_48932,N_48503,N_48556);
and U48933 (N_48933,N_48675,N_48630);
xnor U48934 (N_48934,N_48646,N_48656);
or U48935 (N_48935,N_48579,N_48700);
or U48936 (N_48936,N_48532,N_48547);
nand U48937 (N_48937,N_48606,N_48680);
nor U48938 (N_48938,N_48511,N_48711);
or U48939 (N_48939,N_48718,N_48586);
xor U48940 (N_48940,N_48626,N_48735);
xnor U48941 (N_48941,N_48554,N_48735);
nand U48942 (N_48942,N_48746,N_48692);
xnor U48943 (N_48943,N_48598,N_48560);
nor U48944 (N_48944,N_48722,N_48523);
nand U48945 (N_48945,N_48657,N_48724);
and U48946 (N_48946,N_48625,N_48738);
or U48947 (N_48947,N_48551,N_48591);
nand U48948 (N_48948,N_48651,N_48702);
xnor U48949 (N_48949,N_48569,N_48684);
and U48950 (N_48950,N_48646,N_48663);
nand U48951 (N_48951,N_48730,N_48611);
or U48952 (N_48952,N_48734,N_48557);
or U48953 (N_48953,N_48502,N_48582);
nand U48954 (N_48954,N_48703,N_48651);
xor U48955 (N_48955,N_48722,N_48735);
nand U48956 (N_48956,N_48748,N_48649);
and U48957 (N_48957,N_48532,N_48627);
and U48958 (N_48958,N_48548,N_48620);
xnor U48959 (N_48959,N_48727,N_48600);
nor U48960 (N_48960,N_48586,N_48625);
nor U48961 (N_48961,N_48543,N_48519);
nor U48962 (N_48962,N_48528,N_48558);
or U48963 (N_48963,N_48734,N_48519);
nor U48964 (N_48964,N_48530,N_48687);
and U48965 (N_48965,N_48507,N_48586);
and U48966 (N_48966,N_48684,N_48570);
nand U48967 (N_48967,N_48523,N_48504);
xnor U48968 (N_48968,N_48696,N_48641);
and U48969 (N_48969,N_48677,N_48707);
nand U48970 (N_48970,N_48590,N_48635);
xnor U48971 (N_48971,N_48722,N_48714);
nand U48972 (N_48972,N_48680,N_48645);
and U48973 (N_48973,N_48657,N_48640);
nor U48974 (N_48974,N_48542,N_48584);
nand U48975 (N_48975,N_48583,N_48523);
xnor U48976 (N_48976,N_48501,N_48558);
and U48977 (N_48977,N_48559,N_48653);
or U48978 (N_48978,N_48630,N_48537);
nor U48979 (N_48979,N_48584,N_48667);
nor U48980 (N_48980,N_48506,N_48517);
xor U48981 (N_48981,N_48625,N_48713);
and U48982 (N_48982,N_48576,N_48529);
nand U48983 (N_48983,N_48748,N_48619);
or U48984 (N_48984,N_48704,N_48646);
nand U48985 (N_48985,N_48656,N_48617);
and U48986 (N_48986,N_48565,N_48714);
or U48987 (N_48987,N_48600,N_48553);
and U48988 (N_48988,N_48734,N_48614);
or U48989 (N_48989,N_48700,N_48740);
xor U48990 (N_48990,N_48525,N_48749);
or U48991 (N_48991,N_48608,N_48607);
nor U48992 (N_48992,N_48515,N_48609);
nand U48993 (N_48993,N_48613,N_48539);
xnor U48994 (N_48994,N_48749,N_48663);
or U48995 (N_48995,N_48603,N_48524);
nor U48996 (N_48996,N_48582,N_48561);
nor U48997 (N_48997,N_48742,N_48704);
nor U48998 (N_48998,N_48502,N_48697);
and U48999 (N_48999,N_48696,N_48520);
nor U49000 (N_49000,N_48911,N_48775);
nor U49001 (N_49001,N_48791,N_48910);
nand U49002 (N_49002,N_48840,N_48919);
xor U49003 (N_49003,N_48795,N_48852);
nor U49004 (N_49004,N_48947,N_48777);
xor U49005 (N_49005,N_48930,N_48962);
and U49006 (N_49006,N_48819,N_48996);
nand U49007 (N_49007,N_48994,N_48943);
xnor U49008 (N_49008,N_48813,N_48968);
nor U49009 (N_49009,N_48965,N_48891);
or U49010 (N_49010,N_48948,N_48763);
or U49011 (N_49011,N_48983,N_48826);
nor U49012 (N_49012,N_48766,N_48885);
xor U49013 (N_49013,N_48917,N_48796);
or U49014 (N_49014,N_48824,N_48873);
xnor U49015 (N_49015,N_48990,N_48771);
xor U49016 (N_49016,N_48834,N_48982);
or U49017 (N_49017,N_48854,N_48933);
and U49018 (N_49018,N_48970,N_48963);
nor U49019 (N_49019,N_48822,N_48935);
nand U49020 (N_49020,N_48905,N_48750);
nand U49021 (N_49021,N_48960,N_48801);
and U49022 (N_49022,N_48799,N_48877);
xor U49023 (N_49023,N_48876,N_48986);
nand U49024 (N_49024,N_48850,N_48894);
or U49025 (N_49025,N_48918,N_48853);
and U49026 (N_49026,N_48913,N_48835);
nor U49027 (N_49027,N_48764,N_48769);
xnor U49028 (N_49028,N_48912,N_48859);
nor U49029 (N_49029,N_48939,N_48808);
and U49030 (N_49030,N_48838,N_48780);
nor U49031 (N_49031,N_48847,N_48855);
and U49032 (N_49032,N_48787,N_48793);
nor U49033 (N_49033,N_48844,N_48800);
or U49034 (N_49034,N_48762,N_48839);
nand U49035 (N_49035,N_48991,N_48936);
or U49036 (N_49036,N_48971,N_48938);
nand U49037 (N_49037,N_48862,N_48833);
nor U49038 (N_49038,N_48765,N_48900);
nand U49039 (N_49039,N_48881,N_48916);
or U49040 (N_49040,N_48898,N_48928);
xor U49041 (N_49041,N_48779,N_48836);
xnor U49042 (N_49042,N_48878,N_48992);
nand U49043 (N_49043,N_48893,N_48999);
xor U49044 (N_49044,N_48806,N_48987);
nor U49045 (N_49045,N_48782,N_48906);
or U49046 (N_49046,N_48774,N_48792);
and U49047 (N_49047,N_48997,N_48786);
and U49048 (N_49048,N_48818,N_48976);
and U49049 (N_49049,N_48958,N_48890);
or U49050 (N_49050,N_48816,N_48810);
nor U49051 (N_49051,N_48925,N_48924);
xnor U49052 (N_49052,N_48944,N_48820);
or U49053 (N_49053,N_48773,N_48914);
xnor U49054 (N_49054,N_48904,N_48989);
nor U49055 (N_49055,N_48942,N_48887);
nand U49056 (N_49056,N_48888,N_48874);
nand U49057 (N_49057,N_48940,N_48995);
xor U49058 (N_49058,N_48831,N_48897);
nor U49059 (N_49059,N_48998,N_48978);
and U49060 (N_49060,N_48929,N_48814);
or U49061 (N_49061,N_48975,N_48953);
nand U49062 (N_49062,N_48883,N_48974);
nor U49063 (N_49063,N_48803,N_48949);
nor U49064 (N_49064,N_48776,N_48896);
nand U49065 (N_49065,N_48927,N_48790);
xnor U49066 (N_49066,N_48909,N_48849);
nor U49067 (N_49067,N_48770,N_48842);
nand U49068 (N_49068,N_48809,N_48895);
and U49069 (N_49069,N_48817,N_48972);
and U49070 (N_49070,N_48926,N_48952);
or U49071 (N_49071,N_48977,N_48969);
nand U49072 (N_49072,N_48950,N_48941);
nor U49073 (N_49073,N_48880,N_48922);
nand U49074 (N_49074,N_48867,N_48931);
or U49075 (N_49075,N_48879,N_48828);
and U49076 (N_49076,N_48758,N_48892);
or U49077 (N_49077,N_48753,N_48937);
or U49078 (N_49078,N_48954,N_48884);
or U49079 (N_49079,N_48805,N_48848);
nand U49080 (N_49080,N_48993,N_48945);
nor U49081 (N_49081,N_48860,N_48811);
nand U49082 (N_49082,N_48869,N_48872);
xor U49083 (N_49083,N_48882,N_48851);
nand U49084 (N_49084,N_48798,N_48985);
and U49085 (N_49085,N_48837,N_48812);
nor U49086 (N_49086,N_48961,N_48756);
nor U49087 (N_49087,N_48823,N_48956);
and U49088 (N_49088,N_48856,N_48966);
nor U49089 (N_49089,N_48752,N_48923);
or U49090 (N_49090,N_48870,N_48807);
nor U49091 (N_49091,N_48825,N_48901);
or U49092 (N_49092,N_48751,N_48757);
or U49093 (N_49093,N_48864,N_48934);
or U49094 (N_49094,N_48868,N_48951);
xnor U49095 (N_49095,N_48754,N_48964);
nor U49096 (N_49096,N_48981,N_48832);
and U49097 (N_49097,N_48979,N_48984);
xor U49098 (N_49098,N_48830,N_48783);
xor U49099 (N_49099,N_48755,N_48778);
xnor U49100 (N_49100,N_48784,N_48788);
xor U49101 (N_49101,N_48785,N_48772);
and U49102 (N_49102,N_48858,N_48797);
xnor U49103 (N_49103,N_48841,N_48959);
or U49104 (N_49104,N_48866,N_48760);
and U49105 (N_49105,N_48957,N_48908);
or U49106 (N_49106,N_48857,N_48980);
nor U49107 (N_49107,N_48932,N_48946);
nand U49108 (N_49108,N_48789,N_48915);
or U49109 (N_49109,N_48921,N_48804);
nor U49110 (N_49110,N_48967,N_48827);
nor U49111 (N_49111,N_48829,N_48902);
and U49112 (N_49112,N_48794,N_48865);
xnor U49113 (N_49113,N_48903,N_48886);
nand U49114 (N_49114,N_48889,N_48846);
nand U49115 (N_49115,N_48875,N_48920);
nor U49116 (N_49116,N_48871,N_48955);
xnor U49117 (N_49117,N_48861,N_48815);
nand U49118 (N_49118,N_48988,N_48845);
xor U49119 (N_49119,N_48973,N_48759);
nand U49120 (N_49120,N_48821,N_48843);
nor U49121 (N_49121,N_48767,N_48899);
or U49122 (N_49122,N_48863,N_48802);
xor U49123 (N_49123,N_48768,N_48761);
xnor U49124 (N_49124,N_48781,N_48907);
or U49125 (N_49125,N_48901,N_48830);
nand U49126 (N_49126,N_48755,N_48952);
xor U49127 (N_49127,N_48968,N_48927);
xor U49128 (N_49128,N_48960,N_48851);
nand U49129 (N_49129,N_48948,N_48986);
nor U49130 (N_49130,N_48867,N_48846);
nor U49131 (N_49131,N_48946,N_48884);
or U49132 (N_49132,N_48776,N_48772);
xnor U49133 (N_49133,N_48893,N_48965);
and U49134 (N_49134,N_48886,N_48959);
xnor U49135 (N_49135,N_48941,N_48757);
and U49136 (N_49136,N_48764,N_48904);
xor U49137 (N_49137,N_48899,N_48975);
xnor U49138 (N_49138,N_48978,N_48789);
nor U49139 (N_49139,N_48983,N_48902);
nand U49140 (N_49140,N_48885,N_48796);
nor U49141 (N_49141,N_48974,N_48819);
nor U49142 (N_49142,N_48915,N_48867);
and U49143 (N_49143,N_48938,N_48759);
and U49144 (N_49144,N_48954,N_48804);
and U49145 (N_49145,N_48972,N_48992);
and U49146 (N_49146,N_48944,N_48847);
nor U49147 (N_49147,N_48983,N_48878);
or U49148 (N_49148,N_48865,N_48982);
xor U49149 (N_49149,N_48870,N_48886);
nand U49150 (N_49150,N_48932,N_48791);
xnor U49151 (N_49151,N_48751,N_48879);
xor U49152 (N_49152,N_48807,N_48848);
xor U49153 (N_49153,N_48906,N_48771);
xnor U49154 (N_49154,N_48875,N_48961);
nand U49155 (N_49155,N_48946,N_48993);
nand U49156 (N_49156,N_48794,N_48868);
nand U49157 (N_49157,N_48985,N_48780);
or U49158 (N_49158,N_48753,N_48955);
or U49159 (N_49159,N_48960,N_48816);
xnor U49160 (N_49160,N_48766,N_48813);
nand U49161 (N_49161,N_48940,N_48985);
nor U49162 (N_49162,N_48794,N_48783);
xnor U49163 (N_49163,N_48857,N_48908);
nor U49164 (N_49164,N_48777,N_48943);
or U49165 (N_49165,N_48905,N_48859);
nor U49166 (N_49166,N_48995,N_48751);
or U49167 (N_49167,N_48899,N_48820);
or U49168 (N_49168,N_48969,N_48825);
or U49169 (N_49169,N_48945,N_48831);
or U49170 (N_49170,N_48775,N_48857);
nor U49171 (N_49171,N_48886,N_48820);
or U49172 (N_49172,N_48781,N_48868);
or U49173 (N_49173,N_48958,N_48868);
nor U49174 (N_49174,N_48799,N_48808);
nor U49175 (N_49175,N_48800,N_48833);
nor U49176 (N_49176,N_48930,N_48945);
and U49177 (N_49177,N_48927,N_48912);
xor U49178 (N_49178,N_48884,N_48880);
or U49179 (N_49179,N_48815,N_48865);
and U49180 (N_49180,N_48824,N_48854);
or U49181 (N_49181,N_48923,N_48991);
or U49182 (N_49182,N_48971,N_48758);
xor U49183 (N_49183,N_48863,N_48953);
or U49184 (N_49184,N_48912,N_48898);
and U49185 (N_49185,N_48818,N_48773);
and U49186 (N_49186,N_48865,N_48808);
nor U49187 (N_49187,N_48799,N_48902);
and U49188 (N_49188,N_48840,N_48981);
and U49189 (N_49189,N_48818,N_48858);
or U49190 (N_49190,N_48828,N_48810);
xnor U49191 (N_49191,N_48881,N_48985);
xnor U49192 (N_49192,N_48829,N_48751);
or U49193 (N_49193,N_48889,N_48908);
or U49194 (N_49194,N_48766,N_48841);
nor U49195 (N_49195,N_48934,N_48822);
or U49196 (N_49196,N_48926,N_48810);
nor U49197 (N_49197,N_48871,N_48858);
or U49198 (N_49198,N_48755,N_48811);
and U49199 (N_49199,N_48973,N_48788);
nand U49200 (N_49200,N_48943,N_48870);
or U49201 (N_49201,N_48781,N_48931);
nand U49202 (N_49202,N_48798,N_48792);
nor U49203 (N_49203,N_48879,N_48961);
nand U49204 (N_49204,N_48980,N_48788);
and U49205 (N_49205,N_48871,N_48845);
and U49206 (N_49206,N_48955,N_48873);
nor U49207 (N_49207,N_48949,N_48924);
nand U49208 (N_49208,N_48781,N_48761);
nand U49209 (N_49209,N_48963,N_48796);
nand U49210 (N_49210,N_48826,N_48912);
and U49211 (N_49211,N_48814,N_48963);
and U49212 (N_49212,N_48845,N_48923);
or U49213 (N_49213,N_48859,N_48964);
nand U49214 (N_49214,N_48810,N_48940);
nand U49215 (N_49215,N_48905,N_48790);
or U49216 (N_49216,N_48756,N_48944);
xor U49217 (N_49217,N_48932,N_48973);
nand U49218 (N_49218,N_48793,N_48928);
and U49219 (N_49219,N_48879,N_48932);
or U49220 (N_49220,N_48870,N_48815);
xor U49221 (N_49221,N_48923,N_48807);
nand U49222 (N_49222,N_48750,N_48780);
xnor U49223 (N_49223,N_48774,N_48970);
nand U49224 (N_49224,N_48873,N_48845);
or U49225 (N_49225,N_48790,N_48808);
nand U49226 (N_49226,N_48811,N_48830);
xnor U49227 (N_49227,N_48862,N_48951);
and U49228 (N_49228,N_48756,N_48996);
xnor U49229 (N_49229,N_48982,N_48856);
and U49230 (N_49230,N_48769,N_48836);
xor U49231 (N_49231,N_48752,N_48972);
and U49232 (N_49232,N_48753,N_48959);
nand U49233 (N_49233,N_48929,N_48884);
xnor U49234 (N_49234,N_48959,N_48909);
and U49235 (N_49235,N_48845,N_48924);
nor U49236 (N_49236,N_48856,N_48899);
xor U49237 (N_49237,N_48889,N_48844);
nor U49238 (N_49238,N_48884,N_48791);
nand U49239 (N_49239,N_48906,N_48986);
nor U49240 (N_49240,N_48757,N_48957);
nor U49241 (N_49241,N_48908,N_48781);
xnor U49242 (N_49242,N_48814,N_48861);
xnor U49243 (N_49243,N_48870,N_48866);
nand U49244 (N_49244,N_48915,N_48820);
and U49245 (N_49245,N_48973,N_48857);
nand U49246 (N_49246,N_48805,N_48798);
nand U49247 (N_49247,N_48982,N_48750);
nand U49248 (N_49248,N_48917,N_48892);
xor U49249 (N_49249,N_48938,N_48906);
xnor U49250 (N_49250,N_49192,N_49049);
nand U49251 (N_49251,N_49052,N_49038);
nand U49252 (N_49252,N_49028,N_49200);
nand U49253 (N_49253,N_49187,N_49001);
xnor U49254 (N_49254,N_49220,N_49176);
or U49255 (N_49255,N_49046,N_49058);
or U49256 (N_49256,N_49054,N_49122);
nor U49257 (N_49257,N_49033,N_49068);
and U49258 (N_49258,N_49152,N_49197);
nor U49259 (N_49259,N_49130,N_49199);
nand U49260 (N_49260,N_49036,N_49222);
nor U49261 (N_49261,N_49237,N_49006);
and U49262 (N_49262,N_49171,N_49218);
and U49263 (N_49263,N_49047,N_49208);
nor U49264 (N_49264,N_49243,N_49221);
or U49265 (N_49265,N_49149,N_49075);
xor U49266 (N_49266,N_49190,N_49105);
nand U49267 (N_49267,N_49037,N_49183);
nand U49268 (N_49268,N_49115,N_49048);
nand U49269 (N_49269,N_49085,N_49113);
xor U49270 (N_49270,N_49163,N_49029);
and U49271 (N_49271,N_49186,N_49181);
and U49272 (N_49272,N_49024,N_49018);
and U49273 (N_49273,N_49177,N_49012);
nand U49274 (N_49274,N_49219,N_49155);
xor U49275 (N_49275,N_49193,N_49069);
and U49276 (N_49276,N_49030,N_49143);
or U49277 (N_49277,N_49232,N_49245);
nor U49278 (N_49278,N_49051,N_49227);
and U49279 (N_49279,N_49156,N_49019);
nor U49280 (N_49280,N_49229,N_49242);
xnor U49281 (N_49281,N_49191,N_49008);
xor U49282 (N_49282,N_49248,N_49147);
and U49283 (N_49283,N_49158,N_49166);
or U49284 (N_49284,N_49127,N_49040);
nor U49285 (N_49285,N_49133,N_49150);
xnor U49286 (N_49286,N_49060,N_49080);
and U49287 (N_49287,N_49004,N_49076);
nand U49288 (N_49288,N_49139,N_49043);
xnor U49289 (N_49289,N_49223,N_49022);
xnor U49290 (N_49290,N_49074,N_49111);
nor U49291 (N_49291,N_49185,N_49057);
or U49292 (N_49292,N_49198,N_49135);
nor U49293 (N_49293,N_49121,N_49228);
nor U49294 (N_49294,N_49134,N_49096);
and U49295 (N_49295,N_49234,N_49039);
nand U49296 (N_49296,N_49138,N_49102);
and U49297 (N_49297,N_49165,N_49194);
nand U49298 (N_49298,N_49010,N_49050);
or U49299 (N_49299,N_49117,N_49009);
nor U49300 (N_49300,N_49241,N_49086);
and U49301 (N_49301,N_49173,N_49097);
nor U49302 (N_49302,N_49116,N_49065);
nand U49303 (N_49303,N_49114,N_49209);
and U49304 (N_49304,N_49083,N_49240);
nand U49305 (N_49305,N_49178,N_49126);
xnor U49306 (N_49306,N_49045,N_49168);
xor U49307 (N_49307,N_49109,N_49099);
and U49308 (N_49308,N_49002,N_49140);
or U49309 (N_49309,N_49160,N_49095);
xor U49310 (N_49310,N_49124,N_49182);
xor U49311 (N_49311,N_49169,N_49106);
nand U49312 (N_49312,N_49180,N_49053);
or U49313 (N_49313,N_49128,N_49204);
or U49314 (N_49314,N_49094,N_49247);
and U49315 (N_49315,N_49013,N_49077);
nor U49316 (N_49316,N_49132,N_49091);
nand U49317 (N_49317,N_49017,N_49161);
or U49318 (N_49318,N_49172,N_49101);
nor U49319 (N_49319,N_49201,N_49151);
nand U49320 (N_49320,N_49020,N_49144);
and U49321 (N_49321,N_49062,N_49202);
nand U49322 (N_49322,N_49066,N_49023);
or U49323 (N_49323,N_49104,N_49196);
xnor U49324 (N_49324,N_49112,N_49032);
or U49325 (N_49325,N_49000,N_49103);
and U49326 (N_49326,N_49189,N_49210);
xor U49327 (N_49327,N_49146,N_49215);
xnor U49328 (N_49328,N_49175,N_49107);
nor U49329 (N_49329,N_49061,N_49225);
xnor U49330 (N_49330,N_49031,N_49063);
nor U49331 (N_49331,N_49005,N_49011);
and U49332 (N_49332,N_49174,N_49067);
nand U49333 (N_49333,N_49082,N_49081);
nand U49334 (N_49334,N_49213,N_49016);
nor U49335 (N_49335,N_49238,N_49188);
xor U49336 (N_49336,N_49071,N_49145);
xor U49337 (N_49337,N_49233,N_49136);
nand U49338 (N_49338,N_49206,N_49170);
and U49339 (N_49339,N_49044,N_49093);
xor U49340 (N_49340,N_49129,N_49021);
or U49341 (N_49341,N_49217,N_49056);
or U49342 (N_49342,N_49110,N_49137);
nand U49343 (N_49343,N_49098,N_49131);
xnor U49344 (N_49344,N_49087,N_49153);
xnor U49345 (N_49345,N_49035,N_49236);
nand U49346 (N_49346,N_49239,N_49142);
and U49347 (N_49347,N_49205,N_49090);
xnor U49348 (N_49348,N_49230,N_49154);
nor U49349 (N_49349,N_49207,N_49118);
nor U49350 (N_49350,N_49064,N_49100);
nand U49351 (N_49351,N_49141,N_49212);
xnor U49352 (N_49352,N_49148,N_49157);
and U49353 (N_49353,N_49108,N_49184);
xor U49354 (N_49354,N_49072,N_49027);
and U49355 (N_49355,N_49179,N_49007);
nor U49356 (N_49356,N_49078,N_49235);
nand U49357 (N_49357,N_49092,N_49014);
or U49358 (N_49358,N_49159,N_49231);
nand U49359 (N_49359,N_49226,N_49123);
xnor U49360 (N_49360,N_49089,N_49120);
nand U49361 (N_49361,N_49079,N_49015);
nor U49362 (N_49362,N_49055,N_49244);
and U49363 (N_49363,N_49119,N_49026);
nor U49364 (N_49364,N_49088,N_49167);
xnor U49365 (N_49365,N_49214,N_49003);
nand U49366 (N_49366,N_49034,N_49084);
and U49367 (N_49367,N_49162,N_49025);
and U49368 (N_49368,N_49249,N_49042);
nor U49369 (N_49369,N_49070,N_49073);
or U49370 (N_49370,N_49211,N_49125);
nor U49371 (N_49371,N_49203,N_49216);
and U49372 (N_49372,N_49059,N_49224);
and U49373 (N_49373,N_49195,N_49164);
nor U49374 (N_49374,N_49041,N_49246);
and U49375 (N_49375,N_49021,N_49026);
xnor U49376 (N_49376,N_49040,N_49111);
and U49377 (N_49377,N_49032,N_49109);
and U49378 (N_49378,N_49002,N_49193);
nand U49379 (N_49379,N_49007,N_49017);
nor U49380 (N_49380,N_49092,N_49232);
and U49381 (N_49381,N_49071,N_49023);
nor U49382 (N_49382,N_49151,N_49135);
nand U49383 (N_49383,N_49238,N_49231);
nor U49384 (N_49384,N_49137,N_49023);
xnor U49385 (N_49385,N_49234,N_49228);
nand U49386 (N_49386,N_49001,N_49089);
nand U49387 (N_49387,N_49210,N_49018);
and U49388 (N_49388,N_49228,N_49147);
and U49389 (N_49389,N_49028,N_49148);
nand U49390 (N_49390,N_49171,N_49240);
nor U49391 (N_49391,N_49071,N_49246);
nand U49392 (N_49392,N_49238,N_49113);
or U49393 (N_49393,N_49069,N_49175);
nor U49394 (N_49394,N_49198,N_49162);
nor U49395 (N_49395,N_49073,N_49138);
xnor U49396 (N_49396,N_49134,N_49131);
xnor U49397 (N_49397,N_49097,N_49088);
nand U49398 (N_49398,N_49109,N_49152);
xnor U49399 (N_49399,N_49036,N_49107);
nor U49400 (N_49400,N_49149,N_49030);
and U49401 (N_49401,N_49012,N_49154);
or U49402 (N_49402,N_49030,N_49132);
xor U49403 (N_49403,N_49058,N_49042);
and U49404 (N_49404,N_49220,N_49058);
and U49405 (N_49405,N_49226,N_49026);
and U49406 (N_49406,N_49047,N_49018);
xor U49407 (N_49407,N_49111,N_49173);
or U49408 (N_49408,N_49193,N_49221);
nand U49409 (N_49409,N_49224,N_49219);
or U49410 (N_49410,N_49179,N_49188);
nor U49411 (N_49411,N_49103,N_49084);
or U49412 (N_49412,N_49063,N_49126);
or U49413 (N_49413,N_49147,N_49237);
or U49414 (N_49414,N_49156,N_49185);
nor U49415 (N_49415,N_49213,N_49132);
or U49416 (N_49416,N_49137,N_49174);
and U49417 (N_49417,N_49087,N_49110);
nand U49418 (N_49418,N_49084,N_49068);
or U49419 (N_49419,N_49211,N_49068);
nor U49420 (N_49420,N_49075,N_49156);
nand U49421 (N_49421,N_49248,N_49235);
xnor U49422 (N_49422,N_49029,N_49011);
or U49423 (N_49423,N_49152,N_49249);
xor U49424 (N_49424,N_49067,N_49081);
or U49425 (N_49425,N_49073,N_49204);
nand U49426 (N_49426,N_49160,N_49238);
and U49427 (N_49427,N_49141,N_49055);
xnor U49428 (N_49428,N_49109,N_49227);
nor U49429 (N_49429,N_49029,N_49244);
xor U49430 (N_49430,N_49189,N_49092);
nand U49431 (N_49431,N_49216,N_49193);
and U49432 (N_49432,N_49152,N_49203);
or U49433 (N_49433,N_49180,N_49141);
and U49434 (N_49434,N_49163,N_49083);
and U49435 (N_49435,N_49007,N_49238);
and U49436 (N_49436,N_49093,N_49034);
xor U49437 (N_49437,N_49147,N_49171);
nor U49438 (N_49438,N_49020,N_49171);
xor U49439 (N_49439,N_49039,N_49000);
xor U49440 (N_49440,N_49218,N_49074);
and U49441 (N_49441,N_49211,N_49167);
nand U49442 (N_49442,N_49090,N_49155);
xor U49443 (N_49443,N_49103,N_49045);
or U49444 (N_49444,N_49243,N_49181);
xnor U49445 (N_49445,N_49217,N_49165);
nor U49446 (N_49446,N_49171,N_49146);
nand U49447 (N_49447,N_49067,N_49017);
or U49448 (N_49448,N_49174,N_49046);
xnor U49449 (N_49449,N_49144,N_49069);
nand U49450 (N_49450,N_49228,N_49106);
and U49451 (N_49451,N_49119,N_49139);
or U49452 (N_49452,N_49090,N_49006);
or U49453 (N_49453,N_49110,N_49194);
xor U49454 (N_49454,N_49001,N_49116);
and U49455 (N_49455,N_49008,N_49028);
xnor U49456 (N_49456,N_49171,N_49045);
and U49457 (N_49457,N_49106,N_49115);
or U49458 (N_49458,N_49038,N_49101);
nor U49459 (N_49459,N_49129,N_49172);
xnor U49460 (N_49460,N_49219,N_49196);
nor U49461 (N_49461,N_49225,N_49152);
and U49462 (N_49462,N_49220,N_49175);
xnor U49463 (N_49463,N_49198,N_49212);
nand U49464 (N_49464,N_49238,N_49240);
or U49465 (N_49465,N_49098,N_49096);
and U49466 (N_49466,N_49127,N_49184);
nor U49467 (N_49467,N_49026,N_49044);
nand U49468 (N_49468,N_49053,N_49016);
nand U49469 (N_49469,N_49026,N_49033);
and U49470 (N_49470,N_49023,N_49029);
and U49471 (N_49471,N_49208,N_49127);
nand U49472 (N_49472,N_49174,N_49148);
nand U49473 (N_49473,N_49152,N_49015);
nor U49474 (N_49474,N_49112,N_49050);
nor U49475 (N_49475,N_49034,N_49204);
and U49476 (N_49476,N_49039,N_49018);
or U49477 (N_49477,N_49049,N_49212);
and U49478 (N_49478,N_49066,N_49022);
or U49479 (N_49479,N_49243,N_49120);
nand U49480 (N_49480,N_49075,N_49001);
or U49481 (N_49481,N_49047,N_49120);
xnor U49482 (N_49482,N_49132,N_49225);
nor U49483 (N_49483,N_49198,N_49159);
xnor U49484 (N_49484,N_49107,N_49206);
nand U49485 (N_49485,N_49242,N_49130);
nor U49486 (N_49486,N_49077,N_49151);
or U49487 (N_49487,N_49005,N_49057);
nand U49488 (N_49488,N_49148,N_49064);
and U49489 (N_49489,N_49208,N_49109);
and U49490 (N_49490,N_49084,N_49018);
xor U49491 (N_49491,N_49098,N_49073);
and U49492 (N_49492,N_49142,N_49146);
xor U49493 (N_49493,N_49222,N_49246);
and U49494 (N_49494,N_49196,N_49113);
and U49495 (N_49495,N_49011,N_49244);
or U49496 (N_49496,N_49131,N_49018);
xor U49497 (N_49497,N_49063,N_49034);
nand U49498 (N_49498,N_49202,N_49004);
nor U49499 (N_49499,N_49055,N_49124);
or U49500 (N_49500,N_49415,N_49485);
xor U49501 (N_49501,N_49388,N_49286);
nand U49502 (N_49502,N_49253,N_49431);
xor U49503 (N_49503,N_49397,N_49296);
nor U49504 (N_49504,N_49292,N_49479);
nor U49505 (N_49505,N_49260,N_49288);
or U49506 (N_49506,N_49449,N_49360);
nor U49507 (N_49507,N_49314,N_49337);
xor U49508 (N_49508,N_49311,N_49460);
nor U49509 (N_49509,N_49406,N_49313);
or U49510 (N_49510,N_49328,N_49250);
nand U49511 (N_49511,N_49486,N_49488);
and U49512 (N_49512,N_49496,N_49299);
xor U49513 (N_49513,N_49257,N_49374);
nand U49514 (N_49514,N_49394,N_49342);
and U49515 (N_49515,N_49282,N_49295);
nor U49516 (N_49516,N_49421,N_49484);
or U49517 (N_49517,N_49437,N_49335);
or U49518 (N_49518,N_49381,N_49396);
and U49519 (N_49519,N_49489,N_49266);
nor U49520 (N_49520,N_49316,N_49472);
or U49521 (N_49521,N_49482,N_49344);
or U49522 (N_49522,N_49332,N_49252);
nor U49523 (N_49523,N_49317,N_49474);
and U49524 (N_49524,N_49309,N_49445);
and U49525 (N_49525,N_49259,N_49270);
xnor U49526 (N_49526,N_49410,N_49477);
or U49527 (N_49527,N_49346,N_49458);
xor U49528 (N_49528,N_49379,N_49436);
nand U49529 (N_49529,N_49378,N_49354);
xnor U49530 (N_49530,N_49255,N_49340);
and U49531 (N_49531,N_49461,N_49305);
nand U49532 (N_49532,N_49476,N_49447);
nor U49533 (N_49533,N_49256,N_49352);
nor U49534 (N_49534,N_49365,N_49369);
nand U49535 (N_49535,N_49363,N_49450);
or U49536 (N_49536,N_49425,N_49469);
xor U49537 (N_49537,N_49339,N_49426);
or U49538 (N_49538,N_49376,N_49399);
and U49539 (N_49539,N_49446,N_49412);
and U49540 (N_49540,N_49383,N_49251);
xor U49541 (N_49541,N_49326,N_49261);
nand U49542 (N_49542,N_49366,N_49343);
xnor U49543 (N_49543,N_49275,N_49478);
nor U49544 (N_49544,N_49320,N_49432);
nand U49545 (N_49545,N_49416,N_49293);
xnor U49546 (N_49546,N_49278,N_49407);
or U49547 (N_49547,N_49404,N_49429);
or U49548 (N_49548,N_49440,N_49418);
and U49549 (N_49549,N_49338,N_49439);
nor U49550 (N_49550,N_49254,N_49468);
or U49551 (N_49551,N_49303,N_49327);
or U49552 (N_49552,N_49398,N_49465);
or U49553 (N_49553,N_49463,N_49427);
xnor U49554 (N_49554,N_49464,N_49393);
xor U49555 (N_49555,N_49308,N_49443);
nand U49556 (N_49556,N_49280,N_49359);
xor U49557 (N_49557,N_49413,N_49435);
and U49558 (N_49558,N_49492,N_49321);
or U49559 (N_49559,N_49298,N_49297);
or U49560 (N_49560,N_49263,N_49470);
xnor U49561 (N_49561,N_49487,N_49361);
xor U49562 (N_49562,N_49294,N_49276);
and U49563 (N_49563,N_49301,N_49371);
nand U49564 (N_49564,N_49457,N_49353);
and U49565 (N_49565,N_49385,N_49284);
xor U49566 (N_49566,N_49265,N_49409);
nand U49567 (N_49567,N_49264,N_49258);
nor U49568 (N_49568,N_49331,N_49430);
and U49569 (N_49569,N_49370,N_49362);
and U49570 (N_49570,N_49373,N_49355);
and U49571 (N_49571,N_49389,N_49411);
nand U49572 (N_49572,N_49467,N_49315);
nand U49573 (N_49573,N_49341,N_49333);
xor U49574 (N_49574,N_49456,N_49272);
and U49575 (N_49575,N_49330,N_49455);
or U49576 (N_49576,N_49358,N_49277);
xnor U49577 (N_49577,N_49279,N_49438);
xnor U49578 (N_49578,N_49312,N_49310);
xnor U49579 (N_49579,N_49267,N_49364);
nand U49580 (N_49580,N_49300,N_49377);
xor U49581 (N_49581,N_49356,N_49307);
nand U49582 (N_49582,N_49483,N_49375);
xor U49583 (N_49583,N_49382,N_49471);
nand U49584 (N_49584,N_49268,N_49283);
xor U49585 (N_49585,N_49290,N_49281);
xnor U49586 (N_49586,N_49451,N_49387);
nor U49587 (N_49587,N_49490,N_49448);
nand U49588 (N_49588,N_49481,N_49420);
nor U49589 (N_49589,N_49271,N_49304);
nor U49590 (N_49590,N_49499,N_49306);
or U49591 (N_49591,N_49324,N_49274);
nand U49592 (N_49592,N_49414,N_49493);
xnor U49593 (N_49593,N_49494,N_49480);
nand U49594 (N_49594,N_49424,N_49495);
and U49595 (N_49595,N_49401,N_49269);
or U49596 (N_49596,N_49302,N_49405);
and U49597 (N_49597,N_49462,N_49386);
and U49598 (N_49598,N_49318,N_49289);
nand U49599 (N_49599,N_49395,N_49403);
nand U49600 (N_49600,N_49287,N_49349);
and U49601 (N_49601,N_49444,N_49345);
nor U49602 (N_49602,N_49441,N_49475);
xor U49603 (N_49603,N_49473,N_49336);
and U49604 (N_49604,N_49422,N_49498);
or U49605 (N_49605,N_49319,N_49417);
nand U49606 (N_49606,N_49497,N_49368);
and U49607 (N_49607,N_49434,N_49428);
xor U49608 (N_49608,N_49350,N_49367);
nand U49609 (N_49609,N_49453,N_49348);
nor U49610 (N_49610,N_49322,N_49391);
or U49611 (N_49611,N_49262,N_49459);
xor U49612 (N_49612,N_49384,N_49452);
nor U49613 (N_49613,N_49273,N_49372);
and U49614 (N_49614,N_49380,N_49491);
nand U49615 (N_49615,N_49433,N_49347);
nand U49616 (N_49616,N_49423,N_49402);
or U49617 (N_49617,N_49329,N_49325);
or U49618 (N_49618,N_49390,N_49408);
nand U49619 (N_49619,N_49442,N_49454);
xnor U49620 (N_49620,N_49357,N_49351);
nand U49621 (N_49621,N_49291,N_49323);
xor U49622 (N_49622,N_49285,N_49466);
xnor U49623 (N_49623,N_49400,N_49392);
xnor U49624 (N_49624,N_49419,N_49334);
or U49625 (N_49625,N_49373,N_49406);
nor U49626 (N_49626,N_49313,N_49426);
nor U49627 (N_49627,N_49308,N_49330);
or U49628 (N_49628,N_49281,N_49498);
xnor U49629 (N_49629,N_49428,N_49420);
or U49630 (N_49630,N_49293,N_49258);
and U49631 (N_49631,N_49433,N_49354);
nor U49632 (N_49632,N_49381,N_49378);
and U49633 (N_49633,N_49369,N_49430);
xor U49634 (N_49634,N_49327,N_49328);
nand U49635 (N_49635,N_49380,N_49317);
nand U49636 (N_49636,N_49465,N_49321);
xor U49637 (N_49637,N_49293,N_49420);
or U49638 (N_49638,N_49399,N_49289);
nor U49639 (N_49639,N_49483,N_49332);
xor U49640 (N_49640,N_49331,N_49344);
or U49641 (N_49641,N_49465,N_49274);
xnor U49642 (N_49642,N_49384,N_49413);
nand U49643 (N_49643,N_49467,N_49280);
nand U49644 (N_49644,N_49473,N_49458);
nand U49645 (N_49645,N_49449,N_49451);
nor U49646 (N_49646,N_49391,N_49401);
or U49647 (N_49647,N_49342,N_49316);
nor U49648 (N_49648,N_49394,N_49298);
xor U49649 (N_49649,N_49311,N_49321);
and U49650 (N_49650,N_49369,N_49472);
nand U49651 (N_49651,N_49325,N_49321);
nand U49652 (N_49652,N_49356,N_49391);
and U49653 (N_49653,N_49307,N_49447);
or U49654 (N_49654,N_49258,N_49288);
nand U49655 (N_49655,N_49320,N_49463);
nor U49656 (N_49656,N_49463,N_49457);
or U49657 (N_49657,N_49275,N_49330);
or U49658 (N_49658,N_49345,N_49294);
or U49659 (N_49659,N_49424,N_49311);
xnor U49660 (N_49660,N_49284,N_49281);
or U49661 (N_49661,N_49436,N_49456);
and U49662 (N_49662,N_49409,N_49454);
nor U49663 (N_49663,N_49432,N_49413);
xnor U49664 (N_49664,N_49488,N_49465);
nand U49665 (N_49665,N_49381,N_49285);
nand U49666 (N_49666,N_49331,N_49432);
and U49667 (N_49667,N_49262,N_49393);
xor U49668 (N_49668,N_49347,N_49480);
nand U49669 (N_49669,N_49497,N_49434);
and U49670 (N_49670,N_49458,N_49438);
or U49671 (N_49671,N_49455,N_49394);
or U49672 (N_49672,N_49308,N_49268);
nand U49673 (N_49673,N_49423,N_49327);
nand U49674 (N_49674,N_49416,N_49363);
or U49675 (N_49675,N_49400,N_49314);
nand U49676 (N_49676,N_49351,N_49480);
nand U49677 (N_49677,N_49273,N_49284);
or U49678 (N_49678,N_49388,N_49315);
and U49679 (N_49679,N_49354,N_49426);
and U49680 (N_49680,N_49308,N_49470);
nand U49681 (N_49681,N_49262,N_49414);
nor U49682 (N_49682,N_49328,N_49300);
and U49683 (N_49683,N_49344,N_49476);
nand U49684 (N_49684,N_49459,N_49369);
nand U49685 (N_49685,N_49264,N_49287);
or U49686 (N_49686,N_49425,N_49291);
xnor U49687 (N_49687,N_49260,N_49390);
or U49688 (N_49688,N_49457,N_49320);
nor U49689 (N_49689,N_49270,N_49368);
xnor U49690 (N_49690,N_49346,N_49324);
nor U49691 (N_49691,N_49337,N_49305);
and U49692 (N_49692,N_49490,N_49427);
nor U49693 (N_49693,N_49298,N_49268);
nand U49694 (N_49694,N_49298,N_49318);
or U49695 (N_49695,N_49332,N_49426);
xor U49696 (N_49696,N_49492,N_49425);
and U49697 (N_49697,N_49421,N_49462);
or U49698 (N_49698,N_49313,N_49270);
xnor U49699 (N_49699,N_49257,N_49480);
and U49700 (N_49700,N_49442,N_49251);
and U49701 (N_49701,N_49389,N_49396);
xor U49702 (N_49702,N_49309,N_49277);
nor U49703 (N_49703,N_49476,N_49286);
and U49704 (N_49704,N_49293,N_49386);
nand U49705 (N_49705,N_49319,N_49356);
nor U49706 (N_49706,N_49267,N_49340);
and U49707 (N_49707,N_49271,N_49490);
nor U49708 (N_49708,N_49284,N_49323);
and U49709 (N_49709,N_49274,N_49323);
or U49710 (N_49710,N_49369,N_49438);
nor U49711 (N_49711,N_49345,N_49392);
or U49712 (N_49712,N_49483,N_49308);
nor U49713 (N_49713,N_49485,N_49368);
and U49714 (N_49714,N_49463,N_49359);
nand U49715 (N_49715,N_49351,N_49317);
and U49716 (N_49716,N_49371,N_49446);
nand U49717 (N_49717,N_49341,N_49364);
or U49718 (N_49718,N_49282,N_49494);
nand U49719 (N_49719,N_49281,N_49367);
nand U49720 (N_49720,N_49358,N_49326);
nor U49721 (N_49721,N_49301,N_49468);
or U49722 (N_49722,N_49259,N_49266);
xor U49723 (N_49723,N_49305,N_49398);
nor U49724 (N_49724,N_49333,N_49423);
nor U49725 (N_49725,N_49490,N_49442);
or U49726 (N_49726,N_49434,N_49328);
and U49727 (N_49727,N_49422,N_49337);
xnor U49728 (N_49728,N_49301,N_49335);
and U49729 (N_49729,N_49261,N_49476);
and U49730 (N_49730,N_49408,N_49496);
nor U49731 (N_49731,N_49446,N_49482);
and U49732 (N_49732,N_49447,N_49289);
xnor U49733 (N_49733,N_49371,N_49452);
and U49734 (N_49734,N_49448,N_49429);
or U49735 (N_49735,N_49262,N_49477);
nor U49736 (N_49736,N_49444,N_49469);
nor U49737 (N_49737,N_49270,N_49492);
nor U49738 (N_49738,N_49459,N_49385);
or U49739 (N_49739,N_49357,N_49282);
or U49740 (N_49740,N_49295,N_49362);
nor U49741 (N_49741,N_49288,N_49445);
or U49742 (N_49742,N_49328,N_49485);
xnor U49743 (N_49743,N_49428,N_49450);
nor U49744 (N_49744,N_49324,N_49393);
nor U49745 (N_49745,N_49335,N_49377);
nand U49746 (N_49746,N_49368,N_49369);
nor U49747 (N_49747,N_49382,N_49365);
xor U49748 (N_49748,N_49364,N_49316);
xor U49749 (N_49749,N_49470,N_49440);
nand U49750 (N_49750,N_49692,N_49737);
and U49751 (N_49751,N_49508,N_49687);
xnor U49752 (N_49752,N_49583,N_49728);
nand U49753 (N_49753,N_49559,N_49614);
and U49754 (N_49754,N_49665,N_49732);
and U49755 (N_49755,N_49661,N_49538);
nor U49756 (N_49756,N_49669,N_49564);
or U49757 (N_49757,N_49719,N_49700);
and U49758 (N_49758,N_49552,N_49549);
nor U49759 (N_49759,N_49602,N_49546);
nor U49760 (N_49760,N_49748,N_49528);
or U49761 (N_49761,N_49634,N_49683);
nand U49762 (N_49762,N_49580,N_49658);
xnor U49763 (N_49763,N_49560,N_49671);
or U49764 (N_49764,N_49697,N_49739);
nor U49765 (N_49765,N_49746,N_49749);
xor U49766 (N_49766,N_49734,N_49736);
nand U49767 (N_49767,N_49677,N_49695);
nand U49768 (N_49768,N_49591,N_49500);
nor U49769 (N_49769,N_49711,N_49523);
and U49770 (N_49770,N_49578,N_49557);
xor U49771 (N_49771,N_49551,N_49513);
and U49772 (N_49772,N_49655,N_49527);
and U49773 (N_49773,N_49521,N_49590);
xor U49774 (N_49774,N_49539,N_49621);
nor U49775 (N_49775,N_49526,N_49550);
xnor U49776 (N_49776,N_49558,N_49686);
nor U49777 (N_49777,N_49660,N_49609);
and U49778 (N_49778,N_49627,N_49678);
nand U49779 (N_49779,N_49653,N_49745);
xor U49780 (N_49780,N_49588,N_49501);
xor U49781 (N_49781,N_49503,N_49544);
nor U49782 (N_49782,N_49600,N_49702);
nand U49783 (N_49783,N_49607,N_49531);
nor U49784 (N_49784,N_49515,N_49703);
nor U49785 (N_49785,N_49708,N_49646);
nand U49786 (N_49786,N_49547,N_49636);
xor U49787 (N_49787,N_49645,N_49622);
nor U49788 (N_49788,N_49718,N_49545);
xor U49789 (N_49789,N_49667,N_49596);
and U49790 (N_49790,N_49524,N_49530);
and U49791 (N_49791,N_49556,N_49720);
nor U49792 (N_49792,N_49509,N_49715);
nand U49793 (N_49793,N_49670,N_49575);
nor U49794 (N_49794,N_49642,N_49599);
and U49795 (N_49795,N_49688,N_49684);
and U49796 (N_49796,N_49594,N_49555);
or U49797 (N_49797,N_49504,N_49685);
or U49798 (N_49798,N_49632,N_49561);
xnor U49799 (N_49799,N_49593,N_49512);
xnor U49800 (N_49800,N_49741,N_49704);
xor U49801 (N_49801,N_49525,N_49535);
or U49802 (N_49802,N_49743,N_49542);
xor U49803 (N_49803,N_49666,N_49735);
xor U49804 (N_49804,N_49554,N_49656);
nand U49805 (N_49805,N_49694,N_49563);
or U49806 (N_49806,N_49540,N_49568);
and U49807 (N_49807,N_49681,N_49592);
nor U49808 (N_49808,N_49682,N_49566);
or U49809 (N_49809,N_49582,N_49630);
or U49810 (N_49810,N_49680,N_49603);
nor U49811 (N_49811,N_49618,N_49572);
nor U49812 (N_49812,N_49586,N_49733);
nand U49813 (N_49813,N_49543,N_49577);
nor U49814 (N_49814,N_49673,N_49714);
nand U49815 (N_49815,N_49725,N_49505);
nand U49816 (N_49816,N_49730,N_49571);
xor U49817 (N_49817,N_49519,N_49693);
or U49818 (N_49818,N_49699,N_49514);
nor U49819 (N_49819,N_49573,N_49637);
or U49820 (N_49820,N_49510,N_49705);
nand U49821 (N_49821,N_49713,N_49690);
nor U49822 (N_49822,N_49706,N_49529);
nand U49823 (N_49823,N_49631,N_49518);
nand U49824 (N_49824,N_49574,N_49663);
nor U49825 (N_49825,N_49724,N_49742);
nand U49826 (N_49826,N_49639,N_49701);
or U49827 (N_49827,N_49676,N_49659);
and U49828 (N_49828,N_49712,N_49640);
nand U49829 (N_49829,N_49541,N_49553);
xnor U49830 (N_49830,N_49726,N_49716);
xor U49831 (N_49831,N_49657,N_49643);
nand U49832 (N_49832,N_49598,N_49565);
or U49833 (N_49833,N_49721,N_49648);
or U49834 (N_49834,N_49585,N_49534);
nand U49835 (N_49835,N_49605,N_49604);
nor U49836 (N_49836,N_49517,N_49507);
nor U49837 (N_49837,N_49626,N_49520);
nor U49838 (N_49838,N_49717,N_49650);
nor U49839 (N_49839,N_49672,N_49511);
and U49840 (N_49840,N_49740,N_49709);
nor U49841 (N_49841,N_49579,N_49674);
xnor U49842 (N_49842,N_49710,N_49633);
and U49843 (N_49843,N_49731,N_49722);
nor U49844 (N_49844,N_49652,N_49584);
and U49845 (N_49845,N_49729,N_49615);
nor U49846 (N_49846,N_49562,N_49635);
xnor U49847 (N_49847,N_49625,N_49723);
xor U49848 (N_49848,N_49654,N_49506);
and U49849 (N_49849,N_49589,N_49619);
xor U49850 (N_49850,N_49668,N_49610);
or U49851 (N_49851,N_49698,N_49502);
nand U49852 (N_49852,N_49533,N_49747);
or U49853 (N_49853,N_49597,N_49649);
or U49854 (N_49854,N_49617,N_49576);
and U49855 (N_49855,N_49532,N_49570);
or U49856 (N_49856,N_49612,N_49624);
and U49857 (N_49857,N_49581,N_49623);
nor U49858 (N_49858,N_49522,N_49644);
xnor U49859 (N_49859,N_49569,N_49606);
or U49860 (N_49860,N_49616,N_49638);
nor U49861 (N_49861,N_49679,N_49587);
xor U49862 (N_49862,N_49675,N_49744);
nor U49863 (N_49863,N_49738,N_49727);
nand U49864 (N_49864,N_49707,N_49611);
xor U49865 (N_49865,N_49613,N_49548);
or U49866 (N_49866,N_49689,N_49641);
or U49867 (N_49867,N_49620,N_49595);
xnor U49868 (N_49868,N_49647,N_49691);
nand U49869 (N_49869,N_49628,N_49651);
and U49870 (N_49870,N_49608,N_49536);
and U49871 (N_49871,N_49664,N_49516);
xnor U49872 (N_49872,N_49662,N_49629);
nor U49873 (N_49873,N_49567,N_49537);
xnor U49874 (N_49874,N_49696,N_49601);
or U49875 (N_49875,N_49636,N_49536);
nor U49876 (N_49876,N_49611,N_49733);
xor U49877 (N_49877,N_49535,N_49749);
nand U49878 (N_49878,N_49532,N_49574);
nand U49879 (N_49879,N_49714,N_49651);
or U49880 (N_49880,N_49510,N_49583);
and U49881 (N_49881,N_49513,N_49665);
nor U49882 (N_49882,N_49548,N_49629);
or U49883 (N_49883,N_49694,N_49749);
nand U49884 (N_49884,N_49532,N_49530);
xnor U49885 (N_49885,N_49522,N_49729);
or U49886 (N_49886,N_49702,N_49598);
nor U49887 (N_49887,N_49738,N_49679);
nand U49888 (N_49888,N_49598,N_49520);
or U49889 (N_49889,N_49607,N_49635);
nor U49890 (N_49890,N_49603,N_49608);
nor U49891 (N_49891,N_49573,N_49537);
and U49892 (N_49892,N_49601,N_49665);
and U49893 (N_49893,N_49516,N_49537);
nand U49894 (N_49894,N_49572,N_49709);
nand U49895 (N_49895,N_49636,N_49710);
nand U49896 (N_49896,N_49650,N_49632);
nor U49897 (N_49897,N_49642,N_49506);
and U49898 (N_49898,N_49699,N_49701);
nand U49899 (N_49899,N_49659,N_49610);
or U49900 (N_49900,N_49620,N_49512);
nand U49901 (N_49901,N_49581,N_49727);
nand U49902 (N_49902,N_49561,N_49572);
nor U49903 (N_49903,N_49585,N_49555);
nand U49904 (N_49904,N_49723,N_49504);
nor U49905 (N_49905,N_49719,N_49536);
and U49906 (N_49906,N_49642,N_49539);
or U49907 (N_49907,N_49614,N_49608);
and U49908 (N_49908,N_49666,N_49701);
or U49909 (N_49909,N_49603,N_49510);
or U49910 (N_49910,N_49690,N_49562);
nand U49911 (N_49911,N_49583,N_49737);
and U49912 (N_49912,N_49619,N_49540);
nand U49913 (N_49913,N_49519,N_49516);
or U49914 (N_49914,N_49593,N_49659);
and U49915 (N_49915,N_49503,N_49678);
nor U49916 (N_49916,N_49580,N_49557);
or U49917 (N_49917,N_49566,N_49509);
nand U49918 (N_49918,N_49539,N_49657);
and U49919 (N_49919,N_49704,N_49715);
nand U49920 (N_49920,N_49580,N_49500);
xnor U49921 (N_49921,N_49734,N_49745);
and U49922 (N_49922,N_49614,N_49535);
xnor U49923 (N_49923,N_49603,N_49656);
and U49924 (N_49924,N_49629,N_49746);
and U49925 (N_49925,N_49628,N_49652);
or U49926 (N_49926,N_49737,N_49684);
nand U49927 (N_49927,N_49673,N_49747);
nor U49928 (N_49928,N_49698,N_49741);
xnor U49929 (N_49929,N_49511,N_49548);
and U49930 (N_49930,N_49617,N_49605);
nand U49931 (N_49931,N_49701,N_49510);
nand U49932 (N_49932,N_49652,N_49588);
or U49933 (N_49933,N_49526,N_49707);
or U49934 (N_49934,N_49728,N_49512);
nor U49935 (N_49935,N_49523,N_49742);
or U49936 (N_49936,N_49575,N_49679);
xor U49937 (N_49937,N_49552,N_49649);
or U49938 (N_49938,N_49568,N_49543);
and U49939 (N_49939,N_49601,N_49572);
and U49940 (N_49940,N_49660,N_49506);
xnor U49941 (N_49941,N_49629,N_49708);
and U49942 (N_49942,N_49748,N_49556);
nor U49943 (N_49943,N_49553,N_49669);
nand U49944 (N_49944,N_49531,N_49662);
nand U49945 (N_49945,N_49724,N_49532);
or U49946 (N_49946,N_49503,N_49661);
and U49947 (N_49947,N_49607,N_49637);
and U49948 (N_49948,N_49579,N_49598);
or U49949 (N_49949,N_49580,N_49726);
xor U49950 (N_49950,N_49673,N_49641);
nor U49951 (N_49951,N_49731,N_49680);
xnor U49952 (N_49952,N_49595,N_49583);
nand U49953 (N_49953,N_49519,N_49555);
and U49954 (N_49954,N_49536,N_49656);
nand U49955 (N_49955,N_49615,N_49592);
nor U49956 (N_49956,N_49506,N_49737);
nand U49957 (N_49957,N_49749,N_49544);
nand U49958 (N_49958,N_49640,N_49701);
nor U49959 (N_49959,N_49737,N_49748);
and U49960 (N_49960,N_49566,N_49742);
nor U49961 (N_49961,N_49658,N_49645);
nor U49962 (N_49962,N_49681,N_49718);
or U49963 (N_49963,N_49550,N_49692);
nor U49964 (N_49964,N_49677,N_49713);
nand U49965 (N_49965,N_49719,N_49660);
nor U49966 (N_49966,N_49612,N_49602);
xnor U49967 (N_49967,N_49603,N_49502);
nand U49968 (N_49968,N_49729,N_49727);
or U49969 (N_49969,N_49547,N_49705);
nor U49970 (N_49970,N_49542,N_49598);
nor U49971 (N_49971,N_49655,N_49662);
nand U49972 (N_49972,N_49534,N_49740);
and U49973 (N_49973,N_49518,N_49560);
nand U49974 (N_49974,N_49646,N_49544);
xor U49975 (N_49975,N_49606,N_49607);
xor U49976 (N_49976,N_49571,N_49510);
or U49977 (N_49977,N_49680,N_49667);
or U49978 (N_49978,N_49507,N_49580);
or U49979 (N_49979,N_49617,N_49588);
xnor U49980 (N_49980,N_49587,N_49689);
nor U49981 (N_49981,N_49536,N_49506);
xor U49982 (N_49982,N_49727,N_49665);
nor U49983 (N_49983,N_49711,N_49535);
xnor U49984 (N_49984,N_49715,N_49595);
nor U49985 (N_49985,N_49623,N_49597);
nand U49986 (N_49986,N_49685,N_49718);
xnor U49987 (N_49987,N_49539,N_49694);
nor U49988 (N_49988,N_49520,N_49624);
or U49989 (N_49989,N_49566,N_49678);
nor U49990 (N_49990,N_49545,N_49590);
nor U49991 (N_49991,N_49652,N_49697);
xnor U49992 (N_49992,N_49514,N_49540);
and U49993 (N_49993,N_49582,N_49573);
and U49994 (N_49994,N_49562,N_49602);
nand U49995 (N_49995,N_49601,N_49736);
or U49996 (N_49996,N_49675,N_49703);
nand U49997 (N_49997,N_49580,N_49550);
xor U49998 (N_49998,N_49560,N_49648);
and U49999 (N_49999,N_49595,N_49651);
nand UO_0 (O_0,N_49880,N_49918);
nand UO_1 (O_1,N_49859,N_49909);
xnor UO_2 (O_2,N_49782,N_49994);
xor UO_3 (O_3,N_49813,N_49759);
nor UO_4 (O_4,N_49970,N_49931);
or UO_5 (O_5,N_49905,N_49928);
and UO_6 (O_6,N_49802,N_49965);
nor UO_7 (O_7,N_49915,N_49989);
or UO_8 (O_8,N_49863,N_49819);
or UO_9 (O_9,N_49978,N_49973);
or UO_10 (O_10,N_49779,N_49943);
or UO_11 (O_11,N_49769,N_49860);
nor UO_12 (O_12,N_49812,N_49752);
nand UO_13 (O_13,N_49824,N_49758);
and UO_14 (O_14,N_49969,N_49876);
or UO_15 (O_15,N_49972,N_49976);
or UO_16 (O_16,N_49977,N_49901);
nor UO_17 (O_17,N_49956,N_49887);
xor UO_18 (O_18,N_49883,N_49757);
nand UO_19 (O_19,N_49835,N_49761);
and UO_20 (O_20,N_49766,N_49950);
xnor UO_21 (O_21,N_49933,N_49955);
nand UO_22 (O_22,N_49800,N_49875);
xnor UO_23 (O_23,N_49843,N_49796);
or UO_24 (O_24,N_49958,N_49991);
and UO_25 (O_25,N_49764,N_49889);
and UO_26 (O_26,N_49895,N_49959);
xnor UO_27 (O_27,N_49798,N_49784);
nor UO_28 (O_28,N_49961,N_49948);
xnor UO_29 (O_29,N_49916,N_49847);
nand UO_30 (O_30,N_49775,N_49795);
nor UO_31 (O_31,N_49919,N_49815);
or UO_32 (O_32,N_49832,N_49820);
xor UO_33 (O_33,N_49855,N_49962);
xnor UO_34 (O_34,N_49774,N_49947);
nor UO_35 (O_35,N_49845,N_49938);
and UO_36 (O_36,N_49981,N_49826);
nor UO_37 (O_37,N_49823,N_49792);
xor UO_38 (O_38,N_49987,N_49957);
xor UO_39 (O_39,N_49930,N_49881);
and UO_40 (O_40,N_49790,N_49854);
and UO_41 (O_41,N_49773,N_49874);
nor UO_42 (O_42,N_49982,N_49898);
nor UO_43 (O_43,N_49828,N_49986);
xnor UO_44 (O_44,N_49760,N_49866);
or UO_45 (O_45,N_49971,N_49885);
nand UO_46 (O_46,N_49914,N_49886);
xor UO_47 (O_47,N_49968,N_49979);
nand UO_48 (O_48,N_49829,N_49794);
xnor UO_49 (O_49,N_49809,N_49871);
nand UO_50 (O_50,N_49793,N_49780);
or UO_51 (O_51,N_49903,N_49750);
and UO_52 (O_52,N_49904,N_49830);
xor UO_53 (O_53,N_49906,N_49788);
nand UO_54 (O_54,N_49879,N_49893);
xnor UO_55 (O_55,N_49787,N_49926);
nand UO_56 (O_56,N_49936,N_49917);
and UO_57 (O_57,N_49814,N_49856);
nand UO_58 (O_58,N_49908,N_49964);
or UO_59 (O_59,N_49935,N_49932);
xnor UO_60 (O_60,N_49984,N_49807);
and UO_61 (O_61,N_49852,N_49990);
and UO_62 (O_62,N_49822,N_49877);
and UO_63 (O_63,N_49882,N_49891);
nor UO_64 (O_64,N_49940,N_49840);
and UO_65 (O_65,N_49870,N_49754);
nor UO_66 (O_66,N_49967,N_49833);
or UO_67 (O_67,N_49922,N_49992);
xor UO_68 (O_68,N_49857,N_49864);
or UO_69 (O_69,N_49949,N_49853);
xor UO_70 (O_70,N_49851,N_49786);
and UO_71 (O_71,N_49999,N_49762);
or UO_72 (O_72,N_49923,N_49839);
nand UO_73 (O_73,N_49996,N_49960);
nand UO_74 (O_74,N_49844,N_49921);
nor UO_75 (O_75,N_49806,N_49768);
or UO_76 (O_76,N_49929,N_49912);
and UO_77 (O_77,N_49825,N_49801);
or UO_78 (O_78,N_49805,N_49980);
nor UO_79 (O_79,N_49902,N_49897);
nand UO_80 (O_80,N_49778,N_49963);
or UO_81 (O_81,N_49842,N_49791);
nor UO_82 (O_82,N_49873,N_49827);
nand UO_83 (O_83,N_49983,N_49763);
xnor UO_84 (O_84,N_49900,N_49837);
and UO_85 (O_85,N_49896,N_49767);
and UO_86 (O_86,N_49910,N_49848);
and UO_87 (O_87,N_49783,N_49878);
and UO_88 (O_88,N_49966,N_49765);
or UO_89 (O_89,N_49988,N_49818);
nand UO_90 (O_90,N_49925,N_49838);
or UO_91 (O_91,N_49899,N_49944);
xnor UO_92 (O_92,N_49861,N_49789);
xnor UO_93 (O_93,N_49951,N_49846);
nand UO_94 (O_94,N_49755,N_49834);
nor UO_95 (O_95,N_49945,N_49942);
nand UO_96 (O_96,N_49811,N_49816);
xnor UO_97 (O_97,N_49756,N_49836);
and UO_98 (O_98,N_49975,N_49797);
nand UO_99 (O_99,N_49867,N_49862);
nor UO_100 (O_100,N_49850,N_49821);
and UO_101 (O_101,N_49817,N_49998);
or UO_102 (O_102,N_49884,N_49753);
nand UO_103 (O_103,N_49771,N_49946);
nor UO_104 (O_104,N_49985,N_49927);
xor UO_105 (O_105,N_49894,N_49872);
nor UO_106 (O_106,N_49924,N_49841);
or UO_107 (O_107,N_49913,N_49911);
or UO_108 (O_108,N_49907,N_49772);
nor UO_109 (O_109,N_49781,N_49803);
xnor UO_110 (O_110,N_49751,N_49993);
xor UO_111 (O_111,N_49808,N_49777);
or UO_112 (O_112,N_49785,N_49770);
xnor UO_113 (O_113,N_49939,N_49776);
nor UO_114 (O_114,N_49952,N_49888);
and UO_115 (O_115,N_49934,N_49920);
nand UO_116 (O_116,N_49810,N_49997);
nor UO_117 (O_117,N_49995,N_49869);
nand UO_118 (O_118,N_49849,N_49974);
nor UO_119 (O_119,N_49868,N_49937);
and UO_120 (O_120,N_49799,N_49804);
nand UO_121 (O_121,N_49890,N_49953);
xnor UO_122 (O_122,N_49831,N_49954);
or UO_123 (O_123,N_49858,N_49865);
nor UO_124 (O_124,N_49941,N_49892);
xnor UO_125 (O_125,N_49991,N_49764);
xnor UO_126 (O_126,N_49910,N_49764);
xnor UO_127 (O_127,N_49989,N_49784);
or UO_128 (O_128,N_49774,N_49864);
or UO_129 (O_129,N_49999,N_49950);
and UO_130 (O_130,N_49891,N_49904);
and UO_131 (O_131,N_49813,N_49810);
or UO_132 (O_132,N_49938,N_49873);
or UO_133 (O_133,N_49797,N_49790);
xnor UO_134 (O_134,N_49846,N_49958);
or UO_135 (O_135,N_49908,N_49832);
nand UO_136 (O_136,N_49961,N_49832);
nor UO_137 (O_137,N_49979,N_49997);
or UO_138 (O_138,N_49975,N_49992);
xnor UO_139 (O_139,N_49914,N_49974);
xnor UO_140 (O_140,N_49863,N_49860);
or UO_141 (O_141,N_49887,N_49883);
nand UO_142 (O_142,N_49990,N_49800);
xnor UO_143 (O_143,N_49920,N_49820);
or UO_144 (O_144,N_49819,N_49849);
nor UO_145 (O_145,N_49826,N_49849);
nor UO_146 (O_146,N_49972,N_49938);
xor UO_147 (O_147,N_49759,N_49882);
and UO_148 (O_148,N_49934,N_49921);
nor UO_149 (O_149,N_49790,N_49758);
and UO_150 (O_150,N_49978,N_49851);
nand UO_151 (O_151,N_49966,N_49965);
nand UO_152 (O_152,N_49836,N_49752);
xnor UO_153 (O_153,N_49982,N_49822);
and UO_154 (O_154,N_49931,N_49874);
nor UO_155 (O_155,N_49914,N_49931);
and UO_156 (O_156,N_49751,N_49832);
nand UO_157 (O_157,N_49953,N_49916);
or UO_158 (O_158,N_49777,N_49863);
xnor UO_159 (O_159,N_49993,N_49933);
xnor UO_160 (O_160,N_49998,N_49956);
and UO_161 (O_161,N_49930,N_49794);
and UO_162 (O_162,N_49884,N_49826);
nand UO_163 (O_163,N_49858,N_49831);
xnor UO_164 (O_164,N_49985,N_49771);
and UO_165 (O_165,N_49852,N_49833);
xor UO_166 (O_166,N_49831,N_49823);
and UO_167 (O_167,N_49926,N_49890);
and UO_168 (O_168,N_49880,N_49789);
nand UO_169 (O_169,N_49959,N_49906);
xnor UO_170 (O_170,N_49809,N_49927);
or UO_171 (O_171,N_49915,N_49896);
or UO_172 (O_172,N_49835,N_49825);
and UO_173 (O_173,N_49829,N_49972);
xnor UO_174 (O_174,N_49801,N_49986);
and UO_175 (O_175,N_49805,N_49859);
nor UO_176 (O_176,N_49768,N_49943);
nand UO_177 (O_177,N_49929,N_49878);
nand UO_178 (O_178,N_49930,N_49750);
or UO_179 (O_179,N_49913,N_49884);
and UO_180 (O_180,N_49800,N_49980);
xor UO_181 (O_181,N_49913,N_49907);
xnor UO_182 (O_182,N_49789,N_49846);
nand UO_183 (O_183,N_49921,N_49849);
nand UO_184 (O_184,N_49848,N_49953);
nand UO_185 (O_185,N_49973,N_49896);
xnor UO_186 (O_186,N_49755,N_49777);
and UO_187 (O_187,N_49809,N_49948);
or UO_188 (O_188,N_49842,N_49884);
nand UO_189 (O_189,N_49878,N_49825);
or UO_190 (O_190,N_49772,N_49877);
xnor UO_191 (O_191,N_49977,N_49969);
and UO_192 (O_192,N_49791,N_49890);
or UO_193 (O_193,N_49849,N_49798);
xnor UO_194 (O_194,N_49955,N_49987);
nand UO_195 (O_195,N_49929,N_49778);
nand UO_196 (O_196,N_49913,N_49807);
and UO_197 (O_197,N_49894,N_49784);
nor UO_198 (O_198,N_49802,N_49823);
and UO_199 (O_199,N_49893,N_49995);
nand UO_200 (O_200,N_49973,N_49970);
or UO_201 (O_201,N_49795,N_49954);
xor UO_202 (O_202,N_49966,N_49855);
xnor UO_203 (O_203,N_49957,N_49920);
xor UO_204 (O_204,N_49939,N_49985);
and UO_205 (O_205,N_49840,N_49994);
or UO_206 (O_206,N_49909,N_49877);
nand UO_207 (O_207,N_49937,N_49857);
and UO_208 (O_208,N_49952,N_49998);
and UO_209 (O_209,N_49937,N_49788);
nand UO_210 (O_210,N_49868,N_49813);
nor UO_211 (O_211,N_49836,N_49878);
nand UO_212 (O_212,N_49911,N_49934);
nand UO_213 (O_213,N_49993,N_49761);
nor UO_214 (O_214,N_49796,N_49804);
xnor UO_215 (O_215,N_49852,N_49933);
xnor UO_216 (O_216,N_49947,N_49805);
or UO_217 (O_217,N_49910,N_49933);
xnor UO_218 (O_218,N_49847,N_49876);
nor UO_219 (O_219,N_49939,N_49999);
xnor UO_220 (O_220,N_49757,N_49792);
and UO_221 (O_221,N_49885,N_49974);
xnor UO_222 (O_222,N_49765,N_49927);
xor UO_223 (O_223,N_49960,N_49803);
nor UO_224 (O_224,N_49845,N_49996);
or UO_225 (O_225,N_49989,N_49840);
xor UO_226 (O_226,N_49811,N_49858);
and UO_227 (O_227,N_49785,N_49869);
xor UO_228 (O_228,N_49854,N_49994);
or UO_229 (O_229,N_49912,N_49992);
nor UO_230 (O_230,N_49830,N_49916);
nor UO_231 (O_231,N_49904,N_49902);
nand UO_232 (O_232,N_49879,N_49864);
xnor UO_233 (O_233,N_49945,N_49983);
nor UO_234 (O_234,N_49833,N_49997);
nand UO_235 (O_235,N_49866,N_49951);
or UO_236 (O_236,N_49983,N_49874);
xor UO_237 (O_237,N_49769,N_49792);
or UO_238 (O_238,N_49827,N_49910);
xor UO_239 (O_239,N_49992,N_49957);
xor UO_240 (O_240,N_49830,N_49883);
nor UO_241 (O_241,N_49991,N_49931);
nand UO_242 (O_242,N_49812,N_49834);
and UO_243 (O_243,N_49895,N_49927);
or UO_244 (O_244,N_49801,N_49751);
or UO_245 (O_245,N_49930,N_49802);
nand UO_246 (O_246,N_49931,N_49870);
nand UO_247 (O_247,N_49980,N_49810);
and UO_248 (O_248,N_49823,N_49799);
xnor UO_249 (O_249,N_49883,N_49959);
nand UO_250 (O_250,N_49894,N_49837);
nor UO_251 (O_251,N_49979,N_49969);
nand UO_252 (O_252,N_49942,N_49954);
nor UO_253 (O_253,N_49943,N_49857);
xor UO_254 (O_254,N_49785,N_49939);
nor UO_255 (O_255,N_49862,N_49791);
nand UO_256 (O_256,N_49839,N_49799);
xor UO_257 (O_257,N_49902,N_49779);
and UO_258 (O_258,N_49867,N_49920);
and UO_259 (O_259,N_49799,N_49897);
or UO_260 (O_260,N_49969,N_49858);
xor UO_261 (O_261,N_49764,N_49795);
nor UO_262 (O_262,N_49963,N_49901);
or UO_263 (O_263,N_49791,N_49871);
nor UO_264 (O_264,N_49756,N_49861);
nor UO_265 (O_265,N_49854,N_49769);
xor UO_266 (O_266,N_49851,N_49884);
and UO_267 (O_267,N_49859,N_49892);
xor UO_268 (O_268,N_49933,N_49864);
xnor UO_269 (O_269,N_49889,N_49865);
and UO_270 (O_270,N_49968,N_49839);
nand UO_271 (O_271,N_49894,N_49994);
and UO_272 (O_272,N_49856,N_49799);
or UO_273 (O_273,N_49779,N_49944);
and UO_274 (O_274,N_49981,N_49887);
nand UO_275 (O_275,N_49939,N_49955);
xnor UO_276 (O_276,N_49947,N_49807);
or UO_277 (O_277,N_49958,N_49896);
or UO_278 (O_278,N_49991,N_49877);
nand UO_279 (O_279,N_49945,N_49858);
nand UO_280 (O_280,N_49986,N_49863);
and UO_281 (O_281,N_49873,N_49845);
nor UO_282 (O_282,N_49844,N_49773);
or UO_283 (O_283,N_49971,N_49814);
and UO_284 (O_284,N_49867,N_49856);
and UO_285 (O_285,N_49851,N_49805);
xor UO_286 (O_286,N_49867,N_49767);
nand UO_287 (O_287,N_49767,N_49769);
nor UO_288 (O_288,N_49787,N_49992);
nand UO_289 (O_289,N_49966,N_49920);
and UO_290 (O_290,N_49841,N_49871);
or UO_291 (O_291,N_49900,N_49954);
nor UO_292 (O_292,N_49977,N_49838);
xnor UO_293 (O_293,N_49840,N_49923);
xnor UO_294 (O_294,N_49909,N_49987);
and UO_295 (O_295,N_49863,N_49824);
nand UO_296 (O_296,N_49954,N_49918);
or UO_297 (O_297,N_49947,N_49929);
nand UO_298 (O_298,N_49795,N_49974);
and UO_299 (O_299,N_49937,N_49774);
nand UO_300 (O_300,N_49811,N_49797);
nor UO_301 (O_301,N_49935,N_49793);
or UO_302 (O_302,N_49945,N_49943);
xnor UO_303 (O_303,N_49953,N_49838);
xor UO_304 (O_304,N_49795,N_49767);
and UO_305 (O_305,N_49797,N_49865);
nand UO_306 (O_306,N_49805,N_49867);
nor UO_307 (O_307,N_49795,N_49970);
nor UO_308 (O_308,N_49992,N_49772);
nand UO_309 (O_309,N_49885,N_49782);
or UO_310 (O_310,N_49846,N_49904);
xor UO_311 (O_311,N_49805,N_49971);
or UO_312 (O_312,N_49994,N_49969);
and UO_313 (O_313,N_49804,N_49920);
xor UO_314 (O_314,N_49829,N_49948);
or UO_315 (O_315,N_49890,N_49754);
or UO_316 (O_316,N_49895,N_49770);
and UO_317 (O_317,N_49962,N_49860);
or UO_318 (O_318,N_49984,N_49972);
nand UO_319 (O_319,N_49883,N_49983);
and UO_320 (O_320,N_49795,N_49847);
nand UO_321 (O_321,N_49984,N_49946);
and UO_322 (O_322,N_49862,N_49896);
and UO_323 (O_323,N_49985,N_49844);
or UO_324 (O_324,N_49997,N_49945);
nor UO_325 (O_325,N_49861,N_49855);
nor UO_326 (O_326,N_49928,N_49971);
and UO_327 (O_327,N_49906,N_49793);
xor UO_328 (O_328,N_49846,N_49941);
nand UO_329 (O_329,N_49992,N_49935);
xnor UO_330 (O_330,N_49819,N_49782);
xnor UO_331 (O_331,N_49983,N_49941);
and UO_332 (O_332,N_49961,N_49810);
or UO_333 (O_333,N_49936,N_49948);
xnor UO_334 (O_334,N_49890,N_49848);
nand UO_335 (O_335,N_49943,N_49975);
nor UO_336 (O_336,N_49953,N_49760);
xor UO_337 (O_337,N_49989,N_49978);
or UO_338 (O_338,N_49806,N_49902);
and UO_339 (O_339,N_49992,N_49854);
and UO_340 (O_340,N_49776,N_49788);
nand UO_341 (O_341,N_49774,N_49945);
nand UO_342 (O_342,N_49808,N_49821);
nor UO_343 (O_343,N_49863,N_49996);
xnor UO_344 (O_344,N_49878,N_49828);
and UO_345 (O_345,N_49826,N_49998);
xnor UO_346 (O_346,N_49842,N_49898);
xnor UO_347 (O_347,N_49852,N_49997);
nand UO_348 (O_348,N_49900,N_49986);
and UO_349 (O_349,N_49829,N_49977);
and UO_350 (O_350,N_49807,N_49973);
or UO_351 (O_351,N_49752,N_49932);
and UO_352 (O_352,N_49929,N_49994);
or UO_353 (O_353,N_49935,N_49868);
nand UO_354 (O_354,N_49795,N_49978);
and UO_355 (O_355,N_49884,N_49771);
nand UO_356 (O_356,N_49837,N_49828);
xor UO_357 (O_357,N_49781,N_49857);
or UO_358 (O_358,N_49788,N_49940);
and UO_359 (O_359,N_49778,N_49820);
xnor UO_360 (O_360,N_49843,N_49926);
and UO_361 (O_361,N_49913,N_49843);
or UO_362 (O_362,N_49945,N_49898);
xnor UO_363 (O_363,N_49943,N_49988);
or UO_364 (O_364,N_49937,N_49806);
or UO_365 (O_365,N_49761,N_49876);
xor UO_366 (O_366,N_49801,N_49868);
or UO_367 (O_367,N_49789,N_49943);
xor UO_368 (O_368,N_49851,N_49814);
nor UO_369 (O_369,N_49758,N_49885);
xor UO_370 (O_370,N_49936,N_49873);
and UO_371 (O_371,N_49754,N_49912);
and UO_372 (O_372,N_49765,N_49930);
nor UO_373 (O_373,N_49789,N_49769);
nand UO_374 (O_374,N_49997,N_49859);
xor UO_375 (O_375,N_49804,N_49871);
and UO_376 (O_376,N_49969,N_49773);
or UO_377 (O_377,N_49794,N_49879);
or UO_378 (O_378,N_49751,N_49998);
xnor UO_379 (O_379,N_49997,N_49984);
nand UO_380 (O_380,N_49919,N_49803);
nand UO_381 (O_381,N_49931,N_49898);
xor UO_382 (O_382,N_49980,N_49939);
and UO_383 (O_383,N_49909,N_49908);
xor UO_384 (O_384,N_49905,N_49884);
and UO_385 (O_385,N_49892,N_49947);
or UO_386 (O_386,N_49836,N_49819);
xor UO_387 (O_387,N_49920,N_49861);
and UO_388 (O_388,N_49918,N_49911);
nor UO_389 (O_389,N_49821,N_49773);
and UO_390 (O_390,N_49948,N_49858);
nor UO_391 (O_391,N_49816,N_49819);
and UO_392 (O_392,N_49822,N_49870);
and UO_393 (O_393,N_49889,N_49863);
nand UO_394 (O_394,N_49852,N_49766);
nand UO_395 (O_395,N_49922,N_49928);
or UO_396 (O_396,N_49862,N_49829);
nand UO_397 (O_397,N_49935,N_49837);
and UO_398 (O_398,N_49806,N_49924);
and UO_399 (O_399,N_49946,N_49959);
xnor UO_400 (O_400,N_49928,N_49808);
xnor UO_401 (O_401,N_49983,N_49910);
or UO_402 (O_402,N_49814,N_49794);
or UO_403 (O_403,N_49784,N_49877);
and UO_404 (O_404,N_49799,N_49969);
nor UO_405 (O_405,N_49951,N_49879);
xnor UO_406 (O_406,N_49870,N_49929);
nand UO_407 (O_407,N_49990,N_49841);
nand UO_408 (O_408,N_49867,N_49895);
xor UO_409 (O_409,N_49779,N_49854);
and UO_410 (O_410,N_49980,N_49999);
and UO_411 (O_411,N_49952,N_49866);
and UO_412 (O_412,N_49891,N_49899);
xnor UO_413 (O_413,N_49803,N_49795);
or UO_414 (O_414,N_49916,N_49926);
nand UO_415 (O_415,N_49760,N_49905);
and UO_416 (O_416,N_49849,N_49889);
nor UO_417 (O_417,N_49977,N_49971);
nand UO_418 (O_418,N_49797,N_49819);
nand UO_419 (O_419,N_49871,N_49991);
nor UO_420 (O_420,N_49893,N_49783);
nand UO_421 (O_421,N_49813,N_49779);
nand UO_422 (O_422,N_49788,N_49771);
and UO_423 (O_423,N_49763,N_49856);
nand UO_424 (O_424,N_49770,N_49907);
nor UO_425 (O_425,N_49884,N_49925);
and UO_426 (O_426,N_49953,N_49841);
nand UO_427 (O_427,N_49850,N_49875);
nor UO_428 (O_428,N_49880,N_49968);
xor UO_429 (O_429,N_49988,N_49932);
and UO_430 (O_430,N_49853,N_49810);
and UO_431 (O_431,N_49831,N_49872);
and UO_432 (O_432,N_49974,N_49893);
nor UO_433 (O_433,N_49857,N_49833);
xor UO_434 (O_434,N_49814,N_49972);
xor UO_435 (O_435,N_49764,N_49868);
nand UO_436 (O_436,N_49943,N_49756);
xnor UO_437 (O_437,N_49872,N_49954);
nor UO_438 (O_438,N_49920,N_49803);
and UO_439 (O_439,N_49836,N_49921);
nand UO_440 (O_440,N_49870,N_49987);
nand UO_441 (O_441,N_49888,N_49918);
or UO_442 (O_442,N_49931,N_49889);
nor UO_443 (O_443,N_49864,N_49794);
nor UO_444 (O_444,N_49781,N_49987);
xor UO_445 (O_445,N_49997,N_49839);
and UO_446 (O_446,N_49849,N_49894);
nand UO_447 (O_447,N_49946,N_49795);
nor UO_448 (O_448,N_49976,N_49860);
xnor UO_449 (O_449,N_49975,N_49995);
nor UO_450 (O_450,N_49790,N_49782);
nand UO_451 (O_451,N_49966,N_49986);
nand UO_452 (O_452,N_49886,N_49789);
nor UO_453 (O_453,N_49891,N_49834);
nand UO_454 (O_454,N_49989,N_49865);
nand UO_455 (O_455,N_49799,N_49883);
and UO_456 (O_456,N_49804,N_49817);
nor UO_457 (O_457,N_49953,N_49755);
nand UO_458 (O_458,N_49797,N_49823);
and UO_459 (O_459,N_49930,N_49896);
and UO_460 (O_460,N_49960,N_49933);
nor UO_461 (O_461,N_49789,N_49888);
xor UO_462 (O_462,N_49759,N_49803);
nor UO_463 (O_463,N_49990,N_49862);
xnor UO_464 (O_464,N_49802,N_49813);
and UO_465 (O_465,N_49916,N_49970);
or UO_466 (O_466,N_49945,N_49768);
xor UO_467 (O_467,N_49878,N_49856);
and UO_468 (O_468,N_49896,N_49880);
and UO_469 (O_469,N_49836,N_49804);
and UO_470 (O_470,N_49874,N_49822);
and UO_471 (O_471,N_49968,N_49802);
nor UO_472 (O_472,N_49986,N_49833);
and UO_473 (O_473,N_49879,N_49924);
and UO_474 (O_474,N_49847,N_49903);
xor UO_475 (O_475,N_49827,N_49898);
xnor UO_476 (O_476,N_49930,N_49897);
xnor UO_477 (O_477,N_49967,N_49910);
nand UO_478 (O_478,N_49958,N_49859);
nor UO_479 (O_479,N_49858,N_49927);
nor UO_480 (O_480,N_49908,N_49773);
nand UO_481 (O_481,N_49883,N_49833);
and UO_482 (O_482,N_49790,N_49867);
nand UO_483 (O_483,N_49798,N_49896);
or UO_484 (O_484,N_49930,N_49757);
nand UO_485 (O_485,N_49852,N_49906);
nand UO_486 (O_486,N_49786,N_49808);
xor UO_487 (O_487,N_49937,N_49919);
and UO_488 (O_488,N_49844,N_49769);
nand UO_489 (O_489,N_49879,N_49756);
xor UO_490 (O_490,N_49868,N_49907);
nor UO_491 (O_491,N_49870,N_49927);
or UO_492 (O_492,N_49900,N_49795);
and UO_493 (O_493,N_49889,N_49915);
xor UO_494 (O_494,N_49971,N_49994);
and UO_495 (O_495,N_49755,N_49836);
nor UO_496 (O_496,N_49967,N_49804);
and UO_497 (O_497,N_49825,N_49861);
xor UO_498 (O_498,N_49870,N_49814);
or UO_499 (O_499,N_49782,N_49794);
or UO_500 (O_500,N_49950,N_49811);
nand UO_501 (O_501,N_49922,N_49883);
or UO_502 (O_502,N_49766,N_49922);
nand UO_503 (O_503,N_49953,N_49875);
or UO_504 (O_504,N_49884,N_49843);
and UO_505 (O_505,N_49762,N_49926);
nor UO_506 (O_506,N_49906,N_49875);
or UO_507 (O_507,N_49802,N_49985);
xnor UO_508 (O_508,N_49963,N_49864);
xnor UO_509 (O_509,N_49830,N_49906);
xor UO_510 (O_510,N_49879,N_49801);
and UO_511 (O_511,N_49808,N_49937);
nor UO_512 (O_512,N_49921,N_49915);
xor UO_513 (O_513,N_49997,N_49901);
or UO_514 (O_514,N_49787,N_49994);
and UO_515 (O_515,N_49873,N_49870);
xnor UO_516 (O_516,N_49891,N_49803);
and UO_517 (O_517,N_49890,N_49892);
nand UO_518 (O_518,N_49872,N_49930);
nand UO_519 (O_519,N_49808,N_49920);
nand UO_520 (O_520,N_49954,N_49761);
nand UO_521 (O_521,N_49987,N_49915);
and UO_522 (O_522,N_49781,N_49832);
xor UO_523 (O_523,N_49973,N_49812);
and UO_524 (O_524,N_49782,N_49935);
and UO_525 (O_525,N_49930,N_49936);
xnor UO_526 (O_526,N_49873,N_49969);
and UO_527 (O_527,N_49857,N_49908);
xnor UO_528 (O_528,N_49876,N_49935);
or UO_529 (O_529,N_49894,N_49803);
nor UO_530 (O_530,N_49898,N_49856);
nor UO_531 (O_531,N_49880,N_49863);
or UO_532 (O_532,N_49932,N_49807);
xnor UO_533 (O_533,N_49939,N_49904);
or UO_534 (O_534,N_49846,N_49960);
and UO_535 (O_535,N_49798,N_49933);
xnor UO_536 (O_536,N_49834,N_49777);
xor UO_537 (O_537,N_49933,N_49816);
xor UO_538 (O_538,N_49822,N_49798);
or UO_539 (O_539,N_49985,N_49903);
nor UO_540 (O_540,N_49771,N_49785);
and UO_541 (O_541,N_49890,N_49792);
nor UO_542 (O_542,N_49812,N_49782);
nor UO_543 (O_543,N_49942,N_49824);
xor UO_544 (O_544,N_49815,N_49894);
and UO_545 (O_545,N_49804,N_49874);
xnor UO_546 (O_546,N_49783,N_49929);
and UO_547 (O_547,N_49922,N_49969);
or UO_548 (O_548,N_49988,N_49805);
and UO_549 (O_549,N_49837,N_49829);
and UO_550 (O_550,N_49872,N_49774);
and UO_551 (O_551,N_49806,N_49903);
and UO_552 (O_552,N_49913,N_49835);
and UO_553 (O_553,N_49816,N_49985);
nand UO_554 (O_554,N_49770,N_49886);
or UO_555 (O_555,N_49885,N_49864);
or UO_556 (O_556,N_49889,N_49846);
nand UO_557 (O_557,N_49896,N_49902);
nor UO_558 (O_558,N_49886,N_49966);
nand UO_559 (O_559,N_49980,N_49791);
or UO_560 (O_560,N_49837,N_49943);
or UO_561 (O_561,N_49846,N_49891);
xnor UO_562 (O_562,N_49753,N_49857);
or UO_563 (O_563,N_49939,N_49778);
nand UO_564 (O_564,N_49917,N_49904);
nor UO_565 (O_565,N_49921,N_49777);
xor UO_566 (O_566,N_49858,N_49915);
xor UO_567 (O_567,N_49776,N_49908);
xor UO_568 (O_568,N_49782,N_49881);
nand UO_569 (O_569,N_49878,N_49802);
or UO_570 (O_570,N_49795,N_49811);
nor UO_571 (O_571,N_49801,N_49949);
nand UO_572 (O_572,N_49877,N_49912);
xnor UO_573 (O_573,N_49975,N_49778);
and UO_574 (O_574,N_49882,N_49962);
nor UO_575 (O_575,N_49989,N_49910);
nor UO_576 (O_576,N_49983,N_49778);
nand UO_577 (O_577,N_49946,N_49912);
nor UO_578 (O_578,N_49818,N_49954);
nor UO_579 (O_579,N_49980,N_49912);
xnor UO_580 (O_580,N_49763,N_49839);
nor UO_581 (O_581,N_49986,N_49866);
and UO_582 (O_582,N_49790,N_49789);
nor UO_583 (O_583,N_49994,N_49831);
or UO_584 (O_584,N_49992,N_49885);
and UO_585 (O_585,N_49821,N_49916);
nand UO_586 (O_586,N_49797,N_49812);
or UO_587 (O_587,N_49894,N_49887);
nand UO_588 (O_588,N_49765,N_49969);
or UO_589 (O_589,N_49854,N_49981);
or UO_590 (O_590,N_49805,N_49787);
nor UO_591 (O_591,N_49943,N_49785);
nand UO_592 (O_592,N_49977,N_49849);
nor UO_593 (O_593,N_49929,N_49988);
nor UO_594 (O_594,N_49792,N_49848);
or UO_595 (O_595,N_49781,N_49874);
and UO_596 (O_596,N_49942,N_49868);
nor UO_597 (O_597,N_49769,N_49978);
or UO_598 (O_598,N_49781,N_49977);
nor UO_599 (O_599,N_49824,N_49823);
nand UO_600 (O_600,N_49919,N_49904);
xor UO_601 (O_601,N_49835,N_49850);
xnor UO_602 (O_602,N_49952,N_49968);
and UO_603 (O_603,N_49940,N_49996);
or UO_604 (O_604,N_49824,N_49869);
or UO_605 (O_605,N_49886,N_49762);
xnor UO_606 (O_606,N_49908,N_49969);
xor UO_607 (O_607,N_49767,N_49757);
nand UO_608 (O_608,N_49852,N_49776);
or UO_609 (O_609,N_49926,N_49984);
xnor UO_610 (O_610,N_49822,N_49864);
xnor UO_611 (O_611,N_49773,N_49766);
nor UO_612 (O_612,N_49979,N_49988);
xor UO_613 (O_613,N_49810,N_49917);
xor UO_614 (O_614,N_49766,N_49911);
nand UO_615 (O_615,N_49957,N_49826);
and UO_616 (O_616,N_49870,N_49905);
xnor UO_617 (O_617,N_49872,N_49803);
xnor UO_618 (O_618,N_49978,N_49792);
nor UO_619 (O_619,N_49995,N_49883);
nor UO_620 (O_620,N_49773,N_49840);
nand UO_621 (O_621,N_49892,N_49828);
xor UO_622 (O_622,N_49804,N_49847);
nand UO_623 (O_623,N_49808,N_49985);
xor UO_624 (O_624,N_49981,N_49821);
nor UO_625 (O_625,N_49929,N_49882);
and UO_626 (O_626,N_49771,N_49868);
nor UO_627 (O_627,N_49894,N_49755);
xnor UO_628 (O_628,N_49751,N_49903);
and UO_629 (O_629,N_49760,N_49902);
xnor UO_630 (O_630,N_49755,N_49855);
nand UO_631 (O_631,N_49898,N_49998);
xor UO_632 (O_632,N_49809,N_49864);
xnor UO_633 (O_633,N_49847,N_49819);
nand UO_634 (O_634,N_49942,N_49993);
and UO_635 (O_635,N_49939,N_49927);
nand UO_636 (O_636,N_49926,N_49810);
nand UO_637 (O_637,N_49852,N_49922);
nand UO_638 (O_638,N_49937,N_49942);
nand UO_639 (O_639,N_49814,N_49788);
or UO_640 (O_640,N_49850,N_49954);
nand UO_641 (O_641,N_49793,N_49862);
or UO_642 (O_642,N_49805,N_49820);
or UO_643 (O_643,N_49850,N_49786);
nor UO_644 (O_644,N_49906,N_49805);
or UO_645 (O_645,N_49993,N_49840);
and UO_646 (O_646,N_49830,N_49968);
nor UO_647 (O_647,N_49927,N_49812);
nand UO_648 (O_648,N_49991,N_49825);
and UO_649 (O_649,N_49951,N_49780);
or UO_650 (O_650,N_49990,N_49914);
nand UO_651 (O_651,N_49913,N_49855);
nand UO_652 (O_652,N_49833,N_49940);
or UO_653 (O_653,N_49856,N_49768);
or UO_654 (O_654,N_49901,N_49882);
or UO_655 (O_655,N_49957,N_49752);
or UO_656 (O_656,N_49801,N_49790);
and UO_657 (O_657,N_49774,N_49962);
nand UO_658 (O_658,N_49925,N_49806);
nor UO_659 (O_659,N_49872,N_49864);
nor UO_660 (O_660,N_49785,N_49857);
or UO_661 (O_661,N_49780,N_49998);
nand UO_662 (O_662,N_49827,N_49901);
xor UO_663 (O_663,N_49940,N_49974);
nand UO_664 (O_664,N_49881,N_49750);
and UO_665 (O_665,N_49789,N_49976);
and UO_666 (O_666,N_49883,N_49819);
nand UO_667 (O_667,N_49880,N_49975);
nor UO_668 (O_668,N_49833,N_49920);
xnor UO_669 (O_669,N_49866,N_49942);
xnor UO_670 (O_670,N_49965,N_49983);
nand UO_671 (O_671,N_49893,N_49887);
nand UO_672 (O_672,N_49907,N_49924);
or UO_673 (O_673,N_49880,N_49961);
xor UO_674 (O_674,N_49933,N_49945);
or UO_675 (O_675,N_49882,N_49916);
and UO_676 (O_676,N_49971,N_49936);
xnor UO_677 (O_677,N_49750,N_49915);
xor UO_678 (O_678,N_49764,N_49962);
nor UO_679 (O_679,N_49931,N_49778);
and UO_680 (O_680,N_49844,N_49899);
and UO_681 (O_681,N_49915,N_49845);
xnor UO_682 (O_682,N_49914,N_49894);
nor UO_683 (O_683,N_49998,N_49999);
nand UO_684 (O_684,N_49755,N_49914);
xnor UO_685 (O_685,N_49758,N_49901);
nand UO_686 (O_686,N_49773,N_49783);
and UO_687 (O_687,N_49866,N_49833);
nor UO_688 (O_688,N_49814,N_49764);
nand UO_689 (O_689,N_49991,N_49903);
xnor UO_690 (O_690,N_49986,N_49965);
and UO_691 (O_691,N_49843,N_49970);
nor UO_692 (O_692,N_49873,N_49836);
xor UO_693 (O_693,N_49809,N_49970);
or UO_694 (O_694,N_49866,N_49825);
xnor UO_695 (O_695,N_49926,N_49838);
nand UO_696 (O_696,N_49893,N_49792);
and UO_697 (O_697,N_49999,N_49957);
nor UO_698 (O_698,N_49845,N_49923);
and UO_699 (O_699,N_49897,N_49776);
xor UO_700 (O_700,N_49823,N_49873);
nand UO_701 (O_701,N_49913,N_49803);
nand UO_702 (O_702,N_49935,N_49899);
and UO_703 (O_703,N_49930,N_49809);
and UO_704 (O_704,N_49926,N_49967);
xor UO_705 (O_705,N_49900,N_49752);
or UO_706 (O_706,N_49754,N_49862);
and UO_707 (O_707,N_49796,N_49943);
nor UO_708 (O_708,N_49944,N_49784);
xor UO_709 (O_709,N_49751,N_49780);
or UO_710 (O_710,N_49908,N_49824);
and UO_711 (O_711,N_49946,N_49810);
nor UO_712 (O_712,N_49844,N_49772);
nand UO_713 (O_713,N_49929,N_49838);
nor UO_714 (O_714,N_49797,N_49978);
and UO_715 (O_715,N_49928,N_49890);
xor UO_716 (O_716,N_49945,N_49824);
or UO_717 (O_717,N_49764,N_49832);
or UO_718 (O_718,N_49807,N_49783);
or UO_719 (O_719,N_49949,N_49758);
xnor UO_720 (O_720,N_49908,N_49780);
nor UO_721 (O_721,N_49902,N_49974);
xor UO_722 (O_722,N_49886,N_49890);
and UO_723 (O_723,N_49926,N_49937);
and UO_724 (O_724,N_49854,N_49788);
nand UO_725 (O_725,N_49874,N_49795);
nor UO_726 (O_726,N_49934,N_49867);
xor UO_727 (O_727,N_49969,N_49865);
xnor UO_728 (O_728,N_49967,N_49830);
or UO_729 (O_729,N_49970,N_49910);
or UO_730 (O_730,N_49969,N_49826);
nor UO_731 (O_731,N_49846,N_49860);
nor UO_732 (O_732,N_49982,N_49969);
and UO_733 (O_733,N_49771,N_49885);
or UO_734 (O_734,N_49887,N_49947);
nor UO_735 (O_735,N_49818,N_49761);
or UO_736 (O_736,N_49867,N_49993);
xnor UO_737 (O_737,N_49846,N_49881);
and UO_738 (O_738,N_49790,N_49778);
nand UO_739 (O_739,N_49970,N_49785);
and UO_740 (O_740,N_49841,N_49888);
or UO_741 (O_741,N_49933,N_49857);
xor UO_742 (O_742,N_49982,N_49963);
nor UO_743 (O_743,N_49922,N_49866);
nand UO_744 (O_744,N_49935,N_49796);
and UO_745 (O_745,N_49987,N_49799);
nor UO_746 (O_746,N_49755,N_49890);
or UO_747 (O_747,N_49756,N_49758);
and UO_748 (O_748,N_49763,N_49800);
and UO_749 (O_749,N_49935,N_49953);
and UO_750 (O_750,N_49870,N_49874);
nand UO_751 (O_751,N_49984,N_49995);
nand UO_752 (O_752,N_49995,N_49993);
nor UO_753 (O_753,N_49841,N_49761);
xor UO_754 (O_754,N_49989,N_49977);
nand UO_755 (O_755,N_49830,N_49992);
nor UO_756 (O_756,N_49826,N_49778);
xor UO_757 (O_757,N_49828,N_49933);
xor UO_758 (O_758,N_49768,N_49760);
and UO_759 (O_759,N_49897,N_49994);
and UO_760 (O_760,N_49964,N_49814);
nand UO_761 (O_761,N_49949,N_49802);
xor UO_762 (O_762,N_49867,N_49900);
nand UO_763 (O_763,N_49755,N_49875);
or UO_764 (O_764,N_49766,N_49783);
and UO_765 (O_765,N_49997,N_49844);
or UO_766 (O_766,N_49750,N_49859);
and UO_767 (O_767,N_49927,N_49978);
nor UO_768 (O_768,N_49804,N_49930);
nand UO_769 (O_769,N_49923,N_49834);
xnor UO_770 (O_770,N_49836,N_49856);
nand UO_771 (O_771,N_49963,N_49764);
nand UO_772 (O_772,N_49994,N_49778);
or UO_773 (O_773,N_49825,N_49762);
xor UO_774 (O_774,N_49931,N_49784);
nor UO_775 (O_775,N_49882,N_49875);
xnor UO_776 (O_776,N_49812,N_49810);
nor UO_777 (O_777,N_49850,N_49981);
and UO_778 (O_778,N_49941,N_49877);
nor UO_779 (O_779,N_49849,N_49908);
or UO_780 (O_780,N_49906,N_49967);
and UO_781 (O_781,N_49778,N_49885);
nand UO_782 (O_782,N_49911,N_49942);
xor UO_783 (O_783,N_49808,N_49785);
and UO_784 (O_784,N_49836,N_49950);
or UO_785 (O_785,N_49921,N_49891);
nand UO_786 (O_786,N_49992,N_49934);
and UO_787 (O_787,N_49823,N_49858);
nand UO_788 (O_788,N_49839,N_49838);
and UO_789 (O_789,N_49924,N_49829);
nand UO_790 (O_790,N_49901,N_49786);
and UO_791 (O_791,N_49884,N_49881);
or UO_792 (O_792,N_49819,N_49891);
or UO_793 (O_793,N_49944,N_49900);
and UO_794 (O_794,N_49852,N_49750);
and UO_795 (O_795,N_49877,N_49870);
nand UO_796 (O_796,N_49780,N_49964);
and UO_797 (O_797,N_49853,N_49920);
nand UO_798 (O_798,N_49923,N_49978);
or UO_799 (O_799,N_49957,N_49809);
and UO_800 (O_800,N_49951,N_49862);
nor UO_801 (O_801,N_49977,N_49885);
nand UO_802 (O_802,N_49835,N_49896);
and UO_803 (O_803,N_49956,N_49779);
or UO_804 (O_804,N_49988,N_49830);
nand UO_805 (O_805,N_49940,N_49928);
xor UO_806 (O_806,N_49909,N_49770);
xor UO_807 (O_807,N_49851,N_49953);
nand UO_808 (O_808,N_49764,N_49752);
or UO_809 (O_809,N_49772,N_49934);
nand UO_810 (O_810,N_49935,N_49895);
and UO_811 (O_811,N_49766,N_49951);
nand UO_812 (O_812,N_49981,N_49845);
nand UO_813 (O_813,N_49874,N_49793);
or UO_814 (O_814,N_49889,N_49811);
xnor UO_815 (O_815,N_49930,N_49766);
and UO_816 (O_816,N_49781,N_49810);
nand UO_817 (O_817,N_49818,N_49876);
and UO_818 (O_818,N_49798,N_49869);
xor UO_819 (O_819,N_49784,N_49778);
and UO_820 (O_820,N_49883,N_49823);
xor UO_821 (O_821,N_49829,N_49783);
nand UO_822 (O_822,N_49895,N_49864);
and UO_823 (O_823,N_49828,N_49895);
xnor UO_824 (O_824,N_49810,N_49847);
nand UO_825 (O_825,N_49845,N_49896);
xor UO_826 (O_826,N_49947,N_49904);
and UO_827 (O_827,N_49935,N_49750);
nand UO_828 (O_828,N_49833,N_49964);
xor UO_829 (O_829,N_49997,N_49868);
nand UO_830 (O_830,N_49753,N_49788);
or UO_831 (O_831,N_49812,N_49799);
nor UO_832 (O_832,N_49781,N_49973);
and UO_833 (O_833,N_49974,N_49995);
and UO_834 (O_834,N_49964,N_49855);
and UO_835 (O_835,N_49802,N_49755);
or UO_836 (O_836,N_49789,N_49752);
and UO_837 (O_837,N_49831,N_49875);
nor UO_838 (O_838,N_49844,N_49981);
or UO_839 (O_839,N_49948,N_49926);
nand UO_840 (O_840,N_49832,N_49824);
xor UO_841 (O_841,N_49881,N_49826);
nor UO_842 (O_842,N_49905,N_49843);
or UO_843 (O_843,N_49781,N_49865);
and UO_844 (O_844,N_49863,N_49813);
xnor UO_845 (O_845,N_49802,N_49854);
nand UO_846 (O_846,N_49792,N_49803);
nor UO_847 (O_847,N_49949,N_49904);
or UO_848 (O_848,N_49964,N_49784);
xnor UO_849 (O_849,N_49795,N_49759);
nand UO_850 (O_850,N_49930,N_49958);
and UO_851 (O_851,N_49894,N_49965);
and UO_852 (O_852,N_49987,N_49910);
nand UO_853 (O_853,N_49971,N_49856);
xnor UO_854 (O_854,N_49963,N_49924);
nand UO_855 (O_855,N_49937,N_49972);
nand UO_856 (O_856,N_49815,N_49836);
and UO_857 (O_857,N_49885,N_49858);
and UO_858 (O_858,N_49848,N_49957);
nor UO_859 (O_859,N_49777,N_49790);
and UO_860 (O_860,N_49970,N_49805);
nor UO_861 (O_861,N_49788,N_49993);
and UO_862 (O_862,N_49956,N_49949);
or UO_863 (O_863,N_49927,N_49991);
nand UO_864 (O_864,N_49842,N_49853);
nor UO_865 (O_865,N_49882,N_49831);
and UO_866 (O_866,N_49850,N_49931);
or UO_867 (O_867,N_49937,N_49904);
and UO_868 (O_868,N_49842,N_49875);
and UO_869 (O_869,N_49876,N_49797);
nand UO_870 (O_870,N_49829,N_49856);
and UO_871 (O_871,N_49893,N_49924);
nor UO_872 (O_872,N_49890,N_49833);
xnor UO_873 (O_873,N_49885,N_49793);
or UO_874 (O_874,N_49797,N_49894);
and UO_875 (O_875,N_49846,N_49864);
nand UO_876 (O_876,N_49991,N_49834);
or UO_877 (O_877,N_49966,N_49758);
nor UO_878 (O_878,N_49892,N_49909);
nand UO_879 (O_879,N_49758,N_49964);
xnor UO_880 (O_880,N_49851,N_49837);
xor UO_881 (O_881,N_49827,N_49837);
nand UO_882 (O_882,N_49948,N_49974);
nand UO_883 (O_883,N_49884,N_49980);
nor UO_884 (O_884,N_49973,N_49810);
nand UO_885 (O_885,N_49899,N_49975);
nand UO_886 (O_886,N_49848,N_49811);
xnor UO_887 (O_887,N_49775,N_49796);
nand UO_888 (O_888,N_49850,N_49788);
nor UO_889 (O_889,N_49898,N_49826);
nand UO_890 (O_890,N_49997,N_49798);
nand UO_891 (O_891,N_49934,N_49990);
nand UO_892 (O_892,N_49934,N_49918);
xor UO_893 (O_893,N_49866,N_49813);
xnor UO_894 (O_894,N_49895,N_49998);
and UO_895 (O_895,N_49911,N_49763);
xor UO_896 (O_896,N_49990,N_49913);
and UO_897 (O_897,N_49995,N_49839);
xnor UO_898 (O_898,N_49891,N_49858);
xnor UO_899 (O_899,N_49826,N_49940);
or UO_900 (O_900,N_49886,N_49763);
xnor UO_901 (O_901,N_49918,N_49776);
xnor UO_902 (O_902,N_49924,N_49864);
nand UO_903 (O_903,N_49948,N_49937);
xnor UO_904 (O_904,N_49891,N_49771);
and UO_905 (O_905,N_49987,N_49854);
and UO_906 (O_906,N_49978,N_49998);
and UO_907 (O_907,N_49911,N_49815);
nor UO_908 (O_908,N_49897,N_49934);
or UO_909 (O_909,N_49898,N_49934);
and UO_910 (O_910,N_49773,N_49880);
nand UO_911 (O_911,N_49833,N_49830);
nor UO_912 (O_912,N_49955,N_49988);
nor UO_913 (O_913,N_49906,N_49820);
nand UO_914 (O_914,N_49919,N_49756);
nand UO_915 (O_915,N_49935,N_49972);
nor UO_916 (O_916,N_49931,N_49955);
or UO_917 (O_917,N_49955,N_49978);
and UO_918 (O_918,N_49889,N_49807);
or UO_919 (O_919,N_49820,N_49817);
and UO_920 (O_920,N_49979,N_49880);
and UO_921 (O_921,N_49957,N_49755);
or UO_922 (O_922,N_49877,N_49933);
xnor UO_923 (O_923,N_49928,N_49858);
xor UO_924 (O_924,N_49792,N_49901);
nor UO_925 (O_925,N_49758,N_49861);
nand UO_926 (O_926,N_49806,N_49949);
or UO_927 (O_927,N_49973,N_49928);
xor UO_928 (O_928,N_49852,N_49850);
nand UO_929 (O_929,N_49999,N_49973);
nor UO_930 (O_930,N_49882,N_49826);
nor UO_931 (O_931,N_49935,N_49989);
xor UO_932 (O_932,N_49919,N_49892);
or UO_933 (O_933,N_49756,N_49901);
nor UO_934 (O_934,N_49989,N_49952);
and UO_935 (O_935,N_49767,N_49840);
and UO_936 (O_936,N_49961,N_49834);
nor UO_937 (O_937,N_49775,N_49753);
nor UO_938 (O_938,N_49830,N_49847);
nor UO_939 (O_939,N_49973,N_49971);
or UO_940 (O_940,N_49897,N_49958);
or UO_941 (O_941,N_49851,N_49826);
and UO_942 (O_942,N_49959,N_49829);
nand UO_943 (O_943,N_49887,N_49881);
nand UO_944 (O_944,N_49844,N_49784);
and UO_945 (O_945,N_49888,N_49805);
and UO_946 (O_946,N_49959,N_49935);
xor UO_947 (O_947,N_49888,N_49990);
nand UO_948 (O_948,N_49872,N_49916);
xnor UO_949 (O_949,N_49840,N_49920);
xor UO_950 (O_950,N_49752,N_49878);
nor UO_951 (O_951,N_49853,N_49952);
and UO_952 (O_952,N_49921,N_49809);
nand UO_953 (O_953,N_49938,N_49812);
xor UO_954 (O_954,N_49849,N_49935);
nor UO_955 (O_955,N_49794,N_49886);
nor UO_956 (O_956,N_49814,N_49887);
and UO_957 (O_957,N_49907,N_49851);
xnor UO_958 (O_958,N_49973,N_49895);
nor UO_959 (O_959,N_49800,N_49993);
nor UO_960 (O_960,N_49973,N_49777);
xnor UO_961 (O_961,N_49814,N_49756);
or UO_962 (O_962,N_49986,N_49755);
xor UO_963 (O_963,N_49835,N_49866);
and UO_964 (O_964,N_49943,N_49907);
and UO_965 (O_965,N_49932,N_49978);
xnor UO_966 (O_966,N_49910,N_49814);
and UO_967 (O_967,N_49866,N_49759);
nor UO_968 (O_968,N_49797,N_49751);
and UO_969 (O_969,N_49890,N_49988);
or UO_970 (O_970,N_49860,N_49814);
and UO_971 (O_971,N_49929,N_49794);
xnor UO_972 (O_972,N_49915,N_49935);
or UO_973 (O_973,N_49969,N_49943);
or UO_974 (O_974,N_49892,N_49767);
nor UO_975 (O_975,N_49764,N_49906);
nand UO_976 (O_976,N_49788,N_49848);
nor UO_977 (O_977,N_49863,N_49757);
or UO_978 (O_978,N_49938,N_49780);
or UO_979 (O_979,N_49967,N_49784);
nand UO_980 (O_980,N_49905,N_49798);
and UO_981 (O_981,N_49862,N_49920);
xor UO_982 (O_982,N_49993,N_49943);
nor UO_983 (O_983,N_49819,N_49801);
or UO_984 (O_984,N_49858,N_49779);
nor UO_985 (O_985,N_49817,N_49994);
and UO_986 (O_986,N_49876,N_49927);
and UO_987 (O_987,N_49875,N_49833);
xor UO_988 (O_988,N_49773,N_49932);
and UO_989 (O_989,N_49940,N_49901);
and UO_990 (O_990,N_49936,N_49755);
nand UO_991 (O_991,N_49898,N_49833);
and UO_992 (O_992,N_49856,N_49961);
and UO_993 (O_993,N_49850,N_49818);
nand UO_994 (O_994,N_49786,N_49831);
nor UO_995 (O_995,N_49825,N_49791);
or UO_996 (O_996,N_49823,N_49947);
xnor UO_997 (O_997,N_49976,N_49991);
nor UO_998 (O_998,N_49808,N_49912);
or UO_999 (O_999,N_49881,N_49879);
nor UO_1000 (O_1000,N_49887,N_49964);
xnor UO_1001 (O_1001,N_49988,N_49843);
or UO_1002 (O_1002,N_49966,N_49960);
nand UO_1003 (O_1003,N_49980,N_49756);
and UO_1004 (O_1004,N_49816,N_49909);
or UO_1005 (O_1005,N_49986,N_49972);
or UO_1006 (O_1006,N_49761,N_49932);
or UO_1007 (O_1007,N_49998,N_49833);
xnor UO_1008 (O_1008,N_49815,N_49807);
nor UO_1009 (O_1009,N_49793,N_49815);
or UO_1010 (O_1010,N_49761,N_49960);
xnor UO_1011 (O_1011,N_49976,N_49894);
and UO_1012 (O_1012,N_49983,N_49930);
or UO_1013 (O_1013,N_49856,N_49921);
xor UO_1014 (O_1014,N_49774,N_49917);
nand UO_1015 (O_1015,N_49840,N_49841);
xnor UO_1016 (O_1016,N_49870,N_49894);
and UO_1017 (O_1017,N_49808,N_49995);
nand UO_1018 (O_1018,N_49793,N_49844);
or UO_1019 (O_1019,N_49963,N_49921);
nor UO_1020 (O_1020,N_49955,N_49779);
or UO_1021 (O_1021,N_49799,N_49869);
nand UO_1022 (O_1022,N_49764,N_49884);
nor UO_1023 (O_1023,N_49846,N_49892);
and UO_1024 (O_1024,N_49957,N_49949);
and UO_1025 (O_1025,N_49754,N_49851);
nand UO_1026 (O_1026,N_49792,N_49873);
or UO_1027 (O_1027,N_49811,N_49879);
xor UO_1028 (O_1028,N_49883,N_49807);
nand UO_1029 (O_1029,N_49757,N_49916);
or UO_1030 (O_1030,N_49972,N_49789);
nand UO_1031 (O_1031,N_49831,N_49979);
and UO_1032 (O_1032,N_49797,N_49752);
xnor UO_1033 (O_1033,N_49830,N_49836);
and UO_1034 (O_1034,N_49923,N_49903);
and UO_1035 (O_1035,N_49970,N_49971);
nand UO_1036 (O_1036,N_49966,N_49818);
xnor UO_1037 (O_1037,N_49804,N_49938);
and UO_1038 (O_1038,N_49972,N_49904);
xnor UO_1039 (O_1039,N_49856,N_49750);
and UO_1040 (O_1040,N_49810,N_49835);
nor UO_1041 (O_1041,N_49956,N_49917);
xnor UO_1042 (O_1042,N_49875,N_49955);
nand UO_1043 (O_1043,N_49881,N_49837);
nand UO_1044 (O_1044,N_49856,N_49769);
or UO_1045 (O_1045,N_49927,N_49963);
or UO_1046 (O_1046,N_49932,N_49859);
xor UO_1047 (O_1047,N_49815,N_49960);
xor UO_1048 (O_1048,N_49941,N_49995);
nand UO_1049 (O_1049,N_49979,N_49839);
nand UO_1050 (O_1050,N_49816,N_49948);
nand UO_1051 (O_1051,N_49889,N_49883);
and UO_1052 (O_1052,N_49859,N_49849);
nor UO_1053 (O_1053,N_49877,N_49832);
nor UO_1054 (O_1054,N_49981,N_49987);
or UO_1055 (O_1055,N_49972,N_49926);
nor UO_1056 (O_1056,N_49798,N_49783);
nor UO_1057 (O_1057,N_49882,N_49811);
xnor UO_1058 (O_1058,N_49907,N_49765);
nand UO_1059 (O_1059,N_49874,N_49758);
nand UO_1060 (O_1060,N_49840,N_49862);
nand UO_1061 (O_1061,N_49794,N_49948);
nand UO_1062 (O_1062,N_49792,N_49754);
nand UO_1063 (O_1063,N_49991,N_49940);
nand UO_1064 (O_1064,N_49813,N_49979);
or UO_1065 (O_1065,N_49812,N_49774);
or UO_1066 (O_1066,N_49773,N_49814);
or UO_1067 (O_1067,N_49882,N_49760);
xnor UO_1068 (O_1068,N_49801,N_49836);
and UO_1069 (O_1069,N_49877,N_49865);
nor UO_1070 (O_1070,N_49911,N_49893);
xor UO_1071 (O_1071,N_49767,N_49963);
nand UO_1072 (O_1072,N_49999,N_49821);
xnor UO_1073 (O_1073,N_49938,N_49844);
and UO_1074 (O_1074,N_49884,N_49908);
xor UO_1075 (O_1075,N_49786,N_49798);
nor UO_1076 (O_1076,N_49998,N_49822);
and UO_1077 (O_1077,N_49774,N_49829);
nand UO_1078 (O_1078,N_49780,N_49932);
xor UO_1079 (O_1079,N_49913,N_49962);
nand UO_1080 (O_1080,N_49862,N_49869);
nand UO_1081 (O_1081,N_49848,N_49869);
or UO_1082 (O_1082,N_49883,N_49818);
and UO_1083 (O_1083,N_49976,N_49890);
nor UO_1084 (O_1084,N_49785,N_49810);
and UO_1085 (O_1085,N_49947,N_49850);
nor UO_1086 (O_1086,N_49918,N_49992);
nand UO_1087 (O_1087,N_49879,N_49856);
nand UO_1088 (O_1088,N_49859,N_49927);
xnor UO_1089 (O_1089,N_49793,N_49931);
nor UO_1090 (O_1090,N_49994,N_49769);
nand UO_1091 (O_1091,N_49980,N_49972);
nand UO_1092 (O_1092,N_49788,N_49956);
nor UO_1093 (O_1093,N_49804,N_49945);
nand UO_1094 (O_1094,N_49961,N_49786);
nand UO_1095 (O_1095,N_49773,N_49922);
xor UO_1096 (O_1096,N_49892,N_49899);
nor UO_1097 (O_1097,N_49889,N_49830);
xnor UO_1098 (O_1098,N_49779,N_49931);
and UO_1099 (O_1099,N_49971,N_49905);
nand UO_1100 (O_1100,N_49864,N_49915);
nor UO_1101 (O_1101,N_49907,N_49938);
and UO_1102 (O_1102,N_49966,N_49801);
or UO_1103 (O_1103,N_49807,N_49925);
or UO_1104 (O_1104,N_49953,N_49947);
nor UO_1105 (O_1105,N_49759,N_49798);
xor UO_1106 (O_1106,N_49903,N_49915);
xor UO_1107 (O_1107,N_49924,N_49825);
nor UO_1108 (O_1108,N_49917,N_49829);
and UO_1109 (O_1109,N_49843,N_49886);
xnor UO_1110 (O_1110,N_49786,N_49822);
nor UO_1111 (O_1111,N_49926,N_49896);
nor UO_1112 (O_1112,N_49791,N_49911);
nand UO_1113 (O_1113,N_49884,N_49929);
xnor UO_1114 (O_1114,N_49879,N_49868);
nand UO_1115 (O_1115,N_49875,N_49904);
and UO_1116 (O_1116,N_49840,N_49854);
or UO_1117 (O_1117,N_49896,N_49904);
xnor UO_1118 (O_1118,N_49833,N_49802);
nor UO_1119 (O_1119,N_49753,N_49895);
or UO_1120 (O_1120,N_49781,N_49789);
and UO_1121 (O_1121,N_49966,N_49992);
or UO_1122 (O_1122,N_49834,N_49784);
and UO_1123 (O_1123,N_49779,N_49918);
xor UO_1124 (O_1124,N_49941,N_49831);
and UO_1125 (O_1125,N_49860,N_49920);
and UO_1126 (O_1126,N_49839,N_49759);
and UO_1127 (O_1127,N_49829,N_49818);
and UO_1128 (O_1128,N_49845,N_49872);
or UO_1129 (O_1129,N_49840,N_49765);
xnor UO_1130 (O_1130,N_49778,N_49936);
or UO_1131 (O_1131,N_49909,N_49797);
and UO_1132 (O_1132,N_49865,N_49988);
or UO_1133 (O_1133,N_49842,N_49838);
nor UO_1134 (O_1134,N_49825,N_49761);
or UO_1135 (O_1135,N_49796,N_49812);
xnor UO_1136 (O_1136,N_49942,N_49875);
nor UO_1137 (O_1137,N_49926,N_49848);
or UO_1138 (O_1138,N_49981,N_49966);
nand UO_1139 (O_1139,N_49824,N_49901);
nor UO_1140 (O_1140,N_49822,N_49928);
nor UO_1141 (O_1141,N_49907,N_49789);
xor UO_1142 (O_1142,N_49771,N_49857);
xor UO_1143 (O_1143,N_49979,N_49856);
and UO_1144 (O_1144,N_49854,N_49900);
and UO_1145 (O_1145,N_49795,N_49884);
nand UO_1146 (O_1146,N_49956,N_49994);
or UO_1147 (O_1147,N_49961,N_49764);
nand UO_1148 (O_1148,N_49794,N_49859);
xnor UO_1149 (O_1149,N_49796,N_49917);
or UO_1150 (O_1150,N_49884,N_49876);
xnor UO_1151 (O_1151,N_49811,N_49840);
nand UO_1152 (O_1152,N_49775,N_49946);
or UO_1153 (O_1153,N_49967,N_49857);
nor UO_1154 (O_1154,N_49936,N_49949);
or UO_1155 (O_1155,N_49896,N_49941);
nor UO_1156 (O_1156,N_49796,N_49851);
or UO_1157 (O_1157,N_49946,N_49831);
nor UO_1158 (O_1158,N_49988,N_49824);
and UO_1159 (O_1159,N_49833,N_49975);
xnor UO_1160 (O_1160,N_49994,N_49800);
and UO_1161 (O_1161,N_49754,N_49784);
nor UO_1162 (O_1162,N_49885,N_49898);
nor UO_1163 (O_1163,N_49968,N_49982);
nor UO_1164 (O_1164,N_49869,N_49803);
nor UO_1165 (O_1165,N_49985,N_49968);
xnor UO_1166 (O_1166,N_49827,N_49971);
nand UO_1167 (O_1167,N_49956,N_49850);
and UO_1168 (O_1168,N_49861,N_49941);
nor UO_1169 (O_1169,N_49829,N_49870);
nor UO_1170 (O_1170,N_49926,N_49808);
and UO_1171 (O_1171,N_49818,N_49985);
nor UO_1172 (O_1172,N_49908,N_49896);
and UO_1173 (O_1173,N_49821,N_49875);
xnor UO_1174 (O_1174,N_49926,N_49897);
or UO_1175 (O_1175,N_49970,N_49757);
xor UO_1176 (O_1176,N_49872,N_49996);
and UO_1177 (O_1177,N_49913,N_49863);
nor UO_1178 (O_1178,N_49805,N_49798);
nor UO_1179 (O_1179,N_49839,N_49976);
xor UO_1180 (O_1180,N_49815,N_49935);
and UO_1181 (O_1181,N_49871,N_49763);
xor UO_1182 (O_1182,N_49817,N_49897);
and UO_1183 (O_1183,N_49961,N_49883);
xnor UO_1184 (O_1184,N_49812,N_49934);
nand UO_1185 (O_1185,N_49858,N_49964);
nand UO_1186 (O_1186,N_49971,N_49931);
xnor UO_1187 (O_1187,N_49756,N_49810);
and UO_1188 (O_1188,N_49869,N_49818);
xor UO_1189 (O_1189,N_49782,N_49927);
or UO_1190 (O_1190,N_49769,N_49926);
or UO_1191 (O_1191,N_49892,N_49992);
or UO_1192 (O_1192,N_49954,N_49810);
xor UO_1193 (O_1193,N_49942,N_49874);
xnor UO_1194 (O_1194,N_49991,N_49993);
or UO_1195 (O_1195,N_49947,N_49758);
or UO_1196 (O_1196,N_49931,N_49877);
nand UO_1197 (O_1197,N_49784,N_49981);
xor UO_1198 (O_1198,N_49914,N_49759);
and UO_1199 (O_1199,N_49758,N_49862);
nor UO_1200 (O_1200,N_49944,N_49897);
xnor UO_1201 (O_1201,N_49794,N_49994);
and UO_1202 (O_1202,N_49957,N_49814);
nor UO_1203 (O_1203,N_49778,N_49875);
nor UO_1204 (O_1204,N_49960,N_49834);
nor UO_1205 (O_1205,N_49881,N_49953);
xor UO_1206 (O_1206,N_49875,N_49985);
xnor UO_1207 (O_1207,N_49959,N_49967);
or UO_1208 (O_1208,N_49852,N_49778);
or UO_1209 (O_1209,N_49775,N_49941);
nand UO_1210 (O_1210,N_49931,N_49883);
nand UO_1211 (O_1211,N_49767,N_49911);
nor UO_1212 (O_1212,N_49769,N_49866);
or UO_1213 (O_1213,N_49797,N_49857);
and UO_1214 (O_1214,N_49986,N_49954);
xor UO_1215 (O_1215,N_49794,N_49983);
or UO_1216 (O_1216,N_49776,N_49949);
xor UO_1217 (O_1217,N_49801,N_49842);
nor UO_1218 (O_1218,N_49896,N_49861);
and UO_1219 (O_1219,N_49883,N_49948);
nand UO_1220 (O_1220,N_49842,N_49836);
xor UO_1221 (O_1221,N_49954,N_49869);
and UO_1222 (O_1222,N_49785,N_49862);
nor UO_1223 (O_1223,N_49853,N_49794);
and UO_1224 (O_1224,N_49753,N_49765);
or UO_1225 (O_1225,N_49905,N_49823);
and UO_1226 (O_1226,N_49821,N_49919);
or UO_1227 (O_1227,N_49996,N_49756);
nand UO_1228 (O_1228,N_49949,N_49810);
nand UO_1229 (O_1229,N_49773,N_49954);
or UO_1230 (O_1230,N_49824,N_49916);
xor UO_1231 (O_1231,N_49889,N_49796);
or UO_1232 (O_1232,N_49848,N_49762);
or UO_1233 (O_1233,N_49787,N_49892);
xnor UO_1234 (O_1234,N_49907,N_49989);
nand UO_1235 (O_1235,N_49929,N_49905);
nor UO_1236 (O_1236,N_49957,N_49795);
or UO_1237 (O_1237,N_49974,N_49918);
xnor UO_1238 (O_1238,N_49819,N_49967);
xnor UO_1239 (O_1239,N_49772,N_49987);
nor UO_1240 (O_1240,N_49771,N_49993);
nand UO_1241 (O_1241,N_49916,N_49840);
nor UO_1242 (O_1242,N_49800,N_49853);
nand UO_1243 (O_1243,N_49929,N_49945);
and UO_1244 (O_1244,N_49753,N_49879);
nand UO_1245 (O_1245,N_49827,N_49751);
xor UO_1246 (O_1246,N_49996,N_49939);
nand UO_1247 (O_1247,N_49875,N_49987);
and UO_1248 (O_1248,N_49854,N_49764);
and UO_1249 (O_1249,N_49967,N_49759);
nor UO_1250 (O_1250,N_49946,N_49806);
or UO_1251 (O_1251,N_49987,N_49852);
nand UO_1252 (O_1252,N_49917,N_49865);
and UO_1253 (O_1253,N_49879,N_49957);
or UO_1254 (O_1254,N_49753,N_49785);
nor UO_1255 (O_1255,N_49946,N_49816);
and UO_1256 (O_1256,N_49895,N_49754);
nor UO_1257 (O_1257,N_49861,N_49810);
nand UO_1258 (O_1258,N_49937,N_49965);
nor UO_1259 (O_1259,N_49787,N_49751);
xnor UO_1260 (O_1260,N_49766,N_49872);
nor UO_1261 (O_1261,N_49877,N_49891);
and UO_1262 (O_1262,N_49924,N_49796);
xor UO_1263 (O_1263,N_49955,N_49864);
and UO_1264 (O_1264,N_49858,N_49892);
nand UO_1265 (O_1265,N_49920,N_49810);
or UO_1266 (O_1266,N_49903,N_49862);
and UO_1267 (O_1267,N_49907,N_49808);
nor UO_1268 (O_1268,N_49771,N_49938);
nand UO_1269 (O_1269,N_49972,N_49903);
nand UO_1270 (O_1270,N_49766,N_49822);
nand UO_1271 (O_1271,N_49861,N_49771);
xor UO_1272 (O_1272,N_49774,N_49916);
and UO_1273 (O_1273,N_49938,N_49889);
nor UO_1274 (O_1274,N_49922,N_49904);
xnor UO_1275 (O_1275,N_49791,N_49782);
or UO_1276 (O_1276,N_49856,N_49944);
xnor UO_1277 (O_1277,N_49898,N_49909);
and UO_1278 (O_1278,N_49804,N_49854);
or UO_1279 (O_1279,N_49817,N_49966);
xor UO_1280 (O_1280,N_49939,N_49782);
nor UO_1281 (O_1281,N_49855,N_49752);
nor UO_1282 (O_1282,N_49766,N_49990);
or UO_1283 (O_1283,N_49817,N_49955);
nand UO_1284 (O_1284,N_49809,N_49918);
nor UO_1285 (O_1285,N_49988,N_49899);
nand UO_1286 (O_1286,N_49826,N_49979);
nand UO_1287 (O_1287,N_49982,N_49974);
xor UO_1288 (O_1288,N_49890,N_49913);
or UO_1289 (O_1289,N_49981,N_49785);
or UO_1290 (O_1290,N_49772,N_49866);
xnor UO_1291 (O_1291,N_49966,N_49777);
nor UO_1292 (O_1292,N_49906,N_49921);
nor UO_1293 (O_1293,N_49815,N_49950);
nor UO_1294 (O_1294,N_49786,N_49887);
xnor UO_1295 (O_1295,N_49964,N_49751);
nor UO_1296 (O_1296,N_49794,N_49855);
nor UO_1297 (O_1297,N_49966,N_49940);
or UO_1298 (O_1298,N_49910,N_49846);
nor UO_1299 (O_1299,N_49923,N_49774);
and UO_1300 (O_1300,N_49872,N_49914);
or UO_1301 (O_1301,N_49772,N_49812);
xnor UO_1302 (O_1302,N_49797,N_49802);
nor UO_1303 (O_1303,N_49977,N_49808);
and UO_1304 (O_1304,N_49788,N_49909);
and UO_1305 (O_1305,N_49996,N_49776);
and UO_1306 (O_1306,N_49979,N_49892);
nor UO_1307 (O_1307,N_49807,N_49904);
nand UO_1308 (O_1308,N_49783,N_49918);
or UO_1309 (O_1309,N_49874,N_49779);
xnor UO_1310 (O_1310,N_49856,N_49868);
nand UO_1311 (O_1311,N_49856,N_49970);
or UO_1312 (O_1312,N_49767,N_49836);
xnor UO_1313 (O_1313,N_49799,N_49886);
nor UO_1314 (O_1314,N_49777,N_49798);
nand UO_1315 (O_1315,N_49860,N_49886);
nand UO_1316 (O_1316,N_49919,N_49780);
xnor UO_1317 (O_1317,N_49853,N_49856);
nor UO_1318 (O_1318,N_49981,N_49884);
or UO_1319 (O_1319,N_49799,N_49790);
and UO_1320 (O_1320,N_49863,N_49932);
nand UO_1321 (O_1321,N_49782,N_49893);
and UO_1322 (O_1322,N_49907,N_49795);
xor UO_1323 (O_1323,N_49854,N_49950);
xnor UO_1324 (O_1324,N_49958,N_49974);
nand UO_1325 (O_1325,N_49885,N_49925);
xor UO_1326 (O_1326,N_49932,N_49820);
nand UO_1327 (O_1327,N_49879,N_49787);
or UO_1328 (O_1328,N_49921,N_49923);
or UO_1329 (O_1329,N_49755,N_49865);
nand UO_1330 (O_1330,N_49933,N_49845);
xnor UO_1331 (O_1331,N_49908,N_49763);
and UO_1332 (O_1332,N_49765,N_49989);
and UO_1333 (O_1333,N_49784,N_49836);
xor UO_1334 (O_1334,N_49788,N_49844);
nand UO_1335 (O_1335,N_49818,N_49888);
nor UO_1336 (O_1336,N_49905,N_49767);
and UO_1337 (O_1337,N_49882,N_49858);
xor UO_1338 (O_1338,N_49895,N_49991);
nand UO_1339 (O_1339,N_49980,N_49933);
and UO_1340 (O_1340,N_49944,N_49921);
and UO_1341 (O_1341,N_49940,N_49995);
nor UO_1342 (O_1342,N_49796,N_49770);
xor UO_1343 (O_1343,N_49781,N_49848);
nand UO_1344 (O_1344,N_49852,N_49947);
or UO_1345 (O_1345,N_49844,N_49861);
nand UO_1346 (O_1346,N_49989,N_49849);
nor UO_1347 (O_1347,N_49857,N_49762);
nand UO_1348 (O_1348,N_49788,N_49935);
or UO_1349 (O_1349,N_49817,N_49871);
nand UO_1350 (O_1350,N_49907,N_49900);
and UO_1351 (O_1351,N_49937,N_49797);
nor UO_1352 (O_1352,N_49921,N_49953);
and UO_1353 (O_1353,N_49954,N_49934);
and UO_1354 (O_1354,N_49784,N_49760);
or UO_1355 (O_1355,N_49884,N_49963);
nor UO_1356 (O_1356,N_49813,N_49984);
nor UO_1357 (O_1357,N_49855,N_49859);
and UO_1358 (O_1358,N_49846,N_49872);
and UO_1359 (O_1359,N_49768,N_49838);
nand UO_1360 (O_1360,N_49788,N_49887);
nand UO_1361 (O_1361,N_49989,N_49883);
and UO_1362 (O_1362,N_49938,N_49783);
and UO_1363 (O_1363,N_49842,N_49775);
nor UO_1364 (O_1364,N_49774,N_49827);
and UO_1365 (O_1365,N_49842,N_49942);
xnor UO_1366 (O_1366,N_49859,N_49862);
xnor UO_1367 (O_1367,N_49803,N_49946);
nand UO_1368 (O_1368,N_49777,N_49769);
and UO_1369 (O_1369,N_49767,N_49843);
and UO_1370 (O_1370,N_49828,N_49951);
or UO_1371 (O_1371,N_49886,N_49935);
nand UO_1372 (O_1372,N_49859,N_49916);
nor UO_1373 (O_1373,N_49951,N_49925);
nand UO_1374 (O_1374,N_49921,N_49788);
and UO_1375 (O_1375,N_49930,N_49921);
xnor UO_1376 (O_1376,N_49938,N_49824);
nand UO_1377 (O_1377,N_49977,N_49852);
or UO_1378 (O_1378,N_49814,N_49998);
nand UO_1379 (O_1379,N_49771,N_49798);
or UO_1380 (O_1380,N_49875,N_49939);
or UO_1381 (O_1381,N_49787,N_49902);
nand UO_1382 (O_1382,N_49892,N_49770);
or UO_1383 (O_1383,N_49915,N_49757);
or UO_1384 (O_1384,N_49768,N_49751);
nand UO_1385 (O_1385,N_49807,N_49839);
and UO_1386 (O_1386,N_49766,N_49755);
or UO_1387 (O_1387,N_49943,N_49922);
and UO_1388 (O_1388,N_49827,N_49943);
xor UO_1389 (O_1389,N_49986,N_49880);
and UO_1390 (O_1390,N_49854,N_49784);
nand UO_1391 (O_1391,N_49792,N_49899);
or UO_1392 (O_1392,N_49820,N_49951);
xor UO_1393 (O_1393,N_49950,N_49949);
xor UO_1394 (O_1394,N_49967,N_49920);
xor UO_1395 (O_1395,N_49852,N_49796);
or UO_1396 (O_1396,N_49927,N_49987);
nor UO_1397 (O_1397,N_49995,N_49899);
and UO_1398 (O_1398,N_49983,N_49942);
and UO_1399 (O_1399,N_49982,N_49938);
nor UO_1400 (O_1400,N_49891,N_49868);
nand UO_1401 (O_1401,N_49835,N_49887);
xnor UO_1402 (O_1402,N_49801,N_49785);
xnor UO_1403 (O_1403,N_49931,N_49885);
or UO_1404 (O_1404,N_49999,N_49958);
and UO_1405 (O_1405,N_49803,N_49874);
and UO_1406 (O_1406,N_49877,N_49800);
nand UO_1407 (O_1407,N_49803,N_49873);
and UO_1408 (O_1408,N_49905,N_49947);
nor UO_1409 (O_1409,N_49880,N_49793);
nor UO_1410 (O_1410,N_49859,N_49846);
nor UO_1411 (O_1411,N_49822,N_49905);
nand UO_1412 (O_1412,N_49931,N_49936);
nand UO_1413 (O_1413,N_49851,N_49937);
nand UO_1414 (O_1414,N_49950,N_49881);
or UO_1415 (O_1415,N_49756,N_49834);
or UO_1416 (O_1416,N_49923,N_49853);
xnor UO_1417 (O_1417,N_49796,N_49936);
nand UO_1418 (O_1418,N_49958,N_49981);
nor UO_1419 (O_1419,N_49961,N_49884);
nor UO_1420 (O_1420,N_49862,N_49786);
nand UO_1421 (O_1421,N_49833,N_49945);
nand UO_1422 (O_1422,N_49796,N_49938);
and UO_1423 (O_1423,N_49824,N_49979);
xor UO_1424 (O_1424,N_49806,N_49881);
xnor UO_1425 (O_1425,N_49871,N_49833);
xnor UO_1426 (O_1426,N_49875,N_49862);
or UO_1427 (O_1427,N_49817,N_49799);
and UO_1428 (O_1428,N_49869,N_49887);
and UO_1429 (O_1429,N_49964,N_49992);
and UO_1430 (O_1430,N_49845,N_49963);
and UO_1431 (O_1431,N_49932,N_49836);
nor UO_1432 (O_1432,N_49821,N_49974);
nand UO_1433 (O_1433,N_49848,N_49927);
xor UO_1434 (O_1434,N_49965,N_49763);
nand UO_1435 (O_1435,N_49876,N_49897);
nor UO_1436 (O_1436,N_49999,N_49925);
nor UO_1437 (O_1437,N_49932,N_49879);
xor UO_1438 (O_1438,N_49922,N_49769);
nor UO_1439 (O_1439,N_49760,N_49940);
or UO_1440 (O_1440,N_49975,N_49767);
nor UO_1441 (O_1441,N_49997,N_49829);
or UO_1442 (O_1442,N_49850,N_49983);
xnor UO_1443 (O_1443,N_49986,N_49961);
nor UO_1444 (O_1444,N_49754,N_49924);
and UO_1445 (O_1445,N_49999,N_49802);
nor UO_1446 (O_1446,N_49799,N_49944);
and UO_1447 (O_1447,N_49756,N_49933);
and UO_1448 (O_1448,N_49783,N_49985);
or UO_1449 (O_1449,N_49801,N_49874);
and UO_1450 (O_1450,N_49854,N_49908);
nor UO_1451 (O_1451,N_49794,N_49901);
nor UO_1452 (O_1452,N_49852,N_49953);
nand UO_1453 (O_1453,N_49956,N_49826);
and UO_1454 (O_1454,N_49847,N_49973);
nor UO_1455 (O_1455,N_49857,N_49988);
nor UO_1456 (O_1456,N_49909,N_49937);
nor UO_1457 (O_1457,N_49922,N_49940);
and UO_1458 (O_1458,N_49820,N_49801);
nor UO_1459 (O_1459,N_49983,N_49814);
nor UO_1460 (O_1460,N_49862,N_49962);
xnor UO_1461 (O_1461,N_49902,N_49809);
or UO_1462 (O_1462,N_49850,N_49776);
and UO_1463 (O_1463,N_49909,N_49869);
nor UO_1464 (O_1464,N_49957,N_49846);
or UO_1465 (O_1465,N_49819,N_49840);
and UO_1466 (O_1466,N_49783,N_49933);
nand UO_1467 (O_1467,N_49968,N_49969);
and UO_1468 (O_1468,N_49849,N_49943);
xor UO_1469 (O_1469,N_49785,N_49991);
nor UO_1470 (O_1470,N_49854,N_49834);
or UO_1471 (O_1471,N_49763,N_49985);
or UO_1472 (O_1472,N_49757,N_49828);
xnor UO_1473 (O_1473,N_49856,N_49947);
nand UO_1474 (O_1474,N_49974,N_49891);
nor UO_1475 (O_1475,N_49949,N_49838);
nand UO_1476 (O_1476,N_49984,N_49893);
nor UO_1477 (O_1477,N_49974,N_49921);
nor UO_1478 (O_1478,N_49958,N_49946);
xor UO_1479 (O_1479,N_49897,N_49919);
or UO_1480 (O_1480,N_49949,N_49756);
xor UO_1481 (O_1481,N_49952,N_49950);
or UO_1482 (O_1482,N_49928,N_49816);
nor UO_1483 (O_1483,N_49837,N_49977);
nand UO_1484 (O_1484,N_49903,N_49963);
or UO_1485 (O_1485,N_49919,N_49911);
xor UO_1486 (O_1486,N_49785,N_49853);
nor UO_1487 (O_1487,N_49824,N_49887);
xnor UO_1488 (O_1488,N_49843,N_49874);
nand UO_1489 (O_1489,N_49768,N_49810);
and UO_1490 (O_1490,N_49841,N_49999);
xnor UO_1491 (O_1491,N_49845,N_49917);
xnor UO_1492 (O_1492,N_49952,N_49860);
xnor UO_1493 (O_1493,N_49976,N_49772);
or UO_1494 (O_1494,N_49770,N_49902);
nand UO_1495 (O_1495,N_49892,N_49926);
nor UO_1496 (O_1496,N_49871,N_49872);
and UO_1497 (O_1497,N_49848,N_49936);
xnor UO_1498 (O_1498,N_49779,N_49859);
and UO_1499 (O_1499,N_49975,N_49979);
or UO_1500 (O_1500,N_49909,N_49953);
and UO_1501 (O_1501,N_49853,N_49845);
xnor UO_1502 (O_1502,N_49881,N_49906);
and UO_1503 (O_1503,N_49920,N_49896);
xor UO_1504 (O_1504,N_49969,N_49963);
or UO_1505 (O_1505,N_49992,N_49891);
and UO_1506 (O_1506,N_49978,N_49929);
or UO_1507 (O_1507,N_49877,N_49848);
or UO_1508 (O_1508,N_49933,N_49811);
or UO_1509 (O_1509,N_49931,N_49771);
nor UO_1510 (O_1510,N_49901,N_49876);
and UO_1511 (O_1511,N_49871,N_49919);
nand UO_1512 (O_1512,N_49911,N_49932);
or UO_1513 (O_1513,N_49884,N_49819);
xnor UO_1514 (O_1514,N_49761,N_49908);
xnor UO_1515 (O_1515,N_49925,N_49802);
xor UO_1516 (O_1516,N_49789,N_49808);
xor UO_1517 (O_1517,N_49932,N_49852);
nand UO_1518 (O_1518,N_49922,N_49884);
or UO_1519 (O_1519,N_49894,N_49773);
and UO_1520 (O_1520,N_49948,N_49768);
and UO_1521 (O_1521,N_49847,N_49873);
and UO_1522 (O_1522,N_49820,N_49780);
nand UO_1523 (O_1523,N_49935,N_49798);
xnor UO_1524 (O_1524,N_49876,N_49889);
and UO_1525 (O_1525,N_49825,N_49925);
and UO_1526 (O_1526,N_49752,N_49814);
and UO_1527 (O_1527,N_49922,N_49809);
or UO_1528 (O_1528,N_49945,N_49756);
or UO_1529 (O_1529,N_49932,N_49855);
xnor UO_1530 (O_1530,N_49814,N_49923);
or UO_1531 (O_1531,N_49752,N_49765);
nor UO_1532 (O_1532,N_49993,N_49959);
xor UO_1533 (O_1533,N_49815,N_49760);
nor UO_1534 (O_1534,N_49871,N_49868);
xnor UO_1535 (O_1535,N_49945,N_49967);
and UO_1536 (O_1536,N_49770,N_49774);
xor UO_1537 (O_1537,N_49946,N_49755);
xnor UO_1538 (O_1538,N_49959,N_49859);
and UO_1539 (O_1539,N_49964,N_49948);
or UO_1540 (O_1540,N_49959,N_49788);
or UO_1541 (O_1541,N_49863,N_49936);
and UO_1542 (O_1542,N_49871,N_49760);
and UO_1543 (O_1543,N_49844,N_49916);
xnor UO_1544 (O_1544,N_49972,N_49754);
xnor UO_1545 (O_1545,N_49937,N_49871);
xnor UO_1546 (O_1546,N_49759,N_49892);
nor UO_1547 (O_1547,N_49944,N_49977);
or UO_1548 (O_1548,N_49782,N_49972);
and UO_1549 (O_1549,N_49846,N_49955);
and UO_1550 (O_1550,N_49999,N_49812);
nand UO_1551 (O_1551,N_49903,N_49925);
xnor UO_1552 (O_1552,N_49833,N_49790);
nor UO_1553 (O_1553,N_49827,N_49765);
or UO_1554 (O_1554,N_49986,N_49818);
or UO_1555 (O_1555,N_49787,N_49769);
or UO_1556 (O_1556,N_49892,N_49928);
nor UO_1557 (O_1557,N_49984,N_49902);
and UO_1558 (O_1558,N_49890,N_49825);
or UO_1559 (O_1559,N_49850,N_49888);
nor UO_1560 (O_1560,N_49981,N_49868);
xnor UO_1561 (O_1561,N_49806,N_49836);
nor UO_1562 (O_1562,N_49803,N_49798);
nor UO_1563 (O_1563,N_49892,N_49798);
nor UO_1564 (O_1564,N_49780,N_49834);
nor UO_1565 (O_1565,N_49767,N_49890);
nor UO_1566 (O_1566,N_49750,N_49819);
nand UO_1567 (O_1567,N_49831,N_49923);
nor UO_1568 (O_1568,N_49770,N_49884);
and UO_1569 (O_1569,N_49885,N_49765);
nor UO_1570 (O_1570,N_49805,N_49893);
and UO_1571 (O_1571,N_49816,N_49806);
and UO_1572 (O_1572,N_49799,N_49798);
and UO_1573 (O_1573,N_49897,N_49832);
nand UO_1574 (O_1574,N_49950,N_49793);
or UO_1575 (O_1575,N_49797,N_49804);
and UO_1576 (O_1576,N_49874,N_49889);
xor UO_1577 (O_1577,N_49964,N_49874);
xor UO_1578 (O_1578,N_49937,N_49914);
or UO_1579 (O_1579,N_49841,N_49942);
nor UO_1580 (O_1580,N_49936,N_49797);
or UO_1581 (O_1581,N_49941,N_49777);
or UO_1582 (O_1582,N_49788,N_49995);
nor UO_1583 (O_1583,N_49989,N_49995);
and UO_1584 (O_1584,N_49899,N_49809);
nand UO_1585 (O_1585,N_49823,N_49808);
xnor UO_1586 (O_1586,N_49970,N_49812);
xor UO_1587 (O_1587,N_49963,N_49804);
and UO_1588 (O_1588,N_49809,N_49812);
nand UO_1589 (O_1589,N_49966,N_49835);
nor UO_1590 (O_1590,N_49845,N_49786);
nor UO_1591 (O_1591,N_49784,N_49792);
nand UO_1592 (O_1592,N_49773,N_49858);
nor UO_1593 (O_1593,N_49894,N_49780);
nand UO_1594 (O_1594,N_49765,N_49757);
nand UO_1595 (O_1595,N_49862,N_49898);
or UO_1596 (O_1596,N_49776,N_49972);
or UO_1597 (O_1597,N_49818,N_49990);
nand UO_1598 (O_1598,N_49849,N_49811);
and UO_1599 (O_1599,N_49933,N_49908);
xnor UO_1600 (O_1600,N_49800,N_49999);
nor UO_1601 (O_1601,N_49993,N_49784);
nand UO_1602 (O_1602,N_49858,N_49828);
xnor UO_1603 (O_1603,N_49926,N_49863);
xor UO_1604 (O_1604,N_49885,N_49873);
xnor UO_1605 (O_1605,N_49751,N_49887);
nand UO_1606 (O_1606,N_49797,N_49994);
xor UO_1607 (O_1607,N_49778,N_49944);
nand UO_1608 (O_1608,N_49834,N_49950);
or UO_1609 (O_1609,N_49966,N_49830);
nor UO_1610 (O_1610,N_49862,N_49936);
xnor UO_1611 (O_1611,N_49870,N_49952);
nand UO_1612 (O_1612,N_49844,N_49992);
or UO_1613 (O_1613,N_49903,N_49983);
or UO_1614 (O_1614,N_49756,N_49893);
nor UO_1615 (O_1615,N_49963,N_49801);
xor UO_1616 (O_1616,N_49907,N_49751);
xor UO_1617 (O_1617,N_49894,N_49806);
nor UO_1618 (O_1618,N_49843,N_49856);
nor UO_1619 (O_1619,N_49955,N_49943);
nor UO_1620 (O_1620,N_49780,N_49777);
nor UO_1621 (O_1621,N_49981,N_49859);
and UO_1622 (O_1622,N_49941,N_49894);
and UO_1623 (O_1623,N_49893,N_49829);
nand UO_1624 (O_1624,N_49775,N_49778);
nor UO_1625 (O_1625,N_49924,N_49933);
or UO_1626 (O_1626,N_49801,N_49811);
or UO_1627 (O_1627,N_49800,N_49801);
nand UO_1628 (O_1628,N_49847,N_49799);
nand UO_1629 (O_1629,N_49851,N_49789);
xor UO_1630 (O_1630,N_49988,N_49914);
nand UO_1631 (O_1631,N_49845,N_49798);
nor UO_1632 (O_1632,N_49949,N_49845);
or UO_1633 (O_1633,N_49888,N_49787);
and UO_1634 (O_1634,N_49965,N_49868);
nor UO_1635 (O_1635,N_49826,N_49824);
nor UO_1636 (O_1636,N_49890,N_49843);
xnor UO_1637 (O_1637,N_49782,N_49971);
and UO_1638 (O_1638,N_49978,N_49996);
and UO_1639 (O_1639,N_49834,N_49833);
or UO_1640 (O_1640,N_49804,N_49917);
nor UO_1641 (O_1641,N_49827,N_49914);
or UO_1642 (O_1642,N_49863,N_49991);
xnor UO_1643 (O_1643,N_49902,N_49866);
nand UO_1644 (O_1644,N_49838,N_49827);
xnor UO_1645 (O_1645,N_49922,N_49925);
and UO_1646 (O_1646,N_49885,N_49792);
or UO_1647 (O_1647,N_49957,N_49990);
xor UO_1648 (O_1648,N_49779,N_49771);
or UO_1649 (O_1649,N_49816,N_49929);
or UO_1650 (O_1650,N_49763,N_49912);
nand UO_1651 (O_1651,N_49940,N_49970);
nand UO_1652 (O_1652,N_49936,N_49782);
xnor UO_1653 (O_1653,N_49837,N_49995);
or UO_1654 (O_1654,N_49939,N_49956);
nor UO_1655 (O_1655,N_49976,N_49936);
or UO_1656 (O_1656,N_49987,N_49903);
xor UO_1657 (O_1657,N_49967,N_49893);
or UO_1658 (O_1658,N_49827,N_49824);
or UO_1659 (O_1659,N_49787,N_49773);
nand UO_1660 (O_1660,N_49920,N_49877);
nor UO_1661 (O_1661,N_49772,N_49977);
xnor UO_1662 (O_1662,N_49979,N_49827);
nor UO_1663 (O_1663,N_49759,N_49874);
xor UO_1664 (O_1664,N_49938,N_49926);
and UO_1665 (O_1665,N_49845,N_49979);
nand UO_1666 (O_1666,N_49790,N_49841);
xnor UO_1667 (O_1667,N_49992,N_49856);
nor UO_1668 (O_1668,N_49910,N_49824);
or UO_1669 (O_1669,N_49751,N_49932);
and UO_1670 (O_1670,N_49833,N_49788);
nor UO_1671 (O_1671,N_49822,N_49873);
and UO_1672 (O_1672,N_49809,N_49947);
or UO_1673 (O_1673,N_49755,N_49762);
nor UO_1674 (O_1674,N_49824,N_49915);
nand UO_1675 (O_1675,N_49871,N_49879);
or UO_1676 (O_1676,N_49897,N_49847);
and UO_1677 (O_1677,N_49943,N_49750);
and UO_1678 (O_1678,N_49837,N_49836);
nor UO_1679 (O_1679,N_49934,N_49838);
nor UO_1680 (O_1680,N_49918,N_49857);
nand UO_1681 (O_1681,N_49888,N_49803);
xor UO_1682 (O_1682,N_49982,N_49858);
and UO_1683 (O_1683,N_49973,N_49820);
and UO_1684 (O_1684,N_49998,N_49874);
and UO_1685 (O_1685,N_49858,N_49802);
nand UO_1686 (O_1686,N_49964,N_49774);
or UO_1687 (O_1687,N_49879,N_49858);
nand UO_1688 (O_1688,N_49766,N_49992);
nor UO_1689 (O_1689,N_49785,N_49880);
and UO_1690 (O_1690,N_49977,N_49947);
and UO_1691 (O_1691,N_49878,N_49843);
xor UO_1692 (O_1692,N_49850,N_49972);
nor UO_1693 (O_1693,N_49770,N_49893);
and UO_1694 (O_1694,N_49794,N_49981);
nand UO_1695 (O_1695,N_49826,N_49750);
nand UO_1696 (O_1696,N_49858,N_49943);
or UO_1697 (O_1697,N_49970,N_49811);
and UO_1698 (O_1698,N_49978,N_49828);
nand UO_1699 (O_1699,N_49760,N_49946);
nand UO_1700 (O_1700,N_49949,N_49789);
and UO_1701 (O_1701,N_49974,N_49826);
nor UO_1702 (O_1702,N_49808,N_49876);
xor UO_1703 (O_1703,N_49897,N_49880);
or UO_1704 (O_1704,N_49858,N_49942);
nor UO_1705 (O_1705,N_49885,N_49995);
nor UO_1706 (O_1706,N_49855,N_49764);
xnor UO_1707 (O_1707,N_49893,N_49906);
and UO_1708 (O_1708,N_49902,N_49773);
nand UO_1709 (O_1709,N_49895,N_49870);
nand UO_1710 (O_1710,N_49825,N_49982);
xnor UO_1711 (O_1711,N_49772,N_49831);
nand UO_1712 (O_1712,N_49868,N_49949);
and UO_1713 (O_1713,N_49803,N_49922);
xor UO_1714 (O_1714,N_49989,N_49750);
xnor UO_1715 (O_1715,N_49913,N_49857);
nor UO_1716 (O_1716,N_49804,N_49751);
xor UO_1717 (O_1717,N_49873,N_49764);
xnor UO_1718 (O_1718,N_49792,N_49812);
xor UO_1719 (O_1719,N_49926,N_49812);
nand UO_1720 (O_1720,N_49821,N_49936);
xnor UO_1721 (O_1721,N_49988,N_49989);
xnor UO_1722 (O_1722,N_49963,N_49896);
and UO_1723 (O_1723,N_49804,N_49811);
and UO_1724 (O_1724,N_49978,N_49758);
and UO_1725 (O_1725,N_49864,N_49908);
and UO_1726 (O_1726,N_49879,N_49848);
xor UO_1727 (O_1727,N_49999,N_49951);
nand UO_1728 (O_1728,N_49801,N_49885);
xor UO_1729 (O_1729,N_49898,N_49860);
and UO_1730 (O_1730,N_49989,N_49816);
xnor UO_1731 (O_1731,N_49832,N_49778);
or UO_1732 (O_1732,N_49820,N_49806);
nor UO_1733 (O_1733,N_49892,N_49935);
xnor UO_1734 (O_1734,N_49987,N_49988);
nand UO_1735 (O_1735,N_49955,N_49805);
and UO_1736 (O_1736,N_49844,N_49856);
and UO_1737 (O_1737,N_49783,N_49865);
xnor UO_1738 (O_1738,N_49838,N_49922);
nor UO_1739 (O_1739,N_49893,N_49797);
nor UO_1740 (O_1740,N_49822,N_49988);
nand UO_1741 (O_1741,N_49782,N_49814);
or UO_1742 (O_1742,N_49946,N_49917);
xnor UO_1743 (O_1743,N_49993,N_49854);
and UO_1744 (O_1744,N_49788,N_49853);
nand UO_1745 (O_1745,N_49885,N_49784);
nand UO_1746 (O_1746,N_49995,N_49828);
xnor UO_1747 (O_1747,N_49991,N_49935);
nand UO_1748 (O_1748,N_49967,N_49780);
nor UO_1749 (O_1749,N_49782,N_49834);
xor UO_1750 (O_1750,N_49915,N_49955);
and UO_1751 (O_1751,N_49941,N_49781);
nand UO_1752 (O_1752,N_49790,N_49932);
and UO_1753 (O_1753,N_49859,N_49811);
nor UO_1754 (O_1754,N_49960,N_49917);
nor UO_1755 (O_1755,N_49803,N_49839);
and UO_1756 (O_1756,N_49806,N_49851);
nor UO_1757 (O_1757,N_49788,N_49905);
nand UO_1758 (O_1758,N_49825,N_49754);
or UO_1759 (O_1759,N_49770,N_49838);
or UO_1760 (O_1760,N_49875,N_49869);
or UO_1761 (O_1761,N_49993,N_49905);
and UO_1762 (O_1762,N_49935,N_49906);
nand UO_1763 (O_1763,N_49966,N_49838);
and UO_1764 (O_1764,N_49819,N_49862);
nor UO_1765 (O_1765,N_49939,N_49832);
nor UO_1766 (O_1766,N_49925,N_49877);
nand UO_1767 (O_1767,N_49986,N_49751);
xor UO_1768 (O_1768,N_49845,N_49903);
nand UO_1769 (O_1769,N_49792,N_49795);
nand UO_1770 (O_1770,N_49861,N_49951);
and UO_1771 (O_1771,N_49985,N_49845);
xor UO_1772 (O_1772,N_49888,N_49963);
xor UO_1773 (O_1773,N_49755,N_49971);
xnor UO_1774 (O_1774,N_49875,N_49883);
nor UO_1775 (O_1775,N_49898,N_49790);
xnor UO_1776 (O_1776,N_49943,N_49770);
nand UO_1777 (O_1777,N_49892,N_49972);
xnor UO_1778 (O_1778,N_49817,N_49768);
nand UO_1779 (O_1779,N_49880,N_49755);
nor UO_1780 (O_1780,N_49896,N_49945);
xnor UO_1781 (O_1781,N_49911,N_49872);
and UO_1782 (O_1782,N_49887,N_49989);
or UO_1783 (O_1783,N_49771,N_49810);
nor UO_1784 (O_1784,N_49961,N_49862);
or UO_1785 (O_1785,N_49809,N_49887);
nor UO_1786 (O_1786,N_49884,N_49798);
and UO_1787 (O_1787,N_49935,N_49984);
xor UO_1788 (O_1788,N_49824,N_49836);
nand UO_1789 (O_1789,N_49868,N_49925);
nand UO_1790 (O_1790,N_49869,N_49880);
or UO_1791 (O_1791,N_49942,N_49752);
xor UO_1792 (O_1792,N_49902,N_49964);
xnor UO_1793 (O_1793,N_49797,N_49771);
and UO_1794 (O_1794,N_49976,N_49794);
or UO_1795 (O_1795,N_49810,N_49815);
and UO_1796 (O_1796,N_49922,N_49921);
xor UO_1797 (O_1797,N_49843,N_49866);
nand UO_1798 (O_1798,N_49820,N_49755);
xor UO_1799 (O_1799,N_49834,N_49783);
and UO_1800 (O_1800,N_49960,N_49774);
nand UO_1801 (O_1801,N_49916,N_49852);
xnor UO_1802 (O_1802,N_49969,N_49896);
and UO_1803 (O_1803,N_49923,N_49805);
and UO_1804 (O_1804,N_49799,N_49891);
or UO_1805 (O_1805,N_49845,N_49891);
nor UO_1806 (O_1806,N_49771,N_49997);
nand UO_1807 (O_1807,N_49889,N_49920);
nand UO_1808 (O_1808,N_49944,N_49769);
nor UO_1809 (O_1809,N_49923,N_49955);
xor UO_1810 (O_1810,N_49908,N_49786);
or UO_1811 (O_1811,N_49858,N_49819);
nand UO_1812 (O_1812,N_49947,N_49939);
and UO_1813 (O_1813,N_49840,N_49796);
nor UO_1814 (O_1814,N_49915,N_49952);
and UO_1815 (O_1815,N_49870,N_49990);
and UO_1816 (O_1816,N_49864,N_49865);
nand UO_1817 (O_1817,N_49858,N_49938);
and UO_1818 (O_1818,N_49798,N_49763);
and UO_1819 (O_1819,N_49750,N_49969);
and UO_1820 (O_1820,N_49968,N_49940);
nand UO_1821 (O_1821,N_49866,N_49860);
or UO_1822 (O_1822,N_49790,N_49979);
and UO_1823 (O_1823,N_49950,N_49816);
xnor UO_1824 (O_1824,N_49780,N_49775);
or UO_1825 (O_1825,N_49905,N_49874);
nand UO_1826 (O_1826,N_49954,N_49793);
or UO_1827 (O_1827,N_49934,N_49927);
or UO_1828 (O_1828,N_49806,N_49807);
and UO_1829 (O_1829,N_49929,N_49818);
nand UO_1830 (O_1830,N_49869,N_49917);
xor UO_1831 (O_1831,N_49975,N_49846);
nor UO_1832 (O_1832,N_49868,N_49880);
or UO_1833 (O_1833,N_49919,N_49889);
xnor UO_1834 (O_1834,N_49863,N_49785);
xnor UO_1835 (O_1835,N_49767,N_49949);
nand UO_1836 (O_1836,N_49791,N_49938);
or UO_1837 (O_1837,N_49887,N_49943);
or UO_1838 (O_1838,N_49900,N_49913);
nand UO_1839 (O_1839,N_49877,N_49815);
nor UO_1840 (O_1840,N_49892,N_49957);
or UO_1841 (O_1841,N_49969,N_49825);
or UO_1842 (O_1842,N_49793,N_49873);
or UO_1843 (O_1843,N_49764,N_49928);
and UO_1844 (O_1844,N_49885,N_49827);
nor UO_1845 (O_1845,N_49900,N_49767);
or UO_1846 (O_1846,N_49856,N_49901);
or UO_1847 (O_1847,N_49978,N_49876);
nor UO_1848 (O_1848,N_49859,N_49988);
nand UO_1849 (O_1849,N_49977,N_49754);
xnor UO_1850 (O_1850,N_49755,N_49952);
nand UO_1851 (O_1851,N_49813,N_49945);
and UO_1852 (O_1852,N_49923,N_49764);
nor UO_1853 (O_1853,N_49860,N_49892);
xor UO_1854 (O_1854,N_49765,N_49964);
nor UO_1855 (O_1855,N_49789,N_49836);
nor UO_1856 (O_1856,N_49845,N_49849);
nand UO_1857 (O_1857,N_49861,N_49950);
and UO_1858 (O_1858,N_49977,N_49785);
nor UO_1859 (O_1859,N_49778,N_49972);
and UO_1860 (O_1860,N_49932,N_49908);
nor UO_1861 (O_1861,N_49774,N_49776);
or UO_1862 (O_1862,N_49824,N_49980);
nor UO_1863 (O_1863,N_49976,N_49959);
or UO_1864 (O_1864,N_49856,N_49858);
nand UO_1865 (O_1865,N_49770,N_49939);
nand UO_1866 (O_1866,N_49769,N_49939);
xnor UO_1867 (O_1867,N_49887,N_49787);
and UO_1868 (O_1868,N_49781,N_49896);
and UO_1869 (O_1869,N_49800,N_49926);
xnor UO_1870 (O_1870,N_49892,N_49872);
xnor UO_1871 (O_1871,N_49812,N_49755);
xnor UO_1872 (O_1872,N_49861,N_49862);
nand UO_1873 (O_1873,N_49839,N_49765);
and UO_1874 (O_1874,N_49859,N_49956);
and UO_1875 (O_1875,N_49813,N_49795);
nor UO_1876 (O_1876,N_49969,N_49835);
nor UO_1877 (O_1877,N_49793,N_49778);
nand UO_1878 (O_1878,N_49908,N_49902);
or UO_1879 (O_1879,N_49910,N_49904);
and UO_1880 (O_1880,N_49797,N_49983);
nand UO_1881 (O_1881,N_49824,N_49937);
or UO_1882 (O_1882,N_49880,N_49867);
and UO_1883 (O_1883,N_49794,N_49793);
and UO_1884 (O_1884,N_49820,N_49912);
nand UO_1885 (O_1885,N_49791,N_49750);
or UO_1886 (O_1886,N_49925,N_49856);
or UO_1887 (O_1887,N_49798,N_49917);
nor UO_1888 (O_1888,N_49978,N_49763);
nor UO_1889 (O_1889,N_49838,N_49913);
nor UO_1890 (O_1890,N_49799,N_49771);
nand UO_1891 (O_1891,N_49801,N_49951);
nand UO_1892 (O_1892,N_49753,N_49862);
nand UO_1893 (O_1893,N_49901,N_49863);
or UO_1894 (O_1894,N_49998,N_49769);
xor UO_1895 (O_1895,N_49898,N_49837);
nor UO_1896 (O_1896,N_49839,N_49961);
nand UO_1897 (O_1897,N_49857,N_49977);
or UO_1898 (O_1898,N_49838,N_49893);
nor UO_1899 (O_1899,N_49822,N_49834);
or UO_1900 (O_1900,N_49782,N_49773);
nand UO_1901 (O_1901,N_49915,N_49821);
or UO_1902 (O_1902,N_49781,N_49986);
nand UO_1903 (O_1903,N_49990,N_49964);
nand UO_1904 (O_1904,N_49815,N_49923);
and UO_1905 (O_1905,N_49761,N_49832);
or UO_1906 (O_1906,N_49859,N_49894);
nand UO_1907 (O_1907,N_49909,N_49775);
and UO_1908 (O_1908,N_49999,N_49905);
nand UO_1909 (O_1909,N_49875,N_49783);
nand UO_1910 (O_1910,N_49991,N_49878);
nor UO_1911 (O_1911,N_49988,N_49848);
or UO_1912 (O_1912,N_49981,N_49788);
nand UO_1913 (O_1913,N_49840,N_49772);
or UO_1914 (O_1914,N_49808,N_49827);
nor UO_1915 (O_1915,N_49944,N_49859);
xnor UO_1916 (O_1916,N_49841,N_49923);
or UO_1917 (O_1917,N_49856,N_49780);
xnor UO_1918 (O_1918,N_49833,N_49888);
and UO_1919 (O_1919,N_49957,N_49841);
or UO_1920 (O_1920,N_49969,N_49751);
nand UO_1921 (O_1921,N_49951,N_49932);
nand UO_1922 (O_1922,N_49869,N_49981);
xor UO_1923 (O_1923,N_49916,N_49812);
nand UO_1924 (O_1924,N_49997,N_49927);
nand UO_1925 (O_1925,N_49783,N_49814);
xor UO_1926 (O_1926,N_49802,N_49844);
and UO_1927 (O_1927,N_49907,N_49819);
nor UO_1928 (O_1928,N_49904,N_49873);
xor UO_1929 (O_1929,N_49971,N_49816);
and UO_1930 (O_1930,N_49963,N_49761);
and UO_1931 (O_1931,N_49841,N_49776);
xnor UO_1932 (O_1932,N_49823,N_49856);
xnor UO_1933 (O_1933,N_49865,N_49856);
xnor UO_1934 (O_1934,N_49961,N_49940);
or UO_1935 (O_1935,N_49768,N_49858);
and UO_1936 (O_1936,N_49920,N_49835);
or UO_1937 (O_1937,N_49985,N_49923);
nor UO_1938 (O_1938,N_49830,N_49840);
nand UO_1939 (O_1939,N_49949,N_49941);
and UO_1940 (O_1940,N_49996,N_49989);
and UO_1941 (O_1941,N_49803,N_49835);
nand UO_1942 (O_1942,N_49886,N_49990);
or UO_1943 (O_1943,N_49965,N_49934);
nor UO_1944 (O_1944,N_49829,N_49821);
nand UO_1945 (O_1945,N_49897,N_49905);
nand UO_1946 (O_1946,N_49756,N_49890);
nor UO_1947 (O_1947,N_49912,N_49769);
and UO_1948 (O_1948,N_49939,N_49786);
xnor UO_1949 (O_1949,N_49801,N_49900);
and UO_1950 (O_1950,N_49995,N_49866);
xor UO_1951 (O_1951,N_49810,N_49881);
or UO_1952 (O_1952,N_49982,N_49925);
nor UO_1953 (O_1953,N_49982,N_49766);
or UO_1954 (O_1954,N_49780,N_49925);
nor UO_1955 (O_1955,N_49965,N_49936);
xnor UO_1956 (O_1956,N_49898,N_49919);
or UO_1957 (O_1957,N_49998,N_49796);
nor UO_1958 (O_1958,N_49751,N_49974);
or UO_1959 (O_1959,N_49974,N_49814);
nand UO_1960 (O_1960,N_49912,N_49957);
nor UO_1961 (O_1961,N_49929,N_49914);
xnor UO_1962 (O_1962,N_49828,N_49804);
and UO_1963 (O_1963,N_49790,N_49800);
nand UO_1964 (O_1964,N_49890,N_49796);
or UO_1965 (O_1965,N_49975,N_49755);
xor UO_1966 (O_1966,N_49793,N_49985);
nor UO_1967 (O_1967,N_49867,N_49986);
nor UO_1968 (O_1968,N_49846,N_49797);
nor UO_1969 (O_1969,N_49975,N_49784);
and UO_1970 (O_1970,N_49763,N_49898);
and UO_1971 (O_1971,N_49970,N_49870);
nor UO_1972 (O_1972,N_49932,N_49757);
nor UO_1973 (O_1973,N_49965,N_49771);
xnor UO_1974 (O_1974,N_49819,N_49971);
xor UO_1975 (O_1975,N_49855,N_49805);
nand UO_1976 (O_1976,N_49893,N_49940);
nor UO_1977 (O_1977,N_49829,N_49970);
and UO_1978 (O_1978,N_49859,N_49895);
nor UO_1979 (O_1979,N_49858,N_49771);
or UO_1980 (O_1980,N_49770,N_49854);
nor UO_1981 (O_1981,N_49950,N_49776);
xor UO_1982 (O_1982,N_49991,N_49888);
or UO_1983 (O_1983,N_49950,N_49863);
nand UO_1984 (O_1984,N_49781,N_49752);
and UO_1985 (O_1985,N_49791,N_49956);
or UO_1986 (O_1986,N_49993,N_49811);
and UO_1987 (O_1987,N_49752,N_49760);
xor UO_1988 (O_1988,N_49961,N_49969);
nor UO_1989 (O_1989,N_49755,N_49769);
xor UO_1990 (O_1990,N_49946,N_49759);
nor UO_1991 (O_1991,N_49779,N_49763);
nor UO_1992 (O_1992,N_49892,N_49969);
and UO_1993 (O_1993,N_49988,N_49947);
nand UO_1994 (O_1994,N_49848,N_49768);
and UO_1995 (O_1995,N_49860,N_49837);
or UO_1996 (O_1996,N_49755,N_49877);
nand UO_1997 (O_1997,N_49982,N_49847);
and UO_1998 (O_1998,N_49804,N_49844);
nand UO_1999 (O_1999,N_49899,N_49827);
and UO_2000 (O_2000,N_49767,N_49992);
nand UO_2001 (O_2001,N_49865,N_49760);
or UO_2002 (O_2002,N_49816,N_49797);
nor UO_2003 (O_2003,N_49865,N_49829);
nor UO_2004 (O_2004,N_49919,N_49984);
or UO_2005 (O_2005,N_49897,N_49981);
and UO_2006 (O_2006,N_49936,N_49996);
and UO_2007 (O_2007,N_49960,N_49861);
nand UO_2008 (O_2008,N_49835,N_49796);
or UO_2009 (O_2009,N_49808,N_49878);
or UO_2010 (O_2010,N_49876,N_49783);
nand UO_2011 (O_2011,N_49953,N_49931);
nor UO_2012 (O_2012,N_49755,N_49754);
nor UO_2013 (O_2013,N_49823,N_49794);
or UO_2014 (O_2014,N_49879,N_49822);
nor UO_2015 (O_2015,N_49879,N_49815);
xnor UO_2016 (O_2016,N_49851,N_49860);
or UO_2017 (O_2017,N_49926,N_49961);
xor UO_2018 (O_2018,N_49965,N_49981);
xor UO_2019 (O_2019,N_49939,N_49787);
nand UO_2020 (O_2020,N_49992,N_49789);
and UO_2021 (O_2021,N_49818,N_49970);
nand UO_2022 (O_2022,N_49801,N_49954);
nor UO_2023 (O_2023,N_49866,N_49904);
xor UO_2024 (O_2024,N_49753,N_49757);
and UO_2025 (O_2025,N_49928,N_49802);
or UO_2026 (O_2026,N_49904,N_49869);
or UO_2027 (O_2027,N_49870,N_49760);
and UO_2028 (O_2028,N_49807,N_49890);
xnor UO_2029 (O_2029,N_49810,N_49983);
nor UO_2030 (O_2030,N_49869,N_49782);
or UO_2031 (O_2031,N_49924,N_49897);
and UO_2032 (O_2032,N_49785,N_49962);
or UO_2033 (O_2033,N_49811,N_49943);
nand UO_2034 (O_2034,N_49816,N_49942);
xnor UO_2035 (O_2035,N_49831,N_49791);
and UO_2036 (O_2036,N_49880,N_49926);
or UO_2037 (O_2037,N_49996,N_49963);
nor UO_2038 (O_2038,N_49781,N_49944);
nand UO_2039 (O_2039,N_49915,N_49960);
xnor UO_2040 (O_2040,N_49917,N_49921);
nand UO_2041 (O_2041,N_49845,N_49881);
and UO_2042 (O_2042,N_49801,N_49937);
nand UO_2043 (O_2043,N_49777,N_49936);
or UO_2044 (O_2044,N_49986,N_49998);
nand UO_2045 (O_2045,N_49805,N_49968);
xnor UO_2046 (O_2046,N_49752,N_49928);
or UO_2047 (O_2047,N_49888,N_49884);
nor UO_2048 (O_2048,N_49824,N_49969);
xor UO_2049 (O_2049,N_49998,N_49883);
and UO_2050 (O_2050,N_49751,N_49997);
nand UO_2051 (O_2051,N_49864,N_49886);
nand UO_2052 (O_2052,N_49878,N_49930);
xnor UO_2053 (O_2053,N_49799,N_49889);
nor UO_2054 (O_2054,N_49967,N_49905);
or UO_2055 (O_2055,N_49915,N_49861);
nor UO_2056 (O_2056,N_49989,N_49804);
xnor UO_2057 (O_2057,N_49979,N_49911);
nand UO_2058 (O_2058,N_49780,N_49868);
xnor UO_2059 (O_2059,N_49986,N_49946);
xor UO_2060 (O_2060,N_49940,N_49808);
nand UO_2061 (O_2061,N_49780,N_49839);
nor UO_2062 (O_2062,N_49911,N_49987);
nor UO_2063 (O_2063,N_49858,N_49893);
nand UO_2064 (O_2064,N_49906,N_49872);
xnor UO_2065 (O_2065,N_49943,N_49961);
nor UO_2066 (O_2066,N_49863,N_49911);
or UO_2067 (O_2067,N_49881,N_49894);
nor UO_2068 (O_2068,N_49917,N_49833);
nand UO_2069 (O_2069,N_49752,N_49770);
xnor UO_2070 (O_2070,N_49783,N_49946);
or UO_2071 (O_2071,N_49982,N_49967);
nand UO_2072 (O_2072,N_49807,N_49750);
nor UO_2073 (O_2073,N_49870,N_49887);
nand UO_2074 (O_2074,N_49788,N_49973);
and UO_2075 (O_2075,N_49961,N_49766);
nor UO_2076 (O_2076,N_49750,N_49855);
nand UO_2077 (O_2077,N_49775,N_49867);
and UO_2078 (O_2078,N_49874,N_49761);
xor UO_2079 (O_2079,N_49976,N_49775);
xnor UO_2080 (O_2080,N_49920,N_49855);
and UO_2081 (O_2081,N_49820,N_49851);
nor UO_2082 (O_2082,N_49915,N_49884);
nor UO_2083 (O_2083,N_49824,N_49867);
and UO_2084 (O_2084,N_49957,N_49958);
and UO_2085 (O_2085,N_49853,N_49784);
or UO_2086 (O_2086,N_49794,N_49836);
and UO_2087 (O_2087,N_49834,N_49830);
xnor UO_2088 (O_2088,N_49825,N_49967);
or UO_2089 (O_2089,N_49926,N_49945);
and UO_2090 (O_2090,N_49801,N_49976);
or UO_2091 (O_2091,N_49852,N_49958);
or UO_2092 (O_2092,N_49789,N_49827);
xor UO_2093 (O_2093,N_49804,N_49813);
xor UO_2094 (O_2094,N_49756,N_49864);
xnor UO_2095 (O_2095,N_49802,N_49893);
xor UO_2096 (O_2096,N_49790,N_49775);
nand UO_2097 (O_2097,N_49776,N_49770);
and UO_2098 (O_2098,N_49961,N_49763);
xor UO_2099 (O_2099,N_49887,N_49962);
and UO_2100 (O_2100,N_49941,N_49782);
or UO_2101 (O_2101,N_49778,N_49877);
and UO_2102 (O_2102,N_49910,N_49755);
nor UO_2103 (O_2103,N_49826,N_49912);
and UO_2104 (O_2104,N_49852,N_49844);
or UO_2105 (O_2105,N_49869,N_49916);
xor UO_2106 (O_2106,N_49920,N_49787);
nand UO_2107 (O_2107,N_49763,N_49939);
and UO_2108 (O_2108,N_49866,N_49794);
xnor UO_2109 (O_2109,N_49930,N_49993);
or UO_2110 (O_2110,N_49767,N_49877);
or UO_2111 (O_2111,N_49867,N_49860);
nand UO_2112 (O_2112,N_49895,N_49892);
nand UO_2113 (O_2113,N_49902,N_49752);
nor UO_2114 (O_2114,N_49862,N_49865);
nand UO_2115 (O_2115,N_49843,N_49784);
or UO_2116 (O_2116,N_49911,N_49994);
or UO_2117 (O_2117,N_49837,N_49965);
nand UO_2118 (O_2118,N_49833,N_49765);
or UO_2119 (O_2119,N_49904,N_49867);
nor UO_2120 (O_2120,N_49869,N_49889);
or UO_2121 (O_2121,N_49896,N_49801);
and UO_2122 (O_2122,N_49855,N_49817);
and UO_2123 (O_2123,N_49843,N_49980);
nor UO_2124 (O_2124,N_49836,N_49800);
xnor UO_2125 (O_2125,N_49782,N_49874);
nand UO_2126 (O_2126,N_49987,N_49977);
nand UO_2127 (O_2127,N_49812,N_49793);
xnor UO_2128 (O_2128,N_49947,N_49776);
nand UO_2129 (O_2129,N_49863,N_49919);
nor UO_2130 (O_2130,N_49763,N_49951);
xnor UO_2131 (O_2131,N_49880,N_49917);
nand UO_2132 (O_2132,N_49777,N_49932);
or UO_2133 (O_2133,N_49852,N_49783);
and UO_2134 (O_2134,N_49784,N_49916);
nand UO_2135 (O_2135,N_49957,N_49925);
or UO_2136 (O_2136,N_49882,N_49974);
xor UO_2137 (O_2137,N_49775,N_49992);
nor UO_2138 (O_2138,N_49790,N_49859);
nand UO_2139 (O_2139,N_49972,N_49950);
nor UO_2140 (O_2140,N_49951,N_49964);
xnor UO_2141 (O_2141,N_49982,N_49878);
and UO_2142 (O_2142,N_49854,N_49996);
nand UO_2143 (O_2143,N_49957,N_49885);
nand UO_2144 (O_2144,N_49790,N_49835);
and UO_2145 (O_2145,N_49994,N_49766);
nand UO_2146 (O_2146,N_49930,N_49890);
xnor UO_2147 (O_2147,N_49786,N_49756);
and UO_2148 (O_2148,N_49920,N_49949);
xnor UO_2149 (O_2149,N_49779,N_49778);
nor UO_2150 (O_2150,N_49994,N_49871);
nor UO_2151 (O_2151,N_49802,N_49938);
and UO_2152 (O_2152,N_49772,N_49933);
nor UO_2153 (O_2153,N_49924,N_49887);
and UO_2154 (O_2154,N_49885,N_49815);
xnor UO_2155 (O_2155,N_49956,N_49782);
and UO_2156 (O_2156,N_49877,N_49808);
and UO_2157 (O_2157,N_49754,N_49985);
or UO_2158 (O_2158,N_49871,N_49803);
nor UO_2159 (O_2159,N_49794,N_49966);
nor UO_2160 (O_2160,N_49947,N_49989);
or UO_2161 (O_2161,N_49990,N_49768);
nand UO_2162 (O_2162,N_49870,N_49759);
nor UO_2163 (O_2163,N_49922,N_49923);
and UO_2164 (O_2164,N_49899,N_49807);
nand UO_2165 (O_2165,N_49850,N_49984);
nor UO_2166 (O_2166,N_49929,N_49773);
xor UO_2167 (O_2167,N_49922,N_49858);
nor UO_2168 (O_2168,N_49777,N_49831);
xnor UO_2169 (O_2169,N_49938,N_49870);
xor UO_2170 (O_2170,N_49768,N_49782);
xnor UO_2171 (O_2171,N_49784,N_49973);
nand UO_2172 (O_2172,N_49871,N_49860);
or UO_2173 (O_2173,N_49901,N_49825);
and UO_2174 (O_2174,N_49784,N_49837);
nand UO_2175 (O_2175,N_49940,N_49914);
and UO_2176 (O_2176,N_49875,N_49860);
and UO_2177 (O_2177,N_49787,N_49864);
xnor UO_2178 (O_2178,N_49773,N_49835);
nand UO_2179 (O_2179,N_49982,N_49889);
nand UO_2180 (O_2180,N_49854,N_49884);
xnor UO_2181 (O_2181,N_49982,N_49998);
xnor UO_2182 (O_2182,N_49949,N_49867);
and UO_2183 (O_2183,N_49862,N_49879);
and UO_2184 (O_2184,N_49789,N_49793);
nor UO_2185 (O_2185,N_49898,N_49948);
nor UO_2186 (O_2186,N_49900,N_49967);
or UO_2187 (O_2187,N_49869,N_49813);
nor UO_2188 (O_2188,N_49843,N_49854);
nor UO_2189 (O_2189,N_49915,N_49990);
nand UO_2190 (O_2190,N_49967,N_49930);
and UO_2191 (O_2191,N_49947,N_49760);
or UO_2192 (O_2192,N_49820,N_49935);
or UO_2193 (O_2193,N_49880,N_49766);
nand UO_2194 (O_2194,N_49898,N_49887);
nand UO_2195 (O_2195,N_49863,N_49864);
and UO_2196 (O_2196,N_49842,N_49777);
or UO_2197 (O_2197,N_49804,N_49756);
xor UO_2198 (O_2198,N_49880,N_49888);
or UO_2199 (O_2199,N_49811,N_49799);
and UO_2200 (O_2200,N_49802,N_49795);
or UO_2201 (O_2201,N_49887,N_49826);
nand UO_2202 (O_2202,N_49771,N_49944);
xnor UO_2203 (O_2203,N_49889,N_49994);
nor UO_2204 (O_2204,N_49827,N_49989);
nor UO_2205 (O_2205,N_49972,N_49968);
nor UO_2206 (O_2206,N_49807,N_49866);
nor UO_2207 (O_2207,N_49764,N_49824);
nand UO_2208 (O_2208,N_49853,N_49944);
nand UO_2209 (O_2209,N_49888,N_49967);
xnor UO_2210 (O_2210,N_49762,N_49873);
nor UO_2211 (O_2211,N_49915,N_49761);
nor UO_2212 (O_2212,N_49842,N_49986);
nor UO_2213 (O_2213,N_49772,N_49875);
nand UO_2214 (O_2214,N_49893,N_49939);
and UO_2215 (O_2215,N_49825,N_49753);
and UO_2216 (O_2216,N_49997,N_49871);
and UO_2217 (O_2217,N_49924,N_49938);
nor UO_2218 (O_2218,N_49917,N_49876);
nor UO_2219 (O_2219,N_49799,N_49843);
and UO_2220 (O_2220,N_49785,N_49895);
nor UO_2221 (O_2221,N_49945,N_49856);
nand UO_2222 (O_2222,N_49769,N_49923);
or UO_2223 (O_2223,N_49878,N_49851);
xnor UO_2224 (O_2224,N_49965,N_49984);
nor UO_2225 (O_2225,N_49852,N_49884);
xor UO_2226 (O_2226,N_49937,N_49833);
nor UO_2227 (O_2227,N_49946,N_49857);
and UO_2228 (O_2228,N_49776,N_49930);
nand UO_2229 (O_2229,N_49981,N_49933);
xnor UO_2230 (O_2230,N_49865,N_49761);
or UO_2231 (O_2231,N_49784,N_49822);
or UO_2232 (O_2232,N_49914,N_49784);
and UO_2233 (O_2233,N_49846,N_49992);
nor UO_2234 (O_2234,N_49889,N_49838);
nor UO_2235 (O_2235,N_49769,N_49772);
xnor UO_2236 (O_2236,N_49930,N_49828);
nand UO_2237 (O_2237,N_49999,N_49899);
nor UO_2238 (O_2238,N_49796,N_49791);
nand UO_2239 (O_2239,N_49917,N_49959);
or UO_2240 (O_2240,N_49787,N_49800);
xnor UO_2241 (O_2241,N_49811,N_49987);
nor UO_2242 (O_2242,N_49919,N_49759);
xor UO_2243 (O_2243,N_49886,N_49932);
or UO_2244 (O_2244,N_49975,N_49947);
nand UO_2245 (O_2245,N_49766,N_49847);
nand UO_2246 (O_2246,N_49925,N_49761);
xnor UO_2247 (O_2247,N_49858,N_49785);
nor UO_2248 (O_2248,N_49838,N_49881);
xor UO_2249 (O_2249,N_49762,N_49864);
or UO_2250 (O_2250,N_49959,N_49876);
nand UO_2251 (O_2251,N_49838,N_49867);
and UO_2252 (O_2252,N_49976,N_49756);
xor UO_2253 (O_2253,N_49783,N_49955);
or UO_2254 (O_2254,N_49827,N_49850);
xnor UO_2255 (O_2255,N_49842,N_49844);
and UO_2256 (O_2256,N_49861,N_49843);
and UO_2257 (O_2257,N_49888,N_49905);
xor UO_2258 (O_2258,N_49764,N_49894);
xnor UO_2259 (O_2259,N_49990,N_49804);
or UO_2260 (O_2260,N_49800,N_49768);
nor UO_2261 (O_2261,N_49844,N_49813);
and UO_2262 (O_2262,N_49841,N_49807);
or UO_2263 (O_2263,N_49888,N_49826);
xor UO_2264 (O_2264,N_49995,N_49964);
xor UO_2265 (O_2265,N_49882,N_49807);
or UO_2266 (O_2266,N_49855,N_49963);
xor UO_2267 (O_2267,N_49952,N_49928);
nor UO_2268 (O_2268,N_49758,N_49970);
nor UO_2269 (O_2269,N_49759,N_49875);
or UO_2270 (O_2270,N_49896,N_49843);
nor UO_2271 (O_2271,N_49856,N_49928);
and UO_2272 (O_2272,N_49806,N_49824);
and UO_2273 (O_2273,N_49847,N_49955);
xnor UO_2274 (O_2274,N_49919,N_49781);
and UO_2275 (O_2275,N_49977,N_49761);
nand UO_2276 (O_2276,N_49767,N_49766);
and UO_2277 (O_2277,N_49867,N_49753);
or UO_2278 (O_2278,N_49795,N_49897);
nand UO_2279 (O_2279,N_49840,N_49981);
nor UO_2280 (O_2280,N_49820,N_49809);
or UO_2281 (O_2281,N_49874,N_49888);
nor UO_2282 (O_2282,N_49820,N_49875);
or UO_2283 (O_2283,N_49947,N_49972);
nor UO_2284 (O_2284,N_49980,N_49842);
xor UO_2285 (O_2285,N_49849,N_49893);
and UO_2286 (O_2286,N_49867,N_49780);
or UO_2287 (O_2287,N_49913,N_49771);
and UO_2288 (O_2288,N_49992,N_49795);
nand UO_2289 (O_2289,N_49861,N_49974);
nand UO_2290 (O_2290,N_49821,N_49767);
nand UO_2291 (O_2291,N_49851,N_49788);
xor UO_2292 (O_2292,N_49964,N_49838);
and UO_2293 (O_2293,N_49988,N_49781);
nor UO_2294 (O_2294,N_49796,N_49991);
or UO_2295 (O_2295,N_49905,N_49991);
xor UO_2296 (O_2296,N_49769,N_49823);
and UO_2297 (O_2297,N_49826,N_49852);
nor UO_2298 (O_2298,N_49867,N_49807);
or UO_2299 (O_2299,N_49933,N_49934);
nor UO_2300 (O_2300,N_49963,N_49873);
xnor UO_2301 (O_2301,N_49910,N_49771);
or UO_2302 (O_2302,N_49915,N_49922);
and UO_2303 (O_2303,N_49959,N_49844);
and UO_2304 (O_2304,N_49775,N_49865);
or UO_2305 (O_2305,N_49921,N_49768);
xor UO_2306 (O_2306,N_49915,N_49940);
nor UO_2307 (O_2307,N_49941,N_49951);
nand UO_2308 (O_2308,N_49796,N_49854);
xnor UO_2309 (O_2309,N_49816,N_49906);
and UO_2310 (O_2310,N_49948,N_49991);
xnor UO_2311 (O_2311,N_49916,N_49828);
or UO_2312 (O_2312,N_49758,N_49956);
nor UO_2313 (O_2313,N_49759,N_49942);
xnor UO_2314 (O_2314,N_49850,N_49847);
or UO_2315 (O_2315,N_49766,N_49953);
xnor UO_2316 (O_2316,N_49799,N_49879);
nand UO_2317 (O_2317,N_49831,N_49770);
nor UO_2318 (O_2318,N_49956,N_49904);
or UO_2319 (O_2319,N_49892,N_49789);
nand UO_2320 (O_2320,N_49842,N_49916);
nand UO_2321 (O_2321,N_49823,N_49874);
xnor UO_2322 (O_2322,N_49825,N_49763);
nor UO_2323 (O_2323,N_49840,N_49961);
xnor UO_2324 (O_2324,N_49912,N_49913);
xor UO_2325 (O_2325,N_49815,N_49752);
and UO_2326 (O_2326,N_49763,N_49758);
or UO_2327 (O_2327,N_49883,N_49957);
and UO_2328 (O_2328,N_49818,N_49915);
nand UO_2329 (O_2329,N_49933,N_49765);
or UO_2330 (O_2330,N_49775,N_49839);
nor UO_2331 (O_2331,N_49960,N_49804);
or UO_2332 (O_2332,N_49955,N_49947);
xnor UO_2333 (O_2333,N_49923,N_49986);
xor UO_2334 (O_2334,N_49755,N_49898);
nand UO_2335 (O_2335,N_49870,N_49866);
xnor UO_2336 (O_2336,N_49900,N_49800);
xnor UO_2337 (O_2337,N_49763,N_49999);
nand UO_2338 (O_2338,N_49839,N_49767);
or UO_2339 (O_2339,N_49903,N_49900);
nor UO_2340 (O_2340,N_49846,N_49906);
or UO_2341 (O_2341,N_49874,N_49880);
nor UO_2342 (O_2342,N_49888,N_49970);
and UO_2343 (O_2343,N_49763,N_49901);
xnor UO_2344 (O_2344,N_49831,N_49785);
nor UO_2345 (O_2345,N_49983,N_49812);
xnor UO_2346 (O_2346,N_49798,N_49843);
or UO_2347 (O_2347,N_49981,N_49990);
and UO_2348 (O_2348,N_49828,N_49920);
and UO_2349 (O_2349,N_49779,N_49970);
and UO_2350 (O_2350,N_49805,N_49763);
or UO_2351 (O_2351,N_49963,N_49971);
or UO_2352 (O_2352,N_49965,N_49964);
or UO_2353 (O_2353,N_49899,N_49781);
xor UO_2354 (O_2354,N_49816,N_49773);
nand UO_2355 (O_2355,N_49898,N_49953);
nand UO_2356 (O_2356,N_49815,N_49845);
nor UO_2357 (O_2357,N_49799,N_49917);
nand UO_2358 (O_2358,N_49765,N_49979);
xor UO_2359 (O_2359,N_49902,N_49826);
nor UO_2360 (O_2360,N_49929,N_49756);
xnor UO_2361 (O_2361,N_49825,N_49883);
nor UO_2362 (O_2362,N_49773,N_49777);
xnor UO_2363 (O_2363,N_49945,N_49875);
and UO_2364 (O_2364,N_49988,N_49763);
and UO_2365 (O_2365,N_49796,N_49968);
nand UO_2366 (O_2366,N_49957,N_49790);
xnor UO_2367 (O_2367,N_49835,N_49823);
xor UO_2368 (O_2368,N_49833,N_49814);
and UO_2369 (O_2369,N_49808,N_49845);
nor UO_2370 (O_2370,N_49763,N_49819);
xnor UO_2371 (O_2371,N_49855,N_49968);
xnor UO_2372 (O_2372,N_49826,N_49755);
xor UO_2373 (O_2373,N_49794,N_49834);
nand UO_2374 (O_2374,N_49786,N_49810);
and UO_2375 (O_2375,N_49802,N_49895);
and UO_2376 (O_2376,N_49998,N_49784);
xor UO_2377 (O_2377,N_49873,N_49817);
xor UO_2378 (O_2378,N_49888,N_49780);
nand UO_2379 (O_2379,N_49933,N_49844);
nor UO_2380 (O_2380,N_49879,N_49796);
or UO_2381 (O_2381,N_49939,N_49957);
and UO_2382 (O_2382,N_49945,N_49848);
and UO_2383 (O_2383,N_49815,N_49861);
xor UO_2384 (O_2384,N_49942,N_49783);
nand UO_2385 (O_2385,N_49936,N_49946);
and UO_2386 (O_2386,N_49888,N_49921);
or UO_2387 (O_2387,N_49888,N_49848);
or UO_2388 (O_2388,N_49973,N_49958);
nor UO_2389 (O_2389,N_49762,N_49838);
or UO_2390 (O_2390,N_49923,N_49980);
nand UO_2391 (O_2391,N_49965,N_49940);
or UO_2392 (O_2392,N_49831,N_49920);
xnor UO_2393 (O_2393,N_49805,N_49886);
xor UO_2394 (O_2394,N_49984,N_49986);
nand UO_2395 (O_2395,N_49784,N_49791);
nor UO_2396 (O_2396,N_49883,N_49856);
xor UO_2397 (O_2397,N_49806,N_49772);
or UO_2398 (O_2398,N_49859,N_49977);
nand UO_2399 (O_2399,N_49848,N_49756);
or UO_2400 (O_2400,N_49899,N_49966);
nand UO_2401 (O_2401,N_49855,N_49896);
xnor UO_2402 (O_2402,N_49777,N_49783);
xor UO_2403 (O_2403,N_49854,N_49921);
xor UO_2404 (O_2404,N_49845,N_49763);
and UO_2405 (O_2405,N_49845,N_49816);
nor UO_2406 (O_2406,N_49858,N_49899);
nand UO_2407 (O_2407,N_49776,N_49924);
nor UO_2408 (O_2408,N_49883,N_49880);
nand UO_2409 (O_2409,N_49812,N_49785);
nand UO_2410 (O_2410,N_49803,N_49928);
nand UO_2411 (O_2411,N_49818,N_49754);
or UO_2412 (O_2412,N_49922,N_49817);
nor UO_2413 (O_2413,N_49942,N_49760);
and UO_2414 (O_2414,N_49816,N_49800);
xor UO_2415 (O_2415,N_49984,N_49870);
nand UO_2416 (O_2416,N_49798,N_49982);
nor UO_2417 (O_2417,N_49848,N_49845);
xor UO_2418 (O_2418,N_49808,N_49936);
nand UO_2419 (O_2419,N_49818,N_49925);
nor UO_2420 (O_2420,N_49985,N_49956);
and UO_2421 (O_2421,N_49962,N_49796);
and UO_2422 (O_2422,N_49798,N_49801);
and UO_2423 (O_2423,N_49764,N_49880);
xor UO_2424 (O_2424,N_49973,N_49830);
and UO_2425 (O_2425,N_49971,N_49863);
nor UO_2426 (O_2426,N_49841,N_49961);
or UO_2427 (O_2427,N_49750,N_49879);
nor UO_2428 (O_2428,N_49750,N_49837);
and UO_2429 (O_2429,N_49951,N_49836);
nor UO_2430 (O_2430,N_49766,N_49882);
xor UO_2431 (O_2431,N_49796,N_49939);
and UO_2432 (O_2432,N_49997,N_49805);
xnor UO_2433 (O_2433,N_49876,N_49782);
nand UO_2434 (O_2434,N_49801,N_49964);
and UO_2435 (O_2435,N_49965,N_49769);
xnor UO_2436 (O_2436,N_49882,N_49857);
and UO_2437 (O_2437,N_49991,N_49929);
xor UO_2438 (O_2438,N_49800,N_49912);
xor UO_2439 (O_2439,N_49847,N_49986);
and UO_2440 (O_2440,N_49808,N_49872);
or UO_2441 (O_2441,N_49952,N_49781);
nor UO_2442 (O_2442,N_49977,N_49919);
nand UO_2443 (O_2443,N_49848,N_49810);
nand UO_2444 (O_2444,N_49756,N_49894);
nand UO_2445 (O_2445,N_49857,N_49987);
xor UO_2446 (O_2446,N_49867,N_49792);
and UO_2447 (O_2447,N_49865,N_49958);
nand UO_2448 (O_2448,N_49867,N_49787);
xnor UO_2449 (O_2449,N_49981,N_49753);
nor UO_2450 (O_2450,N_49908,N_49781);
xor UO_2451 (O_2451,N_49850,N_49756);
or UO_2452 (O_2452,N_49849,N_49991);
xor UO_2453 (O_2453,N_49858,N_49876);
or UO_2454 (O_2454,N_49954,N_49982);
nand UO_2455 (O_2455,N_49946,N_49801);
or UO_2456 (O_2456,N_49873,N_49921);
and UO_2457 (O_2457,N_49927,N_49768);
or UO_2458 (O_2458,N_49783,N_49957);
nor UO_2459 (O_2459,N_49977,N_49753);
nor UO_2460 (O_2460,N_49803,N_49769);
xnor UO_2461 (O_2461,N_49797,N_49809);
nand UO_2462 (O_2462,N_49987,N_49873);
and UO_2463 (O_2463,N_49881,N_49785);
or UO_2464 (O_2464,N_49793,N_49918);
nand UO_2465 (O_2465,N_49988,N_49907);
nor UO_2466 (O_2466,N_49885,N_49819);
xor UO_2467 (O_2467,N_49984,N_49932);
and UO_2468 (O_2468,N_49978,N_49911);
nor UO_2469 (O_2469,N_49800,N_49779);
or UO_2470 (O_2470,N_49851,N_49998);
nand UO_2471 (O_2471,N_49764,N_49965);
nor UO_2472 (O_2472,N_49999,N_49886);
nor UO_2473 (O_2473,N_49948,N_49779);
and UO_2474 (O_2474,N_49940,N_49873);
nand UO_2475 (O_2475,N_49771,N_49888);
and UO_2476 (O_2476,N_49901,N_49919);
xnor UO_2477 (O_2477,N_49846,N_49827);
xor UO_2478 (O_2478,N_49984,N_49864);
nand UO_2479 (O_2479,N_49841,N_49789);
nand UO_2480 (O_2480,N_49857,N_49816);
nor UO_2481 (O_2481,N_49878,N_49765);
xnor UO_2482 (O_2482,N_49945,N_49781);
xnor UO_2483 (O_2483,N_49773,N_49812);
xnor UO_2484 (O_2484,N_49850,N_49883);
nor UO_2485 (O_2485,N_49984,N_49996);
nor UO_2486 (O_2486,N_49794,N_49774);
xnor UO_2487 (O_2487,N_49983,N_49889);
xor UO_2488 (O_2488,N_49912,N_49812);
xnor UO_2489 (O_2489,N_49753,N_49843);
nor UO_2490 (O_2490,N_49756,N_49818);
or UO_2491 (O_2491,N_49817,N_49854);
and UO_2492 (O_2492,N_49969,N_49905);
and UO_2493 (O_2493,N_49809,N_49831);
nor UO_2494 (O_2494,N_49989,N_49920);
xnor UO_2495 (O_2495,N_49913,N_49894);
and UO_2496 (O_2496,N_49756,N_49869);
nor UO_2497 (O_2497,N_49988,N_49909);
or UO_2498 (O_2498,N_49871,N_49985);
xor UO_2499 (O_2499,N_49906,N_49765);
or UO_2500 (O_2500,N_49862,N_49752);
or UO_2501 (O_2501,N_49959,N_49910);
nand UO_2502 (O_2502,N_49845,N_49793);
nor UO_2503 (O_2503,N_49969,N_49915);
nand UO_2504 (O_2504,N_49801,N_49814);
and UO_2505 (O_2505,N_49859,N_49978);
and UO_2506 (O_2506,N_49920,N_49764);
and UO_2507 (O_2507,N_49799,N_49884);
and UO_2508 (O_2508,N_49963,N_49952);
or UO_2509 (O_2509,N_49907,N_49773);
nor UO_2510 (O_2510,N_49751,N_49872);
xnor UO_2511 (O_2511,N_49883,N_49886);
nor UO_2512 (O_2512,N_49982,N_49931);
nand UO_2513 (O_2513,N_49972,N_49835);
nand UO_2514 (O_2514,N_49831,N_49899);
nor UO_2515 (O_2515,N_49974,N_49836);
nand UO_2516 (O_2516,N_49831,N_49966);
or UO_2517 (O_2517,N_49962,N_49754);
or UO_2518 (O_2518,N_49901,N_49971);
or UO_2519 (O_2519,N_49878,N_49793);
and UO_2520 (O_2520,N_49839,N_49853);
nor UO_2521 (O_2521,N_49985,N_49785);
nand UO_2522 (O_2522,N_49938,N_49797);
xnor UO_2523 (O_2523,N_49973,N_49761);
or UO_2524 (O_2524,N_49753,N_49802);
xnor UO_2525 (O_2525,N_49793,N_49864);
or UO_2526 (O_2526,N_49836,N_49807);
nor UO_2527 (O_2527,N_49760,N_49831);
nor UO_2528 (O_2528,N_49886,N_49892);
nor UO_2529 (O_2529,N_49945,N_49770);
and UO_2530 (O_2530,N_49917,N_49772);
xor UO_2531 (O_2531,N_49869,N_49753);
or UO_2532 (O_2532,N_49911,N_49877);
nand UO_2533 (O_2533,N_49771,N_49886);
nor UO_2534 (O_2534,N_49872,N_49816);
or UO_2535 (O_2535,N_49943,N_49863);
nor UO_2536 (O_2536,N_49886,N_49977);
and UO_2537 (O_2537,N_49829,N_49905);
and UO_2538 (O_2538,N_49976,N_49841);
or UO_2539 (O_2539,N_49863,N_49976);
or UO_2540 (O_2540,N_49978,N_49928);
or UO_2541 (O_2541,N_49935,N_49878);
or UO_2542 (O_2542,N_49925,N_49931);
nor UO_2543 (O_2543,N_49844,N_49950);
nor UO_2544 (O_2544,N_49780,N_49805);
nor UO_2545 (O_2545,N_49768,N_49775);
or UO_2546 (O_2546,N_49940,N_49777);
nand UO_2547 (O_2547,N_49990,N_49910);
xor UO_2548 (O_2548,N_49887,N_49986);
nor UO_2549 (O_2549,N_49786,N_49906);
or UO_2550 (O_2550,N_49751,N_49884);
or UO_2551 (O_2551,N_49892,N_49837);
nand UO_2552 (O_2552,N_49941,N_49766);
nor UO_2553 (O_2553,N_49751,N_49912);
nor UO_2554 (O_2554,N_49938,N_49853);
and UO_2555 (O_2555,N_49872,N_49856);
or UO_2556 (O_2556,N_49837,N_49755);
xnor UO_2557 (O_2557,N_49800,N_49850);
nor UO_2558 (O_2558,N_49838,N_49857);
and UO_2559 (O_2559,N_49918,N_49780);
or UO_2560 (O_2560,N_49756,N_49880);
xor UO_2561 (O_2561,N_49938,N_49987);
nor UO_2562 (O_2562,N_49992,N_49890);
or UO_2563 (O_2563,N_49963,N_49995);
or UO_2564 (O_2564,N_49829,N_49909);
xor UO_2565 (O_2565,N_49866,N_49785);
nor UO_2566 (O_2566,N_49990,N_49928);
xnor UO_2567 (O_2567,N_49761,N_49776);
and UO_2568 (O_2568,N_49847,N_49829);
and UO_2569 (O_2569,N_49999,N_49961);
and UO_2570 (O_2570,N_49866,N_49956);
xor UO_2571 (O_2571,N_49937,N_49996);
nor UO_2572 (O_2572,N_49798,N_49914);
xor UO_2573 (O_2573,N_49814,N_49955);
nor UO_2574 (O_2574,N_49990,N_49968);
or UO_2575 (O_2575,N_49998,N_49844);
nand UO_2576 (O_2576,N_49750,N_49988);
or UO_2577 (O_2577,N_49802,N_49856);
or UO_2578 (O_2578,N_49789,N_49905);
nor UO_2579 (O_2579,N_49889,N_49978);
or UO_2580 (O_2580,N_49999,N_49853);
and UO_2581 (O_2581,N_49884,N_49792);
and UO_2582 (O_2582,N_49756,N_49801);
nor UO_2583 (O_2583,N_49929,N_49937);
or UO_2584 (O_2584,N_49778,N_49861);
or UO_2585 (O_2585,N_49881,N_49769);
xor UO_2586 (O_2586,N_49800,N_49750);
xnor UO_2587 (O_2587,N_49752,N_49852);
xor UO_2588 (O_2588,N_49793,N_49805);
xor UO_2589 (O_2589,N_49812,N_49870);
nand UO_2590 (O_2590,N_49885,N_49877);
nor UO_2591 (O_2591,N_49751,N_49848);
xnor UO_2592 (O_2592,N_49975,N_49879);
nand UO_2593 (O_2593,N_49758,N_49950);
or UO_2594 (O_2594,N_49998,N_49759);
nand UO_2595 (O_2595,N_49847,N_49979);
or UO_2596 (O_2596,N_49799,N_49797);
nor UO_2597 (O_2597,N_49802,N_49852);
nand UO_2598 (O_2598,N_49753,N_49792);
or UO_2599 (O_2599,N_49866,N_49821);
and UO_2600 (O_2600,N_49750,N_49937);
or UO_2601 (O_2601,N_49949,N_49813);
nor UO_2602 (O_2602,N_49863,N_49784);
and UO_2603 (O_2603,N_49997,N_49825);
nor UO_2604 (O_2604,N_49981,N_49950);
or UO_2605 (O_2605,N_49772,N_49764);
or UO_2606 (O_2606,N_49868,N_49943);
nand UO_2607 (O_2607,N_49870,N_49979);
or UO_2608 (O_2608,N_49954,N_49855);
and UO_2609 (O_2609,N_49809,N_49775);
xnor UO_2610 (O_2610,N_49801,N_49847);
or UO_2611 (O_2611,N_49826,N_49796);
and UO_2612 (O_2612,N_49844,N_49835);
nor UO_2613 (O_2613,N_49955,N_49976);
nor UO_2614 (O_2614,N_49944,N_49973);
or UO_2615 (O_2615,N_49987,N_49886);
and UO_2616 (O_2616,N_49866,N_49798);
xnor UO_2617 (O_2617,N_49963,N_49919);
and UO_2618 (O_2618,N_49906,N_49868);
and UO_2619 (O_2619,N_49932,N_49861);
nor UO_2620 (O_2620,N_49760,N_49998);
or UO_2621 (O_2621,N_49833,N_49838);
nor UO_2622 (O_2622,N_49853,N_49876);
nor UO_2623 (O_2623,N_49911,N_49970);
nor UO_2624 (O_2624,N_49970,N_49799);
and UO_2625 (O_2625,N_49803,N_49917);
or UO_2626 (O_2626,N_49893,N_49954);
or UO_2627 (O_2627,N_49921,N_49892);
and UO_2628 (O_2628,N_49843,N_49981);
nand UO_2629 (O_2629,N_49772,N_49784);
nor UO_2630 (O_2630,N_49917,N_49973);
or UO_2631 (O_2631,N_49826,N_49799);
and UO_2632 (O_2632,N_49881,N_49996);
or UO_2633 (O_2633,N_49873,N_49751);
nand UO_2634 (O_2634,N_49865,N_49791);
nand UO_2635 (O_2635,N_49777,N_49891);
xnor UO_2636 (O_2636,N_49851,N_49862);
xor UO_2637 (O_2637,N_49784,N_49924);
nand UO_2638 (O_2638,N_49824,N_49799);
xor UO_2639 (O_2639,N_49789,N_49988);
xor UO_2640 (O_2640,N_49832,N_49768);
or UO_2641 (O_2641,N_49770,N_49887);
xnor UO_2642 (O_2642,N_49994,N_49845);
or UO_2643 (O_2643,N_49763,N_49889);
xnor UO_2644 (O_2644,N_49796,N_49907);
or UO_2645 (O_2645,N_49941,N_49841);
xnor UO_2646 (O_2646,N_49785,N_49995);
and UO_2647 (O_2647,N_49802,N_49942);
nor UO_2648 (O_2648,N_49934,N_49828);
nand UO_2649 (O_2649,N_49757,N_49880);
xnor UO_2650 (O_2650,N_49918,N_49802);
nand UO_2651 (O_2651,N_49768,N_49843);
and UO_2652 (O_2652,N_49914,N_49897);
and UO_2653 (O_2653,N_49833,N_49835);
xnor UO_2654 (O_2654,N_49908,N_49900);
nor UO_2655 (O_2655,N_49859,N_49776);
or UO_2656 (O_2656,N_49844,N_49869);
and UO_2657 (O_2657,N_49991,N_49839);
nand UO_2658 (O_2658,N_49754,N_49886);
and UO_2659 (O_2659,N_49944,N_49994);
nor UO_2660 (O_2660,N_49914,N_49915);
nand UO_2661 (O_2661,N_49876,N_49804);
nor UO_2662 (O_2662,N_49872,N_49920);
and UO_2663 (O_2663,N_49961,N_49949);
nor UO_2664 (O_2664,N_49847,N_49957);
or UO_2665 (O_2665,N_49820,N_49772);
nor UO_2666 (O_2666,N_49780,N_49849);
xnor UO_2667 (O_2667,N_49940,N_49804);
nor UO_2668 (O_2668,N_49981,N_49851);
nand UO_2669 (O_2669,N_49842,N_49941);
xnor UO_2670 (O_2670,N_49806,N_49942);
or UO_2671 (O_2671,N_49929,N_49909);
xnor UO_2672 (O_2672,N_49897,N_49790);
and UO_2673 (O_2673,N_49878,N_49757);
nor UO_2674 (O_2674,N_49805,N_49904);
nor UO_2675 (O_2675,N_49803,N_49765);
or UO_2676 (O_2676,N_49827,N_49822);
or UO_2677 (O_2677,N_49983,N_49956);
nand UO_2678 (O_2678,N_49942,N_49853);
nor UO_2679 (O_2679,N_49812,N_49988);
xnor UO_2680 (O_2680,N_49925,N_49829);
xnor UO_2681 (O_2681,N_49764,N_49907);
or UO_2682 (O_2682,N_49905,N_49975);
nand UO_2683 (O_2683,N_49877,N_49918);
or UO_2684 (O_2684,N_49964,N_49775);
and UO_2685 (O_2685,N_49872,N_49801);
nand UO_2686 (O_2686,N_49826,N_49899);
and UO_2687 (O_2687,N_49956,N_49823);
and UO_2688 (O_2688,N_49949,N_49805);
xor UO_2689 (O_2689,N_49931,N_49934);
or UO_2690 (O_2690,N_49947,N_49970);
and UO_2691 (O_2691,N_49977,N_49820);
nand UO_2692 (O_2692,N_49966,N_49754);
or UO_2693 (O_2693,N_49765,N_49889);
xor UO_2694 (O_2694,N_49818,N_49956);
xnor UO_2695 (O_2695,N_49817,N_49843);
nor UO_2696 (O_2696,N_49931,N_49788);
or UO_2697 (O_2697,N_49815,N_49853);
nor UO_2698 (O_2698,N_49994,N_49760);
xor UO_2699 (O_2699,N_49933,N_49867);
and UO_2700 (O_2700,N_49789,N_49878);
nand UO_2701 (O_2701,N_49975,N_49945);
or UO_2702 (O_2702,N_49944,N_49809);
xor UO_2703 (O_2703,N_49895,N_49976);
or UO_2704 (O_2704,N_49907,N_49763);
and UO_2705 (O_2705,N_49772,N_49765);
nand UO_2706 (O_2706,N_49979,N_49853);
or UO_2707 (O_2707,N_49828,N_49820);
nand UO_2708 (O_2708,N_49953,N_49816);
or UO_2709 (O_2709,N_49822,N_49906);
and UO_2710 (O_2710,N_49782,N_49895);
xor UO_2711 (O_2711,N_49775,N_49994);
nand UO_2712 (O_2712,N_49759,N_49766);
and UO_2713 (O_2713,N_49999,N_49865);
xor UO_2714 (O_2714,N_49796,N_49911);
xor UO_2715 (O_2715,N_49813,N_49798);
or UO_2716 (O_2716,N_49977,N_49975);
nand UO_2717 (O_2717,N_49949,N_49850);
and UO_2718 (O_2718,N_49932,N_49926);
nor UO_2719 (O_2719,N_49794,N_49759);
and UO_2720 (O_2720,N_49993,N_49753);
nand UO_2721 (O_2721,N_49797,N_49969);
nor UO_2722 (O_2722,N_49943,N_49824);
xnor UO_2723 (O_2723,N_49791,N_49959);
and UO_2724 (O_2724,N_49770,N_49930);
and UO_2725 (O_2725,N_49876,N_49982);
nor UO_2726 (O_2726,N_49872,N_49829);
nand UO_2727 (O_2727,N_49818,N_49779);
nor UO_2728 (O_2728,N_49865,N_49931);
or UO_2729 (O_2729,N_49974,N_49790);
nand UO_2730 (O_2730,N_49804,N_49885);
xnor UO_2731 (O_2731,N_49852,N_49876);
or UO_2732 (O_2732,N_49890,N_49844);
or UO_2733 (O_2733,N_49787,N_49868);
or UO_2734 (O_2734,N_49888,N_49761);
and UO_2735 (O_2735,N_49812,N_49858);
and UO_2736 (O_2736,N_49914,N_49895);
nand UO_2737 (O_2737,N_49952,N_49880);
nand UO_2738 (O_2738,N_49889,N_49970);
xor UO_2739 (O_2739,N_49795,N_49832);
nand UO_2740 (O_2740,N_49899,N_49837);
nand UO_2741 (O_2741,N_49903,N_49799);
or UO_2742 (O_2742,N_49770,N_49985);
and UO_2743 (O_2743,N_49953,N_49825);
xor UO_2744 (O_2744,N_49801,N_49810);
xor UO_2745 (O_2745,N_49849,N_49863);
or UO_2746 (O_2746,N_49887,N_49931);
xor UO_2747 (O_2747,N_49828,N_49860);
or UO_2748 (O_2748,N_49977,N_49914);
or UO_2749 (O_2749,N_49856,N_49790);
nor UO_2750 (O_2750,N_49770,N_49993);
nand UO_2751 (O_2751,N_49922,N_49881);
nor UO_2752 (O_2752,N_49874,N_49990);
and UO_2753 (O_2753,N_49933,N_49957);
xor UO_2754 (O_2754,N_49882,N_49928);
or UO_2755 (O_2755,N_49803,N_49966);
nand UO_2756 (O_2756,N_49962,N_49921);
nand UO_2757 (O_2757,N_49990,N_49793);
nor UO_2758 (O_2758,N_49964,N_49878);
nand UO_2759 (O_2759,N_49808,N_49895);
xnor UO_2760 (O_2760,N_49992,N_49924);
nor UO_2761 (O_2761,N_49867,N_49768);
nand UO_2762 (O_2762,N_49816,N_49764);
and UO_2763 (O_2763,N_49881,N_49951);
xor UO_2764 (O_2764,N_49934,N_49962);
or UO_2765 (O_2765,N_49861,N_49826);
or UO_2766 (O_2766,N_49820,N_49768);
nand UO_2767 (O_2767,N_49999,N_49818);
nor UO_2768 (O_2768,N_49942,N_49903);
and UO_2769 (O_2769,N_49969,N_49877);
nor UO_2770 (O_2770,N_49919,N_49947);
and UO_2771 (O_2771,N_49842,N_49945);
nor UO_2772 (O_2772,N_49927,N_49988);
xor UO_2773 (O_2773,N_49946,N_49899);
nor UO_2774 (O_2774,N_49793,N_49924);
xor UO_2775 (O_2775,N_49967,N_49978);
nor UO_2776 (O_2776,N_49979,N_49763);
or UO_2777 (O_2777,N_49883,N_49903);
and UO_2778 (O_2778,N_49952,N_49994);
and UO_2779 (O_2779,N_49844,N_49785);
nand UO_2780 (O_2780,N_49896,N_49751);
nor UO_2781 (O_2781,N_49752,N_49929);
nand UO_2782 (O_2782,N_49834,N_49971);
and UO_2783 (O_2783,N_49883,N_49940);
xnor UO_2784 (O_2784,N_49789,N_49866);
nor UO_2785 (O_2785,N_49763,N_49846);
nand UO_2786 (O_2786,N_49910,N_49781);
or UO_2787 (O_2787,N_49866,N_49791);
nor UO_2788 (O_2788,N_49752,N_49799);
nand UO_2789 (O_2789,N_49759,N_49877);
nand UO_2790 (O_2790,N_49904,N_49996);
nand UO_2791 (O_2791,N_49815,N_49778);
nand UO_2792 (O_2792,N_49879,N_49806);
and UO_2793 (O_2793,N_49918,N_49924);
nor UO_2794 (O_2794,N_49952,N_49816);
xnor UO_2795 (O_2795,N_49984,N_49921);
nor UO_2796 (O_2796,N_49919,N_49867);
or UO_2797 (O_2797,N_49956,N_49789);
and UO_2798 (O_2798,N_49941,N_49769);
nor UO_2799 (O_2799,N_49924,N_49815);
and UO_2800 (O_2800,N_49979,N_49950);
nand UO_2801 (O_2801,N_49985,N_49929);
nand UO_2802 (O_2802,N_49986,N_49814);
or UO_2803 (O_2803,N_49886,N_49871);
and UO_2804 (O_2804,N_49931,N_49935);
nand UO_2805 (O_2805,N_49752,N_49953);
nand UO_2806 (O_2806,N_49794,N_49753);
xnor UO_2807 (O_2807,N_49871,N_49953);
nand UO_2808 (O_2808,N_49898,N_49799);
nor UO_2809 (O_2809,N_49766,N_49775);
nand UO_2810 (O_2810,N_49868,N_49966);
nor UO_2811 (O_2811,N_49864,N_49930);
and UO_2812 (O_2812,N_49880,N_49844);
xor UO_2813 (O_2813,N_49925,N_49776);
nor UO_2814 (O_2814,N_49965,N_49943);
or UO_2815 (O_2815,N_49836,N_49851);
nor UO_2816 (O_2816,N_49840,N_49913);
and UO_2817 (O_2817,N_49788,N_49822);
nand UO_2818 (O_2818,N_49977,N_49965);
xor UO_2819 (O_2819,N_49811,N_49763);
nand UO_2820 (O_2820,N_49894,N_49809);
or UO_2821 (O_2821,N_49954,N_49823);
or UO_2822 (O_2822,N_49903,N_49978);
xnor UO_2823 (O_2823,N_49936,N_49805);
nand UO_2824 (O_2824,N_49871,N_49808);
xor UO_2825 (O_2825,N_49853,N_49783);
and UO_2826 (O_2826,N_49825,N_49800);
or UO_2827 (O_2827,N_49914,N_49751);
nand UO_2828 (O_2828,N_49858,N_49897);
and UO_2829 (O_2829,N_49936,N_49828);
nor UO_2830 (O_2830,N_49901,N_49986);
xor UO_2831 (O_2831,N_49891,N_49765);
xnor UO_2832 (O_2832,N_49825,N_49807);
xnor UO_2833 (O_2833,N_49829,N_49976);
nand UO_2834 (O_2834,N_49777,N_49923);
and UO_2835 (O_2835,N_49960,N_49989);
or UO_2836 (O_2836,N_49958,N_49756);
nor UO_2837 (O_2837,N_49950,N_49879);
and UO_2838 (O_2838,N_49851,N_49868);
or UO_2839 (O_2839,N_49821,N_49779);
nor UO_2840 (O_2840,N_49858,N_49939);
nor UO_2841 (O_2841,N_49929,N_49998);
or UO_2842 (O_2842,N_49975,N_49791);
nor UO_2843 (O_2843,N_49869,N_49828);
and UO_2844 (O_2844,N_49964,N_49799);
nor UO_2845 (O_2845,N_49760,N_49849);
and UO_2846 (O_2846,N_49755,N_49872);
or UO_2847 (O_2847,N_49886,N_49807);
and UO_2848 (O_2848,N_49946,N_49988);
nor UO_2849 (O_2849,N_49957,N_49807);
nor UO_2850 (O_2850,N_49891,N_49826);
nand UO_2851 (O_2851,N_49868,N_49961);
or UO_2852 (O_2852,N_49821,N_49910);
nand UO_2853 (O_2853,N_49997,N_49838);
and UO_2854 (O_2854,N_49819,N_49931);
or UO_2855 (O_2855,N_49978,N_49879);
nor UO_2856 (O_2856,N_49901,N_49830);
nand UO_2857 (O_2857,N_49816,N_49975);
nor UO_2858 (O_2858,N_49911,N_49757);
or UO_2859 (O_2859,N_49911,N_49988);
and UO_2860 (O_2860,N_49961,N_49906);
nand UO_2861 (O_2861,N_49862,N_49836);
xnor UO_2862 (O_2862,N_49963,N_49998);
or UO_2863 (O_2863,N_49767,N_49995);
and UO_2864 (O_2864,N_49888,N_49894);
xor UO_2865 (O_2865,N_49962,N_49959);
nor UO_2866 (O_2866,N_49775,N_49765);
nor UO_2867 (O_2867,N_49958,N_49753);
and UO_2868 (O_2868,N_49954,N_49837);
nor UO_2869 (O_2869,N_49979,N_49976);
nand UO_2870 (O_2870,N_49961,N_49833);
nand UO_2871 (O_2871,N_49772,N_49888);
nand UO_2872 (O_2872,N_49929,N_49815);
or UO_2873 (O_2873,N_49881,N_49920);
nor UO_2874 (O_2874,N_49905,N_49932);
and UO_2875 (O_2875,N_49912,N_49878);
nor UO_2876 (O_2876,N_49955,N_49759);
nor UO_2877 (O_2877,N_49836,N_49787);
nor UO_2878 (O_2878,N_49949,N_49914);
xor UO_2879 (O_2879,N_49932,N_49976);
and UO_2880 (O_2880,N_49935,N_49930);
nor UO_2881 (O_2881,N_49856,N_49811);
or UO_2882 (O_2882,N_49896,N_49850);
or UO_2883 (O_2883,N_49961,N_49785);
nand UO_2884 (O_2884,N_49988,N_49753);
and UO_2885 (O_2885,N_49833,N_49851);
nand UO_2886 (O_2886,N_49869,N_49843);
or UO_2887 (O_2887,N_49802,N_49835);
nor UO_2888 (O_2888,N_49894,N_49823);
nor UO_2889 (O_2889,N_49971,N_49884);
and UO_2890 (O_2890,N_49786,N_49922);
nor UO_2891 (O_2891,N_49920,N_49990);
or UO_2892 (O_2892,N_49952,N_49805);
nand UO_2893 (O_2893,N_49800,N_49806);
xnor UO_2894 (O_2894,N_49849,N_49800);
or UO_2895 (O_2895,N_49938,N_49809);
or UO_2896 (O_2896,N_49766,N_49939);
xnor UO_2897 (O_2897,N_49763,N_49866);
or UO_2898 (O_2898,N_49821,N_49920);
nor UO_2899 (O_2899,N_49770,N_49936);
or UO_2900 (O_2900,N_49844,N_49971);
xnor UO_2901 (O_2901,N_49896,N_49774);
nand UO_2902 (O_2902,N_49926,N_49969);
nor UO_2903 (O_2903,N_49873,N_49875);
xor UO_2904 (O_2904,N_49760,N_49962);
nor UO_2905 (O_2905,N_49855,N_49767);
nand UO_2906 (O_2906,N_49812,N_49897);
nor UO_2907 (O_2907,N_49855,N_49987);
xnor UO_2908 (O_2908,N_49816,N_49965);
and UO_2909 (O_2909,N_49848,N_49816);
or UO_2910 (O_2910,N_49807,N_49938);
or UO_2911 (O_2911,N_49752,N_49927);
nand UO_2912 (O_2912,N_49981,N_49813);
and UO_2913 (O_2913,N_49896,N_49867);
xnor UO_2914 (O_2914,N_49989,N_49882);
and UO_2915 (O_2915,N_49801,N_49838);
nor UO_2916 (O_2916,N_49766,N_49962);
and UO_2917 (O_2917,N_49826,N_49915);
nand UO_2918 (O_2918,N_49951,N_49969);
or UO_2919 (O_2919,N_49840,N_49944);
xor UO_2920 (O_2920,N_49753,N_49980);
or UO_2921 (O_2921,N_49763,N_49813);
nor UO_2922 (O_2922,N_49930,N_49947);
xor UO_2923 (O_2923,N_49912,N_49976);
xnor UO_2924 (O_2924,N_49903,N_49872);
and UO_2925 (O_2925,N_49925,N_49939);
nand UO_2926 (O_2926,N_49961,N_49846);
and UO_2927 (O_2927,N_49759,N_49894);
xnor UO_2928 (O_2928,N_49835,N_49978);
xor UO_2929 (O_2929,N_49823,N_49910);
or UO_2930 (O_2930,N_49773,N_49974);
xnor UO_2931 (O_2931,N_49811,N_49773);
xnor UO_2932 (O_2932,N_49915,N_49899);
xor UO_2933 (O_2933,N_49991,N_49805);
and UO_2934 (O_2934,N_49870,N_49804);
nor UO_2935 (O_2935,N_49997,N_49890);
xor UO_2936 (O_2936,N_49948,N_49866);
or UO_2937 (O_2937,N_49793,N_49849);
xor UO_2938 (O_2938,N_49894,N_49910);
nor UO_2939 (O_2939,N_49802,N_49788);
or UO_2940 (O_2940,N_49777,N_49815);
xor UO_2941 (O_2941,N_49956,N_49777);
nor UO_2942 (O_2942,N_49975,N_49914);
and UO_2943 (O_2943,N_49804,N_49993);
or UO_2944 (O_2944,N_49784,N_49796);
xor UO_2945 (O_2945,N_49990,N_49828);
and UO_2946 (O_2946,N_49886,N_49895);
nor UO_2947 (O_2947,N_49769,N_49806);
and UO_2948 (O_2948,N_49872,N_49979);
nor UO_2949 (O_2949,N_49811,N_49952);
nor UO_2950 (O_2950,N_49902,N_49781);
xor UO_2951 (O_2951,N_49761,N_49864);
xnor UO_2952 (O_2952,N_49887,N_49871);
xor UO_2953 (O_2953,N_49827,N_49964);
nand UO_2954 (O_2954,N_49824,N_49814);
and UO_2955 (O_2955,N_49752,N_49987);
xor UO_2956 (O_2956,N_49764,N_49798);
nand UO_2957 (O_2957,N_49813,N_49973);
or UO_2958 (O_2958,N_49755,N_49938);
or UO_2959 (O_2959,N_49850,N_49995);
and UO_2960 (O_2960,N_49996,N_49832);
nand UO_2961 (O_2961,N_49759,N_49951);
nand UO_2962 (O_2962,N_49764,N_49820);
and UO_2963 (O_2963,N_49809,N_49937);
xnor UO_2964 (O_2964,N_49882,N_49982);
nand UO_2965 (O_2965,N_49897,N_49888);
nor UO_2966 (O_2966,N_49993,N_49992);
nand UO_2967 (O_2967,N_49853,N_49870);
nand UO_2968 (O_2968,N_49840,N_49905);
nor UO_2969 (O_2969,N_49801,N_49862);
xor UO_2970 (O_2970,N_49792,N_49790);
nand UO_2971 (O_2971,N_49825,N_49959);
xnor UO_2972 (O_2972,N_49823,N_49879);
xor UO_2973 (O_2973,N_49830,N_49800);
and UO_2974 (O_2974,N_49864,N_49852);
and UO_2975 (O_2975,N_49962,N_49903);
nand UO_2976 (O_2976,N_49903,N_49773);
and UO_2977 (O_2977,N_49872,N_49867);
nand UO_2978 (O_2978,N_49784,N_49899);
and UO_2979 (O_2979,N_49860,N_49792);
xor UO_2980 (O_2980,N_49902,N_49774);
nor UO_2981 (O_2981,N_49896,N_49906);
or UO_2982 (O_2982,N_49778,N_49849);
nor UO_2983 (O_2983,N_49801,N_49850);
nor UO_2984 (O_2984,N_49767,N_49758);
or UO_2985 (O_2985,N_49867,N_49909);
and UO_2986 (O_2986,N_49759,N_49888);
and UO_2987 (O_2987,N_49932,N_49902);
nor UO_2988 (O_2988,N_49882,N_49956);
nand UO_2989 (O_2989,N_49874,N_49883);
and UO_2990 (O_2990,N_49967,N_49866);
and UO_2991 (O_2991,N_49972,N_49951);
xnor UO_2992 (O_2992,N_49938,N_49911);
and UO_2993 (O_2993,N_49824,N_49891);
and UO_2994 (O_2994,N_49942,N_49772);
xor UO_2995 (O_2995,N_49784,N_49917);
or UO_2996 (O_2996,N_49784,N_49978);
xnor UO_2997 (O_2997,N_49970,N_49847);
or UO_2998 (O_2998,N_49921,N_49994);
or UO_2999 (O_2999,N_49828,N_49844);
and UO_3000 (O_3000,N_49910,N_49831);
or UO_3001 (O_3001,N_49833,N_49872);
or UO_3002 (O_3002,N_49763,N_49860);
and UO_3003 (O_3003,N_49846,N_49750);
nand UO_3004 (O_3004,N_49882,N_49822);
and UO_3005 (O_3005,N_49777,N_49874);
and UO_3006 (O_3006,N_49841,N_49788);
nor UO_3007 (O_3007,N_49985,N_49851);
or UO_3008 (O_3008,N_49805,N_49750);
and UO_3009 (O_3009,N_49987,N_49936);
nor UO_3010 (O_3010,N_49963,N_49799);
and UO_3011 (O_3011,N_49842,N_49855);
or UO_3012 (O_3012,N_49930,N_49777);
or UO_3013 (O_3013,N_49946,N_49943);
nor UO_3014 (O_3014,N_49950,N_49764);
and UO_3015 (O_3015,N_49948,N_49808);
and UO_3016 (O_3016,N_49768,N_49985);
xor UO_3017 (O_3017,N_49803,N_49924);
nand UO_3018 (O_3018,N_49946,N_49819);
nor UO_3019 (O_3019,N_49848,N_49823);
xnor UO_3020 (O_3020,N_49754,N_49855);
nor UO_3021 (O_3021,N_49941,N_49922);
nor UO_3022 (O_3022,N_49955,N_49876);
xor UO_3023 (O_3023,N_49918,N_49995);
nand UO_3024 (O_3024,N_49945,N_49798);
xor UO_3025 (O_3025,N_49973,N_49837);
and UO_3026 (O_3026,N_49975,N_49853);
or UO_3027 (O_3027,N_49760,N_49922);
xnor UO_3028 (O_3028,N_49981,N_49763);
or UO_3029 (O_3029,N_49967,N_49970);
or UO_3030 (O_3030,N_49839,N_49909);
and UO_3031 (O_3031,N_49829,N_49765);
nor UO_3032 (O_3032,N_49983,N_49762);
nor UO_3033 (O_3033,N_49785,N_49790);
nand UO_3034 (O_3034,N_49827,N_49804);
nor UO_3035 (O_3035,N_49970,N_49769);
nor UO_3036 (O_3036,N_49985,N_49970);
xor UO_3037 (O_3037,N_49917,N_49900);
nand UO_3038 (O_3038,N_49965,N_49803);
and UO_3039 (O_3039,N_49939,N_49895);
and UO_3040 (O_3040,N_49977,N_49843);
or UO_3041 (O_3041,N_49751,N_49888);
nor UO_3042 (O_3042,N_49753,N_49990);
nand UO_3043 (O_3043,N_49853,N_49875);
nand UO_3044 (O_3044,N_49858,N_49929);
nand UO_3045 (O_3045,N_49891,N_49918);
nor UO_3046 (O_3046,N_49937,N_49843);
xnor UO_3047 (O_3047,N_49925,N_49952);
nand UO_3048 (O_3048,N_49981,N_49998);
or UO_3049 (O_3049,N_49862,N_49771);
or UO_3050 (O_3050,N_49962,N_49964);
nand UO_3051 (O_3051,N_49869,N_49834);
or UO_3052 (O_3052,N_49976,N_49806);
nor UO_3053 (O_3053,N_49963,N_49893);
nor UO_3054 (O_3054,N_49859,N_49906);
xnor UO_3055 (O_3055,N_49817,N_49985);
nor UO_3056 (O_3056,N_49911,N_49914);
or UO_3057 (O_3057,N_49863,N_49855);
nor UO_3058 (O_3058,N_49765,N_49819);
or UO_3059 (O_3059,N_49762,N_49956);
and UO_3060 (O_3060,N_49937,N_49918);
nand UO_3061 (O_3061,N_49944,N_49972);
nand UO_3062 (O_3062,N_49918,N_49811);
xnor UO_3063 (O_3063,N_49871,N_49781);
or UO_3064 (O_3064,N_49949,N_49794);
or UO_3065 (O_3065,N_49800,N_49929);
nor UO_3066 (O_3066,N_49896,N_49856);
nand UO_3067 (O_3067,N_49910,N_49822);
and UO_3068 (O_3068,N_49992,N_49907);
and UO_3069 (O_3069,N_49998,N_49864);
or UO_3070 (O_3070,N_49873,N_49882);
and UO_3071 (O_3071,N_49804,N_49759);
nor UO_3072 (O_3072,N_49900,N_49761);
or UO_3073 (O_3073,N_49885,N_49825);
nand UO_3074 (O_3074,N_49879,N_49762);
xor UO_3075 (O_3075,N_49774,N_49911);
nand UO_3076 (O_3076,N_49916,N_49877);
nand UO_3077 (O_3077,N_49798,N_49912);
xor UO_3078 (O_3078,N_49929,N_49935);
or UO_3079 (O_3079,N_49890,N_49993);
and UO_3080 (O_3080,N_49990,N_49955);
xnor UO_3081 (O_3081,N_49787,N_49855);
nor UO_3082 (O_3082,N_49803,N_49860);
or UO_3083 (O_3083,N_49924,N_49851);
nor UO_3084 (O_3084,N_49793,N_49944);
and UO_3085 (O_3085,N_49935,N_49829);
xnor UO_3086 (O_3086,N_49776,N_49861);
xnor UO_3087 (O_3087,N_49948,N_49793);
nand UO_3088 (O_3088,N_49797,N_49877);
or UO_3089 (O_3089,N_49931,N_49818);
nor UO_3090 (O_3090,N_49942,N_49872);
or UO_3091 (O_3091,N_49878,N_49785);
nor UO_3092 (O_3092,N_49885,N_49834);
xor UO_3093 (O_3093,N_49860,N_49993);
nor UO_3094 (O_3094,N_49897,N_49843);
nand UO_3095 (O_3095,N_49752,N_49893);
nor UO_3096 (O_3096,N_49975,N_49788);
nor UO_3097 (O_3097,N_49820,N_49842);
or UO_3098 (O_3098,N_49756,N_49912);
or UO_3099 (O_3099,N_49888,N_49831);
and UO_3100 (O_3100,N_49783,N_49772);
or UO_3101 (O_3101,N_49766,N_49761);
or UO_3102 (O_3102,N_49890,N_49766);
and UO_3103 (O_3103,N_49812,N_49818);
xnor UO_3104 (O_3104,N_49848,N_49981);
nor UO_3105 (O_3105,N_49791,N_49805);
nor UO_3106 (O_3106,N_49788,N_49842);
nor UO_3107 (O_3107,N_49913,N_49786);
nand UO_3108 (O_3108,N_49950,N_49751);
and UO_3109 (O_3109,N_49852,N_49896);
nor UO_3110 (O_3110,N_49958,N_49857);
nor UO_3111 (O_3111,N_49912,N_49981);
and UO_3112 (O_3112,N_49817,N_49809);
or UO_3113 (O_3113,N_49948,N_49825);
nand UO_3114 (O_3114,N_49810,N_49945);
and UO_3115 (O_3115,N_49828,N_49919);
nor UO_3116 (O_3116,N_49921,N_49910);
nand UO_3117 (O_3117,N_49999,N_49752);
xor UO_3118 (O_3118,N_49792,N_49875);
nor UO_3119 (O_3119,N_49846,N_49999);
xor UO_3120 (O_3120,N_49837,N_49886);
and UO_3121 (O_3121,N_49824,N_49870);
and UO_3122 (O_3122,N_49898,N_49936);
or UO_3123 (O_3123,N_49759,N_49859);
or UO_3124 (O_3124,N_49956,N_49881);
or UO_3125 (O_3125,N_49865,N_49820);
and UO_3126 (O_3126,N_49953,N_49860);
or UO_3127 (O_3127,N_49800,N_49947);
nand UO_3128 (O_3128,N_49907,N_49768);
nor UO_3129 (O_3129,N_49924,N_49945);
xor UO_3130 (O_3130,N_49890,N_49768);
or UO_3131 (O_3131,N_49956,N_49870);
nand UO_3132 (O_3132,N_49812,N_49836);
and UO_3133 (O_3133,N_49829,N_49990);
or UO_3134 (O_3134,N_49989,N_49825);
nor UO_3135 (O_3135,N_49926,N_49875);
or UO_3136 (O_3136,N_49919,N_49755);
nand UO_3137 (O_3137,N_49935,N_49795);
xnor UO_3138 (O_3138,N_49835,N_49993);
nor UO_3139 (O_3139,N_49827,N_49929);
or UO_3140 (O_3140,N_49777,N_49919);
nand UO_3141 (O_3141,N_49829,N_49755);
nor UO_3142 (O_3142,N_49991,N_49926);
nand UO_3143 (O_3143,N_49819,N_49965);
or UO_3144 (O_3144,N_49984,N_49803);
or UO_3145 (O_3145,N_49781,N_49841);
nand UO_3146 (O_3146,N_49861,N_49881);
or UO_3147 (O_3147,N_49775,N_49810);
or UO_3148 (O_3148,N_49780,N_49790);
xor UO_3149 (O_3149,N_49801,N_49907);
xor UO_3150 (O_3150,N_49946,N_49954);
nand UO_3151 (O_3151,N_49883,N_49966);
nand UO_3152 (O_3152,N_49751,N_49959);
or UO_3153 (O_3153,N_49978,N_49949);
or UO_3154 (O_3154,N_49768,N_49971);
nor UO_3155 (O_3155,N_49780,N_49810);
xnor UO_3156 (O_3156,N_49826,N_49820);
or UO_3157 (O_3157,N_49766,N_49835);
nor UO_3158 (O_3158,N_49790,N_49900);
nand UO_3159 (O_3159,N_49883,N_49977);
nand UO_3160 (O_3160,N_49777,N_49933);
nand UO_3161 (O_3161,N_49926,N_49889);
xor UO_3162 (O_3162,N_49844,N_49771);
and UO_3163 (O_3163,N_49759,N_49852);
and UO_3164 (O_3164,N_49975,N_49906);
nand UO_3165 (O_3165,N_49873,N_49760);
nand UO_3166 (O_3166,N_49973,N_49965);
and UO_3167 (O_3167,N_49808,N_49756);
nand UO_3168 (O_3168,N_49942,N_49917);
nor UO_3169 (O_3169,N_49850,N_49771);
nor UO_3170 (O_3170,N_49792,N_49933);
or UO_3171 (O_3171,N_49989,N_49768);
nor UO_3172 (O_3172,N_49982,N_49805);
nor UO_3173 (O_3173,N_49835,N_49921);
nor UO_3174 (O_3174,N_49772,N_49863);
nand UO_3175 (O_3175,N_49947,N_49839);
nor UO_3176 (O_3176,N_49791,N_49859);
nand UO_3177 (O_3177,N_49792,N_49999);
or UO_3178 (O_3178,N_49894,N_49893);
nand UO_3179 (O_3179,N_49989,N_49979);
xor UO_3180 (O_3180,N_49869,N_49991);
or UO_3181 (O_3181,N_49785,N_49904);
and UO_3182 (O_3182,N_49853,N_49809);
nand UO_3183 (O_3183,N_49783,N_49922);
nand UO_3184 (O_3184,N_49912,N_49863);
xor UO_3185 (O_3185,N_49988,N_49891);
and UO_3186 (O_3186,N_49806,N_49877);
and UO_3187 (O_3187,N_49979,N_49964);
nand UO_3188 (O_3188,N_49906,N_49954);
or UO_3189 (O_3189,N_49923,N_49822);
or UO_3190 (O_3190,N_49940,N_49784);
xnor UO_3191 (O_3191,N_49988,N_49949);
or UO_3192 (O_3192,N_49760,N_49776);
nand UO_3193 (O_3193,N_49773,N_49793);
nand UO_3194 (O_3194,N_49797,N_49992);
xor UO_3195 (O_3195,N_49998,N_49797);
xnor UO_3196 (O_3196,N_49890,N_49956);
xnor UO_3197 (O_3197,N_49814,N_49888);
nor UO_3198 (O_3198,N_49954,N_49917);
and UO_3199 (O_3199,N_49751,N_49842);
and UO_3200 (O_3200,N_49995,N_49814);
and UO_3201 (O_3201,N_49943,N_49781);
and UO_3202 (O_3202,N_49928,N_49979);
nand UO_3203 (O_3203,N_49938,N_49949);
xor UO_3204 (O_3204,N_49981,N_49997);
or UO_3205 (O_3205,N_49985,N_49863);
and UO_3206 (O_3206,N_49802,N_49808);
nor UO_3207 (O_3207,N_49875,N_49798);
and UO_3208 (O_3208,N_49795,N_49998);
nor UO_3209 (O_3209,N_49926,N_49858);
nand UO_3210 (O_3210,N_49860,N_49882);
nand UO_3211 (O_3211,N_49805,N_49773);
xnor UO_3212 (O_3212,N_49796,N_49763);
nor UO_3213 (O_3213,N_49828,N_49888);
xor UO_3214 (O_3214,N_49911,N_49775);
nor UO_3215 (O_3215,N_49811,N_49886);
nor UO_3216 (O_3216,N_49835,N_49776);
nor UO_3217 (O_3217,N_49873,N_49784);
or UO_3218 (O_3218,N_49923,N_49758);
nand UO_3219 (O_3219,N_49903,N_49899);
nand UO_3220 (O_3220,N_49976,N_49822);
nor UO_3221 (O_3221,N_49867,N_49865);
xor UO_3222 (O_3222,N_49763,N_49754);
xor UO_3223 (O_3223,N_49756,N_49904);
or UO_3224 (O_3224,N_49823,N_49950);
or UO_3225 (O_3225,N_49787,N_49908);
or UO_3226 (O_3226,N_49773,N_49790);
xnor UO_3227 (O_3227,N_49757,N_49853);
and UO_3228 (O_3228,N_49998,N_49771);
and UO_3229 (O_3229,N_49862,N_49938);
nand UO_3230 (O_3230,N_49914,N_49966);
nand UO_3231 (O_3231,N_49982,N_49759);
nor UO_3232 (O_3232,N_49975,N_49757);
nor UO_3233 (O_3233,N_49908,N_49918);
nand UO_3234 (O_3234,N_49968,N_49752);
or UO_3235 (O_3235,N_49773,N_49934);
and UO_3236 (O_3236,N_49972,N_49924);
xnor UO_3237 (O_3237,N_49975,N_49946);
nor UO_3238 (O_3238,N_49981,N_49983);
xor UO_3239 (O_3239,N_49947,N_49846);
nand UO_3240 (O_3240,N_49846,N_49919);
nor UO_3241 (O_3241,N_49771,N_49793);
nor UO_3242 (O_3242,N_49857,N_49823);
and UO_3243 (O_3243,N_49947,N_49865);
xor UO_3244 (O_3244,N_49785,N_49877);
and UO_3245 (O_3245,N_49790,N_49844);
nand UO_3246 (O_3246,N_49801,N_49855);
xor UO_3247 (O_3247,N_49819,N_49921);
nand UO_3248 (O_3248,N_49989,N_49837);
or UO_3249 (O_3249,N_49978,N_49895);
nand UO_3250 (O_3250,N_49881,N_49751);
nor UO_3251 (O_3251,N_49818,N_49906);
nor UO_3252 (O_3252,N_49844,N_49911);
or UO_3253 (O_3253,N_49768,N_49761);
and UO_3254 (O_3254,N_49903,N_49953);
nor UO_3255 (O_3255,N_49917,N_49943);
xnor UO_3256 (O_3256,N_49960,N_49860);
nand UO_3257 (O_3257,N_49787,N_49896);
nand UO_3258 (O_3258,N_49987,N_49791);
and UO_3259 (O_3259,N_49762,N_49774);
nand UO_3260 (O_3260,N_49995,N_49829);
nand UO_3261 (O_3261,N_49751,N_49861);
nand UO_3262 (O_3262,N_49982,N_49861);
nand UO_3263 (O_3263,N_49759,N_49846);
and UO_3264 (O_3264,N_49944,N_49986);
and UO_3265 (O_3265,N_49790,N_49783);
nand UO_3266 (O_3266,N_49787,N_49778);
nand UO_3267 (O_3267,N_49768,N_49859);
nand UO_3268 (O_3268,N_49844,N_49853);
xnor UO_3269 (O_3269,N_49791,N_49832);
nand UO_3270 (O_3270,N_49789,N_49965);
nor UO_3271 (O_3271,N_49953,N_49808);
nor UO_3272 (O_3272,N_49863,N_49751);
or UO_3273 (O_3273,N_49773,N_49906);
nor UO_3274 (O_3274,N_49792,N_49942);
or UO_3275 (O_3275,N_49869,N_49984);
or UO_3276 (O_3276,N_49899,N_49923);
xor UO_3277 (O_3277,N_49793,N_49764);
and UO_3278 (O_3278,N_49863,N_49874);
xnor UO_3279 (O_3279,N_49928,N_49878);
nor UO_3280 (O_3280,N_49882,N_49787);
xor UO_3281 (O_3281,N_49964,N_49924);
or UO_3282 (O_3282,N_49923,N_49961);
xor UO_3283 (O_3283,N_49842,N_49854);
nor UO_3284 (O_3284,N_49826,N_49836);
or UO_3285 (O_3285,N_49753,N_49831);
and UO_3286 (O_3286,N_49966,N_49908);
nor UO_3287 (O_3287,N_49801,N_49799);
or UO_3288 (O_3288,N_49950,N_49918);
and UO_3289 (O_3289,N_49936,N_49817);
nor UO_3290 (O_3290,N_49775,N_49897);
and UO_3291 (O_3291,N_49772,N_49768);
nand UO_3292 (O_3292,N_49966,N_49798);
nand UO_3293 (O_3293,N_49995,N_49792);
nor UO_3294 (O_3294,N_49870,N_49948);
nand UO_3295 (O_3295,N_49875,N_49829);
xor UO_3296 (O_3296,N_49802,N_49826);
nor UO_3297 (O_3297,N_49862,N_49952);
nor UO_3298 (O_3298,N_49870,N_49950);
and UO_3299 (O_3299,N_49978,N_49873);
nand UO_3300 (O_3300,N_49859,N_49989);
xnor UO_3301 (O_3301,N_49784,N_49765);
xor UO_3302 (O_3302,N_49795,N_49904);
xor UO_3303 (O_3303,N_49952,N_49908);
or UO_3304 (O_3304,N_49901,N_49921);
nand UO_3305 (O_3305,N_49881,N_49813);
or UO_3306 (O_3306,N_49874,N_49923);
nor UO_3307 (O_3307,N_49955,N_49918);
xor UO_3308 (O_3308,N_49988,N_49856);
and UO_3309 (O_3309,N_49928,N_49805);
nand UO_3310 (O_3310,N_49880,N_49800);
or UO_3311 (O_3311,N_49854,N_49821);
nand UO_3312 (O_3312,N_49849,N_49920);
or UO_3313 (O_3313,N_49974,N_49987);
xnor UO_3314 (O_3314,N_49961,N_49791);
or UO_3315 (O_3315,N_49761,N_49972);
and UO_3316 (O_3316,N_49849,N_49927);
xnor UO_3317 (O_3317,N_49791,N_49849);
nand UO_3318 (O_3318,N_49852,N_49809);
and UO_3319 (O_3319,N_49948,N_49978);
nor UO_3320 (O_3320,N_49969,N_49836);
nor UO_3321 (O_3321,N_49999,N_49849);
xnor UO_3322 (O_3322,N_49756,N_49989);
nand UO_3323 (O_3323,N_49822,N_49875);
xnor UO_3324 (O_3324,N_49802,N_49904);
or UO_3325 (O_3325,N_49989,N_49886);
nand UO_3326 (O_3326,N_49996,N_49790);
or UO_3327 (O_3327,N_49978,N_49772);
nor UO_3328 (O_3328,N_49970,N_49886);
nand UO_3329 (O_3329,N_49754,N_49846);
nor UO_3330 (O_3330,N_49962,N_49884);
nand UO_3331 (O_3331,N_49947,N_49933);
and UO_3332 (O_3332,N_49988,N_49769);
nand UO_3333 (O_3333,N_49895,N_49917);
and UO_3334 (O_3334,N_49996,N_49783);
xor UO_3335 (O_3335,N_49961,N_49776);
xor UO_3336 (O_3336,N_49812,N_49918);
and UO_3337 (O_3337,N_49919,N_49885);
or UO_3338 (O_3338,N_49771,N_49796);
xor UO_3339 (O_3339,N_49944,N_49875);
and UO_3340 (O_3340,N_49916,N_49856);
xnor UO_3341 (O_3341,N_49930,N_49899);
nor UO_3342 (O_3342,N_49832,N_49828);
xor UO_3343 (O_3343,N_49872,N_49997);
and UO_3344 (O_3344,N_49952,N_49984);
nand UO_3345 (O_3345,N_49933,N_49951);
nor UO_3346 (O_3346,N_49858,N_49962);
or UO_3347 (O_3347,N_49987,N_49770);
xnor UO_3348 (O_3348,N_49751,N_49885);
nor UO_3349 (O_3349,N_49884,N_49949);
or UO_3350 (O_3350,N_49811,N_49961);
xor UO_3351 (O_3351,N_49858,N_49852);
xor UO_3352 (O_3352,N_49947,N_49889);
and UO_3353 (O_3353,N_49887,N_49933);
nor UO_3354 (O_3354,N_49962,N_49849);
xor UO_3355 (O_3355,N_49848,N_49997);
nor UO_3356 (O_3356,N_49930,N_49933);
nand UO_3357 (O_3357,N_49784,N_49982);
xnor UO_3358 (O_3358,N_49818,N_49998);
nor UO_3359 (O_3359,N_49792,N_49755);
nor UO_3360 (O_3360,N_49988,N_49823);
or UO_3361 (O_3361,N_49811,N_49957);
nor UO_3362 (O_3362,N_49760,N_49779);
xor UO_3363 (O_3363,N_49895,N_49950);
or UO_3364 (O_3364,N_49818,N_49905);
nor UO_3365 (O_3365,N_49882,N_49892);
and UO_3366 (O_3366,N_49895,N_49798);
nand UO_3367 (O_3367,N_49998,N_49949);
or UO_3368 (O_3368,N_49846,N_49767);
or UO_3369 (O_3369,N_49895,N_49884);
nor UO_3370 (O_3370,N_49928,N_49766);
xor UO_3371 (O_3371,N_49824,N_49861);
and UO_3372 (O_3372,N_49918,N_49800);
and UO_3373 (O_3373,N_49905,N_49990);
xnor UO_3374 (O_3374,N_49842,N_49946);
xor UO_3375 (O_3375,N_49979,N_49782);
xnor UO_3376 (O_3376,N_49792,N_49822);
or UO_3377 (O_3377,N_49783,N_49914);
and UO_3378 (O_3378,N_49752,N_49914);
nor UO_3379 (O_3379,N_49855,N_49760);
xor UO_3380 (O_3380,N_49972,N_49844);
or UO_3381 (O_3381,N_49822,N_49987);
nor UO_3382 (O_3382,N_49885,N_49817);
xnor UO_3383 (O_3383,N_49822,N_49841);
or UO_3384 (O_3384,N_49967,N_49989);
nand UO_3385 (O_3385,N_49940,N_49932);
and UO_3386 (O_3386,N_49808,N_49853);
nand UO_3387 (O_3387,N_49803,N_49868);
or UO_3388 (O_3388,N_49854,N_49859);
xor UO_3389 (O_3389,N_49860,N_49990);
nor UO_3390 (O_3390,N_49941,N_49978);
and UO_3391 (O_3391,N_49842,N_49771);
nor UO_3392 (O_3392,N_49889,N_49784);
and UO_3393 (O_3393,N_49970,N_49753);
or UO_3394 (O_3394,N_49759,N_49930);
and UO_3395 (O_3395,N_49850,N_49784);
and UO_3396 (O_3396,N_49843,N_49889);
and UO_3397 (O_3397,N_49900,N_49788);
or UO_3398 (O_3398,N_49935,N_49850);
or UO_3399 (O_3399,N_49941,N_49935);
and UO_3400 (O_3400,N_49763,N_49963);
nor UO_3401 (O_3401,N_49971,N_49847);
nor UO_3402 (O_3402,N_49954,N_49927);
or UO_3403 (O_3403,N_49956,N_49889);
and UO_3404 (O_3404,N_49853,N_49834);
nor UO_3405 (O_3405,N_49791,N_49780);
or UO_3406 (O_3406,N_49956,N_49936);
and UO_3407 (O_3407,N_49812,N_49775);
and UO_3408 (O_3408,N_49948,N_49910);
nor UO_3409 (O_3409,N_49832,N_49906);
nor UO_3410 (O_3410,N_49903,N_49811);
or UO_3411 (O_3411,N_49929,N_49936);
nor UO_3412 (O_3412,N_49896,N_49772);
nand UO_3413 (O_3413,N_49811,N_49978);
or UO_3414 (O_3414,N_49752,N_49838);
and UO_3415 (O_3415,N_49920,N_49980);
nand UO_3416 (O_3416,N_49951,N_49803);
nand UO_3417 (O_3417,N_49997,N_49843);
xnor UO_3418 (O_3418,N_49822,N_49878);
nor UO_3419 (O_3419,N_49955,N_49867);
xor UO_3420 (O_3420,N_49788,N_49954);
nand UO_3421 (O_3421,N_49976,N_49989);
nor UO_3422 (O_3422,N_49944,N_49926);
nor UO_3423 (O_3423,N_49815,N_49920);
or UO_3424 (O_3424,N_49865,N_49997);
and UO_3425 (O_3425,N_49885,N_49800);
xnor UO_3426 (O_3426,N_49787,N_49775);
and UO_3427 (O_3427,N_49758,N_49907);
and UO_3428 (O_3428,N_49977,N_49784);
xnor UO_3429 (O_3429,N_49889,N_49814);
nand UO_3430 (O_3430,N_49842,N_49754);
or UO_3431 (O_3431,N_49753,N_49870);
nand UO_3432 (O_3432,N_49798,N_49840);
nor UO_3433 (O_3433,N_49824,N_49875);
nor UO_3434 (O_3434,N_49927,N_49873);
nor UO_3435 (O_3435,N_49805,N_49898);
nand UO_3436 (O_3436,N_49774,N_49798);
or UO_3437 (O_3437,N_49980,N_49815);
nor UO_3438 (O_3438,N_49954,N_49988);
nand UO_3439 (O_3439,N_49883,N_49930);
nor UO_3440 (O_3440,N_49798,N_49760);
xnor UO_3441 (O_3441,N_49824,N_49930);
nand UO_3442 (O_3442,N_49885,N_49944);
and UO_3443 (O_3443,N_49829,N_49949);
or UO_3444 (O_3444,N_49805,N_49871);
and UO_3445 (O_3445,N_49945,N_49993);
nor UO_3446 (O_3446,N_49785,N_49993);
or UO_3447 (O_3447,N_49827,N_49792);
nor UO_3448 (O_3448,N_49962,N_49833);
or UO_3449 (O_3449,N_49772,N_49817);
nand UO_3450 (O_3450,N_49985,N_49777);
nand UO_3451 (O_3451,N_49994,N_49804);
nand UO_3452 (O_3452,N_49877,N_49926);
nand UO_3453 (O_3453,N_49896,N_49909);
nor UO_3454 (O_3454,N_49810,N_49814);
nand UO_3455 (O_3455,N_49898,N_49789);
or UO_3456 (O_3456,N_49998,N_49804);
and UO_3457 (O_3457,N_49799,N_49763);
or UO_3458 (O_3458,N_49950,N_49882);
xor UO_3459 (O_3459,N_49992,N_49893);
nor UO_3460 (O_3460,N_49969,N_49804);
and UO_3461 (O_3461,N_49853,N_49934);
and UO_3462 (O_3462,N_49896,N_49770);
or UO_3463 (O_3463,N_49885,N_49983);
nor UO_3464 (O_3464,N_49871,N_49796);
and UO_3465 (O_3465,N_49815,N_49914);
nor UO_3466 (O_3466,N_49784,N_49871);
nor UO_3467 (O_3467,N_49966,N_49824);
and UO_3468 (O_3468,N_49815,N_49999);
and UO_3469 (O_3469,N_49960,N_49911);
nand UO_3470 (O_3470,N_49752,N_49807);
or UO_3471 (O_3471,N_49820,N_49894);
xnor UO_3472 (O_3472,N_49766,N_49976);
and UO_3473 (O_3473,N_49998,N_49793);
and UO_3474 (O_3474,N_49963,N_49791);
and UO_3475 (O_3475,N_49928,N_49968);
nor UO_3476 (O_3476,N_49899,N_49882);
or UO_3477 (O_3477,N_49801,N_49952);
and UO_3478 (O_3478,N_49754,N_49960);
nor UO_3479 (O_3479,N_49790,N_49878);
nor UO_3480 (O_3480,N_49814,N_49772);
and UO_3481 (O_3481,N_49789,N_49824);
nand UO_3482 (O_3482,N_49902,N_49762);
nor UO_3483 (O_3483,N_49960,N_49807);
nand UO_3484 (O_3484,N_49975,N_49841);
xnor UO_3485 (O_3485,N_49992,N_49954);
nand UO_3486 (O_3486,N_49793,N_49822);
nor UO_3487 (O_3487,N_49926,N_49796);
xnor UO_3488 (O_3488,N_49922,N_49770);
nand UO_3489 (O_3489,N_49858,N_49979);
or UO_3490 (O_3490,N_49896,N_49803);
xor UO_3491 (O_3491,N_49973,N_49795);
xnor UO_3492 (O_3492,N_49842,N_49988);
and UO_3493 (O_3493,N_49964,N_49905);
xnor UO_3494 (O_3494,N_49789,N_49869);
nor UO_3495 (O_3495,N_49987,N_49761);
nor UO_3496 (O_3496,N_49918,N_49894);
nor UO_3497 (O_3497,N_49999,N_49774);
or UO_3498 (O_3498,N_49998,N_49762);
or UO_3499 (O_3499,N_49897,N_49827);
and UO_3500 (O_3500,N_49782,N_49900);
nor UO_3501 (O_3501,N_49758,N_49806);
xnor UO_3502 (O_3502,N_49774,N_49899);
nor UO_3503 (O_3503,N_49968,N_49861);
xnor UO_3504 (O_3504,N_49856,N_49826);
xor UO_3505 (O_3505,N_49814,N_49951);
nand UO_3506 (O_3506,N_49832,N_49750);
and UO_3507 (O_3507,N_49804,N_49818);
or UO_3508 (O_3508,N_49790,N_49826);
xnor UO_3509 (O_3509,N_49767,N_49880);
and UO_3510 (O_3510,N_49816,N_49977);
or UO_3511 (O_3511,N_49818,N_49885);
nor UO_3512 (O_3512,N_49890,N_49771);
xor UO_3513 (O_3513,N_49778,N_49802);
xor UO_3514 (O_3514,N_49902,N_49874);
and UO_3515 (O_3515,N_49860,N_49774);
nor UO_3516 (O_3516,N_49894,N_49775);
nand UO_3517 (O_3517,N_49857,N_49951);
and UO_3518 (O_3518,N_49912,N_49759);
and UO_3519 (O_3519,N_49915,N_49851);
nand UO_3520 (O_3520,N_49807,N_49834);
nor UO_3521 (O_3521,N_49750,N_49790);
nor UO_3522 (O_3522,N_49765,N_49758);
nor UO_3523 (O_3523,N_49969,N_49920);
xor UO_3524 (O_3524,N_49870,N_49823);
or UO_3525 (O_3525,N_49920,N_49752);
nand UO_3526 (O_3526,N_49948,N_49788);
or UO_3527 (O_3527,N_49963,N_49974);
nor UO_3528 (O_3528,N_49914,N_49987);
nor UO_3529 (O_3529,N_49857,N_49808);
xor UO_3530 (O_3530,N_49871,N_49799);
or UO_3531 (O_3531,N_49766,N_49812);
xnor UO_3532 (O_3532,N_49916,N_49760);
nor UO_3533 (O_3533,N_49951,N_49947);
and UO_3534 (O_3534,N_49890,N_49920);
nand UO_3535 (O_3535,N_49945,N_49807);
and UO_3536 (O_3536,N_49943,N_49995);
and UO_3537 (O_3537,N_49940,N_49909);
nand UO_3538 (O_3538,N_49770,N_49932);
nor UO_3539 (O_3539,N_49973,N_49863);
or UO_3540 (O_3540,N_49907,N_49810);
and UO_3541 (O_3541,N_49795,N_49757);
xor UO_3542 (O_3542,N_49950,N_49856);
and UO_3543 (O_3543,N_49785,N_49963);
or UO_3544 (O_3544,N_49792,N_49830);
nor UO_3545 (O_3545,N_49828,N_49754);
nand UO_3546 (O_3546,N_49910,N_49767);
nand UO_3547 (O_3547,N_49925,N_49960);
or UO_3548 (O_3548,N_49892,N_49781);
nor UO_3549 (O_3549,N_49758,N_49896);
or UO_3550 (O_3550,N_49897,N_49844);
nor UO_3551 (O_3551,N_49805,N_49899);
xor UO_3552 (O_3552,N_49760,N_49836);
xnor UO_3553 (O_3553,N_49764,N_49997);
nand UO_3554 (O_3554,N_49767,N_49986);
nor UO_3555 (O_3555,N_49935,N_49826);
nand UO_3556 (O_3556,N_49949,N_49754);
xor UO_3557 (O_3557,N_49907,N_49881);
or UO_3558 (O_3558,N_49765,N_49843);
or UO_3559 (O_3559,N_49909,N_49964);
and UO_3560 (O_3560,N_49788,N_49772);
and UO_3561 (O_3561,N_49887,N_49953);
and UO_3562 (O_3562,N_49836,N_49785);
nor UO_3563 (O_3563,N_49989,N_49751);
or UO_3564 (O_3564,N_49883,N_49904);
or UO_3565 (O_3565,N_49888,N_49941);
or UO_3566 (O_3566,N_49948,N_49906);
xnor UO_3567 (O_3567,N_49918,N_49873);
xor UO_3568 (O_3568,N_49971,N_49975);
nand UO_3569 (O_3569,N_49880,N_49914);
or UO_3570 (O_3570,N_49812,N_49982);
and UO_3571 (O_3571,N_49769,N_49996);
nor UO_3572 (O_3572,N_49783,N_49848);
nand UO_3573 (O_3573,N_49968,N_49981);
xnor UO_3574 (O_3574,N_49849,N_49769);
nand UO_3575 (O_3575,N_49871,N_49851);
nor UO_3576 (O_3576,N_49866,N_49926);
xnor UO_3577 (O_3577,N_49755,N_49922);
xor UO_3578 (O_3578,N_49750,N_49981);
nand UO_3579 (O_3579,N_49840,N_49938);
and UO_3580 (O_3580,N_49757,N_49918);
nor UO_3581 (O_3581,N_49829,N_49751);
nor UO_3582 (O_3582,N_49965,N_49792);
or UO_3583 (O_3583,N_49933,N_49931);
xor UO_3584 (O_3584,N_49814,N_49853);
nor UO_3585 (O_3585,N_49985,N_49997);
nor UO_3586 (O_3586,N_49956,N_49766);
xor UO_3587 (O_3587,N_49906,N_49761);
xnor UO_3588 (O_3588,N_49970,N_49974);
and UO_3589 (O_3589,N_49985,N_49979);
xnor UO_3590 (O_3590,N_49828,N_49863);
nand UO_3591 (O_3591,N_49840,N_49926);
and UO_3592 (O_3592,N_49919,N_49949);
nand UO_3593 (O_3593,N_49956,N_49937);
or UO_3594 (O_3594,N_49902,N_49884);
or UO_3595 (O_3595,N_49917,N_49855);
nor UO_3596 (O_3596,N_49879,N_49928);
nor UO_3597 (O_3597,N_49793,N_49917);
nor UO_3598 (O_3598,N_49790,N_49820);
or UO_3599 (O_3599,N_49775,N_49922);
nand UO_3600 (O_3600,N_49751,N_49818);
nor UO_3601 (O_3601,N_49996,N_49761);
and UO_3602 (O_3602,N_49762,N_49895);
nand UO_3603 (O_3603,N_49839,N_49863);
nand UO_3604 (O_3604,N_49946,N_49937);
and UO_3605 (O_3605,N_49936,N_49999);
and UO_3606 (O_3606,N_49813,N_49897);
nor UO_3607 (O_3607,N_49858,N_49911);
nor UO_3608 (O_3608,N_49898,N_49802);
and UO_3609 (O_3609,N_49960,N_49897);
or UO_3610 (O_3610,N_49815,N_49875);
nand UO_3611 (O_3611,N_49985,N_49883);
and UO_3612 (O_3612,N_49941,N_49972);
xnor UO_3613 (O_3613,N_49782,N_49886);
nor UO_3614 (O_3614,N_49951,N_49991);
nand UO_3615 (O_3615,N_49842,N_49835);
or UO_3616 (O_3616,N_49854,N_49932);
nor UO_3617 (O_3617,N_49881,N_49940);
nor UO_3618 (O_3618,N_49978,N_49807);
and UO_3619 (O_3619,N_49780,N_49761);
nor UO_3620 (O_3620,N_49762,N_49793);
or UO_3621 (O_3621,N_49995,N_49925);
xor UO_3622 (O_3622,N_49776,N_49946);
or UO_3623 (O_3623,N_49869,N_49840);
xnor UO_3624 (O_3624,N_49774,N_49918);
or UO_3625 (O_3625,N_49871,N_49911);
or UO_3626 (O_3626,N_49844,N_49904);
xor UO_3627 (O_3627,N_49991,N_49923);
nand UO_3628 (O_3628,N_49910,N_49819);
nand UO_3629 (O_3629,N_49824,N_49878);
nor UO_3630 (O_3630,N_49958,N_49916);
nand UO_3631 (O_3631,N_49931,N_49792);
and UO_3632 (O_3632,N_49962,N_49994);
nor UO_3633 (O_3633,N_49852,N_49935);
nand UO_3634 (O_3634,N_49799,N_49902);
xor UO_3635 (O_3635,N_49916,N_49892);
xor UO_3636 (O_3636,N_49992,N_49910);
xnor UO_3637 (O_3637,N_49839,N_49784);
nand UO_3638 (O_3638,N_49868,N_49980);
xnor UO_3639 (O_3639,N_49791,N_49997);
nand UO_3640 (O_3640,N_49760,N_49827);
xnor UO_3641 (O_3641,N_49844,N_49936);
or UO_3642 (O_3642,N_49917,N_49785);
or UO_3643 (O_3643,N_49892,N_49938);
or UO_3644 (O_3644,N_49860,N_49918);
or UO_3645 (O_3645,N_49929,N_49805);
or UO_3646 (O_3646,N_49897,N_49855);
nand UO_3647 (O_3647,N_49824,N_49812);
xnor UO_3648 (O_3648,N_49905,N_49948);
nand UO_3649 (O_3649,N_49869,N_49910);
xor UO_3650 (O_3650,N_49935,N_49937);
nor UO_3651 (O_3651,N_49826,N_49791);
nor UO_3652 (O_3652,N_49945,N_49979);
or UO_3653 (O_3653,N_49780,N_49845);
nand UO_3654 (O_3654,N_49861,N_49836);
nor UO_3655 (O_3655,N_49908,N_49811);
or UO_3656 (O_3656,N_49856,N_49855);
and UO_3657 (O_3657,N_49851,N_49834);
xnor UO_3658 (O_3658,N_49989,N_49998);
or UO_3659 (O_3659,N_49835,N_49893);
nor UO_3660 (O_3660,N_49818,N_49775);
nor UO_3661 (O_3661,N_49782,N_49763);
nor UO_3662 (O_3662,N_49823,N_49855);
xnor UO_3663 (O_3663,N_49767,N_49893);
xnor UO_3664 (O_3664,N_49933,N_49917);
nand UO_3665 (O_3665,N_49816,N_49843);
nor UO_3666 (O_3666,N_49907,N_49939);
or UO_3667 (O_3667,N_49803,N_49824);
nor UO_3668 (O_3668,N_49953,N_49922);
nand UO_3669 (O_3669,N_49881,N_49811);
and UO_3670 (O_3670,N_49928,N_49953);
xor UO_3671 (O_3671,N_49908,N_49797);
and UO_3672 (O_3672,N_49826,N_49913);
or UO_3673 (O_3673,N_49836,N_49960);
xor UO_3674 (O_3674,N_49891,N_49768);
nand UO_3675 (O_3675,N_49858,N_49894);
nor UO_3676 (O_3676,N_49987,N_49777);
or UO_3677 (O_3677,N_49837,N_49852);
nor UO_3678 (O_3678,N_49972,N_49773);
nor UO_3679 (O_3679,N_49896,N_49789);
xor UO_3680 (O_3680,N_49787,N_49831);
nor UO_3681 (O_3681,N_49869,N_49962);
or UO_3682 (O_3682,N_49799,N_49784);
nand UO_3683 (O_3683,N_49947,N_49921);
and UO_3684 (O_3684,N_49965,N_49972);
xnor UO_3685 (O_3685,N_49843,N_49971);
or UO_3686 (O_3686,N_49822,N_49813);
and UO_3687 (O_3687,N_49900,N_49813);
nor UO_3688 (O_3688,N_49894,N_49886);
or UO_3689 (O_3689,N_49938,N_49818);
or UO_3690 (O_3690,N_49887,N_49950);
or UO_3691 (O_3691,N_49843,N_49805);
xor UO_3692 (O_3692,N_49833,N_49757);
and UO_3693 (O_3693,N_49862,N_49976);
and UO_3694 (O_3694,N_49869,N_49846);
and UO_3695 (O_3695,N_49819,N_49903);
and UO_3696 (O_3696,N_49923,N_49761);
and UO_3697 (O_3697,N_49924,N_49816);
nand UO_3698 (O_3698,N_49859,N_49863);
and UO_3699 (O_3699,N_49966,N_49791);
and UO_3700 (O_3700,N_49800,N_49919);
and UO_3701 (O_3701,N_49957,N_49891);
and UO_3702 (O_3702,N_49823,N_49780);
xnor UO_3703 (O_3703,N_49776,N_49878);
nand UO_3704 (O_3704,N_49754,N_49779);
and UO_3705 (O_3705,N_49991,N_49811);
xnor UO_3706 (O_3706,N_49870,N_49860);
nor UO_3707 (O_3707,N_49754,N_49920);
xnor UO_3708 (O_3708,N_49944,N_49824);
nor UO_3709 (O_3709,N_49860,N_49777);
nor UO_3710 (O_3710,N_49999,N_49895);
xnor UO_3711 (O_3711,N_49824,N_49772);
nor UO_3712 (O_3712,N_49789,N_49768);
nor UO_3713 (O_3713,N_49818,N_49912);
nand UO_3714 (O_3714,N_49976,N_49777);
and UO_3715 (O_3715,N_49872,N_49909);
nor UO_3716 (O_3716,N_49823,N_49980);
nand UO_3717 (O_3717,N_49883,N_49756);
nand UO_3718 (O_3718,N_49894,N_49983);
nand UO_3719 (O_3719,N_49768,N_49837);
and UO_3720 (O_3720,N_49811,N_49753);
and UO_3721 (O_3721,N_49875,N_49936);
or UO_3722 (O_3722,N_49768,N_49993);
and UO_3723 (O_3723,N_49895,N_49888);
and UO_3724 (O_3724,N_49841,N_49794);
xnor UO_3725 (O_3725,N_49912,N_49861);
nand UO_3726 (O_3726,N_49885,N_49786);
nor UO_3727 (O_3727,N_49850,N_49857);
nor UO_3728 (O_3728,N_49955,N_49768);
xnor UO_3729 (O_3729,N_49987,N_49859);
nor UO_3730 (O_3730,N_49936,N_49953);
nor UO_3731 (O_3731,N_49945,N_49801);
and UO_3732 (O_3732,N_49856,N_49894);
xnor UO_3733 (O_3733,N_49985,N_49829);
nand UO_3734 (O_3734,N_49894,N_49835);
or UO_3735 (O_3735,N_49803,N_49762);
xnor UO_3736 (O_3736,N_49979,N_49823);
and UO_3737 (O_3737,N_49942,N_49924);
and UO_3738 (O_3738,N_49982,N_49802);
xor UO_3739 (O_3739,N_49890,N_49859);
xor UO_3740 (O_3740,N_49788,N_49860);
nor UO_3741 (O_3741,N_49940,N_49786);
xnor UO_3742 (O_3742,N_49880,N_49905);
xnor UO_3743 (O_3743,N_49950,N_49940);
xor UO_3744 (O_3744,N_49994,N_49990);
or UO_3745 (O_3745,N_49808,N_49761);
nand UO_3746 (O_3746,N_49870,N_49767);
xnor UO_3747 (O_3747,N_49875,N_49872);
and UO_3748 (O_3748,N_49756,N_49851);
nand UO_3749 (O_3749,N_49794,N_49751);
and UO_3750 (O_3750,N_49801,N_49992);
nor UO_3751 (O_3751,N_49798,N_49943);
nand UO_3752 (O_3752,N_49772,N_49762);
or UO_3753 (O_3753,N_49949,N_49991);
xor UO_3754 (O_3754,N_49785,N_49987);
nor UO_3755 (O_3755,N_49894,N_49980);
xnor UO_3756 (O_3756,N_49953,N_49810);
or UO_3757 (O_3757,N_49923,N_49949);
and UO_3758 (O_3758,N_49751,N_49785);
nand UO_3759 (O_3759,N_49945,N_49866);
nand UO_3760 (O_3760,N_49836,N_49775);
and UO_3761 (O_3761,N_49845,N_49945);
or UO_3762 (O_3762,N_49943,N_49974);
nand UO_3763 (O_3763,N_49854,N_49970);
xor UO_3764 (O_3764,N_49815,N_49944);
nand UO_3765 (O_3765,N_49963,N_49820);
xor UO_3766 (O_3766,N_49889,N_49868);
and UO_3767 (O_3767,N_49798,N_49944);
nor UO_3768 (O_3768,N_49842,N_49793);
nand UO_3769 (O_3769,N_49965,N_49832);
and UO_3770 (O_3770,N_49965,N_49798);
nand UO_3771 (O_3771,N_49974,N_49879);
or UO_3772 (O_3772,N_49758,N_49802);
nand UO_3773 (O_3773,N_49829,N_49968);
and UO_3774 (O_3774,N_49944,N_49829);
and UO_3775 (O_3775,N_49832,N_49807);
nor UO_3776 (O_3776,N_49932,N_49823);
nor UO_3777 (O_3777,N_49991,N_49853);
xor UO_3778 (O_3778,N_49788,N_49924);
nor UO_3779 (O_3779,N_49945,N_49851);
nand UO_3780 (O_3780,N_49848,N_49758);
nand UO_3781 (O_3781,N_49762,N_49829);
xor UO_3782 (O_3782,N_49775,N_49969);
xnor UO_3783 (O_3783,N_49969,N_49960);
or UO_3784 (O_3784,N_49771,N_49879);
and UO_3785 (O_3785,N_49895,N_49932);
and UO_3786 (O_3786,N_49841,N_49885);
xor UO_3787 (O_3787,N_49977,N_49913);
xor UO_3788 (O_3788,N_49997,N_49960);
nor UO_3789 (O_3789,N_49872,N_49977);
nor UO_3790 (O_3790,N_49758,N_49951);
nand UO_3791 (O_3791,N_49938,N_49900);
and UO_3792 (O_3792,N_49864,N_49937);
xnor UO_3793 (O_3793,N_49950,N_49941);
or UO_3794 (O_3794,N_49960,N_49870);
or UO_3795 (O_3795,N_49889,N_49788);
and UO_3796 (O_3796,N_49761,N_49757);
or UO_3797 (O_3797,N_49951,N_49880);
and UO_3798 (O_3798,N_49808,N_49787);
xor UO_3799 (O_3799,N_49782,N_49777);
and UO_3800 (O_3800,N_49987,N_49908);
nand UO_3801 (O_3801,N_49828,N_49976);
nor UO_3802 (O_3802,N_49823,N_49977);
or UO_3803 (O_3803,N_49962,N_49927);
xnor UO_3804 (O_3804,N_49961,N_49965);
nand UO_3805 (O_3805,N_49782,N_49933);
nand UO_3806 (O_3806,N_49938,N_49916);
nor UO_3807 (O_3807,N_49953,N_49812);
xnor UO_3808 (O_3808,N_49931,N_49926);
and UO_3809 (O_3809,N_49871,N_49931);
nor UO_3810 (O_3810,N_49783,N_49959);
nor UO_3811 (O_3811,N_49815,N_49907);
nand UO_3812 (O_3812,N_49872,N_49785);
nand UO_3813 (O_3813,N_49899,N_49963);
or UO_3814 (O_3814,N_49848,N_49854);
nand UO_3815 (O_3815,N_49898,N_49990);
and UO_3816 (O_3816,N_49871,N_49895);
nor UO_3817 (O_3817,N_49857,N_49869);
and UO_3818 (O_3818,N_49785,N_49796);
and UO_3819 (O_3819,N_49764,N_49869);
xor UO_3820 (O_3820,N_49949,N_49940);
and UO_3821 (O_3821,N_49951,N_49916);
or UO_3822 (O_3822,N_49949,N_49862);
or UO_3823 (O_3823,N_49934,N_49780);
nor UO_3824 (O_3824,N_49831,N_49940);
or UO_3825 (O_3825,N_49919,N_49971);
xnor UO_3826 (O_3826,N_49797,N_49883);
and UO_3827 (O_3827,N_49750,N_49794);
nand UO_3828 (O_3828,N_49825,N_49853);
xnor UO_3829 (O_3829,N_49755,N_49966);
nor UO_3830 (O_3830,N_49961,N_49821);
nor UO_3831 (O_3831,N_49970,N_49838);
xnor UO_3832 (O_3832,N_49853,N_49971);
nor UO_3833 (O_3833,N_49808,N_49967);
nor UO_3834 (O_3834,N_49873,N_49824);
and UO_3835 (O_3835,N_49806,N_49897);
nand UO_3836 (O_3836,N_49815,N_49878);
or UO_3837 (O_3837,N_49848,N_49878);
nand UO_3838 (O_3838,N_49912,N_49880);
and UO_3839 (O_3839,N_49902,N_49920);
and UO_3840 (O_3840,N_49982,N_49793);
or UO_3841 (O_3841,N_49877,N_49839);
xor UO_3842 (O_3842,N_49835,N_49762);
nand UO_3843 (O_3843,N_49789,N_49968);
or UO_3844 (O_3844,N_49858,N_49889);
or UO_3845 (O_3845,N_49962,N_49898);
nand UO_3846 (O_3846,N_49934,N_49816);
or UO_3847 (O_3847,N_49971,N_49759);
nand UO_3848 (O_3848,N_49790,N_49868);
nand UO_3849 (O_3849,N_49881,N_49779);
and UO_3850 (O_3850,N_49897,N_49786);
nand UO_3851 (O_3851,N_49867,N_49829);
or UO_3852 (O_3852,N_49999,N_49860);
and UO_3853 (O_3853,N_49767,N_49807);
or UO_3854 (O_3854,N_49982,N_49977);
nor UO_3855 (O_3855,N_49870,N_49878);
xor UO_3856 (O_3856,N_49886,N_49950);
nor UO_3857 (O_3857,N_49966,N_49944);
or UO_3858 (O_3858,N_49992,N_49865);
nor UO_3859 (O_3859,N_49893,N_49824);
and UO_3860 (O_3860,N_49887,N_49929);
or UO_3861 (O_3861,N_49796,N_49825);
and UO_3862 (O_3862,N_49838,N_49931);
nor UO_3863 (O_3863,N_49986,N_49936);
nand UO_3864 (O_3864,N_49830,N_49801);
and UO_3865 (O_3865,N_49778,N_49773);
nand UO_3866 (O_3866,N_49837,N_49823);
or UO_3867 (O_3867,N_49989,N_49838);
and UO_3868 (O_3868,N_49832,N_49982);
nor UO_3869 (O_3869,N_49906,N_49931);
xor UO_3870 (O_3870,N_49775,N_49757);
nand UO_3871 (O_3871,N_49928,N_49956);
nand UO_3872 (O_3872,N_49940,N_49983);
or UO_3873 (O_3873,N_49836,N_49791);
or UO_3874 (O_3874,N_49845,N_49784);
xor UO_3875 (O_3875,N_49983,N_49967);
or UO_3876 (O_3876,N_49807,N_49907);
xnor UO_3877 (O_3877,N_49804,N_49762);
nand UO_3878 (O_3878,N_49968,N_49781);
nor UO_3879 (O_3879,N_49942,N_49960);
xnor UO_3880 (O_3880,N_49796,N_49773);
or UO_3881 (O_3881,N_49819,N_49968);
or UO_3882 (O_3882,N_49778,N_49951);
and UO_3883 (O_3883,N_49765,N_49787);
nor UO_3884 (O_3884,N_49977,N_49869);
xnor UO_3885 (O_3885,N_49941,N_49774);
nand UO_3886 (O_3886,N_49966,N_49851);
nand UO_3887 (O_3887,N_49929,N_49881);
or UO_3888 (O_3888,N_49763,N_49958);
or UO_3889 (O_3889,N_49782,N_49861);
and UO_3890 (O_3890,N_49758,N_49811);
xor UO_3891 (O_3891,N_49846,N_49953);
and UO_3892 (O_3892,N_49926,N_49837);
and UO_3893 (O_3893,N_49880,N_49922);
or UO_3894 (O_3894,N_49866,N_49876);
or UO_3895 (O_3895,N_49952,N_49821);
or UO_3896 (O_3896,N_49936,N_49858);
nand UO_3897 (O_3897,N_49979,N_49948);
or UO_3898 (O_3898,N_49936,N_49852);
and UO_3899 (O_3899,N_49801,N_49863);
or UO_3900 (O_3900,N_49770,N_49889);
nand UO_3901 (O_3901,N_49922,N_49779);
and UO_3902 (O_3902,N_49965,N_49820);
xnor UO_3903 (O_3903,N_49768,N_49790);
and UO_3904 (O_3904,N_49818,N_49877);
xor UO_3905 (O_3905,N_49938,N_49906);
nor UO_3906 (O_3906,N_49799,N_49968);
xor UO_3907 (O_3907,N_49766,N_49985);
or UO_3908 (O_3908,N_49950,N_49794);
nand UO_3909 (O_3909,N_49869,N_49835);
or UO_3910 (O_3910,N_49923,N_49856);
and UO_3911 (O_3911,N_49928,N_49984);
xnor UO_3912 (O_3912,N_49823,N_49942);
nand UO_3913 (O_3913,N_49811,N_49855);
nor UO_3914 (O_3914,N_49851,N_49968);
nor UO_3915 (O_3915,N_49950,N_49762);
nor UO_3916 (O_3916,N_49766,N_49809);
nand UO_3917 (O_3917,N_49883,N_49771);
or UO_3918 (O_3918,N_49916,N_49834);
nand UO_3919 (O_3919,N_49917,N_49935);
or UO_3920 (O_3920,N_49922,N_49867);
and UO_3921 (O_3921,N_49773,N_49993);
nand UO_3922 (O_3922,N_49813,N_49768);
nand UO_3923 (O_3923,N_49904,N_49797);
or UO_3924 (O_3924,N_49961,N_49915);
nand UO_3925 (O_3925,N_49880,N_49989);
nand UO_3926 (O_3926,N_49792,N_49781);
or UO_3927 (O_3927,N_49769,N_49958);
xor UO_3928 (O_3928,N_49995,N_49761);
xor UO_3929 (O_3929,N_49881,N_49896);
nand UO_3930 (O_3930,N_49884,N_49781);
or UO_3931 (O_3931,N_49953,N_49942);
nor UO_3932 (O_3932,N_49902,N_49994);
nor UO_3933 (O_3933,N_49966,N_49995);
nor UO_3934 (O_3934,N_49980,N_49944);
or UO_3935 (O_3935,N_49830,N_49952);
nand UO_3936 (O_3936,N_49867,N_49869);
or UO_3937 (O_3937,N_49776,N_49976);
nor UO_3938 (O_3938,N_49929,N_49864);
and UO_3939 (O_3939,N_49880,N_49759);
nor UO_3940 (O_3940,N_49914,N_49825);
and UO_3941 (O_3941,N_49830,N_49756);
xor UO_3942 (O_3942,N_49961,N_49877);
nor UO_3943 (O_3943,N_49987,N_49902);
nor UO_3944 (O_3944,N_49839,N_49890);
xor UO_3945 (O_3945,N_49759,N_49940);
nor UO_3946 (O_3946,N_49769,N_49753);
nor UO_3947 (O_3947,N_49772,N_49997);
or UO_3948 (O_3948,N_49935,N_49947);
nand UO_3949 (O_3949,N_49812,N_49867);
nand UO_3950 (O_3950,N_49880,N_49935);
nor UO_3951 (O_3951,N_49900,N_49768);
and UO_3952 (O_3952,N_49922,N_49910);
nand UO_3953 (O_3953,N_49843,N_49825);
nand UO_3954 (O_3954,N_49923,N_49809);
and UO_3955 (O_3955,N_49806,N_49939);
xor UO_3956 (O_3956,N_49814,N_49961);
xor UO_3957 (O_3957,N_49790,N_49928);
or UO_3958 (O_3958,N_49907,N_49771);
nor UO_3959 (O_3959,N_49985,N_49779);
nand UO_3960 (O_3960,N_49863,N_49806);
xnor UO_3961 (O_3961,N_49853,N_49866);
and UO_3962 (O_3962,N_49764,N_49887);
xnor UO_3963 (O_3963,N_49829,N_49971);
and UO_3964 (O_3964,N_49898,N_49978);
nand UO_3965 (O_3965,N_49877,N_49998);
nand UO_3966 (O_3966,N_49933,N_49936);
and UO_3967 (O_3967,N_49918,N_49865);
xor UO_3968 (O_3968,N_49777,N_49965);
xor UO_3969 (O_3969,N_49803,N_49825);
xnor UO_3970 (O_3970,N_49856,N_49983);
nand UO_3971 (O_3971,N_49903,N_49758);
nor UO_3972 (O_3972,N_49971,N_49809);
nor UO_3973 (O_3973,N_49912,N_49952);
nand UO_3974 (O_3974,N_49846,N_49870);
nand UO_3975 (O_3975,N_49974,N_49906);
nor UO_3976 (O_3976,N_49993,N_49990);
nor UO_3977 (O_3977,N_49792,N_49926);
and UO_3978 (O_3978,N_49897,N_49801);
or UO_3979 (O_3979,N_49775,N_49885);
nor UO_3980 (O_3980,N_49866,N_49827);
nor UO_3981 (O_3981,N_49813,N_49962);
nor UO_3982 (O_3982,N_49890,N_49778);
nor UO_3983 (O_3983,N_49968,N_49815);
or UO_3984 (O_3984,N_49982,N_49817);
xor UO_3985 (O_3985,N_49992,N_49806);
nor UO_3986 (O_3986,N_49864,N_49883);
and UO_3987 (O_3987,N_49891,N_49914);
or UO_3988 (O_3988,N_49935,N_49807);
nand UO_3989 (O_3989,N_49842,N_49784);
nor UO_3990 (O_3990,N_49999,N_49781);
nor UO_3991 (O_3991,N_49934,N_49974);
xnor UO_3992 (O_3992,N_49996,N_49771);
nor UO_3993 (O_3993,N_49888,N_49920);
nor UO_3994 (O_3994,N_49899,N_49950);
nor UO_3995 (O_3995,N_49824,N_49888);
nor UO_3996 (O_3996,N_49845,N_49911);
and UO_3997 (O_3997,N_49805,N_49815);
xor UO_3998 (O_3998,N_49899,N_49799);
nand UO_3999 (O_3999,N_49904,N_49798);
or UO_4000 (O_4000,N_49776,N_49802);
nand UO_4001 (O_4001,N_49944,N_49906);
xnor UO_4002 (O_4002,N_49907,N_49779);
nand UO_4003 (O_4003,N_49896,N_49956);
nor UO_4004 (O_4004,N_49793,N_49986);
and UO_4005 (O_4005,N_49815,N_49870);
nand UO_4006 (O_4006,N_49890,N_49955);
xor UO_4007 (O_4007,N_49873,N_49981);
and UO_4008 (O_4008,N_49816,N_49847);
xnor UO_4009 (O_4009,N_49780,N_49884);
nor UO_4010 (O_4010,N_49993,N_49816);
xnor UO_4011 (O_4011,N_49967,N_49782);
nand UO_4012 (O_4012,N_49965,N_49761);
xor UO_4013 (O_4013,N_49863,N_49942);
nor UO_4014 (O_4014,N_49876,N_49802);
xor UO_4015 (O_4015,N_49980,N_49848);
or UO_4016 (O_4016,N_49859,N_49788);
nand UO_4017 (O_4017,N_49940,N_49944);
nor UO_4018 (O_4018,N_49914,N_49772);
xor UO_4019 (O_4019,N_49778,N_49987);
nand UO_4020 (O_4020,N_49911,N_49990);
nor UO_4021 (O_4021,N_49929,N_49976);
nor UO_4022 (O_4022,N_49891,N_49931);
or UO_4023 (O_4023,N_49874,N_49783);
nand UO_4024 (O_4024,N_49916,N_49987);
nor UO_4025 (O_4025,N_49856,N_49754);
or UO_4026 (O_4026,N_49865,N_49830);
or UO_4027 (O_4027,N_49983,N_49872);
nand UO_4028 (O_4028,N_49770,N_49979);
or UO_4029 (O_4029,N_49847,N_49825);
xor UO_4030 (O_4030,N_49779,N_49897);
nand UO_4031 (O_4031,N_49847,N_49909);
and UO_4032 (O_4032,N_49808,N_49846);
xor UO_4033 (O_4033,N_49863,N_49814);
and UO_4034 (O_4034,N_49937,N_49978);
nand UO_4035 (O_4035,N_49788,N_49979);
xnor UO_4036 (O_4036,N_49980,N_49947);
nor UO_4037 (O_4037,N_49923,N_49833);
nor UO_4038 (O_4038,N_49786,N_49807);
nand UO_4039 (O_4039,N_49832,N_49941);
and UO_4040 (O_4040,N_49895,N_49961);
and UO_4041 (O_4041,N_49960,N_49974);
and UO_4042 (O_4042,N_49990,N_49865);
xnor UO_4043 (O_4043,N_49988,N_49976);
xnor UO_4044 (O_4044,N_49947,N_49786);
nand UO_4045 (O_4045,N_49819,N_49920);
xor UO_4046 (O_4046,N_49917,N_49908);
nand UO_4047 (O_4047,N_49759,N_49979);
nand UO_4048 (O_4048,N_49751,N_49910);
nand UO_4049 (O_4049,N_49837,N_49942);
and UO_4050 (O_4050,N_49766,N_49757);
nand UO_4051 (O_4051,N_49760,N_49761);
nor UO_4052 (O_4052,N_49913,N_49961);
nor UO_4053 (O_4053,N_49879,N_49958);
nand UO_4054 (O_4054,N_49810,N_49795);
xor UO_4055 (O_4055,N_49753,N_49878);
nand UO_4056 (O_4056,N_49930,N_49962);
nand UO_4057 (O_4057,N_49894,N_49832);
and UO_4058 (O_4058,N_49936,N_49951);
xor UO_4059 (O_4059,N_49959,N_49832);
xor UO_4060 (O_4060,N_49983,N_49876);
and UO_4061 (O_4061,N_49898,N_49852);
nor UO_4062 (O_4062,N_49800,N_49889);
nor UO_4063 (O_4063,N_49988,N_49886);
nor UO_4064 (O_4064,N_49790,N_49828);
xor UO_4065 (O_4065,N_49854,N_49961);
nor UO_4066 (O_4066,N_49766,N_49816);
or UO_4067 (O_4067,N_49805,N_49795);
and UO_4068 (O_4068,N_49779,N_49936);
and UO_4069 (O_4069,N_49846,N_49774);
nand UO_4070 (O_4070,N_49893,N_49869);
xnor UO_4071 (O_4071,N_49863,N_49809);
and UO_4072 (O_4072,N_49838,N_49866);
nor UO_4073 (O_4073,N_49895,N_49969);
and UO_4074 (O_4074,N_49774,N_49951);
nor UO_4075 (O_4075,N_49931,N_49975);
nand UO_4076 (O_4076,N_49932,N_49969);
nor UO_4077 (O_4077,N_49789,N_49946);
nor UO_4078 (O_4078,N_49977,N_49909);
or UO_4079 (O_4079,N_49908,N_49856);
or UO_4080 (O_4080,N_49918,N_49821);
nor UO_4081 (O_4081,N_49964,N_49927);
nor UO_4082 (O_4082,N_49965,N_49974);
and UO_4083 (O_4083,N_49903,N_49980);
and UO_4084 (O_4084,N_49965,N_49892);
or UO_4085 (O_4085,N_49825,N_49839);
xnor UO_4086 (O_4086,N_49854,N_49877);
xor UO_4087 (O_4087,N_49839,N_49795);
xor UO_4088 (O_4088,N_49793,N_49930);
or UO_4089 (O_4089,N_49989,N_49894);
xor UO_4090 (O_4090,N_49902,N_49829);
nor UO_4091 (O_4091,N_49869,N_49822);
nand UO_4092 (O_4092,N_49858,N_49978);
or UO_4093 (O_4093,N_49773,N_49762);
or UO_4094 (O_4094,N_49841,N_49817);
xnor UO_4095 (O_4095,N_49829,N_49788);
nand UO_4096 (O_4096,N_49818,N_49859);
nor UO_4097 (O_4097,N_49895,N_49794);
nand UO_4098 (O_4098,N_49850,N_49817);
or UO_4099 (O_4099,N_49833,N_49854);
nor UO_4100 (O_4100,N_49994,N_49934);
and UO_4101 (O_4101,N_49849,N_49973);
or UO_4102 (O_4102,N_49933,N_49953);
xnor UO_4103 (O_4103,N_49822,N_49794);
nand UO_4104 (O_4104,N_49962,N_49890);
xnor UO_4105 (O_4105,N_49977,N_49759);
and UO_4106 (O_4106,N_49871,N_49987);
nor UO_4107 (O_4107,N_49971,N_49760);
or UO_4108 (O_4108,N_49778,N_49750);
xor UO_4109 (O_4109,N_49907,N_49816);
xnor UO_4110 (O_4110,N_49864,N_49858);
nor UO_4111 (O_4111,N_49771,N_49787);
nor UO_4112 (O_4112,N_49892,N_49845);
nor UO_4113 (O_4113,N_49824,N_49975);
and UO_4114 (O_4114,N_49991,N_49845);
xnor UO_4115 (O_4115,N_49793,N_49881);
and UO_4116 (O_4116,N_49811,N_49812);
nand UO_4117 (O_4117,N_49856,N_49831);
xor UO_4118 (O_4118,N_49858,N_49995);
or UO_4119 (O_4119,N_49810,N_49918);
xor UO_4120 (O_4120,N_49807,N_49894);
xor UO_4121 (O_4121,N_49965,N_49883);
and UO_4122 (O_4122,N_49979,N_49871);
nor UO_4123 (O_4123,N_49876,N_49764);
nor UO_4124 (O_4124,N_49828,N_49947);
nand UO_4125 (O_4125,N_49975,N_49920);
nor UO_4126 (O_4126,N_49798,N_49927);
xor UO_4127 (O_4127,N_49870,N_49851);
xor UO_4128 (O_4128,N_49917,N_49835);
and UO_4129 (O_4129,N_49791,N_49845);
or UO_4130 (O_4130,N_49838,N_49780);
and UO_4131 (O_4131,N_49775,N_49923);
nand UO_4132 (O_4132,N_49859,N_49857);
and UO_4133 (O_4133,N_49832,N_49873);
nand UO_4134 (O_4134,N_49836,N_49952);
nand UO_4135 (O_4135,N_49773,N_49772);
nor UO_4136 (O_4136,N_49848,N_49933);
nand UO_4137 (O_4137,N_49817,N_49753);
nor UO_4138 (O_4138,N_49961,N_49874);
or UO_4139 (O_4139,N_49839,N_49777);
and UO_4140 (O_4140,N_49966,N_49998);
nor UO_4141 (O_4141,N_49859,N_49774);
or UO_4142 (O_4142,N_49962,N_49968);
nand UO_4143 (O_4143,N_49919,N_49778);
nand UO_4144 (O_4144,N_49853,N_49994);
nand UO_4145 (O_4145,N_49920,N_49904);
or UO_4146 (O_4146,N_49963,N_49853);
nand UO_4147 (O_4147,N_49990,N_49850);
and UO_4148 (O_4148,N_49934,N_49822);
and UO_4149 (O_4149,N_49946,N_49770);
nand UO_4150 (O_4150,N_49926,N_49814);
xnor UO_4151 (O_4151,N_49965,N_49887);
or UO_4152 (O_4152,N_49766,N_49959);
or UO_4153 (O_4153,N_49824,N_49810);
and UO_4154 (O_4154,N_49879,N_49941);
nor UO_4155 (O_4155,N_49785,N_49864);
xor UO_4156 (O_4156,N_49929,N_49811);
or UO_4157 (O_4157,N_49780,N_49994);
nand UO_4158 (O_4158,N_49925,N_49753);
nand UO_4159 (O_4159,N_49833,N_49933);
or UO_4160 (O_4160,N_49816,N_49751);
or UO_4161 (O_4161,N_49828,N_49957);
nand UO_4162 (O_4162,N_49998,N_49893);
xor UO_4163 (O_4163,N_49887,N_49810);
nand UO_4164 (O_4164,N_49979,N_49803);
nand UO_4165 (O_4165,N_49870,N_49919);
xor UO_4166 (O_4166,N_49833,N_49895);
or UO_4167 (O_4167,N_49767,N_49915);
nand UO_4168 (O_4168,N_49861,N_49852);
xor UO_4169 (O_4169,N_49916,N_49930);
nor UO_4170 (O_4170,N_49774,N_49786);
or UO_4171 (O_4171,N_49817,N_49900);
or UO_4172 (O_4172,N_49801,N_49943);
nand UO_4173 (O_4173,N_49847,N_49785);
and UO_4174 (O_4174,N_49803,N_49750);
nor UO_4175 (O_4175,N_49906,N_49883);
and UO_4176 (O_4176,N_49918,N_49997);
nand UO_4177 (O_4177,N_49991,N_49982);
nor UO_4178 (O_4178,N_49755,N_49797);
or UO_4179 (O_4179,N_49763,N_49849);
nand UO_4180 (O_4180,N_49911,N_49750);
nand UO_4181 (O_4181,N_49968,N_49766);
or UO_4182 (O_4182,N_49921,N_49837);
or UO_4183 (O_4183,N_49920,N_49922);
nand UO_4184 (O_4184,N_49831,N_49950);
or UO_4185 (O_4185,N_49907,N_49859);
nor UO_4186 (O_4186,N_49926,N_49900);
nand UO_4187 (O_4187,N_49908,N_49865);
nor UO_4188 (O_4188,N_49890,N_49804);
nor UO_4189 (O_4189,N_49793,N_49755);
nor UO_4190 (O_4190,N_49905,N_49858);
xor UO_4191 (O_4191,N_49848,N_49808);
xor UO_4192 (O_4192,N_49940,N_49816);
nor UO_4193 (O_4193,N_49771,N_49962);
and UO_4194 (O_4194,N_49803,N_49794);
xor UO_4195 (O_4195,N_49985,N_49750);
nor UO_4196 (O_4196,N_49809,N_49859);
nor UO_4197 (O_4197,N_49979,N_49987);
or UO_4198 (O_4198,N_49855,N_49967);
or UO_4199 (O_4199,N_49928,N_49926);
nor UO_4200 (O_4200,N_49864,N_49848);
nand UO_4201 (O_4201,N_49913,N_49812);
and UO_4202 (O_4202,N_49875,N_49908);
xnor UO_4203 (O_4203,N_49928,N_49777);
nor UO_4204 (O_4204,N_49876,N_49995);
or UO_4205 (O_4205,N_49893,N_49986);
nor UO_4206 (O_4206,N_49997,N_49759);
xnor UO_4207 (O_4207,N_49994,N_49953);
and UO_4208 (O_4208,N_49948,N_49917);
or UO_4209 (O_4209,N_49809,N_49849);
and UO_4210 (O_4210,N_49969,N_49941);
and UO_4211 (O_4211,N_49766,N_49866);
xor UO_4212 (O_4212,N_49752,N_49936);
or UO_4213 (O_4213,N_49814,N_49884);
and UO_4214 (O_4214,N_49917,N_49888);
and UO_4215 (O_4215,N_49839,N_49779);
or UO_4216 (O_4216,N_49889,N_49969);
xor UO_4217 (O_4217,N_49894,N_49833);
and UO_4218 (O_4218,N_49883,N_49849);
or UO_4219 (O_4219,N_49759,N_49921);
or UO_4220 (O_4220,N_49976,N_49906);
and UO_4221 (O_4221,N_49913,N_49845);
nor UO_4222 (O_4222,N_49786,N_49891);
nand UO_4223 (O_4223,N_49822,N_49881);
and UO_4224 (O_4224,N_49971,N_49825);
xor UO_4225 (O_4225,N_49921,N_49816);
xnor UO_4226 (O_4226,N_49844,N_49872);
nand UO_4227 (O_4227,N_49946,N_49756);
nand UO_4228 (O_4228,N_49995,N_49817);
nor UO_4229 (O_4229,N_49967,N_49836);
nor UO_4230 (O_4230,N_49916,N_49896);
nor UO_4231 (O_4231,N_49907,N_49874);
nor UO_4232 (O_4232,N_49834,N_49892);
xnor UO_4233 (O_4233,N_49864,N_49898);
xnor UO_4234 (O_4234,N_49981,N_49751);
or UO_4235 (O_4235,N_49876,N_49977);
nor UO_4236 (O_4236,N_49956,N_49773);
and UO_4237 (O_4237,N_49895,N_49838);
and UO_4238 (O_4238,N_49928,N_49844);
or UO_4239 (O_4239,N_49785,N_49908);
or UO_4240 (O_4240,N_49813,N_49774);
or UO_4241 (O_4241,N_49911,N_49811);
and UO_4242 (O_4242,N_49964,N_49752);
or UO_4243 (O_4243,N_49788,N_49890);
and UO_4244 (O_4244,N_49805,N_49866);
xor UO_4245 (O_4245,N_49787,N_49804);
nand UO_4246 (O_4246,N_49935,N_49865);
and UO_4247 (O_4247,N_49752,N_49853);
nor UO_4248 (O_4248,N_49930,N_49754);
and UO_4249 (O_4249,N_49877,N_49952);
nor UO_4250 (O_4250,N_49766,N_49860);
or UO_4251 (O_4251,N_49877,N_49853);
or UO_4252 (O_4252,N_49895,N_49990);
xnor UO_4253 (O_4253,N_49931,N_49781);
xor UO_4254 (O_4254,N_49835,N_49829);
or UO_4255 (O_4255,N_49759,N_49751);
nand UO_4256 (O_4256,N_49759,N_49904);
and UO_4257 (O_4257,N_49766,N_49758);
nand UO_4258 (O_4258,N_49757,N_49787);
or UO_4259 (O_4259,N_49863,N_49899);
xnor UO_4260 (O_4260,N_49826,N_49844);
nor UO_4261 (O_4261,N_49995,N_49973);
and UO_4262 (O_4262,N_49907,N_49791);
nor UO_4263 (O_4263,N_49886,N_49893);
nand UO_4264 (O_4264,N_49954,N_49867);
nor UO_4265 (O_4265,N_49808,N_49773);
or UO_4266 (O_4266,N_49993,N_49809);
xnor UO_4267 (O_4267,N_49958,N_49812);
nor UO_4268 (O_4268,N_49911,N_49906);
xnor UO_4269 (O_4269,N_49927,N_49818);
and UO_4270 (O_4270,N_49833,N_49918);
and UO_4271 (O_4271,N_49985,N_49864);
nor UO_4272 (O_4272,N_49904,N_49834);
or UO_4273 (O_4273,N_49835,N_49858);
nor UO_4274 (O_4274,N_49964,N_49769);
nand UO_4275 (O_4275,N_49893,N_49975);
nand UO_4276 (O_4276,N_49948,N_49800);
nand UO_4277 (O_4277,N_49865,N_49981);
and UO_4278 (O_4278,N_49805,N_49849);
nand UO_4279 (O_4279,N_49831,N_49822);
xnor UO_4280 (O_4280,N_49880,N_49827);
xor UO_4281 (O_4281,N_49978,N_49846);
nor UO_4282 (O_4282,N_49966,N_49878);
nor UO_4283 (O_4283,N_49900,N_49973);
or UO_4284 (O_4284,N_49798,N_49781);
nand UO_4285 (O_4285,N_49976,N_49877);
xor UO_4286 (O_4286,N_49796,N_49830);
and UO_4287 (O_4287,N_49784,N_49807);
xor UO_4288 (O_4288,N_49838,N_49767);
xnor UO_4289 (O_4289,N_49956,N_49987);
nand UO_4290 (O_4290,N_49813,N_49838);
or UO_4291 (O_4291,N_49797,N_49902);
nor UO_4292 (O_4292,N_49911,N_49849);
nor UO_4293 (O_4293,N_49852,N_49910);
xnor UO_4294 (O_4294,N_49986,N_49791);
nand UO_4295 (O_4295,N_49776,N_49922);
nand UO_4296 (O_4296,N_49897,N_49889);
nand UO_4297 (O_4297,N_49937,N_49784);
or UO_4298 (O_4298,N_49917,N_49878);
nor UO_4299 (O_4299,N_49756,N_49813);
nor UO_4300 (O_4300,N_49810,N_49886);
or UO_4301 (O_4301,N_49966,N_49993);
nand UO_4302 (O_4302,N_49934,N_49799);
nand UO_4303 (O_4303,N_49953,N_49889);
and UO_4304 (O_4304,N_49763,N_49862);
nor UO_4305 (O_4305,N_49997,N_49757);
nand UO_4306 (O_4306,N_49916,N_49855);
or UO_4307 (O_4307,N_49759,N_49907);
nand UO_4308 (O_4308,N_49957,N_49971);
nand UO_4309 (O_4309,N_49781,N_49976);
or UO_4310 (O_4310,N_49869,N_49907);
and UO_4311 (O_4311,N_49945,N_49965);
nand UO_4312 (O_4312,N_49851,N_49819);
nor UO_4313 (O_4313,N_49842,N_49876);
nor UO_4314 (O_4314,N_49903,N_49792);
nor UO_4315 (O_4315,N_49872,N_49752);
and UO_4316 (O_4316,N_49946,N_49823);
xor UO_4317 (O_4317,N_49975,N_49829);
and UO_4318 (O_4318,N_49982,N_49934);
and UO_4319 (O_4319,N_49791,N_49807);
nor UO_4320 (O_4320,N_49806,N_49883);
and UO_4321 (O_4321,N_49967,N_49816);
or UO_4322 (O_4322,N_49884,N_49849);
and UO_4323 (O_4323,N_49943,N_49876);
nand UO_4324 (O_4324,N_49947,N_49824);
nor UO_4325 (O_4325,N_49833,N_49907);
nand UO_4326 (O_4326,N_49838,N_49754);
nor UO_4327 (O_4327,N_49929,N_49819);
and UO_4328 (O_4328,N_49954,N_49947);
nor UO_4329 (O_4329,N_49759,N_49935);
or UO_4330 (O_4330,N_49841,N_49995);
xor UO_4331 (O_4331,N_49812,N_49762);
or UO_4332 (O_4332,N_49813,N_49875);
xnor UO_4333 (O_4333,N_49783,N_49756);
nor UO_4334 (O_4334,N_49820,N_49927);
and UO_4335 (O_4335,N_49771,N_49775);
nor UO_4336 (O_4336,N_49915,N_49909);
xnor UO_4337 (O_4337,N_49763,N_49775);
and UO_4338 (O_4338,N_49861,N_49807);
or UO_4339 (O_4339,N_49941,N_49847);
and UO_4340 (O_4340,N_49900,N_49769);
nor UO_4341 (O_4341,N_49914,N_49810);
and UO_4342 (O_4342,N_49889,N_49761);
nor UO_4343 (O_4343,N_49962,N_49955);
xnor UO_4344 (O_4344,N_49961,N_49887);
and UO_4345 (O_4345,N_49752,N_49943);
xor UO_4346 (O_4346,N_49931,N_49835);
and UO_4347 (O_4347,N_49984,N_49987);
or UO_4348 (O_4348,N_49841,N_49842);
and UO_4349 (O_4349,N_49986,N_49850);
nor UO_4350 (O_4350,N_49925,N_49792);
or UO_4351 (O_4351,N_49787,N_49997);
nand UO_4352 (O_4352,N_49960,N_49822);
or UO_4353 (O_4353,N_49787,N_49940);
nand UO_4354 (O_4354,N_49877,N_49878);
nand UO_4355 (O_4355,N_49839,N_49818);
nand UO_4356 (O_4356,N_49811,N_49875);
nand UO_4357 (O_4357,N_49825,N_49795);
or UO_4358 (O_4358,N_49827,N_49754);
or UO_4359 (O_4359,N_49837,N_49800);
nand UO_4360 (O_4360,N_49968,N_49833);
or UO_4361 (O_4361,N_49766,N_49781);
nor UO_4362 (O_4362,N_49942,N_49867);
nand UO_4363 (O_4363,N_49784,N_49804);
or UO_4364 (O_4364,N_49811,N_49788);
nand UO_4365 (O_4365,N_49935,N_49973);
xor UO_4366 (O_4366,N_49807,N_49992);
nand UO_4367 (O_4367,N_49845,N_49756);
nor UO_4368 (O_4368,N_49898,N_49794);
xor UO_4369 (O_4369,N_49907,N_49875);
nand UO_4370 (O_4370,N_49890,N_49980);
or UO_4371 (O_4371,N_49801,N_49970);
and UO_4372 (O_4372,N_49923,N_49894);
or UO_4373 (O_4373,N_49889,N_49961);
or UO_4374 (O_4374,N_49905,N_49989);
and UO_4375 (O_4375,N_49992,N_49883);
xnor UO_4376 (O_4376,N_49950,N_49948);
nand UO_4377 (O_4377,N_49957,N_49820);
or UO_4378 (O_4378,N_49808,N_49794);
and UO_4379 (O_4379,N_49927,N_49751);
xor UO_4380 (O_4380,N_49949,N_49994);
nor UO_4381 (O_4381,N_49823,N_49786);
and UO_4382 (O_4382,N_49823,N_49897);
nor UO_4383 (O_4383,N_49898,N_49756);
and UO_4384 (O_4384,N_49939,N_49881);
or UO_4385 (O_4385,N_49959,N_49808);
or UO_4386 (O_4386,N_49937,N_49873);
or UO_4387 (O_4387,N_49866,N_49897);
and UO_4388 (O_4388,N_49848,N_49884);
or UO_4389 (O_4389,N_49852,N_49830);
xor UO_4390 (O_4390,N_49808,N_49779);
nor UO_4391 (O_4391,N_49982,N_49873);
or UO_4392 (O_4392,N_49751,N_49810);
xnor UO_4393 (O_4393,N_49994,N_49836);
and UO_4394 (O_4394,N_49878,N_49891);
nand UO_4395 (O_4395,N_49985,N_49891);
xnor UO_4396 (O_4396,N_49948,N_49876);
nor UO_4397 (O_4397,N_49843,N_49984);
and UO_4398 (O_4398,N_49757,N_49886);
and UO_4399 (O_4399,N_49994,N_49941);
nor UO_4400 (O_4400,N_49952,N_49897);
nand UO_4401 (O_4401,N_49930,N_49762);
or UO_4402 (O_4402,N_49797,N_49863);
or UO_4403 (O_4403,N_49889,N_49756);
or UO_4404 (O_4404,N_49832,N_49802);
xnor UO_4405 (O_4405,N_49880,N_49851);
nand UO_4406 (O_4406,N_49967,N_49976);
nor UO_4407 (O_4407,N_49759,N_49827);
nand UO_4408 (O_4408,N_49987,N_49922);
nand UO_4409 (O_4409,N_49885,N_49796);
nand UO_4410 (O_4410,N_49905,N_49914);
and UO_4411 (O_4411,N_49828,N_49893);
or UO_4412 (O_4412,N_49972,N_49788);
xnor UO_4413 (O_4413,N_49893,N_49902);
nor UO_4414 (O_4414,N_49773,N_49901);
or UO_4415 (O_4415,N_49978,N_49759);
xor UO_4416 (O_4416,N_49782,N_49965);
xor UO_4417 (O_4417,N_49862,N_49918);
or UO_4418 (O_4418,N_49967,N_49826);
nor UO_4419 (O_4419,N_49826,N_49883);
nor UO_4420 (O_4420,N_49942,N_49795);
xnor UO_4421 (O_4421,N_49860,N_49980);
nor UO_4422 (O_4422,N_49786,N_49995);
nor UO_4423 (O_4423,N_49911,N_49957);
or UO_4424 (O_4424,N_49835,N_49926);
and UO_4425 (O_4425,N_49752,N_49913);
xnor UO_4426 (O_4426,N_49924,N_49765);
nand UO_4427 (O_4427,N_49857,N_49901);
xnor UO_4428 (O_4428,N_49944,N_49888);
xor UO_4429 (O_4429,N_49816,N_49774);
and UO_4430 (O_4430,N_49764,N_49951);
nand UO_4431 (O_4431,N_49866,N_49975);
and UO_4432 (O_4432,N_49837,N_49918);
xnor UO_4433 (O_4433,N_49981,N_49909);
nand UO_4434 (O_4434,N_49785,N_49897);
nand UO_4435 (O_4435,N_49773,N_49920);
nor UO_4436 (O_4436,N_49906,N_49950);
nor UO_4437 (O_4437,N_49975,N_49787);
nand UO_4438 (O_4438,N_49754,N_49848);
or UO_4439 (O_4439,N_49955,N_49788);
and UO_4440 (O_4440,N_49899,N_49770);
and UO_4441 (O_4441,N_49879,N_49920);
nand UO_4442 (O_4442,N_49926,N_49993);
nor UO_4443 (O_4443,N_49910,N_49880);
nor UO_4444 (O_4444,N_49934,N_49923);
or UO_4445 (O_4445,N_49803,N_49789);
nand UO_4446 (O_4446,N_49821,N_49899);
xor UO_4447 (O_4447,N_49816,N_49825);
nand UO_4448 (O_4448,N_49811,N_49945);
nor UO_4449 (O_4449,N_49910,N_49812);
or UO_4450 (O_4450,N_49798,N_49848);
nand UO_4451 (O_4451,N_49784,N_49999);
or UO_4452 (O_4452,N_49832,N_49874);
and UO_4453 (O_4453,N_49778,N_49926);
nand UO_4454 (O_4454,N_49887,N_49803);
or UO_4455 (O_4455,N_49783,N_49913);
nand UO_4456 (O_4456,N_49940,N_49750);
nand UO_4457 (O_4457,N_49814,N_49931);
nor UO_4458 (O_4458,N_49860,N_49779);
or UO_4459 (O_4459,N_49824,N_49992);
nor UO_4460 (O_4460,N_49980,N_49776);
nor UO_4461 (O_4461,N_49792,N_49906);
and UO_4462 (O_4462,N_49750,N_49873);
and UO_4463 (O_4463,N_49835,N_49992);
or UO_4464 (O_4464,N_49830,N_49869);
nor UO_4465 (O_4465,N_49920,N_49851);
nand UO_4466 (O_4466,N_49980,N_49759);
xor UO_4467 (O_4467,N_49961,N_49851);
and UO_4468 (O_4468,N_49882,N_49998);
nand UO_4469 (O_4469,N_49871,N_49932);
nor UO_4470 (O_4470,N_49915,N_49879);
and UO_4471 (O_4471,N_49898,N_49991);
and UO_4472 (O_4472,N_49758,N_49878);
nor UO_4473 (O_4473,N_49864,N_49959);
or UO_4474 (O_4474,N_49908,N_49955);
xor UO_4475 (O_4475,N_49903,N_49924);
nand UO_4476 (O_4476,N_49943,N_49851);
nand UO_4477 (O_4477,N_49763,N_49902);
or UO_4478 (O_4478,N_49986,N_49953);
nand UO_4479 (O_4479,N_49926,N_49771);
xnor UO_4480 (O_4480,N_49906,N_49956);
or UO_4481 (O_4481,N_49912,N_49991);
or UO_4482 (O_4482,N_49760,N_49987);
xnor UO_4483 (O_4483,N_49911,N_49885);
or UO_4484 (O_4484,N_49894,N_49932);
or UO_4485 (O_4485,N_49789,N_49961);
or UO_4486 (O_4486,N_49909,N_49957);
xor UO_4487 (O_4487,N_49901,N_49994);
nor UO_4488 (O_4488,N_49910,N_49926);
and UO_4489 (O_4489,N_49787,N_49972);
xor UO_4490 (O_4490,N_49770,N_49877);
nand UO_4491 (O_4491,N_49931,N_49840);
nand UO_4492 (O_4492,N_49967,N_49773);
xnor UO_4493 (O_4493,N_49869,N_49948);
and UO_4494 (O_4494,N_49972,N_49994);
nand UO_4495 (O_4495,N_49893,N_49999);
nand UO_4496 (O_4496,N_49856,N_49803);
nor UO_4497 (O_4497,N_49891,N_49930);
and UO_4498 (O_4498,N_49760,N_49975);
or UO_4499 (O_4499,N_49810,N_49935);
or UO_4500 (O_4500,N_49912,N_49971);
xnor UO_4501 (O_4501,N_49791,N_49846);
nor UO_4502 (O_4502,N_49947,N_49916);
xnor UO_4503 (O_4503,N_49852,N_49771);
nand UO_4504 (O_4504,N_49866,N_49783);
or UO_4505 (O_4505,N_49848,N_49976);
and UO_4506 (O_4506,N_49899,N_49846);
or UO_4507 (O_4507,N_49998,N_49754);
nand UO_4508 (O_4508,N_49817,N_49952);
xnor UO_4509 (O_4509,N_49867,N_49859);
nor UO_4510 (O_4510,N_49769,N_49995);
nor UO_4511 (O_4511,N_49907,N_49871);
xor UO_4512 (O_4512,N_49783,N_49964);
nor UO_4513 (O_4513,N_49929,N_49934);
and UO_4514 (O_4514,N_49840,N_49980);
and UO_4515 (O_4515,N_49918,N_49936);
nand UO_4516 (O_4516,N_49843,N_49892);
and UO_4517 (O_4517,N_49961,N_49800);
nand UO_4518 (O_4518,N_49975,N_49839);
nor UO_4519 (O_4519,N_49827,N_49942);
xnor UO_4520 (O_4520,N_49928,N_49891);
and UO_4521 (O_4521,N_49824,N_49776);
and UO_4522 (O_4522,N_49881,N_49967);
or UO_4523 (O_4523,N_49830,N_49837);
and UO_4524 (O_4524,N_49911,N_49949);
nand UO_4525 (O_4525,N_49936,N_49950);
xnor UO_4526 (O_4526,N_49980,N_49940);
nand UO_4527 (O_4527,N_49953,N_49805);
xor UO_4528 (O_4528,N_49842,N_49806);
nor UO_4529 (O_4529,N_49838,N_49868);
nor UO_4530 (O_4530,N_49754,N_49794);
or UO_4531 (O_4531,N_49815,N_49849);
or UO_4532 (O_4532,N_49907,N_49752);
nand UO_4533 (O_4533,N_49778,N_49957);
nand UO_4534 (O_4534,N_49961,N_49838);
nor UO_4535 (O_4535,N_49765,N_49788);
nor UO_4536 (O_4536,N_49939,N_49931);
or UO_4537 (O_4537,N_49933,N_49871);
nor UO_4538 (O_4538,N_49763,N_49760);
xor UO_4539 (O_4539,N_49845,N_49894);
and UO_4540 (O_4540,N_49924,N_49842);
nand UO_4541 (O_4541,N_49785,N_49901);
and UO_4542 (O_4542,N_49879,N_49942);
xor UO_4543 (O_4543,N_49934,N_49850);
nor UO_4544 (O_4544,N_49869,N_49780);
and UO_4545 (O_4545,N_49853,N_49939);
nor UO_4546 (O_4546,N_49977,N_49976);
nor UO_4547 (O_4547,N_49848,N_49834);
nor UO_4548 (O_4548,N_49872,N_49849);
nor UO_4549 (O_4549,N_49941,N_49844);
nand UO_4550 (O_4550,N_49808,N_49818);
xnor UO_4551 (O_4551,N_49935,N_49997);
or UO_4552 (O_4552,N_49967,N_49904);
nand UO_4553 (O_4553,N_49979,N_49793);
nor UO_4554 (O_4554,N_49764,N_49895);
xor UO_4555 (O_4555,N_49754,N_49861);
and UO_4556 (O_4556,N_49759,N_49945);
and UO_4557 (O_4557,N_49773,N_49924);
and UO_4558 (O_4558,N_49766,N_49837);
nand UO_4559 (O_4559,N_49997,N_49957);
and UO_4560 (O_4560,N_49895,N_49759);
nor UO_4561 (O_4561,N_49989,N_49931);
xor UO_4562 (O_4562,N_49964,N_49985);
nor UO_4563 (O_4563,N_49988,N_49767);
and UO_4564 (O_4564,N_49942,N_49843);
nor UO_4565 (O_4565,N_49883,N_49822);
and UO_4566 (O_4566,N_49758,N_49914);
xnor UO_4567 (O_4567,N_49846,N_49830);
or UO_4568 (O_4568,N_49826,N_49811);
or UO_4569 (O_4569,N_49770,N_49947);
nor UO_4570 (O_4570,N_49915,N_49763);
nand UO_4571 (O_4571,N_49797,N_49964);
nand UO_4572 (O_4572,N_49829,N_49871);
and UO_4573 (O_4573,N_49793,N_49826);
or UO_4574 (O_4574,N_49790,N_49918);
or UO_4575 (O_4575,N_49844,N_49949);
xnor UO_4576 (O_4576,N_49983,N_49966);
nand UO_4577 (O_4577,N_49857,N_49982);
xnor UO_4578 (O_4578,N_49972,N_49750);
and UO_4579 (O_4579,N_49945,N_49869);
xnor UO_4580 (O_4580,N_49974,N_49857);
and UO_4581 (O_4581,N_49881,N_49974);
nand UO_4582 (O_4582,N_49938,N_49902);
and UO_4583 (O_4583,N_49751,N_49892);
and UO_4584 (O_4584,N_49770,N_49820);
nand UO_4585 (O_4585,N_49873,N_49931);
xor UO_4586 (O_4586,N_49984,N_49856);
nor UO_4587 (O_4587,N_49987,N_49784);
and UO_4588 (O_4588,N_49900,N_49894);
and UO_4589 (O_4589,N_49971,N_49838);
and UO_4590 (O_4590,N_49974,N_49764);
xor UO_4591 (O_4591,N_49989,N_49831);
nor UO_4592 (O_4592,N_49882,N_49861);
and UO_4593 (O_4593,N_49890,N_49985);
nor UO_4594 (O_4594,N_49887,N_49995);
or UO_4595 (O_4595,N_49882,N_49971);
and UO_4596 (O_4596,N_49986,N_49864);
or UO_4597 (O_4597,N_49891,N_49915);
or UO_4598 (O_4598,N_49997,N_49942);
and UO_4599 (O_4599,N_49878,N_49764);
xor UO_4600 (O_4600,N_49966,N_49957);
nand UO_4601 (O_4601,N_49954,N_49916);
nor UO_4602 (O_4602,N_49917,N_49765);
and UO_4603 (O_4603,N_49795,N_49763);
or UO_4604 (O_4604,N_49862,N_49790);
and UO_4605 (O_4605,N_49970,N_49826);
and UO_4606 (O_4606,N_49764,N_49796);
xor UO_4607 (O_4607,N_49897,N_49815);
nor UO_4608 (O_4608,N_49829,N_49915);
nand UO_4609 (O_4609,N_49891,N_49934);
or UO_4610 (O_4610,N_49843,N_49901);
nand UO_4611 (O_4611,N_49787,N_49761);
xnor UO_4612 (O_4612,N_49845,N_49878);
and UO_4613 (O_4613,N_49901,N_49911);
xnor UO_4614 (O_4614,N_49828,N_49973);
nand UO_4615 (O_4615,N_49790,N_49901);
or UO_4616 (O_4616,N_49795,N_49823);
nand UO_4617 (O_4617,N_49847,N_49838);
xnor UO_4618 (O_4618,N_49910,N_49930);
or UO_4619 (O_4619,N_49849,N_49869);
nand UO_4620 (O_4620,N_49989,N_49819);
nor UO_4621 (O_4621,N_49818,N_49921);
or UO_4622 (O_4622,N_49804,N_49806);
nand UO_4623 (O_4623,N_49861,N_49857);
nor UO_4624 (O_4624,N_49791,N_49883);
and UO_4625 (O_4625,N_49984,N_49939);
nor UO_4626 (O_4626,N_49904,N_49957);
and UO_4627 (O_4627,N_49879,N_49786);
nand UO_4628 (O_4628,N_49804,N_49925);
and UO_4629 (O_4629,N_49971,N_49951);
nand UO_4630 (O_4630,N_49831,N_49803);
or UO_4631 (O_4631,N_49978,N_49788);
xnor UO_4632 (O_4632,N_49781,N_49821);
xor UO_4633 (O_4633,N_49935,N_49916);
nor UO_4634 (O_4634,N_49788,N_49806);
nand UO_4635 (O_4635,N_49991,N_49792);
or UO_4636 (O_4636,N_49912,N_49810);
and UO_4637 (O_4637,N_49750,N_49998);
nand UO_4638 (O_4638,N_49892,N_49996);
or UO_4639 (O_4639,N_49973,N_49764);
nand UO_4640 (O_4640,N_49757,N_49810);
and UO_4641 (O_4641,N_49868,N_49751);
xnor UO_4642 (O_4642,N_49877,N_49840);
nor UO_4643 (O_4643,N_49802,N_49820);
nor UO_4644 (O_4644,N_49850,N_49765);
nand UO_4645 (O_4645,N_49879,N_49875);
or UO_4646 (O_4646,N_49982,N_49776);
xnor UO_4647 (O_4647,N_49925,N_49852);
or UO_4648 (O_4648,N_49850,N_49792);
nand UO_4649 (O_4649,N_49986,N_49761);
xor UO_4650 (O_4650,N_49986,N_49902);
nor UO_4651 (O_4651,N_49876,N_49921);
or UO_4652 (O_4652,N_49819,N_49762);
nor UO_4653 (O_4653,N_49792,N_49816);
or UO_4654 (O_4654,N_49888,N_49775);
nor UO_4655 (O_4655,N_49821,N_49845);
nor UO_4656 (O_4656,N_49804,N_49809);
xnor UO_4657 (O_4657,N_49903,N_49805);
nor UO_4658 (O_4658,N_49886,N_49852);
nand UO_4659 (O_4659,N_49959,N_49880);
and UO_4660 (O_4660,N_49774,N_49887);
nand UO_4661 (O_4661,N_49980,N_49882);
and UO_4662 (O_4662,N_49912,N_49801);
or UO_4663 (O_4663,N_49831,N_49963);
xnor UO_4664 (O_4664,N_49949,N_49963);
or UO_4665 (O_4665,N_49993,N_49936);
or UO_4666 (O_4666,N_49913,N_49754);
nand UO_4667 (O_4667,N_49756,N_49942);
xnor UO_4668 (O_4668,N_49986,N_49808);
and UO_4669 (O_4669,N_49803,N_49880);
xor UO_4670 (O_4670,N_49986,N_49892);
nand UO_4671 (O_4671,N_49849,N_49877);
xor UO_4672 (O_4672,N_49896,N_49955);
nor UO_4673 (O_4673,N_49917,N_49978);
xor UO_4674 (O_4674,N_49885,N_49820);
nand UO_4675 (O_4675,N_49828,N_49904);
xnor UO_4676 (O_4676,N_49862,N_49872);
and UO_4677 (O_4677,N_49786,N_49924);
or UO_4678 (O_4678,N_49960,N_49751);
or UO_4679 (O_4679,N_49756,N_49951);
and UO_4680 (O_4680,N_49944,N_49845);
or UO_4681 (O_4681,N_49923,N_49770);
and UO_4682 (O_4682,N_49941,N_49806);
or UO_4683 (O_4683,N_49809,N_49875);
and UO_4684 (O_4684,N_49804,N_49798);
nand UO_4685 (O_4685,N_49933,N_49962);
nand UO_4686 (O_4686,N_49829,N_49889);
nor UO_4687 (O_4687,N_49856,N_49784);
nand UO_4688 (O_4688,N_49849,N_49983);
and UO_4689 (O_4689,N_49969,N_49754);
and UO_4690 (O_4690,N_49783,N_49858);
nand UO_4691 (O_4691,N_49793,N_49915);
xnor UO_4692 (O_4692,N_49842,N_49866);
nor UO_4693 (O_4693,N_49924,N_49799);
nand UO_4694 (O_4694,N_49761,N_49939);
nor UO_4695 (O_4695,N_49954,N_49821);
or UO_4696 (O_4696,N_49819,N_49802);
xor UO_4697 (O_4697,N_49918,N_49853);
and UO_4698 (O_4698,N_49808,N_49882);
and UO_4699 (O_4699,N_49850,N_49978);
and UO_4700 (O_4700,N_49932,N_49779);
and UO_4701 (O_4701,N_49786,N_49967);
nor UO_4702 (O_4702,N_49829,N_49838);
nand UO_4703 (O_4703,N_49954,N_49885);
xnor UO_4704 (O_4704,N_49786,N_49985);
nor UO_4705 (O_4705,N_49757,N_49893);
or UO_4706 (O_4706,N_49883,N_49913);
xor UO_4707 (O_4707,N_49812,N_49842);
nor UO_4708 (O_4708,N_49988,N_49941);
nor UO_4709 (O_4709,N_49784,N_49800);
and UO_4710 (O_4710,N_49970,N_49903);
nor UO_4711 (O_4711,N_49853,N_49817);
nand UO_4712 (O_4712,N_49989,N_49932);
and UO_4713 (O_4713,N_49833,N_49827);
nor UO_4714 (O_4714,N_49831,N_49959);
xor UO_4715 (O_4715,N_49923,N_49888);
xor UO_4716 (O_4716,N_49993,N_49833);
or UO_4717 (O_4717,N_49816,N_49833);
or UO_4718 (O_4718,N_49938,N_49850);
and UO_4719 (O_4719,N_49862,N_49889);
xnor UO_4720 (O_4720,N_49980,N_49974);
nor UO_4721 (O_4721,N_49785,N_49784);
nand UO_4722 (O_4722,N_49822,N_49826);
or UO_4723 (O_4723,N_49921,N_49865);
xor UO_4724 (O_4724,N_49886,N_49778);
and UO_4725 (O_4725,N_49959,N_49994);
or UO_4726 (O_4726,N_49922,N_49932);
and UO_4727 (O_4727,N_49813,N_49997);
or UO_4728 (O_4728,N_49794,N_49910);
nand UO_4729 (O_4729,N_49856,N_49974);
and UO_4730 (O_4730,N_49863,N_49988);
or UO_4731 (O_4731,N_49787,N_49986);
and UO_4732 (O_4732,N_49758,N_49814);
xor UO_4733 (O_4733,N_49861,N_49954);
or UO_4734 (O_4734,N_49936,N_49912);
xor UO_4735 (O_4735,N_49961,N_49960);
and UO_4736 (O_4736,N_49820,N_49925);
xor UO_4737 (O_4737,N_49813,N_49990);
nand UO_4738 (O_4738,N_49753,N_49868);
nand UO_4739 (O_4739,N_49783,N_49805);
and UO_4740 (O_4740,N_49858,N_49870);
or UO_4741 (O_4741,N_49794,N_49885);
and UO_4742 (O_4742,N_49935,N_49789);
or UO_4743 (O_4743,N_49799,N_49881);
nand UO_4744 (O_4744,N_49854,N_49925);
xor UO_4745 (O_4745,N_49942,N_49797);
and UO_4746 (O_4746,N_49956,N_49926);
nand UO_4747 (O_4747,N_49927,N_49773);
xor UO_4748 (O_4748,N_49802,N_49843);
xor UO_4749 (O_4749,N_49856,N_49782);
xor UO_4750 (O_4750,N_49787,N_49984);
or UO_4751 (O_4751,N_49916,N_49780);
nor UO_4752 (O_4752,N_49948,N_49918);
and UO_4753 (O_4753,N_49827,N_49954);
nor UO_4754 (O_4754,N_49891,N_49911);
nand UO_4755 (O_4755,N_49872,N_49790);
nand UO_4756 (O_4756,N_49952,N_49826);
xnor UO_4757 (O_4757,N_49853,N_49879);
nand UO_4758 (O_4758,N_49787,N_49796);
nor UO_4759 (O_4759,N_49950,N_49850);
nor UO_4760 (O_4760,N_49761,N_49821);
xor UO_4761 (O_4761,N_49840,N_49833);
and UO_4762 (O_4762,N_49832,N_49944);
or UO_4763 (O_4763,N_49823,N_49791);
and UO_4764 (O_4764,N_49894,N_49814);
and UO_4765 (O_4765,N_49979,N_49908);
nor UO_4766 (O_4766,N_49976,N_49952);
nand UO_4767 (O_4767,N_49856,N_49930);
xnor UO_4768 (O_4768,N_49845,N_49768);
and UO_4769 (O_4769,N_49937,N_49908);
or UO_4770 (O_4770,N_49897,N_49864);
nor UO_4771 (O_4771,N_49803,N_49788);
nor UO_4772 (O_4772,N_49902,N_49835);
or UO_4773 (O_4773,N_49876,N_49831);
and UO_4774 (O_4774,N_49874,N_49778);
nand UO_4775 (O_4775,N_49881,N_49872);
or UO_4776 (O_4776,N_49996,N_49985);
or UO_4777 (O_4777,N_49908,N_49825);
or UO_4778 (O_4778,N_49846,N_49927);
xnor UO_4779 (O_4779,N_49846,N_49850);
and UO_4780 (O_4780,N_49896,N_49823);
or UO_4781 (O_4781,N_49784,N_49915);
or UO_4782 (O_4782,N_49849,N_49779);
nand UO_4783 (O_4783,N_49993,N_49958);
nand UO_4784 (O_4784,N_49857,N_49893);
nor UO_4785 (O_4785,N_49931,N_49912);
or UO_4786 (O_4786,N_49830,N_49995);
nor UO_4787 (O_4787,N_49798,N_49950);
or UO_4788 (O_4788,N_49803,N_49793);
or UO_4789 (O_4789,N_49957,N_49865);
xor UO_4790 (O_4790,N_49851,N_49906);
and UO_4791 (O_4791,N_49909,N_49814);
nand UO_4792 (O_4792,N_49777,N_49859);
or UO_4793 (O_4793,N_49790,N_49769);
and UO_4794 (O_4794,N_49824,N_49876);
nor UO_4795 (O_4795,N_49915,N_49972);
nor UO_4796 (O_4796,N_49821,N_49860);
xnor UO_4797 (O_4797,N_49855,N_49972);
or UO_4798 (O_4798,N_49765,N_49896);
nor UO_4799 (O_4799,N_49801,N_49765);
nand UO_4800 (O_4800,N_49942,N_49981);
nor UO_4801 (O_4801,N_49783,N_49816);
and UO_4802 (O_4802,N_49880,N_49849);
or UO_4803 (O_4803,N_49890,N_49884);
nor UO_4804 (O_4804,N_49909,N_49771);
or UO_4805 (O_4805,N_49883,N_49855);
and UO_4806 (O_4806,N_49854,N_49809);
nor UO_4807 (O_4807,N_49845,N_49899);
or UO_4808 (O_4808,N_49835,N_49988);
nor UO_4809 (O_4809,N_49870,N_49828);
nor UO_4810 (O_4810,N_49880,N_49865);
and UO_4811 (O_4811,N_49767,N_49929);
xnor UO_4812 (O_4812,N_49928,N_49884);
nand UO_4813 (O_4813,N_49756,N_49966);
or UO_4814 (O_4814,N_49819,N_49970);
and UO_4815 (O_4815,N_49757,N_49874);
nand UO_4816 (O_4816,N_49927,N_49769);
or UO_4817 (O_4817,N_49807,N_49853);
nor UO_4818 (O_4818,N_49849,N_49837);
xnor UO_4819 (O_4819,N_49765,N_49856);
xor UO_4820 (O_4820,N_49801,N_49975);
nor UO_4821 (O_4821,N_49998,N_49977);
nand UO_4822 (O_4822,N_49952,N_49993);
or UO_4823 (O_4823,N_49804,N_49832);
or UO_4824 (O_4824,N_49758,N_49850);
xor UO_4825 (O_4825,N_49854,N_49947);
xor UO_4826 (O_4826,N_49939,N_49962);
and UO_4827 (O_4827,N_49805,N_49807);
nand UO_4828 (O_4828,N_49906,N_49942);
xor UO_4829 (O_4829,N_49916,N_49866);
xor UO_4830 (O_4830,N_49929,N_49776);
nor UO_4831 (O_4831,N_49845,N_49910);
xor UO_4832 (O_4832,N_49921,N_49898);
xnor UO_4833 (O_4833,N_49994,N_49922);
nand UO_4834 (O_4834,N_49881,N_49900);
nor UO_4835 (O_4835,N_49943,N_49867);
xnor UO_4836 (O_4836,N_49972,N_49828);
nor UO_4837 (O_4837,N_49869,N_49953);
xnor UO_4838 (O_4838,N_49925,N_49821);
xor UO_4839 (O_4839,N_49995,N_49981);
and UO_4840 (O_4840,N_49829,N_49927);
nand UO_4841 (O_4841,N_49801,N_49890);
or UO_4842 (O_4842,N_49840,N_49964);
or UO_4843 (O_4843,N_49848,N_49852);
xnor UO_4844 (O_4844,N_49827,N_49916);
nand UO_4845 (O_4845,N_49827,N_49983);
nand UO_4846 (O_4846,N_49970,N_49835);
nor UO_4847 (O_4847,N_49766,N_49850);
and UO_4848 (O_4848,N_49844,N_49943);
xnor UO_4849 (O_4849,N_49898,N_49894);
nor UO_4850 (O_4850,N_49788,N_49750);
and UO_4851 (O_4851,N_49886,N_49908);
xnor UO_4852 (O_4852,N_49919,N_49820);
nand UO_4853 (O_4853,N_49827,N_49836);
nor UO_4854 (O_4854,N_49966,N_49858);
nor UO_4855 (O_4855,N_49987,N_49935);
nand UO_4856 (O_4856,N_49833,N_49991);
or UO_4857 (O_4857,N_49944,N_49960);
nor UO_4858 (O_4858,N_49762,N_49841);
nor UO_4859 (O_4859,N_49981,N_49931);
nand UO_4860 (O_4860,N_49973,N_49923);
nand UO_4861 (O_4861,N_49836,N_49865);
nand UO_4862 (O_4862,N_49839,N_49774);
xor UO_4863 (O_4863,N_49983,N_49936);
nor UO_4864 (O_4864,N_49825,N_49787);
xnor UO_4865 (O_4865,N_49795,N_49968);
or UO_4866 (O_4866,N_49890,N_49911);
or UO_4867 (O_4867,N_49851,N_49773);
xor UO_4868 (O_4868,N_49976,N_49957);
nor UO_4869 (O_4869,N_49821,N_49798);
and UO_4870 (O_4870,N_49883,N_49907);
and UO_4871 (O_4871,N_49885,N_49755);
xnor UO_4872 (O_4872,N_49910,N_49896);
and UO_4873 (O_4873,N_49764,N_49783);
nand UO_4874 (O_4874,N_49833,N_49948);
or UO_4875 (O_4875,N_49984,N_49835);
and UO_4876 (O_4876,N_49953,N_49927);
nor UO_4877 (O_4877,N_49788,N_49786);
xor UO_4878 (O_4878,N_49756,N_49982);
or UO_4879 (O_4879,N_49895,N_49955);
and UO_4880 (O_4880,N_49833,N_49903);
or UO_4881 (O_4881,N_49853,N_49824);
or UO_4882 (O_4882,N_49806,N_49795);
nand UO_4883 (O_4883,N_49962,N_49767);
xnor UO_4884 (O_4884,N_49764,N_49995);
nor UO_4885 (O_4885,N_49788,N_49929);
xnor UO_4886 (O_4886,N_49829,N_49911);
or UO_4887 (O_4887,N_49976,N_49994);
and UO_4888 (O_4888,N_49878,N_49767);
or UO_4889 (O_4889,N_49753,N_49848);
xnor UO_4890 (O_4890,N_49905,N_49883);
or UO_4891 (O_4891,N_49986,N_49769);
and UO_4892 (O_4892,N_49972,N_49901);
xnor UO_4893 (O_4893,N_49910,N_49791);
nor UO_4894 (O_4894,N_49961,N_49908);
xor UO_4895 (O_4895,N_49879,N_49865);
nand UO_4896 (O_4896,N_49915,N_49951);
or UO_4897 (O_4897,N_49827,N_49768);
xnor UO_4898 (O_4898,N_49822,N_49860);
and UO_4899 (O_4899,N_49916,N_49862);
nand UO_4900 (O_4900,N_49752,N_49863);
or UO_4901 (O_4901,N_49767,N_49819);
and UO_4902 (O_4902,N_49907,N_49937);
or UO_4903 (O_4903,N_49867,N_49959);
xnor UO_4904 (O_4904,N_49843,N_49850);
xor UO_4905 (O_4905,N_49997,N_49820);
nor UO_4906 (O_4906,N_49937,N_49831);
xnor UO_4907 (O_4907,N_49932,N_49847);
nor UO_4908 (O_4908,N_49762,N_49927);
nand UO_4909 (O_4909,N_49958,N_49893);
xnor UO_4910 (O_4910,N_49766,N_49838);
nand UO_4911 (O_4911,N_49985,N_49922);
and UO_4912 (O_4912,N_49822,N_49770);
xor UO_4913 (O_4913,N_49784,N_49835);
and UO_4914 (O_4914,N_49852,N_49934);
and UO_4915 (O_4915,N_49924,N_49874);
or UO_4916 (O_4916,N_49880,N_49894);
and UO_4917 (O_4917,N_49857,N_49750);
nand UO_4918 (O_4918,N_49840,N_49849);
and UO_4919 (O_4919,N_49993,N_49986);
or UO_4920 (O_4920,N_49859,N_49838);
xor UO_4921 (O_4921,N_49765,N_49846);
or UO_4922 (O_4922,N_49826,N_49960);
xnor UO_4923 (O_4923,N_49994,N_49754);
and UO_4924 (O_4924,N_49841,N_49986);
nor UO_4925 (O_4925,N_49889,N_49979);
or UO_4926 (O_4926,N_49969,N_49874);
or UO_4927 (O_4927,N_49929,N_49980);
or UO_4928 (O_4928,N_49913,N_49842);
nand UO_4929 (O_4929,N_49979,N_49951);
nand UO_4930 (O_4930,N_49960,N_49916);
xor UO_4931 (O_4931,N_49891,N_49892);
nor UO_4932 (O_4932,N_49881,N_49960);
or UO_4933 (O_4933,N_49887,N_49925);
nor UO_4934 (O_4934,N_49780,N_49822);
nor UO_4935 (O_4935,N_49938,N_49905);
nand UO_4936 (O_4936,N_49923,N_49763);
and UO_4937 (O_4937,N_49924,N_49882);
xnor UO_4938 (O_4938,N_49907,N_49858);
nor UO_4939 (O_4939,N_49987,N_49926);
nor UO_4940 (O_4940,N_49829,N_49808);
xnor UO_4941 (O_4941,N_49880,N_49953);
or UO_4942 (O_4942,N_49799,N_49802);
or UO_4943 (O_4943,N_49937,N_49804);
and UO_4944 (O_4944,N_49978,N_49841);
xor UO_4945 (O_4945,N_49784,N_49925);
and UO_4946 (O_4946,N_49907,N_49927);
and UO_4947 (O_4947,N_49883,N_49984);
or UO_4948 (O_4948,N_49801,N_49884);
and UO_4949 (O_4949,N_49986,N_49914);
nor UO_4950 (O_4950,N_49887,N_49791);
xor UO_4951 (O_4951,N_49850,N_49898);
nor UO_4952 (O_4952,N_49916,N_49931);
xnor UO_4953 (O_4953,N_49921,N_49827);
or UO_4954 (O_4954,N_49904,N_49981);
nand UO_4955 (O_4955,N_49943,N_49942);
xnor UO_4956 (O_4956,N_49862,N_49909);
xnor UO_4957 (O_4957,N_49768,N_49931);
nor UO_4958 (O_4958,N_49977,N_49921);
nor UO_4959 (O_4959,N_49752,N_49879);
or UO_4960 (O_4960,N_49946,N_49881);
nand UO_4961 (O_4961,N_49915,N_49779);
and UO_4962 (O_4962,N_49888,N_49998);
nor UO_4963 (O_4963,N_49874,N_49794);
xor UO_4964 (O_4964,N_49800,N_49809);
nor UO_4965 (O_4965,N_49758,N_49817);
or UO_4966 (O_4966,N_49893,N_49843);
and UO_4967 (O_4967,N_49882,N_49761);
nor UO_4968 (O_4968,N_49814,N_49915);
xnor UO_4969 (O_4969,N_49947,N_49976);
or UO_4970 (O_4970,N_49808,N_49751);
or UO_4971 (O_4971,N_49816,N_49772);
and UO_4972 (O_4972,N_49894,N_49778);
nor UO_4973 (O_4973,N_49832,N_49956);
nand UO_4974 (O_4974,N_49802,N_49839);
xor UO_4975 (O_4975,N_49945,N_49839);
or UO_4976 (O_4976,N_49888,N_49935);
nand UO_4977 (O_4977,N_49956,N_49858);
and UO_4978 (O_4978,N_49831,N_49811);
or UO_4979 (O_4979,N_49980,N_49911);
nor UO_4980 (O_4980,N_49817,N_49945);
xor UO_4981 (O_4981,N_49835,N_49851);
nand UO_4982 (O_4982,N_49897,N_49938);
xor UO_4983 (O_4983,N_49833,N_49953);
nand UO_4984 (O_4984,N_49976,N_49889);
and UO_4985 (O_4985,N_49971,N_49948);
xnor UO_4986 (O_4986,N_49949,N_49839);
nor UO_4987 (O_4987,N_49860,N_49772);
xnor UO_4988 (O_4988,N_49983,N_49799);
nand UO_4989 (O_4989,N_49795,N_49867);
nand UO_4990 (O_4990,N_49759,N_49791);
nor UO_4991 (O_4991,N_49866,N_49909);
and UO_4992 (O_4992,N_49871,N_49875);
xnor UO_4993 (O_4993,N_49785,N_49909);
nand UO_4994 (O_4994,N_49774,N_49977);
and UO_4995 (O_4995,N_49781,N_49787);
xnor UO_4996 (O_4996,N_49816,N_49812);
xor UO_4997 (O_4997,N_49882,N_49821);
xnor UO_4998 (O_4998,N_49891,N_49788);
nor UO_4999 (O_4999,N_49988,N_49952);
endmodule