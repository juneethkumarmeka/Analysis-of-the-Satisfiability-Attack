module basic_3000_30000_3500_100_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_560,In_15);
nand U1 (N_1,In_209,In_2725);
and U2 (N_2,In_1160,In_457);
nor U3 (N_3,In_723,In_2555);
nand U4 (N_4,In_2752,In_1204);
or U5 (N_5,In_955,In_2327);
xor U6 (N_6,In_783,In_181);
nand U7 (N_7,In_494,In_1326);
or U8 (N_8,In_472,In_2779);
nor U9 (N_9,In_1230,In_1840);
nor U10 (N_10,In_1596,In_589);
nor U11 (N_11,In_1377,In_978);
nor U12 (N_12,In_902,In_1576);
xnor U13 (N_13,In_1397,In_2584);
and U14 (N_14,In_263,In_2530);
nand U15 (N_15,In_1359,In_2435);
or U16 (N_16,In_1499,In_2583);
xor U17 (N_17,In_1318,In_1121);
xnor U18 (N_18,In_767,In_1093);
xor U19 (N_19,In_2238,In_2589);
or U20 (N_20,In_1563,In_897);
nand U21 (N_21,In_1613,In_56);
nand U22 (N_22,In_657,In_1082);
or U23 (N_23,In_2654,In_1587);
nand U24 (N_24,In_982,In_2223);
nor U25 (N_25,In_1772,In_642);
xnor U26 (N_26,In_1213,In_2153);
or U27 (N_27,In_2791,In_23);
xor U28 (N_28,In_213,In_516);
nand U29 (N_29,In_2684,In_1723);
nor U30 (N_30,In_775,In_1151);
or U31 (N_31,In_1939,In_1429);
nand U32 (N_32,In_1057,In_1663);
and U33 (N_33,In_1292,In_475);
and U34 (N_34,In_1074,In_238);
nand U35 (N_35,In_2813,In_1167);
and U36 (N_36,In_2459,In_561);
nor U37 (N_37,In_2982,In_2449);
and U38 (N_38,In_2298,In_2861);
nand U39 (N_39,In_449,In_2189);
nand U40 (N_40,In_1743,In_1207);
nor U41 (N_41,In_1411,In_1937);
nor U42 (N_42,In_448,In_1741);
and U43 (N_43,In_2048,In_2894);
nor U44 (N_44,In_2321,In_1978);
or U45 (N_45,In_1878,In_490);
nor U46 (N_46,In_761,In_2563);
and U47 (N_47,In_2879,In_113);
nor U48 (N_48,In_1451,In_1693);
nand U49 (N_49,In_2084,In_1822);
xnor U50 (N_50,In_2182,In_1386);
nand U51 (N_51,In_1503,In_1086);
and U52 (N_52,In_1801,In_567);
or U53 (N_53,In_2920,In_2427);
nand U54 (N_54,In_1977,In_1431);
or U55 (N_55,In_308,In_2102);
or U56 (N_56,In_1214,In_2544);
nor U57 (N_57,In_21,In_525);
nor U58 (N_58,In_1242,In_678);
nor U59 (N_59,In_1833,In_752);
xor U60 (N_60,In_2837,In_6);
or U61 (N_61,In_2925,In_931);
nor U62 (N_62,In_2500,In_816);
or U63 (N_63,In_973,In_2436);
and U64 (N_64,In_1385,In_739);
nand U65 (N_65,In_712,In_2440);
and U66 (N_66,In_969,In_1362);
and U67 (N_67,In_1552,In_161);
nor U68 (N_68,In_2383,In_2012);
and U69 (N_69,In_2739,In_1188);
nand U70 (N_70,In_1004,In_2208);
xor U71 (N_71,In_215,In_2319);
or U72 (N_72,In_1845,In_857);
nand U73 (N_73,In_2479,In_764);
and U74 (N_74,In_971,In_252);
nand U75 (N_75,In_1664,In_2411);
xor U76 (N_76,In_915,In_160);
or U77 (N_77,In_1256,In_1967);
nor U78 (N_78,In_2301,In_1756);
or U79 (N_79,In_1487,In_1248);
xnor U80 (N_80,In_1703,In_944);
nor U81 (N_81,In_740,In_2767);
nor U82 (N_82,In_1506,In_48);
nor U83 (N_83,In_429,In_1330);
xor U84 (N_84,In_2745,In_519);
nor U85 (N_85,In_1244,In_1818);
nand U86 (N_86,In_2250,In_1905);
nor U87 (N_87,In_33,In_2805);
nor U88 (N_88,In_706,In_608);
xor U89 (N_89,In_1958,In_1518);
nand U90 (N_90,In_2026,In_2797);
nor U91 (N_91,In_2460,In_937);
nor U92 (N_92,In_2075,In_1372);
or U93 (N_93,In_1044,In_2878);
or U94 (N_94,In_242,In_2986);
nor U95 (N_95,In_2516,In_2082);
nand U96 (N_96,In_929,In_2409);
or U97 (N_97,In_175,In_2807);
nand U98 (N_98,In_63,In_1488);
nand U99 (N_99,In_855,In_2098);
or U100 (N_100,In_1711,In_1562);
xor U101 (N_101,In_2175,In_1025);
or U102 (N_102,In_2509,In_588);
xnor U103 (N_103,In_1989,In_1289);
and U104 (N_104,In_1141,In_2361);
or U105 (N_105,In_1998,In_2672);
nor U106 (N_106,In_866,In_2497);
and U107 (N_107,In_1096,In_940);
xor U108 (N_108,In_1980,In_1863);
xor U109 (N_109,In_627,In_316);
xor U110 (N_110,In_1944,In_2609);
nor U111 (N_111,In_1672,In_822);
xor U112 (N_112,In_2748,In_250);
or U113 (N_113,In_1018,In_1892);
and U114 (N_114,In_2483,In_2425);
or U115 (N_115,In_2498,In_192);
and U116 (N_116,In_687,In_2611);
or U117 (N_117,In_2569,In_2195);
xor U118 (N_118,In_827,In_1106);
nand U119 (N_119,In_1333,In_2836);
xor U120 (N_120,In_795,In_2994);
or U121 (N_121,In_1287,In_1066);
nand U122 (N_122,In_1728,In_2608);
or U123 (N_123,In_1946,In_364);
nor U124 (N_124,In_2707,In_180);
nor U125 (N_125,In_1639,In_1231);
nand U126 (N_126,In_596,In_1056);
or U127 (N_127,In_41,In_1886);
and U128 (N_128,In_1896,In_2822);
nand U129 (N_129,In_2732,In_1625);
nor U130 (N_130,In_1316,In_1675);
or U131 (N_131,In_1669,In_1667);
xnor U132 (N_132,In_653,In_899);
nor U133 (N_133,In_340,In_1183);
or U134 (N_134,In_549,In_2222);
nor U135 (N_135,In_942,In_1280);
or U136 (N_136,In_2272,In_1228);
or U137 (N_137,In_2261,In_2641);
or U138 (N_138,In_2566,In_2741);
and U139 (N_139,In_1714,In_2370);
nor U140 (N_140,In_2667,In_535);
xor U141 (N_141,In_52,In_86);
nor U142 (N_142,In_1810,In_2006);
and U143 (N_143,In_1478,In_2580);
nand U144 (N_144,In_1002,In_1284);
or U145 (N_145,In_1750,In_579);
nor U146 (N_146,In_1238,In_1935);
nand U147 (N_147,In_1904,In_1374);
nor U148 (N_148,In_1995,In_37);
nor U149 (N_149,In_2257,In_468);
xor U150 (N_150,In_436,In_1195);
and U151 (N_151,In_2220,In_2282);
and U152 (N_152,In_2452,In_2535);
nand U153 (N_153,In_1285,In_2088);
nand U154 (N_154,In_677,In_1538);
xnor U155 (N_155,In_1361,In_2558);
and U156 (N_156,In_948,In_2299);
nand U157 (N_157,In_1715,In_2600);
or U158 (N_158,In_2653,In_322);
or U159 (N_159,In_458,In_2709);
or U160 (N_160,In_2011,In_599);
xor U161 (N_161,In_1607,In_2377);
nor U162 (N_162,In_580,In_1708);
xor U163 (N_163,In_1688,In_39);
or U164 (N_164,In_1321,In_2884);
and U165 (N_165,In_1761,In_74);
nand U166 (N_166,In_530,In_2874);
and U167 (N_167,In_2616,In_1334);
nor U168 (N_168,In_652,In_184);
or U169 (N_169,In_2700,In_1090);
or U170 (N_170,In_190,In_1283);
nor U171 (N_171,In_952,In_2806);
nand U172 (N_172,In_1125,In_966);
nor U173 (N_173,In_2587,In_97);
xor U174 (N_174,In_665,In_2306);
nand U175 (N_175,In_2400,In_341);
nand U176 (N_176,In_2079,In_363);
and U177 (N_177,In_2723,In_2447);
nand U178 (N_178,In_1960,In_146);
nor U179 (N_179,In_64,In_2151);
and U180 (N_180,In_504,In_2169);
nor U181 (N_181,In_537,In_1114);
or U182 (N_182,In_1144,In_2163);
nand U183 (N_183,In_2539,In_1145);
nor U184 (N_184,In_1441,In_2338);
xnor U185 (N_185,In_2277,In_2139);
nor U186 (N_186,In_1762,In_498);
nand U187 (N_187,In_2107,In_151);
nand U188 (N_188,In_601,In_566);
nor U189 (N_189,In_2532,In_65);
or U190 (N_190,In_981,In_2283);
and U191 (N_191,In_1665,In_1001);
nand U192 (N_192,In_1521,In_983);
and U193 (N_193,In_2154,In_786);
nand U194 (N_194,In_284,In_426);
xnor U195 (N_195,In_2210,In_1961);
nand U196 (N_196,In_2540,In_2716);
or U197 (N_197,In_1486,In_745);
or U198 (N_198,In_1908,In_1799);
or U199 (N_199,In_1749,In_1268);
and U200 (N_200,In_378,In_1738);
nand U201 (N_201,In_550,In_1040);
nand U202 (N_202,In_1541,In_255);
nor U203 (N_203,In_1132,In_2200);
xor U204 (N_204,In_1449,In_531);
nand U205 (N_205,In_1857,In_1498);
xnor U206 (N_206,In_277,In_2506);
and U207 (N_207,In_1511,In_2938);
xor U208 (N_208,In_828,In_422);
nand U209 (N_209,In_205,In_1555);
nand U210 (N_210,In_546,In_2510);
and U211 (N_211,In_2381,In_751);
nor U212 (N_212,In_2568,In_2003);
xnor U213 (N_213,In_125,In_615);
nand U214 (N_214,In_480,In_2846);
and U215 (N_215,In_1171,In_1468);
or U216 (N_216,In_1924,In_2412);
nand U217 (N_217,In_1437,In_1055);
or U218 (N_218,In_572,In_405);
xnor U219 (N_219,In_829,In_843);
and U220 (N_220,In_1860,In_796);
and U221 (N_221,In_651,In_1861);
and U222 (N_222,In_2696,In_492);
xnor U223 (N_223,In_1088,In_1463);
xnor U224 (N_224,In_2028,In_2731);
xnor U225 (N_225,In_2369,In_1376);
xnor U226 (N_226,In_1770,In_38);
or U227 (N_227,In_844,In_555);
nor U228 (N_228,In_842,In_854);
or U229 (N_229,In_1149,In_1842);
xor U230 (N_230,In_2680,In_1578);
nor U231 (N_231,In_2576,In_2567);
xor U232 (N_232,In_1277,In_1869);
nor U233 (N_233,In_766,In_1829);
nand U234 (N_234,In_401,In_1077);
nor U235 (N_235,In_2475,In_235);
nand U236 (N_236,In_1549,In_76);
nand U237 (N_237,In_109,In_2);
nand U238 (N_238,In_1251,In_2701);
or U239 (N_239,In_600,In_569);
nor U240 (N_240,In_934,In_2534);
nor U241 (N_241,In_179,In_2360);
or U242 (N_242,In_353,In_2749);
nor U243 (N_243,In_434,In_2678);
xor U244 (N_244,In_1673,In_2118);
nor U245 (N_245,In_228,In_619);
nor U246 (N_246,In_2845,In_1514);
or U247 (N_247,In_1666,In_2668);
nor U248 (N_248,In_2166,In_49);
xor U249 (N_249,In_1222,In_1203);
nand U250 (N_250,In_2599,In_1925);
nand U251 (N_251,In_1197,In_2219);
xnor U252 (N_252,In_2478,In_2788);
nand U253 (N_253,In_2236,In_1571);
or U254 (N_254,In_411,In_1296);
or U255 (N_255,In_1982,In_732);
nand U256 (N_256,In_278,In_330);
or U257 (N_257,In_1603,In_2081);
nand U258 (N_258,In_320,In_2197);
nor U259 (N_259,In_2122,In_1101);
xor U260 (N_260,In_836,In_1454);
and U261 (N_261,In_282,In_2126);
or U262 (N_262,In_1279,In_208);
xor U263 (N_263,In_2489,In_2612);
and U264 (N_264,In_1636,In_1765);
xor U265 (N_265,In_2985,In_990);
and U266 (N_266,In_1120,In_464);
and U267 (N_267,In_730,In_243);
nor U268 (N_268,In_486,In_747);
nand U269 (N_269,In_2715,In_2183);
nor U270 (N_270,In_374,In_718);
nand U271 (N_271,In_82,In_2512);
nor U272 (N_272,In_2009,In_609);
and U273 (N_273,In_1992,In_1075);
and U274 (N_274,In_626,In_1147);
nand U275 (N_275,In_1835,In_1718);
or U276 (N_276,In_2954,In_8);
or U277 (N_277,In_1897,In_2055);
and U278 (N_278,In_2018,In_2234);
nand U279 (N_279,In_1970,In_2094);
and U280 (N_280,In_1389,In_2916);
and U281 (N_281,In_1573,In_1480);
or U282 (N_282,In_1575,In_2634);
xor U283 (N_283,In_2691,In_1069);
and U284 (N_284,In_387,In_343);
xor U285 (N_285,In_185,In_384);
and U286 (N_286,In_2975,In_1632);
and U287 (N_287,In_42,In_565);
or U288 (N_288,In_887,In_2217);
nand U289 (N_289,In_80,In_1000);
nand U290 (N_290,In_883,In_2582);
nor U291 (N_291,In_2776,In_1653);
and U292 (N_292,In_2072,In_1061);
or U293 (N_293,In_2988,In_2635);
xnor U294 (N_294,In_595,In_1643);
or U295 (N_295,In_587,In_2621);
nor U296 (N_296,In_1224,In_427);
xor U297 (N_297,In_392,In_2083);
xor U298 (N_298,In_2742,In_1191);
nor U299 (N_299,In_2100,In_197);
and U300 (N_300,In_2466,In_1554);
and U301 (N_301,In_1791,In_512);
and U302 (N_302,In_2665,In_2968);
and U303 (N_303,In_1927,In_168);
xnor U304 (N_304,In_2834,In_1720);
nand U305 (N_305,In_1827,In_2625);
nand U306 (N_306,In_2935,In_1716);
nand U307 (N_307,In_920,In_2112);
nand U308 (N_308,In_2605,In_222);
and U309 (N_309,In_1348,In_2271);
xor U310 (N_310,In_2025,In_989);
and U311 (N_311,In_257,In_1914);
or U312 (N_312,In_892,In_2763);
nor U313 (N_313,In_1966,In_1239);
nor U314 (N_314,In_264,In_1391);
nor U315 (N_315,In_2840,In_123);
or U316 (N_316,In_224,In_1084);
nor U317 (N_317,In_1396,In_1751);
nor U318 (N_318,In_811,In_1852);
or U319 (N_319,In_1559,In_1903);
or U320 (N_320,In_2548,In_1009);
nand U321 (N_321,In_2157,In_2728);
or U322 (N_322,In_499,In_2529);
nor U323 (N_323,In_85,In_253);
nand U324 (N_324,N_2,In_1432);
nor U325 (N_325,In_1792,In_2897);
or U326 (N_326,In_2528,In_852);
and U327 (N_327,In_820,In_1194);
or U328 (N_328,In_2921,In_1803);
or U329 (N_329,In_1634,In_2521);
and U330 (N_330,In_2717,In_961);
xnor U331 (N_331,In_2346,In_2648);
nor U332 (N_332,In_1399,In_2486);
nor U333 (N_333,N_40,In_2291);
nor U334 (N_334,In_221,In_2946);
or U335 (N_335,In_2647,In_945);
or U336 (N_336,In_2775,In_1520);
and U337 (N_337,In_1536,In_2288);
and U338 (N_338,In_638,In_2706);
xnor U339 (N_339,In_1525,In_419);
nor U340 (N_340,In_105,N_282);
and U341 (N_341,N_125,In_1319);
nor U342 (N_342,In_1034,In_342);
or U343 (N_343,In_2434,In_762);
nand U344 (N_344,In_469,In_446);
or U345 (N_345,N_21,In_1107);
nor U346 (N_346,In_1050,In_1041);
nand U347 (N_347,N_243,In_1644);
nor U348 (N_348,In_174,In_2753);
nand U349 (N_349,N_141,In_1948);
or U350 (N_350,In_1199,In_2237);
or U351 (N_351,In_2642,In_2880);
nand U352 (N_352,In_1642,In_742);
or U353 (N_353,In_2646,In_46);
and U354 (N_354,In_61,N_77);
nor U355 (N_355,In_2670,In_2441);
and U356 (N_356,In_1365,In_2977);
and U357 (N_357,In_2829,In_2828);
and U358 (N_358,In_2367,In_515);
nor U359 (N_359,In_1648,In_1164);
and U360 (N_360,In_2146,In_799);
or U361 (N_361,N_117,In_1129);
and U362 (N_362,In_2150,In_846);
and U363 (N_363,In_861,N_79);
and U364 (N_364,In_1601,In_1479);
nand U365 (N_365,In_2565,In_603);
nand U366 (N_366,In_2300,In_1647);
nor U367 (N_367,In_834,In_2825);
nor U368 (N_368,N_236,In_1200);
nor U369 (N_369,In_2315,In_437);
nor U370 (N_370,In_311,In_81);
or U371 (N_371,In_1085,In_2418);
xnor U372 (N_372,In_119,In_510);
and U373 (N_373,In_950,In_2364);
nand U374 (N_374,N_187,In_2172);
xnor U375 (N_375,In_1079,In_2382);
and U376 (N_376,In_418,In_1553);
and U377 (N_377,In_2826,In_2727);
or U378 (N_378,In_2179,In_1260);
or U379 (N_379,In_1704,In_2482);
nor U380 (N_380,In_2631,In_204);
nor U381 (N_381,In_1918,In_1465);
or U382 (N_382,In_780,N_128);
nand U383 (N_383,In_1884,In_104);
and U384 (N_384,In_644,In_880);
or U385 (N_385,In_455,In_593);
nor U386 (N_386,In_1572,In_2135);
or U387 (N_387,In_992,N_258);
or U388 (N_388,In_586,In_1115);
xor U389 (N_389,N_18,In_1007);
xnor U390 (N_390,In_1609,In_2255);
nand U391 (N_391,In_1031,In_1097);
and U392 (N_392,In_2485,In_395);
and U393 (N_393,N_45,In_1133);
xnor U394 (N_394,In_111,In_987);
or U395 (N_395,In_1024,In_1300);
nor U396 (N_396,In_2420,N_171);
nand U397 (N_397,In_688,N_299);
nor U398 (N_398,In_1567,In_1032);
nand U399 (N_399,In_279,In_470);
and U400 (N_400,In_1352,In_2858);
or U401 (N_401,In_2948,In_466);
xnor U402 (N_402,In_777,In_156);
nor U403 (N_403,In_1705,In_126);
nor U404 (N_404,In_2821,In_248);
or U405 (N_405,In_2295,In_518);
and U406 (N_406,In_2765,In_1855);
or U407 (N_407,In_283,In_239);
xnor U408 (N_408,In_882,N_116);
and U409 (N_409,In_2015,In_1127);
or U410 (N_410,In_2689,N_111);
xnor U411 (N_411,In_1118,In_2127);
and U412 (N_412,In_2542,N_53);
and U413 (N_413,In_2450,N_247);
nor U414 (N_414,In_800,In_347);
xnor U415 (N_415,In_1641,In_1460);
nor U416 (N_416,In_947,In_1274);
nor U417 (N_417,In_16,In_1633);
and U418 (N_418,N_127,In_1973);
nand U419 (N_419,In_326,In_157);
nand U420 (N_420,In_219,In_2414);
nand U421 (N_421,In_1304,In_2650);
or U422 (N_422,In_251,In_970);
or U423 (N_423,In_1612,In_121);
and U424 (N_424,In_2093,In_2617);
nand U425 (N_425,In_2125,In_2302);
and U426 (N_426,In_1181,In_986);
and U427 (N_427,In_1654,In_2116);
and U428 (N_428,In_833,In_1885);
nand U429 (N_429,In_2110,In_1325);
and U430 (N_430,In_186,In_2324);
xor U431 (N_431,In_1364,In_417);
nand U432 (N_432,N_25,In_1253);
or U433 (N_433,In_1427,N_238);
and U434 (N_434,In_2761,In_57);
nor U435 (N_435,In_2317,In_1781);
nor U436 (N_436,N_139,In_1452);
nor U437 (N_437,In_2817,In_1193);
nand U438 (N_438,In_2493,In_1635);
or U439 (N_439,In_260,In_1063);
and U440 (N_440,In_1802,N_280);
nor U441 (N_441,In_1393,In_2556);
xor U442 (N_442,In_439,In_527);
xnor U443 (N_443,In_1360,In_1906);
xnor U444 (N_444,In_1866,In_2844);
nor U445 (N_445,In_432,In_200);
nand U446 (N_446,In_2594,N_206);
and U447 (N_447,In_397,In_1136);
or U448 (N_448,In_289,N_178);
and U449 (N_449,In_2071,In_1786);
nand U450 (N_450,In_1698,In_1991);
and U451 (N_451,In_1558,N_24);
or U452 (N_452,In_440,In_443);
xnor U453 (N_453,In_1152,In_2495);
xor U454 (N_454,In_467,In_336);
and U455 (N_455,In_1223,In_576);
and U456 (N_456,In_2827,In_1697);
or U457 (N_457,In_372,In_2269);
xor U458 (N_458,In_2909,N_85);
and U459 (N_459,In_354,In_993);
and U460 (N_460,In_2117,In_1684);
and U461 (N_461,In_592,In_2365);
nor U462 (N_462,In_860,In_605);
nand U463 (N_463,In_1619,In_1282);
and U464 (N_464,In_893,In_136);
nor U465 (N_465,In_112,In_1767);
nor U466 (N_466,N_295,In_621);
or U467 (N_467,In_2129,N_191);
xnor U468 (N_468,In_2962,In_1600);
xnor U469 (N_469,In_2947,In_1546);
nor U470 (N_470,N_63,In_957);
and U471 (N_471,In_2216,N_138);
xor U472 (N_472,In_1509,In_695);
nor U473 (N_473,In_2702,In_2783);
xor U474 (N_474,In_1011,In_1685);
nand U475 (N_475,In_2314,In_202);
nor U476 (N_476,In_921,In_2443);
nor U477 (N_477,In_727,In_2736);
nand U478 (N_478,In_445,In_905);
and U479 (N_479,In_1245,In_1174);
or U480 (N_480,In_2471,In_1547);
or U481 (N_481,N_268,N_66);
nand U482 (N_482,In_726,N_108);
or U483 (N_483,In_1444,In_2134);
xor U484 (N_484,In_1343,N_293);
and U485 (N_485,In_1883,In_2734);
nand U486 (N_486,N_198,In_2148);
and U487 (N_487,N_267,In_210);
or U488 (N_488,In_2972,In_2526);
and U489 (N_489,In_58,In_962);
xor U490 (N_490,In_864,N_194);
xor U491 (N_491,In_998,N_10);
and U492 (N_492,In_801,In_1206);
nand U493 (N_493,N_130,In_1094);
nor U494 (N_494,N_168,In_1272);
nor U495 (N_495,In_2823,In_2659);
xnor U496 (N_496,In_2378,In_1629);
nor U497 (N_497,In_1891,In_1128);
nand U498 (N_498,In_2843,In_1489);
and U499 (N_499,In_1777,In_476);
nand U500 (N_500,In_410,In_1423);
or U501 (N_501,In_2224,In_2682);
nand U502 (N_502,In_1010,In_2898);
nand U503 (N_503,In_1899,In_32);
and U504 (N_504,In_2027,In_2784);
nand U505 (N_505,In_2347,In_187);
or U506 (N_506,N_189,N_106);
nand U507 (N_507,In_2240,N_277);
nor U508 (N_508,In_2405,In_2266);
nor U509 (N_509,In_2256,In_927);
or U510 (N_510,In_69,In_454);
or U511 (N_511,In_101,In_2484);
and U512 (N_512,In_1797,In_148);
nand U513 (N_513,In_2919,In_953);
xor U514 (N_514,In_1113,In_450);
and U515 (N_515,In_867,In_2014);
nor U516 (N_516,In_358,In_2666);
nand U517 (N_517,In_2998,In_13);
xnor U518 (N_518,In_2310,N_215);
or U519 (N_519,In_1344,In_1774);
nand U520 (N_520,In_2900,In_2651);
xor U521 (N_521,In_1651,In_2041);
nand U522 (N_522,N_237,In_2464);
and U523 (N_523,In_329,N_19);
xnor U524 (N_524,In_873,In_165);
nand U525 (N_525,In_1119,In_1261);
nand U526 (N_526,In_2348,In_689);
nand U527 (N_527,In_1033,In_637);
or U528 (N_528,In_2431,In_1130);
xnor U529 (N_529,In_2229,In_2368);
or U530 (N_530,In_1659,In_1065);
or U531 (N_531,In_894,In_2432);
and U532 (N_532,In_2991,In_398);
nand U533 (N_533,In_1126,In_756);
or U534 (N_534,In_1068,In_2652);
nor U535 (N_535,In_2918,In_2243);
and U536 (N_536,In_2944,In_170);
nor U537 (N_537,In_1754,In_217);
and U538 (N_538,In_2669,In_2403);
nand U539 (N_539,In_20,In_1543);
or U540 (N_540,In_2850,In_89);
xnor U541 (N_541,In_488,In_35);
xnor U542 (N_542,In_506,In_416);
nand U543 (N_543,In_681,In_541);
or U544 (N_544,In_994,In_90);
xor U545 (N_545,In_1780,In_1582);
or U546 (N_546,In_106,In_2187);
xor U547 (N_547,In_127,In_444);
nor U548 (N_548,In_1969,In_1436);
or U549 (N_549,In_2054,In_878);
nor U550 (N_550,In_2245,In_1273);
nand U551 (N_551,In_823,In_2588);
nor U552 (N_552,In_536,In_660);
or U553 (N_553,In_2456,In_2437);
nor U554 (N_554,In_2043,In_748);
or U555 (N_555,In_2001,In_1139);
nand U556 (N_556,In_1968,In_2729);
nand U557 (N_557,In_648,In_1358);
nor U558 (N_558,In_2740,In_377);
nor U559 (N_559,In_2010,In_2227);
xor U560 (N_560,N_123,In_1890);
nand U561 (N_561,In_421,In_513);
nor U562 (N_562,In_2326,In_2793);
xor U563 (N_563,N_7,In_1176);
or U564 (N_564,In_613,In_2461);
nor U565 (N_565,In_1327,In_870);
and U566 (N_566,In_362,In_178);
xor U567 (N_567,In_2161,In_1535);
or U568 (N_568,N_155,In_139);
nand U569 (N_569,In_1345,In_2592);
or U570 (N_570,In_2373,In_2688);
nand U571 (N_571,In_802,In_692);
xnor U572 (N_572,In_1800,In_1990);
nand U573 (N_573,In_1134,In_1314);
nor U574 (N_574,In_683,In_1026);
nor U575 (N_575,In_2984,In_290);
nand U576 (N_576,In_107,In_774);
nor U577 (N_577,In_1305,In_2362);
xnor U578 (N_578,In_646,In_2883);
or U579 (N_579,In_1594,In_1166);
or U580 (N_580,In_1768,In_847);
nand U581 (N_581,In_1856,N_131);
nand U582 (N_582,In_2915,In_2839);
nor U583 (N_583,In_1734,In_2671);
nor U584 (N_584,In_2737,In_714);
nor U585 (N_585,In_344,In_924);
xnor U586 (N_586,In_2849,In_2726);
or U587 (N_587,In_1453,In_2862);
and U588 (N_588,In_568,In_1874);
and U589 (N_589,In_1790,In_2375);
and U590 (N_590,In_1154,In_399);
or U591 (N_591,In_604,In_881);
nand U592 (N_592,N_96,N_55);
nand U593 (N_593,In_1604,In_2922);
or U594 (N_594,In_2069,In_386);
nor U595 (N_595,In_2549,In_1313);
and U596 (N_596,In_1182,N_213);
nor U597 (N_597,In_2552,In_913);
xor U598 (N_598,In_1976,In_2387);
nor U599 (N_599,In_1523,In_1551);
nor U600 (N_600,In_1934,In_911);
and U601 (N_601,In_2814,In_2876);
or U602 (N_602,In_169,In_1621);
nor U603 (N_603,N_409,N_140);
nand U604 (N_604,In_2867,In_1306);
or U605 (N_605,In_1917,N_372);
nor U606 (N_606,In_2202,N_84);
and U607 (N_607,In_1219,In_1258);
nor U608 (N_608,In_415,In_2395);
and U609 (N_609,In_832,N_70);
or U610 (N_610,N_441,N_56);
and U611 (N_611,In_214,In_1782);
xnor U612 (N_612,In_2303,N_514);
nor U613 (N_613,In_699,In_794);
nor U614 (N_614,In_1233,In_839);
nor U615 (N_615,In_2002,In_2531);
and U616 (N_616,In_655,In_930);
nor U617 (N_617,N_502,In_1356);
or U618 (N_618,In_7,N_564);
or U619 (N_619,N_520,In_1433);
or U620 (N_620,In_1387,In_1293);
xor U621 (N_621,In_47,In_862);
nor U622 (N_622,In_1534,In_1286);
xnor U623 (N_623,In_1796,In_2074);
nand U624 (N_624,In_1721,In_147);
or U625 (N_625,In_2718,In_367);
nand U626 (N_626,In_2595,In_2092);
nand U627 (N_627,In_532,In_303);
xor U628 (N_628,N_91,In_120);
xnor U629 (N_629,In_158,In_1159);
nand U630 (N_630,N_43,In_1919);
xnor U631 (N_631,In_2490,In_1415);
nand U632 (N_632,N_273,N_150);
and U633 (N_633,N_281,In_1524);
nand U634 (N_634,N_4,In_618);
nor U635 (N_635,N_239,N_590);
xor U636 (N_636,In_2355,In_2713);
and U637 (N_637,In_710,In_1769);
or U638 (N_638,In_487,N_315);
nor U639 (N_639,N_455,In_1528);
or U640 (N_640,In_92,In_1422);
nor U641 (N_641,In_817,In_965);
and U642 (N_642,In_2607,In_545);
and U643 (N_643,N_216,In_1059);
or U644 (N_644,In_227,In_2286);
xnor U645 (N_645,N_344,In_1505);
or U646 (N_646,N_222,In_2772);
and U647 (N_647,N_452,N_510);
and U648 (N_648,In_1657,N_269);
nand U649 (N_649,In_1053,In_685);
and U650 (N_650,In_521,In_79);
nand U651 (N_651,In_2316,In_1017);
xor U652 (N_652,N_588,In_1628);
and U653 (N_653,In_1220,In_2931);
or U654 (N_654,In_465,In_1373);
or U655 (N_655,In_1513,N_229);
nand U656 (N_656,In_223,In_2160);
nor U657 (N_657,In_622,In_2782);
xor U658 (N_658,In_2242,N_580);
or U659 (N_659,In_2708,In_2914);
xor U660 (N_660,In_1472,N_124);
nand U661 (N_661,In_2494,In_722);
or U662 (N_662,N_39,In_2546);
or U663 (N_663,In_2439,In_2020);
nand U664 (N_664,N_22,In_2577);
xor U665 (N_665,In_2337,In_1442);
nand U666 (N_666,In_2724,In_137);
and U667 (N_667,In_1887,N_287);
xnor U668 (N_668,In_988,In_556);
nor U669 (N_669,N_537,In_935);
or U670 (N_670,In_1496,N_148);
nor U671 (N_671,In_564,N_369);
nor U672 (N_672,In_1038,N_184);
or U673 (N_673,In_2407,In_1776);
xor U674 (N_674,In_890,N_188);
nor U675 (N_675,In_431,N_146);
nand U676 (N_676,N_59,N_278);
xor U677 (N_677,In_2799,In_744);
xor U678 (N_678,In_964,In_2164);
and U679 (N_679,In_2560,In_976);
nor U680 (N_680,In_1872,In_2472);
or U681 (N_681,In_1830,In_2000);
or U682 (N_682,In_1854,In_578);
nand U683 (N_683,N_358,In_218);
nor U684 (N_684,In_203,In_1210);
or U685 (N_685,N_120,N_157);
xor U686 (N_686,In_51,In_2868);
and U687 (N_687,In_500,In_1380);
nor U688 (N_688,In_2487,In_1264);
nand U689 (N_689,N_470,N_361);
nand U690 (N_690,N_205,N_363);
nand U691 (N_691,N_418,In_1679);
xor U692 (N_692,In_1589,In_1565);
nor U693 (N_693,In_2533,In_1335);
nand U694 (N_694,In_1375,N_592);
nand U695 (N_695,N_567,In_154);
nand U696 (N_696,N_518,In_2413);
xor U697 (N_697,In_967,In_292);
xor U698 (N_698,N_32,In_28);
nor U699 (N_699,In_503,N_98);
xnor U700 (N_700,In_2643,In_2343);
or U701 (N_701,In_1569,In_1466);
xnor U702 (N_702,In_2031,N_553);
xnor U703 (N_703,N_133,In_1901);
xor U704 (N_704,In_1848,N_383);
nor U705 (N_705,In_690,In_331);
nand U706 (N_706,In_1996,In_2292);
xnor U707 (N_707,In_649,In_420);
or U708 (N_708,In_2996,N_513);
or U709 (N_709,In_1072,In_388);
xnor U710 (N_710,In_731,In_1329);
or U711 (N_711,In_2593,N_469);
nand U712 (N_712,In_803,N_407);
nand U713 (N_713,In_2618,In_1157);
xnor U714 (N_714,N_448,In_1865);
nand U715 (N_715,In_2068,In_481);
and U716 (N_716,In_2564,In_1051);
xnor U717 (N_717,In_337,In_2514);
or U718 (N_718,In_889,In_383);
nor U719 (N_719,N_336,N_540);
xnor U720 (N_720,In_871,N_589);
xnor U721 (N_721,N_596,In_2067);
or U722 (N_722,In_2866,In_704);
nor U723 (N_723,In_575,In_2008);
and U724 (N_724,In_559,In_2750);
and U725 (N_725,N_450,In_298);
and U726 (N_726,In_1205,In_349);
and U727 (N_727,In_1913,In_94);
and U728 (N_728,In_2415,In_2438);
nand U729 (N_729,In_2204,In_54);
xnor U730 (N_730,In_1447,In_2394);
nand U731 (N_731,In_2144,In_300);
xnor U732 (N_732,In_2468,N_387);
and U733 (N_733,In_1317,In_2803);
nand U734 (N_734,In_2626,In_2191);
xnor U735 (N_735,In_376,In_1312);
nor U736 (N_736,In_2505,N_459);
nand U737 (N_737,In_2649,In_916);
nand U738 (N_738,In_1493,In_352);
and U739 (N_739,In_2029,In_1290);
nor U740 (N_740,N_475,In_1353);
nand U741 (N_741,In_2847,In_2557);
nor U742 (N_742,In_691,In_645);
nand U743 (N_743,N_482,In_669);
nand U744 (N_744,In_1828,N_220);
xnor U745 (N_745,In_2692,N_562);
or U746 (N_746,In_1766,In_781);
nor U747 (N_747,In_2332,In_2911);
nor U748 (N_748,In_2352,N_248);
nand U749 (N_749,N_263,In_2989);
nor U750 (N_750,In_2719,In_2804);
nor U751 (N_751,In_2279,In_1021);
nand U752 (N_752,In_2188,N_486);
and U753 (N_753,In_98,In_1142);
nor U754 (N_754,In_167,In_1881);
xor U755 (N_755,In_2396,N_457);
and U756 (N_756,In_2869,N_488);
nor U757 (N_757,N_31,In_382);
and U758 (N_758,In_686,N_473);
nand U759 (N_759,N_454,In_2152);
or U760 (N_760,In_2101,In_1650);
xnor U761 (N_761,In_1083,In_1196);
nand U762 (N_762,In_2681,In_2198);
or U763 (N_763,N_529,In_2596);
and U764 (N_764,In_2185,N_250);
or U765 (N_765,In_2201,In_1947);
nand U766 (N_766,In_2503,In_1254);
nor U767 (N_767,In_2973,In_570);
nor U768 (N_768,In_266,In_2873);
nor U769 (N_769,N_414,In_2630);
xor U770 (N_770,In_850,In_1859);
nor U771 (N_771,In_2176,In_528);
and U772 (N_772,In_509,N_583);
nand U773 (N_773,In_2036,In_1190);
nand U774 (N_774,N_464,N_530);
nand U775 (N_775,In_2320,In_496);
xnor U776 (N_776,In_634,N_3);
or U777 (N_777,In_1240,In_922);
xnor U778 (N_778,In_1515,In_2523);
or U779 (N_779,In_1581,In_939);
or U780 (N_780,In_102,In_1003);
or U781 (N_781,In_24,N_444);
and U782 (N_782,In_2334,In_968);
xnor U783 (N_783,In_1813,N_347);
and U784 (N_784,In_812,In_2392);
and U785 (N_785,In_1081,N_307);
nor U786 (N_786,In_2780,In_1435);
nor U787 (N_787,In_1255,In_538);
nor U788 (N_788,In_1421,N_162);
nand U789 (N_789,In_96,In_1339);
or U790 (N_790,In_2551,In_281);
or U791 (N_791,N_328,In_768);
xnor U792 (N_792,In_414,In_2091);
nor U793 (N_793,In_2059,In_735);
or U794 (N_794,In_1759,In_2927);
nor U795 (N_795,N_221,In_1184);
nor U796 (N_796,N_285,N_192);
xnor U797 (N_797,In_2934,In_424);
and U798 (N_798,N_214,In_2042);
nor U799 (N_799,N_29,In_2980);
and U800 (N_800,In_1178,In_540);
or U801 (N_801,In_1311,In_2639);
nand U802 (N_802,In_684,N_27);
nor U803 (N_803,In_919,In_676);
and U804 (N_804,In_782,In_2065);
or U805 (N_805,In_391,N_5);
and U806 (N_806,In_333,N_461);
xnor U807 (N_807,In_2893,In_1417);
or U808 (N_808,N_371,In_1320);
xor U809 (N_809,In_1952,In_1100);
nor U810 (N_810,N_368,N_538);
xor U811 (N_811,N_115,In_2842);
and U812 (N_812,N_332,In_859);
nand U813 (N_813,In_758,In_2448);
xnor U814 (N_814,In_482,N_442);
nor U815 (N_815,In_1678,In_2391);
xor U816 (N_816,In_507,In_2115);
xor U817 (N_817,In_1030,N_476);
and U818 (N_818,In_447,N_543);
nor U819 (N_819,In_2259,In_1585);
nor U820 (N_820,In_821,In_78);
nand U821 (N_821,N_201,In_452);
or U822 (N_822,N_331,In_173);
nor U823 (N_823,In_738,In_176);
nor U824 (N_824,N_193,N_584);
xnor U825 (N_825,In_327,In_1599);
or U826 (N_826,In_1692,N_367);
xnor U827 (N_827,In_2816,In_2262);
xnor U828 (N_828,In_848,In_11);
and U829 (N_829,N_121,N_81);
nand U830 (N_830,N_337,In_1482);
nor U831 (N_831,In_2309,In_297);
or U832 (N_832,N_547,In_909);
nor U833 (N_833,In_1839,In_1733);
or U834 (N_834,In_2455,In_1707);
and U835 (N_835,In_1138,N_270);
nor U836 (N_836,In_1109,In_1146);
or U837 (N_837,In_2061,In_233);
xnor U838 (N_838,In_381,In_2339);
nor U839 (N_839,In_140,N_154);
nor U840 (N_840,In_31,In_2778);
and U841 (N_841,In_2278,In_1894);
and U842 (N_842,N_14,In_863);
or U843 (N_843,In_1014,In_1590);
nand U844 (N_844,In_1162,In_1170);
xnor U845 (N_845,In_543,In_2225);
and U846 (N_846,N_506,N_404);
nand U847 (N_847,In_44,In_77);
and U848 (N_848,N_451,N_52);
and U849 (N_849,In_495,N_253);
xnor U850 (N_850,In_1087,N_391);
xnor U851 (N_851,N_431,In_2445);
xor U852 (N_852,In_2933,In_664);
xor U853 (N_853,In_1404,In_2585);
nor U854 (N_854,In_368,N_433);
or U855 (N_855,N_305,In_625);
and U856 (N_856,In_2203,In_122);
or U857 (N_857,In_787,In_729);
nor U858 (N_858,In_591,In_1428);
xor U859 (N_859,In_29,In_1804);
nor U860 (N_860,N_260,N_298);
nor U861 (N_861,In_1844,N_88);
and U862 (N_862,N_465,In_1249);
nand U863 (N_863,In_2444,In_2744);
nand U864 (N_864,In_628,In_1825);
or U865 (N_865,In_2598,N_339);
and U866 (N_866,N_217,N_251);
or U867 (N_867,In_355,In_2969);
nand U868 (N_868,N_340,In_1108);
nand U869 (N_869,In_2170,In_1974);
xor U870 (N_870,In_1724,In_2704);
and U871 (N_871,In_598,N_324);
or U872 (N_872,N_129,In_2357);
nor U873 (N_873,N_492,In_2086);
and U874 (N_874,In_772,N_246);
and U875 (N_875,In_2932,In_2623);
or U876 (N_876,In_144,N_227);
and U877 (N_877,In_1882,In_451);
nor U878 (N_878,N_548,In_1512);
nor U879 (N_879,N_185,In_2787);
xor U880 (N_880,In_2264,N_164);
nor U881 (N_881,N_435,In_2318);
xor U882 (N_882,In_310,In_997);
xor U883 (N_883,In_230,In_129);
nand U884 (N_884,In_1997,In_1413);
nand U885 (N_885,In_346,In_1627);
nor U886 (N_886,In_2501,In_760);
nand U887 (N_887,In_1784,In_912);
nand U888 (N_888,In_2852,N_385);
and U889 (N_889,In_189,In_2499);
nand U890 (N_890,In_1342,In_2945);
nor U891 (N_891,In_1446,N_80);
xor U892 (N_892,In_1473,In_366);
nand U893 (N_893,N_101,In_656);
or U894 (N_894,N_528,In_1757);
nor U895 (N_895,In_771,N_137);
nand U896 (N_896,N_423,N_478);
nor U897 (N_897,In_1384,In_1778);
nand U898 (N_898,In_360,In_350);
and U899 (N_899,In_1076,In_2354);
and U900 (N_900,In_1005,In_2290);
or U901 (N_901,In_1706,In_473);
and U902 (N_902,N_884,N_868);
or U903 (N_903,In_2685,In_612);
nand U904 (N_904,N_156,In_2133);
xnor U905 (N_905,N_809,In_1028);
nor U906 (N_906,In_1676,In_1789);
nor U907 (N_907,In_673,In_904);
and U908 (N_908,In_2467,In_269);
xnor U909 (N_909,In_2239,In_2978);
nor U910 (N_910,In_979,N_582);
nand U911 (N_911,In_1942,In_1263);
or U912 (N_912,In_936,In_2143);
nor U913 (N_913,In_2124,In_928);
xor U914 (N_914,In_703,N_438);
xor U915 (N_915,In_299,In_633);
and U916 (N_916,In_2136,In_679);
nand U917 (N_917,In_1158,In_2904);
xnor U918 (N_918,N_390,In_385);
or U919 (N_919,In_1221,In_2024);
nand U920 (N_920,In_1073,N_200);
or U921 (N_921,N_294,In_1938);
or U922 (N_922,In_884,In_552);
nor U923 (N_923,In_563,In_1631);
xor U924 (N_924,In_2507,N_546);
xnor U925 (N_925,N_271,In_2181);
and U926 (N_926,In_810,In_2912);
xnor U927 (N_927,In_1909,In_666);
xor U928 (N_928,In_663,In_2524);
and U929 (N_929,N_571,In_819);
nand U930 (N_930,N_628,In_412);
and U931 (N_931,N_643,In_1022);
xor U932 (N_932,In_1910,N_119);
or U933 (N_933,In_1853,In_2895);
xnor U934 (N_934,N_729,In_2114);
nor U935 (N_935,N_795,In_2940);
and U936 (N_936,In_2928,N_170);
xor U937 (N_937,N_365,In_393);
and U938 (N_938,N_16,In_2308);
and U939 (N_939,In_1351,N_731);
and U940 (N_940,N_110,N_144);
nand U941 (N_941,N_622,N_174);
nor U942 (N_942,N_815,In_2801);
xor U943 (N_943,N_747,In_680);
and U944 (N_944,N_93,In_2419);
nor U945 (N_945,N_388,In_1212);
or U946 (N_946,N_802,In_1155);
or U947 (N_947,In_1533,In_721);
nand U948 (N_948,In_87,In_1211);
and U949 (N_949,In_1652,N_397);
nand U950 (N_950,N_539,In_1725);
nand U951 (N_951,In_1036,N_639);
nor U952 (N_952,N_316,In_114);
nand U953 (N_953,In_357,In_261);
and U954 (N_954,N_578,In_1645);
nand U955 (N_955,N_793,In_150);
nand U956 (N_956,In_2207,N_103);
xor U957 (N_957,In_960,In_2138);
or U958 (N_958,In_2770,In_2206);
and U959 (N_959,In_1089,In_1726);
nor U960 (N_960,In_309,In_2005);
nand U961 (N_961,In_1940,N_655);
nor U962 (N_962,In_390,In_2465);
or U963 (N_963,In_59,In_2047);
or U964 (N_964,In_2964,In_896);
nand U965 (N_965,In_1867,N_75);
or U966 (N_966,N_350,In_792);
and U967 (N_967,N_870,In_2889);
or U968 (N_968,In_1297,N_593);
or U969 (N_969,N_757,In_1674);
and U970 (N_970,In_249,N_427);
nand U971 (N_971,In_2209,In_2212);
and U972 (N_972,In_562,In_1785);
nand U973 (N_973,In_1702,In_1713);
xor U974 (N_974,N_621,N_325);
and U975 (N_975,In_1605,In_2561);
nor U976 (N_976,N_446,In_2802);
nor U977 (N_977,In_2789,In_1624);
xnor U978 (N_978,In_1250,N_195);
nor U979 (N_979,In_765,In_1951);
and U980 (N_980,In_2952,In_2870);
nor U981 (N_981,In_793,N_755);
nor U982 (N_982,N_208,In_571);
nor U983 (N_983,N_663,N_641);
or U984 (N_984,In_2771,In_2331);
xnor U985 (N_985,In_2950,In_876);
nand U986 (N_986,In_2177,In_906);
xor U987 (N_987,In_1987,In_1414);
or U988 (N_988,In_1709,In_2913);
nand U989 (N_989,N_308,N_134);
nor U990 (N_990,In_1691,In_2389);
and U991 (N_991,In_2769,N_694);
xnor U992 (N_992,In_529,N_758);
xnor U993 (N_993,N_591,In_1788);
and U994 (N_994,N_426,In_2049);
xor U995 (N_995,N_889,In_1843);
or U996 (N_996,In_2076,In_1962);
and U997 (N_997,In_1570,N_736);
xor U998 (N_998,In_1722,N_17);
xnor U999 (N_999,N_288,In_36);
xnor U1000 (N_1000,N_725,N_323);
xor U1001 (N_1001,In_66,N_348);
and U1002 (N_1002,N_443,In_514);
and U1003 (N_1003,In_977,N_44);
and U1004 (N_1004,In_2457,In_295);
or U1005 (N_1005,In_2214,In_2356);
nor U1006 (N_1006,In_1815,N_313);
nor U1007 (N_1007,In_1112,N_410);
and U1008 (N_1008,In_30,In_1070);
or U1009 (N_1009,In_1983,In_2743);
xnor U1010 (N_1010,In_95,N_882);
or U1011 (N_1011,N_36,N_609);
nor U1012 (N_1012,In_617,N_668);
and U1013 (N_1013,In_2113,In_2759);
nand U1014 (N_1014,In_1809,In_773);
or U1015 (N_1015,In_1764,In_1753);
or U1016 (N_1016,N_824,In_886);
or U1017 (N_1017,N_175,In_1746);
nand U1018 (N_1018,In_1491,In_256);
nand U1019 (N_1019,N_319,N_58);
or U1020 (N_1020,In_910,In_149);
xnor U1021 (N_1021,In_483,In_2604);
or U1022 (N_1022,In_2832,In_212);
xnor U1023 (N_1023,N_301,N_494);
or U1024 (N_1024,In_2910,N_62);
nand U1025 (N_1025,In_2905,N_183);
nand U1026 (N_1026,In_1656,In_1930);
nand U1027 (N_1027,In_1308,In_2730);
nand U1028 (N_1028,In_2602,In_1366);
nor U1029 (N_1029,In_2863,In_1560);
xor U1030 (N_1030,In_2263,In_750);
nor U1031 (N_1031,N_676,N_64);
nor U1032 (N_1032,In_2178,N_730);
nor U1033 (N_1033,In_853,In_423);
nand U1034 (N_1034,N_437,N_392);
nand U1035 (N_1035,In_2619,In_1871);
nor U1036 (N_1036,In_2774,N_100);
xnor U1037 (N_1037,In_972,N_346);
nand U1038 (N_1038,N_661,In_1208);
xor U1039 (N_1039,N_165,In_2746);
nand U1040 (N_1040,In_1811,N_805);
xnor U1041 (N_1041,In_1347,In_548);
or U1042 (N_1042,In_497,In_2171);
nor U1043 (N_1043,In_2312,In_2384);
nor U1044 (N_1044,N_701,In_1931);
xnor U1045 (N_1045,N_432,N_161);
and U1046 (N_1046,In_1406,N_779);
nand U1047 (N_1047,N_445,N_819);
nand U1048 (N_1048,N_439,N_818);
and U1049 (N_1049,In_285,In_2285);
and U1050 (N_1050,N_523,In_1495);
nand U1051 (N_1051,N_594,N_672);
nor U1052 (N_1052,N_671,In_2410);
and U1053 (N_1053,N_695,In_1779);
nand U1054 (N_1054,In_2857,N_102);
nor U1055 (N_1055,N_774,N_727);
nor U1056 (N_1056,N_751,In_1662);
nand U1057 (N_1057,In_659,In_2800);
or U1058 (N_1058,In_2108,N_688);
xnor U1059 (N_1059,In_2571,In_711);
xor U1060 (N_1060,In_826,In_1202);
and U1061 (N_1061,N_145,N_257);
xnor U1062 (N_1062,In_974,In_858);
xor U1063 (N_1063,In_1270,In_1241);
and U1064 (N_1064,In_18,N_840);
nor U1065 (N_1065,N_720,N_355);
nand U1066 (N_1066,In_93,N_531);
xnor U1067 (N_1067,In_1545,In_103);
and U1068 (N_1068,In_195,In_606);
xnor U1069 (N_1069,In_2374,In_1045);
xnor U1070 (N_1070,In_2663,In_2981);
xor U1071 (N_1071,In_558,N_503);
or U1072 (N_1072,In_1269,In_534);
nor U1073 (N_1073,In_2907,In_1008);
nor U1074 (N_1074,In_1586,In_1368);
xnor U1075 (N_1075,In_166,In_2284);
or U1076 (N_1076,In_2683,N_835);
nor U1077 (N_1077,In_616,N_72);
xnor U1078 (N_1078,In_1965,N_849);
or U1079 (N_1079,In_2104,In_296);
nand U1080 (N_1080,N_581,In_1831);
or U1081 (N_1081,In_1458,N_878);
xnor U1082 (N_1082,In_275,In_668);
xor U1083 (N_1083,N_761,N_899);
and U1084 (N_1084,N_838,N_255);
or U1085 (N_1085,In_2192,N_211);
nor U1086 (N_1086,In_461,In_2268);
and U1087 (N_1087,In_413,In_1837);
nand U1088 (N_1088,In_1457,In_2875);
nor U1089 (N_1089,In_2211,N_69);
xor U1090 (N_1090,N_507,In_1655);
xor U1091 (N_1091,In_724,In_1900);
nor U1092 (N_1092,In_1915,In_797);
or U1093 (N_1093,N_524,In_1851);
and U1094 (N_1094,N_163,In_1189);
nor U1095 (N_1095,N_891,In_885);
nand U1096 (N_1096,N_453,N_781);
nor U1097 (N_1097,In_1793,In_1740);
nor U1098 (N_1098,N_692,N_318);
nand U1099 (N_1099,In_2451,N_796);
or U1100 (N_1100,N_636,N_690);
nand U1101 (N_1101,In_682,N_549);
xor U1102 (N_1102,In_1367,N_631);
or U1103 (N_1103,In_891,N_342);
nand U1104 (N_1104,In_1752,In_83);
xor U1105 (N_1105,In_2426,N_606);
and U1106 (N_1106,N_378,In_321);
and U1107 (N_1107,In_442,N_65);
nand U1108 (N_1108,In_88,N_235);
xor U1109 (N_1109,N_733,In_2287);
and U1110 (N_1110,N_186,N_61);
nor U1111 (N_1111,N_712,In_25);
xnor U1112 (N_1112,N_740,In_313);
or U1113 (N_1113,In_1192,In_2402);
xor U1114 (N_1114,In_2703,In_1060);
and U1115 (N_1115,In_2358,N_225);
nand U1116 (N_1116,In_1588,In_2251);
and U1117 (N_1117,N_78,In_1013);
xor U1118 (N_1118,In_2553,N_569);
xor U1119 (N_1119,In_2993,N_26);
and U1120 (N_1120,N_272,In_84);
nand U1121 (N_1121,N_704,In_1661);
and U1122 (N_1122,N_463,In_1841);
nor U1123 (N_1123,N_573,In_2349);
and U1124 (N_1124,N_196,In_1953);
nor U1125 (N_1125,N_702,N_735);
or U1126 (N_1126,N_673,N_362);
xor U1127 (N_1127,In_1950,In_2103);
nand U1128 (N_1128,In_522,N_491);
and U1129 (N_1129,In_171,In_477);
xnor U1130 (N_1130,In_1445,In_1583);
and U1131 (N_1131,In_2429,In_1440);
xor U1132 (N_1132,N_322,In_2926);
or U1133 (N_1133,N_417,In_55);
nand U1134 (N_1134,In_1755,N_698);
and U1135 (N_1135,In_159,In_2470);
nor U1136 (N_1136,N_0,In_1150);
nor U1137 (N_1137,In_2057,N_159);
nand U1138 (N_1138,N_788,N_877);
or U1139 (N_1139,In_1945,In_635);
nor U1140 (N_1140,In_1439,In_1870);
and U1141 (N_1141,In_1595,In_1388);
or U1142 (N_1142,In_1771,In_736);
and U1143 (N_1143,In_2353,In_2720);
xnor U1144 (N_1144,In_845,N_204);
and U1145 (N_1145,In_2835,In_956);
or U1146 (N_1146,In_2477,In_2831);
or U1147 (N_1147,In_1710,In_901);
xor U1148 (N_1148,N_674,In_1522);
and U1149 (N_1149,In_667,N_585);
nor U1150 (N_1150,N_499,N_291);
or U1151 (N_1151,In_2253,In_1379);
and U1152 (N_1152,N_811,In_1229);
xor U1153 (N_1153,In_791,In_244);
nor U1154 (N_1154,In_1080,N_886);
nor U1155 (N_1155,N_223,In_630);
nand U1156 (N_1156,In_2953,N_74);
nand U1157 (N_1157,In_824,N_421);
nor U1158 (N_1158,In_2891,N_710);
or U1159 (N_1159,In_2882,In_1775);
and U1160 (N_1160,In_641,In_155);
or U1161 (N_1161,N_879,In_2992);
and U1162 (N_1162,N_472,In_1923);
or U1163 (N_1163,In_1879,In_1763);
and U1164 (N_1164,In_2155,In_1880);
or U1165 (N_1165,In_1873,N_458);
or U1166 (N_1166,In_1727,N_791);
or U1167 (N_1167,In_2939,N_481);
xnor U1168 (N_1168,N_82,In_1209);
or U1169 (N_1169,N_801,In_1299);
nand U1170 (N_1170,In_2622,In_2180);
xor U1171 (N_1171,N_334,N_468);
nand U1172 (N_1172,In_2007,N_274);
or U1173 (N_1173,In_813,N_231);
xor U1174 (N_1174,N_551,In_72);
nor U1175 (N_1175,N_489,In_2232);
xnor U1176 (N_1176,In_2351,In_1671);
xnor U1177 (N_1177,In_2053,In_523);
and U1178 (N_1178,In_1928,In_206);
nand U1179 (N_1179,In_943,In_2610);
nor U1180 (N_1180,In_700,N_675);
and U1181 (N_1181,In_2872,In_2517);
and U1182 (N_1182,N_895,In_1338);
or U1183 (N_1183,In_307,In_365);
nor U1184 (N_1184,In_407,N_38);
nor U1185 (N_1185,In_2004,N_603);
and U1186 (N_1186,In_2971,In_2757);
nand U1187 (N_1187,In_2674,In_2342);
nor U1188 (N_1188,In_954,In_68);
xnor U1189 (N_1189,In_1117,N_769);
nand U1190 (N_1190,In_963,N_737);
nor U1191 (N_1191,In_2917,N_780);
xnor U1192 (N_1192,In_2997,N_732);
nor U1193 (N_1193,In_2908,N_449);
and U1194 (N_1194,In_1895,In_2156);
and U1195 (N_1195,N_379,In_268);
nand U1196 (N_1196,In_2442,In_2638);
nor U1197 (N_1197,N_810,In_2656);
and U1198 (N_1198,In_2590,In_2162);
xnor U1199 (N_1199,In_2274,In_2520);
nor U1200 (N_1200,In_2559,N_51);
nand U1201 (N_1201,In_898,N_34);
nand U1202 (N_1202,In_2754,In_1291);
or U1203 (N_1203,In_1098,In_959);
nand U1204 (N_1204,In_2871,In_2230);
nand U1205 (N_1205,In_602,In_1226);
and U1206 (N_1206,In_1424,In_2906);
nand U1207 (N_1207,N_104,N_689);
and U1208 (N_1208,In_1395,N_1123);
nor U1209 (N_1209,In_394,In_2899);
xnor U1210 (N_1210,In_717,N_219);
nand U1211 (N_1211,N_172,N_794);
nand U1212 (N_1212,N_940,In_640);
nor U1213 (N_1213,In_1736,In_1071);
and U1214 (N_1214,In_1542,In_2359);
nand U1215 (N_1215,In_1298,In_2522);
and U1216 (N_1216,N_977,In_1161);
nand U1217 (N_1217,In_814,N_1014);
nand U1218 (N_1218,In_1626,In_225);
and U1219 (N_1219,In_237,In_441);
and U1220 (N_1220,In_2463,N_289);
and U1221 (N_1221,In_338,In_2087);
nor U1222 (N_1222,N_1084,In_26);
nor U1223 (N_1223,In_2675,In_9);
nor U1224 (N_1224,In_1102,N_354);
xor U1225 (N_1225,N_987,In_1739);
nand U1226 (N_1226,In_2109,In_389);
nand U1227 (N_1227,In_1943,N_864);
or U1228 (N_1228,N_841,N_1179);
or U1229 (N_1229,N_825,N_942);
and U1230 (N_1230,N_1002,In_2062);
nor U1231 (N_1231,In_629,N_1049);
or U1232 (N_1232,In_2999,N_1032);
xnor U1233 (N_1233,In_754,In_1955);
xor U1234 (N_1234,N_1180,In_2168);
nor U1235 (N_1235,In_624,N_1166);
and U1236 (N_1236,In_2281,N_635);
or U1237 (N_1237,N_1070,N_773);
xor U1238 (N_1238,N_923,N_1071);
and U1239 (N_1239,N_691,In_900);
and U1240 (N_1240,In_1185,N_297);
xnor U1241 (N_1241,In_1443,N_284);
and U1242 (N_1242,N_1177,In_1826);
xor U1243 (N_1243,In_1532,N_739);
or U1244 (N_1244,In_2581,N_652);
or U1245 (N_1245,In_1064,In_2755);
and U1246 (N_1246,In_1165,In_2344);
or U1247 (N_1247,In_1058,N_1147);
or U1248 (N_1248,N_561,In_1979);
or U1249 (N_1249,In_2957,In_2196);
xnor U1250 (N_1250,In_1037,In_733);
and U1251 (N_1251,N_827,In_2855);
xnor U1252 (N_1252,In_1719,In_2060);
or U1253 (N_1253,N_135,In_2632);
nor U1254 (N_1254,In_1700,In_2023);
or U1255 (N_1255,N_911,In_1929);
or U1256 (N_1256,In_1864,In_324);
nand U1257 (N_1257,In_1467,N_314);
xnor U1258 (N_1258,In_1426,In_611);
and U1259 (N_1259,N_846,In_2690);
nand U1260 (N_1260,In_182,In_2241);
and U1261 (N_1261,In_2574,In_2215);
xnor U1262 (N_1262,In_2637,N_637);
nor U1263 (N_1263,In_273,In_1898);
nor U1264 (N_1264,N_166,In_2792);
nor U1265 (N_1265,N_57,N_839);
or U1266 (N_1266,In_373,In_317);
or U1267 (N_1267,N_556,N_1006);
and U1268 (N_1268,N_726,In_643);
xnor U1269 (N_1269,In_2017,In_1933);
xor U1270 (N_1270,In_2226,In_1288);
nor U1271 (N_1271,N_1149,In_1123);
nand U1272 (N_1272,In_778,N_986);
and U1273 (N_1273,In_2798,In_1156);
xnor U1274 (N_1274,N_338,N_1176);
and U1275 (N_1275,N_1078,N_869);
xnor U1276 (N_1276,In_2265,N_1199);
or U1277 (N_1277,In_2280,In_716);
nor U1278 (N_1278,In_917,In_1608);
nand U1279 (N_1279,N_820,N_95);
xor U1280 (N_1280,In_1042,In_877);
xnor U1281 (N_1281,N_309,In_1510);
nor U1282 (N_1282,In_2838,In_2687);
nor U1283 (N_1283,N_256,In_926);
nand U1284 (N_1284,N_1172,In_2231);
nor U1285 (N_1285,In_287,N_654);
nor U1286 (N_1286,In_348,In_1561);
and U1287 (N_1287,In_2644,In_2379);
or U1288 (N_1288,In_980,N_303);
and U1289 (N_1289,In_1216,N_558);
or U1290 (N_1290,In_177,In_2213);
nor U1291 (N_1291,In_505,In_1095);
or U1292 (N_1292,In_2951,In_2089);
nand U1293 (N_1293,N_722,In_1035);
and U1294 (N_1294,N_743,In_888);
and U1295 (N_1295,In_1019,In_1972);
nand U1296 (N_1296,N_992,N_480);
or U1297 (N_1297,N_113,N_1130);
nor U1298 (N_1298,N_177,In_2070);
and U1299 (N_1299,N_1086,In_1405);
nand U1300 (N_1300,N_349,N_477);
or U1301 (N_1301,N_1195,In_2541);
xor U1302 (N_1302,N_48,N_1089);
and U1303 (N_1303,N_888,In_544);
nand U1304 (N_1304,In_1658,In_319);
xor U1305 (N_1305,N_883,N_623);
or U1306 (N_1306,N_786,In_2399);
nand U1307 (N_1307,In_1806,In_511);
or U1308 (N_1308,In_141,N_1063);
or U1309 (N_1309,In_1135,In_2679);
nand U1310 (N_1310,In_1271,N_1141);
and U1311 (N_1311,In_1646,In_837);
nand U1312 (N_1312,In_2662,In_2603);
or U1313 (N_1313,N_1027,In_1964);
and U1314 (N_1314,In_1975,N_934);
and U1315 (N_1315,In_1849,N_560);
nand U1316 (N_1316,N_787,In_2614);
and U1317 (N_1317,In_1742,N_403);
xnor U1318 (N_1318,In_2660,In_220);
nand U1319 (N_1319,In_1381,In_2056);
and U1320 (N_1320,In_1893,In_1039);
xnor U1321 (N_1321,In_2673,In_91);
nand U1322 (N_1322,N_1190,N_893);
nor U1323 (N_1323,In_2812,N_916);
nor U1324 (N_1324,In_1747,In_270);
xnor U1325 (N_1325,In_2591,In_1907);
nor U1326 (N_1326,In_453,N_926);
or U1327 (N_1327,In_339,In_838);
or U1328 (N_1328,In_1824,N_707);
nand U1329 (N_1329,In_1143,N_151);
xnor U1330 (N_1330,In_132,N_1056);
and U1331 (N_1331,In_2627,N_808);
and U1332 (N_1332,In_805,N_575);
and U1333 (N_1333,N_566,N_865);
and U1334 (N_1334,N_906,In_288);
xnor U1335 (N_1335,In_2492,In_2121);
nand U1336 (N_1336,N_400,In_2233);
xor U1337 (N_1337,In_1731,In_40);
nor U1338 (N_1338,N_629,N_656);
or U1339 (N_1339,N_1036,N_1053);
or U1340 (N_1340,N_357,N_67);
nand U1341 (N_1341,In_636,In_2398);
or U1342 (N_1342,In_705,N_1077);
and U1343 (N_1343,N_842,N_703);
nor U1344 (N_1344,In_2258,In_1544);
nor U1345 (N_1345,N_1096,In_246);
nor U1346 (N_1346,N_1001,N_905);
nor U1347 (N_1347,In_1262,In_2064);
or U1348 (N_1348,N_995,N_424);
nor U1349 (N_1349,In_874,In_1243);
xor U1350 (N_1350,In_2714,N_764);
and U1351 (N_1351,In_1295,N_872);
xor U1352 (N_1352,In_1620,In_1383);
xor U1353 (N_1353,In_356,N_1189);
and U1354 (N_1354,In_1398,In_804);
and U1355 (N_1355,N_76,In_728);
nor U1356 (N_1356,N_713,In_2304);
xor U1357 (N_1357,N_376,In_2694);
nor U1358 (N_1358,In_291,N_706);
or U1359 (N_1359,In_2930,In_2406);
nor U1360 (N_1360,N_552,In_946);
or U1361 (N_1361,In_1623,In_2762);
or U1362 (N_1362,In_757,N_686);
xor U1363 (N_1363,In_788,N_684);
and U1364 (N_1364,In_240,In_2958);
xor U1365 (N_1365,In_741,In_759);
nand U1366 (N_1366,In_2329,In_831);
or U1367 (N_1367,In_1577,In_1092);
and U1368 (N_1368,N_946,N_532);
xor U1369 (N_1369,N_97,In_2294);
nand U1370 (N_1370,N_853,In_100);
nor U1371 (N_1371,In_276,In_34);
and U1372 (N_1372,N_207,In_2888);
or U1373 (N_1373,N_389,In_903);
and U1374 (N_1374,N_927,In_1485);
and U1375 (N_1375,N_6,N_832);
nand U1376 (N_1376,In_1131,In_196);
nor U1377 (N_1377,N_107,N_901);
nor U1378 (N_1378,N_290,N_991);
nor U1379 (N_1379,In_2106,N_1105);
or U1380 (N_1380,N_1008,N_959);
and U1381 (N_1381,In_2246,N_843);
nand U1382 (N_1382,N_1156,In_1412);
nand U1383 (N_1383,In_502,In_2929);
and U1384 (N_1384,N_967,In_2886);
nor U1385 (N_1385,In_2961,In_404);
or U1386 (N_1386,N_311,In_1936);
nand U1387 (N_1387,In_1140,In_1023);
xor U1388 (N_1388,N_863,In_2966);
xnor U1389 (N_1389,N_615,In_743);
nor U1390 (N_1390,N_1020,In_1122);
and U1391 (N_1391,N_579,In_294);
nand U1392 (N_1392,In_1773,In_2820);
xor U1393 (N_1393,N_1058,N_917);
xnor U1394 (N_1394,In_1006,N_829);
and U1395 (N_1395,In_1357,In_1020);
and U1396 (N_1396,N_181,N_696);
and U1397 (N_1397,N_925,In_19);
xor U1398 (N_1398,In_2979,In_1401);
or U1399 (N_1399,N_37,N_885);
or U1400 (N_1400,N_317,N_1112);
and U1401 (N_1401,In_2050,In_1838);
xor U1402 (N_1402,In_1817,N_568);
or U1403 (N_1403,In_1099,In_1760);
xnor U1404 (N_1404,N_1168,N_822);
xnor U1405 (N_1405,In_809,In_2491);
nor U1406 (N_1406,N_152,N_640);
and U1407 (N_1407,N_772,N_495);
xor U1408 (N_1408,In_1902,N_1025);
xor U1409 (N_1409,N_1142,In_985);
xnor U1410 (N_1410,In_707,In_406);
nand U1411 (N_1411,N_613,In_2790);
or U1412 (N_1412,In_2376,N_604);
or U1413 (N_1413,In_1349,In_1111);
nand U1414 (N_1414,In_2606,In_45);
and U1415 (N_1415,N_230,In_2633);
xnor U1416 (N_1416,In_2097,In_594);
nor U1417 (N_1417,N_765,N_861);
and U1418 (N_1418,N_685,N_460);
nand U1419 (N_1419,N_954,In_335);
xnor U1420 (N_1420,In_670,In_2341);
xnor U1421 (N_1421,In_2035,In_991);
or U1422 (N_1422,N_1140,N_874);
nand U1423 (N_1423,N_956,In_216);
and U1424 (N_1424,In_1668,In_784);
or U1425 (N_1425,N_1093,N_742);
and U1426 (N_1426,N_630,N_1035);
and U1427 (N_1427,N_512,In_1823);
nand U1428 (N_1428,N_972,In_2276);
nor U1429 (N_1429,In_1153,In_2416);
or U1430 (N_1430,In_1048,In_746);
nand U1431 (N_1431,In_2902,N_611);
or U1432 (N_1432,N_1088,In_1180);
nand U1433 (N_1433,In_351,In_75);
or U1434 (N_1434,In_2760,N_1083);
nand U1435 (N_1435,N_173,N_525);
or U1436 (N_1436,In_2385,N_782);
nand U1437 (N_1437,In_14,N_777);
nor U1438 (N_1438,N_1171,N_914);
xnor U1439 (N_1439,N_677,N_1158);
nor U1440 (N_1440,In_73,In_201);
or U1441 (N_1441,N_908,N_1162);
xor U1442 (N_1442,N_1074,In_2474);
nand U1443 (N_1443,In_2423,N_544);
nand U1444 (N_1444,In_2942,In_1683);
and U1445 (N_1445,N_687,In_2458);
xor U1446 (N_1446,N_15,In_2824);
nand U1447 (N_1447,In_2661,N_607);
xnor U1448 (N_1448,N_1151,N_1047);
xnor U1449 (N_1449,In_584,In_1236);
nor U1450 (N_1450,N_608,In_1148);
and U1451 (N_1451,N_9,N_68);
nand U1452 (N_1452,N_994,In_1794);
nand U1453 (N_1453,In_2401,In_869);
and U1454 (N_1454,In_590,N_226);
and U1455 (N_1455,N_557,In_2404);
and U1456 (N_1456,In_2090,In_2695);
and U1457 (N_1457,In_116,N_373);
nor U1458 (N_1458,N_860,N_826);
nand U1459 (N_1459,N_50,N_190);
xnor U1460 (N_1460,In_2686,N_1110);
nor U1461 (N_1461,In_1186,N_626);
xnor U1462 (N_1462,In_2397,N_1080);
and U1463 (N_1463,In_1888,N_799);
or U1464 (N_1464,In_1516,N_504);
or U1465 (N_1465,In_1169,In_1737);
nand U1466 (N_1466,In_143,In_484);
xor U1467 (N_1467,N_466,In_17);
xor U1468 (N_1468,In_975,In_379);
nand U1469 (N_1469,N_73,In_1294);
or U1470 (N_1470,In_1540,N_377);
xnor U1471 (N_1471,In_1798,N_768);
nand U1472 (N_1472,In_1957,In_2572);
or U1473 (N_1473,N_395,In_380);
and U1474 (N_1474,N_304,N_143);
and U1475 (N_1475,In_2085,N_821);
nand U1476 (N_1476,In_1556,In_526);
nor U1477 (N_1477,N_705,In_1402);
or U1478 (N_1478,N_1108,N_1043);
xnor U1479 (N_1479,N_771,N_23);
and U1480 (N_1480,N_425,In_2052);
or U1481 (N_1481,N_1023,In_539);
or U1482 (N_1482,N_259,In_1531);
or U1483 (N_1483,In_1732,N_859);
nand U1484 (N_1484,N_320,In_2077);
or U1485 (N_1485,In_2132,In_2527);
nor U1486 (N_1486,N_981,N_1065);
or U1487 (N_1487,In_2096,N_812);
or U1488 (N_1488,In_130,In_1419);
and U1489 (N_1489,In_2149,In_1430);
nor U1490 (N_1490,N_909,N_1038);
nand U1491 (N_1491,In_163,N_245);
nand U1492 (N_1492,N_158,N_862);
or U1493 (N_1493,In_2881,In_2819);
nor U1494 (N_1494,N_875,N_975);
nor U1495 (N_1495,N_784,In_557);
nor U1496 (N_1496,In_2586,In_2408);
nor U1497 (N_1497,In_2335,In_996);
xnor U1498 (N_1498,N_667,N_382);
or U1499 (N_1499,In_1816,In_1787);
or U1500 (N_1500,N_715,N_1098);
nand U1501 (N_1501,N_498,N_1336);
or U1502 (N_1502,In_402,N_1460);
nor U1503 (N_1503,N_1005,N_1224);
nor U1504 (N_1504,In_128,N_1320);
nand U1505 (N_1505,In_456,In_1748);
and U1506 (N_1506,N_345,N_612);
nor U1507 (N_1507,N_1415,In_301);
nor U1508 (N_1508,In_779,N_904);
or U1509 (N_1509,In_574,In_172);
or U1510 (N_1510,N_852,In_207);
nor U1511 (N_1511,N_1253,N_1432);
or U1512 (N_1512,In_2615,N_1359);
and U1513 (N_1513,N_1291,N_1144);
nor U1514 (N_1514,N_1353,In_2311);
or U1515 (N_1515,In_304,N_1303);
or U1516 (N_1516,N_326,In_2896);
and U1517 (N_1517,In_2751,N_650);
xor U1518 (N_1518,N_709,N_1013);
xnor U1519 (N_1519,In_693,N_1218);
xor U1520 (N_1520,N_1449,In_1690);
xnor U1521 (N_1521,N_234,N_647);
and U1522 (N_1522,N_1393,In_835);
nand U1523 (N_1523,In_1527,N_1424);
nand U1524 (N_1524,In_1922,N_996);
xnor U1525 (N_1525,N_1297,In_1985);
nand U1526 (N_1526,N_330,N_1092);
and U1527 (N_1527,In_53,N_988);
nand U1528 (N_1528,N_112,N_638);
or U1529 (N_1529,N_1378,N_900);
and U1530 (N_1530,N_572,In_50);
or U1531 (N_1531,In_851,In_755);
and U1532 (N_1532,In_280,N_642);
or U1533 (N_1533,In_675,In_403);
xor U1534 (N_1534,N_1325,In_1550);
or U1535 (N_1535,N_1427,N_816);
nor U1536 (N_1536,N_678,N_935);
nand U1537 (N_1537,In_607,In_2903);
xnor U1538 (N_1538,In_2597,In_1615);
nor U1539 (N_1539,N_1069,In_1201);
xor U1540 (N_1540,N_952,N_1411);
xor U1541 (N_1541,In_2421,In_1921);
and U1542 (N_1542,N_1055,In_2424);
or U1543 (N_1543,In_2270,N_1293);
nor U1544 (N_1544,In_334,In_697);
or U1545 (N_1545,N_327,N_1492);
or U1546 (N_1546,In_0,In_2851);
or U1547 (N_1547,N_1028,In_1469);
or U1548 (N_1548,N_479,N_1045);
nor U1549 (N_1549,In_1911,In_1941);
or U1550 (N_1550,N_399,In_1834);
nand U1551 (N_1551,N_1388,N_980);
nor U1552 (N_1552,N_1455,N_1066);
nor U1553 (N_1553,In_533,N_847);
and U1554 (N_1554,In_672,In_325);
and U1555 (N_1555,In_1232,In_696);
xnor U1556 (N_1556,N_1135,N_1232);
xnor U1557 (N_1557,In_737,N_1081);
and U1558 (N_1558,N_406,N_1316);
and U1559 (N_1559,N_614,N_1302);
or U1560 (N_1560,In_1354,In_2545);
xnor U1561 (N_1561,N_1277,N_1075);
or U1562 (N_1562,In_1889,In_1371);
nand U1563 (N_1563,N_533,In_234);
xnor U1564 (N_1564,N_1015,N_405);
nor U1565 (N_1565,N_1438,N_577);
or U1566 (N_1566,In_2570,N_1317);
or U1567 (N_1567,N_719,N_997);
xnor U1568 (N_1568,In_1218,In_1434);
xor U1569 (N_1569,N_1343,In_211);
and U1570 (N_1570,N_517,In_2345);
or U1571 (N_1571,In_1593,In_117);
xor U1572 (N_1572,N_402,N_149);
xnor U1573 (N_1573,N_1287,In_1920);
nor U1574 (N_1574,In_2887,In_1858);
nor U1575 (N_1575,N_1265,N_71);
nand U1576 (N_1576,N_806,In_1548);
nand U1577 (N_1577,In_1500,N_1389);
xnor U1578 (N_1578,In_2073,N_1472);
nand U1579 (N_1579,N_1207,N_565);
nor U1580 (N_1580,In_785,N_1379);
xnor U1581 (N_1581,In_2454,N_1368);
and U1582 (N_1582,In_2145,N_1402);
and U1583 (N_1583,In_1876,N_1399);
nand U1584 (N_1584,In_43,N_401);
xor U1585 (N_1585,In_1455,N_1496);
nand U1586 (N_1586,N_487,In_715);
nand U1587 (N_1587,N_1082,N_501);
nor U1588 (N_1588,In_194,In_1579);
or U1589 (N_1589,In_12,N_1364);
or U1590 (N_1590,In_2811,In_2924);
or U1591 (N_1591,In_1614,N_1436);
and U1592 (N_1592,N_598,In_1670);
nor U1593 (N_1593,N_1220,In_2785);
or U1594 (N_1594,In_2601,In_2865);
xnor U1595 (N_1595,In_2289,N_1187);
and U1596 (N_1596,N_13,In_2194);
xor U1597 (N_1597,N_711,N_1309);
nand U1598 (N_1598,In_1598,In_258);
xor U1599 (N_1599,In_489,N_1017);
or U1600 (N_1600,N_1248,N_550);
xnor U1601 (N_1601,N_1128,In_2140);
nor U1602 (N_1602,In_1795,N_1252);
nor U1603 (N_1603,In_1340,In_1916);
nor U1604 (N_1604,In_1682,In_1805);
and U1605 (N_1605,N_264,N_47);
nor U1606 (N_1606,In_2547,N_965);
xnor U1607 (N_1607,N_1004,N_1228);
nor U1608 (N_1608,N_1103,N_1000);
nor U1609 (N_1609,N_1373,In_2158);
xnor U1610 (N_1610,N_961,In_856);
or U1611 (N_1611,N_915,N_898);
nor U1612 (N_1612,N_1163,N_1229);
xnor U1613 (N_1613,N_1266,N_1113);
or U1614 (N_1614,N_343,N_1136);
nand U1615 (N_1615,In_1416,N_982);
xor U1616 (N_1616,N_430,N_798);
nand U1617 (N_1617,In_1302,N_597);
or U1618 (N_1618,N_1283,N_1137);
or U1619 (N_1619,N_1249,N_351);
nand U1620 (N_1620,In_849,In_2244);
xnor U1621 (N_1621,N_1387,N_1227);
nand U1622 (N_1622,In_597,N_1381);
nand U1623 (N_1623,N_1246,In_908);
or U1624 (N_1624,N_1160,In_1418);
xnor U1625 (N_1625,N_60,In_2167);
nand U1626 (N_1626,N_310,In_1504);
nand U1627 (N_1627,N_1118,In_1257);
nor U1628 (N_1628,In_583,N_1164);
nand U1629 (N_1629,In_1276,N_1264);
nand U1630 (N_1630,In_131,N_1219);
or U1631 (N_1631,N_1121,N_1263);
and U1632 (N_1632,In_474,In_2579);
xnor U1633 (N_1633,N_1288,N_854);
nor U1634 (N_1634,In_2710,In_1812);
and U1635 (N_1635,N_951,N_1471);
xor U1636 (N_1636,N_658,In_2051);
nor U1637 (N_1637,In_1862,N_1324);
and U1638 (N_1638,In_332,N_770);
xnor U1639 (N_1639,N_1299,In_254);
or U1640 (N_1640,N_1247,N_105);
and U1641 (N_1641,N_1429,In_2030);
xnor U1642 (N_1642,N_1462,N_1244);
nor U1643 (N_1643,N_1405,In_1476);
nor U1644 (N_1644,In_577,N_1120);
and U1645 (N_1645,N_254,In_1963);
xor U1646 (N_1646,N_610,N_962);
xnor U1647 (N_1647,N_576,N_1426);
or U1648 (N_1648,N_1476,In_2305);
or U1649 (N_1649,N_41,N_1250);
and U1650 (N_1650,In_2960,In_547);
and U1651 (N_1651,N_984,N_644);
or U1652 (N_1652,In_1875,In_702);
or U1653 (N_1653,N_697,In_60);
or U1654 (N_1654,In_1337,N_218);
nor U1655 (N_1655,N_823,N_394);
and U1656 (N_1656,N_1012,N_800);
and U1657 (N_1657,N_797,N_1242);
nor U1658 (N_1658,N_1461,In_1410);
xnor U1659 (N_1659,N_1243,N_1280);
or U1660 (N_1660,In_2099,In_1745);
xor U1661 (N_1661,N_1363,In_2372);
xor U1662 (N_1662,N_505,N_364);
nor U1663 (N_1663,In_1052,N_716);
and U1664 (N_1664,N_202,N_1167);
nor U1665 (N_1665,N_1463,In_2340);
nor U1666 (N_1666,N_1451,In_2080);
or U1667 (N_1667,In_371,In_995);
nand U1668 (N_1668,In_1215,In_2044);
or U1669 (N_1669,N_970,N_1477);
nand U1670 (N_1670,In_508,N_760);
or U1671 (N_1671,N_1361,In_749);
nor U1672 (N_1672,In_1382,In_2699);
nor U1673 (N_1673,N_286,N_1205);
xor U1674 (N_1674,N_837,In_2515);
xor U1675 (N_1675,In_2795,In_2677);
and U1676 (N_1676,In_1328,N_957);
or U1677 (N_1677,In_581,In_1012);
nor U1678 (N_1678,In_1622,N_46);
or U1679 (N_1679,N_1458,N_1124);
nand U1680 (N_1680,In_459,In_479);
or U1681 (N_1681,N_1338,N_1094);
or U1682 (N_1682,In_2796,In_226);
nand U1683 (N_1683,In_520,N_527);
nor U1684 (N_1684,In_2640,In_918);
nand U1685 (N_1685,N_1441,N_1327);
nor U1686 (N_1686,N_1374,In_553);
or U1687 (N_1687,N_1221,In_2794);
xor U1688 (N_1688,N_1307,In_694);
xnor U1689 (N_1689,In_2628,N_1109);
and U1690 (N_1690,N_867,N_1370);
and U1691 (N_1691,N_375,N_28);
nor U1692 (N_1692,In_2033,N_485);
and U1693 (N_1693,N_976,In_2711);
nand U1694 (N_1694,N_1145,N_1403);
xor U1695 (N_1695,In_2810,In_938);
nor U1696 (N_1696,N_1259,N_646);
and U1697 (N_1697,N_851,N_496);
nand U1698 (N_1698,In_1,N_857);
or U1699 (N_1699,In_430,In_2738);
nor U1700 (N_1700,N_1328,In_2693);
or U1701 (N_1701,N_1334,In_1699);
or U1702 (N_1702,In_907,N_1273);
nand U1703 (N_1703,In_198,N_1398);
nor U1704 (N_1704,In_2046,In_2856);
nor U1705 (N_1705,In_2193,N_209);
xnor U1706 (N_1706,N_92,In_713);
nand U1707 (N_1707,In_4,In_1574);
and U1708 (N_1708,N_1465,In_1564);
nor U1709 (N_1709,In_725,N_1060);
nor U1710 (N_1710,In_2959,N_1192);
or U1711 (N_1711,N_356,N_1367);
or U1712 (N_1712,In_425,N_1200);
nor U1713 (N_1713,N_1467,In_2063);
xnor U1714 (N_1714,In_1477,N_1054);
or U1715 (N_1715,In_2508,N_625);
or U1716 (N_1716,N_1159,In_1744);
and U1717 (N_1717,N_292,N_420);
and U1718 (N_1718,N_352,N_817);
xnor U1719 (N_1719,N_1480,In_1956);
nor U1720 (N_1720,N_1425,In_542);
nand U1721 (N_1721,N_943,In_1246);
xor U1722 (N_1722,N_276,N_1256);
nand U1723 (N_1723,N_990,N_160);
nand U1724 (N_1724,In_925,N_312);
and U1725 (N_1725,In_872,N_813);
and U1726 (N_1726,N_1418,N_30);
nand U1727 (N_1727,N_176,N_1042);
or U1728 (N_1728,N_620,In_865);
nand U1729 (N_1729,N_1057,In_293);
and U1730 (N_1730,N_718,N_422);
or U1731 (N_1731,In_2624,N_434);
and U1732 (N_1732,N_708,In_2330);
and U1733 (N_1733,N_1499,In_662);
xnor U1734 (N_1734,N_83,N_738);
or U1735 (N_1735,N_1443,In_306);
nand U1736 (N_1736,In_2987,In_2205);
xor U1737 (N_1737,In_1484,N_902);
xnor U1738 (N_1738,In_1105,N_1464);
and U1739 (N_1739,N_1148,N_880);
xor U1740 (N_1740,In_2141,In_1369);
or U1741 (N_1741,N_664,In_1448);
nand U1742 (N_1742,In_1307,N_1107);
nand U1743 (N_1743,N_1341,N_828);
and U1744 (N_1744,In_1462,In_2039);
or U1745 (N_1745,N_1413,N_1421);
xnor U1746 (N_1746,In_1267,N_1430);
or U1747 (N_1747,In_2664,In_2267);
nor U1748 (N_1748,In_265,In_1681);
nor U1749 (N_1749,In_361,In_2941);
xnor U1750 (N_1750,In_2890,In_2885);
nor U1751 (N_1751,In_2697,N_903);
nand U1752 (N_1752,N_1064,N_212);
xor U1753 (N_1753,In_1868,In_2186);
nor U1754 (N_1754,N_1234,N_1258);
nor U1755 (N_1755,In_1350,N_871);
or U1756 (N_1756,In_2562,In_2658);
and U1757 (N_1757,In_247,N_700);
xor U1758 (N_1758,In_1492,N_645);
and U1759 (N_1759,In_1461,N_744);
and U1760 (N_1760,N_627,N_1236);
or U1761 (N_1761,N_1493,N_1181);
nor U1762 (N_1762,In_2184,In_134);
or U1763 (N_1763,N_634,In_1729);
and U1764 (N_1764,N_1122,In_2764);
nand U1765 (N_1765,N_1301,In_262);
xor U1766 (N_1766,N_785,In_2536);
nor U1767 (N_1767,In_554,N_1260);
nand U1768 (N_1768,N_1437,N_971);
nand U1769 (N_1769,N_924,N_1375);
and U1770 (N_1770,In_2513,N_993);
and U1771 (N_1771,N_1059,In_1701);
xor U1772 (N_1772,In_999,In_1597);
or U1773 (N_1773,In_3,In_2481);
nor U1774 (N_1774,In_639,In_1584);
xor U1775 (N_1775,N_1448,N_559);
nor U1776 (N_1776,N_699,N_866);
nand U1777 (N_1777,N_1340,N_1208);
or U1778 (N_1778,N_921,N_618);
nand U1779 (N_1779,N_1486,N_762);
or U1780 (N_1780,N_1029,N_429);
xor U1781 (N_1781,N_1030,In_1237);
and U1782 (N_1782,In_815,In_1758);
or U1783 (N_1783,N_1010,N_1223);
and U1784 (N_1784,In_1456,N_398);
nor U1785 (N_1785,In_2655,N_814);
or U1786 (N_1786,In_2573,In_932);
xor U1787 (N_1787,N_1298,In_2892);
nor U1788 (N_1788,In_259,In_1819);
nor U1789 (N_1789,In_2841,N_1240);
nand U1790 (N_1790,N_1048,In_2058);
nand U1791 (N_1791,In_1062,N_1041);
nor U1792 (N_1792,In_232,In_2095);
nand U1793 (N_1793,N_804,N_87);
and U1794 (N_1794,In_2350,N_941);
nor U1795 (N_1795,N_1169,N_1268);
xor U1796 (N_1796,In_2147,N_750);
or U1797 (N_1797,N_1211,N_1222);
nor U1798 (N_1798,N_1183,In_709);
xor U1799 (N_1799,In_435,In_1557);
and U1800 (N_1800,N_950,N_497);
xor U1801 (N_1801,N_1628,N_1592);
and U1802 (N_1802,N_1611,N_600);
or U1803 (N_1803,N_1789,N_1686);
and U1804 (N_1804,In_798,N_1522);
nand U1805 (N_1805,N_396,N_1276);
xnor U1806 (N_1806,In_305,N_1292);
nor U1807 (N_1807,N_1531,N_169);
nand U1808 (N_1808,N_228,N_1745);
or U1809 (N_1809,In_2518,N_1355);
nor U1810 (N_1810,N_1743,N_858);
and U1811 (N_1811,N_1459,N_1535);
nand U1812 (N_1812,N_1795,N_1216);
and U1813 (N_1813,N_1683,In_1323);
nand U1814 (N_1814,In_1049,N_1623);
nand U1815 (N_1815,N_1210,N_1605);
xnor U1816 (N_1816,N_1021,In_582);
and U1817 (N_1817,N_1651,N_1371);
nand U1818 (N_1818,N_1569,N_1670);
and U1819 (N_1819,In_286,N_660);
xor U1820 (N_1820,N_845,In_1993);
nor U1821 (N_1821,N_1665,N_522);
nand U1822 (N_1822,N_1062,In_2297);
xnor U1823 (N_1823,N_1618,N_1597);
and U1824 (N_1824,N_1763,N_999);
nor U1825 (N_1825,N_1346,In_1846);
xnor U1826 (N_1826,In_1474,N_109);
nor U1827 (N_1827,N_1420,N_1502);
nor U1828 (N_1828,N_745,In_314);
or U1829 (N_1829,In_2019,N_1290);
and U1830 (N_1830,N_807,In_2128);
or U1831 (N_1831,In_1507,N_1284);
nand U1832 (N_1832,N_1706,In_790);
nor U1833 (N_1833,N_1617,N_1274);
xnor U1834 (N_1834,In_517,N_1560);
xor U1835 (N_1835,In_1877,In_145);
and U1836 (N_1836,N_1677,In_2937);
and U1837 (N_1837,N_570,In_585);
nand U1838 (N_1838,N_682,N_958);
nor U1839 (N_1839,N_1488,N_1282);
nand U1840 (N_1840,In_1999,N_1680);
nand U1841 (N_1841,N_1390,N_1294);
nor U1842 (N_1842,N_1690,N_659);
xor U1843 (N_1843,In_2120,In_267);
and U1844 (N_1844,N_1742,In_1332);
nor U1845 (N_1845,N_1357,N_302);
xor U1846 (N_1846,N_1599,In_2747);
nand U1847 (N_1847,N_1197,N_1018);
nor U1848 (N_1848,N_619,N_33);
and U1849 (N_1849,N_1395,N_922);
nand U1850 (N_1850,N_1215,N_536);
nand U1851 (N_1851,In_841,In_720);
and U1852 (N_1852,N_973,N_1688);
xnor U1853 (N_1853,N_1554,N_1385);
and U1854 (N_1854,In_1592,In_110);
nor U1855 (N_1855,In_369,N_132);
nor U1856 (N_1856,N_1225,N_632);
xor U1857 (N_1857,N_1760,N_1481);
and U1858 (N_1858,N_1409,N_416);
or U1859 (N_1859,N_1286,In_647);
or U1860 (N_1860,N_966,N_1279);
nor U1861 (N_1861,In_701,In_840);
nand U1862 (N_1862,In_2756,N_1691);
and U1863 (N_1863,N_1725,In_2393);
nor U1864 (N_1864,In_152,N_978);
and U1865 (N_1865,N_1175,N_1667);
nor U1866 (N_1866,N_1609,N_1798);
nor U1867 (N_1867,In_1116,N_1559);
and U1868 (N_1868,N_554,N_1703);
nand U1869 (N_1869,In_2313,N_669);
nand U1870 (N_1870,N_1410,N_1408);
xor U1871 (N_1871,In_2901,In_895);
nor U1872 (N_1872,N_1727,N_633);
or U1873 (N_1873,In_1471,N_147);
and U1874 (N_1874,N_844,N_1487);
and U1875 (N_1875,In_345,In_1981);
nor U1876 (N_1876,In_1694,N_1571);
or U1877 (N_1877,N_1085,N_1510);
or U1878 (N_1878,N_892,N_1619);
and U1879 (N_1879,In_5,N_836);
and U1880 (N_1880,N_1335,In_2519);
xor U1881 (N_1881,N_1567,N_1272);
and U1882 (N_1882,N_436,N_1031);
nor U1883 (N_1883,In_138,N_1295);
xor U1884 (N_1884,In_2864,N_500);
and U1885 (N_1885,In_193,N_1668);
nand U1886 (N_1886,N_126,N_833);
and U1887 (N_1887,N_1692,In_162);
nand U1888 (N_1888,N_1506,N_1549);
xor U1889 (N_1889,N_605,In_328);
nand U1890 (N_1890,N_366,N_1217);
nor U1891 (N_1891,N_180,In_315);
nor U1892 (N_1892,N_912,N_1539);
nand U1893 (N_1893,N_1596,N_887);
xor U1894 (N_1894,In_879,In_1618);
nor U1895 (N_1895,In_2645,N_1518);
or U1896 (N_1896,N_386,In_2469);
or U1897 (N_1897,N_341,N_1052);
or U1898 (N_1898,In_2554,N_1634);
and U1899 (N_1899,N_380,N_1152);
and U1900 (N_1900,N_890,N_1257);
nand U1901 (N_1901,N_1514,N_1321);
nor U1902 (N_1902,N_1521,In_698);
and U1903 (N_1903,In_2735,N_462);
xor U1904 (N_1904,N_1358,N_1262);
xnor U1905 (N_1905,N_511,In_2818);
and U1906 (N_1906,N_1528,N_1654);
and U1907 (N_1907,In_1163,In_1303);
xnor U1908 (N_1908,N_944,N_1664);
nor U1909 (N_1909,In_1046,In_1266);
and U1910 (N_1910,In_2228,In_183);
or U1911 (N_1911,In_2859,In_2021);
or U1912 (N_1912,N_1719,In_2473);
nand U1913 (N_1913,In_551,N_1475);
nor U1914 (N_1914,N_515,N_1129);
nand U1915 (N_1915,In_2766,In_272);
or U1916 (N_1916,In_2496,In_868);
nand U1917 (N_1917,N_1423,N_1659);
nor U1918 (N_1918,N_1633,N_1450);
nand U1919 (N_1919,N_1601,N_1350);
nor U1920 (N_1920,N_1333,In_135);
and U1921 (N_1921,N_1604,In_1959);
and U1922 (N_1922,N_1759,In_1494);
nand U1923 (N_1923,N_1422,In_2142);
xnor U1924 (N_1924,N_1174,N_1776);
nor U1925 (N_1925,In_2965,N_1482);
nand U1926 (N_1926,N_1769,N_1626);
or U1927 (N_1927,N_1587,N_122);
or U1928 (N_1928,N_415,N_1792);
and U1929 (N_1929,In_1225,In_610);
or U1930 (N_1930,In_2712,N_1115);
xor U1931 (N_1931,N_778,In_1110);
or U1932 (N_1932,N_983,N_1442);
nand U1933 (N_1933,N_1235,N_1645);
or U1934 (N_1934,In_830,N_969);
or U1935 (N_1935,N_1434,N_574);
xor U1936 (N_1936,N_876,N_1785);
and U1937 (N_1937,N_928,N_1099);
nand U1938 (N_1938,In_2676,In_1677);
nor U1939 (N_1939,N_1527,In_2296);
nand U1940 (N_1940,In_806,In_2066);
nor U1941 (N_1941,N_1332,N_763);
or U1942 (N_1942,N_1782,N_1037);
xnor U1943 (N_1943,N_1356,N_670);
xnor U1944 (N_1944,N_1530,N_1369);
and U1945 (N_1945,N_381,In_1591);
and U1946 (N_1946,In_2371,N_1412);
xnor U1947 (N_1947,N_931,N_1533);
nor U1948 (N_1948,N_1313,N_1641);
and U1949 (N_1949,N_907,N_1453);
xnor U1950 (N_1950,N_483,N_1657);
or U1951 (N_1951,N_1739,N_1490);
or U1952 (N_1952,In_2249,In_2809);
or U1953 (N_1953,N_1768,In_2322);
and U1954 (N_1954,In_1301,N_1362);
xor U1955 (N_1955,In_2833,In_2955);
and U1956 (N_1956,N_1612,N_1104);
nand U1957 (N_1957,In_789,N_653);
and U1958 (N_1958,In_1265,N_803);
nor U1959 (N_1959,N_683,N_1564);
xnor U1960 (N_1960,N_359,In_2446);
nand U1961 (N_1961,N_275,In_1278);
nand U1962 (N_1962,In_1392,In_623);
xnor U1963 (N_1963,N_1024,In_1530);
xor U1964 (N_1964,N_1044,In_2325);
xnor U1965 (N_1965,N_179,N_1687);
or U1966 (N_1966,N_1788,N_1568);
xor U1967 (N_1967,In_2504,N_467);
xnor U1968 (N_1968,N_1050,N_834);
xnor U1969 (N_1969,In_1602,In_1137);
or U1970 (N_1970,N_1756,N_1689);
nor U1971 (N_1971,In_2502,N_86);
or U1972 (N_1972,N_1076,In_438);
and U1973 (N_1973,In_2786,N_1090);
nor U1974 (N_1974,N_419,N_1753);
nor U1975 (N_1975,N_1454,N_1119);
and U1976 (N_1976,N_1555,N_1532);
nor U1977 (N_1977,N_1067,In_1175);
nor U1978 (N_1978,N_519,N_1360);
nand U1979 (N_1979,In_396,N_1643);
xor U1980 (N_1980,In_501,In_2386);
or U1981 (N_1981,N_1775,In_614);
xor U1982 (N_1982,N_508,N_1695);
or U1983 (N_1983,N_1016,N_1003);
nor U1984 (N_1984,In_471,N_1733);
xor U1985 (N_1985,In_2032,N_1625);
nand U1986 (N_1986,N_1019,N_240);
and U1987 (N_1987,N_1310,In_2307);
and U1988 (N_1988,N_1401,In_409);
nor U1989 (N_1989,In_62,N_1548);
or U1990 (N_1990,N_1161,N_509);
or U1991 (N_1991,N_741,In_2768);
or U1992 (N_1992,N_35,N_759);
nand U1993 (N_1993,N_1285,In_2967);
nand U1994 (N_1994,N_20,In_2218);
and U1995 (N_1995,In_188,N_1400);
nand U1996 (N_1996,N_1233,N_1696);
and U1997 (N_1997,N_1590,N_1201);
or U1998 (N_1998,In_231,In_984);
or U1999 (N_1999,N_54,N_1073);
xor U2000 (N_2000,N_1794,In_2248);
and U2001 (N_2001,In_1932,N_1331);
and U2002 (N_2002,In_2538,N_1666);
nand U2003 (N_2003,N_1447,In_2252);
nor U2004 (N_2004,In_763,N_1711);
nand U2005 (N_2005,N_856,N_1675);
and U2006 (N_2006,N_1577,In_2105);
nand U2007 (N_2007,N_1735,N_1730);
and U2008 (N_2008,N_1777,N_1676);
and U2009 (N_2009,In_2417,N_1241);
nand U2010 (N_2010,N_1143,N_1646);
or U2011 (N_2011,N_1383,N_1278);
and U2012 (N_2012,N_1524,In_2808);
and U2013 (N_2013,In_1610,In_573);
nor U2014 (N_2014,N_1586,N_1570);
and U2015 (N_2015,In_2575,N_929);
nand U2016 (N_2016,N_1407,N_1540);
nor U2017 (N_2017,N_913,N_1717);
nand U2018 (N_2018,N_783,N_1007);
and U2019 (N_2019,In_2273,In_1680);
and U2020 (N_2020,In_2159,N_955);
nor U2021 (N_2021,N_1536,N_749);
nor U2022 (N_2022,N_1598,N_1589);
or U2023 (N_2023,In_318,In_1640);
nor U2024 (N_2024,N_1193,In_1526);
nand U2025 (N_2025,In_400,N_1684);
and U2026 (N_2026,N_1519,In_1501);
or U2027 (N_2027,N_1079,N_1757);
and U2028 (N_2028,N_1314,In_2275);
xor U2029 (N_2029,N_1541,In_2480);
nand U2030 (N_2030,N_1610,N_728);
nor U2031 (N_2031,N_12,N_1600);
xnor U2032 (N_2032,In_2877,In_2199);
or U2033 (N_2033,N_936,N_1131);
xor U2034 (N_2034,N_1470,In_2613);
nor U2035 (N_2035,N_265,In_1814);
nand U2036 (N_2036,N_1431,In_463);
or U2037 (N_2037,In_2119,N_1380);
or U2038 (N_2038,N_1673,N_998);
nand U2039 (N_2039,In_2990,N_1563);
nand U2040 (N_2040,N_1572,N_1653);
xor U2041 (N_2041,In_2963,In_1459);
xnor U2042 (N_2042,N_1671,In_478);
nor U2043 (N_2043,N_1127,N_1515);
xnor U2044 (N_2044,N_136,N_1652);
and U2045 (N_2045,N_1551,In_2976);
nand U2046 (N_2046,N_1747,N_1588);
or U2047 (N_2047,N_1765,N_963);
or U2048 (N_2048,N_1382,N_1751);
and U2049 (N_2049,N_1312,In_485);
nor U2050 (N_2050,N_665,N_1255);
or U2051 (N_2051,N_1774,N_210);
nor U2052 (N_2052,N_516,In_1355);
nor U2053 (N_2053,N_1428,N_1138);
nand U2054 (N_2054,N_1663,N_1494);
and U2055 (N_2055,N_1153,N_681);
xor U2056 (N_2056,N_1699,N_114);
and U2057 (N_2057,In_1438,N_649);
and U2058 (N_2058,N_118,N_1543);
nor U2059 (N_2059,In_2636,N_1483);
nor U2060 (N_2060,N_1649,In_2137);
and U2061 (N_2061,N_1584,N_1102);
xor U2062 (N_2062,In_1730,N_1009);
or U2063 (N_2063,In_2705,In_2781);
or U2064 (N_2064,In_632,In_493);
or U2065 (N_2065,N_1329,N_534);
nor U2066 (N_2066,N_8,In_1630);
xor U2067 (N_2067,N_1749,N_233);
or U2068 (N_2068,N_724,In_1617);
or U2069 (N_2069,N_1446,N_1230);
xor U2070 (N_2070,In_2525,N_1758);
nand U2071 (N_2071,N_1155,N_1701);
and U2072 (N_2072,N_197,N_1779);
nand U2073 (N_2073,In_108,N_321);
nand U2074 (N_2074,N_1658,In_1394);
xnor U2075 (N_2075,In_524,N_1238);
or U2076 (N_2076,In_2543,N_1270);
nand U2077 (N_2077,N_1661,In_2974);
nor U2078 (N_2078,In_10,N_300);
xnor U2079 (N_2079,N_1752,N_447);
and U2080 (N_2080,N_1616,In_825);
xor U2081 (N_2081,N_1040,In_2388);
nor U2082 (N_2082,In_1808,In_2537);
xnor U2083 (N_2083,N_1330,N_1178);
nor U2084 (N_2084,In_2221,N_1126);
or U2085 (N_2085,In_142,In_245);
or U2086 (N_2086,In_462,N_651);
nand U2087 (N_2087,In_620,N_1615);
nor U2088 (N_2088,In_2462,N_1117);
xnor U2089 (N_2089,N_1698,N_374);
or U2090 (N_2090,N_1396,In_654);
nand U2091 (N_2091,N_601,N_1269);
xor U2092 (N_2092,N_1150,N_1170);
and U2093 (N_2093,N_1582,In_2123);
and U2094 (N_2094,N_266,In_2983);
nor U2095 (N_2095,In_1187,N_1558);
or U2096 (N_2096,N_384,N_471);
nand U2097 (N_2097,N_1738,In_631);
and U2098 (N_2098,N_1712,N_1744);
xor U2099 (N_2099,N_1580,In_1687);
and U2100 (N_2100,N_1444,N_1839);
nand U2101 (N_2101,N_2038,N_1553);
nand U2102 (N_2102,N_1724,N_1960);
nor U2103 (N_2103,N_1296,N_1996);
xnor U2104 (N_2104,N_1202,N_1904);
nand U2105 (N_2105,In_2620,N_1022);
nand U2106 (N_2106,In_1047,N_1838);
xnor U2107 (N_2107,N_1566,N_1352);
xnor U2108 (N_2108,N_680,N_1503);
nand U2109 (N_2109,In_1336,N_1479);
and U2110 (N_2110,N_329,In_1015);
or U2111 (N_2111,N_1644,N_1557);
nor U2112 (N_2112,N_1583,N_2030);
xor U2113 (N_2113,N_2070,N_244);
and U2114 (N_2114,N_1803,N_2005);
nand U2115 (N_2115,In_1497,N_1198);
nor U2116 (N_2116,In_1712,In_2722);
nand U2117 (N_2117,N_1840,In_2995);
xnor U2118 (N_2118,N_1778,N_2071);
nand U2119 (N_2119,N_1846,N_1831);
or U2120 (N_2120,N_850,N_790);
nor U2121 (N_2121,N_1916,In_2336);
xor U2122 (N_2122,N_2076,N_1809);
or U2123 (N_2123,In_769,N_99);
xor U2124 (N_2124,N_1565,N_1704);
nand U2125 (N_2125,N_1998,N_1498);
or U2126 (N_2126,N_1534,N_2063);
or U2127 (N_2127,N_393,N_1941);
or U2128 (N_2128,N_1964,N_1517);
xnor U2129 (N_2129,N_964,In_1198);
nor U2130 (N_2130,In_27,N_1812);
nor U2131 (N_2131,N_456,N_1949);
nand U2132 (N_2132,In_1179,N_1974);
or U2133 (N_2133,N_1715,In_1954);
nor U2134 (N_2134,N_2057,N_1800);
and U2135 (N_2135,N_1837,N_1134);
or U2136 (N_2136,In_1783,N_1955);
nor U2137 (N_2137,In_2293,N_1877);
xor U2138 (N_2138,In_1409,N_831);
nor U2139 (N_2139,N_1489,N_1245);
or U2140 (N_2140,In_1986,N_1709);
and U2141 (N_2141,N_1970,In_1281);
and U2142 (N_2142,In_1450,N_2064);
nand U2143 (N_2143,N_1905,N_1948);
and U2144 (N_2144,N_1863,In_2016);
nand U2145 (N_2145,N_408,In_1481);
or U2146 (N_2146,In_1984,N_1397);
and U2147 (N_2147,N_1440,N_1376);
or U2148 (N_2148,In_2550,N_1907);
nor U2149 (N_2149,In_2476,N_1754);
nand U2150 (N_2150,In_274,N_1726);
nor U2151 (N_2151,N_1869,N_1836);
or U2152 (N_2152,In_1408,N_1811);
nand U2153 (N_2153,N_1880,N_1550);
and U2154 (N_2154,N_2023,N_2042);
or U2155 (N_2155,N_1516,N_1716);
xor U2156 (N_2156,N_199,N_1975);
nor U2157 (N_2157,N_1906,N_985);
or U2158 (N_2158,N_662,N_1821);
nand U2159 (N_2159,N_1114,N_1908);
xnor U2160 (N_2160,N_1856,N_1624);
and U2161 (N_2161,N_1622,N_1354);
xnor U2162 (N_2162,N_1801,N_1457);
or U2163 (N_2163,N_1992,In_2758);
and U2164 (N_2164,N_1304,N_1844);
nor U2165 (N_2165,N_1116,In_1043);
or U2166 (N_2166,N_1607,N_1594);
xor U2167 (N_2167,N_756,N_873);
nor U2168 (N_2168,N_1714,N_1165);
and U2169 (N_2169,N_1468,N_296);
xor U2170 (N_2170,N_1918,N_1982);
xor U2171 (N_2171,N_1919,In_133);
xor U2172 (N_2172,N_1191,N_2029);
xor U2173 (N_2173,N_1849,N_1870);
or U2174 (N_2174,In_2333,In_2430);
nor U2175 (N_2175,In_271,N_2079);
nand U2176 (N_2176,N_624,N_2008);
xor U2177 (N_2177,N_2036,N_1456);
or U2178 (N_2178,In_2131,N_1780);
or U2179 (N_2179,In_2328,N_2098);
xnor U2180 (N_2180,N_42,In_914);
nand U2181 (N_2181,N_1705,In_71);
nor U2182 (N_2182,N_1988,N_1741);
nand U2183 (N_2183,N_1816,N_1755);
nand U2184 (N_2184,N_2020,N_1231);
or U2185 (N_2185,N_1886,N_1993);
nor U2186 (N_2186,In_1483,N_1942);
nand U2187 (N_2187,In_2488,In_1502);
nor U2188 (N_2188,N_1342,N_90);
nand U2189 (N_2189,N_1614,In_1324);
xor U2190 (N_2190,In_671,N_2016);
nor U2191 (N_2191,N_1348,N_1347);
or U2192 (N_2192,N_2091,N_1945);
nor U2193 (N_2193,N_2026,N_1636);
and U2194 (N_2194,N_1608,N_979);
and U2195 (N_2195,N_1656,N_1545);
nor U2196 (N_2196,N_545,N_413);
xnor U2197 (N_2197,In_2366,N_1635);
and U2198 (N_2198,In_191,N_1936);
nand U2199 (N_2199,N_1921,N_1884);
nand U2200 (N_2200,N_1185,N_1186);
or U2201 (N_2201,N_1497,N_2022);
and U2202 (N_2202,N_1933,In_1378);
nor U2203 (N_2203,N_2049,N_1983);
nand U2204 (N_2204,N_2003,N_1072);
nor U2205 (N_2205,N_1491,N_1061);
nor U2206 (N_2206,N_1306,In_1425);
or U2207 (N_2207,N_1950,N_1237);
and U2208 (N_2208,N_2072,In_2578);
nand U2209 (N_2209,N_563,N_1365);
and U2210 (N_2210,N_2089,N_948);
nor U2211 (N_2211,N_1386,In_1259);
xor U2212 (N_2212,N_595,In_1717);
xor U2213 (N_2213,N_1377,In_2854);
and U2214 (N_2214,N_1969,N_1319);
or U2215 (N_2215,N_1899,N_1261);
and U2216 (N_2216,N_1372,In_808);
or U2217 (N_2217,In_1177,In_1310);
nand U2218 (N_2218,N_1326,N_1281);
or U2219 (N_2219,N_949,N_1925);
xor U2220 (N_2220,N_974,In_2923);
nand U2221 (N_2221,N_1784,N_142);
nand U2222 (N_2222,In_1407,N_616);
and U2223 (N_2223,In_1949,N_1639);
xor U2224 (N_2224,N_1300,In_2428);
and U2225 (N_2225,N_2031,N_1814);
or U2226 (N_2226,N_1790,N_1962);
and U2227 (N_2227,N_1602,In_153);
or U2228 (N_2228,N_1834,N_1987);
xor U2229 (N_2229,N_1184,N_945);
and U2230 (N_2230,N_335,N_1817);
xor U2231 (N_2231,In_302,In_2078);
and U2232 (N_2232,N_1909,In_67);
and U2233 (N_2233,N_1209,N_1526);
xnor U2234 (N_2234,N_2006,N_1648);
and U2235 (N_2235,In_1735,N_2062);
or U2236 (N_2236,N_766,N_2033);
nor U2237 (N_2237,N_2028,In_753);
and U2238 (N_2238,In_923,N_262);
nand U2239 (N_2239,In_1638,N_1896);
or U2240 (N_2240,N_1890,In_1227);
or U2241 (N_2241,N_938,N_1125);
and U2242 (N_2242,In_1400,N_1394);
nor U2243 (N_2243,In_1054,N_1384);
nand U2244 (N_2244,In_1912,N_1928);
and U2245 (N_2245,N_1958,In_949);
or U2246 (N_2246,N_1512,N_2019);
nand U2247 (N_2247,N_1843,In_1537);
or U2248 (N_2248,In_1252,N_1581);
nor U2249 (N_2249,N_1318,N_1729);
or U2250 (N_2250,N_1842,N_1943);
xnor U2251 (N_2251,N_1630,N_1647);
nor U2252 (N_2252,N_1832,N_2021);
and U2253 (N_2253,N_1999,N_1953);
nand U2254 (N_2254,N_1111,N_1473);
nor U2255 (N_2255,In_1247,N_1157);
or U2256 (N_2256,In_2038,N_493);
and U2257 (N_2257,N_2082,N_1852);
nor U2258 (N_2258,In_951,N_602);
nor U2259 (N_2259,N_1866,N_1087);
nand U2260 (N_2260,In_1926,N_1097);
or U2261 (N_2261,N_1511,N_1026);
or U2262 (N_2262,In_2853,N_1961);
nand U2263 (N_2263,N_1315,N_1824);
xor U2264 (N_2264,In_2848,In_2390);
xor U2265 (N_2265,N_1101,N_1980);
xnor U2266 (N_2266,N_930,N_920);
nand U2267 (N_2267,N_1721,N_919);
and U2268 (N_2268,N_2058,In_1390);
and U2269 (N_2269,N_2010,N_1967);
or U2270 (N_2270,N_1154,In_1027);
and U2271 (N_2271,N_2040,N_1973);
nand U2272 (N_2272,N_1930,N_648);
nor U2273 (N_2273,In_1832,In_1275);
xor U2274 (N_2274,N_1959,N_881);
nor U2275 (N_2275,In_2173,In_312);
nand U2276 (N_2276,N_1011,In_2433);
nor U2277 (N_2277,N_714,N_1806);
and U2278 (N_2278,In_650,N_1954);
and U2279 (N_2279,N_370,N_1708);
or U2280 (N_2280,In_115,N_775);
xnor U2281 (N_2281,N_897,N_1881);
or U2282 (N_2282,N_2090,In_2773);
xnor U2283 (N_2283,N_1766,N_1947);
nand U2284 (N_2284,N_1914,N_776);
nor U2285 (N_2285,N_1417,N_1537);
or U2286 (N_2286,N_1818,N_2051);
nor U2287 (N_2287,N_1485,N_1344);
nand U2288 (N_2288,N_830,In_241);
xor U2289 (N_2289,N_2045,N_1786);
nor U2290 (N_2290,N_1323,N_1860);
or U2291 (N_2291,N_1620,N_1366);
nand U2292 (N_2292,In_2733,N_1561);
nand U2293 (N_2293,N_1046,In_1616);
nor U2294 (N_2294,N_666,N_1872);
nor U2295 (N_2295,In_875,In_2034);
xor U2296 (N_2296,In_818,N_1203);
and U2297 (N_2297,In_734,N_1915);
nor U2298 (N_2298,N_1938,N_723);
nor U2299 (N_2299,In_1988,N_1414);
or U2300 (N_2300,N_1133,In_460);
and U2301 (N_2301,In_2040,N_2099);
nand U2302 (N_2302,In_1850,N_693);
nor U2303 (N_2303,In_359,N_1182);
nor U2304 (N_2304,N_1469,N_1547);
nor U2305 (N_2305,N_1433,N_2055);
nand U2306 (N_2306,In_1403,N_1173);
nand U2307 (N_2307,N_1638,N_1416);
or U2308 (N_2308,N_521,N_2011);
or U2309 (N_2309,N_953,N_1764);
xor U2310 (N_2310,N_261,N_1833);
nor U2311 (N_2311,N_1823,N_1351);
nor U2312 (N_2312,N_1868,N_1951);
nor U2313 (N_2313,N_1934,N_910);
nor U2314 (N_2314,N_1681,N_1682);
or U2315 (N_2315,In_22,N_2004);
and U2316 (N_2316,N_555,N_2001);
nor U2317 (N_2317,N_1585,In_428);
and U2318 (N_2318,N_2086,In_1078);
nor U2319 (N_2319,N_1807,N_1897);
nand U2320 (N_2320,N_1864,N_2000);
nand U2321 (N_2321,In_1235,N_1805);
xor U2322 (N_2322,N_2009,N_1576);
nor U2323 (N_2323,N_1781,In_1470);
xnor U2324 (N_2324,N_717,N_1466);
nor U2325 (N_2325,N_1693,N_1650);
nor U2326 (N_2326,N_1815,N_2017);
and U2327 (N_2327,N_2068,N_249);
or U2328 (N_2328,In_661,N_894);
nand U2329 (N_2329,N_1761,N_94);
or U2330 (N_2330,N_1989,In_1539);
and U2331 (N_2331,In_1807,N_2034);
nand U2332 (N_2332,N_1929,N_2081);
xnor U2333 (N_2333,In_2860,N_252);
nor U2334 (N_2334,N_1642,N_1893);
or U2335 (N_2335,N_411,N_490);
or U2336 (N_2336,N_2037,N_2092);
nor U2337 (N_2337,In_1173,N_1674);
nand U2338 (N_2338,N_1509,N_1593);
or U2339 (N_2339,N_1937,N_1804);
nor U2340 (N_2340,N_1848,N_1700);
xor U2341 (N_2341,N_1132,N_1939);
or U2342 (N_2342,N_1902,In_1994);
xor U2343 (N_2343,N_2027,N_1068);
nand U2344 (N_2344,N_2069,In_1637);
nor U2345 (N_2345,N_1051,N_1986);
or U2346 (N_2346,N_1971,In_1475);
and U2347 (N_2347,N_1513,N_2056);
xnor U2348 (N_2348,N_1722,N_1);
and U2349 (N_2349,N_333,In_2956);
or U2350 (N_2350,N_1520,N_167);
and U2351 (N_2351,In_1820,N_1917);
or U2352 (N_2352,In_1696,N_1891);
or U2353 (N_2353,N_2012,N_1573);
and U2354 (N_2354,N_1629,N_1501);
and U2355 (N_2355,N_1484,N_1799);
xnor U2356 (N_2356,In_2698,N_789);
xor U2357 (N_2357,In_229,N_1994);
or U2358 (N_2358,N_599,N_1885);
nor U2359 (N_2359,N_1544,In_1490);
nor U2360 (N_2360,N_1637,N_2080);
nor U2361 (N_2361,N_1139,In_118);
nand U2362 (N_2362,N_1963,N_1591);
nor U2363 (N_2363,In_2013,In_2045);
nor U2364 (N_2364,N_1275,N_1750);
xor U2365 (N_2365,In_770,N_1810);
nand U2366 (N_2366,N_1226,In_1686);
and U2367 (N_2367,In_1104,N_1196);
nor U2368 (N_2368,N_1740,N_767);
nor U2369 (N_2369,In_708,N_2025);
nor U2370 (N_2370,N_1851,N_1662);
and U2371 (N_2371,N_203,In_2511);
nor U2372 (N_2372,N_1746,N_1640);
xor U2373 (N_2373,In_674,N_1271);
nor U2374 (N_2374,N_1911,In_1016);
and U2375 (N_2375,N_1845,N_1927);
nand U2376 (N_2376,In_1649,N_1793);
nor U2377 (N_2377,In_2111,N_1091);
and U2378 (N_2378,N_968,N_526);
or U2379 (N_2379,N_1595,N_792);
xor U2380 (N_2380,In_2165,In_1217);
nand U2381 (N_2381,N_2096,N_232);
nor U2382 (N_2382,N_2061,N_1865);
nand U2383 (N_2383,In_1309,N_1808);
or U2384 (N_2384,In_1580,N_1874);
or U2385 (N_2385,N_939,N_1146);
or U2386 (N_2386,N_1830,In_70);
nand U2387 (N_2387,N_2007,N_1841);
nand U2388 (N_2388,In_1322,In_1689);
nand U2389 (N_2389,In_1464,N_752);
nor U2390 (N_2390,In_1566,N_2067);
xor U2391 (N_2391,N_1305,N_1391);
or U2392 (N_2392,N_1718,N_412);
nor U2393 (N_2393,N_2032,N_2078);
nand U2394 (N_2394,In_2380,In_1168);
nand U2395 (N_2395,N_1578,N_1966);
or U2396 (N_2396,N_1940,N_1952);
or U2397 (N_2397,N_1737,N_1552);
nor U2398 (N_2398,N_1529,N_2077);
and U2399 (N_2399,N_1828,In_1234);
nand U2400 (N_2400,N_2074,N_2278);
xnor U2401 (N_2401,N_1748,N_2174);
xnor U2402 (N_2402,N_1888,N_1728);
and U2403 (N_2403,N_1627,N_2340);
xor U2404 (N_2404,N_2161,N_440);
and U2405 (N_2405,In_124,N_855);
nand U2406 (N_2406,N_1538,In_776);
and U2407 (N_2407,N_2313,N_1773);
nand U2408 (N_2408,N_2154,In_408);
or U2409 (N_2409,N_2211,N_2139);
nand U2410 (N_2410,N_2275,N_2263);
xor U2411 (N_2411,N_1546,N_989);
xnor U2412 (N_2412,N_1827,N_2163);
and U2413 (N_2413,N_1697,N_2052);
and U2414 (N_2414,N_1979,N_1452);
or U2415 (N_2415,N_1505,N_1206);
nor U2416 (N_2416,N_1308,N_2272);
and U2417 (N_2417,N_1889,N_2054);
nor U2418 (N_2418,N_2230,N_1495);
and U2419 (N_2419,N_1802,N_1857);
xor U2420 (N_2420,N_1685,N_2227);
xnor U2421 (N_2421,N_617,N_1990);
nand U2422 (N_2422,N_2323,In_1508);
and U2423 (N_2423,N_1900,N_1694);
and U2424 (N_2424,N_2150,N_2359);
nor U2425 (N_2425,N_2267,In_1029);
xnor U2426 (N_2426,N_1349,N_586);
xor U2427 (N_2427,N_1669,N_2083);
or U2428 (N_2428,N_1935,N_753);
or U2429 (N_2429,N_2186,N_2237);
nand U2430 (N_2430,N_279,N_2308);
or U2431 (N_2431,N_1474,N_535);
or U2432 (N_2432,N_224,N_1772);
and U2433 (N_2433,N_2367,N_1820);
nor U2434 (N_2434,In_323,In_2815);
xnor U2435 (N_2435,N_1504,N_1095);
nor U2436 (N_2436,N_2286,N_2046);
xor U2437 (N_2437,N_1862,N_1034);
nor U2438 (N_2438,N_2357,N_1106);
nor U2439 (N_2439,N_1556,N_2260);
and U2440 (N_2440,N_2247,N_2118);
nor U2441 (N_2441,N_2382,N_947);
nor U2442 (N_2442,N_2132,N_1825);
nand U2443 (N_2443,N_2379,In_1341);
nand U2444 (N_2444,N_1214,N_2166);
or U2445 (N_2445,N_2130,N_2370);
nor U2446 (N_2446,N_2351,N_2141);
and U2447 (N_2447,N_1419,N_1910);
nand U2448 (N_2448,N_241,N_1508);
xnor U2449 (N_2449,In_2949,N_2330);
xnor U2450 (N_2450,N_2144,N_2183);
and U2451 (N_2451,N_2344,N_2238);
nor U2452 (N_2452,N_2122,In_2174);
and U2453 (N_2453,N_1100,N_1932);
nand U2454 (N_2454,N_1813,N_2371);
and U2455 (N_2455,In_1370,N_2354);
nand U2456 (N_2456,N_2116,N_1858);
or U2457 (N_2457,N_1562,N_2264);
or U2458 (N_2458,N_2172,N_2281);
nor U2459 (N_2459,In_370,N_918);
nor U2460 (N_2460,N_2232,N_2196);
and U2461 (N_2461,N_1613,N_2372);
nand U2462 (N_2462,N_2266,N_1926);
xor U2463 (N_2463,N_2321,N_2366);
or U2464 (N_2464,N_2121,N_2242);
xor U2465 (N_2465,N_1879,N_2383);
or U2466 (N_2466,In_1529,In_2830);
and U2467 (N_2467,N_2293,N_2035);
nand U2468 (N_2468,N_2066,N_2131);
xor U2469 (N_2469,N_2393,N_2255);
nor U2470 (N_2470,N_2059,N_2295);
xnor U2471 (N_2471,N_932,N_587);
xnor U2472 (N_2472,N_1575,N_1039);
nor U2473 (N_2473,In_2629,N_2104);
xnor U2474 (N_2474,N_2223,N_2041);
or U2475 (N_2475,N_2214,N_2151);
nor U2476 (N_2476,N_2322,N_2390);
nand U2477 (N_2477,N_2360,N_2363);
xnor U2478 (N_2478,N_746,N_2169);
or U2479 (N_2479,N_2053,N_2252);
or U2480 (N_2480,N_2369,N_1991);
xor U2481 (N_2481,N_2348,N_1895);
nand U2482 (N_2482,In_1517,In_1420);
nor U2483 (N_2483,N_2332,N_2145);
xor U2484 (N_2484,N_2365,N_1542);
xnor U2485 (N_2485,N_2125,N_2297);
nand U2486 (N_2486,In_2657,N_2270);
xnor U2487 (N_2487,N_933,N_2375);
nor U2488 (N_2488,In_933,N_2094);
or U2489 (N_2489,N_2338,N_1875);
xnor U2490 (N_2490,N_2229,N_2342);
nor U2491 (N_2491,N_2381,N_1723);
nand U2492 (N_2492,N_2129,N_2105);
nor U2493 (N_2493,N_1923,N_2327);
nand U2494 (N_2494,N_2362,N_2251);
or U2495 (N_2495,N_1867,N_2084);
and U2496 (N_2496,N_2356,In_2247);
or U2497 (N_2497,N_1876,N_2294);
and U2498 (N_2498,N_1445,N_2050);
and U2499 (N_2499,N_2138,N_937);
and U2500 (N_2500,N_2093,N_2198);
and U2501 (N_2501,N_2111,N_1702);
xor U2502 (N_2502,N_2268,N_2135);
and U2503 (N_2503,N_2143,N_2222);
and U2504 (N_2504,N_1859,N_2220);
xor U2505 (N_2505,N_2326,N_2218);
xor U2506 (N_2506,N_2065,N_2194);
xnor U2507 (N_2507,N_2142,N_2103);
xnor U2508 (N_2508,N_2221,N_2216);
or U2509 (N_2509,In_1611,N_2231);
nor U2510 (N_2510,N_1579,In_1660);
or U2511 (N_2511,N_1977,N_2347);
xnor U2512 (N_2512,N_1337,N_1901);
and U2513 (N_2513,N_1606,N_2107);
xnor U2514 (N_2514,N_2289,N_2155);
or U2515 (N_2515,N_1322,N_2088);
and U2516 (N_2516,N_1878,N_11);
and U2517 (N_2517,N_848,N_2269);
nand U2518 (N_2518,N_1713,N_2208);
nor U2519 (N_2519,N_2178,N_1855);
or U2520 (N_2520,N_2292,N_2241);
or U2521 (N_2521,In_164,N_1345);
nor U2522 (N_2522,N_2047,N_1212);
and U2523 (N_2523,N_2179,N_2180);
or U2524 (N_2524,N_2235,N_153);
and U2525 (N_2525,N_2378,In_2363);
nand U2526 (N_2526,N_2244,N_2243);
and U2527 (N_2527,N_2245,N_2336);
xnor U2528 (N_2528,N_2337,N_1892);
xnor U2529 (N_2529,N_2282,In_1331);
and U2530 (N_2530,In_199,N_542);
or U2531 (N_2531,N_2246,N_1981);
or U2532 (N_2532,N_2259,N_2133);
and U2533 (N_2533,N_2291,In_2130);
nor U2534 (N_2534,N_2306,N_2152);
or U2535 (N_2535,N_2262,N_2182);
or U2536 (N_2536,N_1339,N_2397);
nand U2537 (N_2537,N_1311,N_2140);
or U2538 (N_2538,In_2970,N_2325);
and U2539 (N_2539,N_2239,N_1439);
xnor U2540 (N_2540,N_2044,N_541);
nor U2541 (N_2541,N_2395,N_2346);
or U2542 (N_2542,N_2361,N_2276);
nand U2543 (N_2543,N_2157,N_1767);
nor U2544 (N_2544,N_2097,In_2453);
or U2545 (N_2545,N_2102,N_2335);
nor U2546 (N_2546,N_1882,N_2331);
nor U2547 (N_2547,N_1791,N_2324);
nand U2548 (N_2548,N_1770,N_2167);
nor U2549 (N_2549,N_2358,N_2317);
or U2550 (N_2550,In_1315,N_1033);
xnor U2551 (N_2551,N_2181,N_2373);
xnor U2552 (N_2552,N_2316,N_734);
nor U2553 (N_2553,In_1067,N_2279);
and U2554 (N_2554,N_2043,N_1679);
nand U2555 (N_2555,N_2318,N_2018);
nor U2556 (N_2556,N_2380,N_2250);
and U2557 (N_2557,N_2085,N_1984);
or U2558 (N_2558,N_2160,N_1621);
nand U2559 (N_2559,In_2254,N_1995);
or U2560 (N_2560,In_1346,N_2101);
xnor U2561 (N_2561,In_1836,N_1965);
xnor U2562 (N_2562,N_748,N_1289);
and U2563 (N_2563,N_2117,N_721);
or U2564 (N_2564,N_1239,N_2193);
nor U2565 (N_2565,N_2201,N_2328);
or U2566 (N_2566,N_2368,In_958);
nor U2567 (N_2567,N_896,N_2024);
nand U2568 (N_2568,N_1660,N_2320);
nand U2569 (N_2569,N_1736,N_2014);
nor U2570 (N_2570,N_1731,N_2396);
nor U2571 (N_2571,N_2341,N_2234);
xnor U2572 (N_2572,N_2389,N_2333);
nor U2573 (N_2573,N_2120,N_1946);
xnor U2574 (N_2574,N_2203,N_1435);
xor U2575 (N_2575,N_2128,N_2177);
nand U2576 (N_2576,N_2146,N_2307);
and U2577 (N_2577,N_1732,In_1172);
nand U2578 (N_2578,N_1204,N_2205);
or U2579 (N_2579,N_2219,N_1887);
and U2580 (N_2580,N_1922,N_2388);
xor U2581 (N_2581,In_2260,In_2037);
nor U2582 (N_2582,In_2022,In_2235);
nor U2583 (N_2583,N_2249,N_2349);
xnor U2584 (N_2584,N_2265,N_1972);
and U2585 (N_2585,In_2777,N_1655);
or U2586 (N_2586,N_2213,N_2100);
or U2587 (N_2587,N_2303,In_658);
xor U2588 (N_2588,N_2285,N_2185);
and U2589 (N_2589,N_2187,N_2287);
xnor U2590 (N_2590,In_2936,N_1213);
nor U2591 (N_2591,N_2299,N_1797);
nand U2592 (N_2592,N_2304,N_2253);
nor U2593 (N_2593,N_1920,N_2153);
xor U2594 (N_2594,N_1957,N_2197);
or U2595 (N_2595,N_1847,N_2184);
nor U2596 (N_2596,N_1251,N_1672);
xnor U2597 (N_2597,N_1873,N_2314);
nand U2598 (N_2598,N_1603,N_2110);
nand U2599 (N_2599,N_1796,N_306);
xor U2600 (N_2600,N_1404,N_2164);
xor U2601 (N_2601,N_2204,N_2191);
nor U2602 (N_2602,N_2039,N_2217);
or U2603 (N_2603,N_1392,N_2127);
nor U2604 (N_2604,N_2114,In_1124);
and U2605 (N_2605,N_2195,N_49);
nor U2606 (N_2606,N_2060,N_353);
nand U2607 (N_2607,N_2329,N_657);
xor U2608 (N_2608,N_2106,N_2176);
nand U2609 (N_2609,N_2392,N_1574);
and U2610 (N_2610,N_2199,N_1194);
and U2611 (N_2611,N_960,N_2170);
nand U2612 (N_2612,N_2256,N_2352);
xor U2613 (N_2613,N_2394,N_1861);
nor U2614 (N_2614,N_2048,N_1850);
xnor U2615 (N_2615,N_2206,N_428);
and U2616 (N_2616,N_1997,In_1971);
and U2617 (N_2617,In_1091,N_2345);
xor U2618 (N_2618,N_2073,N_2280);
nor U2619 (N_2619,N_2283,N_2188);
and U2620 (N_2620,N_2355,N_2148);
and U2621 (N_2621,N_2386,N_1968);
or U2622 (N_2622,N_2305,N_2192);
xor U2623 (N_2623,N_1883,N_2126);
or U2624 (N_2624,In_807,N_1771);
or U2625 (N_2625,In_99,N_182);
nand U2626 (N_2626,In_941,N_1523);
nand U2627 (N_2627,N_2296,N_2168);
xor U2628 (N_2628,N_2202,N_2136);
xnor U2629 (N_2629,N_1976,In_491);
nand U2630 (N_2630,N_1822,N_2190);
and U2631 (N_2631,N_2311,N_1720);
xnor U2632 (N_2632,In_2190,N_2261);
xnor U2633 (N_2633,N_2288,N_2257);
or U2634 (N_2634,N_2258,N_1854);
nand U2635 (N_2635,N_2209,N_2309);
nor U2636 (N_2636,In_2721,N_679);
xnor U2637 (N_2637,N_2387,N_2290);
xor U2638 (N_2638,In_1847,In_1606);
nand U2639 (N_2639,In_1568,N_2087);
xor U2640 (N_2640,N_2159,N_1835);
nand U2641 (N_2641,N_2149,N_2399);
nand U2642 (N_2642,N_2124,N_2384);
nor U2643 (N_2643,N_242,N_1500);
nand U2644 (N_2644,N_2233,N_2212);
and U2645 (N_2645,N_2240,N_2385);
and U2646 (N_2646,N_2343,In_2943);
xnor U2647 (N_2647,In_1103,N_1254);
nor U2648 (N_2648,N_2075,N_2119);
or U2649 (N_2649,N_1829,N_2113);
nand U2650 (N_2650,N_1406,N_2002);
or U2651 (N_2651,In_1519,N_1787);
xor U2652 (N_2652,N_2226,N_484);
nor U2653 (N_2653,N_2236,N_2189);
xnor U2654 (N_2654,N_2319,N_2228);
nor U2655 (N_2655,N_2391,N_2175);
or U2656 (N_2656,N_1985,N_2200);
nand U2657 (N_2657,N_2109,N_1267);
xor U2658 (N_2658,N_1826,N_1525);
nand U2659 (N_2659,In_2323,N_1188);
and U2660 (N_2660,N_1944,N_2224);
xnor U2661 (N_2661,N_2147,N_2173);
nor U2662 (N_2662,N_1734,N_2376);
nand U2663 (N_2663,In_1363,N_2225);
xor U2664 (N_2664,In_375,N_360);
or U2665 (N_2665,N_2377,N_2248);
nor U2666 (N_2666,N_2210,N_2254);
nand U2667 (N_2667,N_2312,N_1783);
nor U2668 (N_2668,N_2350,N_2207);
or U2669 (N_2669,N_2298,N_2112);
nor U2670 (N_2670,N_2301,N_2013);
and U2671 (N_2671,N_1913,N_1912);
or U2672 (N_2672,N_1762,In_1821);
xnor U2673 (N_2673,N_2158,N_2374);
or U2674 (N_2674,N_2315,N_1978);
xor U2675 (N_2675,N_1871,N_2310);
nor U2676 (N_2676,N_2137,N_1956);
nand U2677 (N_2677,N_2284,N_754);
nand U2678 (N_2678,N_1707,In_433);
and U2679 (N_2679,N_2273,N_1894);
nand U2680 (N_2680,In_236,N_1898);
xor U2681 (N_2681,N_2134,N_1631);
nor U2682 (N_2682,N_1632,N_2274);
or U2683 (N_2683,N_2156,N_2015);
or U2684 (N_2684,In_1695,In_719);
nand U2685 (N_2685,N_2165,N_2277);
xnor U2686 (N_2686,N_2162,N_2108);
and U2687 (N_2687,N_1924,N_2123);
and U2688 (N_2688,N_1710,N_2353);
nor U2689 (N_2689,In_2422,N_1507);
nand U2690 (N_2690,N_2339,N_2271);
xor U2691 (N_2691,N_2171,N_2115);
nor U2692 (N_2692,N_283,N_2302);
or U2693 (N_2693,N_2364,N_1853);
xnor U2694 (N_2694,N_2215,N_2334);
xor U2695 (N_2695,N_1931,N_2398);
or U2696 (N_2696,N_1478,N_2095);
nand U2697 (N_2697,N_1903,N_89);
or U2698 (N_2698,N_1678,N_1819);
nor U2699 (N_2699,N_2300,N_474);
xnor U2700 (N_2700,N_2438,N_2622);
or U2701 (N_2701,N_2568,N_2515);
nand U2702 (N_2702,N_2592,N_2558);
nand U2703 (N_2703,N_2452,N_2435);
nand U2704 (N_2704,N_2544,N_2470);
and U2705 (N_2705,N_2425,N_2522);
or U2706 (N_2706,N_2514,N_2698);
and U2707 (N_2707,N_2513,N_2631);
xnor U2708 (N_2708,N_2647,N_2693);
and U2709 (N_2709,N_2623,N_2617);
or U2710 (N_2710,N_2492,N_2696);
nor U2711 (N_2711,N_2599,N_2535);
and U2712 (N_2712,N_2642,N_2468);
nor U2713 (N_2713,N_2602,N_2684);
nor U2714 (N_2714,N_2585,N_2621);
nand U2715 (N_2715,N_2507,N_2628);
and U2716 (N_2716,N_2675,N_2538);
nand U2717 (N_2717,N_2671,N_2660);
xor U2718 (N_2718,N_2584,N_2530);
or U2719 (N_2719,N_2594,N_2606);
and U2720 (N_2720,N_2624,N_2497);
xor U2721 (N_2721,N_2483,N_2625);
or U2722 (N_2722,N_2419,N_2550);
or U2723 (N_2723,N_2542,N_2595);
nor U2724 (N_2724,N_2469,N_2478);
nand U2725 (N_2725,N_2678,N_2467);
and U2726 (N_2726,N_2429,N_2600);
xnor U2727 (N_2727,N_2499,N_2569);
nor U2728 (N_2728,N_2521,N_2489);
and U2729 (N_2729,N_2677,N_2466);
nand U2730 (N_2730,N_2432,N_2519);
xnor U2731 (N_2731,N_2412,N_2486);
and U2732 (N_2732,N_2635,N_2646);
nand U2733 (N_2733,N_2460,N_2563);
xor U2734 (N_2734,N_2655,N_2504);
xor U2735 (N_2735,N_2643,N_2554);
nand U2736 (N_2736,N_2472,N_2444);
xor U2737 (N_2737,N_2539,N_2512);
xor U2738 (N_2738,N_2630,N_2598);
nor U2739 (N_2739,N_2638,N_2402);
or U2740 (N_2740,N_2682,N_2587);
nor U2741 (N_2741,N_2508,N_2657);
or U2742 (N_2742,N_2431,N_2440);
nand U2743 (N_2743,N_2577,N_2560);
xnor U2744 (N_2744,N_2581,N_2498);
nor U2745 (N_2745,N_2667,N_2523);
nand U2746 (N_2746,N_2679,N_2495);
and U2747 (N_2747,N_2520,N_2656);
nor U2748 (N_2748,N_2426,N_2494);
nand U2749 (N_2749,N_2593,N_2681);
or U2750 (N_2750,N_2491,N_2511);
xnor U2751 (N_2751,N_2571,N_2518);
nand U2752 (N_2752,N_2404,N_2551);
nor U2753 (N_2753,N_2451,N_2529);
nor U2754 (N_2754,N_2588,N_2505);
and U2755 (N_2755,N_2579,N_2414);
and U2756 (N_2756,N_2528,N_2670);
xnor U2757 (N_2757,N_2596,N_2688);
and U2758 (N_2758,N_2610,N_2651);
nand U2759 (N_2759,N_2540,N_2533);
nor U2760 (N_2760,N_2666,N_2479);
xor U2761 (N_2761,N_2685,N_2436);
xor U2762 (N_2762,N_2537,N_2446);
and U2763 (N_2763,N_2644,N_2524);
and U2764 (N_2764,N_2510,N_2634);
xor U2765 (N_2765,N_2405,N_2603);
and U2766 (N_2766,N_2553,N_2632);
or U2767 (N_2767,N_2601,N_2663);
or U2768 (N_2768,N_2570,N_2475);
or U2769 (N_2769,N_2582,N_2417);
or U2770 (N_2770,N_2428,N_2462);
xnor U2771 (N_2771,N_2464,N_2418);
or U2772 (N_2772,N_2609,N_2439);
or U2773 (N_2773,N_2420,N_2619);
nand U2774 (N_2774,N_2648,N_2503);
nand U2775 (N_2775,N_2676,N_2673);
nor U2776 (N_2776,N_2641,N_2430);
nor U2777 (N_2777,N_2616,N_2629);
nand U2778 (N_2778,N_2626,N_2664);
and U2779 (N_2779,N_2456,N_2516);
and U2780 (N_2780,N_2561,N_2509);
nand U2781 (N_2781,N_2607,N_2672);
xnor U2782 (N_2782,N_2690,N_2604);
nor U2783 (N_2783,N_2662,N_2557);
and U2784 (N_2784,N_2574,N_2454);
and U2785 (N_2785,N_2500,N_2687);
xnor U2786 (N_2786,N_2416,N_2415);
or U2787 (N_2787,N_2562,N_2580);
xor U2788 (N_2788,N_2455,N_2493);
nor U2789 (N_2789,N_2633,N_2659);
nand U2790 (N_2790,N_2408,N_2443);
nand U2791 (N_2791,N_2481,N_2618);
or U2792 (N_2792,N_2527,N_2695);
xor U2793 (N_2793,N_2590,N_2548);
nor U2794 (N_2794,N_2575,N_2477);
xor U2795 (N_2795,N_2611,N_2441);
and U2796 (N_2796,N_2555,N_2547);
and U2797 (N_2797,N_2488,N_2543);
or U2798 (N_2798,N_2683,N_2566);
nand U2799 (N_2799,N_2490,N_2487);
or U2800 (N_2800,N_2526,N_2531);
nand U2801 (N_2801,N_2640,N_2433);
nand U2802 (N_2802,N_2448,N_2445);
nand U2803 (N_2803,N_2669,N_2421);
nand U2804 (N_2804,N_2502,N_2658);
xnor U2805 (N_2805,N_2654,N_2457);
nor U2806 (N_2806,N_2556,N_2565);
and U2807 (N_2807,N_2665,N_2442);
xnor U2808 (N_2808,N_2639,N_2689);
nor U2809 (N_2809,N_2620,N_2567);
xor U2810 (N_2810,N_2597,N_2501);
nor U2811 (N_2811,N_2471,N_2482);
nor U2812 (N_2812,N_2583,N_2552);
xor U2813 (N_2813,N_2564,N_2485);
or U2814 (N_2814,N_2546,N_2573);
xnor U2815 (N_2815,N_2545,N_2637);
nor U2816 (N_2816,N_2668,N_2627);
nand U2817 (N_2817,N_2463,N_2532);
or U2818 (N_2818,N_2541,N_2536);
xnor U2819 (N_2819,N_2615,N_2401);
xnor U2820 (N_2820,N_2534,N_2465);
or U2821 (N_2821,N_2559,N_2458);
nand U2822 (N_2822,N_2591,N_2413);
and U2823 (N_2823,N_2605,N_2434);
or U2824 (N_2824,N_2423,N_2453);
and U2825 (N_2825,N_2649,N_2400);
xor U2826 (N_2826,N_2525,N_2650);
nand U2827 (N_2827,N_2613,N_2409);
or U2828 (N_2828,N_2407,N_2614);
nor U2829 (N_2829,N_2450,N_2636);
xor U2830 (N_2830,N_2449,N_2480);
nor U2831 (N_2831,N_2473,N_2447);
nand U2832 (N_2832,N_2691,N_2411);
or U2833 (N_2833,N_2586,N_2578);
and U2834 (N_2834,N_2461,N_2437);
nor U2835 (N_2835,N_2694,N_2680);
and U2836 (N_2836,N_2661,N_2427);
and U2837 (N_2837,N_2424,N_2459);
nor U2838 (N_2838,N_2422,N_2506);
xnor U2839 (N_2839,N_2652,N_2410);
xor U2840 (N_2840,N_2692,N_2645);
nand U2841 (N_2841,N_2549,N_2686);
or U2842 (N_2842,N_2572,N_2699);
nor U2843 (N_2843,N_2484,N_2403);
and U2844 (N_2844,N_2476,N_2576);
nor U2845 (N_2845,N_2608,N_2653);
xnor U2846 (N_2846,N_2474,N_2674);
nand U2847 (N_2847,N_2406,N_2612);
and U2848 (N_2848,N_2589,N_2517);
xor U2849 (N_2849,N_2697,N_2496);
nand U2850 (N_2850,N_2622,N_2573);
xnor U2851 (N_2851,N_2430,N_2623);
xnor U2852 (N_2852,N_2492,N_2611);
nor U2853 (N_2853,N_2596,N_2511);
or U2854 (N_2854,N_2553,N_2459);
nor U2855 (N_2855,N_2568,N_2682);
or U2856 (N_2856,N_2630,N_2553);
and U2857 (N_2857,N_2414,N_2413);
nand U2858 (N_2858,N_2616,N_2589);
or U2859 (N_2859,N_2647,N_2603);
or U2860 (N_2860,N_2646,N_2670);
nand U2861 (N_2861,N_2682,N_2653);
nand U2862 (N_2862,N_2624,N_2678);
nand U2863 (N_2863,N_2678,N_2593);
nand U2864 (N_2864,N_2470,N_2636);
xnor U2865 (N_2865,N_2583,N_2615);
or U2866 (N_2866,N_2621,N_2531);
or U2867 (N_2867,N_2694,N_2615);
and U2868 (N_2868,N_2467,N_2403);
nor U2869 (N_2869,N_2469,N_2638);
xor U2870 (N_2870,N_2409,N_2627);
or U2871 (N_2871,N_2485,N_2569);
nand U2872 (N_2872,N_2510,N_2454);
nand U2873 (N_2873,N_2424,N_2412);
nand U2874 (N_2874,N_2436,N_2539);
and U2875 (N_2875,N_2504,N_2442);
and U2876 (N_2876,N_2485,N_2699);
xnor U2877 (N_2877,N_2438,N_2525);
xnor U2878 (N_2878,N_2568,N_2581);
and U2879 (N_2879,N_2478,N_2543);
nor U2880 (N_2880,N_2472,N_2696);
and U2881 (N_2881,N_2431,N_2551);
nand U2882 (N_2882,N_2592,N_2499);
xor U2883 (N_2883,N_2622,N_2515);
and U2884 (N_2884,N_2640,N_2484);
or U2885 (N_2885,N_2443,N_2645);
xor U2886 (N_2886,N_2460,N_2543);
nand U2887 (N_2887,N_2699,N_2570);
or U2888 (N_2888,N_2470,N_2581);
nor U2889 (N_2889,N_2558,N_2521);
nor U2890 (N_2890,N_2424,N_2675);
xor U2891 (N_2891,N_2591,N_2694);
or U2892 (N_2892,N_2415,N_2685);
or U2893 (N_2893,N_2494,N_2653);
nand U2894 (N_2894,N_2659,N_2530);
nor U2895 (N_2895,N_2677,N_2496);
and U2896 (N_2896,N_2418,N_2682);
and U2897 (N_2897,N_2527,N_2690);
or U2898 (N_2898,N_2699,N_2480);
and U2899 (N_2899,N_2511,N_2534);
nand U2900 (N_2900,N_2603,N_2506);
or U2901 (N_2901,N_2507,N_2540);
nand U2902 (N_2902,N_2679,N_2450);
and U2903 (N_2903,N_2441,N_2417);
xor U2904 (N_2904,N_2522,N_2472);
and U2905 (N_2905,N_2428,N_2692);
and U2906 (N_2906,N_2422,N_2480);
and U2907 (N_2907,N_2669,N_2510);
or U2908 (N_2908,N_2512,N_2404);
or U2909 (N_2909,N_2589,N_2667);
and U2910 (N_2910,N_2411,N_2432);
xnor U2911 (N_2911,N_2417,N_2454);
or U2912 (N_2912,N_2656,N_2487);
nor U2913 (N_2913,N_2650,N_2551);
xnor U2914 (N_2914,N_2543,N_2518);
or U2915 (N_2915,N_2634,N_2405);
or U2916 (N_2916,N_2453,N_2631);
and U2917 (N_2917,N_2645,N_2629);
nand U2918 (N_2918,N_2515,N_2656);
nor U2919 (N_2919,N_2507,N_2672);
xnor U2920 (N_2920,N_2572,N_2471);
and U2921 (N_2921,N_2504,N_2520);
or U2922 (N_2922,N_2614,N_2501);
nor U2923 (N_2923,N_2688,N_2621);
nand U2924 (N_2924,N_2614,N_2489);
xnor U2925 (N_2925,N_2537,N_2464);
or U2926 (N_2926,N_2629,N_2628);
or U2927 (N_2927,N_2541,N_2469);
xor U2928 (N_2928,N_2508,N_2622);
or U2929 (N_2929,N_2535,N_2483);
or U2930 (N_2930,N_2496,N_2572);
or U2931 (N_2931,N_2402,N_2469);
or U2932 (N_2932,N_2439,N_2518);
or U2933 (N_2933,N_2596,N_2570);
or U2934 (N_2934,N_2652,N_2496);
and U2935 (N_2935,N_2498,N_2405);
nand U2936 (N_2936,N_2432,N_2624);
nand U2937 (N_2937,N_2500,N_2502);
or U2938 (N_2938,N_2640,N_2480);
nor U2939 (N_2939,N_2504,N_2477);
or U2940 (N_2940,N_2564,N_2677);
nor U2941 (N_2941,N_2416,N_2606);
nand U2942 (N_2942,N_2513,N_2496);
and U2943 (N_2943,N_2638,N_2492);
or U2944 (N_2944,N_2405,N_2437);
or U2945 (N_2945,N_2440,N_2676);
and U2946 (N_2946,N_2650,N_2460);
or U2947 (N_2947,N_2469,N_2575);
xnor U2948 (N_2948,N_2600,N_2644);
xor U2949 (N_2949,N_2476,N_2615);
nand U2950 (N_2950,N_2604,N_2615);
nor U2951 (N_2951,N_2638,N_2649);
or U2952 (N_2952,N_2620,N_2680);
nor U2953 (N_2953,N_2612,N_2529);
or U2954 (N_2954,N_2547,N_2418);
nand U2955 (N_2955,N_2558,N_2653);
xor U2956 (N_2956,N_2442,N_2568);
or U2957 (N_2957,N_2411,N_2650);
or U2958 (N_2958,N_2654,N_2695);
nand U2959 (N_2959,N_2636,N_2549);
nand U2960 (N_2960,N_2544,N_2416);
nor U2961 (N_2961,N_2441,N_2561);
or U2962 (N_2962,N_2420,N_2500);
and U2963 (N_2963,N_2686,N_2604);
nor U2964 (N_2964,N_2612,N_2570);
nand U2965 (N_2965,N_2451,N_2431);
nor U2966 (N_2966,N_2536,N_2428);
nand U2967 (N_2967,N_2514,N_2405);
and U2968 (N_2968,N_2513,N_2568);
or U2969 (N_2969,N_2510,N_2604);
or U2970 (N_2970,N_2687,N_2631);
xor U2971 (N_2971,N_2644,N_2538);
and U2972 (N_2972,N_2539,N_2623);
or U2973 (N_2973,N_2483,N_2641);
nand U2974 (N_2974,N_2480,N_2514);
nand U2975 (N_2975,N_2577,N_2665);
or U2976 (N_2976,N_2578,N_2583);
xor U2977 (N_2977,N_2520,N_2471);
nand U2978 (N_2978,N_2603,N_2627);
xor U2979 (N_2979,N_2405,N_2689);
xnor U2980 (N_2980,N_2465,N_2491);
nor U2981 (N_2981,N_2431,N_2510);
nor U2982 (N_2982,N_2685,N_2644);
xor U2983 (N_2983,N_2545,N_2665);
xor U2984 (N_2984,N_2584,N_2528);
or U2985 (N_2985,N_2598,N_2405);
nand U2986 (N_2986,N_2598,N_2515);
nor U2987 (N_2987,N_2613,N_2616);
and U2988 (N_2988,N_2542,N_2505);
nand U2989 (N_2989,N_2464,N_2632);
nand U2990 (N_2990,N_2689,N_2511);
xor U2991 (N_2991,N_2481,N_2452);
nor U2992 (N_2992,N_2583,N_2591);
nand U2993 (N_2993,N_2460,N_2673);
and U2994 (N_2994,N_2614,N_2435);
or U2995 (N_2995,N_2575,N_2465);
nor U2996 (N_2996,N_2574,N_2466);
or U2997 (N_2997,N_2602,N_2559);
and U2998 (N_2998,N_2438,N_2643);
or U2999 (N_2999,N_2560,N_2579);
and U3000 (N_3000,N_2813,N_2851);
and U3001 (N_3001,N_2973,N_2810);
and U3002 (N_3002,N_2882,N_2902);
nor U3003 (N_3003,N_2945,N_2883);
and U3004 (N_3004,N_2730,N_2792);
or U3005 (N_3005,N_2840,N_2827);
nor U3006 (N_3006,N_2885,N_2962);
nor U3007 (N_3007,N_2826,N_2930);
and U3008 (N_3008,N_2905,N_2992);
and U3009 (N_3009,N_2816,N_2887);
nor U3010 (N_3010,N_2971,N_2859);
nand U3011 (N_3011,N_2763,N_2900);
nand U3012 (N_3012,N_2764,N_2766);
or U3013 (N_3013,N_2932,N_2839);
nor U3014 (N_3014,N_2856,N_2939);
and U3015 (N_3015,N_2830,N_2963);
and U3016 (N_3016,N_2967,N_2817);
xnor U3017 (N_3017,N_2768,N_2872);
xnor U3018 (N_3018,N_2958,N_2964);
nand U3019 (N_3019,N_2780,N_2809);
nand U3020 (N_3020,N_2742,N_2977);
and U3021 (N_3021,N_2732,N_2999);
xor U3022 (N_3022,N_2800,N_2854);
or U3023 (N_3023,N_2990,N_2740);
and U3024 (N_3024,N_2980,N_2953);
xnor U3025 (N_3025,N_2925,N_2741);
nand U3026 (N_3026,N_2794,N_2767);
nor U3027 (N_3027,N_2751,N_2702);
nand U3028 (N_3028,N_2874,N_2719);
or U3029 (N_3029,N_2968,N_2750);
or U3030 (N_3030,N_2748,N_2950);
or U3031 (N_3031,N_2713,N_2841);
xor U3032 (N_3032,N_2818,N_2749);
and U3033 (N_3033,N_2998,N_2829);
nor U3034 (N_3034,N_2825,N_2831);
nand U3035 (N_3035,N_2850,N_2888);
nor U3036 (N_3036,N_2848,N_2790);
nor U3037 (N_3037,N_2879,N_2704);
nand U3038 (N_3038,N_2847,N_2937);
xnor U3039 (N_3039,N_2868,N_2737);
and U3040 (N_3040,N_2994,N_2778);
nand U3041 (N_3041,N_2771,N_2947);
nand U3042 (N_3042,N_2983,N_2869);
and U3043 (N_3043,N_2772,N_2711);
and U3044 (N_3044,N_2891,N_2837);
nor U3045 (N_3045,N_2791,N_2821);
nand U3046 (N_3046,N_2870,N_2795);
nand U3047 (N_3047,N_2842,N_2933);
xor U3048 (N_3048,N_2708,N_2918);
and U3049 (N_3049,N_2960,N_2784);
xor U3050 (N_3050,N_2709,N_2982);
nor U3051 (N_3051,N_2736,N_2823);
nand U3052 (N_3052,N_2781,N_2735);
nand U3053 (N_3053,N_2996,N_2917);
xor U3054 (N_3054,N_2815,N_2775);
and U3055 (N_3055,N_2914,N_2836);
and U3056 (N_3056,N_2910,N_2878);
and U3057 (N_3057,N_2812,N_2701);
or U3058 (N_3058,N_2700,N_2715);
or U3059 (N_3059,N_2716,N_2832);
nand U3060 (N_3060,N_2731,N_2776);
and U3061 (N_3061,N_2822,N_2796);
nor U3062 (N_3062,N_2975,N_2838);
xnor U3063 (N_3063,N_2717,N_2940);
nor U3064 (N_3064,N_2824,N_2912);
nand U3065 (N_3065,N_2904,N_2976);
xnor U3066 (N_3066,N_2927,N_2819);
and U3067 (N_3067,N_2849,N_2961);
xnor U3068 (N_3068,N_2738,N_2804);
xnor U3069 (N_3069,N_2943,N_2745);
nor U3070 (N_3070,N_2769,N_2889);
and U3071 (N_3071,N_2928,N_2863);
and U3072 (N_3072,N_2846,N_2987);
xor U3073 (N_3073,N_2941,N_2903);
nand U3074 (N_3074,N_2858,N_2788);
or U3075 (N_3075,N_2981,N_2942);
nand U3076 (N_3076,N_2834,N_2959);
xor U3077 (N_3077,N_2753,N_2876);
nand U3078 (N_3078,N_2864,N_2844);
nor U3079 (N_3079,N_2979,N_2934);
nor U3080 (N_3080,N_2703,N_2728);
xnor U3081 (N_3081,N_2759,N_2797);
nand U3082 (N_3082,N_2965,N_2931);
nor U3083 (N_3083,N_2801,N_2919);
nor U3084 (N_3084,N_2922,N_2762);
xor U3085 (N_3085,N_2787,N_2866);
xnor U3086 (N_3086,N_2957,N_2894);
xor U3087 (N_3087,N_2721,N_2843);
or U3088 (N_3088,N_2916,N_2757);
xnor U3089 (N_3089,N_2743,N_2755);
nor U3090 (N_3090,N_2820,N_2938);
or U3091 (N_3091,N_2779,N_2993);
nor U3092 (N_3092,N_2972,N_2871);
nand U3093 (N_3093,N_2777,N_2899);
and U3094 (N_3094,N_2734,N_2714);
and U3095 (N_3095,N_2896,N_2802);
or U3096 (N_3096,N_2722,N_2718);
or U3097 (N_3097,N_2966,N_2952);
and U3098 (N_3098,N_2770,N_2760);
xnor U3099 (N_3099,N_2954,N_2956);
or U3100 (N_3100,N_2974,N_2706);
xnor U3101 (N_3101,N_2712,N_2989);
xnor U3102 (N_3102,N_2936,N_2873);
xnor U3103 (N_3103,N_2985,N_2806);
xnor U3104 (N_3104,N_2913,N_2752);
xnor U3105 (N_3105,N_2898,N_2901);
nand U3106 (N_3106,N_2988,N_2929);
or U3107 (N_3107,N_2855,N_2835);
and U3108 (N_3108,N_2948,N_2786);
or U3109 (N_3109,N_2915,N_2782);
nand U3110 (N_3110,N_2853,N_2725);
nor U3111 (N_3111,N_2978,N_2793);
or U3112 (N_3112,N_2923,N_2808);
nor U3113 (N_3113,N_2970,N_2893);
and U3114 (N_3114,N_2921,N_2811);
and U3115 (N_3115,N_2724,N_2733);
nor U3116 (N_3116,N_2860,N_2805);
nand U3117 (N_3117,N_2884,N_2908);
nand U3118 (N_3118,N_2997,N_2880);
or U3119 (N_3119,N_2785,N_2991);
nand U3120 (N_3120,N_2814,N_2906);
or U3121 (N_3121,N_2783,N_2739);
nand U3122 (N_3122,N_2944,N_2886);
or U3123 (N_3123,N_2746,N_2707);
or U3124 (N_3124,N_2949,N_2897);
nand U3125 (N_3125,N_2969,N_2833);
nor U3126 (N_3126,N_2865,N_2761);
nor U3127 (N_3127,N_2924,N_2909);
or U3128 (N_3128,N_2935,N_2828);
or U3129 (N_3129,N_2720,N_2926);
and U3130 (N_3130,N_2744,N_2798);
xnor U3131 (N_3131,N_2807,N_2726);
nor U3132 (N_3132,N_2773,N_2911);
xor U3133 (N_3133,N_2881,N_2747);
xor U3134 (N_3134,N_2986,N_2867);
nand U3135 (N_3135,N_2995,N_2765);
nand U3136 (N_3136,N_2955,N_2861);
nand U3137 (N_3137,N_2710,N_2803);
nand U3138 (N_3138,N_2756,N_2852);
nor U3139 (N_3139,N_2727,N_2729);
and U3140 (N_3140,N_2895,N_2723);
or U3141 (N_3141,N_2890,N_2789);
nand U3142 (N_3142,N_2799,N_2892);
nand U3143 (N_3143,N_2875,N_2946);
or U3144 (N_3144,N_2845,N_2705);
xnor U3145 (N_3145,N_2907,N_2951);
xnor U3146 (N_3146,N_2754,N_2984);
nor U3147 (N_3147,N_2920,N_2758);
or U3148 (N_3148,N_2877,N_2862);
nand U3149 (N_3149,N_2857,N_2774);
or U3150 (N_3150,N_2713,N_2819);
nand U3151 (N_3151,N_2768,N_2948);
and U3152 (N_3152,N_2978,N_2852);
nand U3153 (N_3153,N_2909,N_2832);
nor U3154 (N_3154,N_2715,N_2804);
nand U3155 (N_3155,N_2930,N_2859);
xnor U3156 (N_3156,N_2745,N_2711);
nor U3157 (N_3157,N_2704,N_2768);
xnor U3158 (N_3158,N_2931,N_2974);
xor U3159 (N_3159,N_2845,N_2733);
nor U3160 (N_3160,N_2751,N_2704);
or U3161 (N_3161,N_2842,N_2893);
nor U3162 (N_3162,N_2826,N_2992);
and U3163 (N_3163,N_2962,N_2749);
or U3164 (N_3164,N_2882,N_2901);
nor U3165 (N_3165,N_2862,N_2718);
nor U3166 (N_3166,N_2795,N_2958);
nor U3167 (N_3167,N_2903,N_2997);
and U3168 (N_3168,N_2912,N_2896);
nand U3169 (N_3169,N_2799,N_2789);
nand U3170 (N_3170,N_2852,N_2846);
xnor U3171 (N_3171,N_2920,N_2778);
or U3172 (N_3172,N_2966,N_2847);
nand U3173 (N_3173,N_2990,N_2779);
or U3174 (N_3174,N_2705,N_2900);
nor U3175 (N_3175,N_2844,N_2742);
nor U3176 (N_3176,N_2881,N_2949);
and U3177 (N_3177,N_2763,N_2757);
and U3178 (N_3178,N_2771,N_2797);
nor U3179 (N_3179,N_2895,N_2711);
nand U3180 (N_3180,N_2990,N_2706);
and U3181 (N_3181,N_2880,N_2916);
nand U3182 (N_3182,N_2786,N_2912);
nand U3183 (N_3183,N_2911,N_2785);
nor U3184 (N_3184,N_2894,N_2917);
or U3185 (N_3185,N_2811,N_2992);
or U3186 (N_3186,N_2920,N_2937);
nor U3187 (N_3187,N_2946,N_2884);
xor U3188 (N_3188,N_2719,N_2730);
xnor U3189 (N_3189,N_2997,N_2959);
or U3190 (N_3190,N_2731,N_2983);
nor U3191 (N_3191,N_2981,N_2990);
or U3192 (N_3192,N_2953,N_2793);
nand U3193 (N_3193,N_2705,N_2717);
xor U3194 (N_3194,N_2999,N_2789);
and U3195 (N_3195,N_2918,N_2910);
and U3196 (N_3196,N_2732,N_2779);
nor U3197 (N_3197,N_2971,N_2862);
nor U3198 (N_3198,N_2943,N_2904);
nor U3199 (N_3199,N_2749,N_2848);
nor U3200 (N_3200,N_2938,N_2804);
xor U3201 (N_3201,N_2961,N_2745);
nor U3202 (N_3202,N_2702,N_2808);
xnor U3203 (N_3203,N_2761,N_2748);
and U3204 (N_3204,N_2903,N_2822);
nand U3205 (N_3205,N_2922,N_2898);
xor U3206 (N_3206,N_2980,N_2962);
and U3207 (N_3207,N_2943,N_2934);
or U3208 (N_3208,N_2709,N_2824);
xnor U3209 (N_3209,N_2863,N_2862);
xor U3210 (N_3210,N_2855,N_2826);
or U3211 (N_3211,N_2838,N_2731);
or U3212 (N_3212,N_2923,N_2753);
xor U3213 (N_3213,N_2768,N_2840);
nor U3214 (N_3214,N_2878,N_2939);
and U3215 (N_3215,N_2705,N_2973);
xor U3216 (N_3216,N_2958,N_2797);
nand U3217 (N_3217,N_2873,N_2960);
nand U3218 (N_3218,N_2770,N_2813);
or U3219 (N_3219,N_2900,N_2751);
nand U3220 (N_3220,N_2814,N_2910);
nor U3221 (N_3221,N_2892,N_2917);
nand U3222 (N_3222,N_2992,N_2904);
nand U3223 (N_3223,N_2718,N_2956);
or U3224 (N_3224,N_2802,N_2743);
nor U3225 (N_3225,N_2803,N_2738);
nor U3226 (N_3226,N_2772,N_2976);
nand U3227 (N_3227,N_2797,N_2744);
or U3228 (N_3228,N_2727,N_2906);
nor U3229 (N_3229,N_2945,N_2747);
and U3230 (N_3230,N_2906,N_2922);
and U3231 (N_3231,N_2739,N_2723);
nor U3232 (N_3232,N_2969,N_2771);
or U3233 (N_3233,N_2877,N_2901);
xnor U3234 (N_3234,N_2979,N_2723);
and U3235 (N_3235,N_2742,N_2702);
or U3236 (N_3236,N_2904,N_2829);
and U3237 (N_3237,N_2724,N_2838);
and U3238 (N_3238,N_2887,N_2755);
xnor U3239 (N_3239,N_2861,N_2823);
nor U3240 (N_3240,N_2876,N_2864);
or U3241 (N_3241,N_2917,N_2919);
nor U3242 (N_3242,N_2948,N_2796);
and U3243 (N_3243,N_2883,N_2963);
and U3244 (N_3244,N_2959,N_2947);
xor U3245 (N_3245,N_2949,N_2858);
xnor U3246 (N_3246,N_2723,N_2933);
and U3247 (N_3247,N_2742,N_2970);
nand U3248 (N_3248,N_2849,N_2778);
and U3249 (N_3249,N_2818,N_2827);
xnor U3250 (N_3250,N_2814,N_2768);
nand U3251 (N_3251,N_2907,N_2768);
and U3252 (N_3252,N_2849,N_2851);
xnor U3253 (N_3253,N_2805,N_2717);
xor U3254 (N_3254,N_2772,N_2782);
nor U3255 (N_3255,N_2790,N_2944);
xor U3256 (N_3256,N_2814,N_2747);
xnor U3257 (N_3257,N_2864,N_2967);
nand U3258 (N_3258,N_2933,N_2977);
nand U3259 (N_3259,N_2925,N_2889);
xnor U3260 (N_3260,N_2887,N_2809);
nor U3261 (N_3261,N_2924,N_2922);
and U3262 (N_3262,N_2929,N_2958);
xor U3263 (N_3263,N_2854,N_2773);
and U3264 (N_3264,N_2736,N_2832);
or U3265 (N_3265,N_2924,N_2804);
or U3266 (N_3266,N_2861,N_2919);
xnor U3267 (N_3267,N_2798,N_2965);
or U3268 (N_3268,N_2955,N_2820);
nor U3269 (N_3269,N_2922,N_2775);
xnor U3270 (N_3270,N_2953,N_2725);
nor U3271 (N_3271,N_2984,N_2979);
nor U3272 (N_3272,N_2708,N_2898);
nor U3273 (N_3273,N_2977,N_2841);
nand U3274 (N_3274,N_2891,N_2804);
and U3275 (N_3275,N_2810,N_2955);
xnor U3276 (N_3276,N_2966,N_2744);
nor U3277 (N_3277,N_2817,N_2794);
nand U3278 (N_3278,N_2970,N_2847);
xnor U3279 (N_3279,N_2975,N_2711);
xnor U3280 (N_3280,N_2785,N_2971);
nand U3281 (N_3281,N_2780,N_2960);
xnor U3282 (N_3282,N_2972,N_2817);
xor U3283 (N_3283,N_2772,N_2978);
and U3284 (N_3284,N_2908,N_2704);
and U3285 (N_3285,N_2805,N_2986);
nand U3286 (N_3286,N_2812,N_2968);
nor U3287 (N_3287,N_2727,N_2991);
xnor U3288 (N_3288,N_2781,N_2900);
and U3289 (N_3289,N_2833,N_2935);
or U3290 (N_3290,N_2986,N_2729);
nor U3291 (N_3291,N_2723,N_2984);
nand U3292 (N_3292,N_2835,N_2708);
or U3293 (N_3293,N_2995,N_2734);
nor U3294 (N_3294,N_2993,N_2945);
and U3295 (N_3295,N_2971,N_2937);
and U3296 (N_3296,N_2907,N_2863);
and U3297 (N_3297,N_2717,N_2798);
nor U3298 (N_3298,N_2738,N_2747);
and U3299 (N_3299,N_2860,N_2704);
xor U3300 (N_3300,N_3036,N_3290);
or U3301 (N_3301,N_3081,N_3118);
and U3302 (N_3302,N_3229,N_3145);
and U3303 (N_3303,N_3245,N_3020);
and U3304 (N_3304,N_3021,N_3164);
or U3305 (N_3305,N_3051,N_3117);
xnor U3306 (N_3306,N_3057,N_3016);
nand U3307 (N_3307,N_3082,N_3131);
xor U3308 (N_3308,N_3142,N_3029);
and U3309 (N_3309,N_3122,N_3225);
xnor U3310 (N_3310,N_3003,N_3182);
xnor U3311 (N_3311,N_3188,N_3234);
or U3312 (N_3312,N_3150,N_3072);
or U3313 (N_3313,N_3185,N_3125);
xor U3314 (N_3314,N_3212,N_3048);
nand U3315 (N_3315,N_3222,N_3124);
and U3316 (N_3316,N_3062,N_3022);
nand U3317 (N_3317,N_3152,N_3272);
xnor U3318 (N_3318,N_3217,N_3066);
nor U3319 (N_3319,N_3095,N_3269);
nand U3320 (N_3320,N_3006,N_3058);
and U3321 (N_3321,N_3141,N_3154);
and U3322 (N_3322,N_3250,N_3059);
xnor U3323 (N_3323,N_3278,N_3251);
or U3324 (N_3324,N_3069,N_3293);
xor U3325 (N_3325,N_3107,N_3135);
xor U3326 (N_3326,N_3194,N_3296);
xnor U3327 (N_3327,N_3127,N_3249);
nor U3328 (N_3328,N_3071,N_3247);
or U3329 (N_3329,N_3077,N_3119);
or U3330 (N_3330,N_3094,N_3284);
nor U3331 (N_3331,N_3261,N_3139);
xor U3332 (N_3332,N_3049,N_3056);
xnor U3333 (N_3333,N_3063,N_3252);
and U3334 (N_3334,N_3240,N_3092);
nor U3335 (N_3335,N_3074,N_3209);
and U3336 (N_3336,N_3040,N_3253);
or U3337 (N_3337,N_3091,N_3153);
or U3338 (N_3338,N_3009,N_3024);
and U3339 (N_3339,N_3047,N_3170);
and U3340 (N_3340,N_3130,N_3243);
and U3341 (N_3341,N_3045,N_3149);
or U3342 (N_3342,N_3086,N_3255);
xnor U3343 (N_3343,N_3044,N_3023);
nor U3344 (N_3344,N_3041,N_3033);
nor U3345 (N_3345,N_3210,N_3053);
or U3346 (N_3346,N_3004,N_3148);
nand U3347 (N_3347,N_3208,N_3111);
xnor U3348 (N_3348,N_3183,N_3147);
nand U3349 (N_3349,N_3032,N_3256);
or U3350 (N_3350,N_3181,N_3027);
and U3351 (N_3351,N_3075,N_3060);
xnor U3352 (N_3352,N_3031,N_3159);
nor U3353 (N_3353,N_3179,N_3115);
xnor U3354 (N_3354,N_3203,N_3246);
or U3355 (N_3355,N_3175,N_3166);
nand U3356 (N_3356,N_3097,N_3035);
nor U3357 (N_3357,N_3237,N_3223);
xor U3358 (N_3358,N_3200,N_3151);
xor U3359 (N_3359,N_3242,N_3224);
and U3360 (N_3360,N_3076,N_3191);
nand U3361 (N_3361,N_3120,N_3177);
nor U3362 (N_3362,N_3167,N_3002);
nor U3363 (N_3363,N_3132,N_3068);
nand U3364 (N_3364,N_3171,N_3015);
xor U3365 (N_3365,N_3282,N_3163);
nor U3366 (N_3366,N_3158,N_3143);
nand U3367 (N_3367,N_3258,N_3079);
or U3368 (N_3368,N_3043,N_3114);
nor U3369 (N_3369,N_3219,N_3128);
xor U3370 (N_3370,N_3112,N_3244);
and U3371 (N_3371,N_3264,N_3226);
nor U3372 (N_3372,N_3106,N_3197);
nor U3373 (N_3373,N_3103,N_3270);
or U3374 (N_3374,N_3105,N_3227);
or U3375 (N_3375,N_3206,N_3100);
xnor U3376 (N_3376,N_3201,N_3214);
nor U3377 (N_3377,N_3134,N_3078);
and U3378 (N_3378,N_3241,N_3202);
nand U3379 (N_3379,N_3207,N_3133);
or U3380 (N_3380,N_3236,N_3018);
nor U3381 (N_3381,N_3285,N_3013);
nand U3382 (N_3382,N_3146,N_3101);
or U3383 (N_3383,N_3129,N_3279);
xnor U3384 (N_3384,N_3001,N_3187);
and U3385 (N_3385,N_3108,N_3287);
and U3386 (N_3386,N_3291,N_3157);
and U3387 (N_3387,N_3088,N_3289);
nand U3388 (N_3388,N_3233,N_3087);
nand U3389 (N_3389,N_3011,N_3030);
nand U3390 (N_3390,N_3230,N_3294);
nor U3391 (N_3391,N_3160,N_3039);
or U3392 (N_3392,N_3121,N_3268);
and U3393 (N_3393,N_3262,N_3277);
xnor U3394 (N_3394,N_3073,N_3138);
nand U3395 (N_3395,N_3162,N_3000);
or U3396 (N_3396,N_3025,N_3235);
nor U3397 (N_3397,N_3070,N_3050);
nand U3398 (N_3398,N_3273,N_3193);
or U3399 (N_3399,N_3099,N_3257);
nor U3400 (N_3400,N_3144,N_3172);
and U3401 (N_3401,N_3218,N_3288);
and U3402 (N_3402,N_3017,N_3228);
or U3403 (N_3403,N_3123,N_3054);
nor U3404 (N_3404,N_3104,N_3010);
and U3405 (N_3405,N_3026,N_3007);
xnor U3406 (N_3406,N_3174,N_3110);
nor U3407 (N_3407,N_3263,N_3028);
nor U3408 (N_3408,N_3037,N_3140);
or U3409 (N_3409,N_3090,N_3038);
xnor U3410 (N_3410,N_3176,N_3042);
xor U3411 (N_3411,N_3286,N_3168);
nand U3412 (N_3412,N_3136,N_3098);
xnor U3413 (N_3413,N_3267,N_3216);
or U3414 (N_3414,N_3085,N_3213);
nand U3415 (N_3415,N_3067,N_3126);
xor U3416 (N_3416,N_3232,N_3276);
xor U3417 (N_3417,N_3292,N_3199);
nor U3418 (N_3418,N_3005,N_3109);
nor U3419 (N_3419,N_3283,N_3161);
xnor U3420 (N_3420,N_3297,N_3196);
nand U3421 (N_3421,N_3178,N_3184);
nand U3422 (N_3422,N_3084,N_3019);
and U3423 (N_3423,N_3231,N_3254);
nand U3424 (N_3424,N_3198,N_3204);
and U3425 (N_3425,N_3211,N_3266);
and U3426 (N_3426,N_3064,N_3093);
or U3427 (N_3427,N_3173,N_3281);
nor U3428 (N_3428,N_3186,N_3052);
nand U3429 (N_3429,N_3155,N_3295);
or U3430 (N_3430,N_3061,N_3260);
or U3431 (N_3431,N_3205,N_3298);
or U3432 (N_3432,N_3280,N_3034);
nand U3433 (N_3433,N_3089,N_3113);
nand U3434 (N_3434,N_3248,N_3169);
nor U3435 (N_3435,N_3220,N_3065);
xnor U3436 (N_3436,N_3215,N_3299);
nor U3437 (N_3437,N_3238,N_3180);
nor U3438 (N_3438,N_3055,N_3271);
xor U3439 (N_3439,N_3190,N_3274);
xnor U3440 (N_3440,N_3265,N_3008);
nor U3441 (N_3441,N_3102,N_3275);
nor U3442 (N_3442,N_3137,N_3156);
and U3443 (N_3443,N_3080,N_3195);
nand U3444 (N_3444,N_3012,N_3192);
and U3445 (N_3445,N_3189,N_3083);
nor U3446 (N_3446,N_3096,N_3239);
nand U3447 (N_3447,N_3259,N_3165);
nor U3448 (N_3448,N_3116,N_3014);
nor U3449 (N_3449,N_3046,N_3221);
or U3450 (N_3450,N_3073,N_3103);
nor U3451 (N_3451,N_3197,N_3245);
xor U3452 (N_3452,N_3071,N_3223);
nand U3453 (N_3453,N_3293,N_3025);
nand U3454 (N_3454,N_3250,N_3224);
nand U3455 (N_3455,N_3042,N_3294);
nand U3456 (N_3456,N_3215,N_3001);
and U3457 (N_3457,N_3119,N_3260);
and U3458 (N_3458,N_3157,N_3034);
and U3459 (N_3459,N_3076,N_3146);
or U3460 (N_3460,N_3282,N_3125);
nor U3461 (N_3461,N_3001,N_3188);
nor U3462 (N_3462,N_3298,N_3037);
or U3463 (N_3463,N_3299,N_3221);
nand U3464 (N_3464,N_3045,N_3239);
nand U3465 (N_3465,N_3287,N_3052);
nor U3466 (N_3466,N_3217,N_3044);
or U3467 (N_3467,N_3264,N_3119);
xnor U3468 (N_3468,N_3128,N_3163);
nor U3469 (N_3469,N_3003,N_3289);
or U3470 (N_3470,N_3047,N_3034);
or U3471 (N_3471,N_3043,N_3138);
nand U3472 (N_3472,N_3023,N_3031);
xnor U3473 (N_3473,N_3058,N_3020);
and U3474 (N_3474,N_3070,N_3221);
and U3475 (N_3475,N_3008,N_3188);
nor U3476 (N_3476,N_3117,N_3238);
xor U3477 (N_3477,N_3170,N_3036);
nor U3478 (N_3478,N_3157,N_3045);
nor U3479 (N_3479,N_3241,N_3189);
xnor U3480 (N_3480,N_3206,N_3233);
and U3481 (N_3481,N_3175,N_3034);
nand U3482 (N_3482,N_3041,N_3014);
nand U3483 (N_3483,N_3161,N_3235);
and U3484 (N_3484,N_3183,N_3136);
nor U3485 (N_3485,N_3229,N_3191);
nand U3486 (N_3486,N_3172,N_3127);
and U3487 (N_3487,N_3246,N_3292);
and U3488 (N_3488,N_3259,N_3227);
or U3489 (N_3489,N_3181,N_3246);
nand U3490 (N_3490,N_3042,N_3257);
xnor U3491 (N_3491,N_3114,N_3160);
nor U3492 (N_3492,N_3191,N_3023);
nand U3493 (N_3493,N_3051,N_3080);
and U3494 (N_3494,N_3007,N_3027);
or U3495 (N_3495,N_3109,N_3192);
and U3496 (N_3496,N_3210,N_3273);
or U3497 (N_3497,N_3068,N_3176);
and U3498 (N_3498,N_3093,N_3218);
nand U3499 (N_3499,N_3193,N_3205);
xnor U3500 (N_3500,N_3190,N_3203);
or U3501 (N_3501,N_3211,N_3018);
and U3502 (N_3502,N_3144,N_3150);
nand U3503 (N_3503,N_3161,N_3020);
xor U3504 (N_3504,N_3252,N_3077);
or U3505 (N_3505,N_3163,N_3219);
and U3506 (N_3506,N_3240,N_3161);
xnor U3507 (N_3507,N_3287,N_3050);
nor U3508 (N_3508,N_3241,N_3262);
or U3509 (N_3509,N_3279,N_3169);
and U3510 (N_3510,N_3269,N_3215);
xnor U3511 (N_3511,N_3089,N_3151);
xor U3512 (N_3512,N_3127,N_3219);
nor U3513 (N_3513,N_3101,N_3100);
nand U3514 (N_3514,N_3025,N_3282);
nor U3515 (N_3515,N_3074,N_3176);
xor U3516 (N_3516,N_3287,N_3163);
xor U3517 (N_3517,N_3090,N_3203);
and U3518 (N_3518,N_3189,N_3138);
and U3519 (N_3519,N_3112,N_3137);
xor U3520 (N_3520,N_3207,N_3153);
and U3521 (N_3521,N_3233,N_3194);
or U3522 (N_3522,N_3236,N_3243);
and U3523 (N_3523,N_3288,N_3252);
or U3524 (N_3524,N_3136,N_3051);
nor U3525 (N_3525,N_3001,N_3212);
xor U3526 (N_3526,N_3197,N_3297);
nor U3527 (N_3527,N_3285,N_3052);
nor U3528 (N_3528,N_3218,N_3000);
xnor U3529 (N_3529,N_3034,N_3087);
nor U3530 (N_3530,N_3046,N_3200);
xnor U3531 (N_3531,N_3180,N_3155);
xor U3532 (N_3532,N_3085,N_3273);
xnor U3533 (N_3533,N_3052,N_3235);
xnor U3534 (N_3534,N_3060,N_3299);
nand U3535 (N_3535,N_3196,N_3010);
and U3536 (N_3536,N_3064,N_3204);
nand U3537 (N_3537,N_3085,N_3183);
nor U3538 (N_3538,N_3151,N_3096);
nand U3539 (N_3539,N_3110,N_3089);
nand U3540 (N_3540,N_3029,N_3038);
or U3541 (N_3541,N_3176,N_3284);
and U3542 (N_3542,N_3025,N_3097);
nand U3543 (N_3543,N_3039,N_3007);
or U3544 (N_3544,N_3118,N_3255);
and U3545 (N_3545,N_3239,N_3137);
nand U3546 (N_3546,N_3232,N_3164);
and U3547 (N_3547,N_3169,N_3185);
nand U3548 (N_3548,N_3091,N_3211);
nand U3549 (N_3549,N_3160,N_3075);
xnor U3550 (N_3550,N_3131,N_3243);
and U3551 (N_3551,N_3094,N_3040);
nor U3552 (N_3552,N_3128,N_3236);
or U3553 (N_3553,N_3267,N_3016);
nor U3554 (N_3554,N_3196,N_3210);
and U3555 (N_3555,N_3295,N_3148);
nand U3556 (N_3556,N_3120,N_3124);
nand U3557 (N_3557,N_3290,N_3171);
or U3558 (N_3558,N_3092,N_3294);
nand U3559 (N_3559,N_3177,N_3030);
nand U3560 (N_3560,N_3143,N_3025);
xnor U3561 (N_3561,N_3076,N_3288);
and U3562 (N_3562,N_3239,N_3017);
xor U3563 (N_3563,N_3011,N_3071);
and U3564 (N_3564,N_3064,N_3168);
nor U3565 (N_3565,N_3256,N_3207);
xnor U3566 (N_3566,N_3126,N_3223);
nor U3567 (N_3567,N_3291,N_3092);
xnor U3568 (N_3568,N_3134,N_3107);
xnor U3569 (N_3569,N_3291,N_3059);
xnor U3570 (N_3570,N_3294,N_3244);
xnor U3571 (N_3571,N_3016,N_3167);
nor U3572 (N_3572,N_3035,N_3258);
nand U3573 (N_3573,N_3093,N_3026);
nor U3574 (N_3574,N_3218,N_3256);
nor U3575 (N_3575,N_3284,N_3133);
nor U3576 (N_3576,N_3256,N_3288);
nand U3577 (N_3577,N_3220,N_3010);
nor U3578 (N_3578,N_3111,N_3166);
nor U3579 (N_3579,N_3016,N_3269);
nor U3580 (N_3580,N_3159,N_3161);
or U3581 (N_3581,N_3173,N_3205);
xor U3582 (N_3582,N_3178,N_3007);
and U3583 (N_3583,N_3056,N_3244);
xor U3584 (N_3584,N_3220,N_3287);
xor U3585 (N_3585,N_3046,N_3192);
nand U3586 (N_3586,N_3167,N_3125);
nand U3587 (N_3587,N_3263,N_3072);
or U3588 (N_3588,N_3004,N_3218);
and U3589 (N_3589,N_3279,N_3240);
nand U3590 (N_3590,N_3100,N_3014);
and U3591 (N_3591,N_3121,N_3132);
nor U3592 (N_3592,N_3148,N_3040);
nand U3593 (N_3593,N_3235,N_3122);
nand U3594 (N_3594,N_3004,N_3253);
nor U3595 (N_3595,N_3167,N_3213);
nand U3596 (N_3596,N_3157,N_3160);
or U3597 (N_3597,N_3243,N_3009);
and U3598 (N_3598,N_3020,N_3033);
nor U3599 (N_3599,N_3272,N_3004);
or U3600 (N_3600,N_3468,N_3374);
or U3601 (N_3601,N_3422,N_3312);
nor U3602 (N_3602,N_3471,N_3524);
or U3603 (N_3603,N_3516,N_3318);
nand U3604 (N_3604,N_3529,N_3511);
and U3605 (N_3605,N_3456,N_3587);
or U3606 (N_3606,N_3444,N_3419);
xnor U3607 (N_3607,N_3326,N_3405);
or U3608 (N_3608,N_3310,N_3591);
nor U3609 (N_3609,N_3599,N_3499);
or U3610 (N_3610,N_3396,N_3391);
or U3611 (N_3611,N_3433,N_3497);
nand U3612 (N_3612,N_3306,N_3596);
and U3613 (N_3613,N_3439,N_3340);
and U3614 (N_3614,N_3465,N_3362);
and U3615 (N_3615,N_3530,N_3515);
or U3616 (N_3616,N_3555,N_3570);
xor U3617 (N_3617,N_3552,N_3531);
and U3618 (N_3618,N_3490,N_3407);
nand U3619 (N_3619,N_3474,N_3546);
or U3620 (N_3620,N_3417,N_3428);
nand U3621 (N_3621,N_3375,N_3452);
nor U3622 (N_3622,N_3356,N_3408);
nor U3623 (N_3623,N_3455,N_3593);
nor U3624 (N_3624,N_3431,N_3486);
nor U3625 (N_3625,N_3594,N_3496);
xnor U3626 (N_3626,N_3342,N_3321);
or U3627 (N_3627,N_3527,N_3475);
or U3628 (N_3628,N_3350,N_3392);
xor U3629 (N_3629,N_3488,N_3506);
nand U3630 (N_3630,N_3373,N_3371);
nor U3631 (N_3631,N_3369,N_3335);
and U3632 (N_3632,N_3443,N_3410);
nand U3633 (N_3633,N_3359,N_3545);
or U3634 (N_3634,N_3432,N_3418);
xnor U3635 (N_3635,N_3595,N_3523);
nand U3636 (N_3636,N_3331,N_3532);
or U3637 (N_3637,N_3420,N_3353);
xnor U3638 (N_3638,N_3470,N_3401);
and U3639 (N_3639,N_3507,N_3569);
or U3640 (N_3640,N_3317,N_3493);
and U3641 (N_3641,N_3332,N_3548);
xor U3642 (N_3642,N_3320,N_3505);
nand U3643 (N_3643,N_3333,N_3438);
xnor U3644 (N_3644,N_3361,N_3365);
nor U3645 (N_3645,N_3514,N_3416);
nand U3646 (N_3646,N_3400,N_3517);
and U3647 (N_3647,N_3550,N_3462);
or U3648 (N_3648,N_3313,N_3352);
nand U3649 (N_3649,N_3349,N_3502);
nand U3650 (N_3650,N_3351,N_3492);
or U3651 (N_3651,N_3344,N_3554);
nand U3652 (N_3652,N_3380,N_3571);
nor U3653 (N_3653,N_3576,N_3328);
and U3654 (N_3654,N_3458,N_3397);
nand U3655 (N_3655,N_3539,N_3543);
nand U3656 (N_3656,N_3437,N_3453);
xnor U3657 (N_3657,N_3466,N_3575);
nor U3658 (N_3658,N_3395,N_3322);
and U3659 (N_3659,N_3533,N_3343);
or U3660 (N_3660,N_3482,N_3304);
and U3661 (N_3661,N_3513,N_3363);
xor U3662 (N_3662,N_3557,N_3327);
xnor U3663 (N_3663,N_3491,N_3519);
or U3664 (N_3664,N_3580,N_3319);
nand U3665 (N_3665,N_3556,N_3479);
xnor U3666 (N_3666,N_3553,N_3518);
nand U3667 (N_3667,N_3354,N_3338);
xnor U3668 (N_3668,N_3325,N_3414);
xnor U3669 (N_3669,N_3478,N_3525);
or U3670 (N_3670,N_3307,N_3551);
or U3671 (N_3671,N_3430,N_3508);
nand U3672 (N_3672,N_3538,N_3549);
and U3673 (N_3673,N_3314,N_3563);
nor U3674 (N_3674,N_3454,N_3447);
xnor U3675 (N_3675,N_3572,N_3330);
nor U3676 (N_3676,N_3542,N_3535);
or U3677 (N_3677,N_3584,N_3489);
xnor U3678 (N_3678,N_3472,N_3436);
nor U3679 (N_3679,N_3526,N_3510);
and U3680 (N_3680,N_3381,N_3337);
or U3681 (N_3681,N_3302,N_3567);
nand U3682 (N_3682,N_3540,N_3463);
nor U3683 (N_3683,N_3329,N_3424);
nand U3684 (N_3684,N_3429,N_3503);
nor U3685 (N_3685,N_3303,N_3480);
nor U3686 (N_3686,N_3585,N_3435);
or U3687 (N_3687,N_3394,N_3485);
xor U3688 (N_3688,N_3562,N_3347);
and U3689 (N_3689,N_3323,N_3382);
nor U3690 (N_3690,N_3426,N_3387);
nand U3691 (N_3691,N_3441,N_3481);
or U3692 (N_3692,N_3520,N_3425);
or U3693 (N_3693,N_3390,N_3592);
and U3694 (N_3694,N_3528,N_3364);
or U3695 (N_3695,N_3477,N_3577);
nand U3696 (N_3696,N_3336,N_3589);
nand U3697 (N_3697,N_3367,N_3504);
or U3698 (N_3698,N_3383,N_3560);
and U3699 (N_3699,N_3366,N_3574);
or U3700 (N_3700,N_3389,N_3355);
xor U3701 (N_3701,N_3579,N_3469);
nand U3702 (N_3702,N_3464,N_3566);
and U3703 (N_3703,N_3451,N_3348);
or U3704 (N_3704,N_3427,N_3370);
or U3705 (N_3705,N_3568,N_3402);
nor U3706 (N_3706,N_3590,N_3301);
nand U3707 (N_3707,N_3399,N_3376);
nand U3708 (N_3708,N_3403,N_3345);
and U3709 (N_3709,N_3309,N_3598);
nand U3710 (N_3710,N_3597,N_3457);
xnor U3711 (N_3711,N_3440,N_3421);
and U3712 (N_3712,N_3448,N_3386);
nor U3713 (N_3713,N_3565,N_3413);
nor U3714 (N_3714,N_3522,N_3467);
and U3715 (N_3715,N_3368,N_3498);
or U3716 (N_3716,N_3442,N_3379);
and U3717 (N_3717,N_3377,N_3358);
nand U3718 (N_3718,N_3446,N_3583);
or U3719 (N_3719,N_3393,N_3547);
xnor U3720 (N_3720,N_3459,N_3536);
and U3721 (N_3721,N_3558,N_3385);
xnor U3722 (N_3722,N_3494,N_3315);
nor U3723 (N_3723,N_3450,N_3384);
nand U3724 (N_3724,N_3308,N_3341);
xor U3725 (N_3725,N_3483,N_3564);
or U3726 (N_3726,N_3324,N_3509);
and U3727 (N_3727,N_3588,N_3300);
and U3728 (N_3728,N_3512,N_3473);
nand U3729 (N_3729,N_3521,N_3360);
and U3730 (N_3730,N_3409,N_3541);
nor U3731 (N_3731,N_3500,N_3411);
and U3732 (N_3732,N_3460,N_3561);
and U3733 (N_3733,N_3484,N_3388);
nor U3734 (N_3734,N_3487,N_3501);
nand U3735 (N_3735,N_3559,N_3461);
and U3736 (N_3736,N_3412,N_3404);
and U3737 (N_3737,N_3581,N_3406);
nor U3738 (N_3738,N_3573,N_3316);
nor U3739 (N_3739,N_3346,N_3305);
nand U3740 (N_3740,N_3544,N_3378);
and U3741 (N_3741,N_3398,N_3445);
xnor U3742 (N_3742,N_3586,N_3339);
xor U3743 (N_3743,N_3415,N_3495);
nor U3744 (N_3744,N_3582,N_3476);
nor U3745 (N_3745,N_3311,N_3537);
and U3746 (N_3746,N_3423,N_3372);
and U3747 (N_3747,N_3434,N_3534);
nand U3748 (N_3748,N_3357,N_3449);
or U3749 (N_3749,N_3578,N_3334);
nor U3750 (N_3750,N_3355,N_3365);
nor U3751 (N_3751,N_3448,N_3377);
nor U3752 (N_3752,N_3445,N_3493);
nand U3753 (N_3753,N_3596,N_3349);
nand U3754 (N_3754,N_3466,N_3411);
or U3755 (N_3755,N_3463,N_3495);
and U3756 (N_3756,N_3496,N_3335);
nand U3757 (N_3757,N_3348,N_3394);
xnor U3758 (N_3758,N_3370,N_3411);
and U3759 (N_3759,N_3543,N_3540);
or U3760 (N_3760,N_3383,N_3324);
nor U3761 (N_3761,N_3390,N_3376);
xnor U3762 (N_3762,N_3337,N_3329);
and U3763 (N_3763,N_3462,N_3388);
nor U3764 (N_3764,N_3411,N_3328);
xnor U3765 (N_3765,N_3539,N_3328);
nand U3766 (N_3766,N_3390,N_3324);
xnor U3767 (N_3767,N_3562,N_3566);
or U3768 (N_3768,N_3525,N_3357);
or U3769 (N_3769,N_3432,N_3406);
and U3770 (N_3770,N_3586,N_3450);
nand U3771 (N_3771,N_3450,N_3403);
nand U3772 (N_3772,N_3490,N_3592);
nor U3773 (N_3773,N_3329,N_3472);
xor U3774 (N_3774,N_3479,N_3551);
or U3775 (N_3775,N_3546,N_3395);
nor U3776 (N_3776,N_3545,N_3426);
and U3777 (N_3777,N_3534,N_3467);
nor U3778 (N_3778,N_3513,N_3472);
or U3779 (N_3779,N_3472,N_3509);
nand U3780 (N_3780,N_3529,N_3415);
nor U3781 (N_3781,N_3357,N_3345);
and U3782 (N_3782,N_3414,N_3436);
or U3783 (N_3783,N_3384,N_3523);
or U3784 (N_3784,N_3362,N_3459);
nor U3785 (N_3785,N_3350,N_3356);
and U3786 (N_3786,N_3355,N_3516);
nor U3787 (N_3787,N_3539,N_3385);
or U3788 (N_3788,N_3533,N_3490);
nand U3789 (N_3789,N_3526,N_3373);
or U3790 (N_3790,N_3500,N_3418);
nor U3791 (N_3791,N_3335,N_3483);
nand U3792 (N_3792,N_3306,N_3463);
nand U3793 (N_3793,N_3413,N_3570);
and U3794 (N_3794,N_3404,N_3564);
nand U3795 (N_3795,N_3386,N_3430);
nor U3796 (N_3796,N_3551,N_3382);
nor U3797 (N_3797,N_3446,N_3562);
and U3798 (N_3798,N_3437,N_3573);
xor U3799 (N_3799,N_3456,N_3411);
nand U3800 (N_3800,N_3347,N_3510);
and U3801 (N_3801,N_3429,N_3489);
xor U3802 (N_3802,N_3422,N_3350);
nand U3803 (N_3803,N_3545,N_3365);
xnor U3804 (N_3804,N_3302,N_3576);
and U3805 (N_3805,N_3531,N_3328);
nand U3806 (N_3806,N_3387,N_3459);
xor U3807 (N_3807,N_3414,N_3499);
xnor U3808 (N_3808,N_3343,N_3404);
or U3809 (N_3809,N_3428,N_3492);
and U3810 (N_3810,N_3339,N_3454);
nand U3811 (N_3811,N_3430,N_3573);
or U3812 (N_3812,N_3448,N_3432);
and U3813 (N_3813,N_3443,N_3380);
nor U3814 (N_3814,N_3444,N_3425);
nand U3815 (N_3815,N_3415,N_3534);
or U3816 (N_3816,N_3477,N_3358);
or U3817 (N_3817,N_3332,N_3514);
and U3818 (N_3818,N_3591,N_3319);
xnor U3819 (N_3819,N_3484,N_3409);
or U3820 (N_3820,N_3360,N_3377);
and U3821 (N_3821,N_3305,N_3425);
xor U3822 (N_3822,N_3336,N_3382);
nor U3823 (N_3823,N_3469,N_3382);
xnor U3824 (N_3824,N_3454,N_3338);
and U3825 (N_3825,N_3361,N_3359);
or U3826 (N_3826,N_3587,N_3489);
and U3827 (N_3827,N_3470,N_3321);
nor U3828 (N_3828,N_3438,N_3595);
nand U3829 (N_3829,N_3477,N_3351);
and U3830 (N_3830,N_3566,N_3574);
and U3831 (N_3831,N_3514,N_3476);
nor U3832 (N_3832,N_3405,N_3589);
nand U3833 (N_3833,N_3341,N_3548);
nand U3834 (N_3834,N_3548,N_3599);
xor U3835 (N_3835,N_3397,N_3596);
nor U3836 (N_3836,N_3414,N_3353);
nor U3837 (N_3837,N_3424,N_3480);
xor U3838 (N_3838,N_3461,N_3394);
nand U3839 (N_3839,N_3598,N_3384);
nand U3840 (N_3840,N_3443,N_3581);
nand U3841 (N_3841,N_3427,N_3564);
nand U3842 (N_3842,N_3487,N_3345);
nor U3843 (N_3843,N_3568,N_3476);
or U3844 (N_3844,N_3389,N_3415);
nor U3845 (N_3845,N_3569,N_3598);
and U3846 (N_3846,N_3388,N_3510);
nand U3847 (N_3847,N_3414,N_3530);
nand U3848 (N_3848,N_3504,N_3579);
nor U3849 (N_3849,N_3463,N_3494);
or U3850 (N_3850,N_3581,N_3419);
or U3851 (N_3851,N_3513,N_3522);
xnor U3852 (N_3852,N_3443,N_3574);
and U3853 (N_3853,N_3432,N_3551);
or U3854 (N_3854,N_3321,N_3411);
nand U3855 (N_3855,N_3377,N_3510);
or U3856 (N_3856,N_3403,N_3400);
or U3857 (N_3857,N_3595,N_3594);
nor U3858 (N_3858,N_3509,N_3519);
xnor U3859 (N_3859,N_3518,N_3337);
and U3860 (N_3860,N_3408,N_3313);
nand U3861 (N_3861,N_3439,N_3455);
and U3862 (N_3862,N_3453,N_3485);
xor U3863 (N_3863,N_3316,N_3371);
or U3864 (N_3864,N_3405,N_3544);
or U3865 (N_3865,N_3548,N_3580);
nor U3866 (N_3866,N_3515,N_3510);
nand U3867 (N_3867,N_3310,N_3476);
xor U3868 (N_3868,N_3306,N_3377);
xnor U3869 (N_3869,N_3402,N_3405);
or U3870 (N_3870,N_3347,N_3305);
xnor U3871 (N_3871,N_3491,N_3486);
or U3872 (N_3872,N_3586,N_3476);
or U3873 (N_3873,N_3519,N_3365);
and U3874 (N_3874,N_3442,N_3374);
or U3875 (N_3875,N_3522,N_3561);
and U3876 (N_3876,N_3532,N_3311);
nand U3877 (N_3877,N_3322,N_3388);
xor U3878 (N_3878,N_3335,N_3503);
xor U3879 (N_3879,N_3521,N_3435);
nand U3880 (N_3880,N_3542,N_3544);
xor U3881 (N_3881,N_3578,N_3474);
and U3882 (N_3882,N_3382,N_3535);
nand U3883 (N_3883,N_3488,N_3525);
nor U3884 (N_3884,N_3450,N_3368);
nand U3885 (N_3885,N_3355,N_3480);
and U3886 (N_3886,N_3388,N_3381);
nand U3887 (N_3887,N_3332,N_3418);
nor U3888 (N_3888,N_3429,N_3389);
or U3889 (N_3889,N_3513,N_3329);
or U3890 (N_3890,N_3484,N_3458);
xnor U3891 (N_3891,N_3332,N_3559);
or U3892 (N_3892,N_3484,N_3583);
and U3893 (N_3893,N_3489,N_3469);
nor U3894 (N_3894,N_3368,N_3438);
and U3895 (N_3895,N_3522,N_3360);
nand U3896 (N_3896,N_3400,N_3585);
or U3897 (N_3897,N_3399,N_3559);
xnor U3898 (N_3898,N_3429,N_3588);
or U3899 (N_3899,N_3490,N_3316);
or U3900 (N_3900,N_3774,N_3790);
nand U3901 (N_3901,N_3702,N_3777);
xor U3902 (N_3902,N_3886,N_3826);
nor U3903 (N_3903,N_3779,N_3854);
nor U3904 (N_3904,N_3791,N_3718);
nand U3905 (N_3905,N_3861,N_3683);
nor U3906 (N_3906,N_3698,N_3661);
xnor U3907 (N_3907,N_3612,N_3682);
nand U3908 (N_3908,N_3807,N_3782);
nor U3909 (N_3909,N_3789,N_3755);
or U3910 (N_3910,N_3655,N_3831);
xnor U3911 (N_3911,N_3768,N_3868);
and U3912 (N_3912,N_3762,N_3756);
nor U3913 (N_3913,N_3644,N_3838);
nand U3914 (N_3914,N_3764,N_3712);
or U3915 (N_3915,N_3647,N_3643);
or U3916 (N_3916,N_3851,N_3641);
or U3917 (N_3917,N_3651,N_3728);
and U3918 (N_3918,N_3634,N_3800);
xnor U3919 (N_3919,N_3658,N_3897);
or U3920 (N_3920,N_3846,N_3862);
nor U3921 (N_3921,N_3687,N_3827);
or U3922 (N_3922,N_3686,N_3860);
nor U3923 (N_3923,N_3738,N_3781);
and U3924 (N_3924,N_3714,N_3732);
nand U3925 (N_3925,N_3867,N_3637);
or U3926 (N_3926,N_3803,N_3614);
xor U3927 (N_3927,N_3872,N_3741);
and U3928 (N_3928,N_3815,N_3623);
nand U3929 (N_3929,N_3674,N_3848);
and U3930 (N_3930,N_3734,N_3694);
xor U3931 (N_3931,N_3716,N_3692);
nand U3932 (N_3932,N_3783,N_3684);
and U3933 (N_3933,N_3725,N_3744);
xor U3934 (N_3934,N_3875,N_3631);
and U3935 (N_3935,N_3776,N_3746);
and U3936 (N_3936,N_3881,N_3856);
nand U3937 (N_3937,N_3677,N_3652);
nor U3938 (N_3938,N_3710,N_3666);
nand U3939 (N_3939,N_3703,N_3757);
nand U3940 (N_3940,N_3742,N_3608);
or U3941 (N_3941,N_3770,N_3660);
nor U3942 (N_3942,N_3720,N_3681);
xor U3943 (N_3943,N_3855,N_3813);
or U3944 (N_3944,N_3695,N_3898);
or U3945 (N_3945,N_3794,N_3676);
nor U3946 (N_3946,N_3765,N_3858);
xnor U3947 (N_3947,N_3622,N_3606);
xnor U3948 (N_3948,N_3893,N_3834);
nor U3949 (N_3949,N_3825,N_3638);
nor U3950 (N_3950,N_3602,N_3615);
nor U3951 (N_3951,N_3653,N_3849);
or U3952 (N_3952,N_3625,N_3662);
nand U3953 (N_3953,N_3894,N_3880);
nor U3954 (N_3954,N_3735,N_3889);
and U3955 (N_3955,N_3633,N_3717);
xor U3956 (N_3956,N_3648,N_3727);
and U3957 (N_3957,N_3721,N_3624);
xnor U3958 (N_3958,N_3729,N_3773);
or U3959 (N_3959,N_3796,N_3837);
and U3960 (N_3960,N_3621,N_3816);
or U3961 (N_3961,N_3784,N_3785);
or U3962 (N_3962,N_3767,N_3832);
and U3963 (N_3963,N_3751,N_3795);
nand U3964 (N_3964,N_3759,N_3891);
nor U3965 (N_3965,N_3670,N_3866);
xor U3966 (N_3966,N_3873,N_3845);
nand U3967 (N_3967,N_3739,N_3769);
nand U3968 (N_3968,N_3899,N_3678);
nor U3969 (N_3969,N_3863,N_3693);
xor U3970 (N_3970,N_3616,N_3724);
xor U3971 (N_3971,N_3731,N_3814);
xor U3972 (N_3972,N_3664,N_3707);
nor U3973 (N_3973,N_3610,N_3749);
or U3974 (N_3974,N_3824,N_3645);
and U3975 (N_3975,N_3799,N_3806);
nor U3976 (N_3976,N_3745,N_3890);
nand U3977 (N_3977,N_3792,N_3805);
and U3978 (N_3978,N_3819,N_3705);
nor U3979 (N_3979,N_3828,N_3619);
nand U3980 (N_3980,N_3667,N_3704);
nor U3981 (N_3981,N_3669,N_3723);
or U3982 (N_3982,N_3696,N_3766);
nand U3983 (N_3983,N_3620,N_3627);
and U3984 (N_3984,N_3771,N_3689);
and U3985 (N_3985,N_3715,N_3758);
nand U3986 (N_3986,N_3857,N_3787);
nand U3987 (N_3987,N_3752,N_3663);
and U3988 (N_3988,N_3874,N_3690);
or U3989 (N_3989,N_3844,N_3812);
nand U3990 (N_3990,N_3871,N_3895);
nand U3991 (N_3991,N_3668,N_3835);
xor U3992 (N_3992,N_3811,N_3671);
or U3993 (N_3993,N_3869,N_3865);
and U3994 (N_3994,N_3630,N_3659);
nand U3995 (N_3995,N_3760,N_3743);
and U3996 (N_3996,N_3642,N_3804);
and U3997 (N_3997,N_3892,N_3818);
or U3998 (N_3998,N_3636,N_3798);
nand U3999 (N_3999,N_3793,N_3836);
nor U4000 (N_4000,N_3635,N_3822);
xor U4001 (N_4001,N_3656,N_3737);
and U4002 (N_4002,N_3650,N_3801);
or U4003 (N_4003,N_3639,N_3699);
xnor U4004 (N_4004,N_3605,N_3809);
nand U4005 (N_4005,N_3680,N_3879);
nor U4006 (N_4006,N_3778,N_3883);
nor U4007 (N_4007,N_3709,N_3888);
nor U4008 (N_4008,N_3697,N_3685);
xnor U4009 (N_4009,N_3706,N_3673);
xnor U4010 (N_4010,N_3618,N_3607);
xor U4011 (N_4011,N_3646,N_3839);
or U4012 (N_4012,N_3701,N_3802);
and U4013 (N_4013,N_3842,N_3754);
nand U4014 (N_4014,N_3859,N_3613);
xor U4015 (N_4015,N_3821,N_3654);
or U4016 (N_4016,N_3877,N_3786);
xor U4017 (N_4017,N_3665,N_3626);
or U4018 (N_4018,N_3876,N_3688);
xnor U4019 (N_4019,N_3600,N_3850);
nor U4020 (N_4020,N_3611,N_3708);
xnor U4021 (N_4021,N_3808,N_3853);
xor U4022 (N_4022,N_3640,N_3843);
or U4023 (N_4023,N_3864,N_3719);
and U4024 (N_4024,N_3657,N_3617);
or U4025 (N_4025,N_3840,N_3884);
nor U4026 (N_4026,N_3733,N_3736);
nand U4027 (N_4027,N_3629,N_3823);
or U4028 (N_4028,N_3740,N_3753);
or U4029 (N_4029,N_3722,N_3604);
nor U4030 (N_4030,N_3780,N_3628);
and U4031 (N_4031,N_3887,N_3830);
nand U4032 (N_4032,N_3870,N_3748);
xor U4033 (N_4033,N_3713,N_3885);
nor U4034 (N_4034,N_3847,N_3675);
and U4035 (N_4035,N_3711,N_3761);
nor U4036 (N_4036,N_3797,N_3882);
nor U4037 (N_4037,N_3603,N_3730);
or U4038 (N_4038,N_3750,N_3649);
nand U4039 (N_4039,N_3772,N_3817);
and U4040 (N_4040,N_3852,N_3775);
nor U4041 (N_4041,N_3820,N_3763);
xnor U4042 (N_4042,N_3833,N_3841);
and U4043 (N_4043,N_3878,N_3601);
nor U4044 (N_4044,N_3747,N_3726);
nand U4045 (N_4045,N_3896,N_3609);
or U4046 (N_4046,N_3672,N_3679);
nor U4047 (N_4047,N_3810,N_3632);
nor U4048 (N_4048,N_3829,N_3788);
xor U4049 (N_4049,N_3691,N_3700);
nor U4050 (N_4050,N_3634,N_3708);
nand U4051 (N_4051,N_3647,N_3723);
nor U4052 (N_4052,N_3669,N_3860);
or U4053 (N_4053,N_3719,N_3645);
xor U4054 (N_4054,N_3668,N_3802);
xor U4055 (N_4055,N_3732,N_3606);
nor U4056 (N_4056,N_3771,N_3761);
nor U4057 (N_4057,N_3698,N_3827);
nand U4058 (N_4058,N_3855,N_3893);
and U4059 (N_4059,N_3745,N_3646);
xor U4060 (N_4060,N_3609,N_3811);
or U4061 (N_4061,N_3856,N_3871);
and U4062 (N_4062,N_3656,N_3630);
nand U4063 (N_4063,N_3617,N_3815);
and U4064 (N_4064,N_3815,N_3690);
and U4065 (N_4065,N_3875,N_3847);
xor U4066 (N_4066,N_3642,N_3861);
xor U4067 (N_4067,N_3796,N_3809);
xor U4068 (N_4068,N_3823,N_3826);
or U4069 (N_4069,N_3881,N_3794);
nor U4070 (N_4070,N_3817,N_3805);
and U4071 (N_4071,N_3802,N_3899);
or U4072 (N_4072,N_3679,N_3685);
and U4073 (N_4073,N_3634,N_3702);
nor U4074 (N_4074,N_3803,N_3898);
or U4075 (N_4075,N_3822,N_3889);
and U4076 (N_4076,N_3876,N_3745);
xnor U4077 (N_4077,N_3781,N_3850);
nand U4078 (N_4078,N_3805,N_3625);
nand U4079 (N_4079,N_3776,N_3726);
or U4080 (N_4080,N_3678,N_3615);
nand U4081 (N_4081,N_3824,N_3896);
xnor U4082 (N_4082,N_3879,N_3802);
and U4083 (N_4083,N_3897,N_3605);
or U4084 (N_4084,N_3744,N_3872);
xnor U4085 (N_4085,N_3666,N_3626);
nand U4086 (N_4086,N_3622,N_3811);
nor U4087 (N_4087,N_3618,N_3830);
nor U4088 (N_4088,N_3642,N_3789);
and U4089 (N_4089,N_3694,N_3709);
nor U4090 (N_4090,N_3625,N_3655);
nand U4091 (N_4091,N_3792,N_3611);
nor U4092 (N_4092,N_3644,N_3729);
and U4093 (N_4093,N_3639,N_3773);
nand U4094 (N_4094,N_3890,N_3639);
nand U4095 (N_4095,N_3744,N_3807);
nor U4096 (N_4096,N_3673,N_3855);
and U4097 (N_4097,N_3673,N_3721);
nor U4098 (N_4098,N_3813,N_3744);
and U4099 (N_4099,N_3621,N_3635);
nand U4100 (N_4100,N_3797,N_3686);
nor U4101 (N_4101,N_3791,N_3689);
xnor U4102 (N_4102,N_3630,N_3631);
nor U4103 (N_4103,N_3748,N_3690);
and U4104 (N_4104,N_3849,N_3824);
nor U4105 (N_4105,N_3671,N_3698);
or U4106 (N_4106,N_3737,N_3864);
or U4107 (N_4107,N_3838,N_3849);
or U4108 (N_4108,N_3653,N_3638);
nand U4109 (N_4109,N_3715,N_3835);
or U4110 (N_4110,N_3893,N_3616);
nand U4111 (N_4111,N_3723,N_3875);
and U4112 (N_4112,N_3709,N_3711);
and U4113 (N_4113,N_3790,N_3636);
nand U4114 (N_4114,N_3793,N_3639);
nand U4115 (N_4115,N_3773,N_3698);
nor U4116 (N_4116,N_3867,N_3701);
or U4117 (N_4117,N_3669,N_3857);
xnor U4118 (N_4118,N_3676,N_3729);
or U4119 (N_4119,N_3833,N_3643);
nor U4120 (N_4120,N_3713,N_3721);
or U4121 (N_4121,N_3691,N_3740);
nand U4122 (N_4122,N_3638,N_3840);
xor U4123 (N_4123,N_3695,N_3702);
xor U4124 (N_4124,N_3805,N_3722);
xnor U4125 (N_4125,N_3696,N_3823);
nor U4126 (N_4126,N_3694,N_3835);
or U4127 (N_4127,N_3814,N_3879);
nor U4128 (N_4128,N_3846,N_3672);
and U4129 (N_4129,N_3702,N_3803);
or U4130 (N_4130,N_3742,N_3806);
xnor U4131 (N_4131,N_3700,N_3802);
xor U4132 (N_4132,N_3638,N_3776);
nor U4133 (N_4133,N_3676,N_3891);
or U4134 (N_4134,N_3686,N_3740);
nand U4135 (N_4135,N_3696,N_3717);
or U4136 (N_4136,N_3890,N_3817);
and U4137 (N_4137,N_3611,N_3699);
nor U4138 (N_4138,N_3621,N_3612);
xor U4139 (N_4139,N_3851,N_3833);
nor U4140 (N_4140,N_3790,N_3835);
xor U4141 (N_4141,N_3836,N_3830);
nand U4142 (N_4142,N_3855,N_3738);
or U4143 (N_4143,N_3723,N_3718);
or U4144 (N_4144,N_3610,N_3801);
or U4145 (N_4145,N_3708,N_3776);
nor U4146 (N_4146,N_3681,N_3848);
or U4147 (N_4147,N_3779,N_3606);
nand U4148 (N_4148,N_3850,N_3713);
or U4149 (N_4149,N_3742,N_3856);
or U4150 (N_4150,N_3659,N_3709);
or U4151 (N_4151,N_3823,N_3860);
xor U4152 (N_4152,N_3635,N_3876);
nand U4153 (N_4153,N_3856,N_3843);
nor U4154 (N_4154,N_3857,N_3628);
nand U4155 (N_4155,N_3620,N_3864);
nand U4156 (N_4156,N_3613,N_3815);
nand U4157 (N_4157,N_3607,N_3768);
nand U4158 (N_4158,N_3680,N_3754);
and U4159 (N_4159,N_3727,N_3825);
or U4160 (N_4160,N_3719,N_3646);
and U4161 (N_4161,N_3619,N_3831);
xnor U4162 (N_4162,N_3634,N_3772);
and U4163 (N_4163,N_3650,N_3840);
and U4164 (N_4164,N_3867,N_3829);
xnor U4165 (N_4165,N_3893,N_3674);
nor U4166 (N_4166,N_3858,N_3718);
nor U4167 (N_4167,N_3695,N_3639);
nand U4168 (N_4168,N_3816,N_3855);
xor U4169 (N_4169,N_3681,N_3649);
or U4170 (N_4170,N_3817,N_3876);
or U4171 (N_4171,N_3834,N_3822);
nand U4172 (N_4172,N_3601,N_3774);
nand U4173 (N_4173,N_3844,N_3746);
and U4174 (N_4174,N_3897,N_3757);
xor U4175 (N_4175,N_3742,N_3765);
and U4176 (N_4176,N_3761,N_3803);
nand U4177 (N_4177,N_3608,N_3804);
xor U4178 (N_4178,N_3630,N_3834);
nor U4179 (N_4179,N_3685,N_3724);
xor U4180 (N_4180,N_3810,N_3741);
xnor U4181 (N_4181,N_3763,N_3767);
nand U4182 (N_4182,N_3674,N_3680);
nand U4183 (N_4183,N_3605,N_3702);
nor U4184 (N_4184,N_3759,N_3784);
or U4185 (N_4185,N_3613,N_3871);
or U4186 (N_4186,N_3831,N_3761);
nand U4187 (N_4187,N_3818,N_3845);
nand U4188 (N_4188,N_3775,N_3689);
and U4189 (N_4189,N_3614,N_3881);
or U4190 (N_4190,N_3856,N_3704);
nor U4191 (N_4191,N_3728,N_3750);
nor U4192 (N_4192,N_3682,N_3816);
xnor U4193 (N_4193,N_3878,N_3818);
xnor U4194 (N_4194,N_3606,N_3777);
or U4195 (N_4195,N_3685,N_3769);
xnor U4196 (N_4196,N_3704,N_3675);
nand U4197 (N_4197,N_3741,N_3612);
and U4198 (N_4198,N_3744,N_3833);
xnor U4199 (N_4199,N_3763,N_3611);
nor U4200 (N_4200,N_4190,N_4015);
nand U4201 (N_4201,N_4003,N_4146);
nand U4202 (N_4202,N_4184,N_3987);
nor U4203 (N_4203,N_3910,N_4171);
nor U4204 (N_4204,N_3920,N_4187);
or U4205 (N_4205,N_4051,N_4045);
and U4206 (N_4206,N_3946,N_4151);
or U4207 (N_4207,N_4122,N_4150);
xor U4208 (N_4208,N_4042,N_3962);
nor U4209 (N_4209,N_3943,N_4070);
nand U4210 (N_4210,N_3961,N_4049);
and U4211 (N_4211,N_4170,N_4031);
nor U4212 (N_4212,N_4163,N_4054);
or U4213 (N_4213,N_4059,N_3921);
nand U4214 (N_4214,N_4176,N_4009);
nand U4215 (N_4215,N_4172,N_3908);
xnor U4216 (N_4216,N_4126,N_4188);
nand U4217 (N_4217,N_4008,N_3902);
and U4218 (N_4218,N_3918,N_4021);
and U4219 (N_4219,N_4037,N_3979);
or U4220 (N_4220,N_4086,N_4032);
nor U4221 (N_4221,N_3948,N_4127);
nor U4222 (N_4222,N_4134,N_4084);
nor U4223 (N_4223,N_4101,N_3939);
or U4224 (N_4224,N_3985,N_4061);
nor U4225 (N_4225,N_4191,N_3960);
xor U4226 (N_4226,N_3942,N_3906);
nand U4227 (N_4227,N_4073,N_4135);
and U4228 (N_4228,N_3991,N_3933);
and U4229 (N_4229,N_4067,N_4006);
xnor U4230 (N_4230,N_4131,N_4095);
nand U4231 (N_4231,N_3974,N_4169);
nor U4232 (N_4232,N_4088,N_4099);
nand U4233 (N_4233,N_4133,N_4090);
xnor U4234 (N_4234,N_4089,N_4182);
nor U4235 (N_4235,N_4155,N_4194);
or U4236 (N_4236,N_3988,N_3938);
and U4237 (N_4237,N_3953,N_3941);
nand U4238 (N_4238,N_4076,N_4192);
nand U4239 (N_4239,N_4068,N_4043);
or U4240 (N_4240,N_3975,N_4082);
xnor U4241 (N_4241,N_3931,N_3956);
or U4242 (N_4242,N_4077,N_3903);
xnor U4243 (N_4243,N_4193,N_4110);
nand U4244 (N_4244,N_4121,N_3955);
nor U4245 (N_4245,N_3925,N_3992);
xnor U4246 (N_4246,N_4039,N_3909);
nand U4247 (N_4247,N_4142,N_4013);
xnor U4248 (N_4248,N_4166,N_4103);
xor U4249 (N_4249,N_3937,N_3935);
or U4250 (N_4250,N_4114,N_3919);
or U4251 (N_4251,N_4138,N_3923);
nor U4252 (N_4252,N_3989,N_4036);
nor U4253 (N_4253,N_3994,N_4041);
or U4254 (N_4254,N_4012,N_3949);
xor U4255 (N_4255,N_3978,N_3922);
xnor U4256 (N_4256,N_4152,N_3957);
nand U4257 (N_4257,N_4034,N_3976);
nor U4258 (N_4258,N_3998,N_4112);
and U4259 (N_4259,N_4143,N_4145);
and U4260 (N_4260,N_4071,N_3984);
nor U4261 (N_4261,N_3914,N_3940);
and U4262 (N_4262,N_4024,N_4100);
or U4263 (N_4263,N_3905,N_4074);
xnor U4264 (N_4264,N_4018,N_3970);
and U4265 (N_4265,N_3916,N_4029);
nand U4266 (N_4266,N_3969,N_4186);
xnor U4267 (N_4267,N_4026,N_4157);
or U4268 (N_4268,N_4149,N_3934);
or U4269 (N_4269,N_4047,N_4053);
nor U4270 (N_4270,N_4109,N_4046);
nor U4271 (N_4271,N_4102,N_4028);
nor U4272 (N_4272,N_3930,N_4132);
nor U4273 (N_4273,N_4130,N_4107);
nor U4274 (N_4274,N_3911,N_4069);
nor U4275 (N_4275,N_4137,N_4136);
nor U4276 (N_4276,N_3980,N_4123);
xor U4277 (N_4277,N_4104,N_4196);
or U4278 (N_4278,N_3965,N_4129);
nor U4279 (N_4279,N_4128,N_4162);
nor U4280 (N_4280,N_4033,N_4080);
and U4281 (N_4281,N_4173,N_3981);
and U4282 (N_4282,N_3993,N_3977);
nor U4283 (N_4283,N_4183,N_3959);
nor U4284 (N_4284,N_3954,N_4139);
nand U4285 (N_4285,N_4017,N_4000);
and U4286 (N_4286,N_4091,N_4010);
nor U4287 (N_4287,N_4081,N_4087);
xnor U4288 (N_4288,N_3968,N_3966);
nand U4289 (N_4289,N_4085,N_4159);
nor U4290 (N_4290,N_4165,N_4199);
and U4291 (N_4291,N_3929,N_4167);
nand U4292 (N_4292,N_3982,N_4058);
nand U4293 (N_4293,N_4065,N_4001);
and U4294 (N_4294,N_4140,N_4092);
and U4295 (N_4295,N_4118,N_3983);
or U4296 (N_4296,N_4063,N_4156);
or U4297 (N_4297,N_4105,N_4016);
nand U4298 (N_4298,N_4004,N_4083);
or U4299 (N_4299,N_3945,N_4055);
nor U4300 (N_4300,N_4161,N_3973);
nor U4301 (N_4301,N_4064,N_4005);
nand U4302 (N_4302,N_3944,N_3901);
or U4303 (N_4303,N_3951,N_4189);
nor U4304 (N_4304,N_4197,N_4062);
and U4305 (N_4305,N_4124,N_4175);
nor U4306 (N_4306,N_4060,N_3995);
xor U4307 (N_4307,N_4030,N_4177);
or U4308 (N_4308,N_4106,N_3924);
and U4309 (N_4309,N_4025,N_4050);
xor U4310 (N_4310,N_4115,N_3936);
and U4311 (N_4311,N_4164,N_4160);
or U4312 (N_4312,N_3904,N_4044);
or U4313 (N_4313,N_4111,N_4093);
xor U4314 (N_4314,N_3986,N_4116);
nand U4315 (N_4315,N_4078,N_3932);
nor U4316 (N_4316,N_3915,N_4108);
or U4317 (N_4317,N_4185,N_4040);
or U4318 (N_4318,N_3927,N_4098);
xor U4319 (N_4319,N_4180,N_4148);
and U4320 (N_4320,N_4096,N_4168);
or U4321 (N_4321,N_4014,N_4141);
xor U4322 (N_4322,N_3971,N_3952);
or U4323 (N_4323,N_3926,N_4048);
nor U4324 (N_4324,N_4057,N_3996);
nand U4325 (N_4325,N_4181,N_4020);
or U4326 (N_4326,N_4153,N_4079);
nor U4327 (N_4327,N_4154,N_4022);
or U4328 (N_4328,N_3999,N_3928);
nor U4329 (N_4329,N_3964,N_4120);
nand U4330 (N_4330,N_4158,N_4125);
or U4331 (N_4331,N_3917,N_4027);
or U4332 (N_4332,N_4011,N_4002);
nand U4333 (N_4333,N_4097,N_4066);
and U4334 (N_4334,N_3907,N_4094);
or U4335 (N_4335,N_4117,N_4198);
nor U4336 (N_4336,N_4179,N_4056);
xnor U4337 (N_4337,N_3950,N_3912);
nor U4338 (N_4338,N_4119,N_3947);
nor U4339 (N_4339,N_3997,N_4144);
or U4340 (N_4340,N_4019,N_4075);
xnor U4341 (N_4341,N_3900,N_4038);
nand U4342 (N_4342,N_4007,N_4174);
and U4343 (N_4343,N_3990,N_4072);
nand U4344 (N_4344,N_3967,N_3958);
xnor U4345 (N_4345,N_4178,N_4023);
or U4346 (N_4346,N_3963,N_4113);
and U4347 (N_4347,N_3913,N_4147);
xnor U4348 (N_4348,N_4195,N_4052);
and U4349 (N_4349,N_4035,N_3972);
or U4350 (N_4350,N_4134,N_4058);
nor U4351 (N_4351,N_3984,N_3921);
and U4352 (N_4352,N_3932,N_4152);
and U4353 (N_4353,N_4068,N_4114);
nor U4354 (N_4354,N_4073,N_3966);
or U4355 (N_4355,N_4051,N_4124);
or U4356 (N_4356,N_4181,N_4155);
xor U4357 (N_4357,N_3998,N_4082);
nand U4358 (N_4358,N_3982,N_4092);
xnor U4359 (N_4359,N_3970,N_3994);
and U4360 (N_4360,N_3999,N_4149);
xor U4361 (N_4361,N_3980,N_4183);
nand U4362 (N_4362,N_3902,N_4037);
xnor U4363 (N_4363,N_4026,N_4154);
xor U4364 (N_4364,N_3991,N_3941);
or U4365 (N_4365,N_3979,N_4175);
or U4366 (N_4366,N_4053,N_4061);
nand U4367 (N_4367,N_4072,N_4067);
nand U4368 (N_4368,N_4172,N_3929);
xnor U4369 (N_4369,N_3963,N_4147);
and U4370 (N_4370,N_4000,N_3970);
and U4371 (N_4371,N_4183,N_4028);
xnor U4372 (N_4372,N_4054,N_4051);
and U4373 (N_4373,N_4005,N_3964);
nand U4374 (N_4374,N_3954,N_3937);
xnor U4375 (N_4375,N_3975,N_4114);
nand U4376 (N_4376,N_4036,N_4121);
or U4377 (N_4377,N_4110,N_4146);
or U4378 (N_4378,N_4035,N_4147);
xor U4379 (N_4379,N_4034,N_4126);
or U4380 (N_4380,N_4072,N_4145);
nand U4381 (N_4381,N_4129,N_4077);
xnor U4382 (N_4382,N_4075,N_4093);
or U4383 (N_4383,N_4046,N_4102);
nor U4384 (N_4384,N_4068,N_3967);
or U4385 (N_4385,N_4145,N_4178);
nor U4386 (N_4386,N_3921,N_3963);
or U4387 (N_4387,N_4096,N_3993);
or U4388 (N_4388,N_3958,N_3937);
nor U4389 (N_4389,N_3992,N_4005);
and U4390 (N_4390,N_4171,N_4077);
nand U4391 (N_4391,N_4182,N_3949);
nor U4392 (N_4392,N_4060,N_4180);
nor U4393 (N_4393,N_4150,N_4154);
xnor U4394 (N_4394,N_4143,N_4114);
nand U4395 (N_4395,N_4029,N_3938);
xnor U4396 (N_4396,N_3994,N_3995);
nor U4397 (N_4397,N_3923,N_4195);
or U4398 (N_4398,N_3932,N_4048);
or U4399 (N_4399,N_3948,N_3975);
nand U4400 (N_4400,N_4086,N_4069);
xnor U4401 (N_4401,N_4074,N_3947);
xor U4402 (N_4402,N_4018,N_4109);
xnor U4403 (N_4403,N_4048,N_4007);
or U4404 (N_4404,N_4196,N_4103);
nor U4405 (N_4405,N_4140,N_3973);
and U4406 (N_4406,N_3992,N_4145);
or U4407 (N_4407,N_4031,N_4092);
nand U4408 (N_4408,N_3985,N_4032);
and U4409 (N_4409,N_3939,N_4109);
nand U4410 (N_4410,N_4155,N_4197);
xnor U4411 (N_4411,N_3917,N_4067);
nand U4412 (N_4412,N_3942,N_3916);
nor U4413 (N_4413,N_4117,N_4176);
or U4414 (N_4414,N_3989,N_3908);
nor U4415 (N_4415,N_4052,N_4093);
and U4416 (N_4416,N_4096,N_4003);
nand U4417 (N_4417,N_4077,N_3957);
or U4418 (N_4418,N_4081,N_3926);
nand U4419 (N_4419,N_4034,N_4042);
nand U4420 (N_4420,N_4041,N_4129);
or U4421 (N_4421,N_4167,N_3966);
nor U4422 (N_4422,N_4002,N_4061);
xor U4423 (N_4423,N_4032,N_4195);
and U4424 (N_4424,N_3958,N_4148);
xor U4425 (N_4425,N_4143,N_4141);
or U4426 (N_4426,N_4136,N_4025);
or U4427 (N_4427,N_3952,N_4146);
or U4428 (N_4428,N_4045,N_4142);
xor U4429 (N_4429,N_4139,N_4033);
nor U4430 (N_4430,N_4160,N_3937);
or U4431 (N_4431,N_4198,N_3972);
nor U4432 (N_4432,N_4147,N_4198);
xnor U4433 (N_4433,N_4182,N_3970);
and U4434 (N_4434,N_4118,N_4143);
nand U4435 (N_4435,N_4187,N_3965);
nand U4436 (N_4436,N_4077,N_3985);
nor U4437 (N_4437,N_3982,N_4020);
nor U4438 (N_4438,N_4105,N_4178);
and U4439 (N_4439,N_4094,N_4014);
xor U4440 (N_4440,N_3932,N_4036);
or U4441 (N_4441,N_3920,N_4099);
nor U4442 (N_4442,N_4014,N_4032);
or U4443 (N_4443,N_4103,N_4165);
nor U4444 (N_4444,N_4005,N_4000);
or U4445 (N_4445,N_4139,N_4058);
xnor U4446 (N_4446,N_4035,N_3965);
nor U4447 (N_4447,N_4101,N_3912);
nor U4448 (N_4448,N_4197,N_4079);
and U4449 (N_4449,N_4028,N_3930);
nor U4450 (N_4450,N_3997,N_4120);
or U4451 (N_4451,N_3977,N_4080);
and U4452 (N_4452,N_3942,N_4015);
nor U4453 (N_4453,N_4193,N_4125);
and U4454 (N_4454,N_4182,N_4051);
and U4455 (N_4455,N_4031,N_3995);
xnor U4456 (N_4456,N_4017,N_4030);
and U4457 (N_4457,N_4076,N_3929);
nor U4458 (N_4458,N_3918,N_3986);
or U4459 (N_4459,N_3922,N_4081);
and U4460 (N_4460,N_4050,N_3921);
xnor U4461 (N_4461,N_4180,N_4057);
and U4462 (N_4462,N_3987,N_3917);
and U4463 (N_4463,N_4006,N_4073);
or U4464 (N_4464,N_4045,N_4029);
xnor U4465 (N_4465,N_4052,N_4013);
nand U4466 (N_4466,N_4067,N_4057);
nor U4467 (N_4467,N_3979,N_3911);
and U4468 (N_4468,N_4179,N_4159);
xnor U4469 (N_4469,N_3927,N_4025);
nand U4470 (N_4470,N_4172,N_4041);
or U4471 (N_4471,N_3997,N_4159);
nand U4472 (N_4472,N_3934,N_4084);
or U4473 (N_4473,N_4147,N_4073);
nand U4474 (N_4474,N_4177,N_4075);
xnor U4475 (N_4475,N_3919,N_3907);
nor U4476 (N_4476,N_4098,N_3994);
nor U4477 (N_4477,N_3996,N_4114);
and U4478 (N_4478,N_4069,N_3936);
and U4479 (N_4479,N_3963,N_4099);
or U4480 (N_4480,N_4118,N_4114);
xor U4481 (N_4481,N_3971,N_4199);
xor U4482 (N_4482,N_3963,N_3993);
xor U4483 (N_4483,N_4101,N_4155);
nand U4484 (N_4484,N_4190,N_4048);
or U4485 (N_4485,N_4034,N_4051);
or U4486 (N_4486,N_3947,N_4086);
nand U4487 (N_4487,N_3946,N_3997);
nor U4488 (N_4488,N_4066,N_4073);
xnor U4489 (N_4489,N_4060,N_3991);
nand U4490 (N_4490,N_4126,N_4060);
nand U4491 (N_4491,N_4083,N_3908);
nand U4492 (N_4492,N_4037,N_3932);
and U4493 (N_4493,N_4180,N_4049);
nand U4494 (N_4494,N_3973,N_4107);
nor U4495 (N_4495,N_4053,N_4100);
and U4496 (N_4496,N_3963,N_3923);
nand U4497 (N_4497,N_4035,N_4106);
or U4498 (N_4498,N_3987,N_4110);
and U4499 (N_4499,N_3966,N_4012);
nand U4500 (N_4500,N_4313,N_4464);
nor U4501 (N_4501,N_4367,N_4370);
nand U4502 (N_4502,N_4491,N_4223);
and U4503 (N_4503,N_4454,N_4272);
xor U4504 (N_4504,N_4455,N_4387);
or U4505 (N_4505,N_4280,N_4218);
xor U4506 (N_4506,N_4214,N_4257);
nand U4507 (N_4507,N_4476,N_4470);
and U4508 (N_4508,N_4279,N_4399);
xnor U4509 (N_4509,N_4406,N_4262);
or U4510 (N_4510,N_4232,N_4288);
and U4511 (N_4511,N_4376,N_4267);
and U4512 (N_4512,N_4353,N_4445);
and U4513 (N_4513,N_4438,N_4215);
nand U4514 (N_4514,N_4447,N_4497);
or U4515 (N_4515,N_4268,N_4263);
xor U4516 (N_4516,N_4326,N_4322);
xor U4517 (N_4517,N_4243,N_4248);
nor U4518 (N_4518,N_4211,N_4308);
and U4519 (N_4519,N_4297,N_4256);
nand U4520 (N_4520,N_4207,N_4479);
or U4521 (N_4521,N_4361,N_4221);
nand U4522 (N_4522,N_4316,N_4246);
or U4523 (N_4523,N_4385,N_4252);
nand U4524 (N_4524,N_4286,N_4315);
and U4525 (N_4525,N_4443,N_4337);
or U4526 (N_4526,N_4465,N_4359);
nor U4527 (N_4527,N_4331,N_4425);
and U4528 (N_4528,N_4404,N_4349);
nand U4529 (N_4529,N_4436,N_4206);
and U4530 (N_4530,N_4369,N_4449);
nand U4531 (N_4531,N_4383,N_4453);
nor U4532 (N_4532,N_4309,N_4451);
nand U4533 (N_4533,N_4356,N_4234);
nor U4534 (N_4534,N_4224,N_4293);
nor U4535 (N_4535,N_4238,N_4499);
and U4536 (N_4536,N_4466,N_4396);
or U4537 (N_4537,N_4490,N_4474);
xnor U4538 (N_4538,N_4434,N_4420);
nor U4539 (N_4539,N_4446,N_4303);
and U4540 (N_4540,N_4304,N_4384);
nand U4541 (N_4541,N_4249,N_4422);
nand U4542 (N_4542,N_4428,N_4273);
xor U4543 (N_4543,N_4284,N_4358);
xnor U4544 (N_4544,N_4324,N_4202);
nand U4545 (N_4545,N_4365,N_4299);
xnor U4546 (N_4546,N_4336,N_4258);
or U4547 (N_4547,N_4203,N_4416);
xor U4548 (N_4548,N_4329,N_4302);
nand U4549 (N_4549,N_4255,N_4220);
nand U4550 (N_4550,N_4435,N_4318);
xor U4551 (N_4551,N_4333,N_4291);
nand U4552 (N_4552,N_4362,N_4292);
nand U4553 (N_4553,N_4397,N_4418);
nand U4554 (N_4554,N_4317,N_4282);
nor U4555 (N_4555,N_4244,N_4250);
nand U4556 (N_4556,N_4412,N_4261);
and U4557 (N_4557,N_4290,N_4419);
or U4558 (N_4558,N_4401,N_4495);
and U4559 (N_4559,N_4378,N_4323);
nor U4560 (N_4560,N_4433,N_4442);
nor U4561 (N_4561,N_4368,N_4482);
or U4562 (N_4562,N_4450,N_4347);
nor U4563 (N_4563,N_4265,N_4469);
nand U4564 (N_4564,N_4216,N_4366);
or U4565 (N_4565,N_4415,N_4269);
nor U4566 (N_4566,N_4372,N_4287);
nor U4567 (N_4567,N_4311,N_4254);
or U4568 (N_4568,N_4364,N_4374);
nand U4569 (N_4569,N_4410,N_4431);
and U4570 (N_4570,N_4421,N_4334);
or U4571 (N_4571,N_4430,N_4320);
and U4572 (N_4572,N_4295,N_4427);
nand U4573 (N_4573,N_4205,N_4237);
nand U4574 (N_4574,N_4266,N_4457);
nand U4575 (N_4575,N_4306,N_4341);
nand U4576 (N_4576,N_4325,N_4448);
nand U4577 (N_4577,N_4228,N_4283);
or U4578 (N_4578,N_4225,N_4432);
or U4579 (N_4579,N_4312,N_4231);
nor U4580 (N_4580,N_4478,N_4350);
or U4581 (N_4581,N_4407,N_4363);
nand U4582 (N_4582,N_4354,N_4245);
and U4583 (N_4583,N_4371,N_4239);
or U4584 (N_4584,N_4296,N_4226);
and U4585 (N_4585,N_4379,N_4242);
and U4586 (N_4586,N_4417,N_4227);
and U4587 (N_4587,N_4241,N_4305);
nand U4588 (N_4588,N_4314,N_4213);
and U4589 (N_4589,N_4204,N_4332);
nand U4590 (N_4590,N_4395,N_4480);
or U4591 (N_4591,N_4328,N_4209);
nor U4592 (N_4592,N_4392,N_4487);
nand U4593 (N_4593,N_4408,N_4230);
and U4594 (N_4594,N_4473,N_4348);
nor U4595 (N_4595,N_4467,N_4437);
nand U4596 (N_4596,N_4319,N_4452);
xnor U4597 (N_4597,N_4461,N_4253);
or U4598 (N_4598,N_4298,N_4310);
xnor U4599 (N_4599,N_4471,N_4342);
nor U4600 (N_4600,N_4389,N_4247);
xor U4601 (N_4601,N_4496,N_4259);
nand U4602 (N_4602,N_4468,N_4498);
or U4603 (N_4603,N_4278,N_4210);
and U4604 (N_4604,N_4441,N_4338);
and U4605 (N_4605,N_4346,N_4380);
xor U4606 (N_4606,N_4403,N_4274);
xnor U4607 (N_4607,N_4373,N_4251);
xor U4608 (N_4608,N_4413,N_4344);
nor U4609 (N_4609,N_4382,N_4472);
nand U4610 (N_4610,N_4330,N_4294);
xnor U4611 (N_4611,N_4388,N_4477);
nor U4612 (N_4612,N_4393,N_4307);
nand U4613 (N_4613,N_4456,N_4201);
xnor U4614 (N_4614,N_4212,N_4300);
nand U4615 (N_4615,N_4475,N_4377);
or U4616 (N_4616,N_4460,N_4481);
and U4617 (N_4617,N_4277,N_4405);
xor U4618 (N_4618,N_4208,N_4381);
nor U4619 (N_4619,N_4375,N_4285);
or U4620 (N_4620,N_4235,N_4343);
nor U4621 (N_4621,N_4335,N_4494);
nand U4622 (N_4622,N_4394,N_4345);
nor U4623 (N_4623,N_4357,N_4236);
xnor U4624 (N_4624,N_4409,N_4264);
xnor U4625 (N_4625,N_4462,N_4458);
or U4626 (N_4626,N_4327,N_4483);
or U4627 (N_4627,N_4400,N_4423);
nand U4628 (N_4628,N_4429,N_4492);
xor U4629 (N_4629,N_4355,N_4402);
xnor U4630 (N_4630,N_4222,N_4391);
nand U4631 (N_4631,N_4289,N_4352);
and U4632 (N_4632,N_4270,N_4233);
xor U4633 (N_4633,N_4281,N_4489);
or U4634 (N_4634,N_4240,N_4484);
nand U4635 (N_4635,N_4275,N_4459);
nand U4636 (N_4636,N_4351,N_4424);
nand U4637 (N_4637,N_4229,N_4440);
nand U4638 (N_4638,N_4276,N_4426);
and U4639 (N_4639,N_4463,N_4493);
or U4640 (N_4640,N_4439,N_4386);
and U4641 (N_4641,N_4217,N_4219);
and U4642 (N_4642,N_4485,N_4411);
and U4643 (N_4643,N_4271,N_4398);
or U4644 (N_4644,N_4444,N_4301);
nor U4645 (N_4645,N_4200,N_4488);
xor U4646 (N_4646,N_4414,N_4260);
or U4647 (N_4647,N_4339,N_4360);
nor U4648 (N_4648,N_4340,N_4390);
xor U4649 (N_4649,N_4486,N_4321);
or U4650 (N_4650,N_4497,N_4202);
nand U4651 (N_4651,N_4409,N_4211);
nand U4652 (N_4652,N_4230,N_4312);
nand U4653 (N_4653,N_4356,N_4266);
nand U4654 (N_4654,N_4358,N_4441);
xnor U4655 (N_4655,N_4401,N_4413);
nor U4656 (N_4656,N_4456,N_4277);
and U4657 (N_4657,N_4457,N_4359);
or U4658 (N_4658,N_4340,N_4252);
xnor U4659 (N_4659,N_4308,N_4361);
or U4660 (N_4660,N_4418,N_4476);
or U4661 (N_4661,N_4367,N_4463);
nor U4662 (N_4662,N_4277,N_4373);
nand U4663 (N_4663,N_4304,N_4489);
nand U4664 (N_4664,N_4304,N_4378);
nor U4665 (N_4665,N_4255,N_4365);
nor U4666 (N_4666,N_4426,N_4255);
xnor U4667 (N_4667,N_4217,N_4475);
and U4668 (N_4668,N_4227,N_4449);
nor U4669 (N_4669,N_4351,N_4245);
and U4670 (N_4670,N_4246,N_4227);
or U4671 (N_4671,N_4338,N_4224);
nor U4672 (N_4672,N_4413,N_4292);
and U4673 (N_4673,N_4331,N_4273);
xnor U4674 (N_4674,N_4293,N_4351);
nor U4675 (N_4675,N_4395,N_4235);
xor U4676 (N_4676,N_4327,N_4352);
nand U4677 (N_4677,N_4321,N_4364);
or U4678 (N_4678,N_4233,N_4495);
xor U4679 (N_4679,N_4228,N_4281);
nand U4680 (N_4680,N_4439,N_4350);
or U4681 (N_4681,N_4229,N_4218);
nand U4682 (N_4682,N_4427,N_4345);
nand U4683 (N_4683,N_4421,N_4314);
or U4684 (N_4684,N_4268,N_4312);
xor U4685 (N_4685,N_4334,N_4294);
nor U4686 (N_4686,N_4489,N_4490);
or U4687 (N_4687,N_4222,N_4471);
xnor U4688 (N_4688,N_4279,N_4307);
nor U4689 (N_4689,N_4230,N_4300);
and U4690 (N_4690,N_4404,N_4287);
nand U4691 (N_4691,N_4206,N_4453);
nand U4692 (N_4692,N_4331,N_4342);
or U4693 (N_4693,N_4417,N_4239);
nand U4694 (N_4694,N_4415,N_4247);
or U4695 (N_4695,N_4485,N_4364);
nand U4696 (N_4696,N_4234,N_4430);
nor U4697 (N_4697,N_4236,N_4271);
nor U4698 (N_4698,N_4400,N_4341);
nand U4699 (N_4699,N_4398,N_4227);
and U4700 (N_4700,N_4296,N_4493);
nor U4701 (N_4701,N_4488,N_4293);
nand U4702 (N_4702,N_4432,N_4276);
xor U4703 (N_4703,N_4223,N_4203);
and U4704 (N_4704,N_4201,N_4397);
or U4705 (N_4705,N_4316,N_4227);
nor U4706 (N_4706,N_4378,N_4485);
or U4707 (N_4707,N_4489,N_4403);
nand U4708 (N_4708,N_4298,N_4329);
xnor U4709 (N_4709,N_4377,N_4384);
nor U4710 (N_4710,N_4439,N_4304);
xnor U4711 (N_4711,N_4407,N_4300);
xnor U4712 (N_4712,N_4399,N_4270);
xnor U4713 (N_4713,N_4338,N_4291);
xnor U4714 (N_4714,N_4219,N_4332);
and U4715 (N_4715,N_4216,N_4350);
xor U4716 (N_4716,N_4327,N_4210);
nand U4717 (N_4717,N_4419,N_4375);
xnor U4718 (N_4718,N_4352,N_4316);
and U4719 (N_4719,N_4461,N_4232);
nor U4720 (N_4720,N_4457,N_4462);
and U4721 (N_4721,N_4324,N_4441);
xor U4722 (N_4722,N_4314,N_4251);
nor U4723 (N_4723,N_4320,N_4331);
xor U4724 (N_4724,N_4228,N_4463);
nand U4725 (N_4725,N_4246,N_4239);
xor U4726 (N_4726,N_4459,N_4202);
xor U4727 (N_4727,N_4235,N_4391);
and U4728 (N_4728,N_4496,N_4219);
xnor U4729 (N_4729,N_4214,N_4260);
nand U4730 (N_4730,N_4234,N_4483);
or U4731 (N_4731,N_4485,N_4312);
or U4732 (N_4732,N_4230,N_4478);
nor U4733 (N_4733,N_4453,N_4425);
or U4734 (N_4734,N_4279,N_4309);
and U4735 (N_4735,N_4265,N_4374);
nor U4736 (N_4736,N_4321,N_4427);
nand U4737 (N_4737,N_4253,N_4434);
and U4738 (N_4738,N_4245,N_4272);
xnor U4739 (N_4739,N_4474,N_4377);
or U4740 (N_4740,N_4489,N_4373);
nor U4741 (N_4741,N_4389,N_4447);
or U4742 (N_4742,N_4444,N_4278);
nor U4743 (N_4743,N_4264,N_4462);
nor U4744 (N_4744,N_4344,N_4226);
and U4745 (N_4745,N_4450,N_4249);
xor U4746 (N_4746,N_4314,N_4245);
nor U4747 (N_4747,N_4310,N_4489);
nor U4748 (N_4748,N_4381,N_4490);
and U4749 (N_4749,N_4432,N_4285);
xor U4750 (N_4750,N_4211,N_4216);
xor U4751 (N_4751,N_4318,N_4212);
nor U4752 (N_4752,N_4339,N_4273);
xnor U4753 (N_4753,N_4236,N_4470);
nor U4754 (N_4754,N_4320,N_4243);
and U4755 (N_4755,N_4325,N_4242);
nor U4756 (N_4756,N_4333,N_4433);
or U4757 (N_4757,N_4353,N_4425);
and U4758 (N_4758,N_4427,N_4475);
or U4759 (N_4759,N_4296,N_4215);
xor U4760 (N_4760,N_4492,N_4300);
or U4761 (N_4761,N_4417,N_4260);
or U4762 (N_4762,N_4251,N_4297);
nand U4763 (N_4763,N_4379,N_4212);
xor U4764 (N_4764,N_4339,N_4262);
and U4765 (N_4765,N_4292,N_4210);
nor U4766 (N_4766,N_4499,N_4386);
and U4767 (N_4767,N_4232,N_4327);
and U4768 (N_4768,N_4215,N_4434);
xnor U4769 (N_4769,N_4338,N_4492);
nand U4770 (N_4770,N_4480,N_4230);
xnor U4771 (N_4771,N_4444,N_4335);
xor U4772 (N_4772,N_4445,N_4407);
and U4773 (N_4773,N_4330,N_4466);
and U4774 (N_4774,N_4201,N_4308);
nand U4775 (N_4775,N_4293,N_4424);
nor U4776 (N_4776,N_4263,N_4423);
xnor U4777 (N_4777,N_4477,N_4464);
xnor U4778 (N_4778,N_4433,N_4218);
xnor U4779 (N_4779,N_4269,N_4273);
nand U4780 (N_4780,N_4375,N_4495);
or U4781 (N_4781,N_4243,N_4382);
nor U4782 (N_4782,N_4459,N_4376);
and U4783 (N_4783,N_4368,N_4454);
and U4784 (N_4784,N_4496,N_4265);
or U4785 (N_4785,N_4337,N_4263);
nand U4786 (N_4786,N_4330,N_4430);
and U4787 (N_4787,N_4497,N_4441);
and U4788 (N_4788,N_4482,N_4441);
nor U4789 (N_4789,N_4488,N_4276);
or U4790 (N_4790,N_4367,N_4459);
nor U4791 (N_4791,N_4411,N_4434);
or U4792 (N_4792,N_4333,N_4232);
nor U4793 (N_4793,N_4293,N_4470);
or U4794 (N_4794,N_4249,N_4230);
nand U4795 (N_4795,N_4447,N_4254);
nor U4796 (N_4796,N_4253,N_4241);
and U4797 (N_4797,N_4308,N_4322);
xnor U4798 (N_4798,N_4498,N_4352);
nand U4799 (N_4799,N_4439,N_4239);
nor U4800 (N_4800,N_4715,N_4503);
or U4801 (N_4801,N_4607,N_4554);
or U4802 (N_4802,N_4587,N_4604);
or U4803 (N_4803,N_4500,N_4752);
xnor U4804 (N_4804,N_4623,N_4627);
xor U4805 (N_4805,N_4726,N_4541);
nor U4806 (N_4806,N_4513,N_4617);
nor U4807 (N_4807,N_4717,N_4711);
nor U4808 (N_4808,N_4507,N_4687);
or U4809 (N_4809,N_4703,N_4534);
and U4810 (N_4810,N_4666,N_4619);
nand U4811 (N_4811,N_4505,N_4542);
xnor U4812 (N_4812,N_4594,N_4519);
nand U4813 (N_4813,N_4560,N_4664);
and U4814 (N_4814,N_4732,N_4581);
nand U4815 (N_4815,N_4660,N_4684);
xnor U4816 (N_4816,N_4657,N_4598);
nor U4817 (N_4817,N_4725,N_4646);
or U4818 (N_4818,N_4788,N_4522);
or U4819 (N_4819,N_4792,N_4536);
nor U4820 (N_4820,N_4764,N_4766);
and U4821 (N_4821,N_4548,N_4694);
xnor U4822 (N_4822,N_4525,N_4596);
nor U4823 (N_4823,N_4678,N_4670);
nor U4824 (N_4824,N_4680,N_4663);
or U4825 (N_4825,N_4693,N_4515);
or U4826 (N_4826,N_4669,N_4785);
or U4827 (N_4827,N_4665,N_4586);
nand U4828 (N_4828,N_4798,N_4674);
nor U4829 (N_4829,N_4620,N_4603);
xor U4830 (N_4830,N_4577,N_4616);
xnor U4831 (N_4831,N_4574,N_4751);
and U4832 (N_4832,N_4593,N_4566);
xnor U4833 (N_4833,N_4786,N_4533);
or U4834 (N_4834,N_4641,N_4777);
nor U4835 (N_4835,N_4696,N_4568);
nand U4836 (N_4836,N_4701,N_4565);
nor U4837 (N_4837,N_4748,N_4768);
and U4838 (N_4838,N_4625,N_4704);
xor U4839 (N_4839,N_4501,N_4649);
or U4840 (N_4840,N_4775,N_4773);
nand U4841 (N_4841,N_4799,N_4588);
or U4842 (N_4842,N_4614,N_4563);
xor U4843 (N_4843,N_4762,N_4747);
nor U4844 (N_4844,N_4714,N_4545);
or U4845 (N_4845,N_4727,N_4564);
or U4846 (N_4846,N_4592,N_4784);
nor U4847 (N_4847,N_4636,N_4612);
nand U4848 (N_4848,N_4742,N_4638);
xnor U4849 (N_4849,N_4756,N_4540);
or U4850 (N_4850,N_4644,N_4793);
or U4851 (N_4851,N_4647,N_4672);
nand U4852 (N_4852,N_4658,N_4632);
nand U4853 (N_4853,N_4523,N_4713);
nand U4854 (N_4854,N_4512,N_4723);
nor U4855 (N_4855,N_4730,N_4610);
xnor U4856 (N_4856,N_4530,N_4741);
nor U4857 (N_4857,N_4561,N_4502);
and U4858 (N_4858,N_4575,N_4780);
nand U4859 (N_4859,N_4640,N_4746);
and U4860 (N_4860,N_4739,N_4705);
and U4861 (N_4861,N_4570,N_4744);
or U4862 (N_4862,N_4690,N_4759);
nand U4863 (N_4863,N_4676,N_4552);
and U4864 (N_4864,N_4655,N_4633);
xor U4865 (N_4865,N_4510,N_4683);
xnor U4866 (N_4866,N_4685,N_4506);
nor U4867 (N_4867,N_4582,N_4584);
nand U4868 (N_4868,N_4629,N_4659);
nor U4869 (N_4869,N_4553,N_4547);
nor U4870 (N_4870,N_4735,N_4538);
and U4871 (N_4871,N_4535,N_4543);
nor U4872 (N_4872,N_4527,N_4528);
xnor U4873 (N_4873,N_4615,N_4776);
xor U4874 (N_4874,N_4681,N_4662);
xnor U4875 (N_4875,N_4661,N_4520);
or U4876 (N_4876,N_4710,N_4731);
xor U4877 (N_4877,N_4763,N_4743);
or U4878 (N_4878,N_4760,N_4618);
nand U4879 (N_4879,N_4645,N_4637);
nor U4880 (N_4880,N_4771,N_4611);
and U4881 (N_4881,N_4537,N_4772);
or U4882 (N_4882,N_4787,N_4555);
xor U4883 (N_4883,N_4654,N_4708);
and U4884 (N_4884,N_4609,N_4740);
nand U4885 (N_4885,N_4724,N_4608);
xnor U4886 (N_4886,N_4692,N_4562);
or U4887 (N_4887,N_4778,N_4688);
and U4888 (N_4888,N_4738,N_4765);
or U4889 (N_4889,N_4511,N_4729);
nor U4890 (N_4890,N_4757,N_4558);
xnor U4891 (N_4891,N_4745,N_4628);
nand U4892 (N_4892,N_4700,N_4789);
nand U4893 (N_4893,N_4576,N_4585);
and U4894 (N_4894,N_4557,N_4597);
xnor U4895 (N_4895,N_4544,N_4516);
and U4896 (N_4896,N_4599,N_4781);
or U4897 (N_4897,N_4758,N_4613);
or U4898 (N_4898,N_4769,N_4720);
or U4899 (N_4899,N_4634,N_4737);
nor U4900 (N_4900,N_4753,N_4567);
nand U4901 (N_4901,N_4754,N_4718);
nor U4902 (N_4902,N_4795,N_4571);
nor U4903 (N_4903,N_4712,N_4755);
nor U4904 (N_4904,N_4702,N_4642);
xnor U4905 (N_4905,N_4695,N_4546);
and U4906 (N_4906,N_4650,N_4606);
xor U4907 (N_4907,N_4697,N_4509);
nor U4908 (N_4908,N_4569,N_4668);
or U4909 (N_4909,N_4539,N_4689);
nand U4910 (N_4910,N_4529,N_4526);
nor U4911 (N_4911,N_4635,N_4589);
or U4912 (N_4912,N_4602,N_4677);
or U4913 (N_4913,N_4691,N_4648);
and U4914 (N_4914,N_4622,N_4524);
nor U4915 (N_4915,N_4631,N_4782);
and U4916 (N_4916,N_4699,N_4770);
or U4917 (N_4917,N_4774,N_4779);
or U4918 (N_4918,N_4508,N_4595);
or U4919 (N_4919,N_4621,N_4749);
or U4920 (N_4920,N_4791,N_4532);
nor U4921 (N_4921,N_4686,N_4790);
nor U4922 (N_4922,N_4590,N_4796);
nand U4923 (N_4923,N_4578,N_4504);
xor U4924 (N_4924,N_4709,N_4656);
nand U4925 (N_4925,N_4531,N_4736);
and U4926 (N_4926,N_4728,N_4783);
or U4927 (N_4927,N_4698,N_4794);
and U4928 (N_4928,N_4722,N_4682);
nand U4929 (N_4929,N_4716,N_4630);
and U4930 (N_4930,N_4675,N_4750);
xor U4931 (N_4931,N_4733,N_4583);
or U4932 (N_4932,N_4572,N_4626);
nor U4933 (N_4933,N_4579,N_4521);
xor U4934 (N_4934,N_4671,N_4679);
nor U4935 (N_4935,N_4667,N_4573);
and U4936 (N_4936,N_4600,N_4517);
or U4937 (N_4937,N_4721,N_4707);
or U4938 (N_4938,N_4719,N_4673);
or U4939 (N_4939,N_4601,N_4797);
nand U4940 (N_4940,N_4643,N_4639);
nand U4941 (N_4941,N_4559,N_4653);
xor U4942 (N_4942,N_4549,N_4652);
and U4943 (N_4943,N_4651,N_4767);
and U4944 (N_4944,N_4518,N_4556);
nor U4945 (N_4945,N_4551,N_4591);
and U4946 (N_4946,N_4550,N_4624);
or U4947 (N_4947,N_4514,N_4734);
nor U4948 (N_4948,N_4706,N_4605);
and U4949 (N_4949,N_4580,N_4761);
nor U4950 (N_4950,N_4634,N_4517);
or U4951 (N_4951,N_4712,N_4710);
or U4952 (N_4952,N_4685,N_4770);
or U4953 (N_4953,N_4780,N_4606);
or U4954 (N_4954,N_4698,N_4681);
or U4955 (N_4955,N_4646,N_4762);
or U4956 (N_4956,N_4501,N_4516);
nor U4957 (N_4957,N_4510,N_4692);
or U4958 (N_4958,N_4577,N_4589);
and U4959 (N_4959,N_4563,N_4679);
nor U4960 (N_4960,N_4729,N_4789);
or U4961 (N_4961,N_4730,N_4712);
nor U4962 (N_4962,N_4598,N_4562);
xor U4963 (N_4963,N_4796,N_4632);
or U4964 (N_4964,N_4734,N_4725);
and U4965 (N_4965,N_4638,N_4720);
xnor U4966 (N_4966,N_4600,N_4700);
or U4967 (N_4967,N_4587,N_4577);
or U4968 (N_4968,N_4677,N_4689);
xor U4969 (N_4969,N_4663,N_4756);
and U4970 (N_4970,N_4702,N_4792);
nand U4971 (N_4971,N_4759,N_4506);
nand U4972 (N_4972,N_4773,N_4683);
nand U4973 (N_4973,N_4719,N_4687);
nor U4974 (N_4974,N_4699,N_4648);
xor U4975 (N_4975,N_4517,N_4740);
and U4976 (N_4976,N_4530,N_4605);
nand U4977 (N_4977,N_4687,N_4554);
or U4978 (N_4978,N_4504,N_4662);
nand U4979 (N_4979,N_4730,N_4523);
xnor U4980 (N_4980,N_4790,N_4765);
xnor U4981 (N_4981,N_4608,N_4535);
nand U4982 (N_4982,N_4657,N_4576);
and U4983 (N_4983,N_4712,N_4665);
nor U4984 (N_4984,N_4594,N_4774);
xor U4985 (N_4985,N_4587,N_4536);
xor U4986 (N_4986,N_4723,N_4594);
and U4987 (N_4987,N_4604,N_4547);
nand U4988 (N_4988,N_4587,N_4692);
nor U4989 (N_4989,N_4677,N_4724);
xor U4990 (N_4990,N_4658,N_4609);
nand U4991 (N_4991,N_4544,N_4778);
and U4992 (N_4992,N_4739,N_4777);
or U4993 (N_4993,N_4728,N_4502);
xor U4994 (N_4994,N_4711,N_4733);
nand U4995 (N_4995,N_4691,N_4700);
nand U4996 (N_4996,N_4748,N_4527);
or U4997 (N_4997,N_4516,N_4512);
and U4998 (N_4998,N_4748,N_4513);
and U4999 (N_4999,N_4614,N_4755);
xnor U5000 (N_5000,N_4764,N_4661);
and U5001 (N_5001,N_4572,N_4740);
and U5002 (N_5002,N_4595,N_4532);
nor U5003 (N_5003,N_4669,N_4723);
or U5004 (N_5004,N_4712,N_4791);
nor U5005 (N_5005,N_4526,N_4725);
xor U5006 (N_5006,N_4746,N_4512);
nor U5007 (N_5007,N_4511,N_4536);
xnor U5008 (N_5008,N_4743,N_4610);
nor U5009 (N_5009,N_4644,N_4619);
or U5010 (N_5010,N_4737,N_4562);
xor U5011 (N_5011,N_4727,N_4734);
xor U5012 (N_5012,N_4733,N_4677);
nor U5013 (N_5013,N_4747,N_4741);
xnor U5014 (N_5014,N_4517,N_4683);
nand U5015 (N_5015,N_4673,N_4600);
or U5016 (N_5016,N_4636,N_4631);
and U5017 (N_5017,N_4545,N_4754);
nor U5018 (N_5018,N_4629,N_4568);
and U5019 (N_5019,N_4729,N_4712);
xnor U5020 (N_5020,N_4583,N_4512);
and U5021 (N_5021,N_4707,N_4764);
or U5022 (N_5022,N_4735,N_4540);
xor U5023 (N_5023,N_4512,N_4730);
xnor U5024 (N_5024,N_4566,N_4748);
nand U5025 (N_5025,N_4690,N_4608);
nand U5026 (N_5026,N_4663,N_4537);
nand U5027 (N_5027,N_4504,N_4758);
and U5028 (N_5028,N_4697,N_4674);
xor U5029 (N_5029,N_4591,N_4554);
nand U5030 (N_5030,N_4681,N_4716);
nand U5031 (N_5031,N_4631,N_4508);
or U5032 (N_5032,N_4689,N_4746);
nand U5033 (N_5033,N_4778,N_4792);
xnor U5034 (N_5034,N_4648,N_4664);
xnor U5035 (N_5035,N_4648,N_4672);
or U5036 (N_5036,N_4553,N_4738);
nor U5037 (N_5037,N_4631,N_4741);
nand U5038 (N_5038,N_4794,N_4754);
nand U5039 (N_5039,N_4738,N_4533);
or U5040 (N_5040,N_4606,N_4557);
nor U5041 (N_5041,N_4582,N_4597);
and U5042 (N_5042,N_4675,N_4793);
nor U5043 (N_5043,N_4630,N_4626);
nand U5044 (N_5044,N_4512,N_4547);
xor U5045 (N_5045,N_4781,N_4572);
xnor U5046 (N_5046,N_4595,N_4770);
nor U5047 (N_5047,N_4668,N_4643);
xnor U5048 (N_5048,N_4536,N_4684);
nand U5049 (N_5049,N_4565,N_4603);
and U5050 (N_5050,N_4636,N_4725);
and U5051 (N_5051,N_4665,N_4669);
nor U5052 (N_5052,N_4575,N_4742);
xor U5053 (N_5053,N_4501,N_4571);
or U5054 (N_5054,N_4678,N_4676);
nor U5055 (N_5055,N_4617,N_4657);
xor U5056 (N_5056,N_4712,N_4699);
or U5057 (N_5057,N_4553,N_4504);
and U5058 (N_5058,N_4613,N_4598);
and U5059 (N_5059,N_4751,N_4690);
xnor U5060 (N_5060,N_4530,N_4769);
or U5061 (N_5061,N_4762,N_4743);
and U5062 (N_5062,N_4661,N_4581);
or U5063 (N_5063,N_4785,N_4761);
nand U5064 (N_5064,N_4751,N_4689);
or U5065 (N_5065,N_4663,N_4697);
and U5066 (N_5066,N_4536,N_4789);
and U5067 (N_5067,N_4758,N_4732);
nand U5068 (N_5068,N_4561,N_4558);
or U5069 (N_5069,N_4607,N_4504);
xnor U5070 (N_5070,N_4753,N_4648);
xor U5071 (N_5071,N_4758,N_4627);
nor U5072 (N_5072,N_4661,N_4508);
xnor U5073 (N_5073,N_4507,N_4729);
nand U5074 (N_5074,N_4692,N_4613);
and U5075 (N_5075,N_4732,N_4500);
or U5076 (N_5076,N_4792,N_4520);
or U5077 (N_5077,N_4633,N_4520);
and U5078 (N_5078,N_4512,N_4768);
or U5079 (N_5079,N_4669,N_4673);
nor U5080 (N_5080,N_4593,N_4717);
nor U5081 (N_5081,N_4589,N_4798);
or U5082 (N_5082,N_4791,N_4788);
or U5083 (N_5083,N_4572,N_4623);
nor U5084 (N_5084,N_4627,N_4522);
nand U5085 (N_5085,N_4504,N_4503);
and U5086 (N_5086,N_4590,N_4780);
nand U5087 (N_5087,N_4641,N_4796);
or U5088 (N_5088,N_4649,N_4643);
nand U5089 (N_5089,N_4608,N_4795);
nand U5090 (N_5090,N_4705,N_4791);
or U5091 (N_5091,N_4735,N_4568);
xor U5092 (N_5092,N_4599,N_4564);
and U5093 (N_5093,N_4524,N_4714);
nand U5094 (N_5094,N_4699,N_4736);
and U5095 (N_5095,N_4713,N_4553);
or U5096 (N_5096,N_4640,N_4591);
and U5097 (N_5097,N_4797,N_4786);
and U5098 (N_5098,N_4521,N_4668);
and U5099 (N_5099,N_4569,N_4634);
nand U5100 (N_5100,N_4991,N_5036);
xnor U5101 (N_5101,N_5028,N_4931);
xnor U5102 (N_5102,N_4927,N_5008);
nand U5103 (N_5103,N_4851,N_4836);
or U5104 (N_5104,N_4953,N_4810);
nor U5105 (N_5105,N_5067,N_4907);
and U5106 (N_5106,N_4998,N_4896);
xnor U5107 (N_5107,N_4848,N_4886);
nor U5108 (N_5108,N_5047,N_4857);
xor U5109 (N_5109,N_5022,N_4811);
and U5110 (N_5110,N_5053,N_4838);
nand U5111 (N_5111,N_4855,N_4928);
xor U5112 (N_5112,N_4849,N_4925);
nor U5113 (N_5113,N_4901,N_5045);
xor U5114 (N_5114,N_4913,N_4930);
or U5115 (N_5115,N_4958,N_4912);
nand U5116 (N_5116,N_5016,N_5049);
or U5117 (N_5117,N_4984,N_4936);
nor U5118 (N_5118,N_5011,N_4875);
xnor U5119 (N_5119,N_5078,N_4880);
xnor U5120 (N_5120,N_4996,N_4987);
xnor U5121 (N_5121,N_4847,N_4934);
nand U5122 (N_5122,N_4832,N_5069);
or U5123 (N_5123,N_5020,N_4842);
or U5124 (N_5124,N_5015,N_4844);
nor U5125 (N_5125,N_4878,N_4841);
nor U5126 (N_5126,N_5073,N_4899);
nand U5127 (N_5127,N_4920,N_4973);
xor U5128 (N_5128,N_4948,N_4893);
or U5129 (N_5129,N_4858,N_5039);
nor U5130 (N_5130,N_4982,N_4850);
and U5131 (N_5131,N_4960,N_4883);
and U5132 (N_5132,N_4826,N_4882);
or U5133 (N_5133,N_4820,N_5061);
xnor U5134 (N_5134,N_4877,N_4807);
or U5135 (N_5135,N_4992,N_4852);
or U5136 (N_5136,N_5072,N_4803);
or U5137 (N_5137,N_4827,N_5012);
or U5138 (N_5138,N_5000,N_4846);
and U5139 (N_5139,N_4995,N_4814);
nand U5140 (N_5140,N_4900,N_4809);
or U5141 (N_5141,N_4974,N_4916);
or U5142 (N_5142,N_5026,N_4823);
and U5143 (N_5143,N_4862,N_4994);
and U5144 (N_5144,N_4989,N_4961);
xnor U5145 (N_5145,N_5055,N_5052);
or U5146 (N_5146,N_4921,N_4970);
nand U5147 (N_5147,N_4924,N_5059);
nor U5148 (N_5148,N_4825,N_4819);
and U5149 (N_5149,N_4840,N_5058);
nand U5150 (N_5150,N_4954,N_4902);
nand U5151 (N_5151,N_5034,N_4828);
nand U5152 (N_5152,N_4949,N_4829);
or U5153 (N_5153,N_5032,N_5089);
nand U5154 (N_5154,N_4872,N_4969);
xnor U5155 (N_5155,N_5017,N_4894);
or U5156 (N_5156,N_4843,N_5082);
and U5157 (N_5157,N_4922,N_4835);
or U5158 (N_5158,N_4853,N_4837);
xor U5159 (N_5159,N_5035,N_5019);
or U5160 (N_5160,N_4885,N_4946);
or U5161 (N_5161,N_4932,N_4881);
or U5162 (N_5162,N_5009,N_4915);
xor U5163 (N_5163,N_4867,N_4863);
and U5164 (N_5164,N_4801,N_4892);
or U5165 (N_5165,N_5098,N_5064);
xnor U5166 (N_5166,N_5096,N_4923);
xor U5167 (N_5167,N_4866,N_5041);
nand U5168 (N_5168,N_5063,N_4950);
xnor U5169 (N_5169,N_5087,N_4971);
nand U5170 (N_5170,N_4955,N_4854);
xor U5171 (N_5171,N_4905,N_4968);
and U5172 (N_5172,N_4983,N_4830);
or U5173 (N_5173,N_4890,N_5095);
nand U5174 (N_5174,N_4981,N_4976);
and U5175 (N_5175,N_4914,N_5038);
nand U5176 (N_5176,N_4942,N_4933);
xor U5177 (N_5177,N_5025,N_5068);
xor U5178 (N_5178,N_5062,N_4945);
nand U5179 (N_5179,N_5006,N_5030);
or U5180 (N_5180,N_4940,N_5080);
nor U5181 (N_5181,N_5079,N_4967);
or U5182 (N_5182,N_4839,N_4845);
xor U5183 (N_5183,N_5001,N_5014);
nand U5184 (N_5184,N_5024,N_4941);
nand U5185 (N_5185,N_4963,N_4943);
or U5186 (N_5186,N_4884,N_4904);
nand U5187 (N_5187,N_4833,N_4910);
nor U5188 (N_5188,N_4879,N_4808);
and U5189 (N_5189,N_4966,N_4985);
nand U5190 (N_5190,N_4805,N_5027);
or U5191 (N_5191,N_5076,N_4908);
and U5192 (N_5192,N_4871,N_4802);
nand U5193 (N_5193,N_5084,N_5040);
xnor U5194 (N_5194,N_4997,N_5097);
xor U5195 (N_5195,N_5046,N_5057);
and U5196 (N_5196,N_5013,N_5050);
nor U5197 (N_5197,N_4993,N_4903);
nand U5198 (N_5198,N_4817,N_4999);
nor U5199 (N_5199,N_5004,N_5048);
xor U5200 (N_5200,N_4891,N_4815);
nand U5201 (N_5201,N_5093,N_5033);
or U5202 (N_5202,N_4865,N_5077);
xor U5203 (N_5203,N_5018,N_5054);
nor U5204 (N_5204,N_5042,N_5081);
nand U5205 (N_5205,N_5051,N_5031);
nor U5206 (N_5206,N_4917,N_4868);
nor U5207 (N_5207,N_4957,N_4959);
or U5208 (N_5208,N_4897,N_4918);
nor U5209 (N_5209,N_4834,N_4962);
or U5210 (N_5210,N_4861,N_4972);
and U5211 (N_5211,N_4888,N_4864);
nand U5212 (N_5212,N_5066,N_4937);
and U5213 (N_5213,N_4818,N_4859);
nand U5214 (N_5214,N_5003,N_4978);
or U5215 (N_5215,N_5007,N_5083);
or U5216 (N_5216,N_5043,N_4944);
xor U5217 (N_5217,N_4952,N_4804);
nand U5218 (N_5218,N_4870,N_4980);
nand U5219 (N_5219,N_5023,N_4956);
and U5220 (N_5220,N_4929,N_4986);
and U5221 (N_5221,N_4869,N_4876);
nor U5222 (N_5222,N_4824,N_4889);
xor U5223 (N_5223,N_4975,N_5010);
and U5224 (N_5224,N_5005,N_4813);
xor U5225 (N_5225,N_4856,N_4965);
nand U5226 (N_5226,N_4898,N_4926);
xnor U5227 (N_5227,N_5094,N_4806);
nor U5228 (N_5228,N_4895,N_5021);
nand U5229 (N_5229,N_4964,N_4822);
nor U5230 (N_5230,N_5029,N_4919);
or U5231 (N_5231,N_4939,N_5099);
or U5232 (N_5232,N_5060,N_4821);
or U5233 (N_5233,N_4873,N_5071);
xnor U5234 (N_5234,N_4906,N_5074);
xnor U5235 (N_5235,N_5075,N_5065);
or U5236 (N_5236,N_4812,N_5088);
nor U5237 (N_5237,N_4988,N_4909);
and U5238 (N_5238,N_5085,N_4947);
xnor U5239 (N_5239,N_4938,N_4935);
nand U5240 (N_5240,N_5056,N_5002);
or U5241 (N_5241,N_4887,N_4800);
nand U5242 (N_5242,N_4831,N_4816);
nor U5243 (N_5243,N_5091,N_4979);
xnor U5244 (N_5244,N_4874,N_5070);
and U5245 (N_5245,N_5090,N_5086);
nor U5246 (N_5246,N_5037,N_4990);
nand U5247 (N_5247,N_5044,N_4911);
xnor U5248 (N_5248,N_4977,N_4951);
nor U5249 (N_5249,N_5092,N_4860);
nand U5250 (N_5250,N_4898,N_5010);
nand U5251 (N_5251,N_5045,N_4909);
or U5252 (N_5252,N_5060,N_4946);
nand U5253 (N_5253,N_4892,N_5010);
xor U5254 (N_5254,N_4837,N_4885);
or U5255 (N_5255,N_4932,N_4892);
xnor U5256 (N_5256,N_4997,N_4971);
nand U5257 (N_5257,N_4841,N_4964);
xor U5258 (N_5258,N_4800,N_4996);
xnor U5259 (N_5259,N_5072,N_4947);
and U5260 (N_5260,N_5084,N_5082);
nor U5261 (N_5261,N_4990,N_5000);
and U5262 (N_5262,N_5049,N_4949);
or U5263 (N_5263,N_4918,N_5028);
xnor U5264 (N_5264,N_5009,N_4925);
nor U5265 (N_5265,N_4831,N_4821);
or U5266 (N_5266,N_4953,N_5093);
nor U5267 (N_5267,N_4815,N_4863);
xor U5268 (N_5268,N_4840,N_4948);
xnor U5269 (N_5269,N_4860,N_4995);
nand U5270 (N_5270,N_4925,N_4928);
nand U5271 (N_5271,N_4817,N_5031);
xnor U5272 (N_5272,N_4955,N_4920);
xor U5273 (N_5273,N_4969,N_5077);
xnor U5274 (N_5274,N_4866,N_5098);
nand U5275 (N_5275,N_5078,N_5099);
and U5276 (N_5276,N_4994,N_4886);
and U5277 (N_5277,N_5000,N_4843);
and U5278 (N_5278,N_5077,N_5003);
nand U5279 (N_5279,N_5089,N_4997);
and U5280 (N_5280,N_4900,N_4921);
and U5281 (N_5281,N_4939,N_4913);
xor U5282 (N_5282,N_4860,N_4959);
xor U5283 (N_5283,N_5041,N_5033);
or U5284 (N_5284,N_4983,N_4921);
or U5285 (N_5285,N_4870,N_4985);
and U5286 (N_5286,N_5073,N_4971);
and U5287 (N_5287,N_5014,N_4852);
xnor U5288 (N_5288,N_4859,N_4943);
xor U5289 (N_5289,N_4884,N_4871);
or U5290 (N_5290,N_4957,N_4981);
or U5291 (N_5291,N_5023,N_4934);
and U5292 (N_5292,N_4909,N_4997);
or U5293 (N_5293,N_5066,N_4952);
nor U5294 (N_5294,N_4917,N_5032);
and U5295 (N_5295,N_5066,N_4848);
xnor U5296 (N_5296,N_4825,N_4965);
nor U5297 (N_5297,N_4929,N_5063);
and U5298 (N_5298,N_5002,N_4874);
xor U5299 (N_5299,N_5059,N_4822);
or U5300 (N_5300,N_4944,N_4874);
xor U5301 (N_5301,N_5034,N_4884);
xnor U5302 (N_5302,N_4843,N_5079);
and U5303 (N_5303,N_4976,N_4868);
or U5304 (N_5304,N_5036,N_5083);
nand U5305 (N_5305,N_5084,N_5019);
xor U5306 (N_5306,N_4803,N_4877);
nand U5307 (N_5307,N_4878,N_4903);
xor U5308 (N_5308,N_4960,N_4944);
or U5309 (N_5309,N_4910,N_5073);
or U5310 (N_5310,N_5026,N_5087);
nor U5311 (N_5311,N_5053,N_4956);
nand U5312 (N_5312,N_5073,N_5066);
and U5313 (N_5313,N_4859,N_4995);
and U5314 (N_5314,N_4871,N_5088);
nor U5315 (N_5315,N_4994,N_5030);
and U5316 (N_5316,N_4821,N_5087);
xor U5317 (N_5317,N_4806,N_5058);
nand U5318 (N_5318,N_5059,N_5039);
or U5319 (N_5319,N_4990,N_4977);
or U5320 (N_5320,N_5018,N_4932);
or U5321 (N_5321,N_4934,N_5003);
and U5322 (N_5322,N_4830,N_4891);
or U5323 (N_5323,N_4830,N_4883);
nor U5324 (N_5324,N_4907,N_4854);
or U5325 (N_5325,N_5039,N_5092);
xor U5326 (N_5326,N_4869,N_4883);
nor U5327 (N_5327,N_5001,N_4873);
nor U5328 (N_5328,N_4996,N_4871);
xor U5329 (N_5329,N_5009,N_4840);
and U5330 (N_5330,N_4996,N_4972);
and U5331 (N_5331,N_5088,N_4972);
and U5332 (N_5332,N_4945,N_4891);
xnor U5333 (N_5333,N_5085,N_4846);
or U5334 (N_5334,N_5065,N_4872);
nand U5335 (N_5335,N_4956,N_5040);
nor U5336 (N_5336,N_4806,N_5049);
nor U5337 (N_5337,N_4833,N_4983);
nand U5338 (N_5338,N_5004,N_5028);
nor U5339 (N_5339,N_4925,N_4834);
nor U5340 (N_5340,N_4926,N_5038);
or U5341 (N_5341,N_5019,N_5033);
and U5342 (N_5342,N_4882,N_5070);
xor U5343 (N_5343,N_5039,N_4993);
xnor U5344 (N_5344,N_4848,N_4944);
and U5345 (N_5345,N_4913,N_4931);
and U5346 (N_5346,N_4869,N_4894);
xor U5347 (N_5347,N_5011,N_4918);
nor U5348 (N_5348,N_4947,N_4914);
or U5349 (N_5349,N_4822,N_5036);
nor U5350 (N_5350,N_4870,N_4885);
and U5351 (N_5351,N_5060,N_5072);
xor U5352 (N_5352,N_4885,N_4876);
and U5353 (N_5353,N_4832,N_4818);
and U5354 (N_5354,N_5003,N_4986);
xor U5355 (N_5355,N_4960,N_5005);
nand U5356 (N_5356,N_4961,N_4922);
xor U5357 (N_5357,N_4922,N_5039);
and U5358 (N_5358,N_4853,N_4868);
and U5359 (N_5359,N_4886,N_5011);
nor U5360 (N_5360,N_4954,N_5099);
or U5361 (N_5361,N_5058,N_4958);
nand U5362 (N_5362,N_5076,N_5020);
nand U5363 (N_5363,N_4823,N_4867);
or U5364 (N_5364,N_5077,N_4953);
nand U5365 (N_5365,N_5056,N_4806);
xnor U5366 (N_5366,N_4904,N_4829);
and U5367 (N_5367,N_4973,N_4977);
xor U5368 (N_5368,N_4825,N_4845);
nand U5369 (N_5369,N_5054,N_5093);
and U5370 (N_5370,N_5043,N_5074);
or U5371 (N_5371,N_5014,N_5053);
nor U5372 (N_5372,N_4999,N_4910);
or U5373 (N_5373,N_5066,N_4883);
nand U5374 (N_5374,N_4897,N_4937);
or U5375 (N_5375,N_4854,N_5076);
nand U5376 (N_5376,N_4887,N_4995);
xor U5377 (N_5377,N_4867,N_5086);
nor U5378 (N_5378,N_4818,N_4893);
or U5379 (N_5379,N_5014,N_5082);
xor U5380 (N_5380,N_4950,N_5001);
nor U5381 (N_5381,N_4978,N_4975);
nand U5382 (N_5382,N_4834,N_4878);
nor U5383 (N_5383,N_4918,N_4922);
nand U5384 (N_5384,N_4852,N_4849);
xnor U5385 (N_5385,N_4825,N_4836);
or U5386 (N_5386,N_5018,N_4854);
nor U5387 (N_5387,N_5091,N_4912);
and U5388 (N_5388,N_5074,N_4997);
nand U5389 (N_5389,N_4817,N_4906);
nand U5390 (N_5390,N_4926,N_4967);
and U5391 (N_5391,N_4999,N_4812);
or U5392 (N_5392,N_4982,N_5066);
nor U5393 (N_5393,N_4971,N_5085);
nor U5394 (N_5394,N_5069,N_5030);
nor U5395 (N_5395,N_4856,N_4871);
xor U5396 (N_5396,N_4933,N_5046);
xnor U5397 (N_5397,N_4996,N_4928);
nand U5398 (N_5398,N_5034,N_4912);
xnor U5399 (N_5399,N_4993,N_4875);
and U5400 (N_5400,N_5253,N_5178);
nand U5401 (N_5401,N_5376,N_5364);
xnor U5402 (N_5402,N_5220,N_5327);
or U5403 (N_5403,N_5216,N_5369);
nand U5404 (N_5404,N_5222,N_5256);
and U5405 (N_5405,N_5168,N_5221);
nor U5406 (N_5406,N_5329,N_5223);
and U5407 (N_5407,N_5372,N_5338);
or U5408 (N_5408,N_5363,N_5203);
nand U5409 (N_5409,N_5377,N_5177);
and U5410 (N_5410,N_5116,N_5310);
or U5411 (N_5411,N_5301,N_5226);
xor U5412 (N_5412,N_5340,N_5288);
nand U5413 (N_5413,N_5323,N_5276);
or U5414 (N_5414,N_5279,N_5334);
nand U5415 (N_5415,N_5384,N_5371);
or U5416 (N_5416,N_5175,N_5126);
nor U5417 (N_5417,N_5354,N_5394);
nand U5418 (N_5418,N_5294,N_5196);
or U5419 (N_5419,N_5395,N_5343);
nor U5420 (N_5420,N_5254,N_5118);
or U5421 (N_5421,N_5280,N_5393);
xor U5422 (N_5422,N_5251,N_5399);
or U5423 (N_5423,N_5190,N_5213);
or U5424 (N_5424,N_5103,N_5242);
nor U5425 (N_5425,N_5383,N_5200);
and U5426 (N_5426,N_5305,N_5275);
nand U5427 (N_5427,N_5137,N_5373);
or U5428 (N_5428,N_5125,N_5344);
nand U5429 (N_5429,N_5161,N_5247);
or U5430 (N_5430,N_5237,N_5355);
or U5431 (N_5431,N_5236,N_5139);
xor U5432 (N_5432,N_5181,N_5229);
nand U5433 (N_5433,N_5140,N_5321);
nand U5434 (N_5434,N_5111,N_5123);
nor U5435 (N_5435,N_5353,N_5157);
nand U5436 (N_5436,N_5268,N_5345);
or U5437 (N_5437,N_5101,N_5105);
xnor U5438 (N_5438,N_5154,N_5266);
nand U5439 (N_5439,N_5217,N_5366);
and U5440 (N_5440,N_5389,N_5204);
nand U5441 (N_5441,N_5258,N_5114);
nand U5442 (N_5442,N_5215,N_5102);
and U5443 (N_5443,N_5314,N_5100);
or U5444 (N_5444,N_5360,N_5341);
and U5445 (N_5445,N_5194,N_5121);
and U5446 (N_5446,N_5162,N_5262);
nor U5447 (N_5447,N_5248,N_5244);
or U5448 (N_5448,N_5332,N_5156);
nor U5449 (N_5449,N_5241,N_5183);
or U5450 (N_5450,N_5107,N_5296);
nand U5451 (N_5451,N_5284,N_5198);
xnor U5452 (N_5452,N_5291,N_5325);
xnor U5453 (N_5453,N_5135,N_5238);
or U5454 (N_5454,N_5397,N_5170);
xor U5455 (N_5455,N_5233,N_5386);
or U5456 (N_5456,N_5270,N_5337);
or U5457 (N_5457,N_5388,N_5269);
nor U5458 (N_5458,N_5113,N_5283);
and U5459 (N_5459,N_5250,N_5300);
or U5460 (N_5460,N_5231,N_5335);
and U5461 (N_5461,N_5333,N_5147);
nand U5462 (N_5462,N_5187,N_5272);
and U5463 (N_5463,N_5246,N_5180);
xor U5464 (N_5464,N_5320,N_5218);
and U5465 (N_5465,N_5273,N_5207);
nor U5466 (N_5466,N_5163,N_5176);
nor U5467 (N_5467,N_5295,N_5146);
xnor U5468 (N_5468,N_5368,N_5185);
xor U5469 (N_5469,N_5212,N_5342);
nor U5470 (N_5470,N_5287,N_5141);
nand U5471 (N_5471,N_5227,N_5142);
or U5472 (N_5472,N_5317,N_5186);
xnor U5473 (N_5473,N_5165,N_5130);
or U5474 (N_5474,N_5285,N_5326);
xor U5475 (N_5475,N_5235,N_5390);
xnor U5476 (N_5476,N_5106,N_5138);
and U5477 (N_5477,N_5382,N_5169);
nand U5478 (N_5478,N_5239,N_5136);
nand U5479 (N_5479,N_5145,N_5311);
nand U5480 (N_5480,N_5357,N_5159);
and U5481 (N_5481,N_5265,N_5359);
xnor U5482 (N_5482,N_5166,N_5252);
nor U5483 (N_5483,N_5188,N_5132);
nor U5484 (N_5484,N_5290,N_5303);
nor U5485 (N_5485,N_5119,N_5153);
xor U5486 (N_5486,N_5375,N_5219);
nor U5487 (N_5487,N_5104,N_5362);
nor U5488 (N_5488,N_5324,N_5133);
or U5489 (N_5489,N_5128,N_5199);
nor U5490 (N_5490,N_5308,N_5232);
or U5491 (N_5491,N_5349,N_5352);
xnor U5492 (N_5492,N_5189,N_5228);
or U5493 (N_5493,N_5224,N_5124);
nor U5494 (N_5494,N_5307,N_5292);
xnor U5495 (N_5495,N_5182,N_5361);
and U5496 (N_5496,N_5172,N_5134);
xnor U5497 (N_5497,N_5129,N_5289);
or U5498 (N_5498,N_5346,N_5108);
xnor U5499 (N_5499,N_5110,N_5211);
and U5500 (N_5500,N_5259,N_5282);
xor U5501 (N_5501,N_5356,N_5277);
and U5502 (N_5502,N_5380,N_5312);
and U5503 (N_5503,N_5274,N_5319);
nor U5504 (N_5504,N_5122,N_5309);
and U5505 (N_5505,N_5115,N_5365);
nand U5506 (N_5506,N_5158,N_5316);
and U5507 (N_5507,N_5179,N_5243);
or U5508 (N_5508,N_5120,N_5267);
or U5509 (N_5509,N_5379,N_5358);
or U5510 (N_5510,N_5249,N_5195);
xor U5511 (N_5511,N_5164,N_5143);
and U5512 (N_5512,N_5230,N_5117);
or U5513 (N_5513,N_5260,N_5328);
nand U5514 (N_5514,N_5378,N_5151);
nor U5515 (N_5515,N_5192,N_5144);
nand U5516 (N_5516,N_5315,N_5191);
nor U5517 (N_5517,N_5304,N_5263);
nand U5518 (N_5518,N_5293,N_5240);
nor U5519 (N_5519,N_5264,N_5148);
nand U5520 (N_5520,N_5160,N_5298);
nand U5521 (N_5521,N_5234,N_5214);
or U5522 (N_5522,N_5348,N_5174);
or U5523 (N_5523,N_5313,N_5297);
nor U5524 (N_5524,N_5322,N_5347);
nor U5525 (N_5525,N_5306,N_5350);
nor U5526 (N_5526,N_5131,N_5109);
or U5527 (N_5527,N_5385,N_5167);
nor U5528 (N_5528,N_5184,N_5209);
nor U5529 (N_5529,N_5398,N_5396);
nor U5530 (N_5530,N_5374,N_5206);
nor U5531 (N_5531,N_5173,N_5261);
nor U5532 (N_5532,N_5197,N_5152);
or U5533 (N_5533,N_5281,N_5202);
or U5534 (N_5534,N_5381,N_5370);
and U5535 (N_5535,N_5112,N_5331);
nand U5536 (N_5536,N_5387,N_5392);
nor U5537 (N_5537,N_5255,N_5245);
xor U5538 (N_5538,N_5127,N_5367);
or U5539 (N_5539,N_5171,N_5193);
and U5540 (N_5540,N_5330,N_5210);
and U5541 (N_5541,N_5225,N_5150);
and U5542 (N_5542,N_5318,N_5302);
nor U5543 (N_5543,N_5149,N_5351);
nor U5544 (N_5544,N_5286,N_5336);
nand U5545 (N_5545,N_5201,N_5271);
and U5546 (N_5546,N_5339,N_5391);
nand U5547 (N_5547,N_5208,N_5205);
xor U5548 (N_5548,N_5155,N_5299);
nand U5549 (N_5549,N_5257,N_5278);
and U5550 (N_5550,N_5198,N_5300);
nand U5551 (N_5551,N_5178,N_5154);
nor U5552 (N_5552,N_5207,N_5180);
nand U5553 (N_5553,N_5133,N_5344);
nand U5554 (N_5554,N_5377,N_5236);
and U5555 (N_5555,N_5226,N_5278);
and U5556 (N_5556,N_5197,N_5136);
and U5557 (N_5557,N_5110,N_5335);
xnor U5558 (N_5558,N_5377,N_5397);
or U5559 (N_5559,N_5161,N_5285);
nand U5560 (N_5560,N_5191,N_5266);
nand U5561 (N_5561,N_5333,N_5338);
nor U5562 (N_5562,N_5310,N_5301);
nor U5563 (N_5563,N_5156,N_5381);
xor U5564 (N_5564,N_5343,N_5209);
nand U5565 (N_5565,N_5380,N_5351);
xor U5566 (N_5566,N_5392,N_5138);
xnor U5567 (N_5567,N_5178,N_5168);
nor U5568 (N_5568,N_5395,N_5292);
and U5569 (N_5569,N_5193,N_5298);
and U5570 (N_5570,N_5277,N_5307);
or U5571 (N_5571,N_5369,N_5147);
or U5572 (N_5572,N_5359,N_5124);
or U5573 (N_5573,N_5325,N_5169);
nand U5574 (N_5574,N_5161,N_5336);
xnor U5575 (N_5575,N_5117,N_5165);
or U5576 (N_5576,N_5205,N_5118);
xnor U5577 (N_5577,N_5207,N_5111);
nor U5578 (N_5578,N_5133,N_5309);
xnor U5579 (N_5579,N_5151,N_5184);
nor U5580 (N_5580,N_5340,N_5275);
or U5581 (N_5581,N_5393,N_5171);
and U5582 (N_5582,N_5361,N_5115);
nand U5583 (N_5583,N_5341,N_5117);
or U5584 (N_5584,N_5162,N_5394);
nand U5585 (N_5585,N_5370,N_5126);
nor U5586 (N_5586,N_5160,N_5370);
nand U5587 (N_5587,N_5291,N_5338);
xor U5588 (N_5588,N_5392,N_5179);
nand U5589 (N_5589,N_5218,N_5361);
xor U5590 (N_5590,N_5368,N_5394);
nand U5591 (N_5591,N_5134,N_5372);
nand U5592 (N_5592,N_5149,N_5243);
or U5593 (N_5593,N_5259,N_5296);
nand U5594 (N_5594,N_5120,N_5377);
nor U5595 (N_5595,N_5392,N_5391);
nor U5596 (N_5596,N_5355,N_5190);
nand U5597 (N_5597,N_5255,N_5249);
and U5598 (N_5598,N_5346,N_5246);
or U5599 (N_5599,N_5304,N_5170);
xor U5600 (N_5600,N_5271,N_5204);
nand U5601 (N_5601,N_5282,N_5377);
nand U5602 (N_5602,N_5246,N_5308);
nand U5603 (N_5603,N_5288,N_5214);
nand U5604 (N_5604,N_5211,N_5241);
nand U5605 (N_5605,N_5334,N_5380);
nand U5606 (N_5606,N_5187,N_5343);
and U5607 (N_5607,N_5274,N_5101);
or U5608 (N_5608,N_5304,N_5254);
nor U5609 (N_5609,N_5350,N_5223);
nor U5610 (N_5610,N_5261,N_5179);
nor U5611 (N_5611,N_5337,N_5168);
or U5612 (N_5612,N_5175,N_5331);
or U5613 (N_5613,N_5312,N_5130);
nand U5614 (N_5614,N_5321,N_5273);
nor U5615 (N_5615,N_5244,N_5105);
nor U5616 (N_5616,N_5313,N_5227);
xor U5617 (N_5617,N_5243,N_5379);
xor U5618 (N_5618,N_5363,N_5327);
and U5619 (N_5619,N_5209,N_5179);
xor U5620 (N_5620,N_5365,N_5156);
and U5621 (N_5621,N_5299,N_5337);
or U5622 (N_5622,N_5250,N_5361);
and U5623 (N_5623,N_5296,N_5176);
nor U5624 (N_5624,N_5165,N_5190);
and U5625 (N_5625,N_5380,N_5202);
or U5626 (N_5626,N_5209,N_5114);
nor U5627 (N_5627,N_5243,N_5141);
nand U5628 (N_5628,N_5130,N_5290);
or U5629 (N_5629,N_5350,N_5126);
or U5630 (N_5630,N_5126,N_5335);
xnor U5631 (N_5631,N_5251,N_5289);
and U5632 (N_5632,N_5129,N_5397);
and U5633 (N_5633,N_5225,N_5350);
nor U5634 (N_5634,N_5257,N_5172);
and U5635 (N_5635,N_5293,N_5200);
and U5636 (N_5636,N_5160,N_5354);
xor U5637 (N_5637,N_5359,N_5116);
nand U5638 (N_5638,N_5374,N_5125);
xor U5639 (N_5639,N_5284,N_5331);
nand U5640 (N_5640,N_5359,N_5228);
and U5641 (N_5641,N_5323,N_5269);
and U5642 (N_5642,N_5399,N_5388);
or U5643 (N_5643,N_5324,N_5161);
and U5644 (N_5644,N_5150,N_5248);
nand U5645 (N_5645,N_5176,N_5177);
or U5646 (N_5646,N_5365,N_5222);
or U5647 (N_5647,N_5341,N_5148);
nor U5648 (N_5648,N_5187,N_5118);
or U5649 (N_5649,N_5232,N_5322);
and U5650 (N_5650,N_5272,N_5289);
and U5651 (N_5651,N_5205,N_5138);
nor U5652 (N_5652,N_5324,N_5253);
nor U5653 (N_5653,N_5345,N_5386);
xor U5654 (N_5654,N_5142,N_5102);
xor U5655 (N_5655,N_5138,N_5262);
nor U5656 (N_5656,N_5240,N_5129);
nor U5657 (N_5657,N_5224,N_5219);
xor U5658 (N_5658,N_5327,N_5272);
and U5659 (N_5659,N_5143,N_5377);
and U5660 (N_5660,N_5175,N_5317);
or U5661 (N_5661,N_5385,N_5232);
and U5662 (N_5662,N_5270,N_5142);
or U5663 (N_5663,N_5155,N_5190);
xor U5664 (N_5664,N_5210,N_5339);
nand U5665 (N_5665,N_5369,N_5121);
nand U5666 (N_5666,N_5222,N_5387);
and U5667 (N_5667,N_5265,N_5328);
and U5668 (N_5668,N_5343,N_5392);
nor U5669 (N_5669,N_5267,N_5308);
or U5670 (N_5670,N_5309,N_5193);
xnor U5671 (N_5671,N_5263,N_5138);
nor U5672 (N_5672,N_5253,N_5355);
or U5673 (N_5673,N_5167,N_5277);
or U5674 (N_5674,N_5343,N_5348);
nor U5675 (N_5675,N_5361,N_5255);
nor U5676 (N_5676,N_5388,N_5126);
nand U5677 (N_5677,N_5276,N_5328);
or U5678 (N_5678,N_5271,N_5292);
nor U5679 (N_5679,N_5133,N_5383);
or U5680 (N_5680,N_5120,N_5313);
or U5681 (N_5681,N_5273,N_5210);
nor U5682 (N_5682,N_5127,N_5259);
and U5683 (N_5683,N_5251,N_5331);
nor U5684 (N_5684,N_5268,N_5322);
nor U5685 (N_5685,N_5274,N_5280);
or U5686 (N_5686,N_5183,N_5145);
nor U5687 (N_5687,N_5265,N_5333);
or U5688 (N_5688,N_5299,N_5123);
xor U5689 (N_5689,N_5115,N_5189);
or U5690 (N_5690,N_5150,N_5258);
nand U5691 (N_5691,N_5284,N_5179);
nor U5692 (N_5692,N_5387,N_5276);
nand U5693 (N_5693,N_5212,N_5339);
xnor U5694 (N_5694,N_5367,N_5380);
nand U5695 (N_5695,N_5255,N_5194);
and U5696 (N_5696,N_5216,N_5124);
nand U5697 (N_5697,N_5352,N_5173);
xnor U5698 (N_5698,N_5260,N_5194);
nand U5699 (N_5699,N_5248,N_5165);
xor U5700 (N_5700,N_5613,N_5437);
xnor U5701 (N_5701,N_5548,N_5580);
and U5702 (N_5702,N_5603,N_5678);
or U5703 (N_5703,N_5474,N_5670);
nor U5704 (N_5704,N_5672,N_5524);
or U5705 (N_5705,N_5662,N_5405);
or U5706 (N_5706,N_5594,N_5552);
nand U5707 (N_5707,N_5676,N_5617);
xnor U5708 (N_5708,N_5683,N_5442);
and U5709 (N_5709,N_5458,N_5528);
nand U5710 (N_5710,N_5616,N_5413);
and U5711 (N_5711,N_5596,N_5504);
and U5712 (N_5712,N_5465,N_5411);
xor U5713 (N_5713,N_5673,N_5569);
xor U5714 (N_5714,N_5625,N_5565);
nand U5715 (N_5715,N_5557,N_5534);
xnor U5716 (N_5716,N_5460,N_5637);
or U5717 (N_5717,N_5539,N_5591);
and U5718 (N_5718,N_5681,N_5404);
xnor U5719 (N_5719,N_5449,N_5443);
nor U5720 (N_5720,N_5567,N_5698);
nor U5721 (N_5721,N_5452,N_5506);
nand U5722 (N_5722,N_5497,N_5614);
xor U5723 (N_5723,N_5450,N_5650);
xor U5724 (N_5724,N_5619,N_5559);
xor U5725 (N_5725,N_5517,N_5666);
nand U5726 (N_5726,N_5599,N_5615);
and U5727 (N_5727,N_5521,N_5464);
nor U5728 (N_5728,N_5551,N_5526);
xor U5729 (N_5729,N_5634,N_5501);
or U5730 (N_5730,N_5412,N_5478);
xor U5731 (N_5731,N_5447,N_5572);
xnor U5732 (N_5732,N_5498,N_5518);
xnor U5733 (N_5733,N_5657,N_5571);
xor U5734 (N_5734,N_5632,N_5694);
xnor U5735 (N_5735,N_5495,N_5429);
or U5736 (N_5736,N_5612,N_5527);
nor U5737 (N_5737,N_5476,N_5422);
nand U5738 (N_5738,N_5689,N_5640);
and U5739 (N_5739,N_5410,N_5561);
or U5740 (N_5740,N_5570,N_5626);
xnor U5741 (N_5741,N_5491,N_5618);
and U5742 (N_5742,N_5542,N_5586);
nand U5743 (N_5743,N_5510,N_5461);
and U5744 (N_5744,N_5659,N_5477);
nor U5745 (N_5745,N_5522,N_5469);
nand U5746 (N_5746,N_5558,N_5597);
xnor U5747 (N_5747,N_5585,N_5573);
nor U5748 (N_5748,N_5529,N_5457);
nand U5749 (N_5749,N_5503,N_5674);
nor U5750 (N_5750,N_5691,N_5502);
and U5751 (N_5751,N_5505,N_5562);
and U5752 (N_5752,N_5687,N_5540);
nor U5753 (N_5753,N_5608,N_5611);
and U5754 (N_5754,N_5680,N_5642);
and U5755 (N_5755,N_5686,N_5403);
nor U5756 (N_5756,N_5487,N_5440);
or U5757 (N_5757,N_5622,N_5516);
and U5758 (N_5758,N_5675,N_5610);
and U5759 (N_5759,N_5671,N_5514);
nor U5760 (N_5760,N_5463,N_5554);
or U5761 (N_5761,N_5550,N_5545);
nand U5762 (N_5762,N_5607,N_5584);
nand U5763 (N_5763,N_5576,N_5446);
nand U5764 (N_5764,N_5531,N_5624);
and U5765 (N_5765,N_5647,N_5466);
and U5766 (N_5766,N_5547,N_5525);
or U5767 (N_5767,N_5602,N_5685);
nand U5768 (N_5768,N_5424,N_5668);
and U5769 (N_5769,N_5620,N_5544);
nor U5770 (N_5770,N_5648,N_5445);
xnor U5771 (N_5771,N_5682,N_5451);
nand U5772 (N_5772,N_5605,N_5414);
and U5773 (N_5773,N_5459,N_5423);
nor U5774 (N_5774,N_5665,N_5621);
and U5775 (N_5775,N_5435,N_5669);
or U5776 (N_5776,N_5566,N_5630);
xor U5777 (N_5777,N_5490,N_5646);
and U5778 (N_5778,N_5604,N_5515);
or U5779 (N_5779,N_5651,N_5638);
nand U5780 (N_5780,N_5500,N_5577);
and U5781 (N_5781,N_5588,N_5664);
or U5782 (N_5782,N_5568,N_5587);
nor U5783 (N_5783,N_5472,N_5533);
or U5784 (N_5784,N_5623,N_5695);
nand U5785 (N_5785,N_5541,N_5483);
xor U5786 (N_5786,N_5482,N_5537);
and U5787 (N_5787,N_5627,N_5633);
nor U5788 (N_5788,N_5601,N_5473);
or U5789 (N_5789,N_5661,N_5420);
nor U5790 (N_5790,N_5660,N_5656);
or U5791 (N_5791,N_5643,N_5628);
xnor U5792 (N_5792,N_5635,N_5467);
nor U5793 (N_5793,N_5581,N_5532);
and U5794 (N_5794,N_5654,N_5431);
and U5795 (N_5795,N_5430,N_5639);
xor U5796 (N_5796,N_5593,N_5513);
xnor U5797 (N_5797,N_5693,N_5644);
or U5798 (N_5798,N_5579,N_5439);
and U5799 (N_5799,N_5667,N_5493);
or U5800 (N_5800,N_5699,N_5454);
nand U5801 (N_5801,N_5402,N_5408);
xnor U5802 (N_5802,N_5511,N_5481);
xor U5803 (N_5803,N_5575,N_5592);
and U5804 (N_5804,N_5494,N_5684);
xor U5805 (N_5805,N_5468,N_5574);
xnor U5806 (N_5806,N_5416,N_5471);
and U5807 (N_5807,N_5560,N_5598);
nor U5808 (N_5808,N_5595,N_5535);
nand U5809 (N_5809,N_5629,N_5441);
xnor U5810 (N_5810,N_5649,N_5427);
nand U5811 (N_5811,N_5470,N_5489);
and U5812 (N_5812,N_5523,N_5499);
nand U5813 (N_5813,N_5663,N_5507);
or U5814 (N_5814,N_5563,N_5688);
and U5815 (N_5815,N_5578,N_5406);
xor U5816 (N_5816,N_5509,N_5600);
and U5817 (N_5817,N_5426,N_5486);
or U5818 (N_5818,N_5492,N_5436);
and U5819 (N_5819,N_5453,N_5641);
nor U5820 (N_5820,N_5425,N_5484);
nand U5821 (N_5821,N_5401,N_5583);
or U5822 (N_5822,N_5589,N_5655);
and U5823 (N_5823,N_5555,N_5432);
nor U5824 (N_5824,N_5485,N_5433);
or U5825 (N_5825,N_5543,N_5590);
and U5826 (N_5826,N_5409,N_5609);
nor U5827 (N_5827,N_5679,N_5538);
nand U5828 (N_5828,N_5496,N_5582);
or U5829 (N_5829,N_5419,N_5415);
xor U5830 (N_5830,N_5631,N_5488);
or U5831 (N_5831,N_5549,N_5438);
xnor U5832 (N_5832,N_5696,N_5636);
nor U5833 (N_5833,N_5677,N_5645);
or U5834 (N_5834,N_5456,N_5462);
nand U5835 (N_5835,N_5428,N_5400);
nand U5836 (N_5836,N_5697,N_5692);
nor U5837 (N_5837,N_5407,N_5556);
or U5838 (N_5838,N_5480,N_5444);
or U5839 (N_5839,N_5512,N_5448);
nor U5840 (N_5840,N_5519,N_5652);
and U5841 (N_5841,N_5564,N_5508);
and U5842 (N_5842,N_5418,N_5417);
nor U5843 (N_5843,N_5530,N_5434);
xnor U5844 (N_5844,N_5455,N_5606);
or U5845 (N_5845,N_5475,N_5653);
nand U5846 (N_5846,N_5479,N_5536);
or U5847 (N_5847,N_5421,N_5553);
xor U5848 (N_5848,N_5546,N_5520);
xnor U5849 (N_5849,N_5690,N_5658);
xor U5850 (N_5850,N_5504,N_5437);
xnor U5851 (N_5851,N_5661,N_5649);
nor U5852 (N_5852,N_5588,N_5669);
and U5853 (N_5853,N_5561,N_5402);
and U5854 (N_5854,N_5557,N_5504);
xnor U5855 (N_5855,N_5608,N_5512);
nor U5856 (N_5856,N_5628,N_5471);
xnor U5857 (N_5857,N_5664,N_5465);
nor U5858 (N_5858,N_5590,N_5575);
and U5859 (N_5859,N_5418,N_5570);
or U5860 (N_5860,N_5572,N_5421);
nand U5861 (N_5861,N_5514,N_5506);
nor U5862 (N_5862,N_5675,N_5688);
nand U5863 (N_5863,N_5694,N_5416);
nor U5864 (N_5864,N_5546,N_5460);
nor U5865 (N_5865,N_5460,N_5558);
nor U5866 (N_5866,N_5699,N_5608);
and U5867 (N_5867,N_5697,N_5550);
or U5868 (N_5868,N_5558,N_5559);
nor U5869 (N_5869,N_5623,N_5484);
xnor U5870 (N_5870,N_5656,N_5552);
xor U5871 (N_5871,N_5558,N_5570);
or U5872 (N_5872,N_5478,N_5538);
xnor U5873 (N_5873,N_5636,N_5489);
or U5874 (N_5874,N_5546,N_5667);
nor U5875 (N_5875,N_5609,N_5424);
nand U5876 (N_5876,N_5591,N_5472);
and U5877 (N_5877,N_5562,N_5504);
nor U5878 (N_5878,N_5427,N_5656);
xnor U5879 (N_5879,N_5623,N_5436);
nand U5880 (N_5880,N_5667,N_5453);
xor U5881 (N_5881,N_5503,N_5541);
nor U5882 (N_5882,N_5650,N_5404);
xor U5883 (N_5883,N_5404,N_5645);
or U5884 (N_5884,N_5594,N_5598);
or U5885 (N_5885,N_5696,N_5626);
xnor U5886 (N_5886,N_5620,N_5462);
or U5887 (N_5887,N_5669,N_5686);
and U5888 (N_5888,N_5587,N_5462);
xnor U5889 (N_5889,N_5419,N_5662);
xnor U5890 (N_5890,N_5624,N_5591);
xnor U5891 (N_5891,N_5413,N_5519);
nor U5892 (N_5892,N_5609,N_5512);
nor U5893 (N_5893,N_5469,N_5500);
or U5894 (N_5894,N_5556,N_5531);
or U5895 (N_5895,N_5506,N_5530);
xor U5896 (N_5896,N_5509,N_5526);
nor U5897 (N_5897,N_5489,N_5494);
and U5898 (N_5898,N_5582,N_5544);
nor U5899 (N_5899,N_5667,N_5521);
nand U5900 (N_5900,N_5555,N_5652);
and U5901 (N_5901,N_5583,N_5601);
nand U5902 (N_5902,N_5470,N_5601);
and U5903 (N_5903,N_5493,N_5555);
and U5904 (N_5904,N_5651,N_5526);
and U5905 (N_5905,N_5627,N_5426);
xor U5906 (N_5906,N_5545,N_5483);
nor U5907 (N_5907,N_5426,N_5519);
xnor U5908 (N_5908,N_5594,N_5601);
xnor U5909 (N_5909,N_5543,N_5669);
and U5910 (N_5910,N_5605,N_5613);
or U5911 (N_5911,N_5548,N_5653);
or U5912 (N_5912,N_5540,N_5616);
nor U5913 (N_5913,N_5625,N_5662);
nand U5914 (N_5914,N_5478,N_5465);
xor U5915 (N_5915,N_5560,N_5627);
and U5916 (N_5916,N_5638,N_5431);
and U5917 (N_5917,N_5491,N_5417);
nand U5918 (N_5918,N_5503,N_5570);
xnor U5919 (N_5919,N_5461,N_5411);
xnor U5920 (N_5920,N_5528,N_5436);
nand U5921 (N_5921,N_5454,N_5559);
xor U5922 (N_5922,N_5563,N_5544);
xnor U5923 (N_5923,N_5636,N_5651);
nand U5924 (N_5924,N_5651,N_5514);
and U5925 (N_5925,N_5475,N_5668);
and U5926 (N_5926,N_5533,N_5647);
or U5927 (N_5927,N_5538,N_5530);
nand U5928 (N_5928,N_5685,N_5435);
nor U5929 (N_5929,N_5630,N_5564);
and U5930 (N_5930,N_5484,N_5549);
or U5931 (N_5931,N_5496,N_5577);
and U5932 (N_5932,N_5479,N_5665);
nand U5933 (N_5933,N_5636,N_5407);
nor U5934 (N_5934,N_5518,N_5691);
or U5935 (N_5935,N_5486,N_5485);
or U5936 (N_5936,N_5646,N_5619);
nand U5937 (N_5937,N_5424,N_5680);
nor U5938 (N_5938,N_5579,N_5687);
and U5939 (N_5939,N_5564,N_5405);
nor U5940 (N_5940,N_5670,N_5669);
nor U5941 (N_5941,N_5506,N_5663);
and U5942 (N_5942,N_5467,N_5525);
or U5943 (N_5943,N_5531,N_5509);
nor U5944 (N_5944,N_5580,N_5403);
and U5945 (N_5945,N_5529,N_5597);
nor U5946 (N_5946,N_5615,N_5510);
xnor U5947 (N_5947,N_5446,N_5652);
or U5948 (N_5948,N_5431,N_5573);
xnor U5949 (N_5949,N_5547,N_5579);
nand U5950 (N_5950,N_5694,N_5599);
and U5951 (N_5951,N_5558,N_5693);
or U5952 (N_5952,N_5527,N_5417);
and U5953 (N_5953,N_5510,N_5523);
xor U5954 (N_5954,N_5609,N_5417);
xnor U5955 (N_5955,N_5508,N_5572);
or U5956 (N_5956,N_5461,N_5408);
and U5957 (N_5957,N_5569,N_5614);
and U5958 (N_5958,N_5476,N_5519);
and U5959 (N_5959,N_5566,N_5434);
nand U5960 (N_5960,N_5673,N_5495);
nand U5961 (N_5961,N_5413,N_5424);
nor U5962 (N_5962,N_5558,N_5489);
or U5963 (N_5963,N_5672,N_5417);
xor U5964 (N_5964,N_5401,N_5679);
or U5965 (N_5965,N_5474,N_5673);
xnor U5966 (N_5966,N_5437,N_5643);
or U5967 (N_5967,N_5696,N_5520);
xor U5968 (N_5968,N_5482,N_5530);
and U5969 (N_5969,N_5481,N_5554);
xnor U5970 (N_5970,N_5521,N_5484);
xor U5971 (N_5971,N_5652,N_5505);
nand U5972 (N_5972,N_5554,N_5552);
nor U5973 (N_5973,N_5636,N_5633);
nor U5974 (N_5974,N_5427,N_5629);
nor U5975 (N_5975,N_5662,N_5679);
nor U5976 (N_5976,N_5582,N_5688);
nand U5977 (N_5977,N_5406,N_5455);
xnor U5978 (N_5978,N_5515,N_5656);
nor U5979 (N_5979,N_5578,N_5647);
and U5980 (N_5980,N_5454,N_5585);
nor U5981 (N_5981,N_5680,N_5594);
nor U5982 (N_5982,N_5699,N_5476);
nand U5983 (N_5983,N_5423,N_5586);
or U5984 (N_5984,N_5589,N_5493);
nand U5985 (N_5985,N_5681,N_5418);
nand U5986 (N_5986,N_5407,N_5445);
xor U5987 (N_5987,N_5590,N_5594);
nor U5988 (N_5988,N_5681,N_5467);
nand U5989 (N_5989,N_5538,N_5698);
and U5990 (N_5990,N_5613,N_5473);
nand U5991 (N_5991,N_5502,N_5590);
nand U5992 (N_5992,N_5585,N_5572);
xor U5993 (N_5993,N_5458,N_5407);
xor U5994 (N_5994,N_5431,N_5461);
and U5995 (N_5995,N_5537,N_5601);
xor U5996 (N_5996,N_5683,N_5469);
xnor U5997 (N_5997,N_5516,N_5414);
nand U5998 (N_5998,N_5475,N_5514);
xnor U5999 (N_5999,N_5693,N_5455);
nor U6000 (N_6000,N_5957,N_5905);
and U6001 (N_6001,N_5755,N_5933);
and U6002 (N_6002,N_5798,N_5738);
nand U6003 (N_6003,N_5716,N_5804);
xor U6004 (N_6004,N_5821,N_5947);
nor U6005 (N_6005,N_5747,N_5976);
and U6006 (N_6006,N_5734,N_5937);
nand U6007 (N_6007,N_5774,N_5919);
or U6008 (N_6008,N_5704,N_5971);
nor U6009 (N_6009,N_5801,N_5997);
nor U6010 (N_6010,N_5956,N_5744);
and U6011 (N_6011,N_5784,N_5881);
and U6012 (N_6012,N_5736,N_5940);
or U6013 (N_6013,N_5979,N_5918);
and U6014 (N_6014,N_5944,N_5724);
xor U6015 (N_6015,N_5785,N_5748);
xnor U6016 (N_6016,N_5896,N_5728);
xnor U6017 (N_6017,N_5890,N_5843);
nor U6018 (N_6018,N_5946,N_5838);
or U6019 (N_6019,N_5993,N_5851);
or U6020 (N_6020,N_5799,N_5786);
xnor U6021 (N_6021,N_5833,N_5953);
nand U6022 (N_6022,N_5977,N_5795);
xor U6023 (N_6023,N_5768,N_5968);
nand U6024 (N_6024,N_5846,N_5988);
xnor U6025 (N_6025,N_5875,N_5845);
nor U6026 (N_6026,N_5871,N_5816);
or U6027 (N_6027,N_5809,N_5951);
and U6028 (N_6028,N_5961,N_5818);
or U6029 (N_6029,N_5925,N_5757);
and U6030 (N_6030,N_5745,N_5835);
and U6031 (N_6031,N_5863,N_5797);
and U6032 (N_6032,N_5888,N_5964);
xnor U6033 (N_6033,N_5952,N_5852);
xor U6034 (N_6034,N_5989,N_5751);
and U6035 (N_6035,N_5778,N_5802);
xor U6036 (N_6036,N_5707,N_5730);
nand U6037 (N_6037,N_5939,N_5913);
nor U6038 (N_6038,N_5753,N_5883);
and U6039 (N_6039,N_5858,N_5878);
nand U6040 (N_6040,N_5721,N_5931);
xor U6041 (N_6041,N_5991,N_5741);
or U6042 (N_6042,N_5752,N_5932);
nand U6043 (N_6043,N_5959,N_5763);
and U6044 (N_6044,N_5733,N_5807);
nor U6045 (N_6045,N_5822,N_5897);
nor U6046 (N_6046,N_5782,N_5998);
or U6047 (N_6047,N_5815,N_5781);
and U6048 (N_6048,N_5893,N_5914);
nor U6049 (N_6049,N_5864,N_5805);
nand U6050 (N_6050,N_5826,N_5819);
nor U6051 (N_6051,N_5723,N_5894);
and U6052 (N_6052,N_5916,N_5901);
nor U6053 (N_6053,N_5794,N_5986);
xnor U6054 (N_6054,N_5746,N_5739);
nand U6055 (N_6055,N_5941,N_5963);
nor U6056 (N_6056,N_5907,N_5743);
nor U6057 (N_6057,N_5840,N_5823);
xor U6058 (N_6058,N_5992,N_5856);
nand U6059 (N_6059,N_5985,N_5727);
nand U6060 (N_6060,N_5754,N_5880);
xnor U6061 (N_6061,N_5859,N_5970);
or U6062 (N_6062,N_5814,N_5983);
nand U6063 (N_6063,N_5995,N_5712);
nor U6064 (N_6064,N_5965,N_5892);
and U6065 (N_6065,N_5974,N_5788);
or U6066 (N_6066,N_5836,N_5714);
nand U6067 (N_6067,N_5762,N_5972);
nand U6068 (N_6068,N_5954,N_5761);
nand U6069 (N_6069,N_5708,N_5792);
and U6070 (N_6070,N_5984,N_5866);
nor U6071 (N_6071,N_5975,N_5742);
nand U6072 (N_6072,N_5766,N_5830);
xor U6073 (N_6073,N_5879,N_5718);
nand U6074 (N_6074,N_5829,N_5771);
nand U6075 (N_6075,N_5760,N_5732);
or U6076 (N_6076,N_5839,N_5740);
and U6077 (N_6077,N_5715,N_5719);
nor U6078 (N_6078,N_5924,N_5865);
and U6079 (N_6079,N_5789,N_5872);
or U6080 (N_6080,N_5926,N_5731);
xnor U6081 (N_6081,N_5790,N_5960);
nand U6082 (N_6082,N_5780,N_5834);
nor U6083 (N_6083,N_5831,N_5796);
nor U6084 (N_6084,N_5770,N_5950);
xor U6085 (N_6085,N_5793,N_5729);
xor U6086 (N_6086,N_5713,N_5764);
xor U6087 (N_6087,N_5874,N_5868);
or U6088 (N_6088,N_5806,N_5994);
nand U6089 (N_6089,N_5981,N_5904);
or U6090 (N_6090,N_5756,N_5808);
nor U6091 (N_6091,N_5709,N_5917);
nand U6092 (N_6092,N_5943,N_5767);
nor U6093 (N_6093,N_5921,N_5710);
nor U6094 (N_6094,N_5899,N_5886);
nand U6095 (N_6095,N_5922,N_5870);
xnor U6096 (N_6096,N_5720,N_5955);
nor U6097 (N_6097,N_5777,N_5882);
and U6098 (N_6098,N_5810,N_5895);
or U6099 (N_6099,N_5949,N_5800);
or U6100 (N_6100,N_5999,N_5987);
nor U6101 (N_6101,N_5817,N_5824);
nor U6102 (N_6102,N_5832,N_5735);
nor U6103 (N_6103,N_5759,N_5711);
and U6104 (N_6104,N_5930,N_5705);
xor U6105 (N_6105,N_5854,N_5825);
nor U6106 (N_6106,N_5876,N_5857);
nor U6107 (N_6107,N_5750,N_5844);
nand U6108 (N_6108,N_5702,N_5869);
xnor U6109 (N_6109,N_5722,N_5929);
or U6110 (N_6110,N_5725,N_5912);
xor U6111 (N_6111,N_5841,N_5812);
nand U6112 (N_6112,N_5980,N_5915);
nor U6113 (N_6113,N_5967,N_5966);
or U6114 (N_6114,N_5700,N_5811);
xnor U6115 (N_6115,N_5927,N_5948);
nor U6116 (N_6116,N_5758,N_5920);
or U6117 (N_6117,N_5906,N_5982);
and U6118 (N_6118,N_5820,N_5706);
nor U6119 (N_6119,N_5910,N_5911);
and U6120 (N_6120,N_5884,N_5848);
nand U6121 (N_6121,N_5853,N_5978);
or U6122 (N_6122,N_5773,N_5828);
or U6123 (N_6123,N_5873,N_5934);
nand U6124 (N_6124,N_5779,N_5765);
and U6125 (N_6125,N_5850,N_5887);
nand U6126 (N_6126,N_5737,N_5775);
xor U6127 (N_6127,N_5958,N_5885);
or U6128 (N_6128,N_5772,N_5962);
xnor U6129 (N_6129,N_5776,N_5938);
or U6130 (N_6130,N_5701,N_5726);
xnor U6131 (N_6131,N_5935,N_5849);
nand U6132 (N_6132,N_5827,N_5837);
and U6133 (N_6133,N_5898,N_5889);
nand U6134 (N_6134,N_5791,N_5902);
nand U6135 (N_6135,N_5703,N_5783);
and U6136 (N_6136,N_5909,N_5973);
and U6137 (N_6137,N_5936,N_5945);
nand U6138 (N_6138,N_5903,N_5867);
nor U6139 (N_6139,N_5855,N_5862);
nor U6140 (N_6140,N_5928,N_5717);
nor U6141 (N_6141,N_5996,N_5847);
xnor U6142 (N_6142,N_5813,N_5990);
nor U6143 (N_6143,N_5842,N_5923);
and U6144 (N_6144,N_5803,N_5900);
nor U6145 (N_6145,N_5877,N_5891);
nor U6146 (N_6146,N_5787,N_5749);
xor U6147 (N_6147,N_5942,N_5769);
xnor U6148 (N_6148,N_5860,N_5908);
nand U6149 (N_6149,N_5861,N_5969);
and U6150 (N_6150,N_5768,N_5926);
nor U6151 (N_6151,N_5783,N_5792);
xnor U6152 (N_6152,N_5837,N_5881);
nor U6153 (N_6153,N_5767,N_5935);
and U6154 (N_6154,N_5848,N_5969);
nand U6155 (N_6155,N_5757,N_5870);
nor U6156 (N_6156,N_5740,N_5883);
or U6157 (N_6157,N_5803,N_5738);
nand U6158 (N_6158,N_5776,N_5827);
or U6159 (N_6159,N_5723,N_5926);
xnor U6160 (N_6160,N_5734,N_5777);
nand U6161 (N_6161,N_5811,N_5942);
and U6162 (N_6162,N_5772,N_5750);
or U6163 (N_6163,N_5853,N_5709);
nand U6164 (N_6164,N_5991,N_5719);
nand U6165 (N_6165,N_5752,N_5968);
or U6166 (N_6166,N_5953,N_5881);
and U6167 (N_6167,N_5903,N_5852);
nor U6168 (N_6168,N_5860,N_5918);
xor U6169 (N_6169,N_5891,N_5995);
and U6170 (N_6170,N_5855,N_5816);
nand U6171 (N_6171,N_5976,N_5785);
nand U6172 (N_6172,N_5774,N_5717);
nor U6173 (N_6173,N_5760,N_5803);
nand U6174 (N_6174,N_5742,N_5897);
and U6175 (N_6175,N_5881,N_5942);
nor U6176 (N_6176,N_5829,N_5840);
xnor U6177 (N_6177,N_5765,N_5966);
or U6178 (N_6178,N_5731,N_5794);
nor U6179 (N_6179,N_5915,N_5839);
and U6180 (N_6180,N_5839,N_5714);
and U6181 (N_6181,N_5901,N_5750);
nand U6182 (N_6182,N_5961,N_5791);
or U6183 (N_6183,N_5853,N_5842);
nand U6184 (N_6184,N_5837,N_5924);
and U6185 (N_6185,N_5780,N_5927);
nand U6186 (N_6186,N_5912,N_5965);
nor U6187 (N_6187,N_5733,N_5935);
nand U6188 (N_6188,N_5955,N_5797);
and U6189 (N_6189,N_5865,N_5945);
xnor U6190 (N_6190,N_5942,N_5996);
and U6191 (N_6191,N_5707,N_5720);
nand U6192 (N_6192,N_5872,N_5790);
xnor U6193 (N_6193,N_5732,N_5885);
xor U6194 (N_6194,N_5728,N_5810);
nor U6195 (N_6195,N_5873,N_5955);
nor U6196 (N_6196,N_5701,N_5872);
and U6197 (N_6197,N_5770,N_5889);
or U6198 (N_6198,N_5765,N_5875);
and U6199 (N_6199,N_5880,N_5798);
and U6200 (N_6200,N_5766,N_5818);
xnor U6201 (N_6201,N_5841,N_5915);
or U6202 (N_6202,N_5977,N_5999);
nand U6203 (N_6203,N_5796,N_5801);
and U6204 (N_6204,N_5731,N_5836);
xnor U6205 (N_6205,N_5763,N_5854);
and U6206 (N_6206,N_5827,N_5910);
nand U6207 (N_6207,N_5848,N_5877);
xor U6208 (N_6208,N_5867,N_5949);
or U6209 (N_6209,N_5982,N_5725);
or U6210 (N_6210,N_5915,N_5793);
and U6211 (N_6211,N_5839,N_5930);
xor U6212 (N_6212,N_5774,N_5726);
nor U6213 (N_6213,N_5839,N_5720);
xnor U6214 (N_6214,N_5918,N_5858);
or U6215 (N_6215,N_5890,N_5775);
or U6216 (N_6216,N_5924,N_5841);
nand U6217 (N_6217,N_5823,N_5904);
and U6218 (N_6218,N_5931,N_5978);
xor U6219 (N_6219,N_5818,N_5804);
and U6220 (N_6220,N_5979,N_5976);
or U6221 (N_6221,N_5847,N_5921);
or U6222 (N_6222,N_5915,N_5747);
xor U6223 (N_6223,N_5897,N_5788);
nor U6224 (N_6224,N_5797,N_5834);
or U6225 (N_6225,N_5984,N_5889);
nand U6226 (N_6226,N_5726,N_5979);
and U6227 (N_6227,N_5787,N_5755);
or U6228 (N_6228,N_5763,N_5900);
nand U6229 (N_6229,N_5851,N_5744);
xnor U6230 (N_6230,N_5912,N_5759);
or U6231 (N_6231,N_5959,N_5802);
or U6232 (N_6232,N_5755,N_5712);
xor U6233 (N_6233,N_5876,N_5933);
or U6234 (N_6234,N_5709,N_5948);
nand U6235 (N_6235,N_5703,N_5739);
or U6236 (N_6236,N_5896,N_5836);
xor U6237 (N_6237,N_5769,N_5890);
and U6238 (N_6238,N_5971,N_5950);
xnor U6239 (N_6239,N_5908,N_5958);
xor U6240 (N_6240,N_5839,N_5776);
xnor U6241 (N_6241,N_5987,N_5956);
xnor U6242 (N_6242,N_5748,N_5718);
nor U6243 (N_6243,N_5919,N_5841);
nor U6244 (N_6244,N_5995,N_5808);
nor U6245 (N_6245,N_5864,N_5843);
and U6246 (N_6246,N_5936,N_5732);
nor U6247 (N_6247,N_5962,N_5958);
nand U6248 (N_6248,N_5967,N_5986);
nand U6249 (N_6249,N_5901,N_5919);
or U6250 (N_6250,N_5780,N_5857);
nor U6251 (N_6251,N_5752,N_5971);
xor U6252 (N_6252,N_5860,N_5823);
or U6253 (N_6253,N_5701,N_5953);
or U6254 (N_6254,N_5963,N_5911);
or U6255 (N_6255,N_5749,N_5812);
nor U6256 (N_6256,N_5716,N_5761);
or U6257 (N_6257,N_5703,N_5928);
and U6258 (N_6258,N_5988,N_5927);
xor U6259 (N_6259,N_5923,N_5803);
nand U6260 (N_6260,N_5786,N_5761);
xor U6261 (N_6261,N_5928,N_5793);
nand U6262 (N_6262,N_5921,N_5864);
xor U6263 (N_6263,N_5880,N_5775);
and U6264 (N_6264,N_5936,N_5770);
xor U6265 (N_6265,N_5934,N_5797);
or U6266 (N_6266,N_5936,N_5986);
nand U6267 (N_6267,N_5978,N_5980);
xor U6268 (N_6268,N_5832,N_5894);
and U6269 (N_6269,N_5815,N_5944);
nand U6270 (N_6270,N_5847,N_5750);
nor U6271 (N_6271,N_5967,N_5728);
nand U6272 (N_6272,N_5745,N_5754);
nor U6273 (N_6273,N_5747,N_5918);
nor U6274 (N_6274,N_5882,N_5989);
xnor U6275 (N_6275,N_5943,N_5798);
xnor U6276 (N_6276,N_5757,N_5908);
or U6277 (N_6277,N_5818,N_5997);
nor U6278 (N_6278,N_5895,N_5955);
nand U6279 (N_6279,N_5894,N_5813);
or U6280 (N_6280,N_5732,N_5896);
and U6281 (N_6281,N_5826,N_5762);
nand U6282 (N_6282,N_5703,N_5893);
or U6283 (N_6283,N_5827,N_5768);
nand U6284 (N_6284,N_5845,N_5899);
xor U6285 (N_6285,N_5954,N_5823);
nand U6286 (N_6286,N_5883,N_5832);
nor U6287 (N_6287,N_5805,N_5976);
nand U6288 (N_6288,N_5722,N_5892);
or U6289 (N_6289,N_5916,N_5765);
nand U6290 (N_6290,N_5819,N_5989);
or U6291 (N_6291,N_5830,N_5916);
nand U6292 (N_6292,N_5802,N_5769);
xnor U6293 (N_6293,N_5764,N_5965);
and U6294 (N_6294,N_5892,N_5936);
nand U6295 (N_6295,N_5747,N_5709);
nand U6296 (N_6296,N_5705,N_5986);
nor U6297 (N_6297,N_5979,N_5936);
and U6298 (N_6298,N_5898,N_5803);
nand U6299 (N_6299,N_5825,N_5945);
nand U6300 (N_6300,N_6243,N_6079);
or U6301 (N_6301,N_6042,N_6225);
nor U6302 (N_6302,N_6148,N_6230);
nand U6303 (N_6303,N_6204,N_6144);
xnor U6304 (N_6304,N_6129,N_6086);
nor U6305 (N_6305,N_6299,N_6223);
xor U6306 (N_6306,N_6232,N_6047);
nor U6307 (N_6307,N_6192,N_6116);
xnor U6308 (N_6308,N_6215,N_6155);
nand U6309 (N_6309,N_6081,N_6006);
nand U6310 (N_6310,N_6183,N_6197);
nand U6311 (N_6311,N_6083,N_6007);
and U6312 (N_6312,N_6040,N_6093);
nor U6313 (N_6313,N_6062,N_6017);
or U6314 (N_6314,N_6005,N_6294);
xor U6315 (N_6315,N_6010,N_6201);
xnor U6316 (N_6316,N_6291,N_6246);
or U6317 (N_6317,N_6067,N_6241);
and U6318 (N_6318,N_6198,N_6180);
and U6319 (N_6319,N_6045,N_6173);
xnor U6320 (N_6320,N_6004,N_6031);
nand U6321 (N_6321,N_6100,N_6165);
and U6322 (N_6322,N_6097,N_6018);
or U6323 (N_6323,N_6278,N_6267);
and U6324 (N_6324,N_6207,N_6084);
nor U6325 (N_6325,N_6039,N_6104);
or U6326 (N_6326,N_6150,N_6187);
or U6327 (N_6327,N_6235,N_6111);
nor U6328 (N_6328,N_6221,N_6055);
nor U6329 (N_6329,N_6049,N_6222);
and U6330 (N_6330,N_6191,N_6119);
and U6331 (N_6331,N_6106,N_6022);
and U6332 (N_6332,N_6189,N_6029);
or U6333 (N_6333,N_6174,N_6147);
and U6334 (N_6334,N_6070,N_6082);
and U6335 (N_6335,N_6271,N_6091);
nor U6336 (N_6336,N_6151,N_6098);
nand U6337 (N_6337,N_6186,N_6169);
xnor U6338 (N_6338,N_6156,N_6256);
nor U6339 (N_6339,N_6279,N_6126);
xnor U6340 (N_6340,N_6009,N_6142);
nand U6341 (N_6341,N_6120,N_6238);
and U6342 (N_6342,N_6060,N_6133);
nand U6343 (N_6343,N_6074,N_6273);
xor U6344 (N_6344,N_6185,N_6196);
nor U6345 (N_6345,N_6037,N_6228);
and U6346 (N_6346,N_6208,N_6252);
or U6347 (N_6347,N_6154,N_6131);
nand U6348 (N_6348,N_6143,N_6023);
and U6349 (N_6349,N_6021,N_6167);
nor U6350 (N_6350,N_6063,N_6003);
xor U6351 (N_6351,N_6292,N_6134);
or U6352 (N_6352,N_6193,N_6015);
nor U6353 (N_6353,N_6240,N_6262);
and U6354 (N_6354,N_6001,N_6224);
xor U6355 (N_6355,N_6059,N_6163);
nand U6356 (N_6356,N_6088,N_6212);
and U6357 (N_6357,N_6289,N_6166);
and U6358 (N_6358,N_6188,N_6138);
or U6359 (N_6359,N_6195,N_6056);
nor U6360 (N_6360,N_6213,N_6216);
xnor U6361 (N_6361,N_6094,N_6058);
nand U6362 (N_6362,N_6176,N_6105);
or U6363 (N_6363,N_6096,N_6233);
or U6364 (N_6364,N_6244,N_6264);
or U6365 (N_6365,N_6051,N_6122);
and U6366 (N_6366,N_6219,N_6121);
nand U6367 (N_6367,N_6118,N_6260);
or U6368 (N_6368,N_6234,N_6113);
or U6369 (N_6369,N_6136,N_6046);
nor U6370 (N_6370,N_6229,N_6161);
and U6371 (N_6371,N_6170,N_6175);
and U6372 (N_6372,N_6107,N_6297);
nor U6373 (N_6373,N_6251,N_6130);
or U6374 (N_6374,N_6227,N_6149);
nand U6375 (N_6375,N_6019,N_6044);
nor U6376 (N_6376,N_6011,N_6034);
nor U6377 (N_6377,N_6290,N_6199);
nand U6378 (N_6378,N_6179,N_6135);
or U6379 (N_6379,N_6008,N_6205);
xor U6380 (N_6380,N_6069,N_6050);
or U6381 (N_6381,N_6035,N_6048);
or U6382 (N_6382,N_6024,N_6065);
nand U6383 (N_6383,N_6277,N_6020);
nor U6384 (N_6384,N_6249,N_6068);
or U6385 (N_6385,N_6171,N_6190);
nor U6386 (N_6386,N_6139,N_6128);
xor U6387 (N_6387,N_6092,N_6280);
or U6388 (N_6388,N_6028,N_6200);
or U6389 (N_6389,N_6247,N_6132);
nor U6390 (N_6390,N_6285,N_6209);
nand U6391 (N_6391,N_6159,N_6158);
or U6392 (N_6392,N_6282,N_6080);
xor U6393 (N_6393,N_6057,N_6102);
nand U6394 (N_6394,N_6089,N_6283);
xor U6395 (N_6395,N_6178,N_6101);
nand U6396 (N_6396,N_6265,N_6027);
and U6397 (N_6397,N_6012,N_6239);
or U6398 (N_6398,N_6206,N_6066);
or U6399 (N_6399,N_6014,N_6254);
nand U6400 (N_6400,N_6077,N_6250);
nor U6401 (N_6401,N_6172,N_6274);
and U6402 (N_6402,N_6182,N_6184);
and U6403 (N_6403,N_6153,N_6257);
nand U6404 (N_6404,N_6276,N_6293);
or U6405 (N_6405,N_6090,N_6269);
or U6406 (N_6406,N_6203,N_6054);
nor U6407 (N_6407,N_6259,N_6103);
or U6408 (N_6408,N_6275,N_6125);
nand U6409 (N_6409,N_6085,N_6123);
nand U6410 (N_6410,N_6245,N_6115);
nor U6411 (N_6411,N_6272,N_6127);
and U6412 (N_6412,N_6078,N_6052);
nand U6413 (N_6413,N_6258,N_6016);
or U6414 (N_6414,N_6043,N_6287);
xor U6415 (N_6415,N_6168,N_6137);
or U6416 (N_6416,N_6268,N_6284);
nand U6417 (N_6417,N_6073,N_6164);
and U6418 (N_6418,N_6002,N_6177);
and U6419 (N_6419,N_6095,N_6160);
or U6420 (N_6420,N_6237,N_6236);
nor U6421 (N_6421,N_6072,N_6036);
xnor U6422 (N_6422,N_6162,N_6026);
nand U6423 (N_6423,N_6263,N_6099);
xnor U6424 (N_6424,N_6140,N_6053);
nand U6425 (N_6425,N_6033,N_6087);
nor U6426 (N_6426,N_6261,N_6210);
xnor U6427 (N_6427,N_6226,N_6038);
or U6428 (N_6428,N_6231,N_6194);
or U6429 (N_6429,N_6124,N_6061);
and U6430 (N_6430,N_6266,N_6109);
nand U6431 (N_6431,N_6253,N_6114);
and U6432 (N_6432,N_6220,N_6288);
nor U6433 (N_6433,N_6298,N_6108);
nand U6434 (N_6434,N_6255,N_6286);
nor U6435 (N_6435,N_6157,N_6281);
nor U6436 (N_6436,N_6217,N_6025);
and U6437 (N_6437,N_6202,N_6032);
nor U6438 (N_6438,N_6075,N_6117);
nand U6439 (N_6439,N_6152,N_6141);
and U6440 (N_6440,N_6076,N_6013);
and U6441 (N_6441,N_6218,N_6295);
and U6442 (N_6442,N_6270,N_6242);
nand U6443 (N_6443,N_6145,N_6064);
and U6444 (N_6444,N_6211,N_6146);
nand U6445 (N_6445,N_6112,N_6181);
and U6446 (N_6446,N_6296,N_6248);
or U6447 (N_6447,N_6030,N_6041);
xor U6448 (N_6448,N_6071,N_6000);
and U6449 (N_6449,N_6110,N_6214);
nand U6450 (N_6450,N_6177,N_6045);
and U6451 (N_6451,N_6234,N_6178);
nand U6452 (N_6452,N_6106,N_6029);
and U6453 (N_6453,N_6282,N_6176);
nand U6454 (N_6454,N_6295,N_6191);
and U6455 (N_6455,N_6163,N_6211);
or U6456 (N_6456,N_6096,N_6105);
or U6457 (N_6457,N_6170,N_6200);
xnor U6458 (N_6458,N_6046,N_6267);
nor U6459 (N_6459,N_6093,N_6082);
nor U6460 (N_6460,N_6116,N_6239);
nor U6461 (N_6461,N_6268,N_6250);
xnor U6462 (N_6462,N_6247,N_6060);
xnor U6463 (N_6463,N_6124,N_6048);
or U6464 (N_6464,N_6012,N_6213);
xnor U6465 (N_6465,N_6074,N_6096);
or U6466 (N_6466,N_6036,N_6047);
or U6467 (N_6467,N_6163,N_6298);
nor U6468 (N_6468,N_6165,N_6235);
nor U6469 (N_6469,N_6204,N_6021);
and U6470 (N_6470,N_6152,N_6201);
or U6471 (N_6471,N_6122,N_6081);
and U6472 (N_6472,N_6045,N_6052);
or U6473 (N_6473,N_6152,N_6109);
or U6474 (N_6474,N_6264,N_6108);
nor U6475 (N_6475,N_6049,N_6064);
or U6476 (N_6476,N_6132,N_6288);
and U6477 (N_6477,N_6085,N_6005);
or U6478 (N_6478,N_6267,N_6149);
nor U6479 (N_6479,N_6239,N_6086);
nand U6480 (N_6480,N_6130,N_6112);
or U6481 (N_6481,N_6199,N_6189);
nand U6482 (N_6482,N_6051,N_6054);
or U6483 (N_6483,N_6007,N_6294);
or U6484 (N_6484,N_6248,N_6064);
xor U6485 (N_6485,N_6175,N_6108);
or U6486 (N_6486,N_6143,N_6224);
nand U6487 (N_6487,N_6026,N_6021);
and U6488 (N_6488,N_6091,N_6041);
and U6489 (N_6489,N_6015,N_6026);
nand U6490 (N_6490,N_6191,N_6231);
nor U6491 (N_6491,N_6231,N_6062);
nor U6492 (N_6492,N_6178,N_6027);
or U6493 (N_6493,N_6099,N_6199);
nand U6494 (N_6494,N_6004,N_6092);
xnor U6495 (N_6495,N_6008,N_6075);
xor U6496 (N_6496,N_6067,N_6262);
nand U6497 (N_6497,N_6115,N_6267);
nor U6498 (N_6498,N_6093,N_6253);
nor U6499 (N_6499,N_6181,N_6109);
nor U6500 (N_6500,N_6160,N_6058);
xor U6501 (N_6501,N_6028,N_6088);
and U6502 (N_6502,N_6236,N_6139);
and U6503 (N_6503,N_6218,N_6288);
or U6504 (N_6504,N_6006,N_6230);
xnor U6505 (N_6505,N_6235,N_6249);
nor U6506 (N_6506,N_6098,N_6052);
or U6507 (N_6507,N_6000,N_6271);
or U6508 (N_6508,N_6174,N_6210);
xor U6509 (N_6509,N_6168,N_6052);
or U6510 (N_6510,N_6019,N_6279);
nand U6511 (N_6511,N_6271,N_6027);
or U6512 (N_6512,N_6216,N_6011);
and U6513 (N_6513,N_6262,N_6023);
and U6514 (N_6514,N_6248,N_6264);
nor U6515 (N_6515,N_6240,N_6250);
xor U6516 (N_6516,N_6169,N_6059);
nor U6517 (N_6517,N_6173,N_6242);
or U6518 (N_6518,N_6212,N_6218);
or U6519 (N_6519,N_6065,N_6230);
and U6520 (N_6520,N_6221,N_6001);
or U6521 (N_6521,N_6128,N_6093);
nor U6522 (N_6522,N_6148,N_6155);
xnor U6523 (N_6523,N_6295,N_6129);
or U6524 (N_6524,N_6246,N_6025);
or U6525 (N_6525,N_6202,N_6219);
or U6526 (N_6526,N_6293,N_6167);
and U6527 (N_6527,N_6135,N_6195);
nor U6528 (N_6528,N_6089,N_6032);
or U6529 (N_6529,N_6122,N_6178);
nand U6530 (N_6530,N_6176,N_6109);
nor U6531 (N_6531,N_6132,N_6138);
nand U6532 (N_6532,N_6064,N_6029);
nand U6533 (N_6533,N_6131,N_6058);
xor U6534 (N_6534,N_6091,N_6143);
or U6535 (N_6535,N_6105,N_6117);
nor U6536 (N_6536,N_6215,N_6154);
nor U6537 (N_6537,N_6226,N_6129);
xor U6538 (N_6538,N_6289,N_6085);
xor U6539 (N_6539,N_6118,N_6075);
or U6540 (N_6540,N_6263,N_6255);
and U6541 (N_6541,N_6007,N_6200);
or U6542 (N_6542,N_6149,N_6244);
xor U6543 (N_6543,N_6061,N_6010);
and U6544 (N_6544,N_6012,N_6030);
nor U6545 (N_6545,N_6196,N_6183);
nor U6546 (N_6546,N_6269,N_6150);
or U6547 (N_6547,N_6213,N_6039);
nand U6548 (N_6548,N_6171,N_6282);
nand U6549 (N_6549,N_6290,N_6019);
xnor U6550 (N_6550,N_6086,N_6202);
xor U6551 (N_6551,N_6209,N_6060);
and U6552 (N_6552,N_6138,N_6090);
or U6553 (N_6553,N_6230,N_6144);
and U6554 (N_6554,N_6131,N_6245);
nor U6555 (N_6555,N_6012,N_6194);
or U6556 (N_6556,N_6267,N_6231);
and U6557 (N_6557,N_6008,N_6162);
or U6558 (N_6558,N_6237,N_6032);
or U6559 (N_6559,N_6177,N_6138);
nand U6560 (N_6560,N_6125,N_6212);
and U6561 (N_6561,N_6284,N_6006);
and U6562 (N_6562,N_6245,N_6295);
nor U6563 (N_6563,N_6068,N_6246);
nand U6564 (N_6564,N_6005,N_6213);
nor U6565 (N_6565,N_6146,N_6114);
or U6566 (N_6566,N_6102,N_6293);
or U6567 (N_6567,N_6276,N_6012);
nand U6568 (N_6568,N_6139,N_6168);
xnor U6569 (N_6569,N_6038,N_6248);
xor U6570 (N_6570,N_6219,N_6281);
nand U6571 (N_6571,N_6262,N_6168);
nor U6572 (N_6572,N_6121,N_6009);
or U6573 (N_6573,N_6166,N_6236);
nor U6574 (N_6574,N_6263,N_6161);
xor U6575 (N_6575,N_6248,N_6259);
and U6576 (N_6576,N_6034,N_6277);
nor U6577 (N_6577,N_6272,N_6100);
or U6578 (N_6578,N_6292,N_6285);
and U6579 (N_6579,N_6056,N_6000);
xor U6580 (N_6580,N_6118,N_6093);
or U6581 (N_6581,N_6270,N_6040);
and U6582 (N_6582,N_6049,N_6018);
and U6583 (N_6583,N_6273,N_6149);
and U6584 (N_6584,N_6120,N_6257);
nor U6585 (N_6585,N_6167,N_6160);
and U6586 (N_6586,N_6131,N_6031);
nor U6587 (N_6587,N_6249,N_6124);
and U6588 (N_6588,N_6298,N_6070);
nand U6589 (N_6589,N_6102,N_6028);
and U6590 (N_6590,N_6118,N_6277);
xnor U6591 (N_6591,N_6158,N_6110);
or U6592 (N_6592,N_6016,N_6043);
xnor U6593 (N_6593,N_6065,N_6157);
nand U6594 (N_6594,N_6149,N_6295);
nor U6595 (N_6595,N_6223,N_6227);
xnor U6596 (N_6596,N_6113,N_6252);
nor U6597 (N_6597,N_6065,N_6237);
nor U6598 (N_6598,N_6032,N_6176);
nor U6599 (N_6599,N_6151,N_6099);
xnor U6600 (N_6600,N_6516,N_6572);
nand U6601 (N_6601,N_6519,N_6522);
or U6602 (N_6602,N_6472,N_6323);
nand U6603 (N_6603,N_6509,N_6526);
xnor U6604 (N_6604,N_6448,N_6332);
and U6605 (N_6605,N_6417,N_6442);
or U6606 (N_6606,N_6569,N_6549);
nor U6607 (N_6607,N_6588,N_6508);
and U6608 (N_6608,N_6398,N_6386);
or U6609 (N_6609,N_6401,N_6496);
nand U6610 (N_6610,N_6498,N_6330);
or U6611 (N_6611,N_6358,N_6598);
or U6612 (N_6612,N_6543,N_6435);
or U6613 (N_6613,N_6345,N_6337);
and U6614 (N_6614,N_6438,N_6577);
and U6615 (N_6615,N_6404,N_6445);
nand U6616 (N_6616,N_6385,N_6562);
nand U6617 (N_6617,N_6411,N_6425);
nor U6618 (N_6618,N_6497,N_6314);
xnor U6619 (N_6619,N_6304,N_6322);
nor U6620 (N_6620,N_6461,N_6454);
nor U6621 (N_6621,N_6499,N_6450);
or U6622 (N_6622,N_6372,N_6548);
nand U6623 (N_6623,N_6431,N_6556);
or U6624 (N_6624,N_6343,N_6436);
nand U6625 (N_6625,N_6441,N_6570);
or U6626 (N_6626,N_6467,N_6301);
nand U6627 (N_6627,N_6426,N_6381);
nor U6628 (N_6628,N_6429,N_6432);
and U6629 (N_6629,N_6525,N_6300);
nand U6630 (N_6630,N_6592,N_6527);
nor U6631 (N_6631,N_6453,N_6489);
nand U6632 (N_6632,N_6446,N_6494);
xor U6633 (N_6633,N_6424,N_6511);
xnor U6634 (N_6634,N_6319,N_6303);
xor U6635 (N_6635,N_6483,N_6477);
and U6636 (N_6636,N_6523,N_6528);
nor U6637 (N_6637,N_6479,N_6474);
or U6638 (N_6638,N_6360,N_6574);
xor U6639 (N_6639,N_6334,N_6378);
xnor U6640 (N_6640,N_6542,N_6493);
and U6641 (N_6641,N_6410,N_6469);
or U6642 (N_6642,N_6407,N_6532);
nand U6643 (N_6643,N_6536,N_6544);
and U6644 (N_6644,N_6566,N_6357);
xnor U6645 (N_6645,N_6539,N_6375);
or U6646 (N_6646,N_6503,N_6309);
and U6647 (N_6647,N_6463,N_6590);
nand U6648 (N_6648,N_6355,N_6595);
nor U6649 (N_6649,N_6406,N_6465);
and U6650 (N_6650,N_6328,N_6529);
nand U6651 (N_6651,N_6305,N_6505);
xor U6652 (N_6652,N_6361,N_6338);
or U6653 (N_6653,N_6430,N_6391);
nand U6654 (N_6654,N_6537,N_6356);
nand U6655 (N_6655,N_6437,N_6485);
or U6656 (N_6656,N_6571,N_6374);
xor U6657 (N_6657,N_6473,N_6462);
nor U6658 (N_6658,N_6597,N_6351);
nor U6659 (N_6659,N_6315,N_6513);
nor U6660 (N_6660,N_6333,N_6563);
xnor U6661 (N_6661,N_6444,N_6575);
nor U6662 (N_6662,N_6504,N_6546);
xor U6663 (N_6663,N_6587,N_6501);
nand U6664 (N_6664,N_6383,N_6555);
or U6665 (N_6665,N_6567,N_6524);
and U6666 (N_6666,N_6369,N_6326);
xnor U6667 (N_6667,N_6554,N_6565);
and U6668 (N_6668,N_6584,N_6388);
nand U6669 (N_6669,N_6400,N_6415);
or U6670 (N_6670,N_6558,N_6422);
and U6671 (N_6671,N_6510,N_6413);
nor U6672 (N_6672,N_6327,N_6578);
nor U6673 (N_6673,N_6373,N_6387);
nand U6674 (N_6674,N_6395,N_6346);
xor U6675 (N_6675,N_6390,N_6427);
nand U6676 (N_6676,N_6486,N_6347);
or U6677 (N_6677,N_6311,N_6409);
or U6678 (N_6678,N_6335,N_6443);
and U6679 (N_6679,N_6439,N_6460);
or U6680 (N_6680,N_6302,N_6487);
nand U6681 (N_6681,N_6321,N_6350);
nand U6682 (N_6682,N_6541,N_6568);
nand U6683 (N_6683,N_6371,N_6457);
xnor U6684 (N_6684,N_6405,N_6455);
nor U6685 (N_6685,N_6476,N_6550);
or U6686 (N_6686,N_6582,N_6354);
xor U6687 (N_6687,N_6363,N_6480);
nand U6688 (N_6688,N_6403,N_6515);
xor U6689 (N_6689,N_6530,N_6306);
nor U6690 (N_6690,N_6420,N_6464);
and U6691 (N_6691,N_6557,N_6320);
nand U6692 (N_6692,N_6456,N_6331);
or U6693 (N_6693,N_6325,N_6377);
or U6694 (N_6694,N_6394,N_6312);
or U6695 (N_6695,N_6396,N_6553);
xor U6696 (N_6696,N_6589,N_6397);
nand U6697 (N_6697,N_6418,N_6490);
and U6698 (N_6698,N_6492,N_6561);
and U6699 (N_6699,N_6491,N_6416);
xor U6700 (N_6700,N_6535,N_6352);
or U6701 (N_6701,N_6545,N_6596);
or U6702 (N_6702,N_6339,N_6399);
nand U6703 (N_6703,N_6517,N_6583);
xnor U6704 (N_6704,N_6307,N_6324);
xnor U6705 (N_6705,N_6471,N_6336);
xor U6706 (N_6706,N_6440,N_6580);
and U6707 (N_6707,N_6475,N_6362);
nor U6708 (N_6708,N_6470,N_6507);
and U6709 (N_6709,N_6308,N_6342);
nand U6710 (N_6710,N_6382,N_6359);
xor U6711 (N_6711,N_6534,N_6564);
xor U6712 (N_6712,N_6353,N_6512);
or U6713 (N_6713,N_6593,N_6348);
nor U6714 (N_6714,N_6591,N_6488);
xor U6715 (N_6715,N_6341,N_6468);
nor U6716 (N_6716,N_6484,N_6518);
or U6717 (N_6717,N_6329,N_6364);
and U6718 (N_6718,N_6506,N_6482);
nand U6719 (N_6719,N_6428,N_6559);
xor U6720 (N_6720,N_6586,N_6384);
or U6721 (N_6721,N_6365,N_6318);
or U6722 (N_6722,N_6478,N_6370);
or U6723 (N_6723,N_6316,N_6379);
xor U6724 (N_6724,N_6368,N_6451);
nor U6725 (N_6725,N_6481,N_6367);
or U6726 (N_6726,N_6581,N_6502);
nor U6727 (N_6727,N_6393,N_6576);
and U6728 (N_6728,N_6402,N_6349);
and U6729 (N_6729,N_6452,N_6538);
nor U6730 (N_6730,N_6500,N_6560);
nand U6731 (N_6731,N_6531,N_6423);
nor U6732 (N_6732,N_6344,N_6514);
nor U6733 (N_6733,N_6419,N_6434);
xnor U6734 (N_6734,N_6433,N_6317);
xor U6735 (N_6735,N_6520,N_6466);
or U6736 (N_6736,N_6447,N_6585);
or U6737 (N_6737,N_6594,N_6392);
xnor U6738 (N_6738,N_6389,N_6599);
nor U6739 (N_6739,N_6533,N_6459);
or U6740 (N_6740,N_6573,N_6449);
nand U6741 (N_6741,N_6579,N_6495);
nor U6742 (N_6742,N_6414,N_6540);
and U6743 (N_6743,N_6310,N_6547);
or U6744 (N_6744,N_6380,N_6408);
and U6745 (N_6745,N_6552,N_6521);
xnor U6746 (N_6746,N_6421,N_6458);
nand U6747 (N_6747,N_6376,N_6313);
or U6748 (N_6748,N_6551,N_6412);
xnor U6749 (N_6749,N_6366,N_6340);
nor U6750 (N_6750,N_6335,N_6550);
and U6751 (N_6751,N_6493,N_6308);
and U6752 (N_6752,N_6587,N_6469);
and U6753 (N_6753,N_6426,N_6480);
xnor U6754 (N_6754,N_6484,N_6514);
nor U6755 (N_6755,N_6596,N_6312);
xnor U6756 (N_6756,N_6563,N_6559);
or U6757 (N_6757,N_6311,N_6321);
nor U6758 (N_6758,N_6487,N_6442);
xnor U6759 (N_6759,N_6311,N_6556);
or U6760 (N_6760,N_6510,N_6518);
and U6761 (N_6761,N_6397,N_6342);
and U6762 (N_6762,N_6318,N_6575);
xor U6763 (N_6763,N_6383,N_6514);
nand U6764 (N_6764,N_6457,N_6597);
nor U6765 (N_6765,N_6320,N_6479);
nor U6766 (N_6766,N_6375,N_6569);
xnor U6767 (N_6767,N_6467,N_6596);
xor U6768 (N_6768,N_6595,N_6533);
nor U6769 (N_6769,N_6478,N_6320);
nor U6770 (N_6770,N_6312,N_6483);
nand U6771 (N_6771,N_6544,N_6406);
and U6772 (N_6772,N_6453,N_6514);
xor U6773 (N_6773,N_6480,N_6405);
nor U6774 (N_6774,N_6399,N_6311);
xnor U6775 (N_6775,N_6533,N_6598);
xnor U6776 (N_6776,N_6587,N_6306);
or U6777 (N_6777,N_6550,N_6388);
and U6778 (N_6778,N_6465,N_6502);
nor U6779 (N_6779,N_6507,N_6418);
and U6780 (N_6780,N_6305,N_6439);
nand U6781 (N_6781,N_6519,N_6373);
nor U6782 (N_6782,N_6561,N_6399);
nand U6783 (N_6783,N_6496,N_6529);
nor U6784 (N_6784,N_6517,N_6509);
nor U6785 (N_6785,N_6548,N_6340);
and U6786 (N_6786,N_6302,N_6451);
or U6787 (N_6787,N_6446,N_6529);
or U6788 (N_6788,N_6417,N_6427);
xor U6789 (N_6789,N_6357,N_6474);
nand U6790 (N_6790,N_6492,N_6529);
nor U6791 (N_6791,N_6542,N_6561);
or U6792 (N_6792,N_6488,N_6549);
xor U6793 (N_6793,N_6329,N_6358);
and U6794 (N_6794,N_6330,N_6342);
nand U6795 (N_6795,N_6575,N_6343);
nor U6796 (N_6796,N_6555,N_6493);
xor U6797 (N_6797,N_6467,N_6415);
or U6798 (N_6798,N_6441,N_6333);
or U6799 (N_6799,N_6514,N_6465);
nand U6800 (N_6800,N_6363,N_6376);
nor U6801 (N_6801,N_6582,N_6536);
and U6802 (N_6802,N_6413,N_6386);
or U6803 (N_6803,N_6487,N_6510);
xor U6804 (N_6804,N_6589,N_6505);
and U6805 (N_6805,N_6531,N_6511);
nand U6806 (N_6806,N_6386,N_6587);
or U6807 (N_6807,N_6534,N_6399);
nor U6808 (N_6808,N_6530,N_6373);
and U6809 (N_6809,N_6501,N_6560);
nor U6810 (N_6810,N_6462,N_6536);
or U6811 (N_6811,N_6358,N_6315);
nor U6812 (N_6812,N_6457,N_6456);
nor U6813 (N_6813,N_6582,N_6498);
or U6814 (N_6814,N_6563,N_6362);
nand U6815 (N_6815,N_6329,N_6311);
and U6816 (N_6816,N_6576,N_6586);
nand U6817 (N_6817,N_6473,N_6371);
or U6818 (N_6818,N_6374,N_6427);
or U6819 (N_6819,N_6552,N_6583);
and U6820 (N_6820,N_6507,N_6408);
xor U6821 (N_6821,N_6395,N_6397);
or U6822 (N_6822,N_6466,N_6329);
nor U6823 (N_6823,N_6557,N_6511);
nand U6824 (N_6824,N_6562,N_6363);
and U6825 (N_6825,N_6357,N_6521);
or U6826 (N_6826,N_6567,N_6358);
or U6827 (N_6827,N_6365,N_6439);
nand U6828 (N_6828,N_6523,N_6559);
or U6829 (N_6829,N_6504,N_6583);
xor U6830 (N_6830,N_6499,N_6305);
nor U6831 (N_6831,N_6442,N_6466);
or U6832 (N_6832,N_6527,N_6549);
nand U6833 (N_6833,N_6427,N_6401);
or U6834 (N_6834,N_6331,N_6487);
nor U6835 (N_6835,N_6514,N_6593);
xor U6836 (N_6836,N_6520,N_6526);
and U6837 (N_6837,N_6432,N_6308);
or U6838 (N_6838,N_6535,N_6345);
nor U6839 (N_6839,N_6448,N_6315);
or U6840 (N_6840,N_6416,N_6516);
and U6841 (N_6841,N_6590,N_6542);
or U6842 (N_6842,N_6387,N_6469);
and U6843 (N_6843,N_6579,N_6361);
xnor U6844 (N_6844,N_6477,N_6454);
nor U6845 (N_6845,N_6312,N_6328);
xnor U6846 (N_6846,N_6307,N_6444);
or U6847 (N_6847,N_6403,N_6481);
or U6848 (N_6848,N_6413,N_6542);
nand U6849 (N_6849,N_6513,N_6531);
nor U6850 (N_6850,N_6563,N_6500);
or U6851 (N_6851,N_6546,N_6586);
and U6852 (N_6852,N_6413,N_6543);
and U6853 (N_6853,N_6383,N_6452);
or U6854 (N_6854,N_6430,N_6537);
nand U6855 (N_6855,N_6411,N_6457);
nand U6856 (N_6856,N_6525,N_6569);
nor U6857 (N_6857,N_6490,N_6387);
nand U6858 (N_6858,N_6467,N_6497);
nor U6859 (N_6859,N_6528,N_6519);
or U6860 (N_6860,N_6587,N_6405);
xnor U6861 (N_6861,N_6319,N_6498);
nand U6862 (N_6862,N_6389,N_6321);
or U6863 (N_6863,N_6386,N_6531);
nand U6864 (N_6864,N_6531,N_6584);
nor U6865 (N_6865,N_6313,N_6412);
nand U6866 (N_6866,N_6361,N_6518);
nor U6867 (N_6867,N_6322,N_6435);
xnor U6868 (N_6868,N_6533,N_6396);
or U6869 (N_6869,N_6509,N_6373);
and U6870 (N_6870,N_6531,N_6433);
or U6871 (N_6871,N_6475,N_6336);
or U6872 (N_6872,N_6518,N_6590);
or U6873 (N_6873,N_6461,N_6527);
xor U6874 (N_6874,N_6577,N_6387);
xor U6875 (N_6875,N_6439,N_6335);
or U6876 (N_6876,N_6570,N_6584);
nand U6877 (N_6877,N_6352,N_6551);
xor U6878 (N_6878,N_6576,N_6336);
nor U6879 (N_6879,N_6381,N_6308);
or U6880 (N_6880,N_6367,N_6466);
nand U6881 (N_6881,N_6596,N_6363);
xor U6882 (N_6882,N_6328,N_6434);
or U6883 (N_6883,N_6583,N_6536);
nand U6884 (N_6884,N_6528,N_6386);
and U6885 (N_6885,N_6447,N_6338);
or U6886 (N_6886,N_6373,N_6366);
nor U6887 (N_6887,N_6372,N_6446);
or U6888 (N_6888,N_6322,N_6461);
nor U6889 (N_6889,N_6441,N_6543);
and U6890 (N_6890,N_6570,N_6414);
nand U6891 (N_6891,N_6397,N_6385);
xnor U6892 (N_6892,N_6485,N_6439);
nand U6893 (N_6893,N_6427,N_6534);
xor U6894 (N_6894,N_6577,N_6369);
xnor U6895 (N_6895,N_6329,N_6552);
xnor U6896 (N_6896,N_6322,N_6421);
xor U6897 (N_6897,N_6355,N_6374);
nand U6898 (N_6898,N_6537,N_6492);
nor U6899 (N_6899,N_6450,N_6492);
nand U6900 (N_6900,N_6651,N_6698);
and U6901 (N_6901,N_6782,N_6646);
xnor U6902 (N_6902,N_6826,N_6627);
xnor U6903 (N_6903,N_6787,N_6893);
and U6904 (N_6904,N_6885,N_6899);
or U6905 (N_6905,N_6623,N_6809);
and U6906 (N_6906,N_6880,N_6762);
and U6907 (N_6907,N_6648,N_6664);
and U6908 (N_6908,N_6682,N_6850);
nor U6909 (N_6909,N_6833,N_6712);
xor U6910 (N_6910,N_6605,N_6621);
xor U6911 (N_6911,N_6796,N_6754);
xnor U6912 (N_6912,N_6635,N_6875);
nor U6913 (N_6913,N_6720,N_6670);
nor U6914 (N_6914,N_6843,N_6683);
nor U6915 (N_6915,N_6853,N_6625);
and U6916 (N_6916,N_6748,N_6751);
or U6917 (N_6917,N_6849,N_6689);
or U6918 (N_6918,N_6806,N_6614);
nand U6919 (N_6919,N_6765,N_6821);
xor U6920 (N_6920,N_6679,N_6858);
xnor U6921 (N_6921,N_6700,N_6788);
nand U6922 (N_6922,N_6672,N_6804);
nand U6923 (N_6923,N_6737,N_6686);
nand U6924 (N_6924,N_6791,N_6823);
nor U6925 (N_6925,N_6608,N_6793);
nor U6926 (N_6926,N_6871,N_6836);
or U6927 (N_6927,N_6705,N_6638);
nand U6928 (N_6928,N_6717,N_6668);
nor U6929 (N_6929,N_6667,N_6839);
xor U6930 (N_6930,N_6845,N_6766);
nor U6931 (N_6931,N_6786,N_6852);
xnor U6932 (N_6932,N_6855,N_6758);
nand U6933 (N_6933,N_6657,N_6719);
xnor U6934 (N_6934,N_6835,N_6632);
nor U6935 (N_6935,N_6602,N_6652);
xnor U6936 (N_6936,N_6863,N_6760);
and U6937 (N_6937,N_6897,N_6798);
nand U6938 (N_6938,N_6726,N_6781);
nor U6939 (N_6939,N_6661,N_6671);
nand U6940 (N_6940,N_6862,N_6879);
and U6941 (N_6941,N_6660,N_6658);
and U6942 (N_6942,N_6663,N_6889);
nor U6943 (N_6943,N_6868,N_6644);
nor U6944 (N_6944,N_6801,N_6730);
nand U6945 (N_6945,N_6831,N_6817);
xor U6946 (N_6946,N_6736,N_6763);
nand U6947 (N_6947,N_6629,N_6709);
nor U6948 (N_6948,N_6755,N_6691);
xnor U6949 (N_6949,N_6636,N_6721);
nand U6950 (N_6950,N_6764,N_6684);
or U6951 (N_6951,N_6693,N_6674);
xnor U6952 (N_6952,N_6840,N_6878);
and U6953 (N_6953,N_6659,N_6807);
and U6954 (N_6954,N_6738,N_6877);
nor U6955 (N_6955,N_6665,N_6703);
nor U6956 (N_6956,N_6825,N_6723);
or U6957 (N_6957,N_6779,N_6708);
xor U6958 (N_6958,N_6681,N_6799);
xor U6959 (N_6959,N_6851,N_6733);
nor U6960 (N_6960,N_6604,N_6626);
xor U6961 (N_6961,N_6860,N_6800);
nor U6962 (N_6962,N_6677,N_6607);
or U6963 (N_6963,N_6750,N_6829);
and U6964 (N_6964,N_6856,N_6669);
xnor U6965 (N_6965,N_6715,N_6746);
and U6966 (N_6966,N_6805,N_6848);
or U6967 (N_6967,N_6624,N_6713);
nor U6968 (N_6968,N_6729,N_6847);
nor U6969 (N_6969,N_6743,N_6797);
nand U6970 (N_6970,N_6768,N_6811);
nor U6971 (N_6971,N_6702,N_6859);
nand U6972 (N_6972,N_6710,N_6609);
or U6973 (N_6973,N_6892,N_6774);
nor U6974 (N_6974,N_6706,N_6718);
or U6975 (N_6975,N_6615,N_6767);
and U6976 (N_6976,N_6647,N_6864);
and U6977 (N_6977,N_6611,N_6891);
nor U6978 (N_6978,N_6610,N_6676);
and U6979 (N_6979,N_6612,N_6832);
nor U6980 (N_6980,N_6639,N_6601);
nor U6981 (N_6981,N_6704,N_6634);
nand U6982 (N_6982,N_6792,N_6789);
nand U6983 (N_6983,N_6742,N_6687);
nor U6984 (N_6984,N_6716,N_6830);
or U6985 (N_6985,N_6645,N_6620);
and U6986 (N_6986,N_6769,N_6673);
nand U6987 (N_6987,N_6735,N_6756);
nor U6988 (N_6988,N_6841,N_6834);
and U6989 (N_6989,N_6606,N_6739);
xnor U6990 (N_6990,N_6633,N_6641);
or U6991 (N_6991,N_6816,N_6642);
xnor U6992 (N_6992,N_6753,N_6790);
nand U6993 (N_6993,N_6881,N_6828);
nand U6994 (N_6994,N_6622,N_6744);
nor U6995 (N_6995,N_6740,N_6895);
or U6996 (N_6996,N_6745,N_6867);
or U6997 (N_6997,N_6749,N_6697);
or U6998 (N_6998,N_6694,N_6678);
or U6999 (N_6999,N_6894,N_6810);
nand U7000 (N_7000,N_6780,N_6656);
nor U7001 (N_7001,N_6775,N_6643);
xnor U7002 (N_7002,N_6898,N_6613);
or U7003 (N_7003,N_6603,N_6795);
nor U7004 (N_7004,N_6822,N_6776);
or U7005 (N_7005,N_6616,N_6752);
xnor U7006 (N_7006,N_6734,N_6890);
xnor U7007 (N_7007,N_6820,N_6874);
nor U7008 (N_7008,N_6653,N_6630);
nor U7009 (N_7009,N_6772,N_6887);
nor U7010 (N_7010,N_6619,N_6777);
nor U7011 (N_7011,N_6770,N_6888);
and U7012 (N_7012,N_6650,N_6814);
nand U7013 (N_7013,N_6649,N_6844);
xnor U7014 (N_7014,N_6675,N_6838);
xnor U7015 (N_7015,N_6662,N_6866);
xnor U7016 (N_7016,N_6773,N_6728);
and U7017 (N_7017,N_6883,N_6618);
xnor U7018 (N_7018,N_6815,N_6696);
nand U7019 (N_7019,N_6732,N_6690);
or U7020 (N_7020,N_6783,N_6600);
or U7021 (N_7021,N_6876,N_6695);
nor U7022 (N_7022,N_6707,N_6640);
nand U7023 (N_7023,N_6692,N_6784);
or U7024 (N_7024,N_6631,N_6680);
xnor U7025 (N_7025,N_6688,N_6761);
nor U7026 (N_7026,N_6873,N_6785);
or U7027 (N_7027,N_6699,N_6655);
nor U7028 (N_7028,N_6727,N_6884);
xor U7029 (N_7029,N_6869,N_6827);
or U7030 (N_7030,N_6725,N_6818);
or U7031 (N_7031,N_6714,N_6637);
and U7032 (N_7032,N_6813,N_6794);
nor U7033 (N_7033,N_6628,N_6731);
xor U7034 (N_7034,N_6803,N_6846);
nand U7035 (N_7035,N_6808,N_6617);
and U7036 (N_7036,N_6865,N_6842);
xor U7037 (N_7037,N_6870,N_6857);
xor U7038 (N_7038,N_6757,N_6711);
nor U7039 (N_7039,N_6819,N_6861);
or U7040 (N_7040,N_6896,N_6654);
nor U7041 (N_7041,N_6701,N_6872);
and U7042 (N_7042,N_6722,N_6882);
or U7043 (N_7043,N_6724,N_6854);
xnor U7044 (N_7044,N_6771,N_6824);
xor U7045 (N_7045,N_6685,N_6747);
nand U7046 (N_7046,N_6759,N_6666);
nor U7047 (N_7047,N_6802,N_6886);
nand U7048 (N_7048,N_6778,N_6812);
or U7049 (N_7049,N_6741,N_6837);
nand U7050 (N_7050,N_6892,N_6698);
xor U7051 (N_7051,N_6683,N_6887);
xor U7052 (N_7052,N_6859,N_6637);
and U7053 (N_7053,N_6720,N_6652);
or U7054 (N_7054,N_6836,N_6822);
xnor U7055 (N_7055,N_6625,N_6650);
nand U7056 (N_7056,N_6625,N_6813);
nor U7057 (N_7057,N_6879,N_6660);
or U7058 (N_7058,N_6779,N_6658);
nand U7059 (N_7059,N_6820,N_6802);
nand U7060 (N_7060,N_6673,N_6789);
nand U7061 (N_7061,N_6766,N_6881);
xnor U7062 (N_7062,N_6744,N_6705);
and U7063 (N_7063,N_6844,N_6837);
xor U7064 (N_7064,N_6709,N_6702);
xnor U7065 (N_7065,N_6877,N_6891);
xor U7066 (N_7066,N_6715,N_6826);
or U7067 (N_7067,N_6860,N_6782);
nor U7068 (N_7068,N_6713,N_6871);
nor U7069 (N_7069,N_6639,N_6672);
and U7070 (N_7070,N_6618,N_6821);
nand U7071 (N_7071,N_6766,N_6700);
nor U7072 (N_7072,N_6704,N_6690);
nand U7073 (N_7073,N_6739,N_6690);
nor U7074 (N_7074,N_6892,N_6621);
nor U7075 (N_7075,N_6807,N_6610);
nand U7076 (N_7076,N_6722,N_6836);
xor U7077 (N_7077,N_6771,N_6649);
or U7078 (N_7078,N_6806,N_6685);
xor U7079 (N_7079,N_6650,N_6825);
or U7080 (N_7080,N_6742,N_6624);
and U7081 (N_7081,N_6811,N_6641);
or U7082 (N_7082,N_6690,N_6654);
nand U7083 (N_7083,N_6656,N_6814);
nor U7084 (N_7084,N_6804,N_6770);
nand U7085 (N_7085,N_6895,N_6756);
or U7086 (N_7086,N_6673,N_6767);
nand U7087 (N_7087,N_6651,N_6679);
nor U7088 (N_7088,N_6822,N_6813);
or U7089 (N_7089,N_6810,N_6847);
and U7090 (N_7090,N_6868,N_6717);
nand U7091 (N_7091,N_6679,N_6873);
xor U7092 (N_7092,N_6825,N_6703);
nor U7093 (N_7093,N_6788,N_6696);
nand U7094 (N_7094,N_6771,N_6655);
or U7095 (N_7095,N_6761,N_6693);
xnor U7096 (N_7096,N_6755,N_6787);
and U7097 (N_7097,N_6896,N_6851);
xnor U7098 (N_7098,N_6878,N_6784);
nor U7099 (N_7099,N_6818,N_6761);
nor U7100 (N_7100,N_6765,N_6695);
xnor U7101 (N_7101,N_6871,N_6809);
and U7102 (N_7102,N_6753,N_6679);
or U7103 (N_7103,N_6728,N_6700);
nand U7104 (N_7104,N_6705,N_6665);
or U7105 (N_7105,N_6600,N_6635);
nor U7106 (N_7106,N_6842,N_6612);
and U7107 (N_7107,N_6768,N_6795);
and U7108 (N_7108,N_6832,N_6714);
nor U7109 (N_7109,N_6635,N_6838);
nand U7110 (N_7110,N_6812,N_6746);
nand U7111 (N_7111,N_6880,N_6718);
nor U7112 (N_7112,N_6730,N_6739);
nand U7113 (N_7113,N_6766,N_6737);
xor U7114 (N_7114,N_6741,N_6740);
or U7115 (N_7115,N_6700,N_6630);
nor U7116 (N_7116,N_6733,N_6842);
and U7117 (N_7117,N_6600,N_6794);
nor U7118 (N_7118,N_6697,N_6885);
or U7119 (N_7119,N_6695,N_6758);
or U7120 (N_7120,N_6634,N_6806);
or U7121 (N_7121,N_6678,N_6875);
nand U7122 (N_7122,N_6646,N_6705);
nor U7123 (N_7123,N_6694,N_6887);
nand U7124 (N_7124,N_6765,N_6863);
and U7125 (N_7125,N_6696,N_6600);
or U7126 (N_7126,N_6834,N_6828);
xnor U7127 (N_7127,N_6626,N_6759);
nand U7128 (N_7128,N_6785,N_6802);
and U7129 (N_7129,N_6796,N_6729);
nor U7130 (N_7130,N_6892,N_6792);
xor U7131 (N_7131,N_6823,N_6887);
nand U7132 (N_7132,N_6678,N_6715);
and U7133 (N_7133,N_6734,N_6675);
and U7134 (N_7134,N_6635,N_6750);
nand U7135 (N_7135,N_6691,N_6783);
and U7136 (N_7136,N_6853,N_6623);
and U7137 (N_7137,N_6601,N_6756);
nor U7138 (N_7138,N_6679,N_6752);
and U7139 (N_7139,N_6622,N_6676);
nand U7140 (N_7140,N_6864,N_6645);
xor U7141 (N_7141,N_6754,N_6806);
xor U7142 (N_7142,N_6800,N_6632);
xnor U7143 (N_7143,N_6635,N_6727);
nand U7144 (N_7144,N_6806,N_6788);
and U7145 (N_7145,N_6678,N_6848);
and U7146 (N_7146,N_6868,N_6846);
and U7147 (N_7147,N_6819,N_6754);
or U7148 (N_7148,N_6814,N_6880);
nand U7149 (N_7149,N_6856,N_6663);
and U7150 (N_7150,N_6832,N_6819);
xor U7151 (N_7151,N_6884,N_6823);
or U7152 (N_7152,N_6624,N_6787);
nand U7153 (N_7153,N_6815,N_6755);
nor U7154 (N_7154,N_6829,N_6691);
nand U7155 (N_7155,N_6744,N_6707);
xor U7156 (N_7156,N_6673,N_6827);
or U7157 (N_7157,N_6838,N_6757);
nand U7158 (N_7158,N_6852,N_6875);
and U7159 (N_7159,N_6601,N_6613);
nand U7160 (N_7160,N_6663,N_6659);
or U7161 (N_7161,N_6718,N_6789);
xnor U7162 (N_7162,N_6822,N_6864);
or U7163 (N_7163,N_6782,N_6712);
xor U7164 (N_7164,N_6883,N_6794);
xor U7165 (N_7165,N_6748,N_6774);
xor U7166 (N_7166,N_6614,N_6768);
nand U7167 (N_7167,N_6850,N_6698);
nor U7168 (N_7168,N_6608,N_6738);
xor U7169 (N_7169,N_6632,N_6648);
nor U7170 (N_7170,N_6776,N_6896);
nor U7171 (N_7171,N_6872,N_6602);
nand U7172 (N_7172,N_6750,N_6857);
and U7173 (N_7173,N_6878,N_6747);
xnor U7174 (N_7174,N_6640,N_6755);
or U7175 (N_7175,N_6895,N_6649);
and U7176 (N_7176,N_6624,N_6829);
and U7177 (N_7177,N_6678,N_6847);
nor U7178 (N_7178,N_6667,N_6868);
or U7179 (N_7179,N_6747,N_6724);
nor U7180 (N_7180,N_6843,N_6781);
nor U7181 (N_7181,N_6606,N_6832);
or U7182 (N_7182,N_6763,N_6878);
or U7183 (N_7183,N_6851,N_6721);
and U7184 (N_7184,N_6802,N_6896);
nand U7185 (N_7185,N_6749,N_6683);
and U7186 (N_7186,N_6780,N_6633);
nand U7187 (N_7187,N_6833,N_6891);
nand U7188 (N_7188,N_6818,N_6617);
and U7189 (N_7189,N_6674,N_6850);
nand U7190 (N_7190,N_6679,N_6884);
nor U7191 (N_7191,N_6890,N_6761);
or U7192 (N_7192,N_6806,N_6822);
nor U7193 (N_7193,N_6794,N_6627);
or U7194 (N_7194,N_6770,N_6825);
nand U7195 (N_7195,N_6812,N_6855);
and U7196 (N_7196,N_6711,N_6631);
or U7197 (N_7197,N_6881,N_6680);
xor U7198 (N_7198,N_6754,N_6601);
or U7199 (N_7199,N_6835,N_6821);
xnor U7200 (N_7200,N_7029,N_7148);
or U7201 (N_7201,N_7014,N_7074);
and U7202 (N_7202,N_6915,N_6936);
or U7203 (N_7203,N_6932,N_6954);
nor U7204 (N_7204,N_7159,N_6947);
xor U7205 (N_7205,N_7089,N_7067);
xor U7206 (N_7206,N_6982,N_6996);
and U7207 (N_7207,N_7174,N_6907);
or U7208 (N_7208,N_7168,N_6906);
xor U7209 (N_7209,N_7183,N_7017);
or U7210 (N_7210,N_7035,N_7006);
and U7211 (N_7211,N_6938,N_7123);
nor U7212 (N_7212,N_6918,N_7151);
xor U7213 (N_7213,N_7090,N_7152);
nand U7214 (N_7214,N_7186,N_7120);
nor U7215 (N_7215,N_6998,N_6973);
and U7216 (N_7216,N_7030,N_7107);
nor U7217 (N_7217,N_7114,N_7110);
xnor U7218 (N_7218,N_7113,N_7109);
or U7219 (N_7219,N_6997,N_7082);
or U7220 (N_7220,N_7003,N_6976);
and U7221 (N_7221,N_6922,N_6925);
xor U7222 (N_7222,N_7160,N_6916);
nand U7223 (N_7223,N_6960,N_7095);
or U7224 (N_7224,N_6924,N_6985);
xor U7225 (N_7225,N_7078,N_7004);
xor U7226 (N_7226,N_7162,N_7194);
and U7227 (N_7227,N_7102,N_7116);
nand U7228 (N_7228,N_7064,N_7119);
or U7229 (N_7229,N_7138,N_6902);
or U7230 (N_7230,N_7139,N_6931);
nand U7231 (N_7231,N_7104,N_7173);
nor U7232 (N_7232,N_7187,N_7199);
nor U7233 (N_7233,N_7052,N_7143);
nor U7234 (N_7234,N_7031,N_7028);
xor U7235 (N_7235,N_6991,N_7141);
or U7236 (N_7236,N_6959,N_7103);
xnor U7237 (N_7237,N_7177,N_7079);
nand U7238 (N_7238,N_6964,N_6937);
nand U7239 (N_7239,N_6983,N_7026);
or U7240 (N_7240,N_6957,N_7125);
nor U7241 (N_7241,N_7190,N_7001);
or U7242 (N_7242,N_7155,N_6928);
nand U7243 (N_7243,N_7092,N_7038);
xnor U7244 (N_7244,N_7072,N_7080);
nor U7245 (N_7245,N_6980,N_7053);
or U7246 (N_7246,N_6999,N_7022);
nor U7247 (N_7247,N_7009,N_7045);
nand U7248 (N_7248,N_7179,N_6934);
or U7249 (N_7249,N_7037,N_7083);
nand U7250 (N_7250,N_6940,N_6903);
nor U7251 (N_7251,N_6988,N_7158);
and U7252 (N_7252,N_7129,N_7135);
nor U7253 (N_7253,N_7112,N_7044);
xor U7254 (N_7254,N_6939,N_7153);
nor U7255 (N_7255,N_6910,N_7002);
nor U7256 (N_7256,N_7065,N_7097);
xnor U7257 (N_7257,N_7171,N_7066);
and U7258 (N_7258,N_6901,N_6953);
xor U7259 (N_7259,N_7147,N_7070);
nor U7260 (N_7260,N_6917,N_7106);
nand U7261 (N_7261,N_7164,N_7108);
nand U7262 (N_7262,N_7005,N_7087);
or U7263 (N_7263,N_7027,N_7197);
or U7264 (N_7264,N_7099,N_7051);
nand U7265 (N_7265,N_7055,N_6984);
or U7266 (N_7266,N_7161,N_7165);
or U7267 (N_7267,N_7011,N_7069);
xnor U7268 (N_7268,N_6927,N_7166);
nor U7269 (N_7269,N_7034,N_6944);
xnor U7270 (N_7270,N_6965,N_7189);
nor U7271 (N_7271,N_7073,N_7100);
nand U7272 (N_7272,N_7071,N_6900);
nand U7273 (N_7273,N_7145,N_7056);
xnor U7274 (N_7274,N_7157,N_6970);
or U7275 (N_7275,N_6987,N_7008);
or U7276 (N_7276,N_7000,N_7131);
nand U7277 (N_7277,N_6955,N_7185);
nor U7278 (N_7278,N_7054,N_6911);
and U7279 (N_7279,N_6942,N_7101);
xnor U7280 (N_7280,N_7192,N_7117);
or U7281 (N_7281,N_6920,N_7061);
xor U7282 (N_7282,N_7188,N_6951);
xnor U7283 (N_7283,N_7060,N_7196);
or U7284 (N_7284,N_7012,N_7091);
xor U7285 (N_7285,N_7178,N_6956);
or U7286 (N_7286,N_6990,N_7010);
or U7287 (N_7287,N_6914,N_7016);
and U7288 (N_7288,N_6923,N_7133);
and U7289 (N_7289,N_6930,N_6993);
xnor U7290 (N_7290,N_7059,N_7163);
xnor U7291 (N_7291,N_7094,N_6929);
nand U7292 (N_7292,N_7140,N_6945);
xor U7293 (N_7293,N_7023,N_7181);
xnor U7294 (N_7294,N_6967,N_7118);
nor U7295 (N_7295,N_7042,N_7093);
xor U7296 (N_7296,N_7062,N_6994);
nor U7297 (N_7297,N_7046,N_6943);
xor U7298 (N_7298,N_7024,N_7020);
and U7299 (N_7299,N_6968,N_6913);
nor U7300 (N_7300,N_7050,N_7124);
nor U7301 (N_7301,N_7182,N_7191);
xnor U7302 (N_7302,N_7085,N_7036);
and U7303 (N_7303,N_7057,N_6908);
or U7304 (N_7304,N_7176,N_7098);
xor U7305 (N_7305,N_7105,N_7115);
nand U7306 (N_7306,N_7047,N_7063);
or U7307 (N_7307,N_6981,N_7040);
and U7308 (N_7308,N_6933,N_6952);
and U7309 (N_7309,N_6926,N_6949);
and U7310 (N_7310,N_6989,N_7167);
nand U7311 (N_7311,N_7175,N_7128);
or U7312 (N_7312,N_7043,N_7142);
or U7313 (N_7313,N_7033,N_6975);
nand U7314 (N_7314,N_6966,N_7137);
xor U7315 (N_7315,N_7172,N_6978);
nand U7316 (N_7316,N_6979,N_7013);
xor U7317 (N_7317,N_6977,N_7111);
and U7318 (N_7318,N_7058,N_7088);
nor U7319 (N_7319,N_6904,N_7015);
and U7320 (N_7320,N_7198,N_7049);
and U7321 (N_7321,N_6921,N_7048);
nand U7322 (N_7322,N_6905,N_7041);
nand U7323 (N_7323,N_7149,N_7130);
xnor U7324 (N_7324,N_7121,N_7025);
nor U7325 (N_7325,N_7077,N_6992);
or U7326 (N_7326,N_6950,N_6969);
xnor U7327 (N_7327,N_6919,N_6958);
nor U7328 (N_7328,N_7193,N_7180);
nand U7329 (N_7329,N_7146,N_7154);
xnor U7330 (N_7330,N_7081,N_7134);
nor U7331 (N_7331,N_7122,N_7169);
nor U7332 (N_7332,N_7126,N_7068);
nor U7333 (N_7333,N_7039,N_6971);
nand U7334 (N_7334,N_7144,N_7156);
nor U7335 (N_7335,N_7018,N_6963);
and U7336 (N_7336,N_6946,N_6941);
nor U7337 (N_7337,N_7195,N_7150);
nor U7338 (N_7338,N_7086,N_6961);
nand U7339 (N_7339,N_7075,N_6995);
nand U7340 (N_7340,N_6912,N_7136);
nor U7341 (N_7341,N_7007,N_7127);
and U7342 (N_7342,N_7076,N_7019);
nand U7343 (N_7343,N_7170,N_6962);
nor U7344 (N_7344,N_7132,N_7084);
xor U7345 (N_7345,N_6948,N_7021);
nand U7346 (N_7346,N_7032,N_6935);
and U7347 (N_7347,N_6974,N_7096);
or U7348 (N_7348,N_6986,N_7184);
xnor U7349 (N_7349,N_6972,N_6909);
nand U7350 (N_7350,N_6946,N_6963);
and U7351 (N_7351,N_7093,N_7075);
nand U7352 (N_7352,N_7192,N_7025);
nor U7353 (N_7353,N_6922,N_7152);
or U7354 (N_7354,N_7091,N_6916);
or U7355 (N_7355,N_7041,N_6904);
nor U7356 (N_7356,N_7031,N_6935);
nand U7357 (N_7357,N_6930,N_6999);
nor U7358 (N_7358,N_7047,N_7022);
nor U7359 (N_7359,N_7045,N_7019);
nand U7360 (N_7360,N_7058,N_7011);
nor U7361 (N_7361,N_7129,N_7053);
or U7362 (N_7362,N_7001,N_7096);
xnor U7363 (N_7363,N_7037,N_7084);
nand U7364 (N_7364,N_7048,N_7066);
nor U7365 (N_7365,N_7025,N_7164);
nand U7366 (N_7366,N_7113,N_7038);
and U7367 (N_7367,N_7108,N_7113);
nor U7368 (N_7368,N_6916,N_6918);
nor U7369 (N_7369,N_6961,N_7134);
or U7370 (N_7370,N_6956,N_6992);
nand U7371 (N_7371,N_7126,N_7089);
and U7372 (N_7372,N_6949,N_7050);
and U7373 (N_7373,N_7188,N_7041);
nand U7374 (N_7374,N_6985,N_7171);
or U7375 (N_7375,N_7046,N_6908);
nor U7376 (N_7376,N_7180,N_7119);
xnor U7377 (N_7377,N_7105,N_7194);
nor U7378 (N_7378,N_7168,N_7118);
xor U7379 (N_7379,N_7027,N_6978);
xor U7380 (N_7380,N_7069,N_7054);
and U7381 (N_7381,N_7022,N_6948);
nand U7382 (N_7382,N_7148,N_7198);
nor U7383 (N_7383,N_7126,N_7029);
and U7384 (N_7384,N_6931,N_7018);
xor U7385 (N_7385,N_7104,N_6906);
and U7386 (N_7386,N_7013,N_7043);
nor U7387 (N_7387,N_7012,N_7003);
and U7388 (N_7388,N_7050,N_6916);
nor U7389 (N_7389,N_7162,N_7064);
and U7390 (N_7390,N_7134,N_7176);
and U7391 (N_7391,N_7076,N_7098);
xor U7392 (N_7392,N_7069,N_7152);
nand U7393 (N_7393,N_7127,N_6955);
xor U7394 (N_7394,N_7060,N_6938);
xor U7395 (N_7395,N_6987,N_7104);
nor U7396 (N_7396,N_7039,N_6932);
or U7397 (N_7397,N_6968,N_6907);
nand U7398 (N_7398,N_7057,N_7126);
nor U7399 (N_7399,N_7199,N_7051);
nand U7400 (N_7400,N_7011,N_7020);
or U7401 (N_7401,N_6944,N_7015);
xnor U7402 (N_7402,N_7157,N_7187);
or U7403 (N_7403,N_7116,N_7008);
or U7404 (N_7404,N_7075,N_7085);
and U7405 (N_7405,N_7105,N_7172);
xor U7406 (N_7406,N_7093,N_7153);
or U7407 (N_7407,N_7064,N_6903);
nor U7408 (N_7408,N_6939,N_7088);
or U7409 (N_7409,N_6938,N_7046);
and U7410 (N_7410,N_7037,N_7036);
and U7411 (N_7411,N_7150,N_6972);
nand U7412 (N_7412,N_6957,N_6946);
nand U7413 (N_7413,N_7192,N_6925);
xor U7414 (N_7414,N_7060,N_6998);
nand U7415 (N_7415,N_7038,N_6939);
xor U7416 (N_7416,N_7157,N_7138);
nor U7417 (N_7417,N_7031,N_7021);
or U7418 (N_7418,N_6976,N_7061);
nor U7419 (N_7419,N_7160,N_7069);
nor U7420 (N_7420,N_6995,N_7077);
and U7421 (N_7421,N_6973,N_6919);
nand U7422 (N_7422,N_7007,N_7023);
nand U7423 (N_7423,N_7100,N_7163);
and U7424 (N_7424,N_7066,N_7122);
xor U7425 (N_7425,N_6969,N_7103);
and U7426 (N_7426,N_7016,N_7130);
nand U7427 (N_7427,N_7196,N_7122);
nand U7428 (N_7428,N_6959,N_6934);
xor U7429 (N_7429,N_6955,N_6911);
nor U7430 (N_7430,N_7084,N_7098);
xnor U7431 (N_7431,N_7031,N_6922);
xnor U7432 (N_7432,N_7155,N_7045);
or U7433 (N_7433,N_7011,N_7176);
nor U7434 (N_7434,N_6930,N_7150);
or U7435 (N_7435,N_7149,N_6943);
xnor U7436 (N_7436,N_6960,N_7002);
nand U7437 (N_7437,N_7044,N_6968);
or U7438 (N_7438,N_7002,N_7057);
xor U7439 (N_7439,N_6996,N_7092);
xor U7440 (N_7440,N_6999,N_7039);
xnor U7441 (N_7441,N_7000,N_7167);
nor U7442 (N_7442,N_7091,N_6925);
nor U7443 (N_7443,N_7102,N_7197);
xor U7444 (N_7444,N_6932,N_7075);
nor U7445 (N_7445,N_6970,N_7018);
xnor U7446 (N_7446,N_6996,N_7107);
or U7447 (N_7447,N_6988,N_6987);
nand U7448 (N_7448,N_7074,N_7100);
nand U7449 (N_7449,N_6916,N_7135);
xnor U7450 (N_7450,N_7080,N_6966);
nand U7451 (N_7451,N_6938,N_7192);
nand U7452 (N_7452,N_6948,N_6993);
nor U7453 (N_7453,N_7171,N_7134);
and U7454 (N_7454,N_7167,N_7014);
xor U7455 (N_7455,N_6931,N_6902);
and U7456 (N_7456,N_7030,N_7046);
nor U7457 (N_7457,N_7113,N_6963);
and U7458 (N_7458,N_7193,N_7062);
xnor U7459 (N_7459,N_7187,N_7130);
nor U7460 (N_7460,N_6994,N_7146);
nand U7461 (N_7461,N_7104,N_7066);
xor U7462 (N_7462,N_7134,N_7083);
xor U7463 (N_7463,N_7170,N_7140);
nor U7464 (N_7464,N_6934,N_7160);
and U7465 (N_7465,N_6986,N_7071);
nand U7466 (N_7466,N_7020,N_7197);
xor U7467 (N_7467,N_7111,N_7114);
nor U7468 (N_7468,N_7073,N_7034);
nand U7469 (N_7469,N_7182,N_6957);
or U7470 (N_7470,N_7023,N_7070);
nor U7471 (N_7471,N_6945,N_7114);
and U7472 (N_7472,N_7178,N_6925);
and U7473 (N_7473,N_7174,N_7118);
nand U7474 (N_7474,N_7184,N_7110);
nor U7475 (N_7475,N_6998,N_7011);
nand U7476 (N_7476,N_6917,N_7094);
and U7477 (N_7477,N_6985,N_6932);
or U7478 (N_7478,N_6950,N_7077);
xnor U7479 (N_7479,N_6903,N_6926);
xor U7480 (N_7480,N_7114,N_7053);
nand U7481 (N_7481,N_7091,N_6938);
or U7482 (N_7482,N_7164,N_7031);
nor U7483 (N_7483,N_7106,N_7044);
and U7484 (N_7484,N_6933,N_7069);
or U7485 (N_7485,N_7168,N_7177);
nor U7486 (N_7486,N_7124,N_7048);
or U7487 (N_7487,N_7022,N_7028);
nand U7488 (N_7488,N_7046,N_6904);
nor U7489 (N_7489,N_6935,N_7108);
nor U7490 (N_7490,N_6995,N_7034);
nand U7491 (N_7491,N_6940,N_7192);
and U7492 (N_7492,N_6923,N_6936);
or U7493 (N_7493,N_7104,N_6953);
nor U7494 (N_7494,N_7026,N_7105);
or U7495 (N_7495,N_7034,N_7097);
nor U7496 (N_7496,N_7014,N_7083);
nand U7497 (N_7497,N_6985,N_7188);
xor U7498 (N_7498,N_6921,N_6950);
xnor U7499 (N_7499,N_7048,N_6918);
and U7500 (N_7500,N_7386,N_7452);
nand U7501 (N_7501,N_7205,N_7306);
and U7502 (N_7502,N_7322,N_7438);
nor U7503 (N_7503,N_7432,N_7365);
nand U7504 (N_7504,N_7382,N_7376);
and U7505 (N_7505,N_7499,N_7327);
or U7506 (N_7506,N_7310,N_7319);
and U7507 (N_7507,N_7403,N_7463);
nand U7508 (N_7508,N_7467,N_7406);
nand U7509 (N_7509,N_7426,N_7289);
nand U7510 (N_7510,N_7356,N_7293);
and U7511 (N_7511,N_7381,N_7411);
xor U7512 (N_7512,N_7219,N_7313);
nor U7513 (N_7513,N_7425,N_7216);
and U7514 (N_7514,N_7235,N_7421);
xnor U7515 (N_7515,N_7209,N_7484);
or U7516 (N_7516,N_7245,N_7408);
nand U7517 (N_7517,N_7392,N_7480);
or U7518 (N_7518,N_7343,N_7318);
and U7519 (N_7519,N_7283,N_7455);
nand U7520 (N_7520,N_7460,N_7349);
nor U7521 (N_7521,N_7419,N_7324);
and U7522 (N_7522,N_7331,N_7462);
and U7523 (N_7523,N_7314,N_7494);
xor U7524 (N_7524,N_7336,N_7221);
or U7525 (N_7525,N_7272,N_7423);
nor U7526 (N_7526,N_7237,N_7290);
xnor U7527 (N_7527,N_7291,N_7368);
nor U7528 (N_7528,N_7364,N_7266);
and U7529 (N_7529,N_7263,N_7225);
or U7530 (N_7530,N_7397,N_7475);
nor U7531 (N_7531,N_7371,N_7281);
nor U7532 (N_7532,N_7299,N_7352);
xnor U7533 (N_7533,N_7434,N_7479);
nand U7534 (N_7534,N_7208,N_7278);
xnor U7535 (N_7535,N_7335,N_7451);
nand U7536 (N_7536,N_7442,N_7389);
or U7537 (N_7537,N_7370,N_7354);
nor U7538 (N_7538,N_7413,N_7207);
nand U7539 (N_7539,N_7410,N_7280);
nor U7540 (N_7540,N_7328,N_7301);
and U7541 (N_7541,N_7436,N_7294);
and U7542 (N_7542,N_7270,N_7461);
nor U7543 (N_7543,N_7447,N_7456);
and U7544 (N_7544,N_7353,N_7435);
or U7545 (N_7545,N_7302,N_7362);
or U7546 (N_7546,N_7340,N_7261);
and U7547 (N_7547,N_7418,N_7401);
nor U7548 (N_7548,N_7303,N_7220);
or U7549 (N_7549,N_7407,N_7427);
nand U7550 (N_7550,N_7330,N_7206);
nand U7551 (N_7551,N_7262,N_7342);
xor U7552 (N_7552,N_7396,N_7309);
and U7553 (N_7553,N_7474,N_7443);
nand U7554 (N_7554,N_7471,N_7469);
nand U7555 (N_7555,N_7269,N_7264);
and U7556 (N_7556,N_7444,N_7440);
nor U7557 (N_7557,N_7317,N_7493);
or U7558 (N_7558,N_7488,N_7268);
or U7559 (N_7559,N_7476,N_7372);
nand U7560 (N_7560,N_7402,N_7379);
nand U7561 (N_7561,N_7325,N_7374);
nand U7562 (N_7562,N_7387,N_7405);
nor U7563 (N_7563,N_7449,N_7483);
xor U7564 (N_7564,N_7273,N_7253);
xnor U7565 (N_7565,N_7429,N_7450);
and U7566 (N_7566,N_7229,N_7468);
or U7567 (N_7567,N_7366,N_7250);
nand U7568 (N_7568,N_7399,N_7234);
xor U7569 (N_7569,N_7489,N_7296);
xnor U7570 (N_7570,N_7390,N_7200);
nand U7571 (N_7571,N_7380,N_7276);
nor U7572 (N_7572,N_7217,N_7214);
xnor U7573 (N_7573,N_7428,N_7248);
or U7574 (N_7574,N_7232,N_7358);
or U7575 (N_7575,N_7271,N_7414);
nor U7576 (N_7576,N_7482,N_7497);
or U7577 (N_7577,N_7333,N_7465);
nor U7578 (N_7578,N_7230,N_7385);
xor U7579 (N_7579,N_7348,N_7305);
nand U7580 (N_7580,N_7202,N_7393);
nor U7581 (N_7581,N_7466,N_7252);
xnor U7582 (N_7582,N_7334,N_7367);
or U7583 (N_7583,N_7323,N_7363);
nand U7584 (N_7584,N_7203,N_7255);
and U7585 (N_7585,N_7256,N_7486);
nand U7586 (N_7586,N_7251,N_7312);
nor U7587 (N_7587,N_7490,N_7201);
nor U7588 (N_7588,N_7445,N_7236);
nand U7589 (N_7589,N_7400,N_7424);
xor U7590 (N_7590,N_7260,N_7375);
xnor U7591 (N_7591,N_7254,N_7257);
or U7592 (N_7592,N_7338,N_7388);
or U7593 (N_7593,N_7446,N_7345);
and U7594 (N_7594,N_7258,N_7339);
nand U7595 (N_7595,N_7239,N_7259);
and U7596 (N_7596,N_7391,N_7282);
nand U7597 (N_7597,N_7226,N_7287);
nor U7598 (N_7598,N_7241,N_7240);
and U7599 (N_7599,N_7373,N_7320);
xor U7600 (N_7600,N_7496,N_7265);
nor U7601 (N_7601,N_7224,N_7420);
nand U7602 (N_7602,N_7495,N_7360);
nand U7603 (N_7603,N_7249,N_7341);
and U7604 (N_7604,N_7459,N_7223);
nor U7605 (N_7605,N_7383,N_7404);
nor U7606 (N_7606,N_7298,N_7300);
nor U7607 (N_7607,N_7417,N_7395);
nand U7608 (N_7608,N_7347,N_7398);
or U7609 (N_7609,N_7285,N_7409);
or U7610 (N_7610,N_7277,N_7204);
and U7611 (N_7611,N_7369,N_7377);
and U7612 (N_7612,N_7304,N_7437);
and U7613 (N_7613,N_7321,N_7470);
xor U7614 (N_7614,N_7246,N_7247);
nand U7615 (N_7615,N_7238,N_7337);
or U7616 (N_7616,N_7227,N_7211);
nand U7617 (N_7617,N_7458,N_7233);
nand U7618 (N_7618,N_7498,N_7492);
xor U7619 (N_7619,N_7215,N_7297);
xnor U7620 (N_7620,N_7464,N_7213);
and U7621 (N_7621,N_7457,N_7284);
nor U7622 (N_7622,N_7359,N_7412);
and U7623 (N_7623,N_7448,N_7357);
or U7624 (N_7624,N_7288,N_7415);
xor U7625 (N_7625,N_7441,N_7351);
xnor U7626 (N_7626,N_7267,N_7275);
xnor U7627 (N_7627,N_7311,N_7430);
or U7628 (N_7628,N_7279,N_7286);
or U7629 (N_7629,N_7243,N_7350);
and U7630 (N_7630,N_7487,N_7485);
nand U7631 (N_7631,N_7472,N_7212);
nor U7632 (N_7632,N_7231,N_7422);
and U7633 (N_7633,N_7355,N_7378);
or U7634 (N_7634,N_7394,N_7228);
and U7635 (N_7635,N_7326,N_7361);
and U7636 (N_7636,N_7218,N_7431);
nor U7637 (N_7637,N_7332,N_7344);
nor U7638 (N_7638,N_7346,N_7295);
xor U7639 (N_7639,N_7242,N_7329);
or U7640 (N_7640,N_7481,N_7478);
nand U7641 (N_7641,N_7316,N_7453);
xnor U7642 (N_7642,N_7491,N_7433);
nor U7643 (N_7643,N_7307,N_7477);
and U7644 (N_7644,N_7384,N_7274);
nand U7645 (N_7645,N_7292,N_7439);
and U7646 (N_7646,N_7308,N_7454);
and U7647 (N_7647,N_7416,N_7222);
and U7648 (N_7648,N_7473,N_7315);
xor U7649 (N_7649,N_7210,N_7244);
nor U7650 (N_7650,N_7334,N_7252);
and U7651 (N_7651,N_7447,N_7398);
xnor U7652 (N_7652,N_7309,N_7214);
nor U7653 (N_7653,N_7475,N_7385);
and U7654 (N_7654,N_7443,N_7253);
xor U7655 (N_7655,N_7478,N_7361);
and U7656 (N_7656,N_7221,N_7289);
or U7657 (N_7657,N_7314,N_7498);
or U7658 (N_7658,N_7336,N_7395);
nor U7659 (N_7659,N_7290,N_7447);
nor U7660 (N_7660,N_7238,N_7235);
nor U7661 (N_7661,N_7205,N_7333);
or U7662 (N_7662,N_7367,N_7438);
or U7663 (N_7663,N_7240,N_7259);
nand U7664 (N_7664,N_7284,N_7430);
xor U7665 (N_7665,N_7279,N_7402);
or U7666 (N_7666,N_7382,N_7299);
xnor U7667 (N_7667,N_7439,N_7383);
nor U7668 (N_7668,N_7377,N_7262);
or U7669 (N_7669,N_7413,N_7474);
or U7670 (N_7670,N_7214,N_7359);
nor U7671 (N_7671,N_7379,N_7336);
xor U7672 (N_7672,N_7472,N_7201);
and U7673 (N_7673,N_7477,N_7341);
or U7674 (N_7674,N_7280,N_7324);
nor U7675 (N_7675,N_7290,N_7236);
nand U7676 (N_7676,N_7430,N_7395);
and U7677 (N_7677,N_7450,N_7399);
or U7678 (N_7678,N_7207,N_7224);
or U7679 (N_7679,N_7387,N_7230);
xor U7680 (N_7680,N_7420,N_7470);
xor U7681 (N_7681,N_7301,N_7485);
nor U7682 (N_7682,N_7333,N_7281);
nor U7683 (N_7683,N_7313,N_7286);
xnor U7684 (N_7684,N_7267,N_7328);
or U7685 (N_7685,N_7322,N_7298);
xnor U7686 (N_7686,N_7300,N_7370);
and U7687 (N_7687,N_7261,N_7473);
or U7688 (N_7688,N_7263,N_7403);
nand U7689 (N_7689,N_7286,N_7258);
nand U7690 (N_7690,N_7240,N_7228);
nor U7691 (N_7691,N_7339,N_7341);
xor U7692 (N_7692,N_7374,N_7345);
or U7693 (N_7693,N_7375,N_7252);
nand U7694 (N_7694,N_7207,N_7243);
or U7695 (N_7695,N_7216,N_7448);
nand U7696 (N_7696,N_7437,N_7329);
and U7697 (N_7697,N_7406,N_7474);
nand U7698 (N_7698,N_7231,N_7290);
or U7699 (N_7699,N_7231,N_7230);
or U7700 (N_7700,N_7436,N_7448);
and U7701 (N_7701,N_7476,N_7401);
nor U7702 (N_7702,N_7318,N_7231);
and U7703 (N_7703,N_7488,N_7240);
xnor U7704 (N_7704,N_7251,N_7434);
nand U7705 (N_7705,N_7340,N_7301);
xnor U7706 (N_7706,N_7403,N_7413);
nand U7707 (N_7707,N_7201,N_7483);
nor U7708 (N_7708,N_7378,N_7388);
nor U7709 (N_7709,N_7429,N_7442);
xor U7710 (N_7710,N_7440,N_7350);
or U7711 (N_7711,N_7366,N_7202);
nand U7712 (N_7712,N_7222,N_7378);
nand U7713 (N_7713,N_7400,N_7419);
xor U7714 (N_7714,N_7493,N_7258);
nand U7715 (N_7715,N_7236,N_7394);
nand U7716 (N_7716,N_7269,N_7395);
xor U7717 (N_7717,N_7258,N_7395);
nor U7718 (N_7718,N_7339,N_7289);
nand U7719 (N_7719,N_7475,N_7498);
xnor U7720 (N_7720,N_7424,N_7390);
nand U7721 (N_7721,N_7318,N_7214);
nand U7722 (N_7722,N_7460,N_7490);
nor U7723 (N_7723,N_7371,N_7481);
nand U7724 (N_7724,N_7372,N_7255);
or U7725 (N_7725,N_7209,N_7415);
nand U7726 (N_7726,N_7381,N_7404);
or U7727 (N_7727,N_7468,N_7376);
nand U7728 (N_7728,N_7483,N_7264);
nor U7729 (N_7729,N_7360,N_7331);
nor U7730 (N_7730,N_7419,N_7336);
xor U7731 (N_7731,N_7245,N_7406);
nor U7732 (N_7732,N_7228,N_7209);
nor U7733 (N_7733,N_7362,N_7344);
or U7734 (N_7734,N_7263,N_7281);
xor U7735 (N_7735,N_7495,N_7275);
or U7736 (N_7736,N_7495,N_7249);
and U7737 (N_7737,N_7363,N_7455);
xor U7738 (N_7738,N_7239,N_7348);
and U7739 (N_7739,N_7214,N_7351);
and U7740 (N_7740,N_7323,N_7312);
nand U7741 (N_7741,N_7463,N_7482);
xnor U7742 (N_7742,N_7202,N_7288);
nand U7743 (N_7743,N_7386,N_7210);
or U7744 (N_7744,N_7257,N_7327);
nor U7745 (N_7745,N_7460,N_7462);
and U7746 (N_7746,N_7456,N_7485);
nor U7747 (N_7747,N_7303,N_7271);
nand U7748 (N_7748,N_7280,N_7209);
nand U7749 (N_7749,N_7330,N_7236);
xor U7750 (N_7750,N_7455,N_7421);
and U7751 (N_7751,N_7334,N_7462);
nand U7752 (N_7752,N_7410,N_7225);
xnor U7753 (N_7753,N_7339,N_7407);
xor U7754 (N_7754,N_7398,N_7250);
nand U7755 (N_7755,N_7222,N_7207);
and U7756 (N_7756,N_7483,N_7322);
or U7757 (N_7757,N_7365,N_7335);
xor U7758 (N_7758,N_7475,N_7274);
or U7759 (N_7759,N_7406,N_7361);
or U7760 (N_7760,N_7247,N_7408);
or U7761 (N_7761,N_7304,N_7462);
xnor U7762 (N_7762,N_7394,N_7490);
nor U7763 (N_7763,N_7436,N_7254);
nor U7764 (N_7764,N_7449,N_7408);
and U7765 (N_7765,N_7231,N_7227);
or U7766 (N_7766,N_7357,N_7464);
or U7767 (N_7767,N_7492,N_7493);
nand U7768 (N_7768,N_7378,N_7464);
nand U7769 (N_7769,N_7380,N_7420);
xnor U7770 (N_7770,N_7400,N_7245);
xnor U7771 (N_7771,N_7373,N_7398);
or U7772 (N_7772,N_7380,N_7359);
or U7773 (N_7773,N_7331,N_7470);
or U7774 (N_7774,N_7405,N_7211);
nor U7775 (N_7775,N_7376,N_7425);
nand U7776 (N_7776,N_7329,N_7381);
nor U7777 (N_7777,N_7239,N_7421);
nor U7778 (N_7778,N_7340,N_7418);
nor U7779 (N_7779,N_7244,N_7296);
nor U7780 (N_7780,N_7398,N_7499);
and U7781 (N_7781,N_7315,N_7434);
nor U7782 (N_7782,N_7203,N_7264);
nand U7783 (N_7783,N_7303,N_7446);
nor U7784 (N_7784,N_7306,N_7219);
nand U7785 (N_7785,N_7210,N_7400);
nor U7786 (N_7786,N_7263,N_7430);
and U7787 (N_7787,N_7345,N_7334);
nand U7788 (N_7788,N_7394,N_7312);
and U7789 (N_7789,N_7342,N_7396);
or U7790 (N_7790,N_7338,N_7324);
and U7791 (N_7791,N_7412,N_7283);
nor U7792 (N_7792,N_7243,N_7286);
and U7793 (N_7793,N_7427,N_7251);
xor U7794 (N_7794,N_7468,N_7352);
nor U7795 (N_7795,N_7222,N_7465);
nand U7796 (N_7796,N_7440,N_7400);
nor U7797 (N_7797,N_7351,N_7400);
or U7798 (N_7798,N_7286,N_7242);
or U7799 (N_7799,N_7411,N_7439);
nor U7800 (N_7800,N_7532,N_7551);
xor U7801 (N_7801,N_7716,N_7600);
xor U7802 (N_7802,N_7777,N_7683);
xor U7803 (N_7803,N_7796,N_7688);
and U7804 (N_7804,N_7743,N_7611);
nand U7805 (N_7805,N_7646,N_7511);
or U7806 (N_7806,N_7776,N_7545);
and U7807 (N_7807,N_7571,N_7508);
nand U7808 (N_7808,N_7579,N_7725);
or U7809 (N_7809,N_7710,N_7669);
or U7810 (N_7810,N_7699,N_7558);
nor U7811 (N_7811,N_7542,N_7554);
and U7812 (N_7812,N_7745,N_7513);
nand U7813 (N_7813,N_7754,N_7557);
and U7814 (N_7814,N_7578,N_7589);
nand U7815 (N_7815,N_7649,N_7698);
nor U7816 (N_7816,N_7500,N_7522);
or U7817 (N_7817,N_7735,N_7661);
xor U7818 (N_7818,N_7723,N_7520);
xor U7819 (N_7819,N_7761,N_7679);
nand U7820 (N_7820,N_7676,N_7733);
or U7821 (N_7821,N_7724,N_7657);
or U7822 (N_7822,N_7591,N_7539);
xor U7823 (N_7823,N_7708,N_7531);
xnor U7824 (N_7824,N_7555,N_7598);
xnor U7825 (N_7825,N_7566,N_7622);
and U7826 (N_7826,N_7757,N_7677);
or U7827 (N_7827,N_7643,N_7665);
xor U7828 (N_7828,N_7632,N_7667);
xnor U7829 (N_7829,N_7798,N_7625);
nand U7830 (N_7830,N_7595,N_7626);
nor U7831 (N_7831,N_7652,N_7728);
xnor U7832 (N_7832,N_7516,N_7785);
nand U7833 (N_7833,N_7678,N_7507);
or U7834 (N_7834,N_7592,N_7597);
or U7835 (N_7835,N_7616,N_7529);
and U7836 (N_7836,N_7568,N_7791);
nand U7837 (N_7837,N_7779,N_7506);
nand U7838 (N_7838,N_7707,N_7523);
nor U7839 (N_7839,N_7758,N_7627);
and U7840 (N_7840,N_7730,N_7739);
nor U7841 (N_7841,N_7764,N_7717);
nand U7842 (N_7842,N_7623,N_7561);
xor U7843 (N_7843,N_7590,N_7587);
nor U7844 (N_7844,N_7560,N_7747);
nor U7845 (N_7845,N_7624,N_7521);
xor U7846 (N_7846,N_7713,N_7572);
or U7847 (N_7847,N_7606,N_7570);
xnor U7848 (N_7848,N_7619,N_7547);
nand U7849 (N_7849,N_7629,N_7795);
or U7850 (N_7850,N_7663,N_7709);
xnor U7851 (N_7851,N_7794,N_7505);
nor U7852 (N_7852,N_7656,N_7687);
nor U7853 (N_7853,N_7536,N_7573);
and U7854 (N_7854,N_7650,N_7790);
xnor U7855 (N_7855,N_7690,N_7799);
nor U7856 (N_7856,N_7635,N_7540);
or U7857 (N_7857,N_7773,N_7648);
nor U7858 (N_7858,N_7778,N_7530);
xnor U7859 (N_7859,N_7524,N_7509);
and U7860 (N_7860,N_7565,N_7769);
xor U7861 (N_7861,N_7613,N_7768);
xnor U7862 (N_7862,N_7783,N_7762);
nor U7863 (N_7863,N_7519,N_7527);
nand U7864 (N_7864,N_7670,N_7692);
nor U7865 (N_7865,N_7603,N_7628);
xor U7866 (N_7866,N_7680,N_7740);
or U7867 (N_7867,N_7602,N_7548);
or U7868 (N_7868,N_7546,N_7541);
or U7869 (N_7869,N_7681,N_7689);
and U7870 (N_7870,N_7780,N_7787);
or U7871 (N_7871,N_7766,N_7697);
xnor U7872 (N_7872,N_7515,N_7714);
and U7873 (N_7873,N_7550,N_7720);
nor U7874 (N_7874,N_7782,N_7574);
or U7875 (N_7875,N_7586,N_7731);
xor U7876 (N_7876,N_7615,N_7612);
nand U7877 (N_7877,N_7582,N_7537);
nand U7878 (N_7878,N_7750,N_7746);
and U7879 (N_7879,N_7759,N_7621);
xor U7880 (N_7880,N_7748,N_7775);
or U7881 (N_7881,N_7633,N_7651);
and U7882 (N_7882,N_7771,N_7647);
and U7883 (N_7883,N_7639,N_7577);
nand U7884 (N_7884,N_7696,N_7614);
or U7885 (N_7885,N_7630,N_7672);
or U7886 (N_7886,N_7585,N_7749);
nor U7887 (N_7887,N_7642,N_7772);
or U7888 (N_7888,N_7664,N_7737);
and U7889 (N_7889,N_7559,N_7684);
xnor U7890 (N_7890,N_7788,N_7610);
nor U7891 (N_7891,N_7607,N_7502);
and U7892 (N_7892,N_7556,N_7767);
nand U7893 (N_7893,N_7593,N_7753);
or U7894 (N_7894,N_7755,N_7658);
nand U7895 (N_7895,N_7567,N_7662);
nor U7896 (N_7896,N_7605,N_7534);
xor U7897 (N_7897,N_7752,N_7641);
or U7898 (N_7898,N_7721,N_7793);
nand U7899 (N_7899,N_7514,N_7770);
and U7900 (N_7900,N_7617,N_7654);
nand U7901 (N_7901,N_7640,N_7682);
nor U7902 (N_7902,N_7702,N_7666);
or U7903 (N_7903,N_7715,N_7634);
nand U7904 (N_7904,N_7774,N_7638);
or U7905 (N_7905,N_7580,N_7674);
nor U7906 (N_7906,N_7742,N_7608);
and U7907 (N_7907,N_7694,N_7659);
nor U7908 (N_7908,N_7660,N_7594);
nor U7909 (N_7909,N_7518,N_7562);
nand U7910 (N_7910,N_7789,N_7703);
and U7911 (N_7911,N_7701,N_7576);
and U7912 (N_7912,N_7575,N_7784);
xor U7913 (N_7913,N_7552,N_7538);
and U7914 (N_7914,N_7525,N_7644);
nand U7915 (N_7915,N_7738,N_7792);
nand U7916 (N_7916,N_7706,N_7510);
nand U7917 (N_7917,N_7563,N_7569);
nor U7918 (N_7918,N_7693,N_7726);
or U7919 (N_7919,N_7718,N_7751);
and U7920 (N_7920,N_7655,N_7736);
nand U7921 (N_7921,N_7584,N_7620);
nor U7922 (N_7922,N_7583,N_7704);
or U7923 (N_7923,N_7637,N_7596);
xnor U7924 (N_7924,N_7503,N_7763);
and U7925 (N_7925,N_7671,N_7609);
or U7926 (N_7926,N_7588,N_7744);
and U7927 (N_7927,N_7705,N_7695);
nand U7928 (N_7928,N_7673,N_7734);
nand U7929 (N_7929,N_7544,N_7564);
nor U7930 (N_7930,N_7781,N_7722);
nand U7931 (N_7931,N_7712,N_7711);
or U7932 (N_7932,N_7653,N_7553);
nand U7933 (N_7933,N_7549,N_7691);
nor U7934 (N_7934,N_7517,N_7741);
nand U7935 (N_7935,N_7727,N_7528);
xor U7936 (N_7936,N_7543,N_7645);
nor U7937 (N_7937,N_7760,N_7685);
xnor U7938 (N_7938,N_7604,N_7601);
and U7939 (N_7939,N_7636,N_7535);
xor U7940 (N_7940,N_7631,N_7533);
or U7941 (N_7941,N_7504,N_7618);
and U7942 (N_7942,N_7526,N_7599);
nor U7943 (N_7943,N_7797,N_7668);
nand U7944 (N_7944,N_7732,N_7765);
or U7945 (N_7945,N_7729,N_7786);
and U7946 (N_7946,N_7501,N_7700);
nand U7947 (N_7947,N_7756,N_7581);
nand U7948 (N_7948,N_7512,N_7675);
nand U7949 (N_7949,N_7686,N_7719);
or U7950 (N_7950,N_7630,N_7545);
nand U7951 (N_7951,N_7682,N_7588);
nor U7952 (N_7952,N_7660,N_7627);
nand U7953 (N_7953,N_7744,N_7544);
xnor U7954 (N_7954,N_7593,N_7586);
and U7955 (N_7955,N_7701,N_7666);
nand U7956 (N_7956,N_7610,N_7586);
nor U7957 (N_7957,N_7647,N_7712);
nor U7958 (N_7958,N_7784,N_7780);
nor U7959 (N_7959,N_7556,N_7783);
xor U7960 (N_7960,N_7609,N_7678);
or U7961 (N_7961,N_7653,N_7586);
and U7962 (N_7962,N_7759,N_7597);
or U7963 (N_7963,N_7760,N_7751);
or U7964 (N_7964,N_7520,N_7663);
nor U7965 (N_7965,N_7717,N_7749);
nand U7966 (N_7966,N_7795,N_7639);
or U7967 (N_7967,N_7762,N_7644);
nand U7968 (N_7968,N_7783,N_7715);
nand U7969 (N_7969,N_7580,N_7631);
or U7970 (N_7970,N_7563,N_7500);
or U7971 (N_7971,N_7795,N_7734);
nor U7972 (N_7972,N_7737,N_7569);
nand U7973 (N_7973,N_7718,N_7685);
and U7974 (N_7974,N_7644,N_7628);
nor U7975 (N_7975,N_7774,N_7729);
or U7976 (N_7976,N_7689,N_7793);
and U7977 (N_7977,N_7504,N_7746);
and U7978 (N_7978,N_7645,N_7690);
nand U7979 (N_7979,N_7664,N_7681);
xor U7980 (N_7980,N_7578,N_7795);
and U7981 (N_7981,N_7538,N_7542);
nand U7982 (N_7982,N_7726,N_7512);
nand U7983 (N_7983,N_7566,N_7710);
or U7984 (N_7984,N_7725,N_7661);
xnor U7985 (N_7985,N_7571,N_7674);
nand U7986 (N_7986,N_7607,N_7605);
xor U7987 (N_7987,N_7655,N_7514);
or U7988 (N_7988,N_7636,N_7783);
xnor U7989 (N_7989,N_7561,N_7759);
nand U7990 (N_7990,N_7560,N_7569);
and U7991 (N_7991,N_7632,N_7795);
nor U7992 (N_7992,N_7527,N_7747);
or U7993 (N_7993,N_7555,N_7549);
nand U7994 (N_7994,N_7697,N_7686);
xnor U7995 (N_7995,N_7721,N_7744);
or U7996 (N_7996,N_7775,N_7658);
nor U7997 (N_7997,N_7771,N_7630);
and U7998 (N_7998,N_7591,N_7713);
and U7999 (N_7999,N_7712,N_7523);
nor U8000 (N_8000,N_7623,N_7775);
and U8001 (N_8001,N_7742,N_7700);
xor U8002 (N_8002,N_7519,N_7587);
and U8003 (N_8003,N_7710,N_7571);
nor U8004 (N_8004,N_7550,N_7745);
or U8005 (N_8005,N_7792,N_7615);
xor U8006 (N_8006,N_7777,N_7580);
xnor U8007 (N_8007,N_7717,N_7681);
xnor U8008 (N_8008,N_7629,N_7594);
xor U8009 (N_8009,N_7673,N_7503);
nand U8010 (N_8010,N_7678,N_7578);
nand U8011 (N_8011,N_7694,N_7621);
or U8012 (N_8012,N_7519,N_7592);
xnor U8013 (N_8013,N_7752,N_7767);
xnor U8014 (N_8014,N_7725,N_7608);
xnor U8015 (N_8015,N_7648,N_7664);
xnor U8016 (N_8016,N_7562,N_7550);
or U8017 (N_8017,N_7658,N_7586);
nand U8018 (N_8018,N_7533,N_7536);
and U8019 (N_8019,N_7524,N_7717);
nor U8020 (N_8020,N_7762,N_7538);
xnor U8021 (N_8021,N_7683,N_7603);
nand U8022 (N_8022,N_7689,N_7665);
and U8023 (N_8023,N_7576,N_7724);
or U8024 (N_8024,N_7621,N_7597);
nand U8025 (N_8025,N_7729,N_7512);
nand U8026 (N_8026,N_7559,N_7739);
xnor U8027 (N_8027,N_7727,N_7503);
and U8028 (N_8028,N_7697,N_7663);
nor U8029 (N_8029,N_7770,N_7790);
xnor U8030 (N_8030,N_7655,N_7686);
xnor U8031 (N_8031,N_7749,N_7719);
xor U8032 (N_8032,N_7547,N_7609);
xnor U8033 (N_8033,N_7656,N_7676);
or U8034 (N_8034,N_7585,N_7725);
xnor U8035 (N_8035,N_7658,N_7679);
xnor U8036 (N_8036,N_7611,N_7508);
nor U8037 (N_8037,N_7685,N_7777);
and U8038 (N_8038,N_7523,N_7649);
nor U8039 (N_8039,N_7796,N_7604);
xor U8040 (N_8040,N_7551,N_7649);
xor U8041 (N_8041,N_7678,N_7544);
nor U8042 (N_8042,N_7774,N_7613);
nor U8043 (N_8043,N_7568,N_7665);
xnor U8044 (N_8044,N_7697,N_7605);
and U8045 (N_8045,N_7681,N_7760);
nand U8046 (N_8046,N_7618,N_7657);
nor U8047 (N_8047,N_7794,N_7623);
nor U8048 (N_8048,N_7791,N_7746);
or U8049 (N_8049,N_7551,N_7598);
and U8050 (N_8050,N_7671,N_7677);
nor U8051 (N_8051,N_7525,N_7648);
nand U8052 (N_8052,N_7652,N_7551);
xor U8053 (N_8053,N_7759,N_7583);
nor U8054 (N_8054,N_7777,N_7712);
nand U8055 (N_8055,N_7658,N_7672);
and U8056 (N_8056,N_7688,N_7541);
nor U8057 (N_8057,N_7624,N_7590);
xnor U8058 (N_8058,N_7514,N_7534);
nand U8059 (N_8059,N_7648,N_7574);
xnor U8060 (N_8060,N_7605,N_7764);
and U8061 (N_8061,N_7571,N_7549);
nand U8062 (N_8062,N_7583,N_7610);
or U8063 (N_8063,N_7700,N_7701);
nor U8064 (N_8064,N_7677,N_7737);
or U8065 (N_8065,N_7661,N_7670);
xor U8066 (N_8066,N_7670,N_7709);
nand U8067 (N_8067,N_7535,N_7766);
nand U8068 (N_8068,N_7543,N_7747);
or U8069 (N_8069,N_7526,N_7560);
or U8070 (N_8070,N_7751,N_7765);
and U8071 (N_8071,N_7513,N_7527);
and U8072 (N_8072,N_7782,N_7508);
nor U8073 (N_8073,N_7607,N_7786);
nand U8074 (N_8074,N_7575,N_7501);
and U8075 (N_8075,N_7623,N_7579);
nor U8076 (N_8076,N_7534,N_7677);
and U8077 (N_8077,N_7624,N_7746);
nand U8078 (N_8078,N_7540,N_7553);
and U8079 (N_8079,N_7787,N_7769);
and U8080 (N_8080,N_7560,N_7716);
nand U8081 (N_8081,N_7668,N_7610);
xnor U8082 (N_8082,N_7739,N_7570);
nand U8083 (N_8083,N_7638,N_7740);
xor U8084 (N_8084,N_7650,N_7561);
nand U8085 (N_8085,N_7650,N_7508);
and U8086 (N_8086,N_7572,N_7643);
xor U8087 (N_8087,N_7521,N_7740);
nand U8088 (N_8088,N_7715,N_7598);
xor U8089 (N_8089,N_7758,N_7609);
nor U8090 (N_8090,N_7760,N_7750);
or U8091 (N_8091,N_7567,N_7755);
nor U8092 (N_8092,N_7502,N_7609);
and U8093 (N_8093,N_7723,N_7733);
or U8094 (N_8094,N_7665,N_7769);
nor U8095 (N_8095,N_7540,N_7634);
nand U8096 (N_8096,N_7753,N_7578);
nand U8097 (N_8097,N_7746,N_7758);
or U8098 (N_8098,N_7579,N_7687);
or U8099 (N_8099,N_7728,N_7718);
nor U8100 (N_8100,N_7855,N_8099);
and U8101 (N_8101,N_8052,N_8024);
and U8102 (N_8102,N_8056,N_8074);
nand U8103 (N_8103,N_8044,N_7928);
or U8104 (N_8104,N_7891,N_7997);
or U8105 (N_8105,N_7868,N_8039);
xnor U8106 (N_8106,N_8084,N_7939);
nand U8107 (N_8107,N_8058,N_7989);
xor U8108 (N_8108,N_7859,N_8060);
and U8109 (N_8109,N_8010,N_7958);
nand U8110 (N_8110,N_7892,N_7825);
nand U8111 (N_8111,N_8021,N_7974);
and U8112 (N_8112,N_8059,N_7996);
or U8113 (N_8113,N_7967,N_8098);
xor U8114 (N_8114,N_7986,N_8003);
and U8115 (N_8115,N_7903,N_7879);
and U8116 (N_8116,N_8041,N_8035);
or U8117 (N_8117,N_7864,N_7914);
nor U8118 (N_8118,N_8008,N_8028);
xnor U8119 (N_8119,N_7959,N_7975);
nand U8120 (N_8120,N_7888,N_7810);
nand U8121 (N_8121,N_7957,N_7964);
and U8122 (N_8122,N_8065,N_7883);
xnor U8123 (N_8123,N_7884,N_7893);
nor U8124 (N_8124,N_8081,N_7906);
nand U8125 (N_8125,N_8033,N_7886);
nor U8126 (N_8126,N_7822,N_7937);
nor U8127 (N_8127,N_8034,N_7858);
nand U8128 (N_8128,N_7970,N_8090);
or U8129 (N_8129,N_7932,N_7995);
nor U8130 (N_8130,N_7811,N_7870);
and U8131 (N_8131,N_7815,N_7952);
nor U8132 (N_8132,N_8015,N_7818);
xnor U8133 (N_8133,N_7940,N_7999);
nor U8134 (N_8134,N_7807,N_7934);
and U8135 (N_8135,N_8020,N_8023);
xor U8136 (N_8136,N_7878,N_7808);
nor U8137 (N_8137,N_7968,N_7987);
and U8138 (N_8138,N_8030,N_7881);
nand U8139 (N_8139,N_7911,N_7850);
and U8140 (N_8140,N_8053,N_8091);
nand U8141 (N_8141,N_8050,N_7904);
nand U8142 (N_8142,N_7935,N_8097);
or U8143 (N_8143,N_8018,N_7834);
and U8144 (N_8144,N_8085,N_8040);
and U8145 (N_8145,N_8083,N_7917);
nor U8146 (N_8146,N_8013,N_7889);
or U8147 (N_8147,N_8076,N_7938);
nor U8148 (N_8148,N_7953,N_7946);
nand U8149 (N_8149,N_7988,N_7865);
and U8150 (N_8150,N_7910,N_7947);
or U8151 (N_8151,N_8054,N_7843);
nand U8152 (N_8152,N_7972,N_7844);
and U8153 (N_8153,N_7944,N_8006);
nand U8154 (N_8154,N_8000,N_8075);
nand U8155 (N_8155,N_8066,N_8027);
and U8156 (N_8156,N_7907,N_7824);
nand U8157 (N_8157,N_7916,N_7877);
nand U8158 (N_8158,N_7875,N_7918);
and U8159 (N_8159,N_7821,N_7860);
and U8160 (N_8160,N_7926,N_7924);
xor U8161 (N_8161,N_7949,N_8011);
nand U8162 (N_8162,N_7880,N_7896);
nor U8163 (N_8163,N_7831,N_7913);
and U8164 (N_8164,N_7882,N_7945);
nor U8165 (N_8165,N_8064,N_7902);
nand U8166 (N_8166,N_7846,N_7943);
nor U8167 (N_8167,N_8012,N_8007);
or U8168 (N_8168,N_7998,N_7971);
nor U8169 (N_8169,N_7993,N_7871);
nor U8170 (N_8170,N_7894,N_8094);
xnor U8171 (N_8171,N_8017,N_7941);
or U8172 (N_8172,N_8068,N_8082);
or U8173 (N_8173,N_8048,N_7873);
nor U8174 (N_8174,N_7948,N_7981);
xnor U8175 (N_8175,N_7960,N_7931);
xor U8176 (N_8176,N_8061,N_7956);
and U8177 (N_8177,N_7857,N_7861);
nor U8178 (N_8178,N_7826,N_8080);
and U8179 (N_8179,N_7835,N_7982);
and U8180 (N_8180,N_7827,N_8072);
nand U8181 (N_8181,N_7921,N_8046);
and U8182 (N_8182,N_8049,N_8055);
nand U8183 (N_8183,N_7933,N_8029);
nor U8184 (N_8184,N_7994,N_8073);
nor U8185 (N_8185,N_7830,N_7898);
and U8186 (N_8186,N_7813,N_7900);
nor U8187 (N_8187,N_7923,N_7990);
nand U8188 (N_8188,N_8019,N_7866);
nor U8189 (N_8189,N_7833,N_8042);
or U8190 (N_8190,N_7849,N_8070);
xor U8191 (N_8191,N_7983,N_7980);
xor U8192 (N_8192,N_8038,N_7991);
or U8193 (N_8193,N_7929,N_8096);
or U8194 (N_8194,N_7848,N_7804);
and U8195 (N_8195,N_8002,N_7812);
nor U8196 (N_8196,N_7955,N_8057);
nand U8197 (N_8197,N_8093,N_7867);
xor U8198 (N_8198,N_7836,N_7954);
and U8199 (N_8199,N_8004,N_7806);
or U8200 (N_8200,N_8005,N_7828);
nor U8201 (N_8201,N_7909,N_7969);
nand U8202 (N_8202,N_8022,N_8088);
nor U8203 (N_8203,N_8045,N_7901);
xor U8204 (N_8204,N_7856,N_8026);
or U8205 (N_8205,N_7854,N_7805);
nand U8206 (N_8206,N_8001,N_8031);
xnor U8207 (N_8207,N_7847,N_7962);
xnor U8208 (N_8208,N_7899,N_7800);
or U8209 (N_8209,N_7966,N_7801);
or U8210 (N_8210,N_8087,N_8016);
or U8211 (N_8211,N_8051,N_7973);
or U8212 (N_8212,N_8032,N_7908);
and U8213 (N_8213,N_8069,N_7819);
nor U8214 (N_8214,N_7992,N_8089);
and U8215 (N_8215,N_7837,N_7852);
and U8216 (N_8216,N_7936,N_7927);
or U8217 (N_8217,N_7838,N_8086);
or U8218 (N_8218,N_7885,N_7802);
nor U8219 (N_8219,N_8043,N_7965);
xor U8220 (N_8220,N_8025,N_8037);
and U8221 (N_8221,N_7895,N_8079);
or U8222 (N_8222,N_8036,N_7951);
nand U8223 (N_8223,N_7803,N_8078);
and U8224 (N_8224,N_7984,N_8047);
and U8225 (N_8225,N_7922,N_7905);
xnor U8226 (N_8226,N_7816,N_7920);
xnor U8227 (N_8227,N_7890,N_7842);
xnor U8228 (N_8228,N_8095,N_7829);
xor U8229 (N_8229,N_7851,N_7814);
xnor U8230 (N_8230,N_7853,N_8067);
nor U8231 (N_8231,N_7942,N_7841);
xor U8232 (N_8232,N_8014,N_7977);
nor U8233 (N_8233,N_8062,N_7979);
or U8234 (N_8234,N_8071,N_7930);
and U8235 (N_8235,N_7912,N_8092);
xor U8236 (N_8236,N_7919,N_7978);
nor U8237 (N_8237,N_7872,N_7820);
nand U8238 (N_8238,N_7840,N_7817);
and U8239 (N_8239,N_8077,N_7863);
nor U8240 (N_8240,N_7887,N_8063);
and U8241 (N_8241,N_7862,N_7925);
and U8242 (N_8242,N_7961,N_7823);
nand U8243 (N_8243,N_7976,N_7845);
xnor U8244 (N_8244,N_7897,N_7809);
nand U8245 (N_8245,N_7874,N_7915);
nor U8246 (N_8246,N_8009,N_7839);
xor U8247 (N_8247,N_7869,N_7985);
and U8248 (N_8248,N_7963,N_7876);
nor U8249 (N_8249,N_7950,N_7832);
and U8250 (N_8250,N_7825,N_7885);
or U8251 (N_8251,N_7908,N_7863);
nor U8252 (N_8252,N_8048,N_7944);
xnor U8253 (N_8253,N_7838,N_7904);
nand U8254 (N_8254,N_7902,N_8051);
or U8255 (N_8255,N_7802,N_8050);
nand U8256 (N_8256,N_8041,N_7861);
and U8257 (N_8257,N_8002,N_7801);
xor U8258 (N_8258,N_7894,N_7968);
or U8259 (N_8259,N_7948,N_8080);
xor U8260 (N_8260,N_8011,N_7955);
nor U8261 (N_8261,N_8053,N_7900);
xor U8262 (N_8262,N_7909,N_7984);
and U8263 (N_8263,N_8064,N_7864);
and U8264 (N_8264,N_8093,N_7860);
nand U8265 (N_8265,N_8024,N_7974);
and U8266 (N_8266,N_8095,N_7962);
xnor U8267 (N_8267,N_8081,N_7857);
xor U8268 (N_8268,N_7870,N_8047);
or U8269 (N_8269,N_7880,N_8097);
and U8270 (N_8270,N_7833,N_8053);
xor U8271 (N_8271,N_8054,N_8004);
nor U8272 (N_8272,N_7935,N_7956);
nor U8273 (N_8273,N_7844,N_7837);
or U8274 (N_8274,N_7993,N_7841);
xor U8275 (N_8275,N_7941,N_8085);
or U8276 (N_8276,N_8054,N_7885);
nor U8277 (N_8277,N_7922,N_7957);
nor U8278 (N_8278,N_7854,N_8046);
and U8279 (N_8279,N_8024,N_7963);
nor U8280 (N_8280,N_8064,N_8074);
or U8281 (N_8281,N_7811,N_7854);
or U8282 (N_8282,N_7903,N_8073);
or U8283 (N_8283,N_8071,N_7974);
and U8284 (N_8284,N_8055,N_8048);
nand U8285 (N_8285,N_7953,N_7925);
xor U8286 (N_8286,N_7852,N_7806);
nor U8287 (N_8287,N_7876,N_8046);
xor U8288 (N_8288,N_7967,N_7932);
xnor U8289 (N_8289,N_8056,N_7849);
or U8290 (N_8290,N_7924,N_7854);
nand U8291 (N_8291,N_7968,N_7911);
and U8292 (N_8292,N_7963,N_8074);
xnor U8293 (N_8293,N_7868,N_7995);
nand U8294 (N_8294,N_7960,N_7859);
nand U8295 (N_8295,N_8022,N_7997);
nand U8296 (N_8296,N_7859,N_7874);
nor U8297 (N_8297,N_7835,N_8037);
nor U8298 (N_8298,N_7809,N_7934);
xor U8299 (N_8299,N_7838,N_7952);
nand U8300 (N_8300,N_7902,N_7928);
nand U8301 (N_8301,N_8035,N_7995);
and U8302 (N_8302,N_7946,N_8066);
nor U8303 (N_8303,N_8084,N_8076);
or U8304 (N_8304,N_8017,N_7973);
or U8305 (N_8305,N_8045,N_8029);
nand U8306 (N_8306,N_7848,N_8031);
nand U8307 (N_8307,N_7942,N_8031);
or U8308 (N_8308,N_8001,N_7962);
xor U8309 (N_8309,N_7934,N_7920);
xor U8310 (N_8310,N_8087,N_7819);
xnor U8311 (N_8311,N_8036,N_7949);
or U8312 (N_8312,N_8043,N_7815);
and U8313 (N_8313,N_8082,N_8031);
nor U8314 (N_8314,N_7938,N_7852);
or U8315 (N_8315,N_7973,N_8050);
nor U8316 (N_8316,N_8007,N_7905);
xor U8317 (N_8317,N_8094,N_7900);
nand U8318 (N_8318,N_7815,N_7973);
nor U8319 (N_8319,N_7846,N_8018);
nor U8320 (N_8320,N_7967,N_8086);
or U8321 (N_8321,N_7872,N_7924);
or U8322 (N_8322,N_7995,N_7845);
nor U8323 (N_8323,N_7941,N_7991);
and U8324 (N_8324,N_7845,N_7875);
nor U8325 (N_8325,N_8063,N_7997);
nor U8326 (N_8326,N_7944,N_7967);
and U8327 (N_8327,N_7848,N_7841);
or U8328 (N_8328,N_8050,N_7828);
nand U8329 (N_8329,N_7982,N_8086);
and U8330 (N_8330,N_8051,N_7903);
xor U8331 (N_8331,N_7855,N_7984);
or U8332 (N_8332,N_7906,N_8086);
or U8333 (N_8333,N_7989,N_7893);
xnor U8334 (N_8334,N_8010,N_8003);
and U8335 (N_8335,N_8083,N_7878);
or U8336 (N_8336,N_7863,N_8039);
or U8337 (N_8337,N_8048,N_7863);
nor U8338 (N_8338,N_7926,N_8094);
and U8339 (N_8339,N_7814,N_7876);
or U8340 (N_8340,N_7896,N_7814);
xnor U8341 (N_8341,N_7992,N_8074);
nor U8342 (N_8342,N_7948,N_7919);
nand U8343 (N_8343,N_7878,N_8054);
or U8344 (N_8344,N_8006,N_7883);
or U8345 (N_8345,N_7816,N_8039);
nor U8346 (N_8346,N_7861,N_7841);
xnor U8347 (N_8347,N_7951,N_7926);
nor U8348 (N_8348,N_8001,N_8034);
nand U8349 (N_8349,N_7920,N_8095);
and U8350 (N_8350,N_8099,N_7996);
nand U8351 (N_8351,N_8062,N_7873);
nand U8352 (N_8352,N_8022,N_7891);
and U8353 (N_8353,N_7964,N_7983);
nand U8354 (N_8354,N_8088,N_7912);
nand U8355 (N_8355,N_7959,N_7824);
nand U8356 (N_8356,N_7931,N_7855);
nand U8357 (N_8357,N_7848,N_8068);
xor U8358 (N_8358,N_8005,N_7902);
nor U8359 (N_8359,N_8059,N_8065);
nor U8360 (N_8360,N_8042,N_8014);
xor U8361 (N_8361,N_7850,N_8063);
and U8362 (N_8362,N_8008,N_8075);
and U8363 (N_8363,N_7829,N_7854);
nand U8364 (N_8364,N_7859,N_7970);
or U8365 (N_8365,N_7906,N_7846);
nor U8366 (N_8366,N_8073,N_7935);
nor U8367 (N_8367,N_8023,N_7889);
nand U8368 (N_8368,N_8028,N_8046);
and U8369 (N_8369,N_7837,N_7952);
xor U8370 (N_8370,N_7817,N_7979);
nand U8371 (N_8371,N_8024,N_8006);
and U8372 (N_8372,N_8044,N_7823);
nor U8373 (N_8373,N_8059,N_7934);
or U8374 (N_8374,N_8078,N_7920);
or U8375 (N_8375,N_8087,N_7863);
nor U8376 (N_8376,N_8088,N_8075);
nand U8377 (N_8377,N_8066,N_8073);
and U8378 (N_8378,N_8056,N_7814);
nor U8379 (N_8379,N_8036,N_7872);
or U8380 (N_8380,N_8059,N_7841);
nand U8381 (N_8381,N_7936,N_7977);
xnor U8382 (N_8382,N_8005,N_7905);
nor U8383 (N_8383,N_7885,N_7872);
or U8384 (N_8384,N_7867,N_7905);
xnor U8385 (N_8385,N_7901,N_8009);
and U8386 (N_8386,N_7855,N_7878);
nor U8387 (N_8387,N_7842,N_7827);
xor U8388 (N_8388,N_8032,N_8033);
and U8389 (N_8389,N_8022,N_8077);
nand U8390 (N_8390,N_7977,N_7828);
nand U8391 (N_8391,N_7991,N_7834);
nor U8392 (N_8392,N_8033,N_8078);
nand U8393 (N_8393,N_7959,N_7816);
and U8394 (N_8394,N_8026,N_7839);
or U8395 (N_8395,N_7980,N_8035);
or U8396 (N_8396,N_8062,N_8068);
and U8397 (N_8397,N_8009,N_8073);
nand U8398 (N_8398,N_8076,N_7808);
nand U8399 (N_8399,N_7839,N_7982);
or U8400 (N_8400,N_8262,N_8301);
nand U8401 (N_8401,N_8187,N_8297);
and U8402 (N_8402,N_8215,N_8238);
xnor U8403 (N_8403,N_8380,N_8246);
or U8404 (N_8404,N_8217,N_8237);
xnor U8405 (N_8405,N_8165,N_8328);
nor U8406 (N_8406,N_8386,N_8202);
nor U8407 (N_8407,N_8265,N_8389);
xor U8408 (N_8408,N_8211,N_8343);
xor U8409 (N_8409,N_8213,N_8330);
or U8410 (N_8410,N_8138,N_8371);
nand U8411 (N_8411,N_8180,N_8242);
nor U8412 (N_8412,N_8183,N_8379);
and U8413 (N_8413,N_8295,N_8231);
xor U8414 (N_8414,N_8120,N_8245);
or U8415 (N_8415,N_8333,N_8366);
xnor U8416 (N_8416,N_8164,N_8337);
nand U8417 (N_8417,N_8358,N_8144);
nor U8418 (N_8418,N_8334,N_8152);
and U8419 (N_8419,N_8353,N_8158);
and U8420 (N_8420,N_8241,N_8376);
nor U8421 (N_8421,N_8248,N_8107);
nor U8422 (N_8422,N_8263,N_8361);
nor U8423 (N_8423,N_8106,N_8272);
or U8424 (N_8424,N_8200,N_8378);
nor U8425 (N_8425,N_8126,N_8357);
and U8426 (N_8426,N_8129,N_8275);
or U8427 (N_8427,N_8292,N_8123);
and U8428 (N_8428,N_8336,N_8316);
xor U8429 (N_8429,N_8229,N_8383);
nor U8430 (N_8430,N_8135,N_8173);
xnor U8431 (N_8431,N_8290,N_8312);
nor U8432 (N_8432,N_8385,N_8117);
and U8433 (N_8433,N_8370,N_8104);
xor U8434 (N_8434,N_8184,N_8190);
nor U8435 (N_8435,N_8182,N_8395);
nor U8436 (N_8436,N_8354,N_8273);
nand U8437 (N_8437,N_8388,N_8114);
and U8438 (N_8438,N_8320,N_8198);
nand U8439 (N_8439,N_8191,N_8259);
nor U8440 (N_8440,N_8118,N_8307);
and U8441 (N_8441,N_8225,N_8193);
or U8442 (N_8442,N_8221,N_8270);
nand U8443 (N_8443,N_8319,N_8178);
nand U8444 (N_8444,N_8101,N_8345);
nor U8445 (N_8445,N_8318,N_8257);
nor U8446 (N_8446,N_8236,N_8209);
xnor U8447 (N_8447,N_8360,N_8341);
and U8448 (N_8448,N_8365,N_8244);
nand U8449 (N_8449,N_8186,N_8322);
nand U8450 (N_8450,N_8137,N_8296);
nand U8451 (N_8451,N_8167,N_8102);
xor U8452 (N_8452,N_8340,N_8288);
nor U8453 (N_8453,N_8251,N_8188);
and U8454 (N_8454,N_8181,N_8311);
xnor U8455 (N_8455,N_8304,N_8148);
and U8456 (N_8456,N_8195,N_8313);
xnor U8457 (N_8457,N_8155,N_8299);
xor U8458 (N_8458,N_8367,N_8177);
and U8459 (N_8459,N_8103,N_8342);
or U8460 (N_8460,N_8339,N_8151);
and U8461 (N_8461,N_8287,N_8331);
nand U8462 (N_8462,N_8143,N_8274);
xor U8463 (N_8463,N_8232,N_8344);
xor U8464 (N_8464,N_8206,N_8224);
nand U8465 (N_8465,N_8279,N_8175);
and U8466 (N_8466,N_8210,N_8303);
and U8467 (N_8467,N_8192,N_8223);
xor U8468 (N_8468,N_8194,N_8346);
xor U8469 (N_8469,N_8390,N_8214);
and U8470 (N_8470,N_8141,N_8302);
and U8471 (N_8471,N_8282,N_8127);
or U8472 (N_8472,N_8351,N_8147);
and U8473 (N_8473,N_8134,N_8396);
nand U8474 (N_8474,N_8108,N_8309);
and U8475 (N_8475,N_8199,N_8115);
nor U8476 (N_8476,N_8185,N_8163);
or U8477 (N_8477,N_8154,N_8119);
xnor U8478 (N_8478,N_8222,N_8249);
or U8479 (N_8479,N_8391,N_8169);
nor U8480 (N_8480,N_8364,N_8384);
nand U8481 (N_8481,N_8314,N_8113);
nand U8482 (N_8482,N_8255,N_8124);
xor U8483 (N_8483,N_8277,N_8258);
nand U8484 (N_8484,N_8271,N_8289);
nand U8485 (N_8485,N_8105,N_8269);
xnor U8486 (N_8486,N_8161,N_8176);
or U8487 (N_8487,N_8397,N_8197);
or U8488 (N_8488,N_8382,N_8399);
xor U8489 (N_8489,N_8347,N_8324);
xnor U8490 (N_8490,N_8350,N_8368);
nand U8491 (N_8491,N_8122,N_8363);
xor U8492 (N_8492,N_8305,N_8254);
or U8493 (N_8493,N_8233,N_8323);
xor U8494 (N_8494,N_8373,N_8179);
or U8495 (N_8495,N_8374,N_8130);
nand U8496 (N_8496,N_8146,N_8283);
nor U8497 (N_8497,N_8377,N_8189);
nor U8498 (N_8498,N_8329,N_8170);
nor U8499 (N_8499,N_8261,N_8264);
nand U8500 (N_8500,N_8393,N_8280);
xor U8501 (N_8501,N_8327,N_8293);
nand U8502 (N_8502,N_8260,N_8145);
and U8503 (N_8503,N_8235,N_8300);
and U8504 (N_8504,N_8375,N_8110);
and U8505 (N_8505,N_8136,N_8394);
or U8506 (N_8506,N_8218,N_8125);
nand U8507 (N_8507,N_8153,N_8359);
or U8508 (N_8508,N_8243,N_8208);
xnor U8509 (N_8509,N_8285,N_8203);
xor U8510 (N_8510,N_8398,N_8196);
and U8511 (N_8511,N_8253,N_8308);
xor U8512 (N_8512,N_8326,N_8216);
or U8513 (N_8513,N_8291,N_8139);
xnor U8514 (N_8514,N_8294,N_8234);
nor U8515 (N_8515,N_8369,N_8286);
xor U8516 (N_8516,N_8220,N_8160);
nand U8517 (N_8517,N_8239,N_8230);
or U8518 (N_8518,N_8298,N_8201);
nor U8519 (N_8519,N_8372,N_8306);
or U8520 (N_8520,N_8278,N_8109);
and U8521 (N_8521,N_8166,N_8157);
xor U8522 (N_8522,N_8310,N_8256);
nand U8523 (N_8523,N_8212,N_8267);
nor U8524 (N_8524,N_8321,N_8240);
nand U8525 (N_8525,N_8171,N_8133);
and U8526 (N_8526,N_8335,N_8281);
and U8527 (N_8527,N_8100,N_8227);
xor U8528 (N_8528,N_8156,N_8317);
xor U8529 (N_8529,N_8159,N_8121);
xnor U8530 (N_8530,N_8338,N_8325);
and U8531 (N_8531,N_8276,N_8266);
xor U8532 (N_8532,N_8172,N_8140);
and U8533 (N_8533,N_8284,N_8219);
and U8534 (N_8534,N_8128,N_8112);
nand U8535 (N_8535,N_8247,N_8228);
and U8536 (N_8536,N_8332,N_8348);
nor U8537 (N_8537,N_8252,N_8268);
and U8538 (N_8538,N_8204,N_8315);
nand U8539 (N_8539,N_8207,N_8352);
or U8540 (N_8540,N_8355,N_8356);
or U8541 (N_8541,N_8387,N_8168);
or U8542 (N_8542,N_8132,N_8116);
nor U8543 (N_8543,N_8250,N_8131);
or U8544 (N_8544,N_8162,N_8392);
xnor U8545 (N_8545,N_8381,N_8362);
xnor U8546 (N_8546,N_8149,N_8174);
nor U8547 (N_8547,N_8205,N_8150);
or U8548 (N_8548,N_8349,N_8111);
nor U8549 (N_8549,N_8142,N_8226);
or U8550 (N_8550,N_8285,N_8217);
or U8551 (N_8551,N_8144,N_8317);
or U8552 (N_8552,N_8226,N_8235);
and U8553 (N_8553,N_8256,N_8262);
nor U8554 (N_8554,N_8226,N_8186);
and U8555 (N_8555,N_8254,N_8396);
and U8556 (N_8556,N_8248,N_8262);
xor U8557 (N_8557,N_8279,N_8398);
or U8558 (N_8558,N_8257,N_8135);
nor U8559 (N_8559,N_8158,N_8101);
or U8560 (N_8560,N_8302,N_8369);
xnor U8561 (N_8561,N_8110,N_8322);
xnor U8562 (N_8562,N_8337,N_8133);
xor U8563 (N_8563,N_8343,N_8384);
nor U8564 (N_8564,N_8273,N_8312);
nor U8565 (N_8565,N_8131,N_8255);
and U8566 (N_8566,N_8121,N_8227);
or U8567 (N_8567,N_8166,N_8266);
and U8568 (N_8568,N_8101,N_8295);
and U8569 (N_8569,N_8112,N_8270);
and U8570 (N_8570,N_8362,N_8278);
or U8571 (N_8571,N_8140,N_8353);
xnor U8572 (N_8572,N_8137,N_8204);
and U8573 (N_8573,N_8318,N_8153);
and U8574 (N_8574,N_8356,N_8196);
xnor U8575 (N_8575,N_8310,N_8286);
or U8576 (N_8576,N_8342,N_8308);
and U8577 (N_8577,N_8107,N_8176);
xor U8578 (N_8578,N_8171,N_8279);
nor U8579 (N_8579,N_8201,N_8232);
xnor U8580 (N_8580,N_8373,N_8129);
nand U8581 (N_8581,N_8239,N_8193);
xnor U8582 (N_8582,N_8162,N_8280);
xor U8583 (N_8583,N_8114,N_8303);
or U8584 (N_8584,N_8264,N_8204);
nor U8585 (N_8585,N_8169,N_8320);
nor U8586 (N_8586,N_8331,N_8378);
or U8587 (N_8587,N_8390,N_8229);
and U8588 (N_8588,N_8320,N_8332);
and U8589 (N_8589,N_8160,N_8133);
and U8590 (N_8590,N_8151,N_8235);
xnor U8591 (N_8591,N_8249,N_8133);
nand U8592 (N_8592,N_8148,N_8272);
and U8593 (N_8593,N_8358,N_8200);
xnor U8594 (N_8594,N_8225,N_8348);
or U8595 (N_8595,N_8127,N_8200);
or U8596 (N_8596,N_8307,N_8349);
xor U8597 (N_8597,N_8175,N_8322);
nor U8598 (N_8598,N_8317,N_8373);
or U8599 (N_8599,N_8348,N_8134);
nand U8600 (N_8600,N_8148,N_8170);
and U8601 (N_8601,N_8253,N_8266);
xnor U8602 (N_8602,N_8114,N_8309);
xor U8603 (N_8603,N_8161,N_8273);
xor U8604 (N_8604,N_8319,N_8246);
xor U8605 (N_8605,N_8134,N_8323);
nor U8606 (N_8606,N_8135,N_8365);
xor U8607 (N_8607,N_8125,N_8300);
nand U8608 (N_8608,N_8197,N_8370);
and U8609 (N_8609,N_8218,N_8138);
nand U8610 (N_8610,N_8375,N_8283);
nor U8611 (N_8611,N_8137,N_8241);
nor U8612 (N_8612,N_8296,N_8339);
nand U8613 (N_8613,N_8219,N_8178);
nor U8614 (N_8614,N_8386,N_8236);
xnor U8615 (N_8615,N_8269,N_8117);
nor U8616 (N_8616,N_8276,N_8190);
or U8617 (N_8617,N_8124,N_8106);
or U8618 (N_8618,N_8189,N_8387);
nand U8619 (N_8619,N_8142,N_8337);
or U8620 (N_8620,N_8167,N_8278);
nor U8621 (N_8621,N_8169,N_8135);
xor U8622 (N_8622,N_8201,N_8375);
and U8623 (N_8623,N_8306,N_8198);
nor U8624 (N_8624,N_8363,N_8387);
and U8625 (N_8625,N_8304,N_8190);
nand U8626 (N_8626,N_8210,N_8128);
xor U8627 (N_8627,N_8221,N_8210);
nand U8628 (N_8628,N_8120,N_8102);
and U8629 (N_8629,N_8303,N_8138);
and U8630 (N_8630,N_8249,N_8134);
xnor U8631 (N_8631,N_8366,N_8237);
or U8632 (N_8632,N_8338,N_8346);
nor U8633 (N_8633,N_8126,N_8374);
nand U8634 (N_8634,N_8329,N_8125);
and U8635 (N_8635,N_8220,N_8122);
or U8636 (N_8636,N_8282,N_8129);
or U8637 (N_8637,N_8325,N_8220);
nor U8638 (N_8638,N_8395,N_8345);
nand U8639 (N_8639,N_8210,N_8352);
nand U8640 (N_8640,N_8124,N_8200);
and U8641 (N_8641,N_8278,N_8376);
and U8642 (N_8642,N_8116,N_8192);
and U8643 (N_8643,N_8301,N_8146);
and U8644 (N_8644,N_8287,N_8382);
xnor U8645 (N_8645,N_8132,N_8191);
nor U8646 (N_8646,N_8246,N_8345);
and U8647 (N_8647,N_8163,N_8176);
and U8648 (N_8648,N_8389,N_8284);
nor U8649 (N_8649,N_8178,N_8165);
or U8650 (N_8650,N_8276,N_8169);
xor U8651 (N_8651,N_8139,N_8288);
and U8652 (N_8652,N_8311,N_8355);
and U8653 (N_8653,N_8244,N_8121);
xor U8654 (N_8654,N_8262,N_8372);
or U8655 (N_8655,N_8121,N_8233);
nand U8656 (N_8656,N_8275,N_8380);
nor U8657 (N_8657,N_8158,N_8310);
xor U8658 (N_8658,N_8135,N_8145);
nand U8659 (N_8659,N_8267,N_8381);
or U8660 (N_8660,N_8276,N_8141);
nor U8661 (N_8661,N_8282,N_8333);
nand U8662 (N_8662,N_8115,N_8163);
nand U8663 (N_8663,N_8324,N_8137);
and U8664 (N_8664,N_8248,N_8300);
nand U8665 (N_8665,N_8198,N_8310);
nor U8666 (N_8666,N_8170,N_8101);
or U8667 (N_8667,N_8297,N_8114);
nor U8668 (N_8668,N_8349,N_8232);
xnor U8669 (N_8669,N_8307,N_8372);
nor U8670 (N_8670,N_8133,N_8398);
nor U8671 (N_8671,N_8378,N_8264);
nand U8672 (N_8672,N_8310,N_8368);
xor U8673 (N_8673,N_8270,N_8182);
xor U8674 (N_8674,N_8293,N_8136);
or U8675 (N_8675,N_8381,N_8320);
nand U8676 (N_8676,N_8161,N_8174);
nand U8677 (N_8677,N_8216,N_8264);
xor U8678 (N_8678,N_8269,N_8350);
and U8679 (N_8679,N_8233,N_8385);
nor U8680 (N_8680,N_8188,N_8215);
and U8681 (N_8681,N_8112,N_8152);
xor U8682 (N_8682,N_8335,N_8203);
xor U8683 (N_8683,N_8341,N_8356);
nor U8684 (N_8684,N_8189,N_8104);
or U8685 (N_8685,N_8255,N_8309);
nand U8686 (N_8686,N_8301,N_8360);
xor U8687 (N_8687,N_8302,N_8112);
and U8688 (N_8688,N_8138,N_8284);
nor U8689 (N_8689,N_8100,N_8163);
nor U8690 (N_8690,N_8287,N_8301);
and U8691 (N_8691,N_8278,N_8242);
nand U8692 (N_8692,N_8230,N_8252);
nor U8693 (N_8693,N_8143,N_8392);
xor U8694 (N_8694,N_8183,N_8108);
and U8695 (N_8695,N_8167,N_8195);
nand U8696 (N_8696,N_8381,N_8352);
nor U8697 (N_8697,N_8279,N_8150);
and U8698 (N_8698,N_8213,N_8158);
and U8699 (N_8699,N_8104,N_8206);
or U8700 (N_8700,N_8534,N_8687);
or U8701 (N_8701,N_8644,N_8626);
nor U8702 (N_8702,N_8500,N_8567);
nand U8703 (N_8703,N_8630,N_8596);
xor U8704 (N_8704,N_8527,N_8550);
and U8705 (N_8705,N_8420,N_8469);
xor U8706 (N_8706,N_8425,N_8546);
xnor U8707 (N_8707,N_8681,N_8521);
xnor U8708 (N_8708,N_8647,N_8522);
nor U8709 (N_8709,N_8504,N_8502);
xnor U8710 (N_8710,N_8653,N_8435);
xnor U8711 (N_8711,N_8665,N_8624);
nor U8712 (N_8712,N_8456,N_8528);
and U8713 (N_8713,N_8542,N_8417);
nor U8714 (N_8714,N_8478,N_8498);
xnor U8715 (N_8715,N_8675,N_8558);
and U8716 (N_8716,N_8471,N_8676);
xor U8717 (N_8717,N_8451,N_8540);
xnor U8718 (N_8718,N_8688,N_8605);
xor U8719 (N_8719,N_8621,N_8453);
xor U8720 (N_8720,N_8685,N_8447);
nand U8721 (N_8721,N_8679,N_8496);
xnor U8722 (N_8722,N_8423,N_8610);
and U8723 (N_8723,N_8559,N_8578);
and U8724 (N_8724,N_8422,N_8401);
and U8725 (N_8725,N_8466,N_8672);
nand U8726 (N_8726,N_8432,N_8510);
nand U8727 (N_8727,N_8636,N_8455);
or U8728 (N_8728,N_8538,N_8523);
and U8729 (N_8729,N_8557,N_8622);
and U8730 (N_8730,N_8639,N_8406);
or U8731 (N_8731,N_8571,N_8565);
nand U8732 (N_8732,N_8428,N_8494);
or U8733 (N_8733,N_8572,N_8629);
nand U8734 (N_8734,N_8674,N_8650);
nand U8735 (N_8735,N_8634,N_8547);
nor U8736 (N_8736,N_8461,N_8400);
nor U8737 (N_8737,N_8553,N_8412);
xor U8738 (N_8738,N_8439,N_8529);
nand U8739 (N_8739,N_8591,N_8448);
xnor U8740 (N_8740,N_8518,N_8491);
and U8741 (N_8741,N_8515,N_8641);
nor U8742 (N_8742,N_8444,N_8609);
or U8743 (N_8743,N_8600,N_8590);
xor U8744 (N_8744,N_8696,N_8457);
nor U8745 (N_8745,N_8489,N_8427);
nor U8746 (N_8746,N_8541,N_8415);
xnor U8747 (N_8747,N_8651,N_8564);
xnor U8748 (N_8748,N_8555,N_8434);
xnor U8749 (N_8749,N_8530,N_8450);
nand U8750 (N_8750,N_8483,N_8459);
nand U8751 (N_8751,N_8440,N_8535);
xor U8752 (N_8752,N_8648,N_8631);
xor U8753 (N_8753,N_8536,N_8470);
and U8754 (N_8754,N_8479,N_8566);
or U8755 (N_8755,N_8689,N_8511);
or U8756 (N_8756,N_8671,N_8620);
and U8757 (N_8757,N_8556,N_8577);
or U8758 (N_8758,N_8418,N_8413);
nand U8759 (N_8759,N_8508,N_8582);
nand U8760 (N_8760,N_8516,N_8431);
xnor U8761 (N_8761,N_8691,N_8580);
or U8762 (N_8762,N_8560,N_8658);
nor U8763 (N_8763,N_8669,N_8492);
nor U8764 (N_8764,N_8680,N_8467);
xor U8765 (N_8765,N_8454,N_8437);
nand U8766 (N_8766,N_8632,N_8585);
nor U8767 (N_8767,N_8597,N_8402);
or U8768 (N_8768,N_8615,N_8652);
or U8769 (N_8769,N_8524,N_8633);
nor U8770 (N_8770,N_8586,N_8677);
xor U8771 (N_8771,N_8568,N_8646);
nor U8772 (N_8772,N_8552,N_8592);
xnor U8773 (N_8773,N_8458,N_8690);
and U8774 (N_8774,N_8659,N_8573);
nand U8775 (N_8775,N_8551,N_8404);
nand U8776 (N_8776,N_8561,N_8668);
nand U8777 (N_8777,N_8537,N_8581);
or U8778 (N_8778,N_8576,N_8410);
and U8779 (N_8779,N_8525,N_8611);
xor U8780 (N_8780,N_8664,N_8649);
or U8781 (N_8781,N_8436,N_8548);
xor U8782 (N_8782,N_8438,N_8589);
nand U8783 (N_8783,N_8682,N_8429);
nor U8784 (N_8784,N_8424,N_8554);
xnor U8785 (N_8785,N_8487,N_8638);
nor U8786 (N_8786,N_8619,N_8468);
nand U8787 (N_8787,N_8512,N_8628);
and U8788 (N_8788,N_8587,N_8407);
and U8789 (N_8789,N_8416,N_8403);
nor U8790 (N_8790,N_8627,N_8505);
or U8791 (N_8791,N_8497,N_8462);
nor U8792 (N_8792,N_8488,N_8694);
or U8793 (N_8793,N_8699,N_8563);
and U8794 (N_8794,N_8613,N_8618);
nand U8795 (N_8795,N_8623,N_8442);
or U8796 (N_8796,N_8670,N_8408);
and U8797 (N_8797,N_8607,N_8520);
and U8798 (N_8798,N_8692,N_8608);
or U8799 (N_8799,N_8421,N_8643);
or U8800 (N_8800,N_8472,N_8562);
nor U8801 (N_8801,N_8584,N_8441);
xor U8802 (N_8802,N_8477,N_8601);
xor U8803 (N_8803,N_8635,N_8539);
nor U8804 (N_8804,N_8655,N_8549);
nand U8805 (N_8805,N_8452,N_8603);
xnor U8806 (N_8806,N_8476,N_8493);
xor U8807 (N_8807,N_8532,N_8485);
xor U8808 (N_8808,N_8593,N_8693);
nand U8809 (N_8809,N_8463,N_8663);
nor U8810 (N_8810,N_8545,N_8486);
nand U8811 (N_8811,N_8499,N_8490);
and U8812 (N_8812,N_8509,N_8574);
nor U8813 (N_8813,N_8446,N_8517);
xnor U8814 (N_8814,N_8484,N_8506);
nor U8815 (N_8815,N_8598,N_8531);
xnor U8816 (N_8816,N_8503,N_8433);
and U8817 (N_8817,N_8698,N_8657);
nand U8818 (N_8818,N_8579,N_8570);
nor U8819 (N_8819,N_8612,N_8495);
xor U8820 (N_8820,N_8678,N_8661);
nor U8821 (N_8821,N_8475,N_8697);
nand U8822 (N_8822,N_8637,N_8599);
or U8823 (N_8823,N_8606,N_8686);
nand U8824 (N_8824,N_8617,N_8465);
and U8825 (N_8825,N_8544,N_8480);
nor U8826 (N_8826,N_8667,N_8684);
nand U8827 (N_8827,N_8513,N_8588);
nand U8828 (N_8828,N_8662,N_8474);
nand U8829 (N_8829,N_8501,N_8449);
or U8830 (N_8830,N_8656,N_8583);
nand U8831 (N_8831,N_8519,N_8543);
nor U8832 (N_8832,N_8464,N_8411);
or U8833 (N_8833,N_8673,N_8604);
nor U8834 (N_8834,N_8595,N_8481);
and U8835 (N_8835,N_8614,N_8645);
and U8836 (N_8836,N_8660,N_8683);
or U8837 (N_8837,N_8695,N_8533);
xor U8838 (N_8838,N_8602,N_8514);
xnor U8839 (N_8839,N_8426,N_8482);
nand U8840 (N_8840,N_8473,N_8409);
nand U8841 (N_8841,N_8405,N_8445);
nor U8842 (N_8842,N_8430,N_8616);
or U8843 (N_8843,N_8419,N_8640);
nor U8844 (N_8844,N_8625,N_8594);
and U8845 (N_8845,N_8654,N_8666);
or U8846 (N_8846,N_8460,N_8642);
nand U8847 (N_8847,N_8414,N_8526);
nor U8848 (N_8848,N_8569,N_8507);
and U8849 (N_8849,N_8575,N_8443);
or U8850 (N_8850,N_8509,N_8429);
and U8851 (N_8851,N_8573,N_8699);
nor U8852 (N_8852,N_8517,N_8439);
or U8853 (N_8853,N_8474,N_8683);
or U8854 (N_8854,N_8422,N_8614);
or U8855 (N_8855,N_8643,N_8688);
or U8856 (N_8856,N_8525,N_8670);
and U8857 (N_8857,N_8645,N_8499);
xor U8858 (N_8858,N_8563,N_8543);
xnor U8859 (N_8859,N_8488,N_8470);
or U8860 (N_8860,N_8698,N_8533);
xor U8861 (N_8861,N_8550,N_8586);
nand U8862 (N_8862,N_8542,N_8649);
nand U8863 (N_8863,N_8539,N_8677);
and U8864 (N_8864,N_8587,N_8459);
nor U8865 (N_8865,N_8434,N_8690);
nand U8866 (N_8866,N_8568,N_8642);
and U8867 (N_8867,N_8588,N_8516);
xor U8868 (N_8868,N_8602,N_8470);
nor U8869 (N_8869,N_8528,N_8540);
xnor U8870 (N_8870,N_8472,N_8406);
nand U8871 (N_8871,N_8644,N_8485);
or U8872 (N_8872,N_8460,N_8496);
nand U8873 (N_8873,N_8680,N_8634);
nor U8874 (N_8874,N_8669,N_8652);
or U8875 (N_8875,N_8544,N_8408);
and U8876 (N_8876,N_8691,N_8615);
nor U8877 (N_8877,N_8449,N_8464);
and U8878 (N_8878,N_8486,N_8516);
and U8879 (N_8879,N_8645,N_8404);
xor U8880 (N_8880,N_8597,N_8687);
or U8881 (N_8881,N_8674,N_8414);
nand U8882 (N_8882,N_8620,N_8608);
nor U8883 (N_8883,N_8400,N_8514);
xor U8884 (N_8884,N_8498,N_8544);
xnor U8885 (N_8885,N_8566,N_8526);
nor U8886 (N_8886,N_8573,N_8642);
and U8887 (N_8887,N_8651,N_8474);
and U8888 (N_8888,N_8431,N_8440);
or U8889 (N_8889,N_8562,N_8527);
xnor U8890 (N_8890,N_8605,N_8552);
xnor U8891 (N_8891,N_8520,N_8507);
xnor U8892 (N_8892,N_8442,N_8669);
xor U8893 (N_8893,N_8567,N_8476);
nand U8894 (N_8894,N_8540,N_8534);
nand U8895 (N_8895,N_8571,N_8516);
nand U8896 (N_8896,N_8579,N_8419);
and U8897 (N_8897,N_8445,N_8550);
nand U8898 (N_8898,N_8493,N_8514);
and U8899 (N_8899,N_8640,N_8408);
xnor U8900 (N_8900,N_8503,N_8598);
nand U8901 (N_8901,N_8577,N_8609);
nor U8902 (N_8902,N_8642,N_8636);
nand U8903 (N_8903,N_8578,N_8522);
or U8904 (N_8904,N_8549,N_8609);
xor U8905 (N_8905,N_8693,N_8513);
nor U8906 (N_8906,N_8422,N_8444);
nand U8907 (N_8907,N_8663,N_8640);
and U8908 (N_8908,N_8499,N_8546);
nand U8909 (N_8909,N_8444,N_8558);
nand U8910 (N_8910,N_8568,N_8464);
xor U8911 (N_8911,N_8669,N_8612);
and U8912 (N_8912,N_8425,N_8628);
nor U8913 (N_8913,N_8579,N_8505);
and U8914 (N_8914,N_8493,N_8448);
or U8915 (N_8915,N_8582,N_8695);
and U8916 (N_8916,N_8467,N_8462);
and U8917 (N_8917,N_8693,N_8432);
nand U8918 (N_8918,N_8545,N_8410);
and U8919 (N_8919,N_8660,N_8435);
nor U8920 (N_8920,N_8641,N_8570);
xnor U8921 (N_8921,N_8633,N_8435);
or U8922 (N_8922,N_8642,N_8508);
nand U8923 (N_8923,N_8430,N_8470);
nor U8924 (N_8924,N_8480,N_8486);
or U8925 (N_8925,N_8502,N_8584);
and U8926 (N_8926,N_8598,N_8688);
and U8927 (N_8927,N_8551,N_8453);
xor U8928 (N_8928,N_8487,N_8504);
and U8929 (N_8929,N_8441,N_8565);
or U8930 (N_8930,N_8632,N_8572);
nand U8931 (N_8931,N_8603,N_8482);
or U8932 (N_8932,N_8546,N_8420);
nor U8933 (N_8933,N_8597,N_8541);
nor U8934 (N_8934,N_8696,N_8421);
and U8935 (N_8935,N_8472,N_8627);
xnor U8936 (N_8936,N_8593,N_8607);
xor U8937 (N_8937,N_8665,N_8642);
or U8938 (N_8938,N_8498,N_8411);
nand U8939 (N_8939,N_8406,N_8648);
or U8940 (N_8940,N_8617,N_8528);
or U8941 (N_8941,N_8612,N_8464);
nand U8942 (N_8942,N_8599,N_8536);
or U8943 (N_8943,N_8633,N_8657);
or U8944 (N_8944,N_8634,N_8441);
or U8945 (N_8945,N_8624,N_8692);
nand U8946 (N_8946,N_8685,N_8517);
and U8947 (N_8947,N_8552,N_8556);
nand U8948 (N_8948,N_8492,N_8680);
nand U8949 (N_8949,N_8691,N_8678);
and U8950 (N_8950,N_8697,N_8467);
xor U8951 (N_8951,N_8518,N_8634);
nor U8952 (N_8952,N_8673,N_8549);
and U8953 (N_8953,N_8686,N_8456);
and U8954 (N_8954,N_8570,N_8678);
nor U8955 (N_8955,N_8445,N_8534);
nand U8956 (N_8956,N_8641,N_8651);
and U8957 (N_8957,N_8634,N_8695);
nand U8958 (N_8958,N_8628,N_8576);
nor U8959 (N_8959,N_8511,N_8525);
xor U8960 (N_8960,N_8644,N_8691);
and U8961 (N_8961,N_8483,N_8590);
and U8962 (N_8962,N_8512,N_8401);
and U8963 (N_8963,N_8499,N_8511);
nand U8964 (N_8964,N_8495,N_8522);
and U8965 (N_8965,N_8576,N_8517);
nor U8966 (N_8966,N_8649,N_8608);
and U8967 (N_8967,N_8502,N_8620);
xor U8968 (N_8968,N_8576,N_8468);
xnor U8969 (N_8969,N_8433,N_8637);
and U8970 (N_8970,N_8539,N_8554);
and U8971 (N_8971,N_8432,N_8486);
nand U8972 (N_8972,N_8575,N_8507);
xnor U8973 (N_8973,N_8683,N_8484);
xor U8974 (N_8974,N_8659,N_8407);
or U8975 (N_8975,N_8669,N_8516);
xnor U8976 (N_8976,N_8585,N_8536);
xnor U8977 (N_8977,N_8541,N_8652);
and U8978 (N_8978,N_8577,N_8603);
nor U8979 (N_8979,N_8627,N_8643);
and U8980 (N_8980,N_8530,N_8659);
nand U8981 (N_8981,N_8506,N_8623);
and U8982 (N_8982,N_8696,N_8476);
xor U8983 (N_8983,N_8403,N_8624);
and U8984 (N_8984,N_8552,N_8442);
nand U8985 (N_8985,N_8403,N_8580);
nand U8986 (N_8986,N_8583,N_8652);
nor U8987 (N_8987,N_8646,N_8400);
nor U8988 (N_8988,N_8652,N_8516);
nor U8989 (N_8989,N_8562,N_8585);
and U8990 (N_8990,N_8408,N_8552);
and U8991 (N_8991,N_8437,N_8450);
nand U8992 (N_8992,N_8409,N_8615);
nand U8993 (N_8993,N_8411,N_8539);
nand U8994 (N_8994,N_8624,N_8545);
or U8995 (N_8995,N_8668,N_8509);
and U8996 (N_8996,N_8548,N_8475);
xor U8997 (N_8997,N_8463,N_8448);
nor U8998 (N_8998,N_8471,N_8503);
nor U8999 (N_8999,N_8463,N_8498);
nor U9000 (N_9000,N_8948,N_8716);
nand U9001 (N_9001,N_8781,N_8753);
nand U9002 (N_9002,N_8715,N_8998);
nor U9003 (N_9003,N_8944,N_8936);
nand U9004 (N_9004,N_8794,N_8768);
xor U9005 (N_9005,N_8783,N_8995);
nand U9006 (N_9006,N_8991,N_8876);
or U9007 (N_9007,N_8916,N_8928);
or U9008 (N_9008,N_8717,N_8772);
and U9009 (N_9009,N_8754,N_8925);
nor U9010 (N_9010,N_8725,N_8774);
or U9011 (N_9011,N_8858,N_8735);
or U9012 (N_9012,N_8723,N_8872);
or U9013 (N_9013,N_8849,N_8844);
xnor U9014 (N_9014,N_8977,N_8831);
nor U9015 (N_9015,N_8911,N_8862);
xor U9016 (N_9016,N_8714,N_8878);
xnor U9017 (N_9017,N_8953,N_8861);
or U9018 (N_9018,N_8792,N_8852);
xnor U9019 (N_9019,N_8799,N_8760);
or U9020 (N_9020,N_8898,N_8939);
nor U9021 (N_9021,N_8788,N_8963);
and U9022 (N_9022,N_8839,N_8938);
or U9023 (N_9023,N_8947,N_8810);
or U9024 (N_9024,N_8825,N_8842);
and U9025 (N_9025,N_8943,N_8732);
or U9026 (N_9026,N_8880,N_8869);
or U9027 (N_9027,N_8934,N_8802);
or U9028 (N_9028,N_8736,N_8897);
or U9029 (N_9029,N_8919,N_8988);
and U9030 (N_9030,N_8976,N_8950);
or U9031 (N_9031,N_8859,N_8865);
xnor U9032 (N_9032,N_8955,N_8730);
nor U9033 (N_9033,N_8803,N_8968);
xnor U9034 (N_9034,N_8720,N_8741);
and U9035 (N_9035,N_8800,N_8728);
nand U9036 (N_9036,N_8881,N_8931);
nor U9037 (N_9037,N_8771,N_8910);
and U9038 (N_9038,N_8961,N_8906);
or U9039 (N_9039,N_8796,N_8874);
nor U9040 (N_9040,N_8932,N_8914);
and U9041 (N_9041,N_8752,N_8808);
and U9042 (N_9042,N_8873,N_8828);
xor U9043 (N_9043,N_8763,N_8882);
and U9044 (N_9044,N_8710,N_8727);
nand U9045 (N_9045,N_8922,N_8855);
and U9046 (N_9046,N_8787,N_8966);
and U9047 (N_9047,N_8731,N_8890);
or U9048 (N_9048,N_8702,N_8801);
nor U9049 (N_9049,N_8795,N_8896);
xor U9050 (N_9050,N_8889,N_8982);
xor U9051 (N_9051,N_8811,N_8983);
and U9052 (N_9052,N_8912,N_8979);
or U9053 (N_9053,N_8821,N_8952);
and U9054 (N_9054,N_8917,N_8751);
xor U9055 (N_9055,N_8959,N_8846);
and U9056 (N_9056,N_8822,N_8770);
or U9057 (N_9057,N_8851,N_8778);
nor U9058 (N_9058,N_8969,N_8761);
and U9059 (N_9059,N_8806,N_8818);
and U9060 (N_9060,N_8824,N_8784);
nor U9061 (N_9061,N_8709,N_8701);
nor U9062 (N_9062,N_8738,N_8981);
xor U9063 (N_9063,N_8962,N_8960);
and U9064 (N_9064,N_8815,N_8848);
and U9065 (N_9065,N_8777,N_8748);
nor U9066 (N_9066,N_8989,N_8786);
xor U9067 (N_9067,N_8994,N_8779);
or U9068 (N_9068,N_8703,N_8719);
xor U9069 (N_9069,N_8903,N_8762);
nor U9070 (N_9070,N_8870,N_8765);
xnor U9071 (N_9071,N_8984,N_8750);
nand U9072 (N_9072,N_8899,N_8957);
nand U9073 (N_9073,N_8775,N_8860);
nand U9074 (N_9074,N_8879,N_8904);
nand U9075 (N_9075,N_8758,N_8909);
xor U9076 (N_9076,N_8740,N_8764);
nor U9077 (N_9077,N_8713,N_8940);
xor U9078 (N_9078,N_8743,N_8813);
nor U9079 (N_9079,N_8893,N_8926);
or U9080 (N_9080,N_8868,N_8745);
nor U9081 (N_9081,N_8864,N_8837);
and U9082 (N_9082,N_8964,N_8812);
and U9083 (N_9083,N_8990,N_8830);
xor U9084 (N_9084,N_8946,N_8974);
or U9085 (N_9085,N_8773,N_8835);
nand U9086 (N_9086,N_8907,N_8744);
nor U9087 (N_9087,N_8978,N_8722);
nor U9088 (N_9088,N_8833,N_8883);
xnor U9089 (N_9089,N_8954,N_8756);
xnor U9090 (N_9090,N_8742,N_8843);
nor U9091 (N_9091,N_8973,N_8853);
xor U9092 (N_9092,N_8877,N_8992);
xnor U9093 (N_9093,N_8769,N_8980);
or U9094 (N_9094,N_8965,N_8757);
or U9095 (N_9095,N_8705,N_8700);
nand U9096 (N_9096,N_8891,N_8967);
or U9097 (N_9097,N_8749,N_8892);
and U9098 (N_9098,N_8739,N_8886);
xnor U9099 (N_9099,N_8905,N_8704);
xor U9100 (N_9100,N_8708,N_8945);
and U9101 (N_9101,N_8817,N_8999);
xor U9102 (N_9102,N_8805,N_8724);
and U9103 (N_9103,N_8820,N_8885);
and U9104 (N_9104,N_8789,N_8985);
and U9105 (N_9105,N_8942,N_8930);
xnor U9106 (N_9106,N_8941,N_8819);
and U9107 (N_9107,N_8987,N_8780);
and U9108 (N_9108,N_8733,N_8734);
or U9109 (N_9109,N_8863,N_8921);
and U9110 (N_9110,N_8901,N_8793);
or U9111 (N_9111,N_8997,N_8827);
nand U9112 (N_9112,N_8900,N_8856);
nand U9113 (N_9113,N_8949,N_8746);
xnor U9114 (N_9114,N_8816,N_8721);
nor U9115 (N_9115,N_8785,N_8841);
nor U9116 (N_9116,N_8838,N_8993);
and U9117 (N_9117,N_8804,N_8767);
or U9118 (N_9118,N_8923,N_8755);
xor U9119 (N_9119,N_8927,N_8809);
nand U9120 (N_9120,N_8894,N_8867);
or U9121 (N_9121,N_8970,N_8951);
and U9122 (N_9122,N_8823,N_8986);
nor U9123 (N_9123,N_8924,N_8902);
nor U9124 (N_9124,N_8706,N_8797);
or U9125 (N_9125,N_8711,N_8747);
xnor U9126 (N_9126,N_8972,N_8791);
nor U9127 (N_9127,N_8840,N_8790);
nand U9128 (N_9128,N_8845,N_8908);
nand U9129 (N_9129,N_8834,N_8798);
nand U9130 (N_9130,N_8975,N_8888);
nand U9131 (N_9131,N_8935,N_8895);
nand U9132 (N_9132,N_8996,N_8920);
nor U9133 (N_9133,N_8836,N_8875);
and U9134 (N_9134,N_8971,N_8726);
and U9135 (N_9135,N_8937,N_8854);
and U9136 (N_9136,N_8766,N_8866);
or U9137 (N_9137,N_8956,N_8776);
xor U9138 (N_9138,N_8832,N_8884);
and U9139 (N_9139,N_8871,N_8918);
nor U9140 (N_9140,N_8887,N_8707);
or U9141 (N_9141,N_8850,N_8782);
nor U9142 (N_9142,N_8814,N_8929);
or U9143 (N_9143,N_8729,N_8915);
nor U9144 (N_9144,N_8712,N_8826);
and U9145 (N_9145,N_8857,N_8829);
nor U9146 (N_9146,N_8913,N_8847);
or U9147 (N_9147,N_8718,N_8933);
nor U9148 (N_9148,N_8807,N_8759);
or U9149 (N_9149,N_8958,N_8737);
xnor U9150 (N_9150,N_8780,N_8895);
and U9151 (N_9151,N_8881,N_8964);
nand U9152 (N_9152,N_8767,N_8910);
nand U9153 (N_9153,N_8775,N_8939);
and U9154 (N_9154,N_8840,N_8797);
and U9155 (N_9155,N_8908,N_8911);
nand U9156 (N_9156,N_8988,N_8821);
nor U9157 (N_9157,N_8995,N_8725);
xor U9158 (N_9158,N_8880,N_8736);
nor U9159 (N_9159,N_8985,N_8876);
nand U9160 (N_9160,N_8768,N_8755);
and U9161 (N_9161,N_8897,N_8859);
or U9162 (N_9162,N_8816,N_8894);
or U9163 (N_9163,N_8717,N_8926);
or U9164 (N_9164,N_8949,N_8792);
nand U9165 (N_9165,N_8781,N_8712);
xnor U9166 (N_9166,N_8863,N_8890);
and U9167 (N_9167,N_8927,N_8832);
nand U9168 (N_9168,N_8953,N_8952);
nand U9169 (N_9169,N_8816,N_8702);
nor U9170 (N_9170,N_8958,N_8701);
xor U9171 (N_9171,N_8894,N_8963);
xor U9172 (N_9172,N_8713,N_8741);
and U9173 (N_9173,N_8884,N_8978);
nor U9174 (N_9174,N_8905,N_8934);
xnor U9175 (N_9175,N_8808,N_8938);
and U9176 (N_9176,N_8718,N_8703);
xnor U9177 (N_9177,N_8900,N_8714);
and U9178 (N_9178,N_8896,N_8931);
and U9179 (N_9179,N_8890,N_8802);
nor U9180 (N_9180,N_8936,N_8935);
xor U9181 (N_9181,N_8773,N_8860);
xor U9182 (N_9182,N_8812,N_8813);
nand U9183 (N_9183,N_8900,N_8767);
or U9184 (N_9184,N_8759,N_8980);
and U9185 (N_9185,N_8784,N_8838);
or U9186 (N_9186,N_8895,N_8759);
nor U9187 (N_9187,N_8966,N_8837);
xnor U9188 (N_9188,N_8833,N_8805);
nor U9189 (N_9189,N_8864,N_8993);
xor U9190 (N_9190,N_8919,N_8805);
and U9191 (N_9191,N_8725,N_8756);
or U9192 (N_9192,N_8727,N_8734);
nor U9193 (N_9193,N_8740,N_8804);
nor U9194 (N_9194,N_8969,N_8729);
and U9195 (N_9195,N_8979,N_8920);
xor U9196 (N_9196,N_8920,N_8974);
nor U9197 (N_9197,N_8710,N_8792);
or U9198 (N_9198,N_8836,N_8864);
nand U9199 (N_9199,N_8886,N_8875);
or U9200 (N_9200,N_8869,N_8979);
nor U9201 (N_9201,N_8925,N_8913);
xnor U9202 (N_9202,N_8879,N_8778);
xor U9203 (N_9203,N_8876,N_8907);
or U9204 (N_9204,N_8741,N_8962);
nand U9205 (N_9205,N_8750,N_8916);
and U9206 (N_9206,N_8784,N_8748);
xor U9207 (N_9207,N_8882,N_8924);
xnor U9208 (N_9208,N_8827,N_8835);
nor U9209 (N_9209,N_8972,N_8845);
xnor U9210 (N_9210,N_8824,N_8973);
or U9211 (N_9211,N_8978,N_8721);
xor U9212 (N_9212,N_8799,N_8906);
or U9213 (N_9213,N_8869,N_8718);
or U9214 (N_9214,N_8947,N_8973);
or U9215 (N_9215,N_8937,N_8955);
and U9216 (N_9216,N_8744,N_8817);
nand U9217 (N_9217,N_8885,N_8849);
and U9218 (N_9218,N_8943,N_8720);
and U9219 (N_9219,N_8759,N_8865);
nand U9220 (N_9220,N_8866,N_8813);
nand U9221 (N_9221,N_8768,N_8821);
xnor U9222 (N_9222,N_8709,N_8936);
and U9223 (N_9223,N_8800,N_8903);
xnor U9224 (N_9224,N_8751,N_8910);
nand U9225 (N_9225,N_8895,N_8948);
and U9226 (N_9226,N_8975,N_8771);
nor U9227 (N_9227,N_8737,N_8812);
xnor U9228 (N_9228,N_8823,N_8765);
and U9229 (N_9229,N_8883,N_8767);
and U9230 (N_9230,N_8916,N_8851);
or U9231 (N_9231,N_8706,N_8898);
and U9232 (N_9232,N_8969,N_8747);
nand U9233 (N_9233,N_8949,N_8824);
and U9234 (N_9234,N_8886,N_8703);
and U9235 (N_9235,N_8864,N_8961);
nand U9236 (N_9236,N_8933,N_8917);
nand U9237 (N_9237,N_8947,N_8976);
nand U9238 (N_9238,N_8811,N_8862);
and U9239 (N_9239,N_8800,N_8836);
nor U9240 (N_9240,N_8880,N_8814);
nor U9241 (N_9241,N_8920,N_8933);
and U9242 (N_9242,N_8995,N_8894);
and U9243 (N_9243,N_8904,N_8962);
xor U9244 (N_9244,N_8735,N_8913);
or U9245 (N_9245,N_8774,N_8919);
nor U9246 (N_9246,N_8973,N_8797);
nand U9247 (N_9247,N_8714,N_8832);
and U9248 (N_9248,N_8827,N_8766);
and U9249 (N_9249,N_8704,N_8783);
and U9250 (N_9250,N_8798,N_8980);
nor U9251 (N_9251,N_8888,N_8914);
and U9252 (N_9252,N_8997,N_8744);
or U9253 (N_9253,N_8739,N_8971);
xor U9254 (N_9254,N_8900,N_8742);
and U9255 (N_9255,N_8807,N_8787);
and U9256 (N_9256,N_8728,N_8732);
xor U9257 (N_9257,N_8854,N_8891);
xor U9258 (N_9258,N_8943,N_8960);
and U9259 (N_9259,N_8886,N_8988);
xor U9260 (N_9260,N_8862,N_8832);
nand U9261 (N_9261,N_8843,N_8958);
nor U9262 (N_9262,N_8738,N_8749);
xnor U9263 (N_9263,N_8740,N_8835);
nand U9264 (N_9264,N_8856,N_8843);
nand U9265 (N_9265,N_8923,N_8713);
nor U9266 (N_9266,N_8840,N_8868);
nor U9267 (N_9267,N_8875,N_8850);
and U9268 (N_9268,N_8717,N_8732);
or U9269 (N_9269,N_8788,N_8967);
xor U9270 (N_9270,N_8773,N_8713);
or U9271 (N_9271,N_8856,N_8721);
nand U9272 (N_9272,N_8816,N_8810);
and U9273 (N_9273,N_8776,N_8889);
nor U9274 (N_9274,N_8905,N_8966);
nand U9275 (N_9275,N_8834,N_8931);
and U9276 (N_9276,N_8731,N_8814);
nor U9277 (N_9277,N_8828,N_8955);
nor U9278 (N_9278,N_8910,N_8873);
nand U9279 (N_9279,N_8873,N_8813);
and U9280 (N_9280,N_8839,N_8738);
xor U9281 (N_9281,N_8848,N_8755);
and U9282 (N_9282,N_8757,N_8833);
xnor U9283 (N_9283,N_8942,N_8997);
nor U9284 (N_9284,N_8871,N_8754);
and U9285 (N_9285,N_8885,N_8745);
or U9286 (N_9286,N_8824,N_8875);
or U9287 (N_9287,N_8888,N_8989);
and U9288 (N_9288,N_8950,N_8925);
xnor U9289 (N_9289,N_8775,N_8886);
nand U9290 (N_9290,N_8704,N_8748);
and U9291 (N_9291,N_8997,N_8701);
nor U9292 (N_9292,N_8723,N_8816);
xor U9293 (N_9293,N_8723,N_8935);
xnor U9294 (N_9294,N_8702,N_8913);
nand U9295 (N_9295,N_8823,N_8778);
nor U9296 (N_9296,N_8880,N_8898);
nor U9297 (N_9297,N_8908,N_8838);
xnor U9298 (N_9298,N_8874,N_8711);
nand U9299 (N_9299,N_8726,N_8909);
and U9300 (N_9300,N_9120,N_9148);
nand U9301 (N_9301,N_9095,N_9143);
or U9302 (N_9302,N_9176,N_9062);
or U9303 (N_9303,N_9007,N_9249);
xnor U9304 (N_9304,N_9023,N_9052);
nand U9305 (N_9305,N_9213,N_9097);
or U9306 (N_9306,N_9051,N_9247);
xnor U9307 (N_9307,N_9260,N_9156);
nor U9308 (N_9308,N_9183,N_9189);
and U9309 (N_9309,N_9179,N_9286);
or U9310 (N_9310,N_9207,N_9118);
or U9311 (N_9311,N_9230,N_9240);
xor U9312 (N_9312,N_9231,N_9108);
nand U9313 (N_9313,N_9164,N_9098);
nor U9314 (N_9314,N_9026,N_9194);
nor U9315 (N_9315,N_9001,N_9208);
or U9316 (N_9316,N_9281,N_9129);
nor U9317 (N_9317,N_9201,N_9025);
xor U9318 (N_9318,N_9227,N_9091);
and U9319 (N_9319,N_9288,N_9252);
xor U9320 (N_9320,N_9024,N_9153);
or U9321 (N_9321,N_9071,N_9033);
and U9322 (N_9322,N_9109,N_9256);
and U9323 (N_9323,N_9119,N_9042);
or U9324 (N_9324,N_9152,N_9168);
or U9325 (N_9325,N_9180,N_9289);
nand U9326 (N_9326,N_9293,N_9170);
nor U9327 (N_9327,N_9002,N_9149);
nand U9328 (N_9328,N_9094,N_9057);
nand U9329 (N_9329,N_9237,N_9268);
nor U9330 (N_9330,N_9248,N_9200);
and U9331 (N_9331,N_9244,N_9271);
xnor U9332 (N_9332,N_9262,N_9267);
and U9333 (N_9333,N_9137,N_9117);
nor U9334 (N_9334,N_9299,N_9020);
or U9335 (N_9335,N_9018,N_9241);
and U9336 (N_9336,N_9130,N_9246);
nand U9337 (N_9337,N_9048,N_9272);
nand U9338 (N_9338,N_9245,N_9151);
or U9339 (N_9339,N_9031,N_9105);
and U9340 (N_9340,N_9250,N_9228);
xnor U9341 (N_9341,N_9043,N_9212);
xnor U9342 (N_9342,N_9177,N_9236);
and U9343 (N_9343,N_9096,N_9150);
nand U9344 (N_9344,N_9113,N_9006);
nand U9345 (N_9345,N_9093,N_9044);
nand U9346 (N_9346,N_9079,N_9187);
xnor U9347 (N_9347,N_9142,N_9285);
or U9348 (N_9348,N_9069,N_9084);
nor U9349 (N_9349,N_9054,N_9169);
xor U9350 (N_9350,N_9279,N_9166);
or U9351 (N_9351,N_9263,N_9182);
xnor U9352 (N_9352,N_9221,N_9190);
nand U9353 (N_9353,N_9253,N_9283);
and U9354 (N_9354,N_9021,N_9292);
xnor U9355 (N_9355,N_9030,N_9013);
nand U9356 (N_9356,N_9234,N_9211);
and U9357 (N_9357,N_9005,N_9100);
or U9358 (N_9358,N_9010,N_9046);
nand U9359 (N_9359,N_9214,N_9009);
and U9360 (N_9360,N_9178,N_9027);
or U9361 (N_9361,N_9217,N_9242);
xnor U9362 (N_9362,N_9273,N_9000);
xor U9363 (N_9363,N_9114,N_9162);
nor U9364 (N_9364,N_9070,N_9146);
xnor U9365 (N_9365,N_9274,N_9188);
nand U9366 (N_9366,N_9039,N_9101);
or U9367 (N_9367,N_9073,N_9160);
nand U9368 (N_9368,N_9063,N_9123);
or U9369 (N_9369,N_9019,N_9254);
nor U9370 (N_9370,N_9127,N_9135);
nand U9371 (N_9371,N_9204,N_9064);
nor U9372 (N_9372,N_9011,N_9269);
nor U9373 (N_9373,N_9259,N_9068);
nor U9374 (N_9374,N_9131,N_9297);
nand U9375 (N_9375,N_9028,N_9255);
nor U9376 (N_9376,N_9277,N_9161);
and U9377 (N_9377,N_9174,N_9203);
xor U9378 (N_9378,N_9050,N_9053);
xor U9379 (N_9379,N_9004,N_9121);
and U9380 (N_9380,N_9290,N_9072);
or U9381 (N_9381,N_9229,N_9016);
xnor U9382 (N_9382,N_9076,N_9157);
xor U9383 (N_9383,N_9196,N_9088);
nand U9384 (N_9384,N_9215,N_9115);
xnor U9385 (N_9385,N_9251,N_9265);
xnor U9386 (N_9386,N_9029,N_9116);
or U9387 (N_9387,N_9257,N_9047);
nand U9388 (N_9388,N_9078,N_9243);
or U9389 (N_9389,N_9139,N_9282);
and U9390 (N_9390,N_9081,N_9163);
nand U9391 (N_9391,N_9102,N_9173);
or U9392 (N_9392,N_9099,N_9124);
nand U9393 (N_9393,N_9056,N_9141);
nor U9394 (N_9394,N_9270,N_9083);
or U9395 (N_9395,N_9291,N_9296);
nor U9396 (N_9396,N_9167,N_9144);
nor U9397 (N_9397,N_9037,N_9138);
and U9398 (N_9398,N_9090,N_9125);
nor U9399 (N_9399,N_9239,N_9035);
or U9400 (N_9400,N_9206,N_9225);
nand U9401 (N_9401,N_9014,N_9086);
and U9402 (N_9402,N_9181,N_9038);
and U9403 (N_9403,N_9036,N_9295);
nor U9404 (N_9404,N_9159,N_9220);
or U9405 (N_9405,N_9110,N_9205);
and U9406 (N_9406,N_9085,N_9233);
nor U9407 (N_9407,N_9055,N_9219);
or U9408 (N_9408,N_9165,N_9154);
and U9409 (N_9409,N_9216,N_9195);
or U9410 (N_9410,N_9104,N_9107);
nor U9411 (N_9411,N_9080,N_9075);
and U9412 (N_9412,N_9092,N_9103);
nand U9413 (N_9413,N_9122,N_9186);
nor U9414 (N_9414,N_9278,N_9155);
and U9415 (N_9415,N_9238,N_9012);
and U9416 (N_9416,N_9022,N_9275);
nor U9417 (N_9417,N_9222,N_9202);
nor U9418 (N_9418,N_9049,N_9128);
or U9419 (N_9419,N_9032,N_9066);
nand U9420 (N_9420,N_9264,N_9112);
xnor U9421 (N_9421,N_9224,N_9133);
nand U9422 (N_9422,N_9077,N_9126);
xor U9423 (N_9423,N_9218,N_9034);
nand U9424 (N_9424,N_9145,N_9067);
and U9425 (N_9425,N_9106,N_9040);
xor U9426 (N_9426,N_9223,N_9284);
nand U9427 (N_9427,N_9061,N_9197);
nand U9428 (N_9428,N_9210,N_9136);
or U9429 (N_9429,N_9172,N_9059);
nor U9430 (N_9430,N_9258,N_9082);
xor U9431 (N_9431,N_9132,N_9232);
or U9432 (N_9432,N_9226,N_9158);
xor U9433 (N_9433,N_9045,N_9276);
nor U9434 (N_9434,N_9191,N_9185);
nor U9435 (N_9435,N_9175,N_9147);
nor U9436 (N_9436,N_9171,N_9287);
and U9437 (N_9437,N_9111,N_9294);
or U9438 (N_9438,N_9003,N_9074);
and U9439 (N_9439,N_9134,N_9266);
nor U9440 (N_9440,N_9199,N_9087);
nor U9441 (N_9441,N_9065,N_9017);
xnor U9442 (N_9442,N_9015,N_9235);
nand U9443 (N_9443,N_9184,N_9198);
xor U9444 (N_9444,N_9298,N_9008);
and U9445 (N_9445,N_9193,N_9261);
xnor U9446 (N_9446,N_9209,N_9058);
xnor U9447 (N_9447,N_9140,N_9089);
nor U9448 (N_9448,N_9280,N_9041);
xnor U9449 (N_9449,N_9060,N_9192);
or U9450 (N_9450,N_9239,N_9225);
nor U9451 (N_9451,N_9039,N_9024);
or U9452 (N_9452,N_9269,N_9240);
and U9453 (N_9453,N_9072,N_9067);
nand U9454 (N_9454,N_9053,N_9111);
and U9455 (N_9455,N_9050,N_9207);
xnor U9456 (N_9456,N_9298,N_9260);
and U9457 (N_9457,N_9133,N_9056);
nand U9458 (N_9458,N_9290,N_9124);
xor U9459 (N_9459,N_9083,N_9268);
nand U9460 (N_9460,N_9238,N_9015);
nand U9461 (N_9461,N_9240,N_9097);
xor U9462 (N_9462,N_9085,N_9192);
xor U9463 (N_9463,N_9252,N_9011);
and U9464 (N_9464,N_9103,N_9063);
nand U9465 (N_9465,N_9142,N_9224);
or U9466 (N_9466,N_9270,N_9200);
xor U9467 (N_9467,N_9298,N_9225);
and U9468 (N_9468,N_9246,N_9161);
and U9469 (N_9469,N_9095,N_9027);
nand U9470 (N_9470,N_9027,N_9276);
and U9471 (N_9471,N_9054,N_9296);
and U9472 (N_9472,N_9109,N_9026);
nor U9473 (N_9473,N_9272,N_9279);
nor U9474 (N_9474,N_9050,N_9219);
or U9475 (N_9475,N_9118,N_9089);
and U9476 (N_9476,N_9163,N_9047);
xor U9477 (N_9477,N_9187,N_9239);
nor U9478 (N_9478,N_9168,N_9142);
nor U9479 (N_9479,N_9073,N_9148);
nand U9480 (N_9480,N_9031,N_9123);
xnor U9481 (N_9481,N_9135,N_9161);
nand U9482 (N_9482,N_9131,N_9226);
nand U9483 (N_9483,N_9138,N_9211);
xor U9484 (N_9484,N_9077,N_9244);
xor U9485 (N_9485,N_9230,N_9034);
and U9486 (N_9486,N_9208,N_9093);
or U9487 (N_9487,N_9178,N_9144);
or U9488 (N_9488,N_9046,N_9281);
or U9489 (N_9489,N_9140,N_9228);
nand U9490 (N_9490,N_9110,N_9241);
xor U9491 (N_9491,N_9255,N_9151);
xor U9492 (N_9492,N_9021,N_9269);
or U9493 (N_9493,N_9200,N_9218);
nor U9494 (N_9494,N_9153,N_9151);
nor U9495 (N_9495,N_9075,N_9100);
nand U9496 (N_9496,N_9230,N_9165);
xnor U9497 (N_9497,N_9190,N_9098);
xor U9498 (N_9498,N_9237,N_9193);
nand U9499 (N_9499,N_9148,N_9215);
nand U9500 (N_9500,N_9195,N_9089);
or U9501 (N_9501,N_9058,N_9236);
or U9502 (N_9502,N_9015,N_9072);
or U9503 (N_9503,N_9054,N_9099);
or U9504 (N_9504,N_9110,N_9220);
and U9505 (N_9505,N_9020,N_9273);
nor U9506 (N_9506,N_9225,N_9080);
or U9507 (N_9507,N_9081,N_9284);
nor U9508 (N_9508,N_9273,N_9260);
xor U9509 (N_9509,N_9121,N_9035);
xnor U9510 (N_9510,N_9227,N_9225);
nand U9511 (N_9511,N_9047,N_9023);
or U9512 (N_9512,N_9201,N_9092);
and U9513 (N_9513,N_9079,N_9274);
nor U9514 (N_9514,N_9021,N_9024);
nor U9515 (N_9515,N_9204,N_9059);
xor U9516 (N_9516,N_9059,N_9146);
nor U9517 (N_9517,N_9088,N_9099);
nor U9518 (N_9518,N_9108,N_9063);
nor U9519 (N_9519,N_9226,N_9094);
xor U9520 (N_9520,N_9161,N_9056);
nand U9521 (N_9521,N_9012,N_9045);
or U9522 (N_9522,N_9146,N_9152);
nand U9523 (N_9523,N_9017,N_9213);
nor U9524 (N_9524,N_9275,N_9067);
or U9525 (N_9525,N_9118,N_9295);
xor U9526 (N_9526,N_9157,N_9056);
nor U9527 (N_9527,N_9276,N_9048);
xnor U9528 (N_9528,N_9271,N_9230);
and U9529 (N_9529,N_9223,N_9035);
nor U9530 (N_9530,N_9070,N_9266);
nor U9531 (N_9531,N_9253,N_9298);
nand U9532 (N_9532,N_9274,N_9262);
nand U9533 (N_9533,N_9016,N_9291);
and U9534 (N_9534,N_9129,N_9216);
or U9535 (N_9535,N_9120,N_9033);
and U9536 (N_9536,N_9151,N_9100);
nor U9537 (N_9537,N_9272,N_9297);
nor U9538 (N_9538,N_9199,N_9116);
or U9539 (N_9539,N_9227,N_9023);
or U9540 (N_9540,N_9169,N_9120);
nor U9541 (N_9541,N_9110,N_9169);
xor U9542 (N_9542,N_9225,N_9218);
or U9543 (N_9543,N_9098,N_9020);
or U9544 (N_9544,N_9216,N_9066);
or U9545 (N_9545,N_9250,N_9138);
and U9546 (N_9546,N_9205,N_9149);
nor U9547 (N_9547,N_9042,N_9069);
or U9548 (N_9548,N_9244,N_9224);
and U9549 (N_9549,N_9296,N_9114);
or U9550 (N_9550,N_9035,N_9090);
xnor U9551 (N_9551,N_9184,N_9125);
or U9552 (N_9552,N_9179,N_9161);
and U9553 (N_9553,N_9299,N_9263);
xnor U9554 (N_9554,N_9201,N_9200);
nor U9555 (N_9555,N_9238,N_9203);
or U9556 (N_9556,N_9218,N_9171);
xnor U9557 (N_9557,N_9173,N_9051);
and U9558 (N_9558,N_9184,N_9032);
xnor U9559 (N_9559,N_9282,N_9075);
nor U9560 (N_9560,N_9204,N_9153);
or U9561 (N_9561,N_9191,N_9042);
nor U9562 (N_9562,N_9190,N_9242);
nand U9563 (N_9563,N_9223,N_9048);
or U9564 (N_9564,N_9223,N_9078);
nand U9565 (N_9565,N_9072,N_9171);
or U9566 (N_9566,N_9068,N_9152);
nand U9567 (N_9567,N_9202,N_9110);
and U9568 (N_9568,N_9291,N_9198);
and U9569 (N_9569,N_9260,N_9146);
nor U9570 (N_9570,N_9101,N_9108);
and U9571 (N_9571,N_9041,N_9236);
xnor U9572 (N_9572,N_9017,N_9037);
or U9573 (N_9573,N_9251,N_9232);
nand U9574 (N_9574,N_9187,N_9167);
and U9575 (N_9575,N_9204,N_9250);
nand U9576 (N_9576,N_9289,N_9061);
nor U9577 (N_9577,N_9057,N_9166);
or U9578 (N_9578,N_9160,N_9106);
or U9579 (N_9579,N_9241,N_9010);
nand U9580 (N_9580,N_9193,N_9130);
xor U9581 (N_9581,N_9121,N_9211);
and U9582 (N_9582,N_9282,N_9000);
nor U9583 (N_9583,N_9167,N_9274);
nand U9584 (N_9584,N_9034,N_9044);
nor U9585 (N_9585,N_9174,N_9183);
nor U9586 (N_9586,N_9192,N_9187);
or U9587 (N_9587,N_9190,N_9071);
nor U9588 (N_9588,N_9166,N_9147);
or U9589 (N_9589,N_9036,N_9018);
and U9590 (N_9590,N_9257,N_9213);
and U9591 (N_9591,N_9217,N_9136);
nor U9592 (N_9592,N_9074,N_9120);
nand U9593 (N_9593,N_9096,N_9166);
and U9594 (N_9594,N_9232,N_9152);
or U9595 (N_9595,N_9010,N_9091);
nor U9596 (N_9596,N_9238,N_9270);
nor U9597 (N_9597,N_9274,N_9293);
nor U9598 (N_9598,N_9191,N_9205);
nor U9599 (N_9599,N_9277,N_9207);
and U9600 (N_9600,N_9525,N_9560);
nor U9601 (N_9601,N_9585,N_9402);
and U9602 (N_9602,N_9349,N_9414);
nand U9603 (N_9603,N_9377,N_9447);
and U9604 (N_9604,N_9527,N_9568);
xnor U9605 (N_9605,N_9347,N_9388);
and U9606 (N_9606,N_9567,N_9578);
xnor U9607 (N_9607,N_9301,N_9409);
or U9608 (N_9608,N_9463,N_9589);
or U9609 (N_9609,N_9330,N_9551);
xor U9610 (N_9610,N_9479,N_9577);
nand U9611 (N_9611,N_9472,N_9444);
and U9612 (N_9612,N_9488,N_9493);
xor U9613 (N_9613,N_9338,N_9405);
xor U9614 (N_9614,N_9441,N_9535);
xnor U9615 (N_9615,N_9449,N_9403);
xnor U9616 (N_9616,N_9462,N_9368);
nand U9617 (N_9617,N_9314,N_9324);
and U9618 (N_9618,N_9308,N_9571);
or U9619 (N_9619,N_9336,N_9302);
or U9620 (N_9620,N_9546,N_9573);
and U9621 (N_9621,N_9357,N_9473);
nand U9622 (N_9622,N_9307,N_9396);
and U9623 (N_9623,N_9412,N_9555);
or U9624 (N_9624,N_9325,N_9520);
xnor U9625 (N_9625,N_9529,N_9575);
xor U9626 (N_9626,N_9328,N_9430);
nand U9627 (N_9627,N_9598,N_9374);
and U9628 (N_9628,N_9394,N_9446);
and U9629 (N_9629,N_9508,N_9580);
xor U9630 (N_9630,N_9530,N_9310);
or U9631 (N_9631,N_9376,N_9491);
nor U9632 (N_9632,N_9389,N_9509);
and U9633 (N_9633,N_9458,N_9311);
xnor U9634 (N_9634,N_9465,N_9561);
nor U9635 (N_9635,N_9581,N_9417);
nor U9636 (N_9636,N_9553,N_9353);
nand U9637 (N_9637,N_9326,N_9574);
or U9638 (N_9638,N_9306,N_9536);
xor U9639 (N_9639,N_9316,N_9432);
nand U9640 (N_9640,N_9469,N_9411);
or U9641 (N_9641,N_9315,N_9386);
nand U9642 (N_9642,N_9434,N_9362);
nand U9643 (N_9643,N_9439,N_9399);
or U9644 (N_9644,N_9572,N_9387);
nor U9645 (N_9645,N_9378,N_9576);
nor U9646 (N_9646,N_9517,N_9312);
or U9647 (N_9647,N_9317,N_9437);
or U9648 (N_9648,N_9363,N_9429);
xor U9649 (N_9649,N_9321,N_9599);
nor U9650 (N_9650,N_9340,N_9329);
xnor U9651 (N_9651,N_9408,N_9595);
and U9652 (N_9652,N_9319,N_9483);
nand U9653 (N_9653,N_9523,N_9323);
and U9654 (N_9654,N_9550,N_9511);
nor U9655 (N_9655,N_9344,N_9442);
nor U9656 (N_9656,N_9327,N_9482);
or U9657 (N_9657,N_9369,N_9487);
nor U9658 (N_9658,N_9404,N_9359);
nor U9659 (N_9659,N_9440,N_9486);
nor U9660 (N_9660,N_9416,N_9365);
xnor U9661 (N_9661,N_9438,N_9342);
nand U9662 (N_9662,N_9503,N_9496);
or U9663 (N_9663,N_9562,N_9375);
or U9664 (N_9664,N_9521,N_9596);
nor U9665 (N_9665,N_9385,N_9395);
and U9666 (N_9666,N_9556,N_9500);
nor U9667 (N_9667,N_9569,N_9582);
nand U9668 (N_9668,N_9507,N_9380);
or U9669 (N_9669,N_9354,N_9498);
xor U9670 (N_9670,N_9304,N_9547);
xor U9671 (N_9671,N_9459,N_9300);
xor U9672 (N_9672,N_9345,N_9592);
xor U9673 (N_9673,N_9594,N_9322);
nor U9674 (N_9674,N_9502,N_9348);
or U9675 (N_9675,N_9542,N_9397);
and U9676 (N_9676,N_9370,N_9454);
or U9677 (N_9677,N_9460,N_9343);
nand U9678 (N_9678,N_9597,N_9457);
nor U9679 (N_9679,N_9515,N_9445);
or U9680 (N_9680,N_9383,N_9390);
xor U9681 (N_9681,N_9471,N_9320);
nor U9682 (N_9682,N_9522,N_9590);
xor U9683 (N_9683,N_9564,N_9335);
nand U9684 (N_9684,N_9528,N_9512);
nand U9685 (N_9685,N_9565,N_9514);
nand U9686 (N_9686,N_9519,N_9448);
xnor U9687 (N_9687,N_9540,N_9422);
xor U9688 (N_9688,N_9419,N_9524);
nor U9689 (N_9689,N_9333,N_9518);
nand U9690 (N_9690,N_9453,N_9526);
nand U9691 (N_9691,N_9570,N_9351);
nor U9692 (N_9692,N_9475,N_9464);
xnor U9693 (N_9693,N_9428,N_9421);
or U9694 (N_9694,N_9489,N_9309);
xnor U9695 (N_9695,N_9552,N_9485);
xnor U9696 (N_9696,N_9358,N_9513);
nor U9697 (N_9697,N_9346,N_9313);
or U9698 (N_9698,N_9398,N_9418);
nand U9699 (N_9699,N_9593,N_9558);
xnor U9700 (N_9700,N_9426,N_9533);
or U9701 (N_9701,N_9391,N_9364);
xor U9702 (N_9702,N_9548,N_9456);
or U9703 (N_9703,N_9505,N_9366);
nor U9704 (N_9704,N_9549,N_9531);
nand U9705 (N_9705,N_9379,N_9497);
and U9706 (N_9706,N_9337,N_9356);
nor U9707 (N_9707,N_9587,N_9490);
nand U9708 (N_9708,N_9455,N_9452);
xnor U9709 (N_9709,N_9367,N_9534);
xnor U9710 (N_9710,N_9318,N_9543);
nand U9711 (N_9711,N_9481,N_9478);
nor U9712 (N_9712,N_9371,N_9413);
xnor U9713 (N_9713,N_9360,N_9384);
nor U9714 (N_9714,N_9584,N_9433);
or U9715 (N_9715,N_9427,N_9545);
xor U9716 (N_9716,N_9516,N_9436);
or U9717 (N_9717,N_9420,N_9484);
or U9718 (N_9718,N_9537,N_9470);
or U9719 (N_9719,N_9466,N_9450);
or U9720 (N_9720,N_9476,N_9381);
nor U9721 (N_9721,N_9331,N_9423);
nand U9722 (N_9722,N_9332,N_9451);
or U9723 (N_9723,N_9382,N_9334);
nand U9724 (N_9724,N_9563,N_9393);
and U9725 (N_9725,N_9506,N_9443);
nand U9726 (N_9726,N_9372,N_9504);
and U9727 (N_9727,N_9435,N_9579);
nor U9728 (N_9728,N_9392,N_9559);
or U9729 (N_9729,N_9480,N_9554);
and U9730 (N_9730,N_9400,N_9494);
nor U9731 (N_9731,N_9499,N_9415);
nand U9732 (N_9732,N_9424,N_9361);
xnor U9733 (N_9733,N_9566,N_9468);
xnor U9734 (N_9734,N_9477,N_9583);
nand U9735 (N_9735,N_9350,N_9341);
nor U9736 (N_9736,N_9425,N_9591);
nand U9737 (N_9737,N_9305,N_9352);
and U9738 (N_9738,N_9339,N_9407);
nand U9739 (N_9739,N_9501,N_9539);
xnor U9740 (N_9740,N_9406,N_9588);
and U9741 (N_9741,N_9586,N_9355);
nor U9742 (N_9742,N_9557,N_9461);
or U9743 (N_9743,N_9532,N_9410);
or U9744 (N_9744,N_9541,N_9373);
or U9745 (N_9745,N_9510,N_9544);
or U9746 (N_9746,N_9538,N_9431);
or U9747 (N_9747,N_9467,N_9401);
xor U9748 (N_9748,N_9474,N_9495);
and U9749 (N_9749,N_9492,N_9303);
nor U9750 (N_9750,N_9461,N_9414);
xor U9751 (N_9751,N_9339,N_9496);
or U9752 (N_9752,N_9548,N_9589);
and U9753 (N_9753,N_9446,N_9567);
nor U9754 (N_9754,N_9471,N_9378);
and U9755 (N_9755,N_9322,N_9448);
and U9756 (N_9756,N_9524,N_9599);
nor U9757 (N_9757,N_9554,N_9422);
or U9758 (N_9758,N_9470,N_9332);
nand U9759 (N_9759,N_9400,N_9384);
or U9760 (N_9760,N_9565,N_9593);
nand U9761 (N_9761,N_9330,N_9301);
nand U9762 (N_9762,N_9402,N_9431);
xor U9763 (N_9763,N_9403,N_9453);
and U9764 (N_9764,N_9582,N_9309);
nor U9765 (N_9765,N_9503,N_9418);
nand U9766 (N_9766,N_9384,N_9430);
xor U9767 (N_9767,N_9427,N_9459);
xnor U9768 (N_9768,N_9454,N_9438);
xor U9769 (N_9769,N_9445,N_9516);
xor U9770 (N_9770,N_9318,N_9599);
xnor U9771 (N_9771,N_9575,N_9345);
nor U9772 (N_9772,N_9559,N_9542);
xnor U9773 (N_9773,N_9449,N_9490);
or U9774 (N_9774,N_9460,N_9584);
nor U9775 (N_9775,N_9365,N_9450);
or U9776 (N_9776,N_9381,N_9434);
or U9777 (N_9777,N_9433,N_9425);
and U9778 (N_9778,N_9493,N_9380);
and U9779 (N_9779,N_9392,N_9402);
xor U9780 (N_9780,N_9347,N_9569);
xnor U9781 (N_9781,N_9465,N_9582);
or U9782 (N_9782,N_9347,N_9533);
nand U9783 (N_9783,N_9355,N_9316);
xor U9784 (N_9784,N_9478,N_9346);
xnor U9785 (N_9785,N_9364,N_9305);
and U9786 (N_9786,N_9325,N_9598);
and U9787 (N_9787,N_9392,N_9581);
and U9788 (N_9788,N_9491,N_9351);
nor U9789 (N_9789,N_9460,N_9583);
xor U9790 (N_9790,N_9564,N_9397);
nand U9791 (N_9791,N_9351,N_9535);
and U9792 (N_9792,N_9542,N_9423);
or U9793 (N_9793,N_9405,N_9413);
nor U9794 (N_9794,N_9468,N_9527);
nor U9795 (N_9795,N_9577,N_9574);
nor U9796 (N_9796,N_9378,N_9362);
nand U9797 (N_9797,N_9340,N_9426);
xor U9798 (N_9798,N_9397,N_9483);
nand U9799 (N_9799,N_9467,N_9348);
or U9800 (N_9800,N_9390,N_9567);
and U9801 (N_9801,N_9347,N_9455);
and U9802 (N_9802,N_9407,N_9480);
nand U9803 (N_9803,N_9363,N_9444);
nand U9804 (N_9804,N_9384,N_9501);
and U9805 (N_9805,N_9485,N_9316);
nor U9806 (N_9806,N_9434,N_9492);
nor U9807 (N_9807,N_9569,N_9318);
or U9808 (N_9808,N_9438,N_9551);
and U9809 (N_9809,N_9308,N_9398);
xor U9810 (N_9810,N_9438,N_9404);
nand U9811 (N_9811,N_9483,N_9311);
xnor U9812 (N_9812,N_9512,N_9442);
and U9813 (N_9813,N_9565,N_9586);
or U9814 (N_9814,N_9410,N_9431);
xor U9815 (N_9815,N_9555,N_9494);
xor U9816 (N_9816,N_9434,N_9371);
or U9817 (N_9817,N_9375,N_9513);
nor U9818 (N_9818,N_9500,N_9399);
nor U9819 (N_9819,N_9575,N_9335);
and U9820 (N_9820,N_9507,N_9338);
nand U9821 (N_9821,N_9582,N_9391);
nor U9822 (N_9822,N_9349,N_9321);
nor U9823 (N_9823,N_9541,N_9340);
nor U9824 (N_9824,N_9514,N_9302);
nor U9825 (N_9825,N_9588,N_9538);
nor U9826 (N_9826,N_9333,N_9436);
nor U9827 (N_9827,N_9438,N_9479);
nor U9828 (N_9828,N_9494,N_9405);
and U9829 (N_9829,N_9300,N_9325);
nor U9830 (N_9830,N_9566,N_9549);
and U9831 (N_9831,N_9371,N_9461);
xor U9832 (N_9832,N_9565,N_9404);
nor U9833 (N_9833,N_9390,N_9325);
and U9834 (N_9834,N_9438,N_9582);
nand U9835 (N_9835,N_9453,N_9382);
nand U9836 (N_9836,N_9492,N_9431);
or U9837 (N_9837,N_9511,N_9491);
or U9838 (N_9838,N_9451,N_9402);
nand U9839 (N_9839,N_9480,N_9550);
xor U9840 (N_9840,N_9554,N_9304);
xor U9841 (N_9841,N_9577,N_9386);
and U9842 (N_9842,N_9349,N_9484);
xnor U9843 (N_9843,N_9542,N_9527);
nand U9844 (N_9844,N_9583,N_9401);
nand U9845 (N_9845,N_9592,N_9352);
nand U9846 (N_9846,N_9338,N_9456);
nand U9847 (N_9847,N_9524,N_9494);
nor U9848 (N_9848,N_9375,N_9487);
nand U9849 (N_9849,N_9350,N_9516);
xor U9850 (N_9850,N_9520,N_9446);
or U9851 (N_9851,N_9549,N_9526);
nor U9852 (N_9852,N_9499,N_9536);
nand U9853 (N_9853,N_9306,N_9433);
nand U9854 (N_9854,N_9536,N_9393);
or U9855 (N_9855,N_9599,N_9381);
xor U9856 (N_9856,N_9590,N_9441);
and U9857 (N_9857,N_9571,N_9326);
or U9858 (N_9858,N_9314,N_9446);
xor U9859 (N_9859,N_9359,N_9320);
or U9860 (N_9860,N_9478,N_9354);
xor U9861 (N_9861,N_9552,N_9557);
or U9862 (N_9862,N_9468,N_9367);
and U9863 (N_9863,N_9500,N_9448);
nor U9864 (N_9864,N_9363,N_9338);
nand U9865 (N_9865,N_9388,N_9527);
and U9866 (N_9866,N_9307,N_9301);
and U9867 (N_9867,N_9360,N_9373);
nor U9868 (N_9868,N_9316,N_9340);
and U9869 (N_9869,N_9528,N_9511);
nor U9870 (N_9870,N_9423,N_9488);
and U9871 (N_9871,N_9445,N_9319);
xor U9872 (N_9872,N_9482,N_9414);
nand U9873 (N_9873,N_9488,N_9378);
nand U9874 (N_9874,N_9328,N_9537);
nand U9875 (N_9875,N_9356,N_9427);
nand U9876 (N_9876,N_9497,N_9558);
nor U9877 (N_9877,N_9341,N_9505);
and U9878 (N_9878,N_9310,N_9483);
nor U9879 (N_9879,N_9522,N_9583);
nand U9880 (N_9880,N_9390,N_9439);
and U9881 (N_9881,N_9542,N_9491);
and U9882 (N_9882,N_9573,N_9404);
nand U9883 (N_9883,N_9354,N_9552);
and U9884 (N_9884,N_9542,N_9346);
and U9885 (N_9885,N_9301,N_9389);
and U9886 (N_9886,N_9470,N_9338);
and U9887 (N_9887,N_9362,N_9548);
nor U9888 (N_9888,N_9320,N_9313);
nand U9889 (N_9889,N_9365,N_9370);
or U9890 (N_9890,N_9348,N_9349);
nand U9891 (N_9891,N_9320,N_9333);
nor U9892 (N_9892,N_9386,N_9372);
nand U9893 (N_9893,N_9397,N_9378);
or U9894 (N_9894,N_9472,N_9528);
nor U9895 (N_9895,N_9522,N_9520);
nand U9896 (N_9896,N_9493,N_9592);
nand U9897 (N_9897,N_9319,N_9594);
nand U9898 (N_9898,N_9313,N_9581);
nand U9899 (N_9899,N_9481,N_9411);
and U9900 (N_9900,N_9739,N_9889);
nand U9901 (N_9901,N_9700,N_9804);
nand U9902 (N_9902,N_9668,N_9708);
and U9903 (N_9903,N_9705,N_9670);
nand U9904 (N_9904,N_9816,N_9740);
and U9905 (N_9905,N_9642,N_9659);
xor U9906 (N_9906,N_9701,N_9687);
or U9907 (N_9907,N_9666,N_9695);
and U9908 (N_9908,N_9824,N_9846);
or U9909 (N_9909,N_9671,N_9748);
nand U9910 (N_9910,N_9826,N_9607);
nor U9911 (N_9911,N_9820,N_9733);
nor U9912 (N_9912,N_9847,N_9604);
or U9913 (N_9913,N_9882,N_9858);
nor U9914 (N_9914,N_9602,N_9781);
nor U9915 (N_9915,N_9887,N_9864);
and U9916 (N_9916,N_9627,N_9843);
or U9917 (N_9917,N_9896,N_9807);
nand U9918 (N_9918,N_9694,N_9738);
nor U9919 (N_9919,N_9633,N_9663);
nand U9920 (N_9920,N_9646,N_9898);
nor U9921 (N_9921,N_9706,N_9788);
or U9922 (N_9922,N_9773,N_9692);
nand U9923 (N_9923,N_9874,N_9728);
nor U9924 (N_9924,N_9831,N_9769);
nor U9925 (N_9925,N_9845,N_9745);
xnor U9926 (N_9926,N_9619,N_9837);
and U9927 (N_9927,N_9762,N_9702);
nand U9928 (N_9928,N_9849,N_9703);
or U9929 (N_9929,N_9810,N_9871);
nand U9930 (N_9930,N_9654,N_9632);
or U9931 (N_9931,N_9696,N_9835);
nand U9932 (N_9932,N_9606,N_9852);
nor U9933 (N_9933,N_9774,N_9691);
xnor U9934 (N_9934,N_9658,N_9656);
and U9935 (N_9935,N_9634,N_9812);
or U9936 (N_9936,N_9746,N_9635);
nor U9937 (N_9937,N_9723,N_9711);
xor U9938 (N_9938,N_9661,N_9880);
and U9939 (N_9939,N_9648,N_9736);
nand U9940 (N_9940,N_9877,N_9712);
or U9941 (N_9941,N_9873,N_9870);
and U9942 (N_9942,N_9709,N_9787);
or U9943 (N_9943,N_9611,N_9894);
xor U9944 (N_9944,N_9792,N_9629);
xor U9945 (N_9945,N_9756,N_9662);
or U9946 (N_9946,N_9865,N_9672);
or U9947 (N_9947,N_9798,N_9718);
or U9948 (N_9948,N_9775,N_9675);
xor U9949 (N_9949,N_9893,N_9665);
nor U9950 (N_9950,N_9821,N_9717);
xor U9951 (N_9951,N_9651,N_9688);
nor U9952 (N_9952,N_9710,N_9803);
nor U9953 (N_9953,N_9797,N_9744);
or U9954 (N_9954,N_9737,N_9698);
or U9955 (N_9955,N_9653,N_9872);
nor U9956 (N_9956,N_9895,N_9725);
and U9957 (N_9957,N_9652,N_9650);
xor U9958 (N_9958,N_9776,N_9851);
xnor U9959 (N_9959,N_9763,N_9825);
or U9960 (N_9960,N_9639,N_9721);
or U9961 (N_9961,N_9897,N_9734);
nor U9962 (N_9962,N_9892,N_9809);
nor U9963 (N_9963,N_9795,N_9645);
xnor U9964 (N_9964,N_9743,N_9697);
nor U9965 (N_9965,N_9722,N_9778);
xnor U9966 (N_9966,N_9605,N_9680);
xor U9967 (N_9967,N_9890,N_9868);
and U9968 (N_9968,N_9750,N_9863);
nand U9969 (N_9969,N_9735,N_9823);
xnor U9970 (N_9970,N_9616,N_9626);
nor U9971 (N_9971,N_9764,N_9834);
or U9972 (N_9972,N_9747,N_9677);
xnor U9973 (N_9973,N_9855,N_9856);
or U9974 (N_9974,N_9817,N_9753);
or U9975 (N_9975,N_9789,N_9643);
and U9976 (N_9976,N_9741,N_9610);
nor U9977 (N_9977,N_9600,N_9660);
xor U9978 (N_9978,N_9609,N_9867);
and U9979 (N_9979,N_9777,N_9791);
nor U9980 (N_9980,N_9649,N_9640);
nand U9981 (N_9981,N_9881,N_9760);
xor U9982 (N_9982,N_9742,N_9844);
nand U9983 (N_9983,N_9714,N_9784);
or U9984 (N_9984,N_9876,N_9869);
nor U9985 (N_9985,N_9674,N_9815);
or U9986 (N_9986,N_9793,N_9805);
and U9987 (N_9987,N_9818,N_9765);
and U9988 (N_9988,N_9630,N_9664);
or U9989 (N_9989,N_9685,N_9785);
xnor U9990 (N_9990,N_9850,N_9879);
or U9991 (N_9991,N_9704,N_9608);
xor U9992 (N_9992,N_9836,N_9779);
nand U9993 (N_9993,N_9726,N_9848);
nand U9994 (N_9994,N_9832,N_9819);
and U9995 (N_9995,N_9814,N_9885);
xnor U9996 (N_9996,N_9782,N_9612);
nor U9997 (N_9997,N_9839,N_9647);
or U9998 (N_9998,N_9822,N_9716);
nand U9999 (N_9999,N_9636,N_9833);
or U10000 (N_10000,N_9759,N_9888);
xor U10001 (N_10001,N_9829,N_9799);
nor U10002 (N_10002,N_9808,N_9644);
nor U10003 (N_10003,N_9771,N_9842);
nor U10004 (N_10004,N_9669,N_9813);
xor U10005 (N_10005,N_9811,N_9638);
nand U10006 (N_10006,N_9853,N_9806);
or U10007 (N_10007,N_9783,N_9620);
or U10008 (N_10008,N_9875,N_9715);
or U10009 (N_10009,N_9631,N_9796);
nand U10010 (N_10010,N_9732,N_9621);
or U10011 (N_10011,N_9601,N_9752);
and U10012 (N_10012,N_9828,N_9690);
nor U10013 (N_10013,N_9625,N_9641);
or U10014 (N_10014,N_9628,N_9838);
nor U10015 (N_10015,N_9699,N_9801);
xnor U10016 (N_10016,N_9800,N_9724);
nor U10017 (N_10017,N_9755,N_9682);
nand U10018 (N_10018,N_9891,N_9772);
and U10019 (N_10019,N_9862,N_9827);
or U10020 (N_10020,N_9757,N_9766);
xor U10021 (N_10021,N_9857,N_9684);
nor U10022 (N_10022,N_9786,N_9866);
xor U10023 (N_10023,N_9693,N_9618);
and U10024 (N_10024,N_9758,N_9860);
and U10025 (N_10025,N_9720,N_9667);
xor U10026 (N_10026,N_9683,N_9861);
or U10027 (N_10027,N_9657,N_9730);
and U10028 (N_10028,N_9624,N_9617);
xnor U10029 (N_10029,N_9731,N_9727);
or U10030 (N_10030,N_9878,N_9729);
and U10031 (N_10031,N_9679,N_9754);
nand U10032 (N_10032,N_9719,N_9673);
nor U10033 (N_10033,N_9899,N_9707);
nor U10034 (N_10034,N_9761,N_9623);
and U10035 (N_10035,N_9686,N_9770);
nor U10036 (N_10036,N_9681,N_9767);
nand U10037 (N_10037,N_9622,N_9794);
nand U10038 (N_10038,N_9884,N_9859);
or U10039 (N_10039,N_9840,N_9676);
or U10040 (N_10040,N_9603,N_9637);
xnor U10041 (N_10041,N_9883,N_9749);
or U10042 (N_10042,N_9751,N_9614);
nand U10043 (N_10043,N_9613,N_9802);
and U10044 (N_10044,N_9830,N_9689);
nor U10045 (N_10045,N_9886,N_9678);
nor U10046 (N_10046,N_9780,N_9655);
nor U10047 (N_10047,N_9615,N_9854);
and U10048 (N_10048,N_9713,N_9768);
or U10049 (N_10049,N_9790,N_9841);
nor U10050 (N_10050,N_9738,N_9872);
or U10051 (N_10051,N_9656,N_9804);
nor U10052 (N_10052,N_9697,N_9877);
or U10053 (N_10053,N_9798,N_9843);
nor U10054 (N_10054,N_9789,N_9884);
and U10055 (N_10055,N_9866,N_9859);
nor U10056 (N_10056,N_9894,N_9792);
nor U10057 (N_10057,N_9738,N_9668);
and U10058 (N_10058,N_9868,N_9738);
and U10059 (N_10059,N_9770,N_9745);
nand U10060 (N_10060,N_9809,N_9701);
nand U10061 (N_10061,N_9754,N_9802);
or U10062 (N_10062,N_9816,N_9654);
nand U10063 (N_10063,N_9707,N_9788);
and U10064 (N_10064,N_9693,N_9867);
nand U10065 (N_10065,N_9648,N_9799);
xor U10066 (N_10066,N_9683,N_9866);
nor U10067 (N_10067,N_9883,N_9668);
nor U10068 (N_10068,N_9696,N_9885);
nor U10069 (N_10069,N_9825,N_9799);
and U10070 (N_10070,N_9774,N_9600);
nor U10071 (N_10071,N_9715,N_9783);
and U10072 (N_10072,N_9741,N_9849);
xor U10073 (N_10073,N_9845,N_9637);
nor U10074 (N_10074,N_9880,N_9797);
nand U10075 (N_10075,N_9881,N_9695);
and U10076 (N_10076,N_9639,N_9879);
nor U10077 (N_10077,N_9772,N_9854);
xnor U10078 (N_10078,N_9797,N_9897);
nand U10079 (N_10079,N_9603,N_9764);
xor U10080 (N_10080,N_9660,N_9758);
or U10081 (N_10081,N_9890,N_9775);
xor U10082 (N_10082,N_9830,N_9859);
nand U10083 (N_10083,N_9897,N_9854);
or U10084 (N_10084,N_9896,N_9623);
nor U10085 (N_10085,N_9691,N_9847);
or U10086 (N_10086,N_9633,N_9807);
and U10087 (N_10087,N_9650,N_9857);
and U10088 (N_10088,N_9869,N_9897);
nand U10089 (N_10089,N_9800,N_9623);
nor U10090 (N_10090,N_9619,N_9825);
xor U10091 (N_10091,N_9763,N_9645);
xor U10092 (N_10092,N_9765,N_9746);
nand U10093 (N_10093,N_9708,N_9752);
xor U10094 (N_10094,N_9605,N_9637);
or U10095 (N_10095,N_9605,N_9603);
xor U10096 (N_10096,N_9753,N_9814);
nor U10097 (N_10097,N_9725,N_9811);
or U10098 (N_10098,N_9744,N_9615);
or U10099 (N_10099,N_9875,N_9838);
nor U10100 (N_10100,N_9895,N_9704);
nand U10101 (N_10101,N_9890,N_9850);
xor U10102 (N_10102,N_9662,N_9747);
or U10103 (N_10103,N_9868,N_9641);
and U10104 (N_10104,N_9766,N_9876);
xnor U10105 (N_10105,N_9811,N_9662);
and U10106 (N_10106,N_9894,N_9630);
xnor U10107 (N_10107,N_9663,N_9898);
and U10108 (N_10108,N_9825,N_9623);
and U10109 (N_10109,N_9889,N_9888);
nand U10110 (N_10110,N_9615,N_9890);
nand U10111 (N_10111,N_9670,N_9600);
nand U10112 (N_10112,N_9632,N_9820);
and U10113 (N_10113,N_9774,N_9665);
nor U10114 (N_10114,N_9680,N_9690);
or U10115 (N_10115,N_9674,N_9753);
nor U10116 (N_10116,N_9643,N_9823);
or U10117 (N_10117,N_9725,N_9756);
xor U10118 (N_10118,N_9657,N_9658);
or U10119 (N_10119,N_9898,N_9702);
nand U10120 (N_10120,N_9774,N_9878);
nand U10121 (N_10121,N_9869,N_9808);
nand U10122 (N_10122,N_9690,N_9668);
nor U10123 (N_10123,N_9640,N_9645);
nor U10124 (N_10124,N_9713,N_9781);
and U10125 (N_10125,N_9759,N_9652);
nand U10126 (N_10126,N_9781,N_9823);
xnor U10127 (N_10127,N_9814,N_9730);
xnor U10128 (N_10128,N_9675,N_9754);
nand U10129 (N_10129,N_9795,N_9867);
and U10130 (N_10130,N_9715,N_9633);
nand U10131 (N_10131,N_9790,N_9607);
or U10132 (N_10132,N_9824,N_9665);
or U10133 (N_10133,N_9709,N_9765);
or U10134 (N_10134,N_9648,N_9644);
xor U10135 (N_10135,N_9809,N_9732);
or U10136 (N_10136,N_9667,N_9898);
and U10137 (N_10137,N_9876,N_9737);
nor U10138 (N_10138,N_9798,N_9647);
or U10139 (N_10139,N_9632,N_9613);
nor U10140 (N_10140,N_9704,N_9626);
xor U10141 (N_10141,N_9742,N_9805);
nor U10142 (N_10142,N_9607,N_9830);
and U10143 (N_10143,N_9692,N_9711);
xor U10144 (N_10144,N_9727,N_9712);
nor U10145 (N_10145,N_9692,N_9714);
and U10146 (N_10146,N_9686,N_9846);
or U10147 (N_10147,N_9686,N_9670);
and U10148 (N_10148,N_9883,N_9823);
nand U10149 (N_10149,N_9888,N_9611);
nor U10150 (N_10150,N_9723,N_9702);
nor U10151 (N_10151,N_9792,N_9884);
and U10152 (N_10152,N_9858,N_9837);
xnor U10153 (N_10153,N_9771,N_9758);
or U10154 (N_10154,N_9899,N_9877);
or U10155 (N_10155,N_9759,N_9805);
or U10156 (N_10156,N_9789,N_9684);
xnor U10157 (N_10157,N_9868,N_9721);
or U10158 (N_10158,N_9695,N_9785);
and U10159 (N_10159,N_9841,N_9897);
and U10160 (N_10160,N_9692,N_9650);
nand U10161 (N_10161,N_9890,N_9797);
and U10162 (N_10162,N_9817,N_9805);
xnor U10163 (N_10163,N_9797,N_9689);
or U10164 (N_10164,N_9886,N_9633);
or U10165 (N_10165,N_9632,N_9691);
xor U10166 (N_10166,N_9813,N_9886);
nand U10167 (N_10167,N_9714,N_9830);
nor U10168 (N_10168,N_9835,N_9717);
nor U10169 (N_10169,N_9803,N_9706);
nor U10170 (N_10170,N_9772,N_9685);
nand U10171 (N_10171,N_9875,N_9863);
nor U10172 (N_10172,N_9891,N_9870);
nand U10173 (N_10173,N_9684,N_9773);
and U10174 (N_10174,N_9764,N_9709);
or U10175 (N_10175,N_9890,N_9737);
and U10176 (N_10176,N_9703,N_9722);
and U10177 (N_10177,N_9899,N_9722);
or U10178 (N_10178,N_9750,N_9705);
nor U10179 (N_10179,N_9680,N_9895);
nor U10180 (N_10180,N_9685,N_9728);
nor U10181 (N_10181,N_9761,N_9744);
and U10182 (N_10182,N_9627,N_9819);
xnor U10183 (N_10183,N_9816,N_9650);
or U10184 (N_10184,N_9780,N_9896);
or U10185 (N_10185,N_9819,N_9786);
nor U10186 (N_10186,N_9612,N_9708);
or U10187 (N_10187,N_9869,N_9691);
and U10188 (N_10188,N_9678,N_9818);
nor U10189 (N_10189,N_9887,N_9759);
nor U10190 (N_10190,N_9684,N_9721);
nand U10191 (N_10191,N_9749,N_9882);
nand U10192 (N_10192,N_9802,N_9648);
xnor U10193 (N_10193,N_9738,N_9862);
and U10194 (N_10194,N_9757,N_9618);
nor U10195 (N_10195,N_9884,N_9834);
or U10196 (N_10196,N_9666,N_9735);
and U10197 (N_10197,N_9871,N_9601);
and U10198 (N_10198,N_9613,N_9635);
nand U10199 (N_10199,N_9728,N_9721);
or U10200 (N_10200,N_10153,N_10111);
and U10201 (N_10201,N_10138,N_10022);
nand U10202 (N_10202,N_10118,N_10099);
nand U10203 (N_10203,N_9997,N_10177);
xor U10204 (N_10204,N_10016,N_10082);
nand U10205 (N_10205,N_9932,N_9915);
and U10206 (N_10206,N_9914,N_10131);
nor U10207 (N_10207,N_10133,N_10078);
and U10208 (N_10208,N_9952,N_10002);
and U10209 (N_10209,N_10066,N_10000);
or U10210 (N_10210,N_9937,N_10041);
or U10211 (N_10211,N_10097,N_10019);
nor U10212 (N_10212,N_10156,N_10144);
xnor U10213 (N_10213,N_10071,N_9964);
xnor U10214 (N_10214,N_10180,N_9949);
or U10215 (N_10215,N_10028,N_10146);
or U10216 (N_10216,N_10084,N_9998);
and U10217 (N_10217,N_10158,N_10155);
or U10218 (N_10218,N_10054,N_10074);
or U10219 (N_10219,N_10092,N_10150);
and U10220 (N_10220,N_9991,N_10086);
or U10221 (N_10221,N_10089,N_9917);
nor U10222 (N_10222,N_9906,N_9986);
nand U10223 (N_10223,N_10115,N_10185);
nand U10224 (N_10224,N_9943,N_9990);
and U10225 (N_10225,N_10110,N_10112);
and U10226 (N_10226,N_10073,N_10070);
or U10227 (N_10227,N_10045,N_10102);
or U10228 (N_10228,N_10021,N_10091);
xnor U10229 (N_10229,N_9959,N_10007);
nor U10230 (N_10230,N_9987,N_10108);
nand U10231 (N_10231,N_10173,N_9908);
and U10232 (N_10232,N_10151,N_10004);
xor U10233 (N_10233,N_10159,N_10191);
nor U10234 (N_10234,N_10085,N_9930);
xnor U10235 (N_10235,N_10093,N_9909);
or U10236 (N_10236,N_9948,N_10130);
nor U10237 (N_10237,N_9981,N_9905);
nor U10238 (N_10238,N_9940,N_10032);
and U10239 (N_10239,N_10184,N_10119);
nor U10240 (N_10240,N_10077,N_10051);
and U10241 (N_10241,N_10142,N_9988);
and U10242 (N_10242,N_10178,N_10129);
nand U10243 (N_10243,N_10125,N_10167);
and U10244 (N_10244,N_10080,N_9935);
xor U10245 (N_10245,N_10145,N_9912);
and U10246 (N_10246,N_9926,N_9901);
xnor U10247 (N_10247,N_10047,N_10075);
nand U10248 (N_10248,N_9983,N_10175);
xnor U10249 (N_10249,N_10174,N_9922);
or U10250 (N_10250,N_10043,N_10050);
nor U10251 (N_10251,N_10165,N_10056);
and U10252 (N_10252,N_10098,N_10199);
or U10253 (N_10253,N_10198,N_10096);
or U10254 (N_10254,N_10020,N_10104);
and U10255 (N_10255,N_9907,N_10005);
nor U10256 (N_10256,N_10193,N_10106);
nand U10257 (N_10257,N_10181,N_9962);
or U10258 (N_10258,N_10067,N_10038);
nand U10259 (N_10259,N_10152,N_10029);
nor U10260 (N_10260,N_10189,N_10011);
xor U10261 (N_10261,N_9970,N_10134);
nor U10262 (N_10262,N_9972,N_9984);
and U10263 (N_10263,N_10126,N_9956);
xor U10264 (N_10264,N_9946,N_10079);
nor U10265 (N_10265,N_10109,N_10052);
nand U10266 (N_10266,N_9958,N_10026);
nor U10267 (N_10267,N_9941,N_10059);
and U10268 (N_10268,N_9989,N_10182);
nor U10269 (N_10269,N_10187,N_9978);
and U10270 (N_10270,N_10010,N_10058);
or U10271 (N_10271,N_10140,N_10132);
xnor U10272 (N_10272,N_9900,N_9971);
xor U10273 (N_10273,N_10120,N_10083);
nor U10274 (N_10274,N_10055,N_10117);
xor U10275 (N_10275,N_10035,N_10039);
nor U10276 (N_10276,N_10046,N_9916);
and U10277 (N_10277,N_9961,N_10049);
and U10278 (N_10278,N_9950,N_9927);
or U10279 (N_10279,N_10033,N_10057);
nand U10280 (N_10280,N_9993,N_10061);
nor U10281 (N_10281,N_10122,N_9913);
nand U10282 (N_10282,N_10162,N_9982);
nand U10283 (N_10283,N_10161,N_9976);
or U10284 (N_10284,N_10123,N_10023);
xor U10285 (N_10285,N_9918,N_10068);
xnor U10286 (N_10286,N_10088,N_9992);
xnor U10287 (N_10287,N_10105,N_10176);
nor U10288 (N_10288,N_10149,N_9968);
or U10289 (N_10289,N_10171,N_10069);
and U10290 (N_10290,N_10148,N_10087);
xnor U10291 (N_10291,N_9980,N_9999);
nor U10292 (N_10292,N_10103,N_9920);
nor U10293 (N_10293,N_10034,N_10024);
nor U10294 (N_10294,N_10037,N_9966);
nor U10295 (N_10295,N_10013,N_9934);
and U10296 (N_10296,N_9995,N_10168);
or U10297 (N_10297,N_10114,N_10101);
xnor U10298 (N_10298,N_10141,N_10160);
nor U10299 (N_10299,N_10001,N_10018);
nor U10300 (N_10300,N_9921,N_10014);
nand U10301 (N_10301,N_10192,N_10006);
and U10302 (N_10302,N_9944,N_9969);
nor U10303 (N_10303,N_10015,N_9960);
nor U10304 (N_10304,N_10042,N_10031);
nand U10305 (N_10305,N_9957,N_10128);
and U10306 (N_10306,N_10053,N_10166);
or U10307 (N_10307,N_9951,N_9902);
xor U10308 (N_10308,N_9973,N_9931);
nand U10309 (N_10309,N_10194,N_9911);
nand U10310 (N_10310,N_9923,N_9965);
nand U10311 (N_10311,N_10027,N_10030);
nor U10312 (N_10312,N_9910,N_10044);
nor U10313 (N_10313,N_10137,N_10196);
or U10314 (N_10314,N_9994,N_9977);
and U10315 (N_10315,N_9925,N_10154);
xnor U10316 (N_10316,N_9947,N_9938);
nor U10317 (N_10317,N_10081,N_10025);
or U10318 (N_10318,N_10116,N_10017);
or U10319 (N_10319,N_9928,N_9963);
nor U10320 (N_10320,N_10063,N_10048);
nand U10321 (N_10321,N_10164,N_9953);
xnor U10322 (N_10322,N_9929,N_10107);
nor U10323 (N_10323,N_10195,N_10008);
xnor U10324 (N_10324,N_10147,N_10121);
or U10325 (N_10325,N_10036,N_10183);
nor U10326 (N_10326,N_10064,N_9979);
or U10327 (N_10327,N_10163,N_10060);
nand U10328 (N_10328,N_9919,N_10135);
or U10329 (N_10329,N_10095,N_9942);
xnor U10330 (N_10330,N_10172,N_10124);
nor U10331 (N_10331,N_10186,N_10139);
or U10332 (N_10332,N_9903,N_9945);
or U10333 (N_10333,N_10094,N_10062);
nor U10334 (N_10334,N_10143,N_10179);
or U10335 (N_10335,N_10072,N_10113);
nand U10336 (N_10336,N_10012,N_9939);
nand U10337 (N_10337,N_9996,N_10127);
nor U10338 (N_10338,N_10170,N_10169);
xnor U10339 (N_10339,N_9975,N_10090);
or U10340 (N_10340,N_10100,N_10065);
nor U10341 (N_10341,N_10197,N_9967);
nand U10342 (N_10342,N_10009,N_10076);
and U10343 (N_10343,N_9933,N_9974);
xnor U10344 (N_10344,N_10040,N_10136);
nand U10345 (N_10345,N_10190,N_10188);
nor U10346 (N_10346,N_9954,N_10157);
nand U10347 (N_10347,N_9904,N_9985);
or U10348 (N_10348,N_9936,N_9924);
and U10349 (N_10349,N_10003,N_9955);
xnor U10350 (N_10350,N_9971,N_9915);
or U10351 (N_10351,N_10012,N_10062);
or U10352 (N_10352,N_9902,N_10070);
nand U10353 (N_10353,N_9986,N_10123);
xor U10354 (N_10354,N_10182,N_9963);
nand U10355 (N_10355,N_10113,N_10176);
nand U10356 (N_10356,N_10139,N_9948);
and U10357 (N_10357,N_9941,N_9909);
or U10358 (N_10358,N_10077,N_10068);
nor U10359 (N_10359,N_9914,N_9920);
nor U10360 (N_10360,N_10084,N_10153);
nand U10361 (N_10361,N_9913,N_10065);
xnor U10362 (N_10362,N_10186,N_9931);
nand U10363 (N_10363,N_10185,N_9997);
nand U10364 (N_10364,N_9924,N_9983);
and U10365 (N_10365,N_10154,N_10170);
xor U10366 (N_10366,N_10106,N_10002);
or U10367 (N_10367,N_10169,N_10167);
and U10368 (N_10368,N_10054,N_9996);
xnor U10369 (N_10369,N_10179,N_10055);
and U10370 (N_10370,N_10151,N_9932);
nor U10371 (N_10371,N_10172,N_10022);
nand U10372 (N_10372,N_9914,N_10103);
and U10373 (N_10373,N_10152,N_9985);
and U10374 (N_10374,N_9902,N_10166);
nor U10375 (N_10375,N_10086,N_10041);
or U10376 (N_10376,N_10196,N_10151);
nor U10377 (N_10377,N_10038,N_10104);
or U10378 (N_10378,N_10070,N_9988);
and U10379 (N_10379,N_10173,N_10130);
nand U10380 (N_10380,N_10062,N_9941);
xor U10381 (N_10381,N_9922,N_10003);
xor U10382 (N_10382,N_10049,N_9921);
and U10383 (N_10383,N_10063,N_9959);
nand U10384 (N_10384,N_10092,N_10119);
nor U10385 (N_10385,N_10037,N_10100);
or U10386 (N_10386,N_10089,N_10040);
xor U10387 (N_10387,N_9911,N_10084);
or U10388 (N_10388,N_10184,N_10026);
and U10389 (N_10389,N_10126,N_9940);
or U10390 (N_10390,N_10045,N_10104);
nor U10391 (N_10391,N_10068,N_10106);
nor U10392 (N_10392,N_10085,N_10095);
nor U10393 (N_10393,N_10007,N_9936);
and U10394 (N_10394,N_10067,N_10104);
and U10395 (N_10395,N_10002,N_10136);
and U10396 (N_10396,N_10118,N_10175);
and U10397 (N_10397,N_10071,N_9912);
nand U10398 (N_10398,N_10143,N_10004);
and U10399 (N_10399,N_10019,N_9920);
or U10400 (N_10400,N_10146,N_10069);
nand U10401 (N_10401,N_9917,N_10122);
and U10402 (N_10402,N_10018,N_9906);
nand U10403 (N_10403,N_10166,N_10060);
nand U10404 (N_10404,N_10155,N_10157);
xnor U10405 (N_10405,N_10167,N_9939);
xnor U10406 (N_10406,N_9980,N_9919);
xor U10407 (N_10407,N_10096,N_10116);
nor U10408 (N_10408,N_10153,N_9938);
xor U10409 (N_10409,N_10099,N_10043);
xor U10410 (N_10410,N_10024,N_10131);
nand U10411 (N_10411,N_10027,N_10058);
or U10412 (N_10412,N_10116,N_10005);
nand U10413 (N_10413,N_9958,N_9964);
and U10414 (N_10414,N_10044,N_10183);
nor U10415 (N_10415,N_10157,N_10006);
nor U10416 (N_10416,N_10050,N_10102);
nor U10417 (N_10417,N_10175,N_10191);
nand U10418 (N_10418,N_10053,N_10038);
nand U10419 (N_10419,N_10180,N_9952);
nor U10420 (N_10420,N_10061,N_10047);
and U10421 (N_10421,N_9938,N_10172);
nand U10422 (N_10422,N_9948,N_9955);
and U10423 (N_10423,N_9965,N_10110);
nand U10424 (N_10424,N_10097,N_10060);
or U10425 (N_10425,N_10165,N_10083);
nand U10426 (N_10426,N_10114,N_10094);
xnor U10427 (N_10427,N_10132,N_10155);
nor U10428 (N_10428,N_10193,N_9936);
nand U10429 (N_10429,N_10175,N_10192);
nor U10430 (N_10430,N_9929,N_10081);
xnor U10431 (N_10431,N_9952,N_9911);
xor U10432 (N_10432,N_10089,N_10073);
and U10433 (N_10433,N_10091,N_10167);
nor U10434 (N_10434,N_9933,N_9900);
or U10435 (N_10435,N_10116,N_9967);
and U10436 (N_10436,N_9989,N_10080);
xnor U10437 (N_10437,N_10085,N_9933);
nand U10438 (N_10438,N_10129,N_10056);
xnor U10439 (N_10439,N_10088,N_10067);
xor U10440 (N_10440,N_10159,N_10002);
or U10441 (N_10441,N_10199,N_10071);
xor U10442 (N_10442,N_10000,N_10049);
or U10443 (N_10443,N_10139,N_9954);
xnor U10444 (N_10444,N_10197,N_10053);
nand U10445 (N_10445,N_10192,N_9997);
nor U10446 (N_10446,N_10020,N_10147);
and U10447 (N_10447,N_10079,N_9905);
and U10448 (N_10448,N_10198,N_10103);
xnor U10449 (N_10449,N_10025,N_10023);
or U10450 (N_10450,N_10030,N_9993);
xnor U10451 (N_10451,N_10137,N_10086);
nor U10452 (N_10452,N_10177,N_9952);
or U10453 (N_10453,N_9903,N_10160);
nor U10454 (N_10454,N_10174,N_9945);
nor U10455 (N_10455,N_10022,N_10146);
nand U10456 (N_10456,N_9967,N_9910);
or U10457 (N_10457,N_10155,N_9968);
xnor U10458 (N_10458,N_9982,N_10127);
nor U10459 (N_10459,N_10181,N_10088);
and U10460 (N_10460,N_10002,N_9932);
xor U10461 (N_10461,N_10154,N_9936);
or U10462 (N_10462,N_10017,N_10144);
nor U10463 (N_10463,N_9979,N_10101);
and U10464 (N_10464,N_10000,N_10019);
nand U10465 (N_10465,N_10076,N_10197);
xnor U10466 (N_10466,N_10091,N_9984);
nor U10467 (N_10467,N_10102,N_10017);
xor U10468 (N_10468,N_10137,N_10120);
nor U10469 (N_10469,N_9912,N_10058);
and U10470 (N_10470,N_10046,N_10157);
nor U10471 (N_10471,N_9930,N_10197);
or U10472 (N_10472,N_9923,N_10050);
nor U10473 (N_10473,N_10053,N_10177);
or U10474 (N_10474,N_9946,N_10016);
nand U10475 (N_10475,N_10017,N_9934);
or U10476 (N_10476,N_10057,N_9947);
and U10477 (N_10477,N_10134,N_10004);
nand U10478 (N_10478,N_10135,N_10065);
xnor U10479 (N_10479,N_9960,N_10073);
or U10480 (N_10480,N_10083,N_10098);
nor U10481 (N_10481,N_10136,N_9979);
nor U10482 (N_10482,N_10137,N_10004);
nor U10483 (N_10483,N_10032,N_10104);
nor U10484 (N_10484,N_9907,N_10028);
xnor U10485 (N_10485,N_9944,N_9945);
xnor U10486 (N_10486,N_9950,N_10065);
xnor U10487 (N_10487,N_9933,N_9968);
nand U10488 (N_10488,N_9930,N_10108);
nor U10489 (N_10489,N_9934,N_10151);
nand U10490 (N_10490,N_10178,N_10098);
or U10491 (N_10491,N_9990,N_10179);
or U10492 (N_10492,N_9975,N_10033);
and U10493 (N_10493,N_10047,N_9991);
nor U10494 (N_10494,N_10145,N_10103);
nor U10495 (N_10495,N_10174,N_10117);
and U10496 (N_10496,N_9934,N_9901);
nor U10497 (N_10497,N_10062,N_9911);
xor U10498 (N_10498,N_9908,N_9970);
nand U10499 (N_10499,N_9963,N_10173);
nand U10500 (N_10500,N_10374,N_10324);
or U10501 (N_10501,N_10327,N_10266);
xor U10502 (N_10502,N_10449,N_10293);
nor U10503 (N_10503,N_10397,N_10265);
nand U10504 (N_10504,N_10447,N_10490);
or U10505 (N_10505,N_10310,N_10296);
xor U10506 (N_10506,N_10337,N_10303);
xnor U10507 (N_10507,N_10235,N_10416);
nand U10508 (N_10508,N_10281,N_10285);
and U10509 (N_10509,N_10469,N_10319);
and U10510 (N_10510,N_10220,N_10209);
xnor U10511 (N_10511,N_10345,N_10444);
xor U10512 (N_10512,N_10340,N_10218);
xnor U10513 (N_10513,N_10239,N_10452);
or U10514 (N_10514,N_10255,N_10393);
xnor U10515 (N_10515,N_10390,N_10480);
nor U10516 (N_10516,N_10385,N_10458);
nor U10517 (N_10517,N_10460,N_10495);
nand U10518 (N_10518,N_10422,N_10216);
and U10519 (N_10519,N_10295,N_10233);
nor U10520 (N_10520,N_10427,N_10481);
nor U10521 (N_10521,N_10342,N_10386);
nand U10522 (N_10522,N_10333,N_10367);
nor U10523 (N_10523,N_10377,N_10360);
and U10524 (N_10524,N_10356,N_10232);
xnor U10525 (N_10525,N_10329,N_10365);
or U10526 (N_10526,N_10364,N_10243);
or U10527 (N_10527,N_10446,N_10245);
xor U10528 (N_10528,N_10361,N_10226);
or U10529 (N_10529,N_10299,N_10322);
nand U10530 (N_10530,N_10249,N_10334);
and U10531 (N_10531,N_10475,N_10308);
or U10532 (N_10532,N_10461,N_10463);
or U10533 (N_10533,N_10201,N_10257);
nor U10534 (N_10534,N_10211,N_10395);
nand U10535 (N_10535,N_10371,N_10277);
nand U10536 (N_10536,N_10309,N_10399);
xor U10537 (N_10537,N_10489,N_10445);
or U10538 (N_10538,N_10437,N_10259);
and U10539 (N_10539,N_10407,N_10208);
and U10540 (N_10540,N_10478,N_10331);
xnor U10541 (N_10541,N_10482,N_10264);
nand U10542 (N_10542,N_10392,N_10434);
or U10543 (N_10543,N_10472,N_10251);
xnor U10544 (N_10544,N_10234,N_10230);
or U10545 (N_10545,N_10493,N_10419);
nand U10546 (N_10546,N_10272,N_10453);
and U10547 (N_10547,N_10315,N_10261);
xor U10548 (N_10548,N_10421,N_10219);
and U10549 (N_10549,N_10352,N_10213);
and U10550 (N_10550,N_10273,N_10202);
or U10551 (N_10551,N_10372,N_10498);
nor U10552 (N_10552,N_10236,N_10290);
and U10553 (N_10553,N_10271,N_10450);
nand U10554 (N_10554,N_10237,N_10267);
nor U10555 (N_10555,N_10430,N_10441);
or U10556 (N_10556,N_10387,N_10240);
xnor U10557 (N_10557,N_10438,N_10442);
xor U10558 (N_10558,N_10306,N_10341);
or U10559 (N_10559,N_10274,N_10224);
and U10560 (N_10560,N_10215,N_10379);
or U10561 (N_10561,N_10326,N_10487);
and U10562 (N_10562,N_10276,N_10375);
and U10563 (N_10563,N_10280,N_10436);
nor U10564 (N_10564,N_10486,N_10488);
nor U10565 (N_10565,N_10238,N_10204);
or U10566 (N_10566,N_10250,N_10207);
nor U10567 (N_10567,N_10380,N_10378);
or U10568 (N_10568,N_10203,N_10406);
nand U10569 (N_10569,N_10459,N_10253);
xnor U10570 (N_10570,N_10466,N_10328);
xor U10571 (N_10571,N_10431,N_10321);
or U10572 (N_10572,N_10212,N_10351);
nor U10573 (N_10573,N_10363,N_10394);
xnor U10574 (N_10574,N_10314,N_10343);
nor U10575 (N_10575,N_10214,N_10464);
nand U10576 (N_10576,N_10411,N_10292);
or U10577 (N_10577,N_10366,N_10389);
nand U10578 (N_10578,N_10223,N_10408);
nand U10579 (N_10579,N_10228,N_10476);
and U10580 (N_10580,N_10435,N_10443);
nand U10581 (N_10581,N_10317,N_10382);
or U10582 (N_10582,N_10301,N_10256);
xor U10583 (N_10583,N_10483,N_10418);
xor U10584 (N_10584,N_10451,N_10433);
and U10585 (N_10585,N_10425,N_10404);
nand U10586 (N_10586,N_10325,N_10470);
or U10587 (N_10587,N_10298,N_10323);
xor U10588 (N_10588,N_10396,N_10335);
or U10589 (N_10589,N_10428,N_10294);
xnor U10590 (N_10590,N_10288,N_10354);
and U10591 (N_10591,N_10330,N_10426);
nor U10592 (N_10592,N_10359,N_10350);
nor U10593 (N_10593,N_10391,N_10297);
nor U10594 (N_10594,N_10225,N_10413);
nand U10595 (N_10595,N_10388,N_10227);
xor U10596 (N_10596,N_10222,N_10205);
nand U10597 (N_10597,N_10244,N_10381);
or U10598 (N_10598,N_10468,N_10311);
or U10599 (N_10599,N_10403,N_10275);
nor U10600 (N_10600,N_10362,N_10231);
xor U10601 (N_10601,N_10473,N_10499);
nand U10602 (N_10602,N_10383,N_10344);
and U10603 (N_10603,N_10284,N_10286);
nor U10604 (N_10604,N_10258,N_10304);
nand U10605 (N_10605,N_10440,N_10420);
xor U10606 (N_10606,N_10355,N_10467);
and U10607 (N_10607,N_10313,N_10398);
or U10608 (N_10608,N_10347,N_10348);
nand U10609 (N_10609,N_10217,N_10318);
or U10610 (N_10610,N_10402,N_10312);
nand U10611 (N_10611,N_10405,N_10283);
or U10612 (N_10612,N_10477,N_10263);
nand U10613 (N_10613,N_10279,N_10415);
and U10614 (N_10614,N_10457,N_10494);
nor U10615 (N_10615,N_10492,N_10455);
xnor U10616 (N_10616,N_10496,N_10242);
nor U10617 (N_10617,N_10429,N_10485);
or U10618 (N_10618,N_10357,N_10241);
nor U10619 (N_10619,N_10432,N_10302);
xnor U10620 (N_10620,N_10247,N_10307);
xor U10621 (N_10621,N_10270,N_10474);
or U10622 (N_10622,N_10369,N_10260);
xor U10623 (N_10623,N_10439,N_10454);
and U10624 (N_10624,N_10278,N_10484);
nor U10625 (N_10625,N_10254,N_10368);
or U10626 (N_10626,N_10370,N_10349);
nand U10627 (N_10627,N_10346,N_10262);
or U10628 (N_10628,N_10353,N_10248);
nor U10629 (N_10629,N_10206,N_10462);
or U10630 (N_10630,N_10291,N_10289);
nand U10631 (N_10631,N_10479,N_10423);
nor U10632 (N_10632,N_10497,N_10332);
nand U10633 (N_10633,N_10287,N_10300);
nor U10634 (N_10634,N_10252,N_10376);
nor U10635 (N_10635,N_10338,N_10246);
nor U10636 (N_10636,N_10448,N_10384);
and U10637 (N_10637,N_10414,N_10409);
and U10638 (N_10638,N_10358,N_10401);
and U10639 (N_10639,N_10336,N_10410);
xor U10640 (N_10640,N_10491,N_10339);
xnor U10641 (N_10641,N_10456,N_10373);
nand U10642 (N_10642,N_10320,N_10400);
and U10643 (N_10643,N_10471,N_10229);
nor U10644 (N_10644,N_10305,N_10424);
or U10645 (N_10645,N_10221,N_10268);
or U10646 (N_10646,N_10210,N_10412);
nand U10647 (N_10647,N_10282,N_10200);
xor U10648 (N_10648,N_10417,N_10316);
nor U10649 (N_10649,N_10465,N_10269);
and U10650 (N_10650,N_10208,N_10299);
or U10651 (N_10651,N_10253,N_10328);
or U10652 (N_10652,N_10397,N_10262);
or U10653 (N_10653,N_10358,N_10235);
nor U10654 (N_10654,N_10363,N_10395);
and U10655 (N_10655,N_10388,N_10428);
or U10656 (N_10656,N_10301,N_10494);
nand U10657 (N_10657,N_10499,N_10268);
or U10658 (N_10658,N_10474,N_10393);
or U10659 (N_10659,N_10233,N_10205);
xor U10660 (N_10660,N_10266,N_10255);
or U10661 (N_10661,N_10323,N_10464);
nor U10662 (N_10662,N_10221,N_10315);
and U10663 (N_10663,N_10269,N_10389);
and U10664 (N_10664,N_10214,N_10465);
nor U10665 (N_10665,N_10332,N_10244);
xnor U10666 (N_10666,N_10219,N_10261);
nor U10667 (N_10667,N_10414,N_10280);
and U10668 (N_10668,N_10309,N_10371);
nor U10669 (N_10669,N_10406,N_10261);
nor U10670 (N_10670,N_10459,N_10260);
and U10671 (N_10671,N_10245,N_10479);
and U10672 (N_10672,N_10283,N_10346);
nand U10673 (N_10673,N_10279,N_10338);
nor U10674 (N_10674,N_10204,N_10464);
nor U10675 (N_10675,N_10293,N_10303);
xnor U10676 (N_10676,N_10271,N_10284);
nand U10677 (N_10677,N_10407,N_10316);
xnor U10678 (N_10678,N_10227,N_10431);
nor U10679 (N_10679,N_10263,N_10431);
nor U10680 (N_10680,N_10408,N_10336);
xor U10681 (N_10681,N_10394,N_10494);
xnor U10682 (N_10682,N_10405,N_10359);
or U10683 (N_10683,N_10342,N_10231);
and U10684 (N_10684,N_10437,N_10422);
and U10685 (N_10685,N_10416,N_10413);
or U10686 (N_10686,N_10216,N_10441);
nand U10687 (N_10687,N_10481,N_10229);
xnor U10688 (N_10688,N_10422,N_10203);
nor U10689 (N_10689,N_10332,N_10268);
and U10690 (N_10690,N_10267,N_10222);
xnor U10691 (N_10691,N_10429,N_10487);
or U10692 (N_10692,N_10453,N_10382);
and U10693 (N_10693,N_10459,N_10281);
or U10694 (N_10694,N_10442,N_10278);
or U10695 (N_10695,N_10345,N_10241);
nand U10696 (N_10696,N_10237,N_10259);
nor U10697 (N_10697,N_10348,N_10455);
xnor U10698 (N_10698,N_10416,N_10475);
nand U10699 (N_10699,N_10476,N_10200);
nor U10700 (N_10700,N_10208,N_10373);
or U10701 (N_10701,N_10225,N_10476);
nor U10702 (N_10702,N_10222,N_10410);
nor U10703 (N_10703,N_10354,N_10448);
xnor U10704 (N_10704,N_10212,N_10454);
or U10705 (N_10705,N_10331,N_10217);
nor U10706 (N_10706,N_10293,N_10327);
or U10707 (N_10707,N_10332,N_10407);
and U10708 (N_10708,N_10438,N_10221);
and U10709 (N_10709,N_10228,N_10302);
nor U10710 (N_10710,N_10223,N_10459);
or U10711 (N_10711,N_10492,N_10304);
and U10712 (N_10712,N_10386,N_10364);
and U10713 (N_10713,N_10392,N_10315);
and U10714 (N_10714,N_10261,N_10442);
or U10715 (N_10715,N_10399,N_10236);
or U10716 (N_10716,N_10369,N_10363);
nor U10717 (N_10717,N_10397,N_10437);
nor U10718 (N_10718,N_10421,N_10358);
and U10719 (N_10719,N_10436,N_10324);
or U10720 (N_10720,N_10349,N_10228);
xnor U10721 (N_10721,N_10495,N_10282);
nand U10722 (N_10722,N_10412,N_10349);
or U10723 (N_10723,N_10267,N_10325);
nor U10724 (N_10724,N_10275,N_10393);
nor U10725 (N_10725,N_10251,N_10278);
and U10726 (N_10726,N_10279,N_10305);
or U10727 (N_10727,N_10362,N_10211);
nand U10728 (N_10728,N_10337,N_10497);
and U10729 (N_10729,N_10275,N_10448);
or U10730 (N_10730,N_10384,N_10464);
or U10731 (N_10731,N_10420,N_10480);
or U10732 (N_10732,N_10499,N_10460);
and U10733 (N_10733,N_10258,N_10221);
nor U10734 (N_10734,N_10357,N_10418);
and U10735 (N_10735,N_10453,N_10214);
or U10736 (N_10736,N_10351,N_10302);
nor U10737 (N_10737,N_10248,N_10322);
nand U10738 (N_10738,N_10461,N_10342);
or U10739 (N_10739,N_10425,N_10341);
or U10740 (N_10740,N_10406,N_10264);
nor U10741 (N_10741,N_10376,N_10303);
nor U10742 (N_10742,N_10374,N_10313);
nand U10743 (N_10743,N_10453,N_10266);
nor U10744 (N_10744,N_10400,N_10410);
nor U10745 (N_10745,N_10396,N_10379);
or U10746 (N_10746,N_10486,N_10304);
and U10747 (N_10747,N_10344,N_10245);
xnor U10748 (N_10748,N_10209,N_10280);
nand U10749 (N_10749,N_10274,N_10439);
or U10750 (N_10750,N_10218,N_10361);
xor U10751 (N_10751,N_10299,N_10371);
xor U10752 (N_10752,N_10259,N_10467);
xnor U10753 (N_10753,N_10202,N_10420);
xor U10754 (N_10754,N_10266,N_10416);
nor U10755 (N_10755,N_10476,N_10326);
and U10756 (N_10756,N_10313,N_10252);
nor U10757 (N_10757,N_10493,N_10207);
or U10758 (N_10758,N_10495,N_10479);
nor U10759 (N_10759,N_10386,N_10423);
nor U10760 (N_10760,N_10270,N_10436);
xnor U10761 (N_10761,N_10266,N_10341);
and U10762 (N_10762,N_10253,N_10438);
nand U10763 (N_10763,N_10241,N_10344);
xor U10764 (N_10764,N_10201,N_10273);
nand U10765 (N_10765,N_10371,N_10345);
or U10766 (N_10766,N_10409,N_10424);
xnor U10767 (N_10767,N_10424,N_10383);
and U10768 (N_10768,N_10485,N_10409);
nor U10769 (N_10769,N_10495,N_10231);
nand U10770 (N_10770,N_10298,N_10383);
nand U10771 (N_10771,N_10427,N_10372);
nor U10772 (N_10772,N_10443,N_10250);
nand U10773 (N_10773,N_10296,N_10263);
nand U10774 (N_10774,N_10230,N_10286);
or U10775 (N_10775,N_10297,N_10347);
xnor U10776 (N_10776,N_10489,N_10317);
or U10777 (N_10777,N_10457,N_10404);
nand U10778 (N_10778,N_10330,N_10283);
nand U10779 (N_10779,N_10292,N_10349);
xor U10780 (N_10780,N_10237,N_10305);
nor U10781 (N_10781,N_10226,N_10337);
xor U10782 (N_10782,N_10358,N_10216);
nand U10783 (N_10783,N_10429,N_10415);
xnor U10784 (N_10784,N_10385,N_10434);
or U10785 (N_10785,N_10427,N_10367);
or U10786 (N_10786,N_10436,N_10409);
nor U10787 (N_10787,N_10485,N_10475);
xnor U10788 (N_10788,N_10419,N_10480);
nor U10789 (N_10789,N_10300,N_10321);
xor U10790 (N_10790,N_10472,N_10390);
nor U10791 (N_10791,N_10389,N_10201);
nor U10792 (N_10792,N_10366,N_10307);
nor U10793 (N_10793,N_10447,N_10383);
nor U10794 (N_10794,N_10369,N_10298);
nand U10795 (N_10795,N_10269,N_10296);
nor U10796 (N_10796,N_10386,N_10358);
nor U10797 (N_10797,N_10320,N_10385);
or U10798 (N_10798,N_10375,N_10220);
nand U10799 (N_10799,N_10349,N_10313);
nor U10800 (N_10800,N_10595,N_10646);
nor U10801 (N_10801,N_10681,N_10582);
nand U10802 (N_10802,N_10612,N_10679);
or U10803 (N_10803,N_10773,N_10790);
xnor U10804 (N_10804,N_10641,N_10711);
xnor U10805 (N_10805,N_10705,N_10785);
nand U10806 (N_10806,N_10631,N_10789);
xor U10807 (N_10807,N_10793,N_10558);
or U10808 (N_10808,N_10666,N_10639);
or U10809 (N_10809,N_10556,N_10704);
nand U10810 (N_10810,N_10756,N_10664);
xnor U10811 (N_10811,N_10742,N_10621);
nand U10812 (N_10812,N_10607,N_10682);
nand U10813 (N_10813,N_10555,N_10763);
xor U10814 (N_10814,N_10562,N_10581);
and U10815 (N_10815,N_10799,N_10531);
and U10816 (N_10816,N_10642,N_10616);
and U10817 (N_10817,N_10587,N_10638);
nand U10818 (N_10818,N_10518,N_10514);
and U10819 (N_10819,N_10502,N_10598);
or U10820 (N_10820,N_10659,N_10762);
and U10821 (N_10821,N_10637,N_10569);
and U10822 (N_10822,N_10758,N_10528);
xor U10823 (N_10823,N_10594,N_10606);
and U10824 (N_10824,N_10623,N_10533);
nand U10825 (N_10825,N_10510,N_10584);
nand U10826 (N_10826,N_10733,N_10749);
nand U10827 (N_10827,N_10507,N_10716);
or U10828 (N_10828,N_10599,N_10523);
and U10829 (N_10829,N_10661,N_10532);
or U10830 (N_10830,N_10668,N_10740);
nor U10831 (N_10831,N_10683,N_10747);
nand U10832 (N_10832,N_10709,N_10585);
xor U10833 (N_10833,N_10706,N_10689);
and U10834 (N_10834,N_10560,N_10543);
xor U10835 (N_10835,N_10680,N_10651);
nand U10836 (N_10836,N_10529,N_10794);
nand U10837 (N_10837,N_10624,N_10792);
xor U10838 (N_10838,N_10512,N_10547);
xnor U10839 (N_10839,N_10734,N_10537);
nor U10840 (N_10840,N_10636,N_10563);
or U10841 (N_10841,N_10746,N_10658);
nor U10842 (N_10842,N_10564,N_10571);
and U10843 (N_10843,N_10613,N_10736);
and U10844 (N_10844,N_10630,N_10629);
xnor U10845 (N_10845,N_10513,N_10797);
xor U10846 (N_10846,N_10784,N_10656);
xor U10847 (N_10847,N_10710,N_10534);
and U10848 (N_10848,N_10504,N_10778);
or U10849 (N_10849,N_10772,N_10684);
or U10850 (N_10850,N_10782,N_10687);
or U10851 (N_10851,N_10781,N_10720);
and U10852 (N_10852,N_10753,N_10591);
and U10853 (N_10853,N_10695,N_10660);
or U10854 (N_10854,N_10643,N_10748);
nand U10855 (N_10855,N_10712,N_10501);
xnor U10856 (N_10856,N_10743,N_10718);
or U10857 (N_10857,N_10551,N_10647);
or U10858 (N_10858,N_10751,N_10698);
nor U10859 (N_10859,N_10542,N_10725);
xor U10860 (N_10860,N_10615,N_10634);
nand U10861 (N_10861,N_10674,N_10670);
xnor U10862 (N_10862,N_10541,N_10786);
xor U10863 (N_10863,N_10791,N_10663);
and U10864 (N_10864,N_10685,N_10576);
nand U10865 (N_10865,N_10795,N_10618);
xnor U10866 (N_10866,N_10766,N_10644);
and U10867 (N_10867,N_10506,N_10653);
nand U10868 (N_10868,N_10574,N_10548);
xnor U10869 (N_10869,N_10731,N_10759);
xor U10870 (N_10870,N_10610,N_10538);
and U10871 (N_10871,N_10719,N_10707);
or U10872 (N_10872,N_10774,N_10578);
xor U10873 (N_10873,N_10770,N_10566);
xnor U10874 (N_10874,N_10568,N_10761);
nor U10875 (N_10875,N_10741,N_10667);
nand U10876 (N_10876,N_10527,N_10633);
or U10877 (N_10877,N_10776,N_10605);
and U10878 (N_10878,N_10655,N_10662);
nand U10879 (N_10879,N_10750,N_10767);
nand U10880 (N_10880,N_10696,N_10597);
xor U10881 (N_10881,N_10545,N_10721);
xnor U10882 (N_10882,N_10693,N_10671);
nor U10883 (N_10883,N_10549,N_10602);
or U10884 (N_10884,N_10552,N_10678);
xor U10885 (N_10885,N_10604,N_10783);
nand U10886 (N_10886,N_10596,N_10752);
nand U10887 (N_10887,N_10617,N_10775);
xor U10888 (N_10888,N_10714,N_10620);
or U10889 (N_10889,N_10516,N_10665);
nand U10890 (N_10890,N_10694,N_10760);
nand U10891 (N_10891,N_10652,N_10727);
and U10892 (N_10892,N_10730,N_10544);
xor U10893 (N_10893,N_10798,N_10702);
and U10894 (N_10894,N_10586,N_10757);
nor U10895 (N_10895,N_10713,N_10546);
nor U10896 (N_10896,N_10764,N_10686);
nor U10897 (N_10897,N_10735,N_10567);
xor U10898 (N_10898,N_10708,N_10739);
nand U10899 (N_10899,N_10554,N_10565);
nand U10900 (N_10900,N_10622,N_10508);
xor U10901 (N_10901,N_10614,N_10672);
nor U10902 (N_10902,N_10572,N_10648);
or U10903 (N_10903,N_10559,N_10509);
nor U10904 (N_10904,N_10539,N_10632);
nor U10905 (N_10905,N_10728,N_10522);
nand U10906 (N_10906,N_10654,N_10557);
xnor U10907 (N_10907,N_10524,N_10724);
xor U10908 (N_10908,N_10677,N_10669);
xnor U10909 (N_10909,N_10577,N_10593);
xnor U10910 (N_10910,N_10601,N_10583);
nor U10911 (N_10911,N_10722,N_10779);
xnor U10912 (N_10912,N_10526,N_10777);
xnor U10913 (N_10913,N_10603,N_10521);
xor U10914 (N_10914,N_10625,N_10611);
and U10915 (N_10915,N_10699,N_10505);
nand U10916 (N_10916,N_10561,N_10540);
xor U10917 (N_10917,N_10535,N_10649);
nand U10918 (N_10918,N_10626,N_10676);
xor U10919 (N_10919,N_10744,N_10573);
and U10920 (N_10920,N_10765,N_10675);
nand U10921 (N_10921,N_10738,N_10645);
and U10922 (N_10922,N_10745,N_10723);
nand U10923 (N_10923,N_10517,N_10575);
and U10924 (N_10924,N_10787,N_10697);
nor U10925 (N_10925,N_10768,N_10650);
nor U10926 (N_10926,N_10589,N_10688);
xor U10927 (N_10927,N_10520,N_10619);
nor U10928 (N_10928,N_10703,N_10536);
or U10929 (N_10929,N_10717,N_10550);
nor U10930 (N_10930,N_10754,N_10530);
nor U10931 (N_10931,N_10515,N_10592);
nand U10932 (N_10932,N_10609,N_10580);
nor U10933 (N_10933,N_10588,N_10635);
or U10934 (N_10934,N_10690,N_10780);
or U10935 (N_10935,N_10657,N_10519);
and U10936 (N_10936,N_10640,N_10553);
and U10937 (N_10937,N_10726,N_10590);
nand U10938 (N_10938,N_10796,N_10500);
and U10939 (N_10939,N_10788,N_10570);
xor U10940 (N_10940,N_10692,N_10755);
or U10941 (N_10941,N_10729,N_10769);
nor U10942 (N_10942,N_10628,N_10608);
nand U10943 (N_10943,N_10700,N_10503);
xnor U10944 (N_10944,N_10701,N_10673);
nor U10945 (N_10945,N_10737,N_10715);
nand U10946 (N_10946,N_10511,N_10732);
xor U10947 (N_10947,N_10771,N_10579);
nand U10948 (N_10948,N_10525,N_10600);
or U10949 (N_10949,N_10627,N_10691);
or U10950 (N_10950,N_10654,N_10623);
nor U10951 (N_10951,N_10669,N_10647);
xnor U10952 (N_10952,N_10575,N_10562);
xor U10953 (N_10953,N_10641,N_10506);
nand U10954 (N_10954,N_10716,N_10657);
xnor U10955 (N_10955,N_10567,N_10633);
xnor U10956 (N_10956,N_10526,N_10680);
nand U10957 (N_10957,N_10701,N_10689);
or U10958 (N_10958,N_10738,N_10768);
nand U10959 (N_10959,N_10606,N_10524);
xor U10960 (N_10960,N_10741,N_10586);
xnor U10961 (N_10961,N_10693,N_10719);
or U10962 (N_10962,N_10576,N_10612);
xor U10963 (N_10963,N_10671,N_10659);
and U10964 (N_10964,N_10641,N_10692);
xor U10965 (N_10965,N_10608,N_10549);
xnor U10966 (N_10966,N_10742,N_10760);
or U10967 (N_10967,N_10662,N_10764);
or U10968 (N_10968,N_10567,N_10578);
or U10969 (N_10969,N_10578,N_10620);
xnor U10970 (N_10970,N_10741,N_10519);
and U10971 (N_10971,N_10785,N_10614);
nor U10972 (N_10972,N_10697,N_10774);
or U10973 (N_10973,N_10546,N_10538);
or U10974 (N_10974,N_10629,N_10711);
and U10975 (N_10975,N_10645,N_10565);
or U10976 (N_10976,N_10627,N_10558);
nand U10977 (N_10977,N_10566,N_10540);
nor U10978 (N_10978,N_10771,N_10693);
nor U10979 (N_10979,N_10648,N_10749);
or U10980 (N_10980,N_10620,N_10552);
nand U10981 (N_10981,N_10684,N_10706);
nor U10982 (N_10982,N_10737,N_10630);
or U10983 (N_10983,N_10616,N_10531);
nand U10984 (N_10984,N_10702,N_10680);
and U10985 (N_10985,N_10606,N_10764);
or U10986 (N_10986,N_10609,N_10595);
nand U10987 (N_10987,N_10585,N_10652);
or U10988 (N_10988,N_10797,N_10554);
xnor U10989 (N_10989,N_10598,N_10685);
xor U10990 (N_10990,N_10688,N_10584);
nand U10991 (N_10991,N_10752,N_10733);
nand U10992 (N_10992,N_10667,N_10709);
xnor U10993 (N_10993,N_10793,N_10706);
nand U10994 (N_10994,N_10734,N_10671);
and U10995 (N_10995,N_10686,N_10748);
nor U10996 (N_10996,N_10576,N_10670);
nand U10997 (N_10997,N_10717,N_10627);
nor U10998 (N_10998,N_10756,N_10713);
or U10999 (N_10999,N_10561,N_10706);
and U11000 (N_11000,N_10712,N_10536);
or U11001 (N_11001,N_10700,N_10735);
xnor U11002 (N_11002,N_10773,N_10641);
nor U11003 (N_11003,N_10526,N_10543);
nor U11004 (N_11004,N_10507,N_10595);
nand U11005 (N_11005,N_10794,N_10730);
or U11006 (N_11006,N_10501,N_10634);
nor U11007 (N_11007,N_10745,N_10779);
and U11008 (N_11008,N_10752,N_10736);
xor U11009 (N_11009,N_10583,N_10726);
or U11010 (N_11010,N_10753,N_10695);
nor U11011 (N_11011,N_10605,N_10692);
or U11012 (N_11012,N_10625,N_10678);
nand U11013 (N_11013,N_10767,N_10683);
nor U11014 (N_11014,N_10597,N_10746);
nor U11015 (N_11015,N_10531,N_10789);
nand U11016 (N_11016,N_10766,N_10677);
nor U11017 (N_11017,N_10696,N_10613);
nor U11018 (N_11018,N_10597,N_10522);
nor U11019 (N_11019,N_10677,N_10635);
and U11020 (N_11020,N_10615,N_10643);
nand U11021 (N_11021,N_10603,N_10524);
nor U11022 (N_11022,N_10636,N_10717);
or U11023 (N_11023,N_10689,N_10640);
nor U11024 (N_11024,N_10775,N_10721);
nand U11025 (N_11025,N_10717,N_10707);
xor U11026 (N_11026,N_10640,N_10673);
or U11027 (N_11027,N_10764,N_10584);
nor U11028 (N_11028,N_10757,N_10572);
or U11029 (N_11029,N_10665,N_10709);
or U11030 (N_11030,N_10786,N_10746);
or U11031 (N_11031,N_10542,N_10566);
nand U11032 (N_11032,N_10508,N_10643);
or U11033 (N_11033,N_10685,N_10632);
nand U11034 (N_11034,N_10783,N_10523);
and U11035 (N_11035,N_10708,N_10754);
nor U11036 (N_11036,N_10680,N_10654);
nor U11037 (N_11037,N_10518,N_10696);
or U11038 (N_11038,N_10673,N_10688);
xnor U11039 (N_11039,N_10626,N_10640);
nand U11040 (N_11040,N_10667,N_10511);
or U11041 (N_11041,N_10689,N_10604);
nand U11042 (N_11042,N_10516,N_10722);
xnor U11043 (N_11043,N_10680,N_10606);
or U11044 (N_11044,N_10730,N_10646);
and U11045 (N_11045,N_10773,N_10696);
or U11046 (N_11046,N_10745,N_10736);
or U11047 (N_11047,N_10568,N_10523);
or U11048 (N_11048,N_10560,N_10777);
or U11049 (N_11049,N_10500,N_10690);
and U11050 (N_11050,N_10748,N_10703);
xnor U11051 (N_11051,N_10740,N_10569);
nand U11052 (N_11052,N_10753,N_10784);
and U11053 (N_11053,N_10635,N_10726);
and U11054 (N_11054,N_10683,N_10613);
nor U11055 (N_11055,N_10777,N_10562);
and U11056 (N_11056,N_10535,N_10580);
and U11057 (N_11057,N_10688,N_10773);
and U11058 (N_11058,N_10730,N_10537);
nand U11059 (N_11059,N_10722,N_10730);
xnor U11060 (N_11060,N_10558,N_10690);
or U11061 (N_11061,N_10664,N_10615);
or U11062 (N_11062,N_10723,N_10772);
or U11063 (N_11063,N_10650,N_10593);
or U11064 (N_11064,N_10613,N_10532);
or U11065 (N_11065,N_10764,N_10657);
nor U11066 (N_11066,N_10660,N_10767);
or U11067 (N_11067,N_10753,N_10655);
or U11068 (N_11068,N_10734,N_10788);
nand U11069 (N_11069,N_10503,N_10538);
or U11070 (N_11070,N_10630,N_10573);
nor U11071 (N_11071,N_10553,N_10667);
or U11072 (N_11072,N_10738,N_10678);
and U11073 (N_11073,N_10607,N_10564);
or U11074 (N_11074,N_10793,N_10738);
nor U11075 (N_11075,N_10619,N_10761);
nand U11076 (N_11076,N_10782,N_10704);
and U11077 (N_11077,N_10744,N_10606);
nand U11078 (N_11078,N_10612,N_10785);
or U11079 (N_11079,N_10616,N_10727);
nand U11080 (N_11080,N_10585,N_10710);
nor U11081 (N_11081,N_10642,N_10541);
and U11082 (N_11082,N_10753,N_10622);
or U11083 (N_11083,N_10755,N_10584);
or U11084 (N_11084,N_10689,N_10666);
nor U11085 (N_11085,N_10768,N_10568);
xnor U11086 (N_11086,N_10587,N_10678);
or U11087 (N_11087,N_10568,N_10548);
or U11088 (N_11088,N_10693,N_10533);
and U11089 (N_11089,N_10620,N_10712);
xor U11090 (N_11090,N_10584,N_10622);
nand U11091 (N_11091,N_10697,N_10528);
and U11092 (N_11092,N_10664,N_10730);
or U11093 (N_11093,N_10780,N_10680);
nand U11094 (N_11094,N_10510,N_10621);
or U11095 (N_11095,N_10633,N_10627);
or U11096 (N_11096,N_10595,N_10799);
or U11097 (N_11097,N_10778,N_10792);
and U11098 (N_11098,N_10580,N_10611);
or U11099 (N_11099,N_10641,N_10614);
nor U11100 (N_11100,N_10941,N_10993);
nand U11101 (N_11101,N_10929,N_10875);
xor U11102 (N_11102,N_10907,N_10884);
or U11103 (N_11103,N_10822,N_10834);
nand U11104 (N_11104,N_10931,N_10858);
nor U11105 (N_11105,N_10961,N_10901);
nand U11106 (N_11106,N_10878,N_11056);
xnor U11107 (N_11107,N_11010,N_10898);
and U11108 (N_11108,N_11007,N_10915);
or U11109 (N_11109,N_11066,N_11098);
or U11110 (N_11110,N_10853,N_10843);
nor U11111 (N_11111,N_10977,N_11058);
or U11112 (N_11112,N_11083,N_10954);
or U11113 (N_11113,N_10896,N_10827);
nand U11114 (N_11114,N_10900,N_10897);
xor U11115 (N_11115,N_11065,N_11054);
nor U11116 (N_11116,N_10880,N_10862);
xnor U11117 (N_11117,N_10968,N_11078);
or U11118 (N_11118,N_10824,N_11045);
nand U11119 (N_11119,N_10984,N_11042);
nand U11120 (N_11120,N_10925,N_10821);
nand U11121 (N_11121,N_10937,N_11088);
xor U11122 (N_11122,N_10814,N_10947);
or U11123 (N_11123,N_10994,N_10810);
and U11124 (N_11124,N_11055,N_10879);
or U11125 (N_11125,N_10992,N_10913);
nand U11126 (N_11126,N_11034,N_10930);
nor U11127 (N_11127,N_10806,N_10820);
xor U11128 (N_11128,N_11012,N_10870);
nand U11129 (N_11129,N_11024,N_10831);
and U11130 (N_11130,N_10989,N_10894);
nor U11131 (N_11131,N_11046,N_11074);
xor U11132 (N_11132,N_10815,N_11086);
nor U11133 (N_11133,N_11003,N_11026);
nor U11134 (N_11134,N_10852,N_10948);
xnor U11135 (N_11135,N_11038,N_11095);
nand U11136 (N_11136,N_11033,N_11075);
xor U11137 (N_11137,N_10997,N_10916);
or U11138 (N_11138,N_10914,N_11025);
xnor U11139 (N_11139,N_11017,N_10976);
nand U11140 (N_11140,N_10899,N_10813);
or U11141 (N_11141,N_11051,N_11023);
xnor U11142 (N_11142,N_11022,N_10906);
or U11143 (N_11143,N_11006,N_11014);
and U11144 (N_11144,N_11076,N_10848);
xnor U11145 (N_11145,N_10845,N_11087);
nand U11146 (N_11146,N_10982,N_11080);
nand U11147 (N_11147,N_10847,N_10844);
nand U11148 (N_11148,N_10816,N_10933);
and U11149 (N_11149,N_10952,N_10939);
nor U11150 (N_11150,N_10920,N_11037);
xor U11151 (N_11151,N_10974,N_10936);
xor U11152 (N_11152,N_11020,N_10808);
nand U11153 (N_11153,N_11021,N_11002);
xor U11154 (N_11154,N_11069,N_10932);
or U11155 (N_11155,N_10891,N_11072);
and U11156 (N_11156,N_10927,N_10892);
nor U11157 (N_11157,N_10877,N_10972);
nand U11158 (N_11158,N_10842,N_10832);
nand U11159 (N_11159,N_10865,N_10990);
nor U11160 (N_11160,N_11009,N_10800);
nand U11161 (N_11161,N_11067,N_10838);
or U11162 (N_11162,N_11048,N_11068);
xnor U11163 (N_11163,N_10917,N_11000);
nor U11164 (N_11164,N_10826,N_10846);
nor U11165 (N_11165,N_11079,N_10812);
xor U11166 (N_11166,N_10895,N_10985);
nor U11167 (N_11167,N_10918,N_11035);
nor U11168 (N_11168,N_10979,N_10958);
nor U11169 (N_11169,N_10868,N_10955);
nand U11170 (N_11170,N_10825,N_10829);
or U11171 (N_11171,N_10874,N_10871);
nor U11172 (N_11172,N_10887,N_11008);
nor U11173 (N_11173,N_11092,N_11082);
or U11174 (N_11174,N_10801,N_11089);
or U11175 (N_11175,N_10869,N_10882);
nand U11176 (N_11176,N_10908,N_10857);
nor U11177 (N_11177,N_10975,N_11018);
and U11178 (N_11178,N_11084,N_11053);
nor U11179 (N_11179,N_11027,N_11081);
and U11180 (N_11180,N_11005,N_11030);
xor U11181 (N_11181,N_11070,N_10823);
or U11182 (N_11182,N_10873,N_10904);
xnor U11183 (N_11183,N_10943,N_11049);
nand U11184 (N_11184,N_11062,N_11085);
nor U11185 (N_11185,N_10926,N_11063);
nand U11186 (N_11186,N_10851,N_11041);
and U11187 (N_11187,N_10866,N_10995);
xnor U11188 (N_11188,N_11013,N_11077);
and U11189 (N_11189,N_10905,N_10912);
xnor U11190 (N_11190,N_10854,N_10818);
nand U11191 (N_11191,N_10885,N_10945);
and U11192 (N_11192,N_11059,N_10819);
nor U11193 (N_11193,N_10963,N_10940);
xor U11194 (N_11194,N_10950,N_11016);
or U11195 (N_11195,N_10909,N_10978);
nand U11196 (N_11196,N_10923,N_11031);
or U11197 (N_11197,N_11039,N_10910);
nand U11198 (N_11198,N_11015,N_11019);
nand U11199 (N_11199,N_10859,N_10841);
xor U11200 (N_11200,N_10924,N_10964);
nand U11201 (N_11201,N_11073,N_10861);
and U11202 (N_11202,N_10928,N_11094);
nand U11203 (N_11203,N_10942,N_11096);
nor U11204 (N_11204,N_11044,N_10802);
xor U11205 (N_11205,N_10983,N_10863);
xnor U11206 (N_11206,N_11060,N_10957);
nand U11207 (N_11207,N_10856,N_10888);
xnor U11208 (N_11208,N_10998,N_10803);
xor U11209 (N_11209,N_10999,N_10805);
nor U11210 (N_11210,N_11071,N_10973);
xnor U11211 (N_11211,N_10951,N_10876);
or U11212 (N_11212,N_11029,N_11057);
and U11213 (N_11213,N_11004,N_10902);
nand U11214 (N_11214,N_10956,N_10828);
or U11215 (N_11215,N_10969,N_11011);
or U11216 (N_11216,N_10830,N_10967);
nor U11217 (N_11217,N_11052,N_10817);
nand U11218 (N_11218,N_10807,N_10864);
or U11219 (N_11219,N_10881,N_10981);
nor U11220 (N_11220,N_10836,N_10889);
xnor U11221 (N_11221,N_11061,N_11091);
nor U11222 (N_11222,N_11093,N_11099);
nor U11223 (N_11223,N_11047,N_10921);
or U11224 (N_11224,N_11028,N_10855);
nand U11225 (N_11225,N_11043,N_10867);
xor U11226 (N_11226,N_11032,N_10996);
nor U11227 (N_11227,N_10986,N_10835);
or U11228 (N_11228,N_11050,N_10962);
nor U11229 (N_11229,N_10903,N_11040);
and U11230 (N_11230,N_11036,N_10988);
and U11231 (N_11231,N_10833,N_10893);
nor U11232 (N_11232,N_10971,N_10850);
or U11233 (N_11233,N_10872,N_11090);
or U11234 (N_11234,N_10911,N_11097);
xnor U11235 (N_11235,N_11064,N_10811);
nand U11236 (N_11236,N_10944,N_10934);
xnor U11237 (N_11237,N_10987,N_10839);
or U11238 (N_11238,N_10966,N_10991);
nor U11239 (N_11239,N_10980,N_10922);
or U11240 (N_11240,N_10959,N_10935);
nand U11241 (N_11241,N_10804,N_10946);
and U11242 (N_11242,N_10860,N_10965);
and U11243 (N_11243,N_10960,N_10949);
or U11244 (N_11244,N_10938,N_10953);
xnor U11245 (N_11245,N_10837,N_10890);
nor U11246 (N_11246,N_11001,N_10849);
and U11247 (N_11247,N_10883,N_10970);
nor U11248 (N_11248,N_10840,N_10919);
nor U11249 (N_11249,N_10886,N_10809);
or U11250 (N_11250,N_10897,N_10888);
xnor U11251 (N_11251,N_11012,N_10919);
nand U11252 (N_11252,N_10998,N_10996);
and U11253 (N_11253,N_11092,N_10875);
and U11254 (N_11254,N_11014,N_11007);
nor U11255 (N_11255,N_10898,N_11092);
or U11256 (N_11256,N_11093,N_10856);
nor U11257 (N_11257,N_11007,N_10916);
and U11258 (N_11258,N_10898,N_10931);
nor U11259 (N_11259,N_10895,N_10846);
and U11260 (N_11260,N_10834,N_11094);
nor U11261 (N_11261,N_10843,N_11066);
nor U11262 (N_11262,N_10826,N_10993);
or U11263 (N_11263,N_11027,N_11093);
and U11264 (N_11264,N_10850,N_10947);
nand U11265 (N_11265,N_11018,N_10968);
nor U11266 (N_11266,N_11043,N_10827);
nor U11267 (N_11267,N_10872,N_10846);
xnor U11268 (N_11268,N_10953,N_10872);
and U11269 (N_11269,N_10963,N_11091);
or U11270 (N_11270,N_11063,N_10995);
and U11271 (N_11271,N_10821,N_10957);
or U11272 (N_11272,N_11075,N_10895);
nand U11273 (N_11273,N_10988,N_11014);
nor U11274 (N_11274,N_10815,N_11004);
nand U11275 (N_11275,N_11043,N_11074);
nor U11276 (N_11276,N_10852,N_10966);
nand U11277 (N_11277,N_10940,N_11054);
nand U11278 (N_11278,N_10897,N_10914);
xor U11279 (N_11279,N_10833,N_10902);
xor U11280 (N_11280,N_10894,N_10980);
or U11281 (N_11281,N_11079,N_11006);
xnor U11282 (N_11282,N_10885,N_10840);
xor U11283 (N_11283,N_11042,N_10929);
and U11284 (N_11284,N_10976,N_10834);
or U11285 (N_11285,N_10875,N_10842);
nor U11286 (N_11286,N_11014,N_10991);
or U11287 (N_11287,N_10854,N_11002);
xnor U11288 (N_11288,N_10951,N_10862);
and U11289 (N_11289,N_10900,N_11060);
xnor U11290 (N_11290,N_10979,N_10941);
or U11291 (N_11291,N_11073,N_11021);
nand U11292 (N_11292,N_10847,N_10884);
nand U11293 (N_11293,N_10987,N_10836);
xnor U11294 (N_11294,N_10991,N_10857);
and U11295 (N_11295,N_10858,N_10968);
nand U11296 (N_11296,N_10972,N_11047);
and U11297 (N_11297,N_10904,N_10989);
and U11298 (N_11298,N_10994,N_10905);
or U11299 (N_11299,N_11054,N_10854);
nand U11300 (N_11300,N_11023,N_10837);
and U11301 (N_11301,N_11086,N_10934);
xor U11302 (N_11302,N_10897,N_11081);
or U11303 (N_11303,N_11057,N_10836);
xnor U11304 (N_11304,N_10970,N_11061);
nor U11305 (N_11305,N_11020,N_11074);
xor U11306 (N_11306,N_10850,N_11020);
or U11307 (N_11307,N_10921,N_11096);
xor U11308 (N_11308,N_11023,N_10860);
or U11309 (N_11309,N_11049,N_11062);
nand U11310 (N_11310,N_10974,N_10959);
nor U11311 (N_11311,N_10998,N_11068);
or U11312 (N_11312,N_10851,N_10931);
xnor U11313 (N_11313,N_11032,N_10915);
nor U11314 (N_11314,N_11067,N_10849);
xor U11315 (N_11315,N_10854,N_10809);
nor U11316 (N_11316,N_10955,N_11088);
or U11317 (N_11317,N_10947,N_10864);
and U11318 (N_11318,N_10850,N_11009);
xnor U11319 (N_11319,N_10893,N_11018);
nand U11320 (N_11320,N_10960,N_11006);
xor U11321 (N_11321,N_10812,N_11006);
nand U11322 (N_11322,N_11092,N_10887);
or U11323 (N_11323,N_10864,N_10831);
or U11324 (N_11324,N_11080,N_10868);
and U11325 (N_11325,N_10844,N_10957);
and U11326 (N_11326,N_11096,N_11013);
nand U11327 (N_11327,N_10807,N_10928);
or U11328 (N_11328,N_10936,N_10952);
and U11329 (N_11329,N_11088,N_10832);
or U11330 (N_11330,N_10804,N_10832);
nand U11331 (N_11331,N_11036,N_10814);
or U11332 (N_11332,N_10944,N_11055);
or U11333 (N_11333,N_11088,N_10972);
or U11334 (N_11334,N_10922,N_11007);
and U11335 (N_11335,N_10838,N_10994);
nor U11336 (N_11336,N_10887,N_10993);
nand U11337 (N_11337,N_11006,N_11058);
xnor U11338 (N_11338,N_10822,N_11064);
and U11339 (N_11339,N_10982,N_11045);
and U11340 (N_11340,N_10887,N_10847);
nand U11341 (N_11341,N_10920,N_10886);
nor U11342 (N_11342,N_11097,N_11072);
nand U11343 (N_11343,N_10817,N_11092);
or U11344 (N_11344,N_10879,N_10999);
nor U11345 (N_11345,N_10837,N_10813);
and U11346 (N_11346,N_11056,N_11006);
nor U11347 (N_11347,N_11031,N_10819);
nand U11348 (N_11348,N_11058,N_11075);
or U11349 (N_11349,N_11074,N_10994);
xor U11350 (N_11350,N_10958,N_11065);
nand U11351 (N_11351,N_10992,N_10968);
nand U11352 (N_11352,N_10856,N_11014);
or U11353 (N_11353,N_10930,N_10963);
and U11354 (N_11354,N_11028,N_11000);
or U11355 (N_11355,N_10912,N_11090);
and U11356 (N_11356,N_10836,N_11097);
and U11357 (N_11357,N_10933,N_10985);
nand U11358 (N_11358,N_11025,N_10861);
and U11359 (N_11359,N_10811,N_11005);
nor U11360 (N_11360,N_11057,N_10979);
xnor U11361 (N_11361,N_10941,N_10872);
xnor U11362 (N_11362,N_10987,N_10900);
or U11363 (N_11363,N_11075,N_10896);
nor U11364 (N_11364,N_10854,N_10847);
xnor U11365 (N_11365,N_10930,N_10939);
nor U11366 (N_11366,N_10854,N_11089);
nor U11367 (N_11367,N_10985,N_10880);
nand U11368 (N_11368,N_10923,N_10859);
or U11369 (N_11369,N_10944,N_10901);
or U11370 (N_11370,N_11005,N_10810);
xor U11371 (N_11371,N_10810,N_10912);
and U11372 (N_11372,N_11038,N_10935);
or U11373 (N_11373,N_11031,N_10995);
and U11374 (N_11374,N_10809,N_10897);
or U11375 (N_11375,N_10918,N_10962);
nor U11376 (N_11376,N_11087,N_10987);
nor U11377 (N_11377,N_10808,N_10810);
nand U11378 (N_11378,N_10953,N_10919);
or U11379 (N_11379,N_10813,N_10877);
and U11380 (N_11380,N_10886,N_10869);
or U11381 (N_11381,N_10991,N_10962);
nand U11382 (N_11382,N_10912,N_10824);
xor U11383 (N_11383,N_11090,N_10819);
nand U11384 (N_11384,N_10884,N_10976);
nor U11385 (N_11385,N_10893,N_10806);
xor U11386 (N_11386,N_10900,N_10911);
nor U11387 (N_11387,N_10970,N_10951);
or U11388 (N_11388,N_10913,N_10836);
or U11389 (N_11389,N_11083,N_10820);
nor U11390 (N_11390,N_10937,N_11084);
or U11391 (N_11391,N_11072,N_10955);
and U11392 (N_11392,N_11005,N_10927);
nor U11393 (N_11393,N_11045,N_10803);
xnor U11394 (N_11394,N_11047,N_10908);
xor U11395 (N_11395,N_10974,N_10978);
or U11396 (N_11396,N_10986,N_10915);
or U11397 (N_11397,N_10962,N_11029);
or U11398 (N_11398,N_10880,N_10920);
and U11399 (N_11399,N_11085,N_11079);
nand U11400 (N_11400,N_11384,N_11245);
xnor U11401 (N_11401,N_11382,N_11309);
nor U11402 (N_11402,N_11102,N_11291);
nand U11403 (N_11403,N_11208,N_11319);
or U11404 (N_11404,N_11115,N_11399);
xnor U11405 (N_11405,N_11336,N_11355);
or U11406 (N_11406,N_11130,N_11397);
and U11407 (N_11407,N_11368,N_11188);
xor U11408 (N_11408,N_11190,N_11353);
nand U11409 (N_11409,N_11181,N_11221);
nor U11410 (N_11410,N_11392,N_11119);
xor U11411 (N_11411,N_11395,N_11195);
nand U11412 (N_11412,N_11365,N_11151);
xor U11413 (N_11413,N_11379,N_11199);
nor U11414 (N_11414,N_11204,N_11219);
nor U11415 (N_11415,N_11375,N_11105);
nor U11416 (N_11416,N_11376,N_11152);
xnor U11417 (N_11417,N_11344,N_11150);
xnor U11418 (N_11418,N_11183,N_11369);
nor U11419 (N_11419,N_11374,N_11101);
nand U11420 (N_11420,N_11349,N_11301);
or U11421 (N_11421,N_11142,N_11197);
nor U11422 (N_11422,N_11148,N_11149);
xnor U11423 (N_11423,N_11255,N_11371);
or U11424 (N_11424,N_11345,N_11118);
nand U11425 (N_11425,N_11237,N_11220);
or U11426 (N_11426,N_11233,N_11260);
xnor U11427 (N_11427,N_11316,N_11278);
nor U11428 (N_11428,N_11168,N_11164);
and U11429 (N_11429,N_11347,N_11224);
and U11430 (N_11430,N_11289,N_11339);
xor U11431 (N_11431,N_11109,N_11312);
nor U11432 (N_11432,N_11232,N_11111);
or U11433 (N_11433,N_11308,N_11352);
and U11434 (N_11434,N_11240,N_11236);
or U11435 (N_11435,N_11366,N_11331);
nor U11436 (N_11436,N_11172,N_11185);
xnor U11437 (N_11437,N_11228,N_11292);
xnor U11438 (N_11438,N_11315,N_11244);
xnor U11439 (N_11439,N_11145,N_11385);
nor U11440 (N_11440,N_11297,N_11238);
nand U11441 (N_11441,N_11285,N_11173);
nand U11442 (N_11442,N_11362,N_11126);
xnor U11443 (N_11443,N_11351,N_11174);
nand U11444 (N_11444,N_11192,N_11396);
or U11445 (N_11445,N_11112,N_11265);
and U11446 (N_11446,N_11272,N_11212);
nor U11447 (N_11447,N_11227,N_11129);
or U11448 (N_11448,N_11203,N_11180);
and U11449 (N_11449,N_11155,N_11216);
nor U11450 (N_11450,N_11282,N_11193);
nor U11451 (N_11451,N_11377,N_11288);
and U11452 (N_11452,N_11177,N_11393);
nand U11453 (N_11453,N_11171,N_11122);
xor U11454 (N_11454,N_11159,N_11383);
and U11455 (N_11455,N_11218,N_11106);
or U11456 (N_11456,N_11120,N_11348);
nand U11457 (N_11457,N_11225,N_11242);
nand U11458 (N_11458,N_11223,N_11121);
nand U11459 (N_11459,N_11187,N_11100);
xor U11460 (N_11460,N_11104,N_11141);
nor U11461 (N_11461,N_11133,N_11321);
nand U11462 (N_11462,N_11335,N_11350);
and U11463 (N_11463,N_11103,N_11169);
or U11464 (N_11464,N_11367,N_11184);
or U11465 (N_11465,N_11176,N_11378);
xor U11466 (N_11466,N_11196,N_11311);
or U11467 (N_11467,N_11124,N_11189);
or U11468 (N_11468,N_11284,N_11303);
and U11469 (N_11469,N_11323,N_11156);
and U11470 (N_11470,N_11138,N_11146);
nor U11471 (N_11471,N_11370,N_11209);
nand U11472 (N_11472,N_11337,N_11281);
xnor U11473 (N_11473,N_11234,N_11300);
or U11474 (N_11474,N_11324,N_11107);
and U11475 (N_11475,N_11343,N_11267);
or U11476 (N_11476,N_11143,N_11380);
or U11477 (N_11477,N_11162,N_11389);
xor U11478 (N_11478,N_11249,N_11131);
nand U11479 (N_11479,N_11252,N_11259);
or U11480 (N_11480,N_11266,N_11381);
and U11481 (N_11481,N_11137,N_11123);
xnor U11482 (N_11482,N_11334,N_11361);
and U11483 (N_11483,N_11390,N_11276);
nor U11484 (N_11484,N_11214,N_11313);
or U11485 (N_11485,N_11140,N_11128);
nand U11486 (N_11486,N_11298,N_11153);
nor U11487 (N_11487,N_11191,N_11342);
nor U11488 (N_11488,N_11161,N_11170);
nor U11489 (N_11489,N_11269,N_11239);
or U11490 (N_11490,N_11253,N_11201);
and U11491 (N_11491,N_11229,N_11246);
xor U11492 (N_11492,N_11394,N_11340);
or U11493 (N_11493,N_11318,N_11134);
nor U11494 (N_11494,N_11200,N_11206);
xor U11495 (N_11495,N_11283,N_11108);
nand U11496 (N_11496,N_11186,N_11287);
nor U11497 (N_11497,N_11273,N_11296);
nand U11498 (N_11498,N_11317,N_11166);
nand U11499 (N_11499,N_11363,N_11175);
or U11500 (N_11500,N_11299,N_11182);
nand U11501 (N_11501,N_11290,N_11165);
xor U11502 (N_11502,N_11264,N_11198);
nand U11503 (N_11503,N_11320,N_11388);
and U11504 (N_11504,N_11222,N_11277);
and U11505 (N_11505,N_11127,N_11211);
nand U11506 (N_11506,N_11326,N_11274);
or U11507 (N_11507,N_11325,N_11235);
xor U11508 (N_11508,N_11305,N_11357);
or U11509 (N_11509,N_11160,N_11360);
and U11510 (N_11510,N_11330,N_11241);
xnor U11511 (N_11511,N_11125,N_11167);
nand U11512 (N_11512,N_11215,N_11262);
xor U11513 (N_11513,N_11328,N_11194);
and U11514 (N_11514,N_11387,N_11338);
nor U11515 (N_11515,N_11217,N_11202);
nor U11516 (N_11516,N_11286,N_11250);
or U11517 (N_11517,N_11163,N_11144);
or U11518 (N_11518,N_11207,N_11231);
nand U11519 (N_11519,N_11341,N_11256);
nand U11520 (N_11520,N_11294,N_11327);
and U11521 (N_11521,N_11295,N_11398);
nand U11522 (N_11522,N_11307,N_11293);
or U11523 (N_11523,N_11158,N_11114);
or U11524 (N_11524,N_11205,N_11132);
nand U11525 (N_11525,N_11329,N_11248);
and U11526 (N_11526,N_11364,N_11359);
nand U11527 (N_11527,N_11136,N_11270);
nand U11528 (N_11528,N_11280,N_11243);
nor U11529 (N_11529,N_11391,N_11113);
and U11530 (N_11530,N_11302,N_11373);
and U11531 (N_11531,N_11304,N_11257);
nor U11532 (N_11532,N_11356,N_11110);
xor U11533 (N_11533,N_11268,N_11279);
or U11534 (N_11534,N_11346,N_11213);
xnor U11535 (N_11535,N_11258,N_11310);
nand U11536 (N_11536,N_11263,N_11251);
nand U11537 (N_11537,N_11261,N_11254);
and U11538 (N_11538,N_11179,N_11354);
nor U11539 (N_11539,N_11275,N_11386);
nor U11540 (N_11540,N_11314,N_11154);
and U11541 (N_11541,N_11117,N_11139);
or U11542 (N_11542,N_11271,N_11332);
or U11543 (N_11543,N_11147,N_11157);
xnor U11544 (N_11544,N_11333,N_11178);
nand U11545 (N_11545,N_11210,N_11306);
or U11546 (N_11546,N_11116,N_11226);
xor U11547 (N_11547,N_11322,N_11135);
and U11548 (N_11548,N_11358,N_11230);
nand U11549 (N_11549,N_11372,N_11247);
nor U11550 (N_11550,N_11257,N_11370);
or U11551 (N_11551,N_11174,N_11368);
nor U11552 (N_11552,N_11186,N_11283);
nor U11553 (N_11553,N_11270,N_11391);
nand U11554 (N_11554,N_11314,N_11233);
nand U11555 (N_11555,N_11386,N_11282);
and U11556 (N_11556,N_11221,N_11379);
xnor U11557 (N_11557,N_11294,N_11236);
xnor U11558 (N_11558,N_11349,N_11243);
xor U11559 (N_11559,N_11203,N_11214);
or U11560 (N_11560,N_11318,N_11117);
and U11561 (N_11561,N_11190,N_11196);
nor U11562 (N_11562,N_11190,N_11306);
nand U11563 (N_11563,N_11373,N_11257);
and U11564 (N_11564,N_11251,N_11295);
nand U11565 (N_11565,N_11398,N_11292);
xor U11566 (N_11566,N_11109,N_11150);
nand U11567 (N_11567,N_11209,N_11246);
xor U11568 (N_11568,N_11293,N_11181);
and U11569 (N_11569,N_11361,N_11260);
nor U11570 (N_11570,N_11331,N_11232);
or U11571 (N_11571,N_11207,N_11187);
xnor U11572 (N_11572,N_11164,N_11217);
and U11573 (N_11573,N_11373,N_11380);
nand U11574 (N_11574,N_11281,N_11177);
nand U11575 (N_11575,N_11157,N_11332);
nor U11576 (N_11576,N_11268,N_11121);
or U11577 (N_11577,N_11258,N_11380);
and U11578 (N_11578,N_11298,N_11204);
nor U11579 (N_11579,N_11178,N_11375);
and U11580 (N_11580,N_11380,N_11201);
xnor U11581 (N_11581,N_11149,N_11116);
xor U11582 (N_11582,N_11290,N_11195);
nand U11583 (N_11583,N_11348,N_11109);
nor U11584 (N_11584,N_11255,N_11125);
xor U11585 (N_11585,N_11255,N_11101);
xnor U11586 (N_11586,N_11308,N_11223);
nand U11587 (N_11587,N_11348,N_11134);
xor U11588 (N_11588,N_11194,N_11272);
or U11589 (N_11589,N_11133,N_11123);
xor U11590 (N_11590,N_11252,N_11293);
or U11591 (N_11591,N_11271,N_11156);
and U11592 (N_11592,N_11203,N_11311);
nor U11593 (N_11593,N_11279,N_11126);
xor U11594 (N_11594,N_11354,N_11390);
and U11595 (N_11595,N_11373,N_11162);
or U11596 (N_11596,N_11198,N_11233);
nand U11597 (N_11597,N_11356,N_11249);
nor U11598 (N_11598,N_11327,N_11324);
and U11599 (N_11599,N_11323,N_11106);
nor U11600 (N_11600,N_11210,N_11387);
and U11601 (N_11601,N_11103,N_11163);
nand U11602 (N_11602,N_11185,N_11166);
and U11603 (N_11603,N_11278,N_11178);
xor U11604 (N_11604,N_11263,N_11373);
nor U11605 (N_11605,N_11364,N_11350);
nor U11606 (N_11606,N_11339,N_11107);
and U11607 (N_11607,N_11152,N_11111);
xor U11608 (N_11608,N_11277,N_11324);
nand U11609 (N_11609,N_11254,N_11122);
nor U11610 (N_11610,N_11281,N_11328);
or U11611 (N_11611,N_11352,N_11144);
xnor U11612 (N_11612,N_11180,N_11278);
nor U11613 (N_11613,N_11248,N_11108);
or U11614 (N_11614,N_11244,N_11245);
or U11615 (N_11615,N_11210,N_11159);
nor U11616 (N_11616,N_11318,N_11228);
or U11617 (N_11617,N_11101,N_11175);
and U11618 (N_11618,N_11131,N_11333);
xnor U11619 (N_11619,N_11251,N_11201);
nand U11620 (N_11620,N_11372,N_11385);
xnor U11621 (N_11621,N_11318,N_11391);
nand U11622 (N_11622,N_11101,N_11171);
nand U11623 (N_11623,N_11298,N_11380);
nand U11624 (N_11624,N_11157,N_11235);
nand U11625 (N_11625,N_11157,N_11218);
nand U11626 (N_11626,N_11190,N_11102);
and U11627 (N_11627,N_11210,N_11392);
xor U11628 (N_11628,N_11137,N_11146);
nor U11629 (N_11629,N_11383,N_11277);
nand U11630 (N_11630,N_11357,N_11258);
or U11631 (N_11631,N_11369,N_11153);
or U11632 (N_11632,N_11265,N_11130);
nor U11633 (N_11633,N_11238,N_11247);
or U11634 (N_11634,N_11129,N_11289);
xnor U11635 (N_11635,N_11349,N_11334);
and U11636 (N_11636,N_11324,N_11343);
and U11637 (N_11637,N_11247,N_11329);
xor U11638 (N_11638,N_11221,N_11147);
or U11639 (N_11639,N_11150,N_11201);
nand U11640 (N_11640,N_11351,N_11277);
and U11641 (N_11641,N_11363,N_11330);
or U11642 (N_11642,N_11225,N_11238);
nand U11643 (N_11643,N_11106,N_11160);
or U11644 (N_11644,N_11272,N_11371);
and U11645 (N_11645,N_11339,N_11342);
or U11646 (N_11646,N_11315,N_11291);
and U11647 (N_11647,N_11312,N_11224);
nor U11648 (N_11648,N_11285,N_11384);
nor U11649 (N_11649,N_11289,N_11383);
nor U11650 (N_11650,N_11107,N_11168);
and U11651 (N_11651,N_11346,N_11333);
xor U11652 (N_11652,N_11313,N_11376);
xor U11653 (N_11653,N_11210,N_11274);
and U11654 (N_11654,N_11151,N_11123);
xor U11655 (N_11655,N_11347,N_11121);
or U11656 (N_11656,N_11330,N_11370);
nor U11657 (N_11657,N_11199,N_11120);
and U11658 (N_11658,N_11297,N_11302);
nand U11659 (N_11659,N_11342,N_11242);
or U11660 (N_11660,N_11336,N_11133);
or U11661 (N_11661,N_11367,N_11290);
nand U11662 (N_11662,N_11265,N_11383);
xnor U11663 (N_11663,N_11286,N_11366);
or U11664 (N_11664,N_11332,N_11159);
nor U11665 (N_11665,N_11286,N_11240);
nand U11666 (N_11666,N_11210,N_11267);
and U11667 (N_11667,N_11250,N_11201);
or U11668 (N_11668,N_11128,N_11248);
nand U11669 (N_11669,N_11384,N_11272);
and U11670 (N_11670,N_11397,N_11332);
nor U11671 (N_11671,N_11140,N_11312);
or U11672 (N_11672,N_11387,N_11389);
nor U11673 (N_11673,N_11275,N_11153);
nand U11674 (N_11674,N_11323,N_11181);
nand U11675 (N_11675,N_11112,N_11139);
and U11676 (N_11676,N_11372,N_11371);
nor U11677 (N_11677,N_11210,N_11323);
and U11678 (N_11678,N_11126,N_11118);
nand U11679 (N_11679,N_11221,N_11169);
and U11680 (N_11680,N_11202,N_11274);
or U11681 (N_11681,N_11342,N_11271);
nor U11682 (N_11682,N_11198,N_11148);
nand U11683 (N_11683,N_11159,N_11149);
or U11684 (N_11684,N_11161,N_11105);
xnor U11685 (N_11685,N_11110,N_11173);
or U11686 (N_11686,N_11232,N_11202);
or U11687 (N_11687,N_11328,N_11143);
or U11688 (N_11688,N_11173,N_11306);
xnor U11689 (N_11689,N_11212,N_11274);
or U11690 (N_11690,N_11250,N_11209);
xnor U11691 (N_11691,N_11124,N_11324);
or U11692 (N_11692,N_11388,N_11327);
nand U11693 (N_11693,N_11278,N_11301);
nand U11694 (N_11694,N_11371,N_11390);
or U11695 (N_11695,N_11136,N_11193);
nand U11696 (N_11696,N_11116,N_11386);
or U11697 (N_11697,N_11113,N_11260);
or U11698 (N_11698,N_11226,N_11347);
or U11699 (N_11699,N_11191,N_11312);
or U11700 (N_11700,N_11583,N_11663);
nand U11701 (N_11701,N_11535,N_11656);
nand U11702 (N_11702,N_11690,N_11637);
and U11703 (N_11703,N_11476,N_11633);
or U11704 (N_11704,N_11428,N_11657);
xnor U11705 (N_11705,N_11411,N_11480);
xor U11706 (N_11706,N_11668,N_11551);
nor U11707 (N_11707,N_11413,N_11486);
and U11708 (N_11708,N_11481,N_11563);
nand U11709 (N_11709,N_11602,N_11649);
and U11710 (N_11710,N_11542,N_11555);
or U11711 (N_11711,N_11449,N_11658);
xnor U11712 (N_11712,N_11442,N_11462);
nand U11713 (N_11713,N_11628,N_11433);
or U11714 (N_11714,N_11613,N_11660);
xor U11715 (N_11715,N_11648,N_11463);
nor U11716 (N_11716,N_11482,N_11524);
and U11717 (N_11717,N_11694,N_11582);
nor U11718 (N_11718,N_11445,N_11699);
nand U11719 (N_11719,N_11681,N_11508);
and U11720 (N_11720,N_11483,N_11458);
xor U11721 (N_11721,N_11544,N_11609);
nand U11722 (N_11722,N_11568,N_11651);
or U11723 (N_11723,N_11470,N_11503);
or U11724 (N_11724,N_11403,N_11608);
nor U11725 (N_11725,N_11588,N_11565);
and U11726 (N_11726,N_11557,N_11636);
nand U11727 (N_11727,N_11532,N_11467);
and U11728 (N_11728,N_11536,N_11548);
or U11729 (N_11729,N_11621,N_11506);
xnor U11730 (N_11730,N_11641,N_11598);
xor U11731 (N_11731,N_11487,N_11654);
or U11732 (N_11732,N_11491,N_11454);
or U11733 (N_11733,N_11420,N_11473);
xnor U11734 (N_11734,N_11541,N_11591);
and U11735 (N_11735,N_11610,N_11614);
nand U11736 (N_11736,N_11441,N_11484);
and U11737 (N_11737,N_11566,N_11520);
and U11738 (N_11738,N_11502,N_11434);
or U11739 (N_11739,N_11522,N_11404);
nor U11740 (N_11740,N_11422,N_11642);
and U11741 (N_11741,N_11426,N_11465);
or U11742 (N_11742,N_11407,N_11586);
nor U11743 (N_11743,N_11697,N_11488);
nor U11744 (N_11744,N_11647,N_11571);
xnor U11745 (N_11745,N_11564,N_11468);
and U11746 (N_11746,N_11400,N_11490);
nor U11747 (N_11747,N_11479,N_11616);
nand U11748 (N_11748,N_11691,N_11478);
xnor U11749 (N_11749,N_11471,N_11505);
nand U11750 (N_11750,N_11424,N_11494);
or U11751 (N_11751,N_11553,N_11630);
nor U11752 (N_11752,N_11443,N_11450);
nand U11753 (N_11753,N_11528,N_11440);
nor U11754 (N_11754,N_11526,N_11587);
and U11755 (N_11755,N_11688,N_11592);
nand U11756 (N_11756,N_11423,N_11606);
or U11757 (N_11757,N_11416,N_11509);
xor U11758 (N_11758,N_11569,N_11406);
nand U11759 (N_11759,N_11419,N_11597);
xnor U11760 (N_11760,N_11580,N_11599);
nor U11761 (N_11761,N_11550,N_11518);
and U11762 (N_11762,N_11552,N_11575);
xnor U11763 (N_11763,N_11620,N_11601);
xnor U11764 (N_11764,N_11546,N_11497);
nand U11765 (N_11765,N_11639,N_11650);
nand U11766 (N_11766,N_11638,N_11627);
nor U11767 (N_11767,N_11453,N_11659);
xnor U11768 (N_11768,N_11611,N_11579);
and U11769 (N_11769,N_11489,N_11512);
or U11770 (N_11770,N_11644,N_11612);
or U11771 (N_11771,N_11605,N_11417);
and U11772 (N_11772,N_11593,N_11477);
or U11773 (N_11773,N_11448,N_11698);
or U11774 (N_11774,N_11672,N_11686);
or U11775 (N_11775,N_11452,N_11461);
or U11776 (N_11776,N_11673,N_11600);
or U11777 (N_11777,N_11525,N_11678);
and U11778 (N_11778,N_11455,N_11430);
or U11779 (N_11779,N_11435,N_11515);
and U11780 (N_11780,N_11456,N_11472);
nand U11781 (N_11781,N_11572,N_11560);
nor U11782 (N_11782,N_11594,N_11596);
or U11783 (N_11783,N_11695,N_11573);
and U11784 (N_11784,N_11495,N_11653);
xor U11785 (N_11785,N_11671,N_11436);
and U11786 (N_11786,N_11511,N_11410);
xnor U11787 (N_11787,N_11439,N_11415);
xor U11788 (N_11788,N_11603,N_11676);
xnor U11789 (N_11789,N_11577,N_11501);
xor U11790 (N_11790,N_11684,N_11517);
and U11791 (N_11791,N_11492,N_11558);
or U11792 (N_11792,N_11539,N_11519);
nand U11793 (N_11793,N_11619,N_11632);
nor U11794 (N_11794,N_11409,N_11679);
xor U11795 (N_11795,N_11570,N_11554);
and U11796 (N_11796,N_11421,N_11460);
nor U11797 (N_11797,N_11498,N_11635);
and U11798 (N_11798,N_11696,N_11640);
nor U11799 (N_11799,N_11661,N_11561);
xor U11800 (N_11800,N_11590,N_11578);
or U11801 (N_11801,N_11485,N_11674);
or U11802 (N_11802,N_11670,N_11459);
xor U11803 (N_11803,N_11646,N_11624);
nor U11804 (N_11804,N_11581,N_11504);
nand U11805 (N_11805,N_11618,N_11493);
xnor U11806 (N_11806,N_11510,N_11513);
nor U11807 (N_11807,N_11437,N_11427);
xor U11808 (N_11808,N_11567,N_11543);
and U11809 (N_11809,N_11474,N_11446);
nor U11810 (N_11810,N_11444,N_11408);
or U11811 (N_11811,N_11547,N_11425);
nand U11812 (N_11812,N_11652,N_11669);
xor U11813 (N_11813,N_11665,N_11626);
or U11814 (N_11814,N_11514,N_11692);
xor U11815 (N_11815,N_11469,N_11625);
or U11816 (N_11816,N_11538,N_11682);
nor U11817 (N_11817,N_11418,N_11466);
nand U11818 (N_11818,N_11683,N_11500);
nand U11819 (N_11819,N_11529,N_11629);
xor U11820 (N_11820,N_11677,N_11574);
nand U11821 (N_11821,N_11507,N_11405);
and U11822 (N_11822,N_11595,N_11534);
or U11823 (N_11823,N_11431,N_11662);
nor U11824 (N_11824,N_11604,N_11685);
nor U11825 (N_11825,N_11549,N_11631);
xnor U11826 (N_11826,N_11693,N_11589);
nand U11827 (N_11827,N_11556,N_11576);
and U11828 (N_11828,N_11516,N_11607);
and U11829 (N_11829,N_11521,N_11664);
nor U11830 (N_11830,N_11530,N_11689);
xnor U11831 (N_11831,N_11457,N_11523);
nand U11832 (N_11832,N_11402,N_11401);
xor U11833 (N_11833,N_11655,N_11540);
nand U11834 (N_11834,N_11545,N_11562);
nor U11835 (N_11835,N_11687,N_11623);
or U11836 (N_11836,N_11475,N_11622);
xnor U11837 (N_11837,N_11675,N_11667);
and U11838 (N_11838,N_11680,N_11645);
and U11839 (N_11839,N_11531,N_11412);
xnor U11840 (N_11840,N_11429,N_11533);
nand U11841 (N_11841,N_11464,N_11537);
and U11842 (N_11842,N_11414,N_11617);
nand U11843 (N_11843,N_11499,N_11496);
and U11844 (N_11844,N_11584,N_11634);
and U11845 (N_11845,N_11451,N_11615);
nand U11846 (N_11846,N_11585,N_11666);
xnor U11847 (N_11847,N_11527,N_11447);
nor U11848 (N_11848,N_11559,N_11643);
nor U11849 (N_11849,N_11432,N_11438);
xnor U11850 (N_11850,N_11695,N_11522);
and U11851 (N_11851,N_11586,N_11447);
or U11852 (N_11852,N_11608,N_11445);
xor U11853 (N_11853,N_11419,N_11547);
nand U11854 (N_11854,N_11562,N_11592);
xnor U11855 (N_11855,N_11693,N_11663);
nor U11856 (N_11856,N_11438,N_11490);
and U11857 (N_11857,N_11403,N_11627);
and U11858 (N_11858,N_11687,N_11634);
xor U11859 (N_11859,N_11478,N_11400);
nor U11860 (N_11860,N_11538,N_11571);
xor U11861 (N_11861,N_11484,N_11502);
nor U11862 (N_11862,N_11661,N_11473);
nor U11863 (N_11863,N_11472,N_11636);
nand U11864 (N_11864,N_11485,N_11404);
or U11865 (N_11865,N_11443,N_11485);
xor U11866 (N_11866,N_11632,N_11617);
xnor U11867 (N_11867,N_11593,N_11625);
and U11868 (N_11868,N_11693,N_11513);
xor U11869 (N_11869,N_11601,N_11457);
xnor U11870 (N_11870,N_11635,N_11525);
nor U11871 (N_11871,N_11643,N_11511);
nand U11872 (N_11872,N_11547,N_11540);
nand U11873 (N_11873,N_11557,N_11549);
and U11874 (N_11874,N_11488,N_11523);
and U11875 (N_11875,N_11563,N_11471);
or U11876 (N_11876,N_11601,N_11563);
nand U11877 (N_11877,N_11440,N_11537);
nor U11878 (N_11878,N_11631,N_11600);
and U11879 (N_11879,N_11620,N_11561);
nor U11880 (N_11880,N_11611,N_11690);
or U11881 (N_11881,N_11662,N_11553);
nor U11882 (N_11882,N_11451,N_11631);
nand U11883 (N_11883,N_11458,N_11583);
nor U11884 (N_11884,N_11475,N_11636);
or U11885 (N_11885,N_11576,N_11544);
and U11886 (N_11886,N_11485,N_11575);
nand U11887 (N_11887,N_11535,N_11431);
and U11888 (N_11888,N_11531,N_11512);
and U11889 (N_11889,N_11412,N_11600);
nand U11890 (N_11890,N_11587,N_11507);
or U11891 (N_11891,N_11427,N_11459);
nor U11892 (N_11892,N_11624,N_11653);
nor U11893 (N_11893,N_11677,N_11495);
nor U11894 (N_11894,N_11425,N_11578);
xor U11895 (N_11895,N_11653,N_11403);
or U11896 (N_11896,N_11634,N_11627);
nor U11897 (N_11897,N_11410,N_11565);
xnor U11898 (N_11898,N_11422,N_11558);
and U11899 (N_11899,N_11572,N_11557);
and U11900 (N_11900,N_11520,N_11682);
xor U11901 (N_11901,N_11502,N_11671);
or U11902 (N_11902,N_11432,N_11695);
nor U11903 (N_11903,N_11554,N_11685);
xor U11904 (N_11904,N_11435,N_11627);
and U11905 (N_11905,N_11477,N_11603);
and U11906 (N_11906,N_11496,N_11452);
nor U11907 (N_11907,N_11654,N_11652);
or U11908 (N_11908,N_11647,N_11492);
nor U11909 (N_11909,N_11507,N_11541);
and U11910 (N_11910,N_11434,N_11417);
nor U11911 (N_11911,N_11450,N_11612);
nor U11912 (N_11912,N_11462,N_11674);
xnor U11913 (N_11913,N_11586,N_11682);
and U11914 (N_11914,N_11435,N_11601);
or U11915 (N_11915,N_11537,N_11459);
nand U11916 (N_11916,N_11564,N_11550);
and U11917 (N_11917,N_11675,N_11403);
nor U11918 (N_11918,N_11668,N_11431);
xor U11919 (N_11919,N_11422,N_11664);
and U11920 (N_11920,N_11595,N_11410);
nor U11921 (N_11921,N_11441,N_11436);
nor U11922 (N_11922,N_11562,N_11590);
nor U11923 (N_11923,N_11471,N_11556);
nand U11924 (N_11924,N_11660,N_11605);
nand U11925 (N_11925,N_11430,N_11524);
and U11926 (N_11926,N_11586,N_11610);
nand U11927 (N_11927,N_11642,N_11438);
nand U11928 (N_11928,N_11444,N_11498);
and U11929 (N_11929,N_11595,N_11584);
or U11930 (N_11930,N_11403,N_11543);
or U11931 (N_11931,N_11474,N_11593);
and U11932 (N_11932,N_11687,N_11504);
or U11933 (N_11933,N_11582,N_11621);
or U11934 (N_11934,N_11407,N_11577);
or U11935 (N_11935,N_11475,N_11426);
or U11936 (N_11936,N_11569,N_11493);
or U11937 (N_11937,N_11498,N_11686);
xnor U11938 (N_11938,N_11477,N_11410);
or U11939 (N_11939,N_11412,N_11674);
nor U11940 (N_11940,N_11459,N_11465);
nand U11941 (N_11941,N_11449,N_11644);
or U11942 (N_11942,N_11647,N_11568);
nand U11943 (N_11943,N_11656,N_11612);
and U11944 (N_11944,N_11689,N_11436);
and U11945 (N_11945,N_11678,N_11460);
nand U11946 (N_11946,N_11496,N_11601);
and U11947 (N_11947,N_11547,N_11563);
xnor U11948 (N_11948,N_11487,N_11653);
nor U11949 (N_11949,N_11648,N_11617);
and U11950 (N_11950,N_11515,N_11440);
or U11951 (N_11951,N_11526,N_11611);
or U11952 (N_11952,N_11665,N_11590);
and U11953 (N_11953,N_11599,N_11560);
nor U11954 (N_11954,N_11691,N_11422);
nor U11955 (N_11955,N_11508,N_11662);
nor U11956 (N_11956,N_11469,N_11653);
and U11957 (N_11957,N_11542,N_11620);
or U11958 (N_11958,N_11533,N_11653);
nand U11959 (N_11959,N_11470,N_11562);
and U11960 (N_11960,N_11488,N_11403);
or U11961 (N_11961,N_11521,N_11502);
xnor U11962 (N_11962,N_11509,N_11451);
or U11963 (N_11963,N_11444,N_11591);
or U11964 (N_11964,N_11467,N_11509);
or U11965 (N_11965,N_11581,N_11419);
xor U11966 (N_11966,N_11614,N_11412);
nor U11967 (N_11967,N_11620,N_11584);
xnor U11968 (N_11968,N_11444,N_11594);
or U11969 (N_11969,N_11520,N_11580);
nor U11970 (N_11970,N_11587,N_11699);
xor U11971 (N_11971,N_11458,N_11514);
or U11972 (N_11972,N_11470,N_11548);
or U11973 (N_11973,N_11568,N_11515);
and U11974 (N_11974,N_11609,N_11431);
nor U11975 (N_11975,N_11445,N_11636);
nand U11976 (N_11976,N_11588,N_11558);
nand U11977 (N_11977,N_11681,N_11541);
and U11978 (N_11978,N_11468,N_11505);
and U11979 (N_11979,N_11547,N_11607);
or U11980 (N_11980,N_11416,N_11578);
and U11981 (N_11981,N_11541,N_11576);
and U11982 (N_11982,N_11509,N_11437);
nor U11983 (N_11983,N_11560,N_11608);
xnor U11984 (N_11984,N_11603,N_11423);
nor U11985 (N_11985,N_11690,N_11673);
nand U11986 (N_11986,N_11485,N_11570);
nand U11987 (N_11987,N_11619,N_11608);
nor U11988 (N_11988,N_11497,N_11610);
or U11989 (N_11989,N_11564,N_11646);
nor U11990 (N_11990,N_11650,N_11428);
nand U11991 (N_11991,N_11623,N_11436);
nand U11992 (N_11992,N_11528,N_11438);
nand U11993 (N_11993,N_11459,N_11510);
or U11994 (N_11994,N_11561,N_11490);
and U11995 (N_11995,N_11447,N_11453);
nand U11996 (N_11996,N_11448,N_11561);
nor U11997 (N_11997,N_11487,N_11506);
nor U11998 (N_11998,N_11661,N_11673);
xnor U11999 (N_11999,N_11583,N_11481);
or U12000 (N_12000,N_11853,N_11879);
nand U12001 (N_12001,N_11824,N_11725);
nor U12002 (N_12002,N_11781,N_11757);
nor U12003 (N_12003,N_11842,N_11981);
xnor U12004 (N_12004,N_11791,N_11852);
nor U12005 (N_12005,N_11797,N_11802);
or U12006 (N_12006,N_11943,N_11745);
nor U12007 (N_12007,N_11755,N_11987);
and U12008 (N_12008,N_11900,N_11801);
xnor U12009 (N_12009,N_11936,N_11815);
and U12010 (N_12010,N_11971,N_11773);
nor U12011 (N_12011,N_11800,N_11906);
xor U12012 (N_12012,N_11860,N_11847);
and U12013 (N_12013,N_11929,N_11704);
or U12014 (N_12014,N_11703,N_11778);
nor U12015 (N_12015,N_11828,N_11761);
xor U12016 (N_12016,N_11932,N_11804);
or U12017 (N_12017,N_11765,N_11807);
and U12018 (N_12018,N_11892,N_11876);
and U12019 (N_12019,N_11904,N_11899);
or U12020 (N_12020,N_11786,N_11968);
nand U12021 (N_12021,N_11836,N_11949);
nor U12022 (N_12022,N_11808,N_11708);
nor U12023 (N_12023,N_11877,N_11935);
nor U12024 (N_12024,N_11716,N_11942);
or U12025 (N_12025,N_11731,N_11740);
nor U12026 (N_12026,N_11850,N_11839);
xor U12027 (N_12027,N_11809,N_11978);
nand U12028 (N_12028,N_11792,N_11746);
and U12029 (N_12029,N_11795,N_11894);
or U12030 (N_12030,N_11760,N_11835);
xor U12031 (N_12031,N_11991,N_11827);
nor U12032 (N_12032,N_11796,N_11896);
nor U12033 (N_12033,N_11707,N_11831);
xnor U12034 (N_12034,N_11752,N_11709);
or U12035 (N_12035,N_11771,N_11810);
and U12036 (N_12036,N_11864,N_11714);
and U12037 (N_12037,N_11721,N_11710);
nor U12038 (N_12038,N_11733,N_11735);
nand U12039 (N_12039,N_11812,N_11790);
or U12040 (N_12040,N_11846,N_11724);
nand U12041 (N_12041,N_11838,N_11979);
or U12042 (N_12042,N_11890,N_11861);
xnor U12043 (N_12043,N_11723,N_11889);
xor U12044 (N_12044,N_11893,N_11989);
nor U12045 (N_12045,N_11732,N_11884);
nand U12046 (N_12046,N_11762,N_11905);
nor U12047 (N_12047,N_11953,N_11865);
and U12048 (N_12048,N_11806,N_11830);
and U12049 (N_12049,N_11811,N_11867);
or U12050 (N_12050,N_11938,N_11764);
xnor U12051 (N_12051,N_11798,N_11901);
nand U12052 (N_12052,N_11817,N_11998);
or U12053 (N_12053,N_11832,N_11834);
xor U12054 (N_12054,N_11705,N_11754);
xnor U12055 (N_12055,N_11963,N_11756);
nand U12056 (N_12056,N_11758,N_11910);
xnor U12057 (N_12057,N_11854,N_11726);
or U12058 (N_12058,N_11766,N_11931);
nand U12059 (N_12059,N_11921,N_11925);
xnor U12060 (N_12060,N_11888,N_11779);
xor U12061 (N_12061,N_11780,N_11702);
or U12062 (N_12062,N_11950,N_11886);
xor U12063 (N_12063,N_11734,N_11911);
or U12064 (N_12064,N_11934,N_11916);
nor U12065 (N_12065,N_11883,N_11873);
nand U12066 (N_12066,N_11713,N_11887);
nand U12067 (N_12067,N_11872,N_11819);
nand U12068 (N_12068,N_11818,N_11957);
nor U12069 (N_12069,N_11794,N_11776);
or U12070 (N_12070,N_11772,N_11933);
or U12071 (N_12071,N_11767,N_11717);
nor U12072 (N_12072,N_11782,N_11774);
xor U12073 (N_12073,N_11914,N_11826);
xnor U12074 (N_12074,N_11996,N_11898);
and U12075 (N_12075,N_11958,N_11907);
or U12076 (N_12076,N_11737,N_11980);
nand U12077 (N_12077,N_11727,N_11927);
or U12078 (N_12078,N_11912,N_11816);
and U12079 (N_12079,N_11909,N_11753);
nor U12080 (N_12080,N_11730,N_11833);
xor U12081 (N_12081,N_11969,N_11722);
and U12082 (N_12082,N_11859,N_11701);
nor U12083 (N_12083,N_11928,N_11769);
nand U12084 (N_12084,N_11881,N_11903);
and U12085 (N_12085,N_11982,N_11729);
or U12086 (N_12086,N_11706,N_11744);
xor U12087 (N_12087,N_11777,N_11851);
xnor U12088 (N_12088,N_11885,N_11870);
or U12089 (N_12089,N_11857,N_11895);
nor U12090 (N_12090,N_11937,N_11995);
nor U12091 (N_12091,N_11997,N_11915);
nor U12092 (N_12092,N_11700,N_11858);
and U12093 (N_12093,N_11719,N_11965);
and U12094 (N_12094,N_11820,N_11992);
nand U12095 (N_12095,N_11803,N_11742);
nand U12096 (N_12096,N_11902,N_11952);
or U12097 (N_12097,N_11947,N_11974);
nor U12098 (N_12098,N_11825,N_11941);
nand U12099 (N_12099,N_11964,N_11959);
nand U12100 (N_12100,N_11863,N_11994);
and U12101 (N_12101,N_11967,N_11763);
nor U12102 (N_12102,N_11787,N_11789);
xnor U12103 (N_12103,N_11874,N_11944);
or U12104 (N_12104,N_11954,N_11749);
and U12105 (N_12105,N_11983,N_11882);
or U12106 (N_12106,N_11939,N_11845);
xor U12107 (N_12107,N_11930,N_11720);
xnor U12108 (N_12108,N_11741,N_11821);
nand U12109 (N_12109,N_11750,N_11955);
or U12110 (N_12110,N_11738,N_11822);
nor U12111 (N_12111,N_11948,N_11977);
and U12112 (N_12112,N_11837,N_11962);
nor U12113 (N_12113,N_11813,N_11785);
nor U12114 (N_12114,N_11871,N_11711);
xor U12115 (N_12115,N_11966,N_11926);
nand U12116 (N_12116,N_11840,N_11960);
nand U12117 (N_12117,N_11975,N_11999);
or U12118 (N_12118,N_11751,N_11875);
and U12119 (N_12119,N_11940,N_11951);
and U12120 (N_12120,N_11843,N_11799);
nand U12121 (N_12121,N_11844,N_11759);
nand U12122 (N_12122,N_11973,N_11993);
xor U12123 (N_12123,N_11868,N_11743);
nand U12124 (N_12124,N_11922,N_11918);
xor U12125 (N_12125,N_11985,N_11862);
nand U12126 (N_12126,N_11897,N_11984);
nor U12127 (N_12127,N_11829,N_11793);
or U12128 (N_12128,N_11990,N_11747);
nand U12129 (N_12129,N_11784,N_11768);
nand U12130 (N_12130,N_11972,N_11775);
or U12131 (N_12131,N_11891,N_11823);
nand U12132 (N_12132,N_11748,N_11923);
xnor U12133 (N_12133,N_11986,N_11770);
nand U12134 (N_12134,N_11805,N_11976);
nand U12135 (N_12135,N_11956,N_11783);
or U12136 (N_12136,N_11970,N_11739);
or U12137 (N_12137,N_11924,N_11869);
and U12138 (N_12138,N_11917,N_11878);
nor U12139 (N_12139,N_11961,N_11849);
xnor U12140 (N_12140,N_11841,N_11908);
and U12141 (N_12141,N_11715,N_11736);
and U12142 (N_12142,N_11712,N_11855);
and U12143 (N_12143,N_11880,N_11728);
or U12144 (N_12144,N_11848,N_11919);
and U12145 (N_12145,N_11913,N_11718);
and U12146 (N_12146,N_11945,N_11988);
nand U12147 (N_12147,N_11856,N_11788);
and U12148 (N_12148,N_11946,N_11866);
xnor U12149 (N_12149,N_11814,N_11920);
nor U12150 (N_12150,N_11968,N_11749);
nand U12151 (N_12151,N_11936,N_11917);
and U12152 (N_12152,N_11926,N_11854);
and U12153 (N_12153,N_11762,N_11978);
xnor U12154 (N_12154,N_11977,N_11864);
and U12155 (N_12155,N_11736,N_11931);
nand U12156 (N_12156,N_11722,N_11833);
xor U12157 (N_12157,N_11883,N_11717);
xor U12158 (N_12158,N_11857,N_11878);
and U12159 (N_12159,N_11808,N_11719);
or U12160 (N_12160,N_11853,N_11723);
nand U12161 (N_12161,N_11757,N_11740);
xnor U12162 (N_12162,N_11852,N_11888);
xnor U12163 (N_12163,N_11983,N_11898);
and U12164 (N_12164,N_11943,N_11958);
and U12165 (N_12165,N_11734,N_11841);
and U12166 (N_12166,N_11922,N_11707);
nor U12167 (N_12167,N_11823,N_11864);
nor U12168 (N_12168,N_11830,N_11816);
and U12169 (N_12169,N_11965,N_11928);
and U12170 (N_12170,N_11968,N_11835);
or U12171 (N_12171,N_11824,N_11794);
nand U12172 (N_12172,N_11868,N_11930);
or U12173 (N_12173,N_11809,N_11733);
or U12174 (N_12174,N_11725,N_11726);
and U12175 (N_12175,N_11914,N_11928);
xor U12176 (N_12176,N_11866,N_11822);
or U12177 (N_12177,N_11780,N_11723);
nor U12178 (N_12178,N_11999,N_11925);
nand U12179 (N_12179,N_11905,N_11894);
and U12180 (N_12180,N_11818,N_11811);
and U12181 (N_12181,N_11715,N_11994);
nor U12182 (N_12182,N_11912,N_11808);
and U12183 (N_12183,N_11888,N_11950);
nor U12184 (N_12184,N_11840,N_11714);
or U12185 (N_12185,N_11770,N_11731);
xnor U12186 (N_12186,N_11849,N_11836);
and U12187 (N_12187,N_11910,N_11960);
xnor U12188 (N_12188,N_11910,N_11797);
or U12189 (N_12189,N_11774,N_11909);
or U12190 (N_12190,N_11934,N_11796);
nor U12191 (N_12191,N_11712,N_11844);
nand U12192 (N_12192,N_11792,N_11946);
nand U12193 (N_12193,N_11918,N_11769);
nor U12194 (N_12194,N_11786,N_11959);
or U12195 (N_12195,N_11860,N_11790);
nand U12196 (N_12196,N_11920,N_11707);
xor U12197 (N_12197,N_11740,N_11834);
xor U12198 (N_12198,N_11825,N_11898);
or U12199 (N_12199,N_11849,N_11833);
nand U12200 (N_12200,N_11704,N_11746);
nor U12201 (N_12201,N_11719,N_11701);
or U12202 (N_12202,N_11728,N_11752);
and U12203 (N_12203,N_11819,N_11871);
xor U12204 (N_12204,N_11820,N_11974);
and U12205 (N_12205,N_11872,N_11936);
xor U12206 (N_12206,N_11767,N_11775);
nand U12207 (N_12207,N_11953,N_11788);
nand U12208 (N_12208,N_11727,N_11954);
nor U12209 (N_12209,N_11966,N_11938);
xnor U12210 (N_12210,N_11988,N_11820);
nand U12211 (N_12211,N_11770,N_11873);
and U12212 (N_12212,N_11793,N_11713);
xor U12213 (N_12213,N_11747,N_11807);
nor U12214 (N_12214,N_11749,N_11716);
nand U12215 (N_12215,N_11701,N_11775);
xnor U12216 (N_12216,N_11956,N_11840);
nand U12217 (N_12217,N_11730,N_11961);
and U12218 (N_12218,N_11970,N_11776);
xor U12219 (N_12219,N_11802,N_11813);
xnor U12220 (N_12220,N_11914,N_11866);
and U12221 (N_12221,N_11779,N_11972);
nand U12222 (N_12222,N_11871,N_11747);
or U12223 (N_12223,N_11908,N_11980);
xnor U12224 (N_12224,N_11896,N_11992);
nand U12225 (N_12225,N_11789,N_11859);
nor U12226 (N_12226,N_11848,N_11983);
xnor U12227 (N_12227,N_11742,N_11761);
and U12228 (N_12228,N_11843,N_11885);
xnor U12229 (N_12229,N_11702,N_11819);
nand U12230 (N_12230,N_11756,N_11730);
nor U12231 (N_12231,N_11897,N_11727);
or U12232 (N_12232,N_11801,N_11807);
xor U12233 (N_12233,N_11880,N_11974);
and U12234 (N_12234,N_11792,N_11868);
or U12235 (N_12235,N_11942,N_11856);
or U12236 (N_12236,N_11822,N_11970);
nand U12237 (N_12237,N_11729,N_11977);
or U12238 (N_12238,N_11980,N_11844);
nor U12239 (N_12239,N_11942,N_11971);
nor U12240 (N_12240,N_11849,N_11955);
or U12241 (N_12241,N_11892,N_11950);
nor U12242 (N_12242,N_11955,N_11847);
and U12243 (N_12243,N_11979,N_11937);
nor U12244 (N_12244,N_11963,N_11798);
and U12245 (N_12245,N_11882,N_11869);
or U12246 (N_12246,N_11846,N_11787);
or U12247 (N_12247,N_11975,N_11948);
or U12248 (N_12248,N_11766,N_11904);
nor U12249 (N_12249,N_11792,N_11844);
or U12250 (N_12250,N_11927,N_11728);
nand U12251 (N_12251,N_11797,N_11927);
nor U12252 (N_12252,N_11839,N_11875);
nand U12253 (N_12253,N_11700,N_11975);
and U12254 (N_12254,N_11742,N_11934);
nor U12255 (N_12255,N_11875,N_11739);
or U12256 (N_12256,N_11984,N_11796);
and U12257 (N_12257,N_11998,N_11760);
and U12258 (N_12258,N_11774,N_11804);
nand U12259 (N_12259,N_11715,N_11955);
xor U12260 (N_12260,N_11754,N_11971);
xor U12261 (N_12261,N_11751,N_11802);
nor U12262 (N_12262,N_11834,N_11734);
or U12263 (N_12263,N_11803,N_11798);
or U12264 (N_12264,N_11817,N_11795);
nand U12265 (N_12265,N_11962,N_11752);
nand U12266 (N_12266,N_11744,N_11737);
and U12267 (N_12267,N_11858,N_11854);
or U12268 (N_12268,N_11797,N_11947);
nor U12269 (N_12269,N_11922,N_11957);
and U12270 (N_12270,N_11833,N_11760);
and U12271 (N_12271,N_11797,N_11801);
xnor U12272 (N_12272,N_11932,N_11734);
or U12273 (N_12273,N_11864,N_11881);
and U12274 (N_12274,N_11947,N_11829);
or U12275 (N_12275,N_11879,N_11900);
and U12276 (N_12276,N_11825,N_11815);
or U12277 (N_12277,N_11918,N_11737);
or U12278 (N_12278,N_11755,N_11842);
xnor U12279 (N_12279,N_11988,N_11852);
and U12280 (N_12280,N_11737,N_11960);
nand U12281 (N_12281,N_11800,N_11911);
nor U12282 (N_12282,N_11982,N_11879);
nand U12283 (N_12283,N_11754,N_11944);
nand U12284 (N_12284,N_11900,N_11902);
or U12285 (N_12285,N_11869,N_11839);
or U12286 (N_12286,N_11909,N_11701);
nor U12287 (N_12287,N_11811,N_11873);
and U12288 (N_12288,N_11861,N_11980);
and U12289 (N_12289,N_11951,N_11943);
or U12290 (N_12290,N_11951,N_11892);
nor U12291 (N_12291,N_11749,N_11747);
and U12292 (N_12292,N_11864,N_11880);
nand U12293 (N_12293,N_11913,N_11912);
nor U12294 (N_12294,N_11938,N_11886);
or U12295 (N_12295,N_11711,N_11951);
and U12296 (N_12296,N_11831,N_11778);
nand U12297 (N_12297,N_11786,N_11907);
and U12298 (N_12298,N_11855,N_11982);
nor U12299 (N_12299,N_11767,N_11830);
xnor U12300 (N_12300,N_12266,N_12177);
or U12301 (N_12301,N_12071,N_12053);
and U12302 (N_12302,N_12061,N_12132);
and U12303 (N_12303,N_12058,N_12152);
and U12304 (N_12304,N_12222,N_12005);
and U12305 (N_12305,N_12018,N_12153);
nor U12306 (N_12306,N_12158,N_12011);
nand U12307 (N_12307,N_12259,N_12291);
nor U12308 (N_12308,N_12275,N_12290);
nor U12309 (N_12309,N_12125,N_12032);
xnor U12310 (N_12310,N_12213,N_12164);
nand U12311 (N_12311,N_12134,N_12117);
nand U12312 (N_12312,N_12288,N_12086);
xnor U12313 (N_12313,N_12185,N_12059);
and U12314 (N_12314,N_12150,N_12016);
and U12315 (N_12315,N_12189,N_12127);
xnor U12316 (N_12316,N_12283,N_12039);
xnor U12317 (N_12317,N_12115,N_12129);
or U12318 (N_12318,N_12041,N_12148);
xnor U12319 (N_12319,N_12159,N_12195);
nand U12320 (N_12320,N_12082,N_12237);
and U12321 (N_12321,N_12084,N_12192);
nand U12322 (N_12322,N_12080,N_12253);
xor U12323 (N_12323,N_12285,N_12295);
nor U12324 (N_12324,N_12089,N_12094);
xor U12325 (N_12325,N_12278,N_12293);
and U12326 (N_12326,N_12078,N_12087);
nor U12327 (N_12327,N_12160,N_12104);
or U12328 (N_12328,N_12140,N_12047);
or U12329 (N_12329,N_12157,N_12170);
xor U12330 (N_12330,N_12155,N_12114);
nand U12331 (N_12331,N_12223,N_12046);
nor U12332 (N_12332,N_12135,N_12004);
and U12333 (N_12333,N_12228,N_12179);
or U12334 (N_12334,N_12161,N_12038);
or U12335 (N_12335,N_12027,N_12243);
nor U12336 (N_12336,N_12035,N_12113);
xor U12337 (N_12337,N_12062,N_12050);
and U12338 (N_12338,N_12077,N_12252);
and U12339 (N_12339,N_12128,N_12122);
xor U12340 (N_12340,N_12261,N_12245);
nand U12341 (N_12341,N_12183,N_12240);
nor U12342 (N_12342,N_12067,N_12199);
nand U12343 (N_12343,N_12013,N_12149);
and U12344 (N_12344,N_12001,N_12265);
nand U12345 (N_12345,N_12264,N_12180);
xor U12346 (N_12346,N_12196,N_12145);
xor U12347 (N_12347,N_12219,N_12023);
nor U12348 (N_12348,N_12093,N_12056);
nor U12349 (N_12349,N_12151,N_12028);
xor U12350 (N_12350,N_12099,N_12298);
xor U12351 (N_12351,N_12258,N_12090);
nor U12352 (N_12352,N_12057,N_12108);
or U12353 (N_12353,N_12042,N_12221);
nand U12354 (N_12354,N_12095,N_12244);
and U12355 (N_12355,N_12215,N_12040);
and U12356 (N_12356,N_12015,N_12165);
nor U12357 (N_12357,N_12209,N_12268);
nand U12358 (N_12358,N_12142,N_12247);
or U12359 (N_12359,N_12131,N_12162);
nand U12360 (N_12360,N_12009,N_12019);
or U12361 (N_12361,N_12281,N_12081);
or U12362 (N_12362,N_12097,N_12024);
or U12363 (N_12363,N_12186,N_12141);
nor U12364 (N_12364,N_12200,N_12257);
and U12365 (N_12365,N_12030,N_12188);
xnor U12366 (N_12366,N_12201,N_12230);
nand U12367 (N_12367,N_12226,N_12197);
nand U12368 (N_12368,N_12267,N_12225);
or U12369 (N_12369,N_12103,N_12255);
and U12370 (N_12370,N_12100,N_12048);
or U12371 (N_12371,N_12233,N_12296);
xnor U12372 (N_12372,N_12286,N_12178);
nor U12373 (N_12373,N_12006,N_12212);
xor U12374 (N_12374,N_12144,N_12017);
nand U12375 (N_12375,N_12248,N_12156);
or U12376 (N_12376,N_12294,N_12121);
or U12377 (N_12377,N_12218,N_12075);
nand U12378 (N_12378,N_12069,N_12203);
or U12379 (N_12379,N_12065,N_12064);
nor U12380 (N_12380,N_12014,N_12003);
and U12381 (N_12381,N_12138,N_12169);
nand U12382 (N_12382,N_12299,N_12249);
nor U12383 (N_12383,N_12193,N_12124);
xnor U12384 (N_12384,N_12231,N_12269);
and U12385 (N_12385,N_12175,N_12147);
nand U12386 (N_12386,N_12176,N_12289);
and U12387 (N_12387,N_12284,N_12020);
nand U12388 (N_12388,N_12060,N_12049);
or U12389 (N_12389,N_12098,N_12074);
or U12390 (N_12390,N_12172,N_12234);
nand U12391 (N_12391,N_12068,N_12012);
nor U12392 (N_12392,N_12130,N_12073);
nor U12393 (N_12393,N_12002,N_12214);
xnor U12394 (N_12394,N_12220,N_12119);
and U12395 (N_12395,N_12277,N_12044);
or U12396 (N_12396,N_12204,N_12184);
nand U12397 (N_12397,N_12174,N_12000);
and U12398 (N_12398,N_12292,N_12166);
xnor U12399 (N_12399,N_12181,N_12072);
nor U12400 (N_12400,N_12085,N_12246);
xnor U12401 (N_12401,N_12208,N_12251);
and U12402 (N_12402,N_12045,N_12109);
and U12403 (N_12403,N_12163,N_12139);
and U12404 (N_12404,N_12025,N_12224);
or U12405 (N_12405,N_12271,N_12239);
and U12406 (N_12406,N_12022,N_12194);
or U12407 (N_12407,N_12279,N_12083);
and U12408 (N_12408,N_12173,N_12287);
xnor U12409 (N_12409,N_12101,N_12137);
nor U12410 (N_12410,N_12021,N_12007);
and U12411 (N_12411,N_12182,N_12229);
nor U12412 (N_12412,N_12106,N_12211);
and U12413 (N_12413,N_12051,N_12118);
or U12414 (N_12414,N_12091,N_12054);
nand U12415 (N_12415,N_12241,N_12235);
and U12416 (N_12416,N_12297,N_12254);
nor U12417 (N_12417,N_12205,N_12107);
nand U12418 (N_12418,N_12282,N_12187);
nand U12419 (N_12419,N_12238,N_12043);
nor U12420 (N_12420,N_12171,N_12242);
nand U12421 (N_12421,N_12136,N_12031);
nand U12422 (N_12422,N_12168,N_12262);
nor U12423 (N_12423,N_12273,N_12260);
and U12424 (N_12424,N_12143,N_12198);
nand U12425 (N_12425,N_12102,N_12146);
nor U12426 (N_12426,N_12126,N_12096);
nor U12427 (N_12427,N_12112,N_12088);
nor U12428 (N_12428,N_12008,N_12207);
nor U12429 (N_12429,N_12066,N_12029);
and U12430 (N_12430,N_12116,N_12210);
or U12431 (N_12431,N_12026,N_12133);
and U12432 (N_12432,N_12076,N_12167);
nand U12433 (N_12433,N_12154,N_12010);
xor U12434 (N_12434,N_12274,N_12037);
nand U12435 (N_12435,N_12033,N_12055);
or U12436 (N_12436,N_12227,N_12110);
or U12437 (N_12437,N_12216,N_12280);
and U12438 (N_12438,N_12092,N_12070);
and U12439 (N_12439,N_12111,N_12250);
and U12440 (N_12440,N_12034,N_12206);
nand U12441 (N_12441,N_12191,N_12276);
and U12442 (N_12442,N_12263,N_12052);
nand U12443 (N_12443,N_12236,N_12036);
nand U12444 (N_12444,N_12217,N_12079);
nor U12445 (N_12445,N_12202,N_12256);
nand U12446 (N_12446,N_12123,N_12272);
and U12447 (N_12447,N_12270,N_12105);
nor U12448 (N_12448,N_12120,N_12190);
nand U12449 (N_12449,N_12063,N_12232);
nor U12450 (N_12450,N_12119,N_12219);
and U12451 (N_12451,N_12086,N_12230);
and U12452 (N_12452,N_12035,N_12018);
nand U12453 (N_12453,N_12103,N_12162);
nand U12454 (N_12454,N_12168,N_12012);
nand U12455 (N_12455,N_12174,N_12038);
nor U12456 (N_12456,N_12223,N_12292);
or U12457 (N_12457,N_12023,N_12233);
and U12458 (N_12458,N_12094,N_12261);
xor U12459 (N_12459,N_12206,N_12200);
nor U12460 (N_12460,N_12067,N_12099);
xnor U12461 (N_12461,N_12271,N_12073);
nor U12462 (N_12462,N_12109,N_12024);
xor U12463 (N_12463,N_12002,N_12241);
and U12464 (N_12464,N_12191,N_12104);
or U12465 (N_12465,N_12043,N_12291);
xor U12466 (N_12466,N_12155,N_12158);
or U12467 (N_12467,N_12206,N_12209);
nor U12468 (N_12468,N_12181,N_12273);
nand U12469 (N_12469,N_12216,N_12182);
or U12470 (N_12470,N_12115,N_12159);
and U12471 (N_12471,N_12163,N_12029);
nand U12472 (N_12472,N_12130,N_12179);
or U12473 (N_12473,N_12252,N_12127);
xor U12474 (N_12474,N_12158,N_12137);
and U12475 (N_12475,N_12097,N_12264);
or U12476 (N_12476,N_12254,N_12023);
and U12477 (N_12477,N_12229,N_12177);
nand U12478 (N_12478,N_12008,N_12134);
and U12479 (N_12479,N_12213,N_12137);
nand U12480 (N_12480,N_12289,N_12209);
xor U12481 (N_12481,N_12082,N_12021);
or U12482 (N_12482,N_12207,N_12139);
or U12483 (N_12483,N_12104,N_12209);
or U12484 (N_12484,N_12009,N_12282);
and U12485 (N_12485,N_12047,N_12200);
and U12486 (N_12486,N_12154,N_12173);
xor U12487 (N_12487,N_12118,N_12190);
or U12488 (N_12488,N_12115,N_12009);
xnor U12489 (N_12489,N_12087,N_12005);
nand U12490 (N_12490,N_12157,N_12221);
xor U12491 (N_12491,N_12171,N_12123);
nor U12492 (N_12492,N_12224,N_12218);
and U12493 (N_12493,N_12096,N_12270);
and U12494 (N_12494,N_12116,N_12260);
or U12495 (N_12495,N_12160,N_12126);
or U12496 (N_12496,N_12246,N_12182);
nand U12497 (N_12497,N_12086,N_12060);
or U12498 (N_12498,N_12227,N_12241);
xor U12499 (N_12499,N_12115,N_12256);
xnor U12500 (N_12500,N_12292,N_12209);
and U12501 (N_12501,N_12030,N_12003);
nor U12502 (N_12502,N_12264,N_12268);
or U12503 (N_12503,N_12072,N_12165);
or U12504 (N_12504,N_12166,N_12141);
xor U12505 (N_12505,N_12083,N_12295);
and U12506 (N_12506,N_12064,N_12174);
and U12507 (N_12507,N_12058,N_12168);
or U12508 (N_12508,N_12048,N_12004);
nand U12509 (N_12509,N_12102,N_12085);
xor U12510 (N_12510,N_12020,N_12167);
nand U12511 (N_12511,N_12214,N_12086);
nor U12512 (N_12512,N_12249,N_12175);
or U12513 (N_12513,N_12068,N_12225);
and U12514 (N_12514,N_12227,N_12222);
and U12515 (N_12515,N_12284,N_12001);
nand U12516 (N_12516,N_12011,N_12240);
nor U12517 (N_12517,N_12297,N_12281);
xor U12518 (N_12518,N_12286,N_12203);
nor U12519 (N_12519,N_12096,N_12198);
nor U12520 (N_12520,N_12185,N_12049);
or U12521 (N_12521,N_12115,N_12082);
nor U12522 (N_12522,N_12283,N_12036);
or U12523 (N_12523,N_12292,N_12048);
or U12524 (N_12524,N_12092,N_12034);
and U12525 (N_12525,N_12164,N_12204);
nor U12526 (N_12526,N_12275,N_12112);
and U12527 (N_12527,N_12270,N_12182);
nand U12528 (N_12528,N_12242,N_12265);
xor U12529 (N_12529,N_12209,N_12152);
and U12530 (N_12530,N_12090,N_12048);
xor U12531 (N_12531,N_12166,N_12234);
or U12532 (N_12532,N_12105,N_12127);
xnor U12533 (N_12533,N_12145,N_12042);
xor U12534 (N_12534,N_12243,N_12261);
nand U12535 (N_12535,N_12285,N_12201);
nor U12536 (N_12536,N_12139,N_12013);
or U12537 (N_12537,N_12140,N_12277);
nand U12538 (N_12538,N_12166,N_12238);
nor U12539 (N_12539,N_12181,N_12087);
and U12540 (N_12540,N_12246,N_12159);
xor U12541 (N_12541,N_12290,N_12026);
xnor U12542 (N_12542,N_12114,N_12077);
or U12543 (N_12543,N_12014,N_12287);
or U12544 (N_12544,N_12172,N_12168);
and U12545 (N_12545,N_12020,N_12245);
or U12546 (N_12546,N_12006,N_12070);
nand U12547 (N_12547,N_12158,N_12161);
xnor U12548 (N_12548,N_12270,N_12159);
nand U12549 (N_12549,N_12225,N_12262);
or U12550 (N_12550,N_12230,N_12267);
or U12551 (N_12551,N_12192,N_12167);
nand U12552 (N_12552,N_12271,N_12297);
and U12553 (N_12553,N_12072,N_12244);
or U12554 (N_12554,N_12189,N_12111);
nand U12555 (N_12555,N_12101,N_12230);
xnor U12556 (N_12556,N_12123,N_12092);
nand U12557 (N_12557,N_12145,N_12245);
and U12558 (N_12558,N_12175,N_12018);
xnor U12559 (N_12559,N_12199,N_12068);
xor U12560 (N_12560,N_12099,N_12285);
nor U12561 (N_12561,N_12069,N_12238);
and U12562 (N_12562,N_12205,N_12078);
xor U12563 (N_12563,N_12131,N_12282);
xnor U12564 (N_12564,N_12211,N_12131);
nand U12565 (N_12565,N_12014,N_12063);
nor U12566 (N_12566,N_12292,N_12102);
xnor U12567 (N_12567,N_12154,N_12252);
and U12568 (N_12568,N_12296,N_12054);
or U12569 (N_12569,N_12288,N_12186);
nand U12570 (N_12570,N_12240,N_12190);
or U12571 (N_12571,N_12190,N_12055);
or U12572 (N_12572,N_12228,N_12132);
xor U12573 (N_12573,N_12261,N_12146);
and U12574 (N_12574,N_12002,N_12172);
xnor U12575 (N_12575,N_12057,N_12014);
or U12576 (N_12576,N_12181,N_12020);
and U12577 (N_12577,N_12285,N_12010);
xor U12578 (N_12578,N_12111,N_12038);
xor U12579 (N_12579,N_12014,N_12267);
xnor U12580 (N_12580,N_12031,N_12226);
or U12581 (N_12581,N_12223,N_12050);
xor U12582 (N_12582,N_12182,N_12185);
xnor U12583 (N_12583,N_12021,N_12209);
xnor U12584 (N_12584,N_12181,N_12157);
nand U12585 (N_12585,N_12214,N_12245);
xor U12586 (N_12586,N_12104,N_12111);
and U12587 (N_12587,N_12228,N_12268);
nand U12588 (N_12588,N_12224,N_12195);
or U12589 (N_12589,N_12228,N_12108);
xor U12590 (N_12590,N_12254,N_12136);
or U12591 (N_12591,N_12232,N_12261);
nand U12592 (N_12592,N_12298,N_12115);
or U12593 (N_12593,N_12232,N_12079);
xor U12594 (N_12594,N_12123,N_12217);
nand U12595 (N_12595,N_12054,N_12178);
and U12596 (N_12596,N_12232,N_12120);
nand U12597 (N_12597,N_12030,N_12014);
and U12598 (N_12598,N_12208,N_12010);
nand U12599 (N_12599,N_12057,N_12147);
nor U12600 (N_12600,N_12466,N_12452);
and U12601 (N_12601,N_12430,N_12308);
xor U12602 (N_12602,N_12426,N_12331);
or U12603 (N_12603,N_12310,N_12345);
nand U12604 (N_12604,N_12406,N_12546);
nand U12605 (N_12605,N_12460,N_12459);
xnor U12606 (N_12606,N_12544,N_12312);
xnor U12607 (N_12607,N_12576,N_12375);
nand U12608 (N_12608,N_12487,N_12302);
nor U12609 (N_12609,N_12599,N_12429);
nand U12610 (N_12610,N_12458,N_12450);
or U12611 (N_12611,N_12488,N_12300);
nand U12612 (N_12612,N_12543,N_12314);
nor U12613 (N_12613,N_12542,N_12392);
xnor U12614 (N_12614,N_12579,N_12499);
nor U12615 (N_12615,N_12518,N_12496);
and U12616 (N_12616,N_12322,N_12477);
and U12617 (N_12617,N_12490,N_12573);
nor U12618 (N_12618,N_12332,N_12531);
or U12619 (N_12619,N_12324,N_12386);
xnor U12620 (N_12620,N_12374,N_12507);
and U12621 (N_12621,N_12570,N_12361);
and U12622 (N_12622,N_12524,N_12453);
xnor U12623 (N_12623,N_12328,N_12569);
or U12624 (N_12624,N_12320,N_12355);
or U12625 (N_12625,N_12514,N_12590);
or U12626 (N_12626,N_12319,N_12550);
xnor U12627 (N_12627,N_12420,N_12567);
or U12628 (N_12628,N_12489,N_12306);
and U12629 (N_12629,N_12584,N_12506);
nand U12630 (N_12630,N_12532,N_12373);
and U12631 (N_12631,N_12303,N_12427);
xor U12632 (N_12632,N_12326,N_12538);
nor U12633 (N_12633,N_12582,N_12409);
nor U12634 (N_12634,N_12595,N_12338);
nor U12635 (N_12635,N_12362,N_12365);
xnor U12636 (N_12636,N_12417,N_12434);
or U12637 (N_12637,N_12418,N_12572);
xnor U12638 (N_12638,N_12435,N_12540);
nor U12639 (N_12639,N_12337,N_12333);
nor U12640 (N_12640,N_12554,N_12467);
or U12641 (N_12641,N_12547,N_12335);
nor U12642 (N_12642,N_12353,N_12359);
or U12643 (N_12643,N_12348,N_12433);
xor U12644 (N_12644,N_12393,N_12592);
xor U12645 (N_12645,N_12556,N_12431);
xor U12646 (N_12646,N_12578,N_12405);
nand U12647 (N_12647,N_12384,N_12442);
nand U12648 (N_12648,N_12307,N_12380);
or U12649 (N_12649,N_12372,N_12425);
or U12650 (N_12650,N_12588,N_12415);
and U12651 (N_12651,N_12597,N_12551);
nand U12652 (N_12652,N_12416,N_12493);
or U12653 (N_12653,N_12422,N_12363);
nand U12654 (N_12654,N_12534,N_12457);
xnor U12655 (N_12655,N_12440,N_12502);
xor U12656 (N_12656,N_12521,N_12505);
or U12657 (N_12657,N_12515,N_12399);
nand U12658 (N_12658,N_12545,N_12347);
xor U12659 (N_12659,N_12587,N_12360);
and U12660 (N_12660,N_12456,N_12329);
and U12661 (N_12661,N_12391,N_12471);
and U12662 (N_12662,N_12411,N_12497);
or U12663 (N_12663,N_12321,N_12585);
nor U12664 (N_12664,N_12400,N_12594);
or U12665 (N_12665,N_12313,N_12316);
nor U12666 (N_12666,N_12522,N_12369);
or U12667 (N_12667,N_12356,N_12494);
nand U12668 (N_12668,N_12475,N_12437);
nor U12669 (N_12669,N_12367,N_12454);
xnor U12670 (N_12670,N_12334,N_12473);
nor U12671 (N_12671,N_12564,N_12448);
xnor U12672 (N_12672,N_12401,N_12560);
and U12673 (N_12673,N_12398,N_12589);
or U12674 (N_12674,N_12478,N_12404);
or U12675 (N_12675,N_12461,N_12301);
nand U12676 (N_12676,N_12575,N_12593);
nand U12677 (N_12677,N_12428,N_12526);
nor U12678 (N_12678,N_12424,N_12480);
xor U12679 (N_12679,N_12342,N_12311);
nand U12680 (N_12680,N_12410,N_12346);
or U12681 (N_12681,N_12492,N_12349);
xor U12682 (N_12682,N_12581,N_12381);
nor U12683 (N_12683,N_12451,N_12468);
nand U12684 (N_12684,N_12516,N_12462);
nand U12685 (N_12685,N_12586,N_12414);
or U12686 (N_12686,N_12561,N_12486);
or U12687 (N_12687,N_12533,N_12412);
or U12688 (N_12688,N_12396,N_12423);
xor U12689 (N_12689,N_12555,N_12495);
xor U12690 (N_12690,N_12389,N_12330);
nand U12691 (N_12691,N_12358,N_12571);
or U12692 (N_12692,N_12376,N_12528);
xor U12693 (N_12693,N_12395,N_12541);
xnor U12694 (N_12694,N_12352,N_12583);
nand U12695 (N_12695,N_12323,N_12513);
xor U12696 (N_12696,N_12327,N_12491);
xor U12697 (N_12697,N_12446,N_12336);
nor U12698 (N_12698,N_12378,N_12509);
nand U12699 (N_12699,N_12441,N_12443);
xnor U12700 (N_12700,N_12503,N_12501);
nor U12701 (N_12701,N_12340,N_12383);
xor U12702 (N_12702,N_12562,N_12370);
nor U12703 (N_12703,N_12421,N_12469);
xor U12704 (N_12704,N_12552,N_12481);
and U12705 (N_12705,N_12484,N_12407);
and U12706 (N_12706,N_12563,N_12498);
nor U12707 (N_12707,N_12403,N_12523);
or U12708 (N_12708,N_12596,N_12463);
xor U12709 (N_12709,N_12483,N_12574);
nor U12710 (N_12710,N_12465,N_12402);
nand U12711 (N_12711,N_12485,N_12357);
nand U12712 (N_12712,N_12559,N_12325);
nor U12713 (N_12713,N_12474,N_12510);
nand U12714 (N_12714,N_12444,N_12565);
nor U12715 (N_12715,N_12341,N_12413);
xnor U12716 (N_12716,N_12500,N_12536);
or U12717 (N_12717,N_12476,N_12512);
nand U12718 (N_12718,N_12529,N_12364);
or U12719 (N_12719,N_12371,N_12520);
nand U12720 (N_12720,N_12436,N_12419);
nor U12721 (N_12721,N_12519,N_12504);
or U12722 (N_12722,N_12305,N_12344);
nor U12723 (N_12723,N_12432,N_12447);
and U12724 (N_12724,N_12408,N_12517);
nand U12725 (N_12725,N_12379,N_12598);
nand U12726 (N_12726,N_12455,N_12558);
nor U12727 (N_12727,N_12397,N_12377);
xnor U12728 (N_12728,N_12525,N_12318);
xnor U12729 (N_12729,N_12537,N_12539);
xor U12730 (N_12730,N_12580,N_12354);
or U12731 (N_12731,N_12482,N_12508);
xnor U12732 (N_12732,N_12394,N_12368);
nor U12733 (N_12733,N_12548,N_12350);
or U12734 (N_12734,N_12382,N_12577);
or U12735 (N_12735,N_12464,N_12439);
xor U12736 (N_12736,N_12557,N_12351);
or U12737 (N_12737,N_12472,N_12479);
nor U12738 (N_12738,N_12309,N_12315);
xor U12739 (N_12739,N_12343,N_12449);
and U12740 (N_12740,N_12304,N_12470);
nand U12741 (N_12741,N_12445,N_12390);
nand U12742 (N_12742,N_12530,N_12317);
and U12743 (N_12743,N_12527,N_12366);
nor U12744 (N_12744,N_12438,N_12535);
nor U12745 (N_12745,N_12385,N_12387);
nor U12746 (N_12746,N_12388,N_12566);
nand U12747 (N_12747,N_12511,N_12339);
nor U12748 (N_12748,N_12553,N_12591);
xnor U12749 (N_12749,N_12568,N_12549);
nor U12750 (N_12750,N_12482,N_12464);
nor U12751 (N_12751,N_12330,N_12438);
nor U12752 (N_12752,N_12479,N_12454);
nand U12753 (N_12753,N_12549,N_12590);
or U12754 (N_12754,N_12581,N_12313);
xor U12755 (N_12755,N_12514,N_12303);
or U12756 (N_12756,N_12485,N_12580);
nor U12757 (N_12757,N_12408,N_12380);
xnor U12758 (N_12758,N_12591,N_12377);
or U12759 (N_12759,N_12377,N_12442);
or U12760 (N_12760,N_12457,N_12359);
or U12761 (N_12761,N_12556,N_12490);
nor U12762 (N_12762,N_12560,N_12545);
nand U12763 (N_12763,N_12345,N_12507);
and U12764 (N_12764,N_12502,N_12529);
or U12765 (N_12765,N_12466,N_12519);
and U12766 (N_12766,N_12458,N_12447);
nor U12767 (N_12767,N_12364,N_12325);
or U12768 (N_12768,N_12468,N_12501);
nor U12769 (N_12769,N_12424,N_12470);
nand U12770 (N_12770,N_12562,N_12316);
or U12771 (N_12771,N_12459,N_12349);
nand U12772 (N_12772,N_12499,N_12415);
or U12773 (N_12773,N_12552,N_12528);
nor U12774 (N_12774,N_12525,N_12464);
nor U12775 (N_12775,N_12469,N_12571);
nand U12776 (N_12776,N_12380,N_12365);
nand U12777 (N_12777,N_12329,N_12478);
nand U12778 (N_12778,N_12544,N_12414);
or U12779 (N_12779,N_12568,N_12360);
or U12780 (N_12780,N_12555,N_12499);
or U12781 (N_12781,N_12397,N_12555);
or U12782 (N_12782,N_12479,N_12456);
xor U12783 (N_12783,N_12484,N_12595);
nand U12784 (N_12784,N_12485,N_12510);
or U12785 (N_12785,N_12526,N_12544);
nor U12786 (N_12786,N_12368,N_12504);
xor U12787 (N_12787,N_12488,N_12528);
xor U12788 (N_12788,N_12338,N_12560);
nor U12789 (N_12789,N_12518,N_12388);
or U12790 (N_12790,N_12382,N_12474);
nor U12791 (N_12791,N_12486,N_12339);
or U12792 (N_12792,N_12383,N_12531);
or U12793 (N_12793,N_12520,N_12544);
nand U12794 (N_12794,N_12523,N_12479);
or U12795 (N_12795,N_12329,N_12529);
xor U12796 (N_12796,N_12488,N_12534);
and U12797 (N_12797,N_12487,N_12540);
nor U12798 (N_12798,N_12373,N_12382);
nor U12799 (N_12799,N_12448,N_12477);
and U12800 (N_12800,N_12518,N_12376);
and U12801 (N_12801,N_12359,N_12338);
nand U12802 (N_12802,N_12457,N_12483);
and U12803 (N_12803,N_12316,N_12528);
xor U12804 (N_12804,N_12410,N_12486);
or U12805 (N_12805,N_12351,N_12319);
xor U12806 (N_12806,N_12404,N_12465);
nor U12807 (N_12807,N_12437,N_12425);
nor U12808 (N_12808,N_12510,N_12547);
xor U12809 (N_12809,N_12329,N_12454);
xnor U12810 (N_12810,N_12465,N_12547);
xnor U12811 (N_12811,N_12454,N_12440);
or U12812 (N_12812,N_12529,N_12453);
and U12813 (N_12813,N_12382,N_12566);
or U12814 (N_12814,N_12448,N_12393);
and U12815 (N_12815,N_12488,N_12380);
and U12816 (N_12816,N_12320,N_12526);
xnor U12817 (N_12817,N_12435,N_12414);
nor U12818 (N_12818,N_12501,N_12367);
nor U12819 (N_12819,N_12322,N_12462);
nand U12820 (N_12820,N_12537,N_12374);
xnor U12821 (N_12821,N_12400,N_12396);
xor U12822 (N_12822,N_12317,N_12379);
xnor U12823 (N_12823,N_12350,N_12366);
or U12824 (N_12824,N_12428,N_12382);
nor U12825 (N_12825,N_12334,N_12419);
nand U12826 (N_12826,N_12483,N_12555);
nor U12827 (N_12827,N_12500,N_12433);
or U12828 (N_12828,N_12322,N_12337);
xor U12829 (N_12829,N_12544,N_12461);
xor U12830 (N_12830,N_12568,N_12555);
nor U12831 (N_12831,N_12329,N_12427);
xnor U12832 (N_12832,N_12458,N_12356);
and U12833 (N_12833,N_12589,N_12476);
and U12834 (N_12834,N_12493,N_12464);
nand U12835 (N_12835,N_12530,N_12508);
nor U12836 (N_12836,N_12382,N_12347);
or U12837 (N_12837,N_12302,N_12378);
xnor U12838 (N_12838,N_12469,N_12441);
nor U12839 (N_12839,N_12345,N_12461);
or U12840 (N_12840,N_12473,N_12304);
xnor U12841 (N_12841,N_12480,N_12508);
nor U12842 (N_12842,N_12422,N_12398);
nand U12843 (N_12843,N_12387,N_12533);
and U12844 (N_12844,N_12382,N_12483);
xnor U12845 (N_12845,N_12368,N_12364);
nor U12846 (N_12846,N_12495,N_12519);
and U12847 (N_12847,N_12360,N_12499);
nor U12848 (N_12848,N_12443,N_12335);
nand U12849 (N_12849,N_12560,N_12502);
xor U12850 (N_12850,N_12551,N_12320);
xor U12851 (N_12851,N_12329,N_12564);
xnor U12852 (N_12852,N_12331,N_12455);
or U12853 (N_12853,N_12338,N_12335);
nand U12854 (N_12854,N_12398,N_12321);
nand U12855 (N_12855,N_12310,N_12342);
xnor U12856 (N_12856,N_12495,N_12540);
or U12857 (N_12857,N_12476,N_12354);
xor U12858 (N_12858,N_12535,N_12396);
xor U12859 (N_12859,N_12398,N_12503);
nand U12860 (N_12860,N_12353,N_12365);
nand U12861 (N_12861,N_12552,N_12384);
and U12862 (N_12862,N_12387,N_12451);
nor U12863 (N_12863,N_12377,N_12438);
nand U12864 (N_12864,N_12590,N_12361);
xor U12865 (N_12865,N_12523,N_12496);
xnor U12866 (N_12866,N_12575,N_12567);
and U12867 (N_12867,N_12430,N_12418);
and U12868 (N_12868,N_12558,N_12467);
xor U12869 (N_12869,N_12316,N_12423);
xnor U12870 (N_12870,N_12321,N_12466);
xor U12871 (N_12871,N_12422,N_12508);
nand U12872 (N_12872,N_12451,N_12508);
nand U12873 (N_12873,N_12526,N_12570);
nand U12874 (N_12874,N_12559,N_12445);
nand U12875 (N_12875,N_12445,N_12302);
nor U12876 (N_12876,N_12514,N_12409);
xor U12877 (N_12877,N_12402,N_12316);
xnor U12878 (N_12878,N_12508,N_12426);
nand U12879 (N_12879,N_12410,N_12389);
and U12880 (N_12880,N_12525,N_12455);
xnor U12881 (N_12881,N_12423,N_12438);
nand U12882 (N_12882,N_12527,N_12469);
and U12883 (N_12883,N_12442,N_12443);
xnor U12884 (N_12884,N_12473,N_12324);
xor U12885 (N_12885,N_12429,N_12404);
xor U12886 (N_12886,N_12333,N_12530);
xor U12887 (N_12887,N_12566,N_12350);
nand U12888 (N_12888,N_12319,N_12362);
nand U12889 (N_12889,N_12513,N_12378);
or U12890 (N_12890,N_12344,N_12491);
or U12891 (N_12891,N_12494,N_12592);
and U12892 (N_12892,N_12331,N_12497);
xnor U12893 (N_12893,N_12507,N_12458);
xnor U12894 (N_12894,N_12570,N_12554);
and U12895 (N_12895,N_12595,N_12331);
xnor U12896 (N_12896,N_12580,N_12436);
or U12897 (N_12897,N_12312,N_12457);
nand U12898 (N_12898,N_12348,N_12386);
xor U12899 (N_12899,N_12450,N_12390);
nand U12900 (N_12900,N_12881,N_12632);
nand U12901 (N_12901,N_12743,N_12879);
xnor U12902 (N_12902,N_12660,N_12742);
nor U12903 (N_12903,N_12705,N_12821);
and U12904 (N_12904,N_12624,N_12643);
nand U12905 (N_12905,N_12680,N_12778);
and U12906 (N_12906,N_12806,N_12674);
nor U12907 (N_12907,N_12886,N_12679);
nand U12908 (N_12908,N_12774,N_12759);
nor U12909 (N_12909,N_12761,N_12644);
nor U12910 (N_12910,N_12877,N_12714);
nand U12911 (N_12911,N_12773,N_12736);
or U12912 (N_12912,N_12801,N_12689);
xor U12913 (N_12913,N_12733,N_12861);
or U12914 (N_12914,N_12737,N_12633);
nand U12915 (N_12915,N_12800,N_12809);
nand U12916 (N_12916,N_12751,N_12693);
nand U12917 (N_12917,N_12698,N_12754);
nor U12918 (N_12918,N_12787,N_12716);
and U12919 (N_12919,N_12795,N_12650);
nand U12920 (N_12920,N_12880,N_12889);
nand U12921 (N_12921,N_12649,N_12860);
and U12922 (N_12922,N_12713,N_12615);
xnor U12923 (N_12923,N_12731,N_12709);
or U12924 (N_12924,N_12728,N_12762);
or U12925 (N_12925,N_12882,N_12864);
nor U12926 (N_12926,N_12883,N_12717);
nand U12927 (N_12927,N_12735,N_12625);
nor U12928 (N_12928,N_12600,N_12828);
nor U12929 (N_12929,N_12694,N_12802);
nor U12930 (N_12930,N_12772,N_12617);
nand U12931 (N_12931,N_12606,N_12706);
and U12932 (N_12932,N_12775,N_12872);
xor U12933 (N_12933,N_12642,N_12641);
nor U12934 (N_12934,N_12610,N_12711);
nand U12935 (N_12935,N_12723,N_12843);
and U12936 (N_12936,N_12631,N_12810);
nor U12937 (N_12937,N_12825,N_12760);
nor U12938 (N_12938,N_12823,N_12654);
nor U12939 (N_12939,N_12636,N_12701);
xor U12940 (N_12940,N_12836,N_12747);
xnor U12941 (N_12941,N_12769,N_12893);
xor U12942 (N_12942,N_12620,N_12687);
or U12943 (N_12943,N_12675,N_12831);
and U12944 (N_12944,N_12870,N_12757);
nand U12945 (N_12945,N_12695,N_12673);
xnor U12946 (N_12946,N_12892,N_12653);
and U12947 (N_12947,N_12652,N_12819);
nor U12948 (N_12948,N_12667,N_12637);
nand U12949 (N_12949,N_12865,N_12640);
nor U12950 (N_12950,N_12720,N_12846);
and U12951 (N_12951,N_12797,N_12672);
or U12952 (N_12952,N_12668,N_12876);
xor U12953 (N_12953,N_12718,N_12724);
xor U12954 (N_12954,N_12655,N_12808);
nor U12955 (N_12955,N_12699,N_12715);
or U12956 (N_12956,N_12666,N_12814);
or U12957 (N_12957,N_12692,N_12894);
and U12958 (N_12958,N_12756,N_12722);
nor U12959 (N_12959,N_12734,N_12829);
nand U12960 (N_12960,N_12656,N_12862);
and U12961 (N_12961,N_12885,N_12703);
nor U12962 (N_12962,N_12700,N_12702);
or U12963 (N_12963,N_12779,N_12634);
nor U12964 (N_12964,N_12803,N_12749);
nand U12965 (N_12965,N_12844,N_12868);
xor U12966 (N_12966,N_12837,N_12607);
and U12967 (N_12967,N_12859,N_12627);
and U12968 (N_12968,N_12613,N_12729);
nor U12969 (N_12969,N_12719,N_12758);
nor U12970 (N_12970,N_12708,N_12662);
nand U12971 (N_12971,N_12605,N_12763);
xor U12972 (N_12972,N_12677,N_12875);
and U12973 (N_12973,N_12755,N_12739);
and U12974 (N_12974,N_12834,N_12738);
nor U12975 (N_12975,N_12614,N_12855);
or U12976 (N_12976,N_12852,N_12746);
xor U12977 (N_12977,N_12753,N_12646);
nand U12978 (N_12978,N_12684,N_12833);
xor U12979 (N_12979,N_12826,N_12678);
xnor U12980 (N_12980,N_12616,N_12811);
nand U12981 (N_12981,N_12623,N_12896);
nor U12982 (N_12982,N_12697,N_12847);
nand U12983 (N_12983,N_12869,N_12647);
or U12984 (N_12984,N_12629,N_12794);
and U12985 (N_12985,N_12884,N_12840);
or U12986 (N_12986,N_12820,N_12732);
and U12987 (N_12987,N_12682,N_12845);
nand U12988 (N_12988,N_12765,N_12822);
or U12989 (N_12989,N_12848,N_12804);
nor U12990 (N_12990,N_12628,N_12745);
and U12991 (N_12991,N_12707,N_12665);
or U12992 (N_12992,N_12609,N_12691);
and U12993 (N_12993,N_12657,N_12887);
nor U12994 (N_12994,N_12824,N_12799);
nor U12995 (N_12995,N_12898,N_12807);
or U12996 (N_12996,N_12741,N_12619);
or U12997 (N_12997,N_12663,N_12878);
nor U12998 (N_12998,N_12812,N_12839);
or U12999 (N_12999,N_12788,N_12659);
nor U13000 (N_13000,N_12740,N_12767);
and U13001 (N_13001,N_12651,N_12661);
or U13002 (N_13002,N_12768,N_12770);
xnor U13003 (N_13003,N_12874,N_12602);
and U13004 (N_13004,N_12664,N_12793);
nor U13005 (N_13005,N_12621,N_12601);
xnor U13006 (N_13006,N_12792,N_12780);
and U13007 (N_13007,N_12850,N_12816);
nor U13008 (N_13008,N_12854,N_12781);
nand U13009 (N_13009,N_12842,N_12669);
nand U13010 (N_13010,N_12856,N_12798);
and U13011 (N_13011,N_12863,N_12784);
or U13012 (N_13012,N_12764,N_12890);
and U13013 (N_13013,N_12866,N_12721);
nand U13014 (N_13014,N_12604,N_12608);
nor U13015 (N_13015,N_12670,N_12805);
or U13016 (N_13016,N_12785,N_12766);
or U13017 (N_13017,N_12888,N_12827);
or U13018 (N_13018,N_12899,N_12710);
nand U13019 (N_13019,N_12638,N_12750);
or U13020 (N_13020,N_12635,N_12818);
and U13021 (N_13021,N_12776,N_12838);
nor U13022 (N_13022,N_12835,N_12676);
xnor U13023 (N_13023,N_12752,N_12790);
nand U13024 (N_13024,N_12873,N_12725);
or U13025 (N_13025,N_12671,N_12639);
or U13026 (N_13026,N_12891,N_12832);
and U13027 (N_13027,N_12857,N_12683);
nand U13028 (N_13028,N_12648,N_12696);
xnor U13029 (N_13029,N_12786,N_12690);
nor U13030 (N_13030,N_12688,N_12849);
and U13031 (N_13031,N_12686,N_12871);
and U13032 (N_13032,N_12748,N_12830);
nand U13033 (N_13033,N_12895,N_12685);
nand U13034 (N_13034,N_12853,N_12645);
and U13035 (N_13035,N_12611,N_12841);
xor U13036 (N_13036,N_12727,N_12813);
xnor U13037 (N_13037,N_12771,N_12783);
and U13038 (N_13038,N_12789,N_12817);
or U13039 (N_13039,N_12858,N_12726);
xnor U13040 (N_13040,N_12730,N_12612);
nand U13041 (N_13041,N_12851,N_12782);
or U13042 (N_13042,N_12630,N_12867);
nor U13043 (N_13043,N_12744,N_12681);
or U13044 (N_13044,N_12897,N_12618);
xnor U13045 (N_13045,N_12815,N_12704);
nand U13046 (N_13046,N_12796,N_12658);
nand U13047 (N_13047,N_12712,N_12626);
nor U13048 (N_13048,N_12791,N_12622);
or U13049 (N_13049,N_12777,N_12603);
nor U13050 (N_13050,N_12648,N_12681);
nand U13051 (N_13051,N_12871,N_12865);
xnor U13052 (N_13052,N_12617,N_12802);
xnor U13053 (N_13053,N_12780,N_12685);
or U13054 (N_13054,N_12766,N_12749);
and U13055 (N_13055,N_12795,N_12711);
nor U13056 (N_13056,N_12836,N_12839);
nand U13057 (N_13057,N_12888,N_12697);
and U13058 (N_13058,N_12803,N_12847);
nor U13059 (N_13059,N_12613,N_12823);
nand U13060 (N_13060,N_12626,N_12665);
nand U13061 (N_13061,N_12847,N_12835);
and U13062 (N_13062,N_12677,N_12808);
nand U13063 (N_13063,N_12867,N_12856);
nand U13064 (N_13064,N_12892,N_12870);
nand U13065 (N_13065,N_12666,N_12701);
xor U13066 (N_13066,N_12786,N_12794);
nor U13067 (N_13067,N_12828,N_12741);
and U13068 (N_13068,N_12608,N_12785);
nor U13069 (N_13069,N_12626,N_12722);
nand U13070 (N_13070,N_12775,N_12711);
or U13071 (N_13071,N_12800,N_12885);
or U13072 (N_13072,N_12614,N_12721);
xor U13073 (N_13073,N_12794,N_12622);
nand U13074 (N_13074,N_12650,N_12662);
and U13075 (N_13075,N_12841,N_12886);
nor U13076 (N_13076,N_12886,N_12769);
nor U13077 (N_13077,N_12608,N_12835);
nor U13078 (N_13078,N_12708,N_12644);
nand U13079 (N_13079,N_12859,N_12658);
xor U13080 (N_13080,N_12797,N_12818);
and U13081 (N_13081,N_12729,N_12610);
xor U13082 (N_13082,N_12817,N_12774);
xnor U13083 (N_13083,N_12784,N_12886);
nand U13084 (N_13084,N_12662,N_12702);
or U13085 (N_13085,N_12692,N_12822);
nor U13086 (N_13086,N_12644,N_12635);
xor U13087 (N_13087,N_12746,N_12816);
nand U13088 (N_13088,N_12899,N_12768);
or U13089 (N_13089,N_12832,N_12675);
and U13090 (N_13090,N_12699,N_12745);
nand U13091 (N_13091,N_12694,N_12671);
nand U13092 (N_13092,N_12821,N_12783);
or U13093 (N_13093,N_12779,N_12603);
nor U13094 (N_13094,N_12766,N_12622);
or U13095 (N_13095,N_12778,N_12817);
and U13096 (N_13096,N_12692,N_12823);
or U13097 (N_13097,N_12682,N_12816);
nand U13098 (N_13098,N_12700,N_12736);
or U13099 (N_13099,N_12676,N_12709);
xnor U13100 (N_13100,N_12757,N_12617);
nand U13101 (N_13101,N_12772,N_12782);
nand U13102 (N_13102,N_12625,N_12814);
and U13103 (N_13103,N_12807,N_12733);
or U13104 (N_13104,N_12616,N_12614);
nand U13105 (N_13105,N_12849,N_12791);
nand U13106 (N_13106,N_12609,N_12891);
or U13107 (N_13107,N_12891,N_12656);
and U13108 (N_13108,N_12844,N_12712);
nand U13109 (N_13109,N_12755,N_12849);
nand U13110 (N_13110,N_12887,N_12837);
nor U13111 (N_13111,N_12776,N_12819);
nor U13112 (N_13112,N_12745,N_12851);
xnor U13113 (N_13113,N_12806,N_12845);
nor U13114 (N_13114,N_12809,N_12796);
xor U13115 (N_13115,N_12821,N_12801);
xnor U13116 (N_13116,N_12763,N_12708);
or U13117 (N_13117,N_12629,N_12761);
and U13118 (N_13118,N_12822,N_12768);
nor U13119 (N_13119,N_12620,N_12861);
and U13120 (N_13120,N_12649,N_12620);
or U13121 (N_13121,N_12731,N_12678);
xor U13122 (N_13122,N_12709,N_12740);
and U13123 (N_13123,N_12746,N_12741);
or U13124 (N_13124,N_12730,N_12643);
nor U13125 (N_13125,N_12753,N_12711);
xor U13126 (N_13126,N_12822,N_12796);
xnor U13127 (N_13127,N_12793,N_12622);
xor U13128 (N_13128,N_12862,N_12814);
or U13129 (N_13129,N_12675,N_12694);
or U13130 (N_13130,N_12602,N_12604);
xnor U13131 (N_13131,N_12826,N_12873);
or U13132 (N_13132,N_12664,N_12623);
or U13133 (N_13133,N_12807,N_12773);
nor U13134 (N_13134,N_12636,N_12734);
nor U13135 (N_13135,N_12716,N_12601);
and U13136 (N_13136,N_12686,N_12803);
nor U13137 (N_13137,N_12692,N_12842);
nand U13138 (N_13138,N_12748,N_12757);
and U13139 (N_13139,N_12757,N_12821);
nand U13140 (N_13140,N_12659,N_12813);
or U13141 (N_13141,N_12836,N_12788);
and U13142 (N_13142,N_12628,N_12821);
nor U13143 (N_13143,N_12626,N_12645);
or U13144 (N_13144,N_12751,N_12642);
nor U13145 (N_13145,N_12631,N_12753);
nor U13146 (N_13146,N_12668,N_12715);
xnor U13147 (N_13147,N_12807,N_12863);
or U13148 (N_13148,N_12843,N_12898);
xnor U13149 (N_13149,N_12615,N_12893);
xnor U13150 (N_13150,N_12873,N_12606);
nor U13151 (N_13151,N_12714,N_12602);
and U13152 (N_13152,N_12743,N_12763);
or U13153 (N_13153,N_12620,N_12665);
or U13154 (N_13154,N_12630,N_12784);
or U13155 (N_13155,N_12789,N_12605);
and U13156 (N_13156,N_12822,N_12808);
or U13157 (N_13157,N_12614,N_12895);
and U13158 (N_13158,N_12880,N_12698);
or U13159 (N_13159,N_12828,N_12634);
nor U13160 (N_13160,N_12658,N_12885);
nor U13161 (N_13161,N_12734,N_12768);
or U13162 (N_13162,N_12641,N_12860);
nand U13163 (N_13163,N_12689,N_12879);
nand U13164 (N_13164,N_12794,N_12645);
or U13165 (N_13165,N_12830,N_12633);
nand U13166 (N_13166,N_12811,N_12659);
nand U13167 (N_13167,N_12603,N_12898);
or U13168 (N_13168,N_12791,N_12635);
and U13169 (N_13169,N_12606,N_12790);
nand U13170 (N_13170,N_12665,N_12805);
nand U13171 (N_13171,N_12761,N_12760);
xnor U13172 (N_13172,N_12895,N_12691);
xnor U13173 (N_13173,N_12778,N_12671);
and U13174 (N_13174,N_12865,N_12658);
and U13175 (N_13175,N_12625,N_12801);
or U13176 (N_13176,N_12780,N_12751);
and U13177 (N_13177,N_12692,N_12758);
nand U13178 (N_13178,N_12821,N_12761);
xor U13179 (N_13179,N_12807,N_12748);
nor U13180 (N_13180,N_12852,N_12639);
or U13181 (N_13181,N_12609,N_12762);
nand U13182 (N_13182,N_12773,N_12803);
and U13183 (N_13183,N_12727,N_12797);
and U13184 (N_13184,N_12894,N_12758);
xnor U13185 (N_13185,N_12759,N_12750);
or U13186 (N_13186,N_12785,N_12898);
and U13187 (N_13187,N_12689,N_12830);
and U13188 (N_13188,N_12807,N_12679);
nor U13189 (N_13189,N_12886,N_12891);
nor U13190 (N_13190,N_12839,N_12673);
nand U13191 (N_13191,N_12770,N_12728);
nor U13192 (N_13192,N_12736,N_12878);
or U13193 (N_13193,N_12738,N_12657);
nor U13194 (N_13194,N_12813,N_12683);
xnor U13195 (N_13195,N_12771,N_12852);
or U13196 (N_13196,N_12876,N_12724);
and U13197 (N_13197,N_12669,N_12807);
and U13198 (N_13198,N_12673,N_12819);
or U13199 (N_13199,N_12676,N_12668);
nand U13200 (N_13200,N_13146,N_13129);
nand U13201 (N_13201,N_12990,N_12955);
nor U13202 (N_13202,N_13192,N_12906);
and U13203 (N_13203,N_12975,N_12962);
xnor U13204 (N_13204,N_12945,N_12953);
nor U13205 (N_13205,N_12937,N_12946);
nor U13206 (N_13206,N_12973,N_13041);
xor U13207 (N_13207,N_12986,N_13073);
or U13208 (N_13208,N_13083,N_13104);
nand U13209 (N_13209,N_13124,N_13061);
xnor U13210 (N_13210,N_12964,N_13156);
nor U13211 (N_13211,N_13181,N_13028);
xnor U13212 (N_13212,N_12954,N_13088);
nor U13213 (N_13213,N_12902,N_12949);
and U13214 (N_13214,N_12967,N_13023);
or U13215 (N_13215,N_13021,N_12971);
and U13216 (N_13216,N_13003,N_13172);
nor U13217 (N_13217,N_13011,N_12970);
or U13218 (N_13218,N_12931,N_12935);
or U13219 (N_13219,N_13095,N_12922);
nand U13220 (N_13220,N_13171,N_12929);
xor U13221 (N_13221,N_13043,N_13051);
or U13222 (N_13222,N_13094,N_13036);
and U13223 (N_13223,N_13186,N_13199);
nand U13224 (N_13224,N_12921,N_13064);
nor U13225 (N_13225,N_12996,N_13002);
xnor U13226 (N_13226,N_13044,N_12942);
or U13227 (N_13227,N_12930,N_12920);
or U13228 (N_13228,N_12944,N_13042);
or U13229 (N_13229,N_13089,N_13077);
nor U13230 (N_13230,N_13166,N_12947);
and U13231 (N_13231,N_12941,N_13151);
and U13232 (N_13232,N_12994,N_12968);
nor U13233 (N_13233,N_12903,N_13152);
and U13234 (N_13234,N_12998,N_12991);
nand U13235 (N_13235,N_13062,N_13183);
nor U13236 (N_13236,N_13154,N_13067);
xnor U13237 (N_13237,N_12988,N_13076);
and U13238 (N_13238,N_13001,N_13145);
or U13239 (N_13239,N_13175,N_12983);
or U13240 (N_13240,N_12956,N_13113);
nor U13241 (N_13241,N_13167,N_13159);
nor U13242 (N_13242,N_13096,N_13133);
nand U13243 (N_13243,N_13012,N_13149);
or U13244 (N_13244,N_12904,N_12936);
xor U13245 (N_13245,N_13082,N_13059);
nor U13246 (N_13246,N_13072,N_13138);
or U13247 (N_13247,N_13142,N_13075);
nand U13248 (N_13248,N_13150,N_12976);
or U13249 (N_13249,N_13136,N_13127);
nor U13250 (N_13250,N_12963,N_12982);
or U13251 (N_13251,N_13101,N_13099);
nor U13252 (N_13252,N_12969,N_13045);
nor U13253 (N_13253,N_12995,N_13031);
nor U13254 (N_13254,N_13102,N_13119);
nand U13255 (N_13255,N_13164,N_13087);
nor U13256 (N_13256,N_13126,N_12919);
xor U13257 (N_13257,N_12993,N_13027);
xnor U13258 (N_13258,N_13147,N_12908);
or U13259 (N_13259,N_13118,N_13026);
or U13260 (N_13260,N_13148,N_13110);
or U13261 (N_13261,N_12974,N_13188);
nor U13262 (N_13262,N_12960,N_12959);
nor U13263 (N_13263,N_13141,N_13063);
or U13264 (N_13264,N_13055,N_13137);
or U13265 (N_13265,N_13174,N_13015);
nor U13266 (N_13266,N_13049,N_12957);
nand U13267 (N_13267,N_12928,N_13046);
xor U13268 (N_13268,N_12913,N_13153);
nand U13269 (N_13269,N_13135,N_13013);
nor U13270 (N_13270,N_13157,N_13185);
xnor U13271 (N_13271,N_13165,N_13092);
nand U13272 (N_13272,N_13111,N_13010);
and U13273 (N_13273,N_12992,N_12972);
or U13274 (N_13274,N_12939,N_13018);
nor U13275 (N_13275,N_13070,N_13038);
xor U13276 (N_13276,N_13184,N_13112);
nor U13277 (N_13277,N_13189,N_13019);
or U13278 (N_13278,N_12912,N_13139);
nor U13279 (N_13279,N_13025,N_12905);
nor U13280 (N_13280,N_13056,N_13169);
nand U13281 (N_13281,N_13086,N_13098);
nand U13282 (N_13282,N_13161,N_12977);
nand U13283 (N_13283,N_13140,N_13144);
and U13284 (N_13284,N_13197,N_13080);
or U13285 (N_13285,N_12951,N_13050);
xor U13286 (N_13286,N_13125,N_12984);
nand U13287 (N_13287,N_13115,N_13130);
xnor U13288 (N_13288,N_13106,N_13177);
nor U13289 (N_13289,N_13009,N_13182);
nor U13290 (N_13290,N_13176,N_13120);
nand U13291 (N_13291,N_12926,N_12901);
and U13292 (N_13292,N_13006,N_13093);
nand U13293 (N_13293,N_12943,N_13024);
and U13294 (N_13294,N_12911,N_12938);
nor U13295 (N_13295,N_12979,N_13187);
xnor U13296 (N_13296,N_13065,N_13029);
nand U13297 (N_13297,N_13053,N_13040);
or U13298 (N_13298,N_13179,N_13109);
and U13299 (N_13299,N_13014,N_12989);
nor U13300 (N_13300,N_13100,N_13017);
or U13301 (N_13301,N_12978,N_13091);
nor U13302 (N_13302,N_13121,N_13128);
nor U13303 (N_13303,N_12987,N_12916);
or U13304 (N_13304,N_12910,N_13054);
nor U13305 (N_13305,N_13107,N_13132);
nor U13306 (N_13306,N_13074,N_13016);
and U13307 (N_13307,N_13039,N_13158);
or U13308 (N_13308,N_13057,N_13180);
xnor U13309 (N_13309,N_12914,N_12948);
nand U13310 (N_13310,N_12961,N_13007);
and U13311 (N_13311,N_13020,N_13195);
nor U13312 (N_13312,N_13173,N_13117);
nand U13313 (N_13313,N_13068,N_13162);
or U13314 (N_13314,N_13052,N_13168);
nor U13315 (N_13315,N_13131,N_13170);
nand U13316 (N_13316,N_13097,N_13108);
and U13317 (N_13317,N_13004,N_13078);
or U13318 (N_13318,N_13194,N_13105);
xor U13319 (N_13319,N_12915,N_13060);
and U13320 (N_13320,N_12932,N_13122);
nand U13321 (N_13321,N_12950,N_13033);
nor U13322 (N_13322,N_12981,N_13114);
or U13323 (N_13323,N_13066,N_12907);
nand U13324 (N_13324,N_13035,N_13081);
nor U13325 (N_13325,N_12917,N_13005);
nor U13326 (N_13326,N_13084,N_12927);
nand U13327 (N_13327,N_12918,N_13123);
or U13328 (N_13328,N_12934,N_13103);
nor U13329 (N_13329,N_13193,N_12958);
nor U13330 (N_13330,N_12999,N_13116);
nor U13331 (N_13331,N_12923,N_13032);
nand U13332 (N_13332,N_13178,N_12966);
nand U13333 (N_13333,N_13163,N_12980);
and U13334 (N_13334,N_13022,N_13034);
and U13335 (N_13335,N_13196,N_13000);
or U13336 (N_13336,N_13048,N_12940);
nand U13337 (N_13337,N_13008,N_13198);
or U13338 (N_13338,N_12925,N_13190);
nand U13339 (N_13339,N_13143,N_13134);
nand U13340 (N_13340,N_13160,N_13085);
nand U13341 (N_13341,N_13069,N_12933);
xor U13342 (N_13342,N_12985,N_13155);
or U13343 (N_13343,N_13079,N_12965);
nand U13344 (N_13344,N_12952,N_13047);
nand U13345 (N_13345,N_12997,N_13030);
nor U13346 (N_13346,N_12909,N_13037);
nand U13347 (N_13347,N_12900,N_12924);
or U13348 (N_13348,N_13071,N_13191);
or U13349 (N_13349,N_13090,N_13058);
and U13350 (N_13350,N_13087,N_12909);
and U13351 (N_13351,N_13030,N_13157);
or U13352 (N_13352,N_13116,N_12976);
and U13353 (N_13353,N_12984,N_13028);
and U13354 (N_13354,N_12902,N_12967);
nand U13355 (N_13355,N_13097,N_13189);
and U13356 (N_13356,N_13114,N_12911);
and U13357 (N_13357,N_12999,N_13102);
or U13358 (N_13358,N_13098,N_13067);
nand U13359 (N_13359,N_13120,N_12924);
nand U13360 (N_13360,N_12919,N_13039);
xnor U13361 (N_13361,N_13123,N_12924);
nor U13362 (N_13362,N_13057,N_13124);
nor U13363 (N_13363,N_13113,N_13044);
and U13364 (N_13364,N_13111,N_13047);
or U13365 (N_13365,N_13064,N_13173);
and U13366 (N_13366,N_13162,N_13085);
nor U13367 (N_13367,N_13026,N_13049);
xnor U13368 (N_13368,N_13060,N_13082);
nor U13369 (N_13369,N_13074,N_12926);
nor U13370 (N_13370,N_13190,N_13166);
or U13371 (N_13371,N_13142,N_13020);
nor U13372 (N_13372,N_12924,N_12964);
or U13373 (N_13373,N_12912,N_13025);
and U13374 (N_13374,N_12959,N_12928);
and U13375 (N_13375,N_12955,N_13092);
or U13376 (N_13376,N_13091,N_12970);
nand U13377 (N_13377,N_13154,N_13059);
xnor U13378 (N_13378,N_13175,N_13138);
or U13379 (N_13379,N_13172,N_12913);
nor U13380 (N_13380,N_13093,N_13007);
nor U13381 (N_13381,N_13036,N_12929);
and U13382 (N_13382,N_13112,N_13173);
and U13383 (N_13383,N_12941,N_13092);
and U13384 (N_13384,N_13005,N_13143);
xnor U13385 (N_13385,N_12919,N_12942);
nand U13386 (N_13386,N_13078,N_13157);
nand U13387 (N_13387,N_13157,N_13123);
and U13388 (N_13388,N_13186,N_12979);
nor U13389 (N_13389,N_12946,N_13108);
and U13390 (N_13390,N_13043,N_13166);
and U13391 (N_13391,N_13176,N_12903);
or U13392 (N_13392,N_12985,N_13065);
nand U13393 (N_13393,N_12962,N_13027);
xor U13394 (N_13394,N_13011,N_12982);
nor U13395 (N_13395,N_12908,N_12964);
xor U13396 (N_13396,N_12901,N_12927);
xor U13397 (N_13397,N_13014,N_13070);
and U13398 (N_13398,N_13092,N_13063);
nand U13399 (N_13399,N_13008,N_12997);
nand U13400 (N_13400,N_13112,N_12967);
nor U13401 (N_13401,N_12948,N_13195);
and U13402 (N_13402,N_13157,N_13003);
xnor U13403 (N_13403,N_13004,N_13112);
nor U13404 (N_13404,N_13039,N_13165);
and U13405 (N_13405,N_13180,N_12984);
xnor U13406 (N_13406,N_13030,N_13140);
and U13407 (N_13407,N_13109,N_13077);
and U13408 (N_13408,N_13057,N_13023);
or U13409 (N_13409,N_12954,N_12987);
and U13410 (N_13410,N_12953,N_13122);
nand U13411 (N_13411,N_13053,N_13051);
or U13412 (N_13412,N_13136,N_13163);
and U13413 (N_13413,N_13102,N_13140);
or U13414 (N_13414,N_13042,N_13069);
xnor U13415 (N_13415,N_12999,N_12980);
or U13416 (N_13416,N_13115,N_12912);
or U13417 (N_13417,N_12930,N_12969);
and U13418 (N_13418,N_12951,N_12919);
xnor U13419 (N_13419,N_13064,N_13179);
nand U13420 (N_13420,N_13198,N_13174);
nor U13421 (N_13421,N_13199,N_13054);
nor U13422 (N_13422,N_13139,N_12959);
nand U13423 (N_13423,N_13154,N_13045);
or U13424 (N_13424,N_12915,N_13073);
nor U13425 (N_13425,N_13057,N_12933);
nor U13426 (N_13426,N_13014,N_13163);
xor U13427 (N_13427,N_13017,N_12941);
or U13428 (N_13428,N_13092,N_12982);
or U13429 (N_13429,N_13094,N_13151);
nand U13430 (N_13430,N_13169,N_12925);
nor U13431 (N_13431,N_13041,N_13003);
nor U13432 (N_13432,N_13089,N_13039);
and U13433 (N_13433,N_13190,N_13102);
xnor U13434 (N_13434,N_13155,N_12981);
nand U13435 (N_13435,N_13026,N_13145);
and U13436 (N_13436,N_13085,N_13056);
xnor U13437 (N_13437,N_12925,N_12906);
xor U13438 (N_13438,N_12949,N_13129);
or U13439 (N_13439,N_13010,N_13125);
or U13440 (N_13440,N_13192,N_13006);
xnor U13441 (N_13441,N_13021,N_12989);
nand U13442 (N_13442,N_12931,N_13035);
or U13443 (N_13443,N_13155,N_12972);
xnor U13444 (N_13444,N_12984,N_12975);
nor U13445 (N_13445,N_12916,N_13179);
or U13446 (N_13446,N_13068,N_13143);
and U13447 (N_13447,N_13010,N_12918);
and U13448 (N_13448,N_13091,N_12953);
nor U13449 (N_13449,N_12962,N_13149);
xor U13450 (N_13450,N_12945,N_13012);
or U13451 (N_13451,N_13029,N_13192);
xor U13452 (N_13452,N_13007,N_13010);
and U13453 (N_13453,N_12997,N_13171);
and U13454 (N_13454,N_13067,N_13070);
xor U13455 (N_13455,N_12929,N_12959);
or U13456 (N_13456,N_13027,N_13076);
nand U13457 (N_13457,N_13146,N_13000);
nor U13458 (N_13458,N_13107,N_13129);
nand U13459 (N_13459,N_13079,N_13111);
xnor U13460 (N_13460,N_13035,N_13038);
or U13461 (N_13461,N_12989,N_12933);
or U13462 (N_13462,N_13090,N_13003);
nand U13463 (N_13463,N_13149,N_13128);
xor U13464 (N_13464,N_12967,N_13134);
nor U13465 (N_13465,N_12973,N_13147);
and U13466 (N_13466,N_13034,N_12967);
nand U13467 (N_13467,N_12962,N_13172);
xnor U13468 (N_13468,N_12911,N_13171);
or U13469 (N_13469,N_12930,N_13026);
xnor U13470 (N_13470,N_12938,N_13004);
xnor U13471 (N_13471,N_13173,N_13106);
xor U13472 (N_13472,N_13148,N_12963);
xnor U13473 (N_13473,N_13108,N_12970);
xor U13474 (N_13474,N_12937,N_12961);
xor U13475 (N_13475,N_12995,N_13193);
nor U13476 (N_13476,N_12991,N_12977);
nor U13477 (N_13477,N_12908,N_13044);
xor U13478 (N_13478,N_12934,N_13167);
xor U13479 (N_13479,N_12999,N_12949);
or U13480 (N_13480,N_13023,N_13107);
or U13481 (N_13481,N_13124,N_13019);
or U13482 (N_13482,N_12908,N_13135);
or U13483 (N_13483,N_13137,N_13148);
nor U13484 (N_13484,N_13124,N_13104);
nand U13485 (N_13485,N_13184,N_12948);
and U13486 (N_13486,N_13083,N_12964);
and U13487 (N_13487,N_12964,N_13060);
nor U13488 (N_13488,N_12902,N_12990);
nand U13489 (N_13489,N_13151,N_13153);
nor U13490 (N_13490,N_12913,N_13096);
and U13491 (N_13491,N_12941,N_12919);
and U13492 (N_13492,N_12937,N_13016);
xor U13493 (N_13493,N_13054,N_13036);
or U13494 (N_13494,N_13185,N_13040);
nor U13495 (N_13495,N_13009,N_13199);
xor U13496 (N_13496,N_13052,N_13131);
or U13497 (N_13497,N_13112,N_12926);
or U13498 (N_13498,N_12943,N_12941);
or U13499 (N_13499,N_12912,N_13106);
nand U13500 (N_13500,N_13331,N_13297);
nor U13501 (N_13501,N_13359,N_13279);
nor U13502 (N_13502,N_13233,N_13263);
or U13503 (N_13503,N_13201,N_13282);
xor U13504 (N_13504,N_13290,N_13238);
nor U13505 (N_13505,N_13212,N_13235);
or U13506 (N_13506,N_13473,N_13440);
nand U13507 (N_13507,N_13305,N_13441);
or U13508 (N_13508,N_13484,N_13439);
nand U13509 (N_13509,N_13448,N_13470);
nor U13510 (N_13510,N_13389,N_13291);
xnor U13511 (N_13511,N_13418,N_13320);
nor U13512 (N_13512,N_13458,N_13388);
and U13513 (N_13513,N_13329,N_13343);
nor U13514 (N_13514,N_13295,N_13341);
nor U13515 (N_13515,N_13221,N_13273);
nand U13516 (N_13516,N_13395,N_13365);
xor U13517 (N_13517,N_13317,N_13224);
xor U13518 (N_13518,N_13269,N_13485);
and U13519 (N_13519,N_13385,N_13457);
or U13520 (N_13520,N_13467,N_13299);
xnor U13521 (N_13521,N_13416,N_13257);
xnor U13522 (N_13522,N_13357,N_13475);
or U13523 (N_13523,N_13248,N_13307);
and U13524 (N_13524,N_13276,N_13298);
nand U13525 (N_13525,N_13350,N_13472);
nand U13526 (N_13526,N_13379,N_13227);
xor U13527 (N_13527,N_13446,N_13258);
xor U13528 (N_13528,N_13333,N_13241);
nor U13529 (N_13529,N_13398,N_13362);
xnor U13530 (N_13530,N_13419,N_13351);
xnor U13531 (N_13531,N_13214,N_13391);
nand U13532 (N_13532,N_13490,N_13286);
xnor U13533 (N_13533,N_13468,N_13314);
xnor U13534 (N_13534,N_13427,N_13280);
nor U13535 (N_13535,N_13246,N_13283);
or U13536 (N_13536,N_13355,N_13397);
and U13537 (N_13537,N_13275,N_13219);
and U13538 (N_13538,N_13387,N_13239);
nand U13539 (N_13539,N_13346,N_13431);
or U13540 (N_13540,N_13474,N_13225);
and U13541 (N_13541,N_13375,N_13412);
xnor U13542 (N_13542,N_13373,N_13471);
and U13543 (N_13543,N_13407,N_13464);
nand U13544 (N_13544,N_13376,N_13450);
nor U13545 (N_13545,N_13240,N_13284);
or U13546 (N_13546,N_13211,N_13491);
nand U13547 (N_13547,N_13402,N_13222);
xor U13548 (N_13548,N_13268,N_13368);
nor U13549 (N_13549,N_13361,N_13496);
xnor U13550 (N_13550,N_13334,N_13486);
xor U13551 (N_13551,N_13459,N_13363);
nor U13552 (N_13552,N_13499,N_13344);
nand U13553 (N_13553,N_13330,N_13293);
nor U13554 (N_13554,N_13337,N_13481);
nand U13555 (N_13555,N_13250,N_13345);
xor U13556 (N_13556,N_13444,N_13367);
or U13557 (N_13557,N_13460,N_13423);
xor U13558 (N_13558,N_13281,N_13462);
nor U13559 (N_13559,N_13237,N_13312);
nor U13560 (N_13560,N_13377,N_13354);
xor U13561 (N_13561,N_13452,N_13456);
xnor U13562 (N_13562,N_13213,N_13342);
nor U13563 (N_13563,N_13370,N_13489);
nor U13564 (N_13564,N_13454,N_13466);
nor U13565 (N_13565,N_13498,N_13324);
xnor U13566 (N_13566,N_13302,N_13369);
and U13567 (N_13567,N_13347,N_13242);
xor U13568 (N_13568,N_13495,N_13453);
xnor U13569 (N_13569,N_13469,N_13294);
xor U13570 (N_13570,N_13349,N_13226);
xor U13571 (N_13571,N_13203,N_13374);
xor U13572 (N_13572,N_13479,N_13271);
and U13573 (N_13573,N_13436,N_13209);
nor U13574 (N_13574,N_13447,N_13262);
and U13575 (N_13575,N_13415,N_13332);
nand U13576 (N_13576,N_13383,N_13210);
nand U13577 (N_13577,N_13411,N_13220);
nor U13578 (N_13578,N_13400,N_13287);
nand U13579 (N_13579,N_13352,N_13399);
or U13580 (N_13580,N_13218,N_13482);
or U13581 (N_13581,N_13438,N_13270);
nand U13582 (N_13582,N_13476,N_13492);
xor U13583 (N_13583,N_13202,N_13455);
and U13584 (N_13584,N_13480,N_13336);
and U13585 (N_13585,N_13394,N_13300);
or U13586 (N_13586,N_13404,N_13483);
nor U13587 (N_13587,N_13200,N_13403);
and U13588 (N_13588,N_13356,N_13339);
nor U13589 (N_13589,N_13372,N_13308);
or U13590 (N_13590,N_13267,N_13278);
nand U13591 (N_13591,N_13325,N_13249);
and U13592 (N_13592,N_13223,N_13463);
nand U13593 (N_13593,N_13445,N_13206);
xnor U13594 (N_13594,N_13392,N_13478);
and U13595 (N_13595,N_13430,N_13232);
xor U13596 (N_13596,N_13261,N_13256);
and U13597 (N_13597,N_13244,N_13381);
and U13598 (N_13598,N_13243,N_13292);
or U13599 (N_13599,N_13353,N_13393);
or U13600 (N_13600,N_13254,N_13309);
nor U13601 (N_13601,N_13378,N_13380);
and U13602 (N_13602,N_13236,N_13420);
or U13603 (N_13603,N_13443,N_13396);
or U13604 (N_13604,N_13442,N_13408);
nand U13605 (N_13605,N_13488,N_13449);
nand U13606 (N_13606,N_13310,N_13251);
nand U13607 (N_13607,N_13424,N_13208);
nor U13608 (N_13608,N_13335,N_13461);
xor U13609 (N_13609,N_13422,N_13266);
and U13610 (N_13610,N_13435,N_13234);
or U13611 (N_13611,N_13306,N_13274);
nor U13612 (N_13612,N_13289,N_13487);
nor U13613 (N_13613,N_13410,N_13428);
or U13614 (N_13614,N_13215,N_13322);
or U13615 (N_13615,N_13311,N_13364);
and U13616 (N_13616,N_13272,N_13264);
nor U13617 (N_13617,N_13434,N_13247);
and U13618 (N_13618,N_13360,N_13228);
and U13619 (N_13619,N_13304,N_13245);
or U13620 (N_13620,N_13358,N_13421);
xnor U13621 (N_13621,N_13338,N_13390);
nor U13622 (N_13622,N_13217,N_13340);
nand U13623 (N_13623,N_13230,N_13382);
and U13624 (N_13624,N_13348,N_13465);
or U13625 (N_13625,N_13406,N_13204);
nand U13626 (N_13626,N_13288,N_13437);
and U13627 (N_13627,N_13229,N_13386);
nor U13628 (N_13628,N_13429,N_13285);
nand U13629 (N_13629,N_13366,N_13477);
nand U13630 (N_13630,N_13207,N_13321);
nor U13631 (N_13631,N_13326,N_13384);
nand U13632 (N_13632,N_13432,N_13252);
nor U13633 (N_13633,N_13409,N_13451);
nand U13634 (N_13634,N_13371,N_13277);
xnor U13635 (N_13635,N_13318,N_13319);
xnor U13636 (N_13636,N_13493,N_13497);
or U13637 (N_13637,N_13413,N_13313);
nand U13638 (N_13638,N_13433,N_13259);
nand U13639 (N_13639,N_13253,N_13216);
nor U13640 (N_13640,N_13316,N_13315);
xnor U13641 (N_13641,N_13414,N_13425);
xor U13642 (N_13642,N_13231,N_13265);
or U13643 (N_13643,N_13328,N_13205);
nand U13644 (N_13644,N_13255,N_13405);
xor U13645 (N_13645,N_13327,N_13323);
nor U13646 (N_13646,N_13401,N_13260);
nand U13647 (N_13647,N_13417,N_13426);
nor U13648 (N_13648,N_13494,N_13296);
and U13649 (N_13649,N_13301,N_13303);
or U13650 (N_13650,N_13473,N_13218);
nand U13651 (N_13651,N_13403,N_13373);
nor U13652 (N_13652,N_13220,N_13416);
nor U13653 (N_13653,N_13223,N_13210);
or U13654 (N_13654,N_13224,N_13267);
or U13655 (N_13655,N_13271,N_13435);
and U13656 (N_13656,N_13275,N_13239);
nor U13657 (N_13657,N_13437,N_13362);
xor U13658 (N_13658,N_13490,N_13381);
xnor U13659 (N_13659,N_13488,N_13494);
nand U13660 (N_13660,N_13398,N_13356);
xnor U13661 (N_13661,N_13336,N_13483);
and U13662 (N_13662,N_13319,N_13489);
xnor U13663 (N_13663,N_13291,N_13210);
xor U13664 (N_13664,N_13482,N_13311);
nor U13665 (N_13665,N_13307,N_13348);
or U13666 (N_13666,N_13249,N_13359);
and U13667 (N_13667,N_13348,N_13290);
nand U13668 (N_13668,N_13335,N_13318);
nand U13669 (N_13669,N_13409,N_13276);
xnor U13670 (N_13670,N_13440,N_13239);
xnor U13671 (N_13671,N_13491,N_13206);
xnor U13672 (N_13672,N_13225,N_13436);
or U13673 (N_13673,N_13312,N_13251);
nor U13674 (N_13674,N_13318,N_13431);
and U13675 (N_13675,N_13412,N_13376);
xnor U13676 (N_13676,N_13220,N_13232);
xor U13677 (N_13677,N_13419,N_13220);
nand U13678 (N_13678,N_13485,N_13279);
nand U13679 (N_13679,N_13492,N_13227);
or U13680 (N_13680,N_13282,N_13300);
and U13681 (N_13681,N_13476,N_13351);
xor U13682 (N_13682,N_13437,N_13450);
and U13683 (N_13683,N_13457,N_13281);
or U13684 (N_13684,N_13475,N_13492);
or U13685 (N_13685,N_13418,N_13442);
nand U13686 (N_13686,N_13390,N_13244);
nand U13687 (N_13687,N_13330,N_13401);
xor U13688 (N_13688,N_13305,N_13342);
xor U13689 (N_13689,N_13354,N_13287);
xor U13690 (N_13690,N_13437,N_13431);
or U13691 (N_13691,N_13296,N_13210);
or U13692 (N_13692,N_13478,N_13236);
nor U13693 (N_13693,N_13366,N_13368);
or U13694 (N_13694,N_13273,N_13240);
xnor U13695 (N_13695,N_13486,N_13291);
and U13696 (N_13696,N_13207,N_13388);
xor U13697 (N_13697,N_13241,N_13264);
or U13698 (N_13698,N_13257,N_13273);
and U13699 (N_13699,N_13395,N_13470);
or U13700 (N_13700,N_13451,N_13377);
or U13701 (N_13701,N_13295,N_13281);
nand U13702 (N_13702,N_13461,N_13397);
nand U13703 (N_13703,N_13318,N_13491);
and U13704 (N_13704,N_13377,N_13350);
nor U13705 (N_13705,N_13344,N_13293);
nor U13706 (N_13706,N_13451,N_13237);
and U13707 (N_13707,N_13358,N_13381);
nand U13708 (N_13708,N_13287,N_13281);
xor U13709 (N_13709,N_13356,N_13399);
nand U13710 (N_13710,N_13208,N_13446);
nand U13711 (N_13711,N_13419,N_13436);
and U13712 (N_13712,N_13448,N_13432);
xnor U13713 (N_13713,N_13267,N_13234);
nor U13714 (N_13714,N_13425,N_13255);
xor U13715 (N_13715,N_13268,N_13438);
and U13716 (N_13716,N_13273,N_13250);
nand U13717 (N_13717,N_13374,N_13406);
xor U13718 (N_13718,N_13227,N_13368);
nand U13719 (N_13719,N_13385,N_13335);
or U13720 (N_13720,N_13335,N_13281);
xor U13721 (N_13721,N_13348,N_13471);
nand U13722 (N_13722,N_13492,N_13344);
nor U13723 (N_13723,N_13205,N_13387);
xnor U13724 (N_13724,N_13216,N_13384);
and U13725 (N_13725,N_13410,N_13229);
nor U13726 (N_13726,N_13261,N_13385);
xor U13727 (N_13727,N_13275,N_13305);
and U13728 (N_13728,N_13417,N_13440);
nand U13729 (N_13729,N_13288,N_13330);
nand U13730 (N_13730,N_13365,N_13393);
and U13731 (N_13731,N_13408,N_13317);
nand U13732 (N_13732,N_13285,N_13463);
or U13733 (N_13733,N_13206,N_13457);
nor U13734 (N_13734,N_13323,N_13286);
and U13735 (N_13735,N_13391,N_13475);
and U13736 (N_13736,N_13432,N_13434);
nor U13737 (N_13737,N_13436,N_13456);
nand U13738 (N_13738,N_13460,N_13231);
and U13739 (N_13739,N_13226,N_13318);
nand U13740 (N_13740,N_13298,N_13437);
nand U13741 (N_13741,N_13232,N_13381);
and U13742 (N_13742,N_13255,N_13465);
xor U13743 (N_13743,N_13395,N_13411);
or U13744 (N_13744,N_13266,N_13353);
and U13745 (N_13745,N_13293,N_13361);
xnor U13746 (N_13746,N_13304,N_13368);
nand U13747 (N_13747,N_13354,N_13294);
nand U13748 (N_13748,N_13463,N_13429);
nand U13749 (N_13749,N_13450,N_13322);
nor U13750 (N_13750,N_13261,N_13423);
or U13751 (N_13751,N_13339,N_13351);
nand U13752 (N_13752,N_13435,N_13315);
or U13753 (N_13753,N_13276,N_13349);
and U13754 (N_13754,N_13428,N_13227);
nand U13755 (N_13755,N_13279,N_13460);
xor U13756 (N_13756,N_13217,N_13466);
nand U13757 (N_13757,N_13457,N_13373);
xor U13758 (N_13758,N_13422,N_13375);
nand U13759 (N_13759,N_13411,N_13297);
nand U13760 (N_13760,N_13443,N_13411);
nand U13761 (N_13761,N_13470,N_13365);
and U13762 (N_13762,N_13452,N_13484);
nand U13763 (N_13763,N_13392,N_13296);
xor U13764 (N_13764,N_13474,N_13450);
or U13765 (N_13765,N_13438,N_13461);
xnor U13766 (N_13766,N_13330,N_13305);
nand U13767 (N_13767,N_13268,N_13402);
xnor U13768 (N_13768,N_13260,N_13482);
or U13769 (N_13769,N_13227,N_13202);
and U13770 (N_13770,N_13235,N_13249);
or U13771 (N_13771,N_13436,N_13484);
nor U13772 (N_13772,N_13317,N_13451);
xnor U13773 (N_13773,N_13343,N_13245);
nor U13774 (N_13774,N_13402,N_13399);
nor U13775 (N_13775,N_13300,N_13376);
xor U13776 (N_13776,N_13272,N_13355);
and U13777 (N_13777,N_13244,N_13281);
nor U13778 (N_13778,N_13271,N_13233);
nand U13779 (N_13779,N_13427,N_13457);
and U13780 (N_13780,N_13420,N_13257);
nor U13781 (N_13781,N_13398,N_13337);
or U13782 (N_13782,N_13331,N_13345);
xnor U13783 (N_13783,N_13397,N_13272);
xor U13784 (N_13784,N_13217,N_13313);
nand U13785 (N_13785,N_13450,N_13251);
xnor U13786 (N_13786,N_13306,N_13200);
nor U13787 (N_13787,N_13477,N_13223);
nand U13788 (N_13788,N_13293,N_13421);
nand U13789 (N_13789,N_13325,N_13220);
and U13790 (N_13790,N_13399,N_13218);
nor U13791 (N_13791,N_13465,N_13267);
xor U13792 (N_13792,N_13308,N_13234);
nand U13793 (N_13793,N_13262,N_13409);
and U13794 (N_13794,N_13213,N_13242);
nor U13795 (N_13795,N_13456,N_13358);
nand U13796 (N_13796,N_13400,N_13215);
nor U13797 (N_13797,N_13297,N_13440);
and U13798 (N_13798,N_13290,N_13346);
nand U13799 (N_13799,N_13463,N_13322);
or U13800 (N_13800,N_13571,N_13723);
xnor U13801 (N_13801,N_13554,N_13549);
nand U13802 (N_13802,N_13582,N_13716);
and U13803 (N_13803,N_13614,N_13730);
xor U13804 (N_13804,N_13641,N_13751);
nand U13805 (N_13805,N_13649,N_13588);
xnor U13806 (N_13806,N_13532,N_13510);
or U13807 (N_13807,N_13720,N_13598);
xor U13808 (N_13808,N_13572,N_13706);
and U13809 (N_13809,N_13519,N_13735);
nand U13810 (N_13810,N_13547,N_13692);
or U13811 (N_13811,N_13652,N_13548);
nand U13812 (N_13812,N_13546,N_13690);
and U13813 (N_13813,N_13701,N_13782);
xnor U13814 (N_13814,N_13615,N_13711);
nand U13815 (N_13815,N_13752,N_13778);
nand U13816 (N_13816,N_13528,N_13784);
xor U13817 (N_13817,N_13775,N_13655);
xor U13818 (N_13818,N_13671,N_13677);
nor U13819 (N_13819,N_13639,N_13623);
or U13820 (N_13820,N_13658,N_13590);
or U13821 (N_13821,N_13539,N_13665);
xor U13822 (N_13822,N_13733,N_13724);
nor U13823 (N_13823,N_13798,N_13699);
and U13824 (N_13824,N_13789,N_13584);
nor U13825 (N_13825,N_13587,N_13766);
xor U13826 (N_13826,N_13607,N_13651);
or U13827 (N_13827,N_13553,N_13796);
and U13828 (N_13828,N_13764,N_13648);
nand U13829 (N_13829,N_13786,N_13559);
and U13830 (N_13830,N_13631,N_13626);
nor U13831 (N_13831,N_13656,N_13776);
and U13832 (N_13832,N_13713,N_13630);
xnor U13833 (N_13833,N_13797,N_13540);
xnor U13834 (N_13834,N_13715,N_13684);
xor U13835 (N_13835,N_13524,N_13592);
and U13836 (N_13836,N_13543,N_13505);
xnor U13837 (N_13837,N_13659,N_13676);
xnor U13838 (N_13838,N_13742,N_13602);
xor U13839 (N_13839,N_13507,N_13581);
nand U13840 (N_13840,N_13618,N_13537);
xnor U13841 (N_13841,N_13691,N_13674);
and U13842 (N_13842,N_13653,N_13600);
and U13843 (N_13843,N_13515,N_13617);
nand U13844 (N_13844,N_13749,N_13650);
and U13845 (N_13845,N_13792,N_13574);
and U13846 (N_13846,N_13688,N_13667);
xor U13847 (N_13847,N_13771,N_13710);
nand U13848 (N_13848,N_13603,N_13601);
or U13849 (N_13849,N_13534,N_13702);
xor U13850 (N_13850,N_13568,N_13663);
nand U13851 (N_13851,N_13561,N_13682);
xor U13852 (N_13852,N_13799,N_13616);
nand U13853 (N_13853,N_13596,N_13608);
xnor U13854 (N_13854,N_13683,N_13576);
or U13855 (N_13855,N_13636,N_13502);
nor U13856 (N_13856,N_13625,N_13647);
or U13857 (N_13857,N_13783,N_13753);
and U13858 (N_13858,N_13604,N_13737);
nor U13859 (N_13859,N_13687,N_13666);
or U13860 (N_13860,N_13660,N_13695);
nand U13861 (N_13861,N_13627,N_13506);
and U13862 (N_13862,N_13762,N_13787);
or U13863 (N_13863,N_13678,N_13550);
or U13864 (N_13864,N_13536,N_13545);
nor U13865 (N_13865,N_13769,N_13746);
nand U13866 (N_13866,N_13514,N_13564);
nor U13867 (N_13867,N_13760,N_13673);
xnor U13868 (N_13868,N_13741,N_13714);
xor U13869 (N_13869,N_13694,N_13542);
nor U13870 (N_13870,N_13612,N_13721);
nand U13871 (N_13871,N_13747,N_13529);
or U13872 (N_13872,N_13662,N_13644);
nor U13873 (N_13873,N_13794,N_13585);
nor U13874 (N_13874,N_13521,N_13516);
xnor U13875 (N_13875,N_13734,N_13689);
xor U13876 (N_13876,N_13624,N_13698);
nand U13877 (N_13877,N_13593,N_13704);
or U13878 (N_13878,N_13664,N_13573);
or U13879 (N_13879,N_13729,N_13731);
xor U13880 (N_13880,N_13793,N_13565);
nor U13881 (N_13881,N_13556,N_13541);
nor U13882 (N_13882,N_13504,N_13781);
nand U13883 (N_13883,N_13591,N_13709);
xnor U13884 (N_13884,N_13520,N_13773);
nor U13885 (N_13885,N_13622,N_13739);
nand U13886 (N_13886,N_13597,N_13705);
xnor U13887 (N_13887,N_13745,N_13579);
nand U13888 (N_13888,N_13566,N_13754);
xnor U13889 (N_13889,N_13759,N_13500);
nor U13890 (N_13890,N_13523,N_13661);
nor U13891 (N_13891,N_13578,N_13642);
nand U13892 (N_13892,N_13621,N_13580);
xor U13893 (N_13893,N_13633,N_13672);
xor U13894 (N_13894,N_13606,N_13791);
nand U13895 (N_13895,N_13567,N_13785);
and U13896 (N_13896,N_13562,N_13669);
or U13897 (N_13897,N_13725,N_13728);
xnor U13898 (N_13898,N_13743,N_13646);
nand U13899 (N_13899,N_13605,N_13717);
or U13900 (N_13900,N_13708,N_13732);
nand U13901 (N_13901,N_13635,N_13531);
xnor U13902 (N_13902,N_13718,N_13513);
xor U13903 (N_13903,N_13670,N_13517);
nor U13904 (N_13904,N_13779,N_13696);
or U13905 (N_13905,N_13558,N_13533);
nand U13906 (N_13906,N_13544,N_13595);
nor U13907 (N_13907,N_13628,N_13763);
or U13908 (N_13908,N_13589,N_13509);
or U13909 (N_13909,N_13693,N_13570);
xor U13910 (N_13910,N_13599,N_13563);
nand U13911 (N_13911,N_13557,N_13609);
or U13912 (N_13912,N_13638,N_13680);
or U13913 (N_13913,N_13795,N_13535);
or U13914 (N_13914,N_13640,N_13632);
or U13915 (N_13915,N_13765,N_13757);
and U13916 (N_13916,N_13575,N_13569);
nand U13917 (N_13917,N_13501,N_13768);
nand U13918 (N_13918,N_13707,N_13620);
xnor U13919 (N_13919,N_13512,N_13619);
and U13920 (N_13920,N_13790,N_13645);
or U13921 (N_13921,N_13522,N_13643);
and U13922 (N_13922,N_13726,N_13700);
nand U13923 (N_13923,N_13770,N_13703);
xnor U13924 (N_13924,N_13518,N_13610);
and U13925 (N_13925,N_13679,N_13748);
nor U13926 (N_13926,N_13552,N_13634);
nor U13927 (N_13927,N_13777,N_13750);
and U13928 (N_13928,N_13611,N_13551);
xnor U13929 (N_13929,N_13685,N_13740);
and U13930 (N_13930,N_13668,N_13527);
nand U13931 (N_13931,N_13755,N_13738);
nand U13932 (N_13932,N_13526,N_13613);
nand U13933 (N_13933,N_13511,N_13657);
nand U13934 (N_13934,N_13560,N_13712);
or U13935 (N_13935,N_13530,N_13780);
nand U13936 (N_13936,N_13772,N_13727);
xnor U13937 (N_13937,N_13555,N_13788);
nor U13938 (N_13938,N_13761,N_13681);
xnor U13939 (N_13939,N_13583,N_13719);
nor U13940 (N_13940,N_13722,N_13577);
xor U13941 (N_13941,N_13686,N_13697);
or U13942 (N_13942,N_13525,N_13756);
nand U13943 (N_13943,N_13637,N_13503);
and U13944 (N_13944,N_13629,N_13675);
or U13945 (N_13945,N_13767,N_13774);
xnor U13946 (N_13946,N_13654,N_13736);
and U13947 (N_13947,N_13744,N_13758);
or U13948 (N_13948,N_13586,N_13594);
nor U13949 (N_13949,N_13538,N_13508);
or U13950 (N_13950,N_13657,N_13754);
nand U13951 (N_13951,N_13749,N_13610);
xor U13952 (N_13952,N_13573,N_13781);
nor U13953 (N_13953,N_13589,N_13659);
or U13954 (N_13954,N_13723,N_13586);
and U13955 (N_13955,N_13589,N_13625);
or U13956 (N_13956,N_13517,N_13609);
nand U13957 (N_13957,N_13579,N_13570);
and U13958 (N_13958,N_13706,N_13655);
and U13959 (N_13959,N_13584,N_13620);
and U13960 (N_13960,N_13637,N_13738);
nand U13961 (N_13961,N_13622,N_13751);
or U13962 (N_13962,N_13516,N_13605);
and U13963 (N_13963,N_13601,N_13753);
and U13964 (N_13964,N_13508,N_13767);
and U13965 (N_13965,N_13702,N_13605);
nor U13966 (N_13966,N_13538,N_13671);
and U13967 (N_13967,N_13632,N_13659);
and U13968 (N_13968,N_13612,N_13506);
nor U13969 (N_13969,N_13734,N_13707);
nand U13970 (N_13970,N_13545,N_13505);
and U13971 (N_13971,N_13556,N_13522);
nand U13972 (N_13972,N_13677,N_13576);
or U13973 (N_13973,N_13741,N_13544);
xor U13974 (N_13974,N_13734,N_13744);
nor U13975 (N_13975,N_13779,N_13728);
xnor U13976 (N_13976,N_13640,N_13567);
xnor U13977 (N_13977,N_13639,N_13687);
nand U13978 (N_13978,N_13690,N_13795);
and U13979 (N_13979,N_13738,N_13556);
nand U13980 (N_13980,N_13538,N_13501);
or U13981 (N_13981,N_13628,N_13501);
or U13982 (N_13982,N_13640,N_13558);
nor U13983 (N_13983,N_13537,N_13611);
nand U13984 (N_13984,N_13514,N_13533);
nor U13985 (N_13985,N_13731,N_13672);
or U13986 (N_13986,N_13723,N_13715);
nor U13987 (N_13987,N_13663,N_13646);
or U13988 (N_13988,N_13754,N_13562);
or U13989 (N_13989,N_13519,N_13609);
and U13990 (N_13990,N_13722,N_13758);
nor U13991 (N_13991,N_13640,N_13786);
nand U13992 (N_13992,N_13588,N_13560);
nor U13993 (N_13993,N_13551,N_13747);
or U13994 (N_13994,N_13503,N_13734);
xnor U13995 (N_13995,N_13589,N_13684);
nand U13996 (N_13996,N_13620,N_13647);
and U13997 (N_13997,N_13517,N_13692);
nand U13998 (N_13998,N_13690,N_13646);
nand U13999 (N_13999,N_13744,N_13757);
or U14000 (N_14000,N_13658,N_13750);
nand U14001 (N_14001,N_13502,N_13567);
nor U14002 (N_14002,N_13770,N_13529);
nand U14003 (N_14003,N_13658,N_13760);
or U14004 (N_14004,N_13699,N_13779);
or U14005 (N_14005,N_13682,N_13628);
or U14006 (N_14006,N_13741,N_13633);
and U14007 (N_14007,N_13733,N_13532);
or U14008 (N_14008,N_13537,N_13743);
and U14009 (N_14009,N_13696,N_13543);
xor U14010 (N_14010,N_13798,N_13504);
nor U14011 (N_14011,N_13600,N_13549);
nand U14012 (N_14012,N_13653,N_13648);
and U14013 (N_14013,N_13610,N_13672);
nor U14014 (N_14014,N_13613,N_13689);
xnor U14015 (N_14015,N_13696,N_13770);
or U14016 (N_14016,N_13659,N_13665);
nor U14017 (N_14017,N_13598,N_13567);
and U14018 (N_14018,N_13797,N_13732);
or U14019 (N_14019,N_13784,N_13739);
xor U14020 (N_14020,N_13680,N_13573);
nor U14021 (N_14021,N_13784,N_13771);
or U14022 (N_14022,N_13519,N_13580);
and U14023 (N_14023,N_13613,N_13582);
nand U14024 (N_14024,N_13579,N_13709);
and U14025 (N_14025,N_13641,N_13740);
and U14026 (N_14026,N_13597,N_13620);
or U14027 (N_14027,N_13698,N_13714);
or U14028 (N_14028,N_13576,N_13648);
nor U14029 (N_14029,N_13771,N_13599);
or U14030 (N_14030,N_13770,N_13730);
or U14031 (N_14031,N_13639,N_13706);
nor U14032 (N_14032,N_13503,N_13526);
xnor U14033 (N_14033,N_13787,N_13761);
nand U14034 (N_14034,N_13698,N_13769);
xor U14035 (N_14035,N_13617,N_13598);
xnor U14036 (N_14036,N_13526,N_13523);
or U14037 (N_14037,N_13633,N_13549);
xnor U14038 (N_14038,N_13726,N_13500);
nand U14039 (N_14039,N_13572,N_13527);
xor U14040 (N_14040,N_13766,N_13576);
or U14041 (N_14041,N_13517,N_13570);
or U14042 (N_14042,N_13793,N_13575);
xnor U14043 (N_14043,N_13743,N_13673);
nor U14044 (N_14044,N_13554,N_13656);
nor U14045 (N_14045,N_13697,N_13500);
and U14046 (N_14046,N_13717,N_13675);
or U14047 (N_14047,N_13651,N_13505);
xor U14048 (N_14048,N_13753,N_13618);
or U14049 (N_14049,N_13570,N_13681);
or U14050 (N_14050,N_13503,N_13731);
nand U14051 (N_14051,N_13658,N_13783);
or U14052 (N_14052,N_13729,N_13630);
nand U14053 (N_14053,N_13572,N_13708);
or U14054 (N_14054,N_13539,N_13561);
nor U14055 (N_14055,N_13691,N_13727);
and U14056 (N_14056,N_13544,N_13547);
xor U14057 (N_14057,N_13686,N_13791);
and U14058 (N_14058,N_13696,N_13784);
nand U14059 (N_14059,N_13724,N_13537);
and U14060 (N_14060,N_13754,N_13654);
and U14061 (N_14061,N_13712,N_13555);
xor U14062 (N_14062,N_13766,N_13765);
xor U14063 (N_14063,N_13789,N_13591);
or U14064 (N_14064,N_13779,N_13759);
xnor U14065 (N_14065,N_13600,N_13552);
xor U14066 (N_14066,N_13743,N_13667);
nand U14067 (N_14067,N_13571,N_13766);
nand U14068 (N_14068,N_13567,N_13778);
and U14069 (N_14069,N_13685,N_13512);
and U14070 (N_14070,N_13512,N_13744);
and U14071 (N_14071,N_13779,N_13744);
xor U14072 (N_14072,N_13724,N_13752);
xnor U14073 (N_14073,N_13780,N_13646);
or U14074 (N_14074,N_13587,N_13727);
xnor U14075 (N_14075,N_13563,N_13507);
xnor U14076 (N_14076,N_13607,N_13748);
nand U14077 (N_14077,N_13523,N_13783);
nor U14078 (N_14078,N_13717,N_13577);
and U14079 (N_14079,N_13594,N_13536);
or U14080 (N_14080,N_13778,N_13507);
xor U14081 (N_14081,N_13739,N_13643);
and U14082 (N_14082,N_13659,N_13720);
nor U14083 (N_14083,N_13562,N_13690);
xor U14084 (N_14084,N_13742,N_13767);
xnor U14085 (N_14085,N_13798,N_13676);
xnor U14086 (N_14086,N_13651,N_13754);
xnor U14087 (N_14087,N_13689,N_13770);
xnor U14088 (N_14088,N_13687,N_13563);
nor U14089 (N_14089,N_13703,N_13608);
xnor U14090 (N_14090,N_13690,N_13745);
nand U14091 (N_14091,N_13684,N_13506);
nand U14092 (N_14092,N_13569,N_13548);
or U14093 (N_14093,N_13655,N_13599);
nor U14094 (N_14094,N_13681,N_13638);
nand U14095 (N_14095,N_13638,N_13736);
or U14096 (N_14096,N_13725,N_13533);
nor U14097 (N_14097,N_13564,N_13645);
nand U14098 (N_14098,N_13785,N_13715);
or U14099 (N_14099,N_13706,N_13690);
nand U14100 (N_14100,N_13979,N_13815);
nor U14101 (N_14101,N_13993,N_13983);
xor U14102 (N_14102,N_14054,N_13931);
xnor U14103 (N_14103,N_14026,N_14052);
nand U14104 (N_14104,N_13975,N_14085);
and U14105 (N_14105,N_14075,N_14080);
nand U14106 (N_14106,N_13988,N_14014);
xnor U14107 (N_14107,N_13887,N_13811);
nor U14108 (N_14108,N_13879,N_14017);
nor U14109 (N_14109,N_13850,N_13928);
xnor U14110 (N_14110,N_14003,N_13892);
and U14111 (N_14111,N_13904,N_13933);
nand U14112 (N_14112,N_14057,N_13981);
xor U14113 (N_14113,N_13828,N_13967);
nor U14114 (N_14114,N_13941,N_14048);
nand U14115 (N_14115,N_13821,N_13958);
nor U14116 (N_14116,N_13814,N_13833);
xnor U14117 (N_14117,N_13955,N_13872);
nand U14118 (N_14118,N_13880,N_13991);
nor U14119 (N_14119,N_13905,N_13940);
and U14120 (N_14120,N_13855,N_14068);
and U14121 (N_14121,N_13959,N_13971);
or U14122 (N_14122,N_13921,N_14030);
or U14123 (N_14123,N_13974,N_14033);
xor U14124 (N_14124,N_14099,N_13961);
or U14125 (N_14125,N_13894,N_13836);
and U14126 (N_14126,N_14020,N_13868);
nor U14127 (N_14127,N_13900,N_14044);
or U14128 (N_14128,N_14065,N_14060);
or U14129 (N_14129,N_13823,N_14095);
and U14130 (N_14130,N_14046,N_13875);
xnor U14131 (N_14131,N_14083,N_13890);
and U14132 (N_14132,N_14073,N_13934);
nand U14133 (N_14133,N_13897,N_14088);
xor U14134 (N_14134,N_14031,N_14045);
nand U14135 (N_14135,N_13857,N_13997);
and U14136 (N_14136,N_13965,N_13893);
nand U14137 (N_14137,N_13952,N_13942);
and U14138 (N_14138,N_13970,N_13852);
nand U14139 (N_14139,N_14038,N_13990);
nand U14140 (N_14140,N_14097,N_13946);
nor U14141 (N_14141,N_14079,N_14091);
and U14142 (N_14142,N_13834,N_13989);
or U14143 (N_14143,N_13994,N_14004);
and U14144 (N_14144,N_13935,N_14084);
nand U14145 (N_14145,N_13812,N_13816);
nor U14146 (N_14146,N_13925,N_13851);
and U14147 (N_14147,N_14037,N_14087);
and U14148 (N_14148,N_13891,N_13831);
and U14149 (N_14149,N_13884,N_13976);
nand U14150 (N_14150,N_13865,N_14072);
xnor U14151 (N_14151,N_14090,N_13911);
nand U14152 (N_14152,N_13984,N_14047);
xnor U14153 (N_14153,N_13835,N_14002);
nand U14154 (N_14154,N_13829,N_13949);
or U14155 (N_14155,N_14076,N_13881);
nand U14156 (N_14156,N_13899,N_13830);
nor U14157 (N_14157,N_14066,N_13930);
nor U14158 (N_14158,N_13846,N_13945);
nand U14159 (N_14159,N_13929,N_13987);
and U14160 (N_14160,N_14092,N_13827);
and U14161 (N_14161,N_13882,N_13943);
nor U14162 (N_14162,N_13863,N_13803);
and U14163 (N_14163,N_13801,N_13832);
nand U14164 (N_14164,N_13840,N_14025);
or U14165 (N_14165,N_14067,N_13849);
nand U14166 (N_14166,N_14059,N_13913);
or U14167 (N_14167,N_13922,N_13927);
xnor U14168 (N_14168,N_13847,N_13874);
and U14169 (N_14169,N_14019,N_13844);
or U14170 (N_14170,N_13826,N_13985);
or U14171 (N_14171,N_13895,N_14013);
and U14172 (N_14172,N_14018,N_13995);
nor U14173 (N_14173,N_14042,N_13907);
nor U14174 (N_14174,N_13999,N_13972);
xor U14175 (N_14175,N_14086,N_13838);
and U14176 (N_14176,N_14000,N_14011);
and U14177 (N_14177,N_13918,N_13822);
and U14178 (N_14178,N_13982,N_13804);
or U14179 (N_14179,N_13819,N_13937);
nor U14180 (N_14180,N_14070,N_14034);
nor U14181 (N_14181,N_13861,N_13869);
nand U14182 (N_14182,N_13966,N_14028);
or U14183 (N_14183,N_14082,N_14043);
xor U14184 (N_14184,N_13859,N_13909);
xor U14185 (N_14185,N_14027,N_13992);
or U14186 (N_14186,N_14077,N_13953);
nor U14187 (N_14187,N_14098,N_13998);
or U14188 (N_14188,N_13964,N_14015);
or U14189 (N_14189,N_14062,N_14016);
or U14190 (N_14190,N_14012,N_13843);
and U14191 (N_14191,N_13877,N_13839);
nand U14192 (N_14192,N_13820,N_13978);
xnor U14193 (N_14193,N_13951,N_13807);
xnor U14194 (N_14194,N_13977,N_14022);
xnor U14195 (N_14195,N_14071,N_13932);
nor U14196 (N_14196,N_13876,N_13948);
xnor U14197 (N_14197,N_13906,N_13968);
xnor U14198 (N_14198,N_14049,N_14006);
or U14199 (N_14199,N_13885,N_13825);
and U14200 (N_14200,N_14089,N_13915);
or U14201 (N_14201,N_14055,N_13969);
or U14202 (N_14202,N_14035,N_13947);
nor U14203 (N_14203,N_13806,N_14061);
or U14204 (N_14204,N_13800,N_14007);
and U14205 (N_14205,N_14001,N_14064);
and U14206 (N_14206,N_13908,N_13853);
and U14207 (N_14207,N_13954,N_13886);
nand U14208 (N_14208,N_13986,N_13817);
or U14209 (N_14209,N_14078,N_13802);
xnor U14210 (N_14210,N_14008,N_13837);
nor U14211 (N_14211,N_13856,N_13870);
nand U14212 (N_14212,N_14093,N_13873);
or U14213 (N_14213,N_13923,N_14032);
and U14214 (N_14214,N_13938,N_14029);
and U14215 (N_14215,N_14094,N_13962);
xnor U14216 (N_14216,N_13960,N_13898);
nor U14217 (N_14217,N_13862,N_14053);
xnor U14218 (N_14218,N_13996,N_13864);
or U14219 (N_14219,N_13824,N_13957);
and U14220 (N_14220,N_13936,N_13896);
and U14221 (N_14221,N_13919,N_13866);
nand U14222 (N_14222,N_13858,N_13883);
nand U14223 (N_14223,N_13808,N_13926);
and U14224 (N_14224,N_14039,N_13889);
nor U14225 (N_14225,N_14021,N_14056);
nor U14226 (N_14226,N_13805,N_14024);
nor U14227 (N_14227,N_14051,N_13888);
or U14228 (N_14228,N_13867,N_13980);
xnor U14229 (N_14229,N_13818,N_13912);
nand U14230 (N_14230,N_14074,N_13810);
nor U14231 (N_14231,N_14009,N_13914);
and U14232 (N_14232,N_13956,N_14041);
xor U14233 (N_14233,N_13901,N_13973);
xor U14234 (N_14234,N_14050,N_13924);
and U14235 (N_14235,N_13920,N_13917);
nor U14236 (N_14236,N_14096,N_14058);
or U14237 (N_14237,N_13813,N_13939);
and U14238 (N_14238,N_13860,N_13854);
or U14239 (N_14239,N_14023,N_14069);
or U14240 (N_14240,N_14081,N_13845);
and U14241 (N_14241,N_14005,N_13910);
xnor U14242 (N_14242,N_13903,N_14036);
and U14243 (N_14243,N_13809,N_13842);
nor U14244 (N_14244,N_13871,N_13944);
xor U14245 (N_14245,N_13902,N_14010);
nand U14246 (N_14246,N_13878,N_14040);
and U14247 (N_14247,N_13916,N_13950);
and U14248 (N_14248,N_13963,N_14063);
and U14249 (N_14249,N_13848,N_13841);
and U14250 (N_14250,N_14020,N_13885);
nor U14251 (N_14251,N_14099,N_13817);
nand U14252 (N_14252,N_14042,N_14057);
nand U14253 (N_14253,N_14092,N_14067);
nand U14254 (N_14254,N_13806,N_14052);
and U14255 (N_14255,N_13975,N_14031);
nor U14256 (N_14256,N_13830,N_14070);
xnor U14257 (N_14257,N_13982,N_13860);
nand U14258 (N_14258,N_13972,N_13941);
and U14259 (N_14259,N_14057,N_13869);
xor U14260 (N_14260,N_14025,N_14010);
nor U14261 (N_14261,N_14029,N_13837);
nand U14262 (N_14262,N_13801,N_13999);
nor U14263 (N_14263,N_13823,N_13987);
nand U14264 (N_14264,N_13968,N_14052);
nor U14265 (N_14265,N_13831,N_14076);
and U14266 (N_14266,N_13923,N_13801);
nand U14267 (N_14267,N_13934,N_13953);
nand U14268 (N_14268,N_13870,N_13841);
and U14269 (N_14269,N_13978,N_13805);
and U14270 (N_14270,N_14062,N_13876);
xor U14271 (N_14271,N_13889,N_13905);
nand U14272 (N_14272,N_13820,N_13836);
and U14273 (N_14273,N_13948,N_13857);
or U14274 (N_14274,N_13972,N_13956);
and U14275 (N_14275,N_13934,N_14006);
or U14276 (N_14276,N_13806,N_13842);
xnor U14277 (N_14277,N_13944,N_13978);
nor U14278 (N_14278,N_13955,N_14047);
or U14279 (N_14279,N_13899,N_13837);
nor U14280 (N_14280,N_13839,N_13980);
xor U14281 (N_14281,N_14009,N_13994);
nand U14282 (N_14282,N_13940,N_13960);
xnor U14283 (N_14283,N_13903,N_13879);
nor U14284 (N_14284,N_13997,N_14082);
nor U14285 (N_14285,N_14065,N_13872);
or U14286 (N_14286,N_13995,N_13850);
nand U14287 (N_14287,N_14033,N_13877);
xnor U14288 (N_14288,N_13859,N_13860);
and U14289 (N_14289,N_14070,N_14012);
or U14290 (N_14290,N_13833,N_14078);
or U14291 (N_14291,N_13978,N_13910);
xor U14292 (N_14292,N_13916,N_14044);
and U14293 (N_14293,N_13821,N_14058);
nor U14294 (N_14294,N_14004,N_13935);
and U14295 (N_14295,N_14090,N_13826);
or U14296 (N_14296,N_13989,N_14062);
or U14297 (N_14297,N_13883,N_13907);
or U14298 (N_14298,N_14091,N_14037);
nor U14299 (N_14299,N_14005,N_13902);
nand U14300 (N_14300,N_14033,N_14067);
xnor U14301 (N_14301,N_13985,N_13862);
nand U14302 (N_14302,N_13877,N_13952);
nor U14303 (N_14303,N_14060,N_13818);
and U14304 (N_14304,N_13834,N_13820);
or U14305 (N_14305,N_13861,N_13939);
or U14306 (N_14306,N_13804,N_13892);
or U14307 (N_14307,N_13893,N_13863);
nand U14308 (N_14308,N_13905,N_13845);
and U14309 (N_14309,N_13826,N_13897);
nand U14310 (N_14310,N_13839,N_14021);
xnor U14311 (N_14311,N_13958,N_14045);
xnor U14312 (N_14312,N_13895,N_13965);
nor U14313 (N_14313,N_13885,N_14011);
nand U14314 (N_14314,N_13944,N_14050);
nor U14315 (N_14315,N_13961,N_14047);
or U14316 (N_14316,N_14089,N_13940);
or U14317 (N_14317,N_14092,N_13912);
xor U14318 (N_14318,N_13982,N_13846);
or U14319 (N_14319,N_13939,N_13988);
or U14320 (N_14320,N_13874,N_13972);
nand U14321 (N_14321,N_14085,N_14029);
nand U14322 (N_14322,N_13965,N_13806);
nor U14323 (N_14323,N_13891,N_13858);
xnor U14324 (N_14324,N_13937,N_13922);
nor U14325 (N_14325,N_13846,N_13889);
and U14326 (N_14326,N_14058,N_13886);
and U14327 (N_14327,N_14097,N_13937);
and U14328 (N_14328,N_13997,N_14093);
nand U14329 (N_14329,N_13964,N_13883);
and U14330 (N_14330,N_13879,N_13898);
nor U14331 (N_14331,N_13973,N_13985);
nor U14332 (N_14332,N_13895,N_14050);
xnor U14333 (N_14333,N_13865,N_13896);
xor U14334 (N_14334,N_13924,N_13974);
nand U14335 (N_14335,N_13906,N_14080);
nand U14336 (N_14336,N_13894,N_14050);
and U14337 (N_14337,N_13819,N_13811);
xor U14338 (N_14338,N_14088,N_14028);
or U14339 (N_14339,N_13965,N_14059);
and U14340 (N_14340,N_13827,N_13802);
nand U14341 (N_14341,N_13976,N_13932);
nor U14342 (N_14342,N_13856,N_13951);
and U14343 (N_14343,N_14004,N_14077);
nand U14344 (N_14344,N_13863,N_13946);
nor U14345 (N_14345,N_14037,N_13863);
or U14346 (N_14346,N_13891,N_14078);
and U14347 (N_14347,N_14010,N_13951);
nor U14348 (N_14348,N_13894,N_13964);
xor U14349 (N_14349,N_14027,N_14081);
xnor U14350 (N_14350,N_14035,N_13954);
nor U14351 (N_14351,N_14023,N_14029);
nor U14352 (N_14352,N_13902,N_14097);
or U14353 (N_14353,N_14052,N_13951);
nand U14354 (N_14354,N_13822,N_14006);
xnor U14355 (N_14355,N_14088,N_13848);
or U14356 (N_14356,N_13951,N_13957);
nand U14357 (N_14357,N_13901,N_13847);
and U14358 (N_14358,N_13938,N_14091);
nand U14359 (N_14359,N_13971,N_13938);
xnor U14360 (N_14360,N_14018,N_13865);
nor U14361 (N_14361,N_13949,N_14089);
nand U14362 (N_14362,N_14098,N_13812);
nand U14363 (N_14363,N_13985,N_14087);
nor U14364 (N_14364,N_13950,N_14038);
nor U14365 (N_14365,N_14037,N_14076);
nand U14366 (N_14366,N_13802,N_13899);
nor U14367 (N_14367,N_13836,N_13851);
or U14368 (N_14368,N_13882,N_14099);
nand U14369 (N_14369,N_14055,N_13982);
or U14370 (N_14370,N_14015,N_13960);
nor U14371 (N_14371,N_14019,N_13981);
and U14372 (N_14372,N_14004,N_13947);
or U14373 (N_14373,N_13826,N_14095);
xnor U14374 (N_14374,N_14096,N_13995);
nor U14375 (N_14375,N_13853,N_13817);
and U14376 (N_14376,N_13923,N_13835);
xor U14377 (N_14377,N_14076,N_13816);
or U14378 (N_14378,N_14029,N_13932);
xor U14379 (N_14379,N_13851,N_13835);
nor U14380 (N_14380,N_13819,N_14021);
or U14381 (N_14381,N_13869,N_13945);
nand U14382 (N_14382,N_13972,N_14058);
nor U14383 (N_14383,N_13888,N_14008);
or U14384 (N_14384,N_13880,N_13914);
nor U14385 (N_14385,N_14094,N_14093);
xor U14386 (N_14386,N_13932,N_13882);
and U14387 (N_14387,N_13999,N_13930);
or U14388 (N_14388,N_14015,N_13820);
and U14389 (N_14389,N_13810,N_14046);
nor U14390 (N_14390,N_14004,N_13992);
or U14391 (N_14391,N_14089,N_14000);
or U14392 (N_14392,N_13976,N_13996);
or U14393 (N_14393,N_14055,N_13924);
and U14394 (N_14394,N_13930,N_13802);
and U14395 (N_14395,N_14021,N_13918);
or U14396 (N_14396,N_14001,N_14022);
nand U14397 (N_14397,N_13985,N_14042);
or U14398 (N_14398,N_14078,N_13996);
nor U14399 (N_14399,N_13878,N_13902);
nand U14400 (N_14400,N_14366,N_14273);
nor U14401 (N_14401,N_14337,N_14259);
nor U14402 (N_14402,N_14324,N_14205);
and U14403 (N_14403,N_14393,N_14142);
nor U14404 (N_14404,N_14113,N_14147);
xor U14405 (N_14405,N_14262,N_14208);
nor U14406 (N_14406,N_14159,N_14327);
and U14407 (N_14407,N_14196,N_14272);
nor U14408 (N_14408,N_14108,N_14370);
nor U14409 (N_14409,N_14115,N_14240);
or U14410 (N_14410,N_14198,N_14357);
nor U14411 (N_14411,N_14136,N_14172);
nand U14412 (N_14412,N_14368,N_14251);
or U14413 (N_14413,N_14342,N_14120);
xnor U14414 (N_14414,N_14322,N_14333);
nand U14415 (N_14415,N_14275,N_14107);
nor U14416 (N_14416,N_14177,N_14310);
or U14417 (N_14417,N_14396,N_14188);
or U14418 (N_14418,N_14277,N_14160);
or U14419 (N_14419,N_14307,N_14350);
nand U14420 (N_14420,N_14346,N_14227);
nor U14421 (N_14421,N_14216,N_14110);
or U14422 (N_14422,N_14320,N_14166);
xnor U14423 (N_14423,N_14398,N_14138);
xnor U14424 (N_14424,N_14224,N_14131);
and U14425 (N_14425,N_14291,N_14135);
xor U14426 (N_14426,N_14339,N_14362);
nand U14427 (N_14427,N_14344,N_14399);
xnor U14428 (N_14428,N_14265,N_14116);
and U14429 (N_14429,N_14164,N_14330);
and U14430 (N_14430,N_14132,N_14246);
xnor U14431 (N_14431,N_14329,N_14144);
and U14432 (N_14432,N_14317,N_14239);
xnor U14433 (N_14433,N_14288,N_14193);
nand U14434 (N_14434,N_14112,N_14129);
nand U14435 (N_14435,N_14296,N_14154);
nor U14436 (N_14436,N_14186,N_14230);
xnor U14437 (N_14437,N_14184,N_14309);
xnor U14438 (N_14438,N_14286,N_14157);
nand U14439 (N_14439,N_14345,N_14280);
and U14440 (N_14440,N_14187,N_14347);
xor U14441 (N_14441,N_14343,N_14137);
xor U14442 (N_14442,N_14143,N_14231);
xor U14443 (N_14443,N_14359,N_14348);
nor U14444 (N_14444,N_14352,N_14146);
and U14445 (N_14445,N_14183,N_14255);
nor U14446 (N_14446,N_14395,N_14270);
nand U14447 (N_14447,N_14122,N_14391);
xor U14448 (N_14448,N_14303,N_14292);
and U14449 (N_14449,N_14388,N_14304);
nor U14450 (N_14450,N_14229,N_14338);
and U14451 (N_14451,N_14313,N_14209);
xor U14452 (N_14452,N_14178,N_14336);
and U14453 (N_14453,N_14235,N_14376);
nand U14454 (N_14454,N_14103,N_14390);
xnor U14455 (N_14455,N_14176,N_14109);
or U14456 (N_14456,N_14182,N_14170);
nand U14457 (N_14457,N_14234,N_14269);
xnor U14458 (N_14458,N_14351,N_14213);
and U14459 (N_14459,N_14165,N_14123);
nand U14460 (N_14460,N_14238,N_14295);
xnor U14461 (N_14461,N_14105,N_14278);
and U14462 (N_14462,N_14171,N_14311);
nand U14463 (N_14463,N_14279,N_14181);
xor U14464 (N_14464,N_14378,N_14220);
xnor U14465 (N_14465,N_14335,N_14163);
or U14466 (N_14466,N_14190,N_14195);
or U14467 (N_14467,N_14389,N_14243);
nand U14468 (N_14468,N_14328,N_14191);
or U14469 (N_14469,N_14215,N_14148);
nor U14470 (N_14470,N_14145,N_14194);
nor U14471 (N_14471,N_14212,N_14384);
xor U14472 (N_14472,N_14150,N_14316);
or U14473 (N_14473,N_14247,N_14349);
nand U14474 (N_14474,N_14232,N_14326);
nand U14475 (N_14475,N_14353,N_14218);
and U14476 (N_14476,N_14167,N_14158);
xnor U14477 (N_14477,N_14210,N_14252);
or U14478 (N_14478,N_14211,N_14363);
nand U14479 (N_14479,N_14192,N_14153);
xor U14480 (N_14480,N_14377,N_14169);
and U14481 (N_14481,N_14139,N_14331);
nand U14482 (N_14482,N_14214,N_14284);
or U14483 (N_14483,N_14161,N_14375);
and U14484 (N_14484,N_14175,N_14117);
nand U14485 (N_14485,N_14222,N_14204);
nand U14486 (N_14486,N_14314,N_14245);
or U14487 (N_14487,N_14371,N_14207);
or U14488 (N_14488,N_14127,N_14258);
nand U14489 (N_14489,N_14263,N_14200);
nand U14490 (N_14490,N_14244,N_14372);
nor U14491 (N_14491,N_14130,N_14385);
nand U14492 (N_14492,N_14358,N_14308);
or U14493 (N_14493,N_14367,N_14302);
or U14494 (N_14494,N_14126,N_14134);
xnor U14495 (N_14495,N_14306,N_14260);
or U14496 (N_14496,N_14141,N_14124);
nor U14497 (N_14497,N_14180,N_14174);
xnor U14498 (N_14498,N_14221,N_14397);
nor U14499 (N_14499,N_14394,N_14114);
or U14500 (N_14500,N_14226,N_14276);
xnor U14501 (N_14501,N_14312,N_14217);
nor U14502 (N_14502,N_14111,N_14225);
and U14503 (N_14503,N_14315,N_14380);
nor U14504 (N_14504,N_14267,N_14199);
nand U14505 (N_14505,N_14386,N_14301);
and U14506 (N_14506,N_14383,N_14289);
nor U14507 (N_14507,N_14290,N_14242);
xor U14508 (N_14508,N_14118,N_14360);
nor U14509 (N_14509,N_14354,N_14237);
nor U14510 (N_14510,N_14133,N_14119);
nor U14511 (N_14511,N_14266,N_14274);
nor U14512 (N_14512,N_14128,N_14356);
nor U14513 (N_14513,N_14341,N_14256);
nor U14514 (N_14514,N_14219,N_14228);
nor U14515 (N_14515,N_14374,N_14323);
nand U14516 (N_14516,N_14287,N_14102);
nand U14517 (N_14517,N_14382,N_14355);
or U14518 (N_14518,N_14173,N_14325);
and U14519 (N_14519,N_14285,N_14156);
nor U14520 (N_14520,N_14249,N_14100);
and U14521 (N_14521,N_14340,N_14283);
xor U14522 (N_14522,N_14261,N_14101);
xnor U14523 (N_14523,N_14185,N_14189);
xnor U14524 (N_14524,N_14369,N_14162);
or U14525 (N_14525,N_14155,N_14233);
xor U14526 (N_14526,N_14319,N_14201);
or U14527 (N_14527,N_14179,N_14264);
xor U14528 (N_14528,N_14281,N_14300);
nand U14529 (N_14529,N_14241,N_14294);
or U14530 (N_14530,N_14271,N_14106);
and U14531 (N_14531,N_14248,N_14297);
nor U14532 (N_14532,N_14299,N_14282);
xor U14533 (N_14533,N_14268,N_14197);
nor U14534 (N_14534,N_14254,N_14151);
or U14535 (N_14535,N_14298,N_14381);
and U14536 (N_14536,N_14125,N_14203);
nand U14537 (N_14537,N_14253,N_14318);
nor U14538 (N_14538,N_14152,N_14332);
nand U14539 (N_14539,N_14236,N_14361);
xor U14540 (N_14540,N_14379,N_14121);
nor U14541 (N_14541,N_14392,N_14364);
and U14542 (N_14542,N_14305,N_14334);
nor U14543 (N_14543,N_14387,N_14149);
and U14544 (N_14544,N_14321,N_14223);
nand U14545 (N_14545,N_14365,N_14373);
nand U14546 (N_14546,N_14257,N_14140);
nor U14547 (N_14547,N_14104,N_14202);
and U14548 (N_14548,N_14250,N_14293);
or U14549 (N_14549,N_14168,N_14206);
nor U14550 (N_14550,N_14363,N_14305);
nand U14551 (N_14551,N_14208,N_14203);
and U14552 (N_14552,N_14223,N_14103);
or U14553 (N_14553,N_14198,N_14340);
xnor U14554 (N_14554,N_14260,N_14255);
nand U14555 (N_14555,N_14398,N_14377);
and U14556 (N_14556,N_14304,N_14302);
xor U14557 (N_14557,N_14242,N_14282);
nand U14558 (N_14558,N_14331,N_14209);
and U14559 (N_14559,N_14120,N_14264);
nor U14560 (N_14560,N_14127,N_14269);
and U14561 (N_14561,N_14148,N_14199);
and U14562 (N_14562,N_14103,N_14288);
xnor U14563 (N_14563,N_14102,N_14309);
and U14564 (N_14564,N_14207,N_14329);
nor U14565 (N_14565,N_14203,N_14336);
nor U14566 (N_14566,N_14151,N_14294);
and U14567 (N_14567,N_14330,N_14169);
and U14568 (N_14568,N_14243,N_14207);
or U14569 (N_14569,N_14119,N_14370);
nor U14570 (N_14570,N_14349,N_14151);
nor U14571 (N_14571,N_14168,N_14178);
and U14572 (N_14572,N_14328,N_14113);
nand U14573 (N_14573,N_14390,N_14307);
nand U14574 (N_14574,N_14353,N_14299);
nor U14575 (N_14575,N_14212,N_14164);
xor U14576 (N_14576,N_14244,N_14187);
nand U14577 (N_14577,N_14289,N_14100);
nand U14578 (N_14578,N_14282,N_14106);
nor U14579 (N_14579,N_14325,N_14373);
and U14580 (N_14580,N_14115,N_14340);
or U14581 (N_14581,N_14263,N_14172);
nand U14582 (N_14582,N_14148,N_14176);
nand U14583 (N_14583,N_14398,N_14188);
nor U14584 (N_14584,N_14201,N_14357);
xor U14585 (N_14585,N_14282,N_14195);
nand U14586 (N_14586,N_14242,N_14100);
nand U14587 (N_14587,N_14369,N_14289);
nand U14588 (N_14588,N_14284,N_14250);
or U14589 (N_14589,N_14393,N_14229);
or U14590 (N_14590,N_14361,N_14398);
nand U14591 (N_14591,N_14301,N_14382);
or U14592 (N_14592,N_14229,N_14298);
nand U14593 (N_14593,N_14196,N_14263);
xor U14594 (N_14594,N_14364,N_14195);
and U14595 (N_14595,N_14242,N_14132);
nand U14596 (N_14596,N_14336,N_14377);
or U14597 (N_14597,N_14382,N_14231);
and U14598 (N_14598,N_14245,N_14117);
nor U14599 (N_14599,N_14308,N_14145);
and U14600 (N_14600,N_14336,N_14326);
or U14601 (N_14601,N_14169,N_14286);
nor U14602 (N_14602,N_14396,N_14341);
or U14603 (N_14603,N_14231,N_14287);
nor U14604 (N_14604,N_14320,N_14210);
nor U14605 (N_14605,N_14388,N_14271);
nor U14606 (N_14606,N_14271,N_14278);
and U14607 (N_14607,N_14250,N_14379);
and U14608 (N_14608,N_14244,N_14329);
or U14609 (N_14609,N_14217,N_14351);
and U14610 (N_14610,N_14166,N_14143);
or U14611 (N_14611,N_14222,N_14319);
nand U14612 (N_14612,N_14350,N_14223);
or U14613 (N_14613,N_14244,N_14241);
and U14614 (N_14614,N_14130,N_14184);
and U14615 (N_14615,N_14131,N_14247);
nand U14616 (N_14616,N_14267,N_14127);
and U14617 (N_14617,N_14368,N_14332);
nor U14618 (N_14618,N_14195,N_14262);
xnor U14619 (N_14619,N_14347,N_14339);
nand U14620 (N_14620,N_14207,N_14348);
nor U14621 (N_14621,N_14378,N_14344);
or U14622 (N_14622,N_14324,N_14157);
nand U14623 (N_14623,N_14182,N_14285);
and U14624 (N_14624,N_14257,N_14213);
nor U14625 (N_14625,N_14216,N_14347);
or U14626 (N_14626,N_14218,N_14279);
nand U14627 (N_14627,N_14183,N_14235);
and U14628 (N_14628,N_14381,N_14393);
nand U14629 (N_14629,N_14299,N_14298);
xnor U14630 (N_14630,N_14257,N_14267);
nor U14631 (N_14631,N_14140,N_14227);
nor U14632 (N_14632,N_14108,N_14317);
nor U14633 (N_14633,N_14329,N_14394);
and U14634 (N_14634,N_14139,N_14287);
and U14635 (N_14635,N_14250,N_14214);
nor U14636 (N_14636,N_14290,N_14297);
and U14637 (N_14637,N_14190,N_14123);
nand U14638 (N_14638,N_14208,N_14399);
and U14639 (N_14639,N_14368,N_14214);
nand U14640 (N_14640,N_14227,N_14218);
nor U14641 (N_14641,N_14150,N_14107);
xor U14642 (N_14642,N_14161,N_14387);
nand U14643 (N_14643,N_14286,N_14291);
nand U14644 (N_14644,N_14202,N_14375);
xor U14645 (N_14645,N_14283,N_14181);
xor U14646 (N_14646,N_14183,N_14179);
or U14647 (N_14647,N_14149,N_14252);
and U14648 (N_14648,N_14299,N_14158);
and U14649 (N_14649,N_14213,N_14363);
xor U14650 (N_14650,N_14317,N_14179);
xor U14651 (N_14651,N_14223,N_14228);
nor U14652 (N_14652,N_14158,N_14198);
xor U14653 (N_14653,N_14109,N_14188);
and U14654 (N_14654,N_14359,N_14309);
and U14655 (N_14655,N_14147,N_14221);
and U14656 (N_14656,N_14332,N_14395);
nor U14657 (N_14657,N_14327,N_14263);
and U14658 (N_14658,N_14281,N_14102);
nor U14659 (N_14659,N_14374,N_14320);
nor U14660 (N_14660,N_14214,N_14120);
nor U14661 (N_14661,N_14137,N_14223);
xnor U14662 (N_14662,N_14384,N_14322);
or U14663 (N_14663,N_14127,N_14161);
or U14664 (N_14664,N_14161,N_14278);
or U14665 (N_14665,N_14340,N_14126);
nand U14666 (N_14666,N_14344,N_14104);
nor U14667 (N_14667,N_14304,N_14267);
nor U14668 (N_14668,N_14194,N_14182);
or U14669 (N_14669,N_14159,N_14271);
xor U14670 (N_14670,N_14321,N_14154);
nor U14671 (N_14671,N_14211,N_14325);
xnor U14672 (N_14672,N_14323,N_14177);
nand U14673 (N_14673,N_14147,N_14335);
xnor U14674 (N_14674,N_14134,N_14232);
and U14675 (N_14675,N_14395,N_14365);
and U14676 (N_14676,N_14326,N_14197);
nor U14677 (N_14677,N_14234,N_14385);
nor U14678 (N_14678,N_14155,N_14344);
or U14679 (N_14679,N_14152,N_14158);
xnor U14680 (N_14680,N_14282,N_14152);
and U14681 (N_14681,N_14223,N_14378);
nor U14682 (N_14682,N_14185,N_14126);
nor U14683 (N_14683,N_14395,N_14198);
nor U14684 (N_14684,N_14113,N_14137);
xnor U14685 (N_14685,N_14398,N_14339);
xnor U14686 (N_14686,N_14178,N_14108);
nand U14687 (N_14687,N_14170,N_14343);
and U14688 (N_14688,N_14186,N_14365);
nor U14689 (N_14689,N_14208,N_14151);
nand U14690 (N_14690,N_14161,N_14143);
or U14691 (N_14691,N_14312,N_14303);
or U14692 (N_14692,N_14107,N_14189);
or U14693 (N_14693,N_14346,N_14143);
nor U14694 (N_14694,N_14123,N_14148);
or U14695 (N_14695,N_14155,N_14250);
nand U14696 (N_14696,N_14254,N_14209);
xor U14697 (N_14697,N_14375,N_14211);
and U14698 (N_14698,N_14216,N_14188);
nor U14699 (N_14699,N_14242,N_14199);
and U14700 (N_14700,N_14431,N_14636);
or U14701 (N_14701,N_14417,N_14486);
and U14702 (N_14702,N_14670,N_14504);
and U14703 (N_14703,N_14613,N_14661);
nand U14704 (N_14704,N_14533,N_14526);
or U14705 (N_14705,N_14592,N_14529);
or U14706 (N_14706,N_14691,N_14481);
xor U14707 (N_14707,N_14425,N_14462);
nor U14708 (N_14708,N_14400,N_14472);
xnor U14709 (N_14709,N_14510,N_14513);
or U14710 (N_14710,N_14604,N_14470);
nand U14711 (N_14711,N_14679,N_14685);
xor U14712 (N_14712,N_14469,N_14515);
xnor U14713 (N_14713,N_14508,N_14501);
or U14714 (N_14714,N_14578,N_14642);
nor U14715 (N_14715,N_14505,N_14522);
and U14716 (N_14716,N_14457,N_14506);
nand U14717 (N_14717,N_14421,N_14493);
and U14718 (N_14718,N_14484,N_14408);
nand U14719 (N_14719,N_14488,N_14567);
or U14720 (N_14720,N_14478,N_14581);
nor U14721 (N_14721,N_14420,N_14656);
xnor U14722 (N_14722,N_14518,N_14694);
xor U14723 (N_14723,N_14650,N_14638);
nor U14724 (N_14724,N_14449,N_14673);
xnor U14725 (N_14725,N_14445,N_14614);
xnor U14726 (N_14726,N_14623,N_14659);
xor U14727 (N_14727,N_14627,N_14680);
or U14728 (N_14728,N_14464,N_14626);
and U14729 (N_14729,N_14557,N_14499);
xor U14730 (N_14730,N_14519,N_14692);
xnor U14731 (N_14731,N_14619,N_14559);
xor U14732 (N_14732,N_14476,N_14637);
xor U14733 (N_14733,N_14450,N_14528);
nor U14734 (N_14734,N_14566,N_14612);
xnor U14735 (N_14735,N_14547,N_14647);
nor U14736 (N_14736,N_14418,N_14683);
nand U14737 (N_14737,N_14684,N_14514);
nor U14738 (N_14738,N_14432,N_14439);
nand U14739 (N_14739,N_14536,N_14452);
xor U14740 (N_14740,N_14459,N_14575);
or U14741 (N_14741,N_14410,N_14534);
xnor U14742 (N_14742,N_14532,N_14696);
nand U14743 (N_14743,N_14444,N_14668);
or U14744 (N_14744,N_14453,N_14573);
and U14745 (N_14745,N_14548,N_14468);
and U14746 (N_14746,N_14615,N_14460);
nand U14747 (N_14747,N_14535,N_14690);
and U14748 (N_14748,N_14697,N_14560);
xnor U14749 (N_14749,N_14549,N_14412);
nand U14750 (N_14750,N_14479,N_14561);
or U14751 (N_14751,N_14585,N_14482);
and U14752 (N_14752,N_14599,N_14541);
nor U14753 (N_14753,N_14456,N_14569);
and U14754 (N_14754,N_14563,N_14525);
xnor U14755 (N_14755,N_14667,N_14671);
or U14756 (N_14756,N_14609,N_14674);
nor U14757 (N_14757,N_14631,N_14660);
nand U14758 (N_14758,N_14639,N_14666);
nand U14759 (N_14759,N_14454,N_14562);
or U14760 (N_14760,N_14507,N_14620);
xnor U14761 (N_14761,N_14429,N_14540);
xnor U14762 (N_14762,N_14428,N_14406);
and U14763 (N_14763,N_14583,N_14448);
and U14764 (N_14764,N_14437,N_14698);
nor U14765 (N_14765,N_14648,N_14676);
xnor U14766 (N_14766,N_14570,N_14404);
xor U14767 (N_14767,N_14621,N_14544);
nor U14768 (N_14768,N_14682,N_14628);
nor U14769 (N_14769,N_14577,N_14405);
nor U14770 (N_14770,N_14584,N_14589);
nor U14771 (N_14771,N_14601,N_14531);
xor U14772 (N_14772,N_14490,N_14669);
or U14773 (N_14773,N_14542,N_14603);
nor U14774 (N_14774,N_14530,N_14443);
nand U14775 (N_14775,N_14537,N_14554);
nand U14776 (N_14776,N_14430,N_14538);
and U14777 (N_14777,N_14401,N_14664);
nor U14778 (N_14778,N_14424,N_14641);
nor U14779 (N_14779,N_14672,N_14665);
nor U14780 (N_14780,N_14571,N_14610);
nand U14781 (N_14781,N_14591,N_14632);
and U14782 (N_14782,N_14625,N_14447);
and U14783 (N_14783,N_14624,N_14503);
nand U14784 (N_14784,N_14527,N_14555);
nor U14785 (N_14785,N_14695,N_14588);
nor U14786 (N_14786,N_14477,N_14579);
and U14787 (N_14787,N_14618,N_14416);
xor U14788 (N_14788,N_14442,N_14688);
nor U14789 (N_14789,N_14458,N_14658);
nand U14790 (N_14790,N_14471,N_14580);
and U14791 (N_14791,N_14582,N_14440);
nor U14792 (N_14792,N_14550,N_14596);
nor U14793 (N_14793,N_14500,N_14520);
or U14794 (N_14794,N_14523,N_14423);
nor U14795 (N_14795,N_14643,N_14480);
and U14796 (N_14796,N_14657,N_14556);
or U14797 (N_14797,N_14496,N_14415);
or U14798 (N_14798,N_14494,N_14622);
nand U14799 (N_14799,N_14605,N_14606);
xor U14800 (N_14800,N_14539,N_14646);
xor U14801 (N_14801,N_14644,N_14699);
nand U14802 (N_14802,N_14593,N_14465);
nor U14803 (N_14803,N_14436,N_14433);
nand U14804 (N_14804,N_14630,N_14546);
nor U14805 (N_14805,N_14511,N_14446);
or U14806 (N_14806,N_14524,N_14543);
and U14807 (N_14807,N_14434,N_14497);
or U14808 (N_14808,N_14414,N_14487);
and U14809 (N_14809,N_14597,N_14595);
nand U14810 (N_14810,N_14652,N_14435);
and U14811 (N_14811,N_14427,N_14681);
xnor U14812 (N_14812,N_14586,N_14441);
and U14813 (N_14813,N_14413,N_14655);
nand U14814 (N_14814,N_14675,N_14629);
or U14815 (N_14815,N_14686,N_14576);
or U14816 (N_14816,N_14616,N_14640);
nor U14817 (N_14817,N_14483,N_14634);
and U14818 (N_14818,N_14502,N_14635);
nand U14819 (N_14819,N_14689,N_14426);
and U14820 (N_14820,N_14411,N_14498);
nand U14821 (N_14821,N_14489,N_14617);
or U14822 (N_14822,N_14572,N_14492);
xnor U14823 (N_14823,N_14693,N_14552);
nor U14824 (N_14824,N_14590,N_14565);
xnor U14825 (N_14825,N_14687,N_14466);
or U14826 (N_14826,N_14422,N_14463);
xnor U14827 (N_14827,N_14516,N_14608);
or U14828 (N_14828,N_14568,N_14633);
xor U14829 (N_14829,N_14512,N_14663);
or U14830 (N_14830,N_14600,N_14553);
nand U14831 (N_14831,N_14611,N_14409);
xor U14832 (N_14832,N_14654,N_14677);
nand U14833 (N_14833,N_14594,N_14455);
or U14834 (N_14834,N_14485,N_14509);
nor U14835 (N_14835,N_14587,N_14662);
or U14836 (N_14836,N_14602,N_14473);
nor U14837 (N_14837,N_14545,N_14607);
xnor U14838 (N_14838,N_14419,N_14558);
nand U14839 (N_14839,N_14521,N_14517);
xnor U14840 (N_14840,N_14649,N_14402);
nor U14841 (N_14841,N_14564,N_14491);
and U14842 (N_14842,N_14653,N_14574);
nor U14843 (N_14843,N_14651,N_14678);
and U14844 (N_14844,N_14474,N_14461);
or U14845 (N_14845,N_14467,N_14598);
xnor U14846 (N_14846,N_14645,N_14438);
nand U14847 (N_14847,N_14475,N_14407);
xnor U14848 (N_14848,N_14451,N_14403);
or U14849 (N_14849,N_14551,N_14495);
nand U14850 (N_14850,N_14525,N_14600);
or U14851 (N_14851,N_14587,N_14540);
or U14852 (N_14852,N_14444,N_14412);
or U14853 (N_14853,N_14490,N_14406);
nand U14854 (N_14854,N_14590,N_14474);
and U14855 (N_14855,N_14435,N_14404);
or U14856 (N_14856,N_14655,N_14403);
or U14857 (N_14857,N_14464,N_14452);
nand U14858 (N_14858,N_14555,N_14483);
or U14859 (N_14859,N_14679,N_14483);
or U14860 (N_14860,N_14448,N_14590);
or U14861 (N_14861,N_14597,N_14509);
nand U14862 (N_14862,N_14519,N_14621);
xor U14863 (N_14863,N_14531,N_14425);
or U14864 (N_14864,N_14646,N_14561);
xnor U14865 (N_14865,N_14636,N_14433);
or U14866 (N_14866,N_14420,N_14446);
nor U14867 (N_14867,N_14627,N_14685);
nand U14868 (N_14868,N_14468,N_14400);
and U14869 (N_14869,N_14422,N_14586);
xor U14870 (N_14870,N_14616,N_14650);
or U14871 (N_14871,N_14484,N_14558);
or U14872 (N_14872,N_14494,N_14600);
nor U14873 (N_14873,N_14567,N_14523);
and U14874 (N_14874,N_14450,N_14639);
xnor U14875 (N_14875,N_14671,N_14611);
xnor U14876 (N_14876,N_14432,N_14613);
xor U14877 (N_14877,N_14484,N_14490);
or U14878 (N_14878,N_14515,N_14548);
nand U14879 (N_14879,N_14599,N_14433);
nand U14880 (N_14880,N_14480,N_14569);
and U14881 (N_14881,N_14483,N_14611);
and U14882 (N_14882,N_14430,N_14676);
and U14883 (N_14883,N_14525,N_14581);
or U14884 (N_14884,N_14417,N_14527);
and U14885 (N_14885,N_14576,N_14402);
nor U14886 (N_14886,N_14450,N_14690);
and U14887 (N_14887,N_14546,N_14566);
nand U14888 (N_14888,N_14432,N_14652);
and U14889 (N_14889,N_14411,N_14461);
and U14890 (N_14890,N_14562,N_14648);
nand U14891 (N_14891,N_14622,N_14528);
nor U14892 (N_14892,N_14436,N_14459);
nor U14893 (N_14893,N_14409,N_14509);
xnor U14894 (N_14894,N_14684,N_14564);
xnor U14895 (N_14895,N_14673,N_14650);
nand U14896 (N_14896,N_14688,N_14460);
and U14897 (N_14897,N_14633,N_14550);
or U14898 (N_14898,N_14422,N_14466);
xor U14899 (N_14899,N_14473,N_14506);
or U14900 (N_14900,N_14583,N_14669);
and U14901 (N_14901,N_14657,N_14572);
nand U14902 (N_14902,N_14571,N_14536);
or U14903 (N_14903,N_14663,N_14692);
nor U14904 (N_14904,N_14588,N_14673);
nand U14905 (N_14905,N_14688,N_14648);
nand U14906 (N_14906,N_14567,N_14532);
nor U14907 (N_14907,N_14696,N_14497);
and U14908 (N_14908,N_14482,N_14436);
and U14909 (N_14909,N_14571,N_14503);
and U14910 (N_14910,N_14433,N_14426);
xnor U14911 (N_14911,N_14500,N_14545);
nor U14912 (N_14912,N_14591,N_14522);
xor U14913 (N_14913,N_14574,N_14465);
or U14914 (N_14914,N_14430,N_14695);
or U14915 (N_14915,N_14696,N_14593);
nor U14916 (N_14916,N_14448,N_14497);
xnor U14917 (N_14917,N_14490,N_14530);
or U14918 (N_14918,N_14668,N_14619);
xnor U14919 (N_14919,N_14638,N_14670);
nor U14920 (N_14920,N_14531,N_14658);
or U14921 (N_14921,N_14564,N_14566);
and U14922 (N_14922,N_14541,N_14508);
nand U14923 (N_14923,N_14506,N_14618);
and U14924 (N_14924,N_14462,N_14694);
nand U14925 (N_14925,N_14687,N_14481);
nor U14926 (N_14926,N_14484,N_14628);
xnor U14927 (N_14927,N_14575,N_14460);
or U14928 (N_14928,N_14693,N_14486);
or U14929 (N_14929,N_14427,N_14505);
xor U14930 (N_14930,N_14468,N_14422);
or U14931 (N_14931,N_14563,N_14474);
or U14932 (N_14932,N_14639,N_14577);
nor U14933 (N_14933,N_14546,N_14417);
or U14934 (N_14934,N_14686,N_14605);
xnor U14935 (N_14935,N_14487,N_14567);
and U14936 (N_14936,N_14633,N_14414);
xor U14937 (N_14937,N_14489,N_14447);
nand U14938 (N_14938,N_14514,N_14600);
nand U14939 (N_14939,N_14517,N_14694);
and U14940 (N_14940,N_14504,N_14547);
or U14941 (N_14941,N_14593,N_14420);
nand U14942 (N_14942,N_14593,N_14545);
xnor U14943 (N_14943,N_14622,N_14590);
xnor U14944 (N_14944,N_14673,N_14682);
or U14945 (N_14945,N_14676,N_14569);
nand U14946 (N_14946,N_14647,N_14533);
and U14947 (N_14947,N_14582,N_14588);
and U14948 (N_14948,N_14682,N_14445);
nand U14949 (N_14949,N_14525,N_14604);
or U14950 (N_14950,N_14476,N_14460);
and U14951 (N_14951,N_14648,N_14554);
nor U14952 (N_14952,N_14573,N_14697);
nand U14953 (N_14953,N_14616,N_14486);
nor U14954 (N_14954,N_14495,N_14403);
and U14955 (N_14955,N_14648,N_14691);
xor U14956 (N_14956,N_14637,N_14454);
nand U14957 (N_14957,N_14409,N_14454);
nand U14958 (N_14958,N_14607,N_14658);
nand U14959 (N_14959,N_14441,N_14408);
xor U14960 (N_14960,N_14445,N_14628);
nand U14961 (N_14961,N_14425,N_14541);
nor U14962 (N_14962,N_14565,N_14495);
and U14963 (N_14963,N_14656,N_14673);
nor U14964 (N_14964,N_14582,N_14473);
and U14965 (N_14965,N_14643,N_14662);
xnor U14966 (N_14966,N_14611,N_14402);
or U14967 (N_14967,N_14583,N_14540);
nand U14968 (N_14968,N_14618,N_14552);
or U14969 (N_14969,N_14456,N_14555);
nor U14970 (N_14970,N_14696,N_14610);
or U14971 (N_14971,N_14520,N_14494);
and U14972 (N_14972,N_14695,N_14678);
nor U14973 (N_14973,N_14615,N_14581);
or U14974 (N_14974,N_14448,N_14488);
xor U14975 (N_14975,N_14625,N_14549);
nand U14976 (N_14976,N_14577,N_14687);
and U14977 (N_14977,N_14551,N_14530);
nand U14978 (N_14978,N_14469,N_14651);
and U14979 (N_14979,N_14503,N_14569);
and U14980 (N_14980,N_14614,N_14463);
or U14981 (N_14981,N_14415,N_14536);
nor U14982 (N_14982,N_14578,N_14438);
and U14983 (N_14983,N_14573,N_14689);
nor U14984 (N_14984,N_14516,N_14659);
or U14985 (N_14985,N_14529,N_14621);
nand U14986 (N_14986,N_14437,N_14489);
nor U14987 (N_14987,N_14566,N_14404);
and U14988 (N_14988,N_14428,N_14613);
xor U14989 (N_14989,N_14535,N_14611);
and U14990 (N_14990,N_14403,N_14490);
and U14991 (N_14991,N_14564,N_14426);
and U14992 (N_14992,N_14601,N_14486);
or U14993 (N_14993,N_14697,N_14635);
xor U14994 (N_14994,N_14506,N_14559);
nor U14995 (N_14995,N_14482,N_14598);
nor U14996 (N_14996,N_14571,N_14615);
xnor U14997 (N_14997,N_14543,N_14586);
xor U14998 (N_14998,N_14405,N_14543);
nand U14999 (N_14999,N_14507,N_14634);
or U15000 (N_15000,N_14761,N_14937);
or U15001 (N_15001,N_14791,N_14836);
nor U15002 (N_15002,N_14751,N_14844);
nand U15003 (N_15003,N_14883,N_14725);
or U15004 (N_15004,N_14955,N_14788);
or U15005 (N_15005,N_14927,N_14884);
and U15006 (N_15006,N_14740,N_14821);
nor U15007 (N_15007,N_14799,N_14762);
nor U15008 (N_15008,N_14841,N_14926);
nor U15009 (N_15009,N_14874,N_14909);
nand U15010 (N_15010,N_14940,N_14952);
and U15011 (N_15011,N_14907,N_14916);
xor U15012 (N_15012,N_14819,N_14818);
nor U15013 (N_15013,N_14896,N_14820);
or U15014 (N_15014,N_14864,N_14815);
nand U15015 (N_15015,N_14833,N_14746);
nand U15016 (N_15016,N_14797,N_14950);
nor U15017 (N_15017,N_14806,N_14882);
xor U15018 (N_15018,N_14742,N_14838);
nand U15019 (N_15019,N_14914,N_14880);
nand U15020 (N_15020,N_14856,N_14723);
xor U15021 (N_15021,N_14703,N_14812);
nand U15022 (N_15022,N_14832,N_14890);
nand U15023 (N_15023,N_14973,N_14996);
nand U15024 (N_15024,N_14750,N_14872);
nor U15025 (N_15025,N_14700,N_14911);
nor U15026 (N_15026,N_14803,N_14877);
or U15027 (N_15027,N_14974,N_14736);
and U15028 (N_15028,N_14816,N_14990);
nand U15029 (N_15029,N_14727,N_14928);
and U15030 (N_15030,N_14733,N_14902);
nor U15031 (N_15031,N_14847,N_14886);
nor U15032 (N_15032,N_14991,N_14946);
xor U15033 (N_15033,N_14767,N_14845);
xnor U15034 (N_15034,N_14891,N_14861);
xor U15035 (N_15035,N_14936,N_14830);
nand U15036 (N_15036,N_14867,N_14939);
and U15037 (N_15037,N_14828,N_14855);
or U15038 (N_15038,N_14732,N_14726);
nor U15039 (N_15039,N_14729,N_14715);
nand U15040 (N_15040,N_14905,N_14802);
nor U15041 (N_15041,N_14889,N_14849);
xnor U15042 (N_15042,N_14798,N_14810);
nor U15043 (N_15043,N_14994,N_14941);
or U15044 (N_15044,N_14826,N_14846);
or U15045 (N_15045,N_14784,N_14707);
or U15046 (N_15046,N_14900,N_14717);
or U15047 (N_15047,N_14962,N_14869);
xnor U15048 (N_15048,N_14748,N_14910);
nand U15049 (N_15049,N_14716,N_14858);
and U15050 (N_15050,N_14992,N_14712);
or U15051 (N_15051,N_14702,N_14997);
nand U15052 (N_15052,N_14731,N_14967);
xnor U15053 (N_15053,N_14879,N_14756);
xnor U15054 (N_15054,N_14829,N_14852);
or U15055 (N_15055,N_14888,N_14765);
and U15056 (N_15056,N_14722,N_14839);
nand U15057 (N_15057,N_14972,N_14778);
and U15058 (N_15058,N_14814,N_14876);
xnor U15059 (N_15059,N_14899,N_14737);
xnor U15060 (N_15060,N_14711,N_14921);
and U15061 (N_15061,N_14753,N_14908);
nor U15062 (N_15062,N_14773,N_14948);
nor U15063 (N_15063,N_14998,N_14735);
xnor U15064 (N_15064,N_14957,N_14875);
or U15065 (N_15065,N_14979,N_14837);
xor U15066 (N_15066,N_14929,N_14747);
and U15067 (N_15067,N_14840,N_14989);
and U15068 (N_15068,N_14808,N_14904);
nor U15069 (N_15069,N_14730,N_14713);
nor U15070 (N_15070,N_14906,N_14757);
or U15071 (N_15071,N_14790,N_14924);
or U15072 (N_15072,N_14705,N_14987);
nand U15073 (N_15073,N_14787,N_14878);
nand U15074 (N_15074,N_14734,N_14807);
or U15075 (N_15075,N_14986,N_14817);
nor U15076 (N_15076,N_14918,N_14744);
nor U15077 (N_15077,N_14868,N_14759);
and U15078 (N_15078,N_14776,N_14963);
xnor U15079 (N_15079,N_14801,N_14894);
nand U15080 (N_15080,N_14993,N_14898);
or U15081 (N_15081,N_14981,N_14971);
nand U15082 (N_15082,N_14789,N_14718);
xnor U15083 (N_15083,N_14854,N_14701);
nand U15084 (N_15084,N_14831,N_14745);
nand U15085 (N_15085,N_14942,N_14796);
nand U15086 (N_15086,N_14708,N_14741);
nor U15087 (N_15087,N_14704,N_14755);
nand U15088 (N_15088,N_14983,N_14925);
xor U15089 (N_15089,N_14714,N_14920);
nand U15090 (N_15090,N_14775,N_14811);
nand U15091 (N_15091,N_14724,N_14739);
xnor U15092 (N_15092,N_14822,N_14738);
xnor U15093 (N_15093,N_14842,N_14934);
nand U15094 (N_15094,N_14795,N_14961);
nor U15095 (N_15095,N_14719,N_14785);
or U15096 (N_15096,N_14794,N_14976);
xor U15097 (N_15097,N_14771,N_14786);
or U15098 (N_15098,N_14763,N_14980);
nand U15099 (N_15099,N_14930,N_14871);
and U15100 (N_15100,N_14985,N_14709);
nor U15101 (N_15101,N_14932,N_14706);
nand U15102 (N_15102,N_14827,N_14947);
or U15103 (N_15103,N_14848,N_14922);
xnor U15104 (N_15104,N_14933,N_14804);
xor U15105 (N_15105,N_14768,N_14865);
nor U15106 (N_15106,N_14988,N_14859);
xnor U15107 (N_15107,N_14766,N_14923);
nor U15108 (N_15108,N_14862,N_14721);
nor U15109 (N_15109,N_14968,N_14866);
and U15110 (N_15110,N_14857,N_14720);
xnor U15111 (N_15111,N_14885,N_14792);
xnor U15112 (N_15112,N_14823,N_14728);
and U15113 (N_15113,N_14710,N_14958);
and U15114 (N_15114,N_14938,N_14977);
or U15115 (N_15115,N_14897,N_14964);
nor U15116 (N_15116,N_14944,N_14860);
xnor U15117 (N_15117,N_14999,N_14887);
and U15118 (N_15118,N_14982,N_14893);
or U15119 (N_15119,N_14913,N_14758);
nor U15120 (N_15120,N_14749,N_14912);
and U15121 (N_15121,N_14960,N_14774);
nor U15122 (N_15122,N_14813,N_14824);
and U15123 (N_15123,N_14978,N_14770);
nor U15124 (N_15124,N_14769,N_14805);
nand U15125 (N_15125,N_14892,N_14975);
nor U15126 (N_15126,N_14772,N_14903);
or U15127 (N_15127,N_14943,N_14895);
nor U15128 (N_15128,N_14931,N_14984);
xor U15129 (N_15129,N_14901,N_14835);
and U15130 (N_15130,N_14853,N_14954);
nand U15131 (N_15131,N_14919,N_14870);
nand U15132 (N_15132,N_14969,N_14935);
and U15133 (N_15133,N_14917,N_14953);
and U15134 (N_15134,N_14825,N_14951);
xnor U15135 (N_15135,N_14873,N_14743);
xnor U15136 (N_15136,N_14965,N_14945);
and U15137 (N_15137,N_14959,N_14850);
xor U15138 (N_15138,N_14966,N_14754);
xnor U15139 (N_15139,N_14764,N_14881);
nand U15140 (N_15140,N_14793,N_14777);
nand U15141 (N_15141,N_14843,N_14780);
and U15142 (N_15142,N_14809,N_14781);
or U15143 (N_15143,N_14834,N_14915);
xnor U15144 (N_15144,N_14970,N_14851);
or U15145 (N_15145,N_14783,N_14752);
and U15146 (N_15146,N_14779,N_14949);
xnor U15147 (N_15147,N_14956,N_14863);
xnor U15148 (N_15148,N_14760,N_14995);
and U15149 (N_15149,N_14782,N_14800);
nor U15150 (N_15150,N_14910,N_14962);
nor U15151 (N_15151,N_14737,N_14731);
nor U15152 (N_15152,N_14901,N_14871);
nor U15153 (N_15153,N_14853,N_14725);
xnor U15154 (N_15154,N_14907,N_14708);
xnor U15155 (N_15155,N_14914,N_14930);
nand U15156 (N_15156,N_14759,N_14815);
nor U15157 (N_15157,N_14881,N_14897);
nor U15158 (N_15158,N_14838,N_14961);
nor U15159 (N_15159,N_14852,N_14807);
and U15160 (N_15160,N_14722,N_14761);
nor U15161 (N_15161,N_14763,N_14707);
and U15162 (N_15162,N_14790,N_14862);
nand U15163 (N_15163,N_14889,N_14865);
xnor U15164 (N_15164,N_14763,N_14708);
and U15165 (N_15165,N_14862,N_14831);
nand U15166 (N_15166,N_14761,N_14885);
or U15167 (N_15167,N_14865,N_14946);
or U15168 (N_15168,N_14842,N_14909);
and U15169 (N_15169,N_14772,N_14994);
nor U15170 (N_15170,N_14978,N_14989);
nand U15171 (N_15171,N_14795,N_14774);
nor U15172 (N_15172,N_14856,N_14994);
and U15173 (N_15173,N_14783,N_14833);
xnor U15174 (N_15174,N_14717,N_14765);
nor U15175 (N_15175,N_14774,N_14730);
nand U15176 (N_15176,N_14881,N_14852);
nand U15177 (N_15177,N_14857,N_14951);
xor U15178 (N_15178,N_14743,N_14976);
or U15179 (N_15179,N_14817,N_14718);
nand U15180 (N_15180,N_14890,N_14766);
nor U15181 (N_15181,N_14874,N_14813);
nand U15182 (N_15182,N_14903,N_14702);
and U15183 (N_15183,N_14756,N_14742);
nand U15184 (N_15184,N_14841,N_14824);
nor U15185 (N_15185,N_14902,N_14763);
and U15186 (N_15186,N_14920,N_14872);
xnor U15187 (N_15187,N_14864,N_14843);
and U15188 (N_15188,N_14967,N_14825);
nand U15189 (N_15189,N_14880,N_14769);
xor U15190 (N_15190,N_14744,N_14892);
and U15191 (N_15191,N_14896,N_14753);
xnor U15192 (N_15192,N_14812,N_14918);
nor U15193 (N_15193,N_14758,N_14881);
nand U15194 (N_15194,N_14731,N_14909);
and U15195 (N_15195,N_14956,N_14770);
nor U15196 (N_15196,N_14932,N_14878);
xor U15197 (N_15197,N_14840,N_14996);
nand U15198 (N_15198,N_14993,N_14987);
nand U15199 (N_15199,N_14923,N_14909);
or U15200 (N_15200,N_14997,N_14730);
nor U15201 (N_15201,N_14970,N_14783);
or U15202 (N_15202,N_14836,N_14701);
nand U15203 (N_15203,N_14806,N_14802);
nand U15204 (N_15204,N_14722,N_14978);
or U15205 (N_15205,N_14763,N_14788);
xnor U15206 (N_15206,N_14918,N_14883);
xnor U15207 (N_15207,N_14768,N_14750);
xnor U15208 (N_15208,N_14890,N_14721);
and U15209 (N_15209,N_14948,N_14722);
or U15210 (N_15210,N_14852,N_14817);
nor U15211 (N_15211,N_14747,N_14958);
xor U15212 (N_15212,N_14793,N_14967);
xor U15213 (N_15213,N_14724,N_14747);
or U15214 (N_15214,N_14872,N_14801);
nor U15215 (N_15215,N_14887,N_14953);
nand U15216 (N_15216,N_14802,N_14708);
nand U15217 (N_15217,N_14902,N_14949);
nand U15218 (N_15218,N_14810,N_14814);
or U15219 (N_15219,N_14704,N_14917);
nor U15220 (N_15220,N_14838,N_14754);
or U15221 (N_15221,N_14929,N_14879);
or U15222 (N_15222,N_14907,N_14717);
and U15223 (N_15223,N_14743,N_14988);
and U15224 (N_15224,N_14926,N_14976);
or U15225 (N_15225,N_14932,N_14908);
and U15226 (N_15226,N_14706,N_14813);
xnor U15227 (N_15227,N_14852,N_14911);
or U15228 (N_15228,N_14864,N_14803);
nand U15229 (N_15229,N_14729,N_14918);
or U15230 (N_15230,N_14780,N_14714);
xor U15231 (N_15231,N_14859,N_14930);
nor U15232 (N_15232,N_14877,N_14743);
nor U15233 (N_15233,N_14797,N_14789);
or U15234 (N_15234,N_14990,N_14966);
xnor U15235 (N_15235,N_14705,N_14804);
or U15236 (N_15236,N_14781,N_14808);
and U15237 (N_15237,N_14711,N_14723);
xor U15238 (N_15238,N_14891,N_14789);
nor U15239 (N_15239,N_14909,N_14939);
nand U15240 (N_15240,N_14888,N_14991);
xor U15241 (N_15241,N_14715,N_14786);
nand U15242 (N_15242,N_14933,N_14964);
nor U15243 (N_15243,N_14845,N_14941);
xnor U15244 (N_15244,N_14812,N_14872);
and U15245 (N_15245,N_14943,N_14811);
nor U15246 (N_15246,N_14821,N_14946);
and U15247 (N_15247,N_14747,N_14824);
or U15248 (N_15248,N_14812,N_14855);
and U15249 (N_15249,N_14850,N_14754);
or U15250 (N_15250,N_14743,N_14851);
nor U15251 (N_15251,N_14784,N_14793);
and U15252 (N_15252,N_14806,N_14950);
xor U15253 (N_15253,N_14903,N_14994);
and U15254 (N_15254,N_14845,N_14834);
xnor U15255 (N_15255,N_14939,N_14737);
nor U15256 (N_15256,N_14919,N_14798);
nor U15257 (N_15257,N_14817,N_14803);
nand U15258 (N_15258,N_14792,N_14830);
nor U15259 (N_15259,N_14971,N_14903);
nor U15260 (N_15260,N_14769,N_14841);
xnor U15261 (N_15261,N_14919,N_14878);
nand U15262 (N_15262,N_14864,N_14919);
and U15263 (N_15263,N_14874,N_14953);
xor U15264 (N_15264,N_14935,N_14805);
xnor U15265 (N_15265,N_14972,N_14739);
nand U15266 (N_15266,N_14725,N_14842);
or U15267 (N_15267,N_14862,N_14963);
or U15268 (N_15268,N_14911,N_14930);
nand U15269 (N_15269,N_14714,N_14812);
nand U15270 (N_15270,N_14810,N_14919);
and U15271 (N_15271,N_14867,N_14963);
nor U15272 (N_15272,N_14864,N_14969);
and U15273 (N_15273,N_14794,N_14826);
nand U15274 (N_15274,N_14904,N_14713);
xor U15275 (N_15275,N_14824,N_14878);
and U15276 (N_15276,N_14966,N_14974);
nor U15277 (N_15277,N_14992,N_14871);
nor U15278 (N_15278,N_14915,N_14719);
xor U15279 (N_15279,N_14804,N_14808);
nor U15280 (N_15280,N_14847,N_14990);
and U15281 (N_15281,N_14852,N_14899);
nor U15282 (N_15282,N_14781,N_14991);
xnor U15283 (N_15283,N_14757,N_14883);
xor U15284 (N_15284,N_14833,N_14920);
nand U15285 (N_15285,N_14886,N_14894);
and U15286 (N_15286,N_14727,N_14842);
xnor U15287 (N_15287,N_14880,N_14744);
xnor U15288 (N_15288,N_14828,N_14995);
nand U15289 (N_15289,N_14886,N_14878);
or U15290 (N_15290,N_14779,N_14903);
and U15291 (N_15291,N_14879,N_14903);
nand U15292 (N_15292,N_14993,N_14853);
nor U15293 (N_15293,N_14756,N_14988);
and U15294 (N_15294,N_14894,N_14994);
xor U15295 (N_15295,N_14827,N_14789);
nor U15296 (N_15296,N_14905,N_14932);
or U15297 (N_15297,N_14923,N_14790);
or U15298 (N_15298,N_14965,N_14917);
and U15299 (N_15299,N_14724,N_14718);
nand U15300 (N_15300,N_15165,N_15117);
or U15301 (N_15301,N_15064,N_15191);
nor U15302 (N_15302,N_15183,N_15175);
xnor U15303 (N_15303,N_15144,N_15101);
and U15304 (N_15304,N_15107,N_15015);
or U15305 (N_15305,N_15072,N_15029);
xnor U15306 (N_15306,N_15155,N_15031);
nand U15307 (N_15307,N_15263,N_15267);
nand U15308 (N_15308,N_15289,N_15042);
nand U15309 (N_15309,N_15136,N_15210);
xnor U15310 (N_15310,N_15141,N_15279);
or U15311 (N_15311,N_15185,N_15124);
and U15312 (N_15312,N_15243,N_15250);
nand U15313 (N_15313,N_15028,N_15208);
and U15314 (N_15314,N_15054,N_15036);
xor U15315 (N_15315,N_15195,N_15079);
nor U15316 (N_15316,N_15179,N_15019);
nand U15317 (N_15317,N_15159,N_15190);
nor U15318 (N_15318,N_15080,N_15166);
nor U15319 (N_15319,N_15253,N_15236);
nor U15320 (N_15320,N_15090,N_15286);
or U15321 (N_15321,N_15131,N_15003);
and U15322 (N_15322,N_15041,N_15120);
and U15323 (N_15323,N_15039,N_15094);
nand U15324 (N_15324,N_15017,N_15061);
nand U15325 (N_15325,N_15298,N_15199);
nand U15326 (N_15326,N_15266,N_15034);
and U15327 (N_15327,N_15122,N_15071);
or U15328 (N_15328,N_15239,N_15085);
nor U15329 (N_15329,N_15128,N_15249);
and U15330 (N_15330,N_15035,N_15009);
xnor U15331 (N_15331,N_15073,N_15276);
and U15332 (N_15332,N_15104,N_15097);
nor U15333 (N_15333,N_15145,N_15016);
and U15334 (N_15334,N_15055,N_15212);
and U15335 (N_15335,N_15132,N_15000);
or U15336 (N_15336,N_15065,N_15273);
or U15337 (N_15337,N_15167,N_15007);
nand U15338 (N_15338,N_15126,N_15173);
xor U15339 (N_15339,N_15281,N_15176);
xnor U15340 (N_15340,N_15225,N_15027);
xnor U15341 (N_15341,N_15091,N_15083);
and U15342 (N_15342,N_15271,N_15060);
xnor U15343 (N_15343,N_15115,N_15218);
or U15344 (N_15344,N_15037,N_15069);
nor U15345 (N_15345,N_15088,N_15074);
nand U15346 (N_15346,N_15047,N_15135);
nor U15347 (N_15347,N_15295,N_15113);
and U15348 (N_15348,N_15233,N_15084);
and U15349 (N_15349,N_15274,N_15109);
nor U15350 (N_15350,N_15228,N_15067);
and U15351 (N_15351,N_15138,N_15114);
or U15352 (N_15352,N_15142,N_15100);
nand U15353 (N_15353,N_15052,N_15219);
or U15354 (N_15354,N_15133,N_15174);
and U15355 (N_15355,N_15044,N_15214);
or U15356 (N_15356,N_15201,N_15251);
nand U15357 (N_15357,N_15127,N_15048);
and U15358 (N_15358,N_15032,N_15194);
xor U15359 (N_15359,N_15033,N_15108);
nand U15360 (N_15360,N_15106,N_15170);
and U15361 (N_15361,N_15223,N_15227);
and U15362 (N_15362,N_15207,N_15200);
nor U15363 (N_15363,N_15211,N_15112);
xnor U15364 (N_15364,N_15096,N_15232);
and U15365 (N_15365,N_15062,N_15293);
and U15366 (N_15366,N_15163,N_15224);
and U15367 (N_15367,N_15291,N_15203);
nand U15368 (N_15368,N_15202,N_15238);
nand U15369 (N_15369,N_15257,N_15008);
xor U15370 (N_15370,N_15148,N_15024);
or U15371 (N_15371,N_15150,N_15264);
nor U15372 (N_15372,N_15255,N_15254);
or U15373 (N_15373,N_15018,N_15057);
nor U15374 (N_15374,N_15012,N_15154);
and U15375 (N_15375,N_15043,N_15181);
and U15376 (N_15376,N_15081,N_15050);
or U15377 (N_15377,N_15013,N_15149);
or U15378 (N_15378,N_15193,N_15247);
or U15379 (N_15379,N_15082,N_15152);
nand U15380 (N_15380,N_15262,N_15277);
nor U15381 (N_15381,N_15296,N_15244);
xnor U15382 (N_15382,N_15075,N_15051);
xnor U15383 (N_15383,N_15011,N_15169);
nor U15384 (N_15384,N_15182,N_15280);
or U15385 (N_15385,N_15220,N_15261);
or U15386 (N_15386,N_15235,N_15177);
xnor U15387 (N_15387,N_15282,N_15269);
nand U15388 (N_15388,N_15078,N_15162);
nor U15389 (N_15389,N_15186,N_15087);
and U15390 (N_15390,N_15153,N_15026);
nand U15391 (N_15391,N_15146,N_15021);
xor U15392 (N_15392,N_15038,N_15187);
and U15393 (N_15393,N_15105,N_15092);
xnor U15394 (N_15394,N_15001,N_15030);
and U15395 (N_15395,N_15164,N_15123);
xor U15396 (N_15396,N_15025,N_15198);
or U15397 (N_15397,N_15217,N_15110);
nor U15398 (N_15398,N_15134,N_15077);
nand U15399 (N_15399,N_15005,N_15172);
xor U15400 (N_15400,N_15095,N_15237);
or U15401 (N_15401,N_15229,N_15216);
nand U15402 (N_15402,N_15140,N_15129);
nand U15403 (N_15403,N_15256,N_15066);
nand U15404 (N_15404,N_15290,N_15272);
nor U15405 (N_15405,N_15288,N_15058);
and U15406 (N_15406,N_15215,N_15059);
or U15407 (N_15407,N_15158,N_15045);
nor U15408 (N_15408,N_15197,N_15143);
nand U15409 (N_15409,N_15089,N_15053);
xor U15410 (N_15410,N_15213,N_15068);
or U15411 (N_15411,N_15231,N_15230);
or U15412 (N_15412,N_15184,N_15260);
or U15413 (N_15413,N_15004,N_15161);
and U15414 (N_15414,N_15268,N_15297);
nand U15415 (N_15415,N_15160,N_15192);
nor U15416 (N_15416,N_15168,N_15147);
or U15417 (N_15417,N_15204,N_15285);
and U15418 (N_15418,N_15240,N_15283);
xor U15419 (N_15419,N_15111,N_15252);
nor U15420 (N_15420,N_15292,N_15125);
and U15421 (N_15421,N_15040,N_15278);
nand U15422 (N_15422,N_15002,N_15121);
xor U15423 (N_15423,N_15014,N_15259);
nand U15424 (N_15424,N_15137,N_15206);
or U15425 (N_15425,N_15275,N_15103);
nand U15426 (N_15426,N_15299,N_15245);
nor U15427 (N_15427,N_15178,N_15258);
xnor U15428 (N_15428,N_15226,N_15070);
nor U15429 (N_15429,N_15241,N_15248);
nor U15430 (N_15430,N_15099,N_15151);
and U15431 (N_15431,N_15234,N_15118);
and U15432 (N_15432,N_15221,N_15056);
nand U15433 (N_15433,N_15222,N_15188);
and U15434 (N_15434,N_15139,N_15294);
and U15435 (N_15435,N_15046,N_15205);
and U15436 (N_15436,N_15023,N_15270);
or U15437 (N_15437,N_15063,N_15010);
and U15438 (N_15438,N_15242,N_15022);
xor U15439 (N_15439,N_15006,N_15020);
and U15440 (N_15440,N_15171,N_15209);
or U15441 (N_15441,N_15189,N_15098);
and U15442 (N_15442,N_15086,N_15093);
nor U15443 (N_15443,N_15246,N_15287);
nor U15444 (N_15444,N_15156,N_15180);
nand U15445 (N_15445,N_15157,N_15119);
and U15446 (N_15446,N_15049,N_15265);
nor U15447 (N_15447,N_15284,N_15130);
xor U15448 (N_15448,N_15196,N_15116);
nand U15449 (N_15449,N_15102,N_15076);
xor U15450 (N_15450,N_15210,N_15254);
xnor U15451 (N_15451,N_15039,N_15041);
or U15452 (N_15452,N_15131,N_15265);
or U15453 (N_15453,N_15012,N_15028);
nor U15454 (N_15454,N_15048,N_15005);
xor U15455 (N_15455,N_15030,N_15033);
nand U15456 (N_15456,N_15045,N_15297);
xor U15457 (N_15457,N_15018,N_15035);
xnor U15458 (N_15458,N_15015,N_15127);
or U15459 (N_15459,N_15021,N_15048);
and U15460 (N_15460,N_15278,N_15185);
nor U15461 (N_15461,N_15030,N_15187);
or U15462 (N_15462,N_15002,N_15226);
or U15463 (N_15463,N_15107,N_15188);
nor U15464 (N_15464,N_15167,N_15120);
nor U15465 (N_15465,N_15110,N_15221);
and U15466 (N_15466,N_15192,N_15190);
nand U15467 (N_15467,N_15078,N_15099);
or U15468 (N_15468,N_15022,N_15281);
xnor U15469 (N_15469,N_15089,N_15259);
or U15470 (N_15470,N_15004,N_15231);
or U15471 (N_15471,N_15047,N_15161);
xor U15472 (N_15472,N_15043,N_15286);
or U15473 (N_15473,N_15044,N_15076);
or U15474 (N_15474,N_15250,N_15031);
or U15475 (N_15475,N_15155,N_15149);
nand U15476 (N_15476,N_15063,N_15058);
nand U15477 (N_15477,N_15105,N_15261);
and U15478 (N_15478,N_15139,N_15218);
or U15479 (N_15479,N_15138,N_15135);
and U15480 (N_15480,N_15069,N_15257);
xor U15481 (N_15481,N_15109,N_15272);
and U15482 (N_15482,N_15237,N_15274);
nand U15483 (N_15483,N_15197,N_15270);
nor U15484 (N_15484,N_15208,N_15068);
and U15485 (N_15485,N_15216,N_15249);
xor U15486 (N_15486,N_15151,N_15152);
nand U15487 (N_15487,N_15263,N_15254);
or U15488 (N_15488,N_15018,N_15009);
xnor U15489 (N_15489,N_15116,N_15243);
nor U15490 (N_15490,N_15072,N_15282);
nor U15491 (N_15491,N_15022,N_15006);
xor U15492 (N_15492,N_15095,N_15017);
and U15493 (N_15493,N_15281,N_15141);
nand U15494 (N_15494,N_15231,N_15217);
and U15495 (N_15495,N_15023,N_15192);
nand U15496 (N_15496,N_15111,N_15236);
and U15497 (N_15497,N_15157,N_15206);
and U15498 (N_15498,N_15168,N_15189);
and U15499 (N_15499,N_15042,N_15026);
xor U15500 (N_15500,N_15206,N_15152);
xnor U15501 (N_15501,N_15113,N_15048);
nand U15502 (N_15502,N_15079,N_15029);
nor U15503 (N_15503,N_15086,N_15053);
or U15504 (N_15504,N_15283,N_15161);
nor U15505 (N_15505,N_15057,N_15023);
xor U15506 (N_15506,N_15052,N_15062);
or U15507 (N_15507,N_15213,N_15270);
and U15508 (N_15508,N_15256,N_15059);
xnor U15509 (N_15509,N_15263,N_15159);
nor U15510 (N_15510,N_15020,N_15147);
nand U15511 (N_15511,N_15154,N_15168);
and U15512 (N_15512,N_15092,N_15154);
xor U15513 (N_15513,N_15132,N_15198);
nand U15514 (N_15514,N_15051,N_15111);
nor U15515 (N_15515,N_15116,N_15037);
or U15516 (N_15516,N_15007,N_15032);
xnor U15517 (N_15517,N_15287,N_15062);
nor U15518 (N_15518,N_15161,N_15060);
and U15519 (N_15519,N_15007,N_15048);
nor U15520 (N_15520,N_15027,N_15076);
nand U15521 (N_15521,N_15230,N_15269);
xnor U15522 (N_15522,N_15070,N_15243);
nor U15523 (N_15523,N_15073,N_15161);
xor U15524 (N_15524,N_15086,N_15028);
nand U15525 (N_15525,N_15265,N_15183);
xnor U15526 (N_15526,N_15085,N_15000);
and U15527 (N_15527,N_15211,N_15179);
or U15528 (N_15528,N_15269,N_15164);
xor U15529 (N_15529,N_15218,N_15184);
nor U15530 (N_15530,N_15299,N_15202);
nand U15531 (N_15531,N_15153,N_15223);
and U15532 (N_15532,N_15065,N_15240);
nand U15533 (N_15533,N_15222,N_15058);
nor U15534 (N_15534,N_15233,N_15049);
nor U15535 (N_15535,N_15131,N_15026);
or U15536 (N_15536,N_15080,N_15254);
xnor U15537 (N_15537,N_15084,N_15247);
or U15538 (N_15538,N_15250,N_15242);
and U15539 (N_15539,N_15222,N_15247);
xnor U15540 (N_15540,N_15288,N_15292);
xor U15541 (N_15541,N_15233,N_15114);
and U15542 (N_15542,N_15101,N_15253);
xor U15543 (N_15543,N_15103,N_15247);
nand U15544 (N_15544,N_15140,N_15210);
and U15545 (N_15545,N_15050,N_15007);
or U15546 (N_15546,N_15114,N_15053);
nor U15547 (N_15547,N_15278,N_15235);
or U15548 (N_15548,N_15078,N_15235);
nand U15549 (N_15549,N_15111,N_15141);
and U15550 (N_15550,N_15145,N_15210);
nor U15551 (N_15551,N_15226,N_15177);
or U15552 (N_15552,N_15265,N_15294);
or U15553 (N_15553,N_15116,N_15173);
or U15554 (N_15554,N_15181,N_15267);
xnor U15555 (N_15555,N_15260,N_15053);
xor U15556 (N_15556,N_15117,N_15012);
nand U15557 (N_15557,N_15185,N_15260);
nor U15558 (N_15558,N_15028,N_15048);
nor U15559 (N_15559,N_15292,N_15091);
nand U15560 (N_15560,N_15080,N_15275);
nor U15561 (N_15561,N_15247,N_15272);
nor U15562 (N_15562,N_15107,N_15094);
xor U15563 (N_15563,N_15005,N_15189);
xor U15564 (N_15564,N_15246,N_15095);
xnor U15565 (N_15565,N_15215,N_15000);
nand U15566 (N_15566,N_15181,N_15133);
or U15567 (N_15567,N_15169,N_15091);
nand U15568 (N_15568,N_15207,N_15007);
nand U15569 (N_15569,N_15224,N_15096);
or U15570 (N_15570,N_15171,N_15134);
xnor U15571 (N_15571,N_15024,N_15159);
nor U15572 (N_15572,N_15283,N_15291);
xor U15573 (N_15573,N_15286,N_15099);
and U15574 (N_15574,N_15157,N_15055);
and U15575 (N_15575,N_15250,N_15004);
xnor U15576 (N_15576,N_15119,N_15177);
nor U15577 (N_15577,N_15000,N_15109);
nand U15578 (N_15578,N_15143,N_15140);
nor U15579 (N_15579,N_15040,N_15145);
nand U15580 (N_15580,N_15084,N_15275);
or U15581 (N_15581,N_15190,N_15079);
nand U15582 (N_15582,N_15119,N_15220);
nor U15583 (N_15583,N_15147,N_15200);
nor U15584 (N_15584,N_15042,N_15220);
xor U15585 (N_15585,N_15083,N_15175);
or U15586 (N_15586,N_15259,N_15074);
nand U15587 (N_15587,N_15283,N_15222);
or U15588 (N_15588,N_15035,N_15126);
nor U15589 (N_15589,N_15296,N_15213);
nor U15590 (N_15590,N_15243,N_15277);
and U15591 (N_15591,N_15061,N_15038);
xor U15592 (N_15592,N_15113,N_15039);
or U15593 (N_15593,N_15008,N_15112);
and U15594 (N_15594,N_15274,N_15009);
nand U15595 (N_15595,N_15053,N_15240);
nand U15596 (N_15596,N_15094,N_15153);
nand U15597 (N_15597,N_15252,N_15198);
or U15598 (N_15598,N_15237,N_15201);
or U15599 (N_15599,N_15182,N_15183);
nor U15600 (N_15600,N_15569,N_15579);
nor U15601 (N_15601,N_15467,N_15494);
nor U15602 (N_15602,N_15301,N_15435);
nor U15603 (N_15603,N_15572,N_15482);
or U15604 (N_15604,N_15458,N_15401);
xor U15605 (N_15605,N_15397,N_15518);
or U15606 (N_15606,N_15527,N_15396);
and U15607 (N_15607,N_15588,N_15353);
or U15608 (N_15608,N_15461,N_15495);
nor U15609 (N_15609,N_15575,N_15547);
nand U15610 (N_15610,N_15381,N_15403);
or U15611 (N_15611,N_15311,N_15424);
nand U15612 (N_15612,N_15481,N_15453);
nand U15613 (N_15613,N_15374,N_15326);
nand U15614 (N_15614,N_15509,N_15593);
nand U15615 (N_15615,N_15418,N_15580);
and U15616 (N_15616,N_15306,N_15542);
nor U15617 (N_15617,N_15457,N_15552);
nor U15618 (N_15618,N_15412,N_15528);
nand U15619 (N_15619,N_15422,N_15357);
xnor U15620 (N_15620,N_15420,N_15426);
xnor U15621 (N_15621,N_15477,N_15516);
nor U15622 (N_15622,N_15555,N_15546);
and U15623 (N_15623,N_15567,N_15317);
or U15624 (N_15624,N_15525,N_15466);
or U15625 (N_15625,N_15339,N_15534);
nand U15626 (N_15626,N_15346,N_15394);
xnor U15627 (N_15627,N_15343,N_15596);
xor U15628 (N_15628,N_15562,N_15522);
and U15629 (N_15629,N_15468,N_15393);
xor U15630 (N_15630,N_15553,N_15554);
nand U15631 (N_15631,N_15587,N_15487);
xor U15632 (N_15632,N_15365,N_15450);
xnor U15633 (N_15633,N_15480,N_15406);
nor U15634 (N_15634,N_15307,N_15479);
nor U15635 (N_15635,N_15584,N_15402);
xnor U15636 (N_15636,N_15328,N_15550);
nand U15637 (N_15637,N_15590,N_15498);
nor U15638 (N_15638,N_15576,N_15310);
nor U15639 (N_15639,N_15473,N_15436);
or U15640 (N_15640,N_15463,N_15415);
nand U15641 (N_15641,N_15348,N_15521);
or U15642 (N_15642,N_15427,N_15517);
xnor U15643 (N_15643,N_15421,N_15452);
nor U15644 (N_15644,N_15434,N_15390);
xnor U15645 (N_15645,N_15488,N_15377);
nand U15646 (N_15646,N_15356,N_15548);
nand U15647 (N_15647,N_15563,N_15471);
and U15648 (N_15648,N_15583,N_15352);
xor U15649 (N_15649,N_15386,N_15591);
nor U15650 (N_15650,N_15568,N_15560);
nand U15651 (N_15651,N_15370,N_15520);
nor U15652 (N_15652,N_15313,N_15300);
and U15653 (N_15653,N_15573,N_15582);
nand U15654 (N_15654,N_15380,N_15383);
xnor U15655 (N_15655,N_15581,N_15375);
xor U15656 (N_15656,N_15388,N_15556);
xor U15657 (N_15657,N_15368,N_15442);
nor U15658 (N_15658,N_15496,N_15541);
and U15659 (N_15659,N_15334,N_15536);
nor U15660 (N_15660,N_15333,N_15492);
nor U15661 (N_15661,N_15410,N_15598);
or U15662 (N_15662,N_15533,N_15508);
and U15663 (N_15663,N_15366,N_15379);
xor U15664 (N_15664,N_15409,N_15369);
nand U15665 (N_15665,N_15391,N_15589);
nor U15666 (N_15666,N_15332,N_15344);
and U15667 (N_15667,N_15561,N_15537);
xnor U15668 (N_15668,N_15413,N_15465);
or U15669 (N_15669,N_15305,N_15511);
nand U15670 (N_15670,N_15507,N_15539);
or U15671 (N_15671,N_15423,N_15378);
and U15672 (N_15672,N_15526,N_15485);
and U15673 (N_15673,N_15557,N_15441);
and U15674 (N_15674,N_15430,N_15491);
nand U15675 (N_15675,N_15318,N_15549);
xor U15676 (N_15676,N_15571,N_15405);
xor U15677 (N_15677,N_15564,N_15519);
nand U15678 (N_15678,N_15322,N_15329);
and U15679 (N_15679,N_15565,N_15490);
nor U15680 (N_15680,N_15544,N_15364);
nand U15681 (N_15681,N_15444,N_15428);
xor U15682 (N_15682,N_15502,N_15543);
nor U15683 (N_15683,N_15531,N_15538);
or U15684 (N_15684,N_15345,N_15448);
or U15685 (N_15685,N_15327,N_15330);
or U15686 (N_15686,N_15392,N_15323);
nor U15687 (N_15687,N_15308,N_15304);
and U15688 (N_15688,N_15595,N_15398);
or U15689 (N_15689,N_15338,N_15462);
or U15690 (N_15690,N_15399,N_15505);
and U15691 (N_15691,N_15439,N_15407);
or U15692 (N_15692,N_15419,N_15446);
nor U15693 (N_15693,N_15512,N_15478);
and U15694 (N_15694,N_15417,N_15367);
or U15695 (N_15695,N_15451,N_15504);
or U15696 (N_15696,N_15578,N_15501);
xnor U15697 (N_15697,N_15577,N_15361);
xor U15698 (N_15698,N_15360,N_15325);
xnor U15699 (N_15699,N_15340,N_15470);
or U15700 (N_15700,N_15599,N_15592);
and U15701 (N_15701,N_15350,N_15513);
nor U15702 (N_15702,N_15351,N_15486);
or U15703 (N_15703,N_15408,N_15337);
nor U15704 (N_15704,N_15455,N_15319);
nor U15705 (N_15705,N_15474,N_15445);
xor U15706 (N_15706,N_15483,N_15371);
nand U15707 (N_15707,N_15497,N_15594);
nand U15708 (N_15708,N_15597,N_15535);
xnor U15709 (N_15709,N_15387,N_15532);
xnor U15710 (N_15710,N_15416,N_15384);
xnor U15711 (N_15711,N_15464,N_15449);
xor U15712 (N_15712,N_15341,N_15335);
and U15713 (N_15713,N_15551,N_15404);
nor U15714 (N_15714,N_15523,N_15358);
nand U15715 (N_15715,N_15315,N_15314);
xnor U15716 (N_15716,N_15302,N_15324);
nand U15717 (N_15717,N_15558,N_15429);
nand U15718 (N_15718,N_15506,N_15362);
nor U15719 (N_15719,N_15514,N_15529);
nand U15720 (N_15720,N_15359,N_15347);
nand U15721 (N_15721,N_15355,N_15440);
nand U15722 (N_15722,N_15376,N_15475);
and U15723 (N_15723,N_15570,N_15540);
and U15724 (N_15724,N_15443,N_15574);
and U15725 (N_15725,N_15385,N_15499);
nor U15726 (N_15726,N_15433,N_15545);
nand U15727 (N_15727,N_15476,N_15342);
and U15728 (N_15728,N_15456,N_15515);
or U15729 (N_15729,N_15363,N_15447);
nand U15730 (N_15730,N_15432,N_15316);
xor U15731 (N_15731,N_15493,N_15312);
or U15732 (N_15732,N_15321,N_15460);
or U15733 (N_15733,N_15431,N_15414);
and U15734 (N_15734,N_15389,N_15425);
or U15735 (N_15735,N_15303,N_15411);
or U15736 (N_15736,N_15459,N_15469);
nand U15737 (N_15737,N_15336,N_15510);
xnor U15738 (N_15738,N_15437,N_15354);
nand U15739 (N_15739,N_15503,N_15530);
nor U15740 (N_15740,N_15400,N_15320);
and U15741 (N_15741,N_15489,N_15309);
and U15742 (N_15742,N_15349,N_15331);
nor U15743 (N_15743,N_15585,N_15566);
and U15744 (N_15744,N_15454,N_15484);
and U15745 (N_15745,N_15373,N_15559);
xor U15746 (N_15746,N_15524,N_15472);
nand U15747 (N_15747,N_15500,N_15395);
xor U15748 (N_15748,N_15438,N_15372);
and U15749 (N_15749,N_15382,N_15586);
or U15750 (N_15750,N_15576,N_15457);
xnor U15751 (N_15751,N_15521,N_15485);
xnor U15752 (N_15752,N_15470,N_15362);
xnor U15753 (N_15753,N_15305,N_15442);
nor U15754 (N_15754,N_15353,N_15478);
nand U15755 (N_15755,N_15482,N_15422);
nand U15756 (N_15756,N_15419,N_15535);
and U15757 (N_15757,N_15357,N_15552);
and U15758 (N_15758,N_15467,N_15451);
xor U15759 (N_15759,N_15314,N_15514);
xnor U15760 (N_15760,N_15553,N_15333);
and U15761 (N_15761,N_15318,N_15507);
xnor U15762 (N_15762,N_15588,N_15342);
or U15763 (N_15763,N_15478,N_15565);
or U15764 (N_15764,N_15565,N_15510);
nand U15765 (N_15765,N_15562,N_15381);
nand U15766 (N_15766,N_15324,N_15443);
and U15767 (N_15767,N_15446,N_15399);
or U15768 (N_15768,N_15409,N_15361);
nand U15769 (N_15769,N_15515,N_15546);
nor U15770 (N_15770,N_15444,N_15370);
xnor U15771 (N_15771,N_15405,N_15543);
and U15772 (N_15772,N_15442,N_15498);
nor U15773 (N_15773,N_15440,N_15521);
or U15774 (N_15774,N_15382,N_15505);
or U15775 (N_15775,N_15436,N_15522);
or U15776 (N_15776,N_15585,N_15411);
nor U15777 (N_15777,N_15360,N_15571);
xnor U15778 (N_15778,N_15365,N_15327);
xor U15779 (N_15779,N_15434,N_15410);
nor U15780 (N_15780,N_15596,N_15348);
nor U15781 (N_15781,N_15557,N_15457);
nor U15782 (N_15782,N_15578,N_15473);
or U15783 (N_15783,N_15377,N_15556);
xor U15784 (N_15784,N_15303,N_15309);
or U15785 (N_15785,N_15473,N_15418);
or U15786 (N_15786,N_15489,N_15370);
nor U15787 (N_15787,N_15575,N_15445);
xor U15788 (N_15788,N_15392,N_15577);
or U15789 (N_15789,N_15438,N_15345);
and U15790 (N_15790,N_15315,N_15360);
nor U15791 (N_15791,N_15343,N_15459);
nand U15792 (N_15792,N_15435,N_15388);
or U15793 (N_15793,N_15349,N_15370);
nand U15794 (N_15794,N_15336,N_15332);
and U15795 (N_15795,N_15577,N_15555);
nor U15796 (N_15796,N_15426,N_15395);
nand U15797 (N_15797,N_15370,N_15388);
or U15798 (N_15798,N_15579,N_15383);
nand U15799 (N_15799,N_15304,N_15471);
nor U15800 (N_15800,N_15590,N_15565);
xor U15801 (N_15801,N_15589,N_15552);
nor U15802 (N_15802,N_15558,N_15427);
xnor U15803 (N_15803,N_15366,N_15308);
nor U15804 (N_15804,N_15365,N_15466);
nor U15805 (N_15805,N_15475,N_15565);
xor U15806 (N_15806,N_15486,N_15429);
and U15807 (N_15807,N_15423,N_15409);
xor U15808 (N_15808,N_15324,N_15488);
or U15809 (N_15809,N_15498,N_15515);
or U15810 (N_15810,N_15316,N_15349);
and U15811 (N_15811,N_15393,N_15535);
nor U15812 (N_15812,N_15594,N_15499);
and U15813 (N_15813,N_15498,N_15356);
xnor U15814 (N_15814,N_15546,N_15472);
or U15815 (N_15815,N_15406,N_15357);
or U15816 (N_15816,N_15350,N_15500);
xor U15817 (N_15817,N_15582,N_15399);
and U15818 (N_15818,N_15349,N_15438);
and U15819 (N_15819,N_15492,N_15363);
xnor U15820 (N_15820,N_15319,N_15348);
nor U15821 (N_15821,N_15463,N_15434);
nand U15822 (N_15822,N_15569,N_15474);
or U15823 (N_15823,N_15565,N_15498);
or U15824 (N_15824,N_15431,N_15313);
or U15825 (N_15825,N_15326,N_15452);
nand U15826 (N_15826,N_15431,N_15401);
nor U15827 (N_15827,N_15417,N_15344);
nand U15828 (N_15828,N_15503,N_15567);
xor U15829 (N_15829,N_15310,N_15422);
and U15830 (N_15830,N_15467,N_15310);
or U15831 (N_15831,N_15424,N_15352);
or U15832 (N_15832,N_15368,N_15322);
and U15833 (N_15833,N_15451,N_15365);
or U15834 (N_15834,N_15593,N_15438);
nor U15835 (N_15835,N_15423,N_15306);
and U15836 (N_15836,N_15455,N_15398);
xnor U15837 (N_15837,N_15424,N_15324);
xor U15838 (N_15838,N_15581,N_15317);
nor U15839 (N_15839,N_15515,N_15342);
and U15840 (N_15840,N_15315,N_15477);
and U15841 (N_15841,N_15337,N_15431);
nor U15842 (N_15842,N_15570,N_15529);
nand U15843 (N_15843,N_15507,N_15365);
xor U15844 (N_15844,N_15316,N_15407);
xor U15845 (N_15845,N_15475,N_15351);
xnor U15846 (N_15846,N_15539,N_15595);
nor U15847 (N_15847,N_15305,N_15435);
xnor U15848 (N_15848,N_15414,N_15590);
nand U15849 (N_15849,N_15310,N_15394);
and U15850 (N_15850,N_15561,N_15574);
and U15851 (N_15851,N_15433,N_15342);
nand U15852 (N_15852,N_15351,N_15309);
xnor U15853 (N_15853,N_15432,N_15539);
nor U15854 (N_15854,N_15442,N_15323);
and U15855 (N_15855,N_15448,N_15471);
and U15856 (N_15856,N_15432,N_15441);
and U15857 (N_15857,N_15450,N_15323);
nand U15858 (N_15858,N_15594,N_15526);
xor U15859 (N_15859,N_15463,N_15353);
nand U15860 (N_15860,N_15413,N_15520);
or U15861 (N_15861,N_15598,N_15358);
nand U15862 (N_15862,N_15541,N_15310);
or U15863 (N_15863,N_15496,N_15507);
xnor U15864 (N_15864,N_15435,N_15500);
xor U15865 (N_15865,N_15432,N_15322);
xnor U15866 (N_15866,N_15570,N_15310);
nor U15867 (N_15867,N_15389,N_15465);
and U15868 (N_15868,N_15556,N_15552);
xor U15869 (N_15869,N_15584,N_15378);
and U15870 (N_15870,N_15523,N_15316);
nand U15871 (N_15871,N_15316,N_15340);
nor U15872 (N_15872,N_15301,N_15371);
nor U15873 (N_15873,N_15551,N_15538);
xnor U15874 (N_15874,N_15369,N_15331);
nand U15875 (N_15875,N_15536,N_15441);
and U15876 (N_15876,N_15535,N_15340);
xnor U15877 (N_15877,N_15415,N_15561);
nand U15878 (N_15878,N_15519,N_15513);
xor U15879 (N_15879,N_15570,N_15500);
xor U15880 (N_15880,N_15468,N_15428);
or U15881 (N_15881,N_15581,N_15599);
nor U15882 (N_15882,N_15569,N_15344);
xor U15883 (N_15883,N_15501,N_15476);
nor U15884 (N_15884,N_15329,N_15545);
and U15885 (N_15885,N_15423,N_15560);
nor U15886 (N_15886,N_15506,N_15375);
xnor U15887 (N_15887,N_15447,N_15531);
and U15888 (N_15888,N_15574,N_15501);
xnor U15889 (N_15889,N_15359,N_15309);
or U15890 (N_15890,N_15508,N_15594);
and U15891 (N_15891,N_15352,N_15460);
and U15892 (N_15892,N_15361,N_15436);
and U15893 (N_15893,N_15416,N_15395);
and U15894 (N_15894,N_15556,N_15372);
or U15895 (N_15895,N_15596,N_15530);
and U15896 (N_15896,N_15539,N_15429);
nor U15897 (N_15897,N_15305,N_15570);
nand U15898 (N_15898,N_15475,N_15495);
nor U15899 (N_15899,N_15346,N_15402);
xnor U15900 (N_15900,N_15700,N_15768);
or U15901 (N_15901,N_15631,N_15669);
and U15902 (N_15902,N_15894,N_15743);
and U15903 (N_15903,N_15750,N_15708);
and U15904 (N_15904,N_15694,N_15718);
or U15905 (N_15905,N_15836,N_15723);
and U15906 (N_15906,N_15872,N_15736);
nor U15907 (N_15907,N_15727,N_15706);
xor U15908 (N_15908,N_15739,N_15603);
nor U15909 (N_15909,N_15600,N_15650);
nor U15910 (N_15910,N_15887,N_15849);
xnor U15911 (N_15911,N_15666,N_15711);
xor U15912 (N_15912,N_15730,N_15678);
or U15913 (N_15913,N_15688,N_15837);
xnor U15914 (N_15914,N_15653,N_15876);
nand U15915 (N_15915,N_15851,N_15838);
or U15916 (N_15916,N_15726,N_15693);
xnor U15917 (N_15917,N_15841,N_15873);
nor U15918 (N_15918,N_15659,N_15828);
or U15919 (N_15919,N_15883,N_15702);
and U15920 (N_15920,N_15681,N_15614);
xor U15921 (N_15921,N_15623,N_15608);
nand U15922 (N_15922,N_15673,N_15691);
xnor U15923 (N_15923,N_15618,N_15648);
or U15924 (N_15924,N_15755,N_15870);
or U15925 (N_15925,N_15840,N_15884);
or U15926 (N_15926,N_15630,N_15867);
xor U15927 (N_15927,N_15756,N_15674);
or U15928 (N_15928,N_15764,N_15896);
or U15929 (N_15929,N_15612,N_15720);
or U15930 (N_15930,N_15763,N_15661);
or U15931 (N_15931,N_15626,N_15619);
xnor U15932 (N_15932,N_15759,N_15856);
or U15933 (N_15933,N_15857,N_15719);
nor U15934 (N_15934,N_15819,N_15733);
nor U15935 (N_15935,N_15793,N_15663);
xor U15936 (N_15936,N_15609,N_15795);
nor U15937 (N_15937,N_15656,N_15810);
nor U15938 (N_15938,N_15751,N_15649);
nor U15939 (N_15939,N_15664,N_15748);
nand U15940 (N_15940,N_15826,N_15728);
and U15941 (N_15941,N_15604,N_15622);
xnor U15942 (N_15942,N_15680,N_15738);
xor U15943 (N_15943,N_15697,N_15746);
xor U15944 (N_15944,N_15880,N_15742);
xnor U15945 (N_15945,N_15846,N_15804);
xor U15946 (N_15946,N_15807,N_15606);
nor U15947 (N_15947,N_15620,N_15744);
nor U15948 (N_15948,N_15615,N_15842);
or U15949 (N_15949,N_15658,N_15682);
nand U15950 (N_15950,N_15652,N_15777);
nor U15951 (N_15951,N_15646,N_15799);
nand U15952 (N_15952,N_15601,N_15879);
nor U15953 (N_15953,N_15639,N_15897);
xnor U15954 (N_15954,N_15893,N_15845);
nand U15955 (N_15955,N_15721,N_15613);
or U15956 (N_15956,N_15634,N_15758);
or U15957 (N_15957,N_15797,N_15647);
xnor U15958 (N_15958,N_15813,N_15766);
nor U15959 (N_15959,N_15687,N_15621);
nand U15960 (N_15960,N_15778,N_15817);
or U15961 (N_15961,N_15789,N_15761);
and U15962 (N_15962,N_15705,N_15627);
or U15963 (N_15963,N_15839,N_15651);
xnor U15964 (N_15964,N_15850,N_15660);
and U15965 (N_15965,N_15689,N_15692);
nand U15966 (N_15966,N_15859,N_15735);
nand U15967 (N_15967,N_15668,N_15820);
nand U15968 (N_15968,N_15786,N_15628);
nor U15969 (N_15969,N_15769,N_15731);
nor U15970 (N_15970,N_15854,N_15881);
or U15971 (N_15971,N_15869,N_15865);
and U15972 (N_15972,N_15787,N_15670);
nor U15973 (N_15973,N_15875,N_15716);
nor U15974 (N_15974,N_15864,N_15878);
nor U15975 (N_15975,N_15809,N_15712);
and U15976 (N_15976,N_15632,N_15794);
nor U15977 (N_15977,N_15625,N_15683);
and U15978 (N_15978,N_15657,N_15675);
xor U15979 (N_15979,N_15827,N_15832);
or U15980 (N_15980,N_15862,N_15677);
and U15981 (N_15981,N_15860,N_15815);
or U15982 (N_15982,N_15796,N_15757);
and U15983 (N_15983,N_15818,N_15800);
nand U15984 (N_15984,N_15734,N_15822);
and U15985 (N_15985,N_15858,N_15747);
xor U15986 (N_15986,N_15753,N_15847);
nor U15987 (N_15987,N_15774,N_15785);
nor U15988 (N_15988,N_15624,N_15830);
nand U15989 (N_15989,N_15607,N_15776);
or U15990 (N_15990,N_15821,N_15835);
or U15991 (N_15991,N_15729,N_15672);
nor U15992 (N_15992,N_15767,N_15722);
nand U15993 (N_15993,N_15791,N_15707);
nor U15994 (N_15994,N_15781,N_15635);
nand U15995 (N_15995,N_15814,N_15792);
nand U15996 (N_15996,N_15641,N_15855);
nand U15997 (N_15997,N_15803,N_15829);
nor U15998 (N_15998,N_15802,N_15638);
xnor U15999 (N_15999,N_15642,N_15874);
or U16000 (N_16000,N_15843,N_15699);
xnor U16001 (N_16001,N_15765,N_15833);
nor U16002 (N_16002,N_15741,N_15770);
nand U16003 (N_16003,N_15886,N_15644);
and U16004 (N_16004,N_15898,N_15782);
nand U16005 (N_16005,N_15715,N_15732);
nor U16006 (N_16006,N_15788,N_15816);
nand U16007 (N_16007,N_15637,N_15724);
and U16008 (N_16008,N_15899,N_15801);
nor U16009 (N_16009,N_15667,N_15824);
or U16010 (N_16010,N_15654,N_15698);
or U16011 (N_16011,N_15779,N_15611);
or U16012 (N_16012,N_15617,N_15780);
xor U16013 (N_16013,N_15868,N_15892);
and U16014 (N_16014,N_15848,N_15725);
xnor U16015 (N_16015,N_15629,N_15752);
or U16016 (N_16016,N_15740,N_15633);
nor U16017 (N_16017,N_15852,N_15790);
nand U16018 (N_16018,N_15772,N_15710);
xnor U16019 (N_16019,N_15605,N_15831);
or U16020 (N_16020,N_15640,N_15844);
nor U16021 (N_16021,N_15762,N_15891);
nor U16022 (N_16022,N_15737,N_15895);
and U16023 (N_16023,N_15671,N_15783);
or U16024 (N_16024,N_15889,N_15695);
or U16025 (N_16025,N_15811,N_15871);
nand U16026 (N_16026,N_15771,N_15636);
xnor U16027 (N_16027,N_15704,N_15806);
or U16028 (N_16028,N_15754,N_15882);
or U16029 (N_16029,N_15890,N_15676);
nand U16030 (N_16030,N_15866,N_15662);
nand U16031 (N_16031,N_15834,N_15665);
and U16032 (N_16032,N_15690,N_15616);
xnor U16033 (N_16033,N_15713,N_15610);
and U16034 (N_16034,N_15696,N_15602);
and U16035 (N_16035,N_15645,N_15825);
xor U16036 (N_16036,N_15686,N_15853);
and U16037 (N_16037,N_15812,N_15745);
and U16038 (N_16038,N_15709,N_15798);
nand U16039 (N_16039,N_15701,N_15877);
xnor U16040 (N_16040,N_15888,N_15808);
xnor U16041 (N_16041,N_15823,N_15643);
or U16042 (N_16042,N_15773,N_15805);
or U16043 (N_16043,N_15863,N_15885);
and U16044 (N_16044,N_15684,N_15861);
xnor U16045 (N_16045,N_15679,N_15655);
nand U16046 (N_16046,N_15760,N_15784);
nand U16047 (N_16047,N_15714,N_15685);
or U16048 (N_16048,N_15703,N_15749);
and U16049 (N_16049,N_15717,N_15775);
or U16050 (N_16050,N_15842,N_15811);
xor U16051 (N_16051,N_15871,N_15703);
and U16052 (N_16052,N_15824,N_15863);
nor U16053 (N_16053,N_15678,N_15875);
or U16054 (N_16054,N_15694,N_15715);
and U16055 (N_16055,N_15601,N_15763);
and U16056 (N_16056,N_15654,N_15716);
xnor U16057 (N_16057,N_15869,N_15746);
xor U16058 (N_16058,N_15732,N_15777);
nor U16059 (N_16059,N_15774,N_15719);
or U16060 (N_16060,N_15812,N_15786);
or U16061 (N_16061,N_15879,N_15854);
or U16062 (N_16062,N_15770,N_15815);
or U16063 (N_16063,N_15778,N_15812);
or U16064 (N_16064,N_15774,N_15859);
nand U16065 (N_16065,N_15796,N_15828);
or U16066 (N_16066,N_15763,N_15773);
nand U16067 (N_16067,N_15751,N_15801);
xnor U16068 (N_16068,N_15616,N_15808);
nor U16069 (N_16069,N_15725,N_15724);
or U16070 (N_16070,N_15688,N_15779);
nand U16071 (N_16071,N_15762,N_15864);
xnor U16072 (N_16072,N_15614,N_15781);
nor U16073 (N_16073,N_15812,N_15829);
and U16074 (N_16074,N_15648,N_15660);
nor U16075 (N_16075,N_15749,N_15684);
nor U16076 (N_16076,N_15807,N_15605);
or U16077 (N_16077,N_15630,N_15797);
or U16078 (N_16078,N_15707,N_15660);
nor U16079 (N_16079,N_15648,N_15873);
and U16080 (N_16080,N_15884,N_15835);
or U16081 (N_16081,N_15754,N_15707);
or U16082 (N_16082,N_15617,N_15770);
and U16083 (N_16083,N_15893,N_15638);
or U16084 (N_16084,N_15631,N_15867);
xor U16085 (N_16085,N_15799,N_15833);
nor U16086 (N_16086,N_15894,N_15661);
xor U16087 (N_16087,N_15802,N_15762);
nand U16088 (N_16088,N_15611,N_15606);
nand U16089 (N_16089,N_15892,N_15790);
nor U16090 (N_16090,N_15739,N_15758);
nand U16091 (N_16091,N_15802,N_15749);
nor U16092 (N_16092,N_15889,N_15753);
or U16093 (N_16093,N_15745,N_15824);
and U16094 (N_16094,N_15887,N_15821);
or U16095 (N_16095,N_15689,N_15632);
nand U16096 (N_16096,N_15845,N_15693);
nor U16097 (N_16097,N_15705,N_15885);
and U16098 (N_16098,N_15843,N_15765);
nand U16099 (N_16099,N_15862,N_15678);
nand U16100 (N_16100,N_15765,N_15880);
xor U16101 (N_16101,N_15847,N_15781);
and U16102 (N_16102,N_15685,N_15755);
and U16103 (N_16103,N_15789,N_15687);
nand U16104 (N_16104,N_15660,N_15733);
xor U16105 (N_16105,N_15749,N_15668);
nor U16106 (N_16106,N_15662,N_15844);
and U16107 (N_16107,N_15796,N_15736);
nor U16108 (N_16108,N_15808,N_15846);
nor U16109 (N_16109,N_15677,N_15777);
nor U16110 (N_16110,N_15768,N_15662);
nor U16111 (N_16111,N_15632,N_15873);
nand U16112 (N_16112,N_15885,N_15804);
or U16113 (N_16113,N_15846,N_15889);
nor U16114 (N_16114,N_15828,N_15898);
and U16115 (N_16115,N_15827,N_15792);
or U16116 (N_16116,N_15719,N_15733);
xor U16117 (N_16117,N_15785,N_15700);
nand U16118 (N_16118,N_15625,N_15790);
or U16119 (N_16119,N_15652,N_15647);
nand U16120 (N_16120,N_15689,N_15793);
xor U16121 (N_16121,N_15703,N_15714);
xor U16122 (N_16122,N_15794,N_15761);
and U16123 (N_16123,N_15688,N_15842);
or U16124 (N_16124,N_15798,N_15892);
xnor U16125 (N_16125,N_15827,N_15760);
and U16126 (N_16126,N_15652,N_15616);
and U16127 (N_16127,N_15819,N_15864);
or U16128 (N_16128,N_15669,N_15678);
or U16129 (N_16129,N_15800,N_15712);
nand U16130 (N_16130,N_15669,N_15664);
xor U16131 (N_16131,N_15722,N_15852);
xnor U16132 (N_16132,N_15807,N_15619);
xnor U16133 (N_16133,N_15827,N_15830);
nor U16134 (N_16134,N_15700,N_15777);
xor U16135 (N_16135,N_15606,N_15740);
xnor U16136 (N_16136,N_15762,N_15875);
or U16137 (N_16137,N_15693,N_15616);
or U16138 (N_16138,N_15622,N_15634);
nor U16139 (N_16139,N_15880,N_15796);
and U16140 (N_16140,N_15692,N_15850);
nand U16141 (N_16141,N_15788,N_15611);
or U16142 (N_16142,N_15736,N_15619);
xnor U16143 (N_16143,N_15751,N_15806);
or U16144 (N_16144,N_15880,N_15843);
or U16145 (N_16145,N_15615,N_15711);
and U16146 (N_16146,N_15814,N_15673);
nand U16147 (N_16147,N_15662,N_15716);
and U16148 (N_16148,N_15814,N_15820);
nand U16149 (N_16149,N_15821,N_15816);
nand U16150 (N_16150,N_15856,N_15709);
nor U16151 (N_16151,N_15706,N_15717);
or U16152 (N_16152,N_15662,N_15719);
or U16153 (N_16153,N_15681,N_15641);
or U16154 (N_16154,N_15716,N_15819);
or U16155 (N_16155,N_15624,N_15813);
nor U16156 (N_16156,N_15689,N_15773);
or U16157 (N_16157,N_15862,N_15743);
xnor U16158 (N_16158,N_15702,N_15845);
or U16159 (N_16159,N_15651,N_15836);
nand U16160 (N_16160,N_15681,N_15637);
nand U16161 (N_16161,N_15719,N_15819);
and U16162 (N_16162,N_15651,N_15875);
or U16163 (N_16163,N_15688,N_15776);
nor U16164 (N_16164,N_15805,N_15896);
or U16165 (N_16165,N_15698,N_15668);
and U16166 (N_16166,N_15700,N_15767);
nand U16167 (N_16167,N_15694,N_15753);
nand U16168 (N_16168,N_15782,N_15716);
or U16169 (N_16169,N_15817,N_15656);
xor U16170 (N_16170,N_15623,N_15856);
and U16171 (N_16171,N_15848,N_15603);
xnor U16172 (N_16172,N_15724,N_15606);
and U16173 (N_16173,N_15741,N_15795);
xor U16174 (N_16174,N_15628,N_15673);
and U16175 (N_16175,N_15614,N_15692);
and U16176 (N_16176,N_15810,N_15883);
nor U16177 (N_16177,N_15828,N_15811);
nor U16178 (N_16178,N_15624,N_15723);
or U16179 (N_16179,N_15745,N_15622);
nand U16180 (N_16180,N_15770,N_15851);
nor U16181 (N_16181,N_15647,N_15622);
and U16182 (N_16182,N_15607,N_15665);
and U16183 (N_16183,N_15888,N_15681);
and U16184 (N_16184,N_15783,N_15613);
nor U16185 (N_16185,N_15785,N_15729);
xnor U16186 (N_16186,N_15849,N_15716);
or U16187 (N_16187,N_15771,N_15830);
or U16188 (N_16188,N_15843,N_15783);
and U16189 (N_16189,N_15632,N_15765);
nor U16190 (N_16190,N_15631,N_15858);
nand U16191 (N_16191,N_15647,N_15896);
xnor U16192 (N_16192,N_15787,N_15851);
nand U16193 (N_16193,N_15653,N_15757);
nand U16194 (N_16194,N_15873,N_15870);
xnor U16195 (N_16195,N_15646,N_15872);
xnor U16196 (N_16196,N_15877,N_15757);
xnor U16197 (N_16197,N_15723,N_15784);
and U16198 (N_16198,N_15614,N_15773);
xor U16199 (N_16199,N_15676,N_15871);
or U16200 (N_16200,N_15923,N_16013);
nand U16201 (N_16201,N_16128,N_16024);
nor U16202 (N_16202,N_16188,N_16050);
or U16203 (N_16203,N_16149,N_16021);
xor U16204 (N_16204,N_16085,N_16140);
xnor U16205 (N_16205,N_16196,N_16168);
nand U16206 (N_16206,N_16062,N_16080);
and U16207 (N_16207,N_16078,N_16175);
nor U16208 (N_16208,N_15960,N_15922);
and U16209 (N_16209,N_16167,N_15964);
nor U16210 (N_16210,N_16158,N_16197);
and U16211 (N_16211,N_16042,N_15944);
nand U16212 (N_16212,N_16090,N_15970);
nand U16213 (N_16213,N_16046,N_15908);
or U16214 (N_16214,N_16100,N_15939);
nand U16215 (N_16215,N_15951,N_15974);
and U16216 (N_16216,N_16191,N_16132);
or U16217 (N_16217,N_16065,N_16082);
nor U16218 (N_16218,N_15940,N_16043);
and U16219 (N_16219,N_16162,N_15926);
xnor U16220 (N_16220,N_16155,N_15965);
nand U16221 (N_16221,N_16157,N_16159);
and U16222 (N_16222,N_16186,N_16031);
nor U16223 (N_16223,N_15972,N_16007);
nor U16224 (N_16224,N_16160,N_15904);
xor U16225 (N_16225,N_16093,N_16161);
xnor U16226 (N_16226,N_16067,N_16106);
nor U16227 (N_16227,N_16037,N_16070);
and U16228 (N_16228,N_15935,N_16135);
nand U16229 (N_16229,N_16185,N_16011);
and U16230 (N_16230,N_16116,N_15907);
nor U16231 (N_16231,N_16111,N_15979);
nor U16232 (N_16232,N_16115,N_16079);
nor U16233 (N_16233,N_15941,N_15994);
and U16234 (N_16234,N_16017,N_15906);
nor U16235 (N_16235,N_16027,N_16130);
nand U16236 (N_16236,N_16099,N_16059);
or U16237 (N_16237,N_16156,N_16077);
xnor U16238 (N_16238,N_16081,N_16127);
nor U16239 (N_16239,N_16174,N_16124);
and U16240 (N_16240,N_15966,N_16183);
or U16241 (N_16241,N_16152,N_15985);
and U16242 (N_16242,N_15955,N_16146);
xor U16243 (N_16243,N_15961,N_16038);
or U16244 (N_16244,N_16066,N_15957);
and U16245 (N_16245,N_15924,N_15902);
and U16246 (N_16246,N_15933,N_16154);
xnor U16247 (N_16247,N_16000,N_16045);
xor U16248 (N_16248,N_16069,N_15947);
xnor U16249 (N_16249,N_16060,N_16129);
nor U16250 (N_16250,N_16098,N_16008);
nand U16251 (N_16251,N_15949,N_16187);
and U16252 (N_16252,N_16112,N_15910);
nand U16253 (N_16253,N_16144,N_16118);
and U16254 (N_16254,N_16189,N_16051);
and U16255 (N_16255,N_15946,N_15976);
xnor U16256 (N_16256,N_16166,N_16108);
xnor U16257 (N_16257,N_16094,N_16004);
xor U16258 (N_16258,N_16015,N_16063);
or U16259 (N_16259,N_15988,N_16018);
xnor U16260 (N_16260,N_16057,N_15920);
nand U16261 (N_16261,N_15929,N_16176);
and U16262 (N_16262,N_16073,N_16142);
nand U16263 (N_16263,N_15932,N_16180);
or U16264 (N_16264,N_16109,N_15975);
nor U16265 (N_16265,N_16091,N_15945);
and U16266 (N_16266,N_16055,N_15905);
or U16267 (N_16267,N_16030,N_16138);
nand U16268 (N_16268,N_16010,N_16048);
xnor U16269 (N_16269,N_16170,N_16103);
nand U16270 (N_16270,N_16019,N_16095);
nor U16271 (N_16271,N_15977,N_16029);
xor U16272 (N_16272,N_15934,N_15989);
or U16273 (N_16273,N_16104,N_15900);
nand U16274 (N_16274,N_16044,N_16033);
and U16275 (N_16275,N_15915,N_16068);
nand U16276 (N_16276,N_15986,N_16151);
xnor U16277 (N_16277,N_15981,N_15918);
nand U16278 (N_16278,N_15948,N_15925);
nor U16279 (N_16279,N_16088,N_15928);
nor U16280 (N_16280,N_16198,N_16139);
nand U16281 (N_16281,N_16125,N_16102);
or U16282 (N_16282,N_16133,N_16034);
nand U16283 (N_16283,N_16150,N_16052);
nor U16284 (N_16284,N_15942,N_15987);
nor U16285 (N_16285,N_16041,N_16113);
nor U16286 (N_16286,N_16194,N_16074);
xnor U16287 (N_16287,N_16025,N_15903);
and U16288 (N_16288,N_15962,N_16054);
nor U16289 (N_16289,N_16092,N_16097);
xnor U16290 (N_16290,N_16119,N_15997);
or U16291 (N_16291,N_16153,N_16178);
xnor U16292 (N_16292,N_16141,N_16026);
and U16293 (N_16293,N_16002,N_16136);
and U16294 (N_16294,N_15911,N_16028);
nor U16295 (N_16295,N_16076,N_16184);
nor U16296 (N_16296,N_15950,N_16056);
xnor U16297 (N_16297,N_15992,N_15952);
and U16298 (N_16298,N_15999,N_16173);
or U16299 (N_16299,N_15901,N_16134);
nand U16300 (N_16300,N_16172,N_16163);
and U16301 (N_16301,N_16107,N_16053);
xnor U16302 (N_16302,N_16199,N_15991);
xor U16303 (N_16303,N_16023,N_15938);
nand U16304 (N_16304,N_16039,N_16071);
and U16305 (N_16305,N_15984,N_16001);
or U16306 (N_16306,N_16084,N_16164);
nand U16307 (N_16307,N_16145,N_15930);
nor U16308 (N_16308,N_16020,N_16192);
or U16309 (N_16309,N_16101,N_16003);
xnor U16310 (N_16310,N_16169,N_16012);
xnor U16311 (N_16311,N_16032,N_16058);
nor U16312 (N_16312,N_16123,N_15912);
nor U16313 (N_16313,N_15913,N_15956);
nor U16314 (N_16314,N_16117,N_15963);
and U16315 (N_16315,N_16096,N_16120);
nand U16316 (N_16316,N_16126,N_16009);
or U16317 (N_16317,N_15959,N_16121);
or U16318 (N_16318,N_15971,N_16089);
and U16319 (N_16319,N_15998,N_16110);
or U16320 (N_16320,N_15967,N_15995);
or U16321 (N_16321,N_15943,N_16143);
nand U16322 (N_16322,N_16165,N_16105);
xor U16323 (N_16323,N_15931,N_16040);
nor U16324 (N_16324,N_16122,N_16064);
and U16325 (N_16325,N_16087,N_16179);
or U16326 (N_16326,N_15953,N_15993);
and U16327 (N_16327,N_16182,N_16014);
and U16328 (N_16328,N_16016,N_15973);
and U16329 (N_16329,N_15983,N_16190);
or U16330 (N_16330,N_15927,N_16083);
xnor U16331 (N_16331,N_16148,N_15980);
nand U16332 (N_16332,N_16047,N_15909);
xor U16333 (N_16333,N_15914,N_15937);
and U16334 (N_16334,N_15968,N_15921);
nand U16335 (N_16335,N_16006,N_16195);
nand U16336 (N_16336,N_15916,N_15990);
xnor U16337 (N_16337,N_16147,N_16061);
xor U16338 (N_16338,N_15969,N_16075);
nand U16339 (N_16339,N_16072,N_15936);
nand U16340 (N_16340,N_16049,N_15996);
xnor U16341 (N_16341,N_16171,N_16086);
nor U16342 (N_16342,N_16035,N_16137);
nand U16343 (N_16343,N_15954,N_15982);
and U16344 (N_16344,N_16114,N_16131);
xor U16345 (N_16345,N_15958,N_16193);
and U16346 (N_16346,N_15919,N_16036);
and U16347 (N_16347,N_15917,N_16181);
nand U16348 (N_16348,N_16022,N_16005);
and U16349 (N_16349,N_16177,N_15978);
and U16350 (N_16350,N_15962,N_15982);
nor U16351 (N_16351,N_15920,N_16139);
and U16352 (N_16352,N_16126,N_16138);
and U16353 (N_16353,N_15953,N_15970);
xnor U16354 (N_16354,N_16024,N_15985);
nand U16355 (N_16355,N_16147,N_15908);
nor U16356 (N_16356,N_16077,N_16098);
nor U16357 (N_16357,N_16089,N_16167);
or U16358 (N_16358,N_16051,N_15904);
or U16359 (N_16359,N_16113,N_16150);
nand U16360 (N_16360,N_16094,N_16129);
nand U16361 (N_16361,N_15907,N_16053);
or U16362 (N_16362,N_15954,N_15974);
nor U16363 (N_16363,N_15979,N_16150);
and U16364 (N_16364,N_16053,N_16064);
nor U16365 (N_16365,N_15970,N_15979);
and U16366 (N_16366,N_15998,N_16101);
nor U16367 (N_16367,N_16122,N_16168);
nor U16368 (N_16368,N_16176,N_15945);
nand U16369 (N_16369,N_16166,N_16117);
and U16370 (N_16370,N_16170,N_16027);
nand U16371 (N_16371,N_16199,N_16058);
and U16372 (N_16372,N_16080,N_15918);
or U16373 (N_16373,N_16156,N_15996);
xor U16374 (N_16374,N_16197,N_16127);
or U16375 (N_16375,N_16116,N_16170);
or U16376 (N_16376,N_15916,N_15939);
and U16377 (N_16377,N_15955,N_16114);
or U16378 (N_16378,N_16170,N_15997);
or U16379 (N_16379,N_16003,N_16166);
xnor U16380 (N_16380,N_16040,N_16038);
or U16381 (N_16381,N_16085,N_16027);
nor U16382 (N_16382,N_16144,N_15916);
or U16383 (N_16383,N_15901,N_16142);
or U16384 (N_16384,N_16171,N_16124);
nor U16385 (N_16385,N_16109,N_16167);
and U16386 (N_16386,N_15960,N_15984);
and U16387 (N_16387,N_15900,N_16032);
and U16388 (N_16388,N_16179,N_15926);
nor U16389 (N_16389,N_15953,N_15987);
nand U16390 (N_16390,N_15922,N_16072);
or U16391 (N_16391,N_16015,N_15905);
and U16392 (N_16392,N_15971,N_16062);
and U16393 (N_16393,N_15977,N_15910);
xnor U16394 (N_16394,N_16090,N_16072);
or U16395 (N_16395,N_16000,N_16047);
or U16396 (N_16396,N_16161,N_16010);
xnor U16397 (N_16397,N_15926,N_16126);
and U16398 (N_16398,N_15978,N_16011);
or U16399 (N_16399,N_15944,N_16054);
or U16400 (N_16400,N_16050,N_16061);
and U16401 (N_16401,N_16106,N_16024);
nor U16402 (N_16402,N_15949,N_15937);
nand U16403 (N_16403,N_16122,N_15903);
nand U16404 (N_16404,N_16076,N_16125);
nand U16405 (N_16405,N_16142,N_16144);
nor U16406 (N_16406,N_16005,N_15904);
or U16407 (N_16407,N_16045,N_16169);
nor U16408 (N_16408,N_16014,N_16161);
or U16409 (N_16409,N_16022,N_15938);
xnor U16410 (N_16410,N_15964,N_16035);
and U16411 (N_16411,N_15909,N_16139);
xor U16412 (N_16412,N_15961,N_16013);
nor U16413 (N_16413,N_16105,N_16189);
or U16414 (N_16414,N_16059,N_16052);
nor U16415 (N_16415,N_16070,N_15912);
nand U16416 (N_16416,N_16019,N_16155);
nor U16417 (N_16417,N_16061,N_16153);
or U16418 (N_16418,N_16124,N_16033);
or U16419 (N_16419,N_15962,N_15998);
or U16420 (N_16420,N_15929,N_15947);
nand U16421 (N_16421,N_15983,N_15966);
and U16422 (N_16422,N_16023,N_15906);
nand U16423 (N_16423,N_16041,N_16038);
nor U16424 (N_16424,N_16134,N_16017);
and U16425 (N_16425,N_15999,N_16004);
nand U16426 (N_16426,N_15958,N_15924);
or U16427 (N_16427,N_16123,N_16000);
xnor U16428 (N_16428,N_16092,N_16086);
or U16429 (N_16429,N_16096,N_16129);
or U16430 (N_16430,N_16189,N_16197);
xnor U16431 (N_16431,N_16086,N_16004);
nand U16432 (N_16432,N_15925,N_16083);
or U16433 (N_16433,N_16120,N_16099);
nand U16434 (N_16434,N_16010,N_16047);
xor U16435 (N_16435,N_16124,N_16148);
and U16436 (N_16436,N_16132,N_16128);
or U16437 (N_16437,N_16066,N_15964);
or U16438 (N_16438,N_15927,N_16058);
nand U16439 (N_16439,N_16140,N_16007);
xnor U16440 (N_16440,N_15941,N_15960);
xor U16441 (N_16441,N_16017,N_16090);
nor U16442 (N_16442,N_16090,N_15949);
nor U16443 (N_16443,N_16194,N_15928);
or U16444 (N_16444,N_16054,N_15989);
nand U16445 (N_16445,N_16016,N_15967);
xor U16446 (N_16446,N_16062,N_16176);
xnor U16447 (N_16447,N_16148,N_16069);
nor U16448 (N_16448,N_15983,N_16148);
and U16449 (N_16449,N_16095,N_16148);
xnor U16450 (N_16450,N_15976,N_16125);
and U16451 (N_16451,N_16191,N_16085);
nand U16452 (N_16452,N_16082,N_15974);
or U16453 (N_16453,N_15919,N_15932);
xnor U16454 (N_16454,N_16152,N_15997);
nand U16455 (N_16455,N_16036,N_16186);
nor U16456 (N_16456,N_15902,N_16014);
nor U16457 (N_16457,N_15908,N_16139);
and U16458 (N_16458,N_15922,N_16024);
xor U16459 (N_16459,N_16010,N_16102);
xor U16460 (N_16460,N_16121,N_16157);
nor U16461 (N_16461,N_16059,N_16148);
nand U16462 (N_16462,N_15970,N_16146);
nand U16463 (N_16463,N_16012,N_16097);
nor U16464 (N_16464,N_16145,N_16183);
or U16465 (N_16465,N_16002,N_15957);
or U16466 (N_16466,N_16157,N_15908);
xnor U16467 (N_16467,N_16161,N_15954);
nor U16468 (N_16468,N_15939,N_16178);
or U16469 (N_16469,N_16063,N_15933);
nand U16470 (N_16470,N_16122,N_15902);
or U16471 (N_16471,N_16036,N_15946);
or U16472 (N_16472,N_16040,N_16147);
xor U16473 (N_16473,N_15900,N_15989);
and U16474 (N_16474,N_16119,N_16044);
and U16475 (N_16475,N_16158,N_15950);
or U16476 (N_16476,N_15992,N_16080);
nor U16477 (N_16477,N_16176,N_15951);
nand U16478 (N_16478,N_16065,N_16116);
nor U16479 (N_16479,N_15998,N_15917);
nand U16480 (N_16480,N_16120,N_15917);
or U16481 (N_16481,N_16017,N_16149);
xor U16482 (N_16482,N_15915,N_16081);
and U16483 (N_16483,N_15938,N_16066);
or U16484 (N_16484,N_16055,N_16008);
nand U16485 (N_16485,N_15932,N_16107);
nand U16486 (N_16486,N_16094,N_15932);
or U16487 (N_16487,N_16089,N_15958);
and U16488 (N_16488,N_16107,N_16097);
and U16489 (N_16489,N_16035,N_16112);
nor U16490 (N_16490,N_15971,N_16073);
xnor U16491 (N_16491,N_16151,N_16027);
xnor U16492 (N_16492,N_15959,N_15971);
nand U16493 (N_16493,N_15957,N_16015);
and U16494 (N_16494,N_15927,N_16131);
or U16495 (N_16495,N_16037,N_16149);
and U16496 (N_16496,N_16020,N_16010);
nor U16497 (N_16497,N_15971,N_15967);
xnor U16498 (N_16498,N_16132,N_16030);
nand U16499 (N_16499,N_15925,N_16042);
nor U16500 (N_16500,N_16240,N_16405);
nand U16501 (N_16501,N_16289,N_16312);
nand U16502 (N_16502,N_16403,N_16427);
or U16503 (N_16503,N_16333,N_16447);
xor U16504 (N_16504,N_16202,N_16206);
nand U16505 (N_16505,N_16367,N_16487);
or U16506 (N_16506,N_16421,N_16390);
or U16507 (N_16507,N_16327,N_16249);
nor U16508 (N_16508,N_16244,N_16460);
xor U16509 (N_16509,N_16365,N_16279);
nand U16510 (N_16510,N_16238,N_16478);
nor U16511 (N_16511,N_16247,N_16307);
nand U16512 (N_16512,N_16462,N_16391);
and U16513 (N_16513,N_16356,N_16233);
or U16514 (N_16514,N_16201,N_16393);
or U16515 (N_16515,N_16493,N_16292);
or U16516 (N_16516,N_16474,N_16344);
and U16517 (N_16517,N_16259,N_16329);
and U16518 (N_16518,N_16451,N_16224);
xnor U16519 (N_16519,N_16433,N_16234);
or U16520 (N_16520,N_16271,N_16281);
or U16521 (N_16521,N_16318,N_16334);
xor U16522 (N_16522,N_16383,N_16291);
nand U16523 (N_16523,N_16210,N_16364);
xor U16524 (N_16524,N_16353,N_16430);
nor U16525 (N_16525,N_16243,N_16398);
xor U16526 (N_16526,N_16337,N_16310);
or U16527 (N_16527,N_16453,N_16273);
and U16528 (N_16528,N_16262,N_16440);
nor U16529 (N_16529,N_16228,N_16268);
nor U16530 (N_16530,N_16250,N_16363);
nor U16531 (N_16531,N_16229,N_16217);
xnor U16532 (N_16532,N_16299,N_16283);
xnor U16533 (N_16533,N_16248,N_16261);
nand U16534 (N_16534,N_16282,N_16388);
xor U16535 (N_16535,N_16232,N_16470);
xor U16536 (N_16536,N_16406,N_16270);
nand U16537 (N_16537,N_16293,N_16456);
nor U16538 (N_16538,N_16352,N_16200);
and U16539 (N_16539,N_16392,N_16311);
and U16540 (N_16540,N_16436,N_16414);
xnor U16541 (N_16541,N_16357,N_16226);
and U16542 (N_16542,N_16236,N_16497);
and U16543 (N_16543,N_16449,N_16490);
nand U16544 (N_16544,N_16242,N_16362);
nor U16545 (N_16545,N_16425,N_16439);
nand U16546 (N_16546,N_16286,N_16446);
or U16547 (N_16547,N_16284,N_16339);
xor U16548 (N_16548,N_16251,N_16420);
xor U16549 (N_16549,N_16256,N_16346);
nor U16550 (N_16550,N_16287,N_16417);
nand U16551 (N_16551,N_16389,N_16257);
xor U16552 (N_16552,N_16354,N_16306);
nor U16553 (N_16553,N_16338,N_16272);
xor U16554 (N_16554,N_16237,N_16209);
xor U16555 (N_16555,N_16336,N_16494);
xnor U16556 (N_16556,N_16409,N_16216);
xor U16557 (N_16557,N_16263,N_16486);
nor U16558 (N_16558,N_16467,N_16215);
nand U16559 (N_16559,N_16347,N_16332);
xor U16560 (N_16560,N_16371,N_16258);
xor U16561 (N_16561,N_16401,N_16492);
and U16562 (N_16562,N_16212,N_16375);
or U16563 (N_16563,N_16372,N_16316);
nand U16564 (N_16564,N_16475,N_16431);
nand U16565 (N_16565,N_16472,N_16477);
xnor U16566 (N_16566,N_16351,N_16252);
nand U16567 (N_16567,N_16481,N_16437);
nand U16568 (N_16568,N_16419,N_16264);
and U16569 (N_16569,N_16384,N_16397);
nand U16570 (N_16570,N_16211,N_16276);
nor U16571 (N_16571,N_16319,N_16482);
and U16572 (N_16572,N_16476,N_16359);
xnor U16573 (N_16573,N_16330,N_16426);
or U16574 (N_16574,N_16459,N_16428);
or U16575 (N_16575,N_16345,N_16402);
xor U16576 (N_16576,N_16328,N_16304);
and U16577 (N_16577,N_16214,N_16239);
xnor U16578 (N_16578,N_16408,N_16297);
and U16579 (N_16579,N_16480,N_16277);
or U16580 (N_16580,N_16223,N_16300);
nor U16581 (N_16581,N_16280,N_16416);
nand U16582 (N_16582,N_16320,N_16368);
nand U16583 (N_16583,N_16444,N_16495);
xor U16584 (N_16584,N_16227,N_16413);
or U16585 (N_16585,N_16491,N_16432);
or U16586 (N_16586,N_16213,N_16322);
nor U16587 (N_16587,N_16349,N_16450);
and U16588 (N_16588,N_16458,N_16455);
or U16589 (N_16589,N_16274,N_16222);
xor U16590 (N_16590,N_16381,N_16423);
or U16591 (N_16591,N_16415,N_16204);
or U16592 (N_16592,N_16323,N_16341);
nand U16593 (N_16593,N_16342,N_16246);
nor U16594 (N_16594,N_16241,N_16321);
or U16595 (N_16595,N_16253,N_16385);
xnor U16596 (N_16596,N_16245,N_16317);
and U16597 (N_16597,N_16326,N_16376);
or U16598 (N_16598,N_16411,N_16422);
nor U16599 (N_16599,N_16360,N_16348);
nand U16600 (N_16600,N_16254,N_16361);
and U16601 (N_16601,N_16309,N_16340);
or U16602 (N_16602,N_16255,N_16441);
or U16603 (N_16603,N_16285,N_16448);
or U16604 (N_16604,N_16313,N_16374);
xnor U16605 (N_16605,N_16479,N_16218);
nand U16606 (N_16606,N_16429,N_16366);
xnor U16607 (N_16607,N_16219,N_16463);
nor U16608 (N_16608,N_16335,N_16469);
and U16609 (N_16609,N_16298,N_16395);
nand U16610 (N_16610,N_16373,N_16488);
or U16611 (N_16611,N_16295,N_16260);
and U16612 (N_16612,N_16484,N_16485);
and U16613 (N_16613,N_16308,N_16386);
or U16614 (N_16614,N_16294,N_16434);
nand U16615 (N_16615,N_16331,N_16203);
xnor U16616 (N_16616,N_16466,N_16404);
nand U16617 (N_16617,N_16370,N_16438);
nor U16618 (N_16618,N_16235,N_16305);
nand U16619 (N_16619,N_16424,N_16269);
nor U16620 (N_16620,N_16473,N_16496);
nand U16621 (N_16621,N_16471,N_16394);
nand U16622 (N_16622,N_16208,N_16498);
or U16623 (N_16623,N_16290,N_16457);
nand U16624 (N_16624,N_16303,N_16489);
or U16625 (N_16625,N_16288,N_16358);
nand U16626 (N_16626,N_16343,N_16278);
xor U16627 (N_16627,N_16499,N_16410);
nor U16628 (N_16628,N_16265,N_16207);
and U16629 (N_16629,N_16400,N_16387);
xnor U16630 (N_16630,N_16452,N_16399);
or U16631 (N_16631,N_16396,N_16301);
or U16632 (N_16632,N_16369,N_16266);
xor U16633 (N_16633,N_16454,N_16382);
or U16634 (N_16634,N_16355,N_16483);
nand U16635 (N_16635,N_16314,N_16221);
nor U16636 (N_16636,N_16468,N_16350);
or U16637 (N_16637,N_16220,N_16230);
nor U16638 (N_16638,N_16464,N_16465);
and U16639 (N_16639,N_16378,N_16205);
and U16640 (N_16640,N_16435,N_16418);
nand U16641 (N_16641,N_16412,N_16231);
and U16642 (N_16642,N_16302,N_16267);
or U16643 (N_16643,N_16442,N_16380);
nor U16644 (N_16644,N_16325,N_16445);
and U16645 (N_16645,N_16324,N_16407);
xnor U16646 (N_16646,N_16225,N_16275);
nor U16647 (N_16647,N_16443,N_16377);
nand U16648 (N_16648,N_16461,N_16296);
nand U16649 (N_16649,N_16315,N_16379);
nand U16650 (N_16650,N_16251,N_16234);
or U16651 (N_16651,N_16203,N_16249);
xnor U16652 (N_16652,N_16209,N_16242);
nand U16653 (N_16653,N_16278,N_16355);
xor U16654 (N_16654,N_16457,N_16452);
and U16655 (N_16655,N_16462,N_16316);
xnor U16656 (N_16656,N_16488,N_16424);
xor U16657 (N_16657,N_16310,N_16389);
nand U16658 (N_16658,N_16373,N_16311);
nand U16659 (N_16659,N_16206,N_16354);
nor U16660 (N_16660,N_16475,N_16486);
nor U16661 (N_16661,N_16411,N_16442);
xor U16662 (N_16662,N_16262,N_16370);
xnor U16663 (N_16663,N_16480,N_16300);
nor U16664 (N_16664,N_16484,N_16466);
xnor U16665 (N_16665,N_16304,N_16366);
or U16666 (N_16666,N_16304,N_16204);
nor U16667 (N_16667,N_16488,N_16240);
and U16668 (N_16668,N_16483,N_16309);
and U16669 (N_16669,N_16405,N_16443);
nand U16670 (N_16670,N_16464,N_16254);
xor U16671 (N_16671,N_16378,N_16390);
and U16672 (N_16672,N_16322,N_16342);
nor U16673 (N_16673,N_16374,N_16433);
or U16674 (N_16674,N_16392,N_16336);
and U16675 (N_16675,N_16369,N_16300);
or U16676 (N_16676,N_16310,N_16316);
or U16677 (N_16677,N_16410,N_16279);
xor U16678 (N_16678,N_16391,N_16299);
or U16679 (N_16679,N_16263,N_16489);
xnor U16680 (N_16680,N_16445,N_16415);
or U16681 (N_16681,N_16359,N_16221);
or U16682 (N_16682,N_16335,N_16260);
xor U16683 (N_16683,N_16457,N_16277);
and U16684 (N_16684,N_16208,N_16398);
nand U16685 (N_16685,N_16476,N_16420);
or U16686 (N_16686,N_16271,N_16266);
xor U16687 (N_16687,N_16324,N_16287);
nor U16688 (N_16688,N_16367,N_16484);
nand U16689 (N_16689,N_16403,N_16441);
nor U16690 (N_16690,N_16382,N_16380);
nand U16691 (N_16691,N_16247,N_16262);
nor U16692 (N_16692,N_16351,N_16316);
and U16693 (N_16693,N_16453,N_16439);
or U16694 (N_16694,N_16427,N_16306);
xnor U16695 (N_16695,N_16379,N_16397);
or U16696 (N_16696,N_16315,N_16397);
nand U16697 (N_16697,N_16374,N_16410);
nand U16698 (N_16698,N_16256,N_16227);
and U16699 (N_16699,N_16324,N_16493);
or U16700 (N_16700,N_16450,N_16249);
nor U16701 (N_16701,N_16468,N_16299);
nand U16702 (N_16702,N_16209,N_16325);
nand U16703 (N_16703,N_16468,N_16488);
nand U16704 (N_16704,N_16200,N_16351);
nand U16705 (N_16705,N_16407,N_16251);
or U16706 (N_16706,N_16426,N_16349);
nor U16707 (N_16707,N_16344,N_16370);
xnor U16708 (N_16708,N_16345,N_16295);
nand U16709 (N_16709,N_16457,N_16267);
or U16710 (N_16710,N_16256,N_16339);
and U16711 (N_16711,N_16260,N_16304);
and U16712 (N_16712,N_16440,N_16407);
nand U16713 (N_16713,N_16396,N_16314);
nand U16714 (N_16714,N_16446,N_16476);
nand U16715 (N_16715,N_16407,N_16327);
xor U16716 (N_16716,N_16328,N_16437);
nor U16717 (N_16717,N_16259,N_16285);
nand U16718 (N_16718,N_16263,N_16357);
and U16719 (N_16719,N_16265,N_16385);
xor U16720 (N_16720,N_16291,N_16353);
or U16721 (N_16721,N_16204,N_16370);
nor U16722 (N_16722,N_16496,N_16260);
xnor U16723 (N_16723,N_16290,N_16341);
xor U16724 (N_16724,N_16419,N_16257);
xnor U16725 (N_16725,N_16241,N_16464);
and U16726 (N_16726,N_16234,N_16300);
and U16727 (N_16727,N_16327,N_16238);
and U16728 (N_16728,N_16493,N_16366);
or U16729 (N_16729,N_16268,N_16300);
nand U16730 (N_16730,N_16448,N_16419);
nor U16731 (N_16731,N_16253,N_16312);
and U16732 (N_16732,N_16315,N_16417);
nand U16733 (N_16733,N_16247,N_16356);
xor U16734 (N_16734,N_16370,N_16424);
nand U16735 (N_16735,N_16413,N_16289);
and U16736 (N_16736,N_16288,N_16327);
xor U16737 (N_16737,N_16238,N_16303);
nand U16738 (N_16738,N_16451,N_16237);
xor U16739 (N_16739,N_16443,N_16340);
nor U16740 (N_16740,N_16298,N_16376);
nand U16741 (N_16741,N_16228,N_16232);
and U16742 (N_16742,N_16204,N_16217);
or U16743 (N_16743,N_16335,N_16425);
or U16744 (N_16744,N_16358,N_16423);
or U16745 (N_16745,N_16426,N_16346);
nor U16746 (N_16746,N_16351,N_16335);
nor U16747 (N_16747,N_16331,N_16247);
nand U16748 (N_16748,N_16323,N_16464);
and U16749 (N_16749,N_16390,N_16388);
nand U16750 (N_16750,N_16361,N_16387);
nand U16751 (N_16751,N_16286,N_16400);
xnor U16752 (N_16752,N_16428,N_16432);
nand U16753 (N_16753,N_16477,N_16448);
nand U16754 (N_16754,N_16301,N_16478);
and U16755 (N_16755,N_16277,N_16499);
and U16756 (N_16756,N_16240,N_16397);
xor U16757 (N_16757,N_16318,N_16236);
nor U16758 (N_16758,N_16344,N_16332);
or U16759 (N_16759,N_16250,N_16312);
nor U16760 (N_16760,N_16238,N_16371);
or U16761 (N_16761,N_16202,N_16458);
xnor U16762 (N_16762,N_16425,N_16476);
nand U16763 (N_16763,N_16218,N_16227);
xor U16764 (N_16764,N_16436,N_16206);
xnor U16765 (N_16765,N_16211,N_16361);
nor U16766 (N_16766,N_16289,N_16361);
nor U16767 (N_16767,N_16318,N_16303);
and U16768 (N_16768,N_16301,N_16202);
and U16769 (N_16769,N_16413,N_16264);
xnor U16770 (N_16770,N_16451,N_16418);
nand U16771 (N_16771,N_16225,N_16319);
or U16772 (N_16772,N_16319,N_16481);
xor U16773 (N_16773,N_16266,N_16261);
xor U16774 (N_16774,N_16372,N_16331);
nor U16775 (N_16775,N_16341,N_16470);
or U16776 (N_16776,N_16494,N_16397);
xor U16777 (N_16777,N_16300,N_16211);
nand U16778 (N_16778,N_16204,N_16454);
nor U16779 (N_16779,N_16474,N_16426);
and U16780 (N_16780,N_16240,N_16470);
xor U16781 (N_16781,N_16370,N_16436);
nor U16782 (N_16782,N_16430,N_16444);
or U16783 (N_16783,N_16201,N_16245);
and U16784 (N_16784,N_16242,N_16312);
and U16785 (N_16785,N_16451,N_16236);
nand U16786 (N_16786,N_16237,N_16457);
or U16787 (N_16787,N_16450,N_16418);
and U16788 (N_16788,N_16497,N_16352);
nor U16789 (N_16789,N_16496,N_16326);
nor U16790 (N_16790,N_16392,N_16307);
and U16791 (N_16791,N_16267,N_16226);
xor U16792 (N_16792,N_16430,N_16476);
or U16793 (N_16793,N_16220,N_16390);
nor U16794 (N_16794,N_16382,N_16427);
nor U16795 (N_16795,N_16468,N_16231);
nand U16796 (N_16796,N_16285,N_16201);
xor U16797 (N_16797,N_16492,N_16347);
and U16798 (N_16798,N_16482,N_16237);
nor U16799 (N_16799,N_16477,N_16443);
xnor U16800 (N_16800,N_16628,N_16522);
nor U16801 (N_16801,N_16719,N_16621);
nor U16802 (N_16802,N_16562,N_16701);
xnor U16803 (N_16803,N_16543,N_16713);
and U16804 (N_16804,N_16609,N_16553);
or U16805 (N_16805,N_16512,N_16755);
nor U16806 (N_16806,N_16655,N_16792);
xnor U16807 (N_16807,N_16581,N_16545);
or U16808 (N_16808,N_16574,N_16617);
or U16809 (N_16809,N_16680,N_16767);
or U16810 (N_16810,N_16779,N_16513);
xor U16811 (N_16811,N_16784,N_16747);
nor U16812 (N_16812,N_16537,N_16633);
and U16813 (N_16813,N_16731,N_16644);
and U16814 (N_16814,N_16514,N_16596);
or U16815 (N_16815,N_16673,N_16667);
or U16816 (N_16816,N_16593,N_16651);
nor U16817 (N_16817,N_16729,N_16650);
nand U16818 (N_16818,N_16796,N_16642);
and U16819 (N_16819,N_16653,N_16619);
nand U16820 (N_16820,N_16720,N_16556);
and U16821 (N_16821,N_16561,N_16600);
and U16822 (N_16822,N_16705,N_16631);
xnor U16823 (N_16823,N_16584,N_16590);
or U16824 (N_16824,N_16568,N_16519);
xor U16825 (N_16825,N_16674,N_16761);
xor U16826 (N_16826,N_16782,N_16575);
or U16827 (N_16827,N_16531,N_16723);
nor U16828 (N_16828,N_16640,N_16707);
or U16829 (N_16829,N_16613,N_16757);
and U16830 (N_16830,N_16622,N_16618);
nor U16831 (N_16831,N_16740,N_16589);
nor U16832 (N_16832,N_16550,N_16520);
nand U16833 (N_16833,N_16503,N_16636);
and U16834 (N_16834,N_16534,N_16739);
nand U16835 (N_16835,N_16635,N_16588);
or U16836 (N_16836,N_16547,N_16546);
or U16837 (N_16837,N_16592,N_16746);
xnor U16838 (N_16838,N_16539,N_16741);
and U16839 (N_16839,N_16607,N_16656);
nor U16840 (N_16840,N_16795,N_16742);
or U16841 (N_16841,N_16798,N_16657);
xnor U16842 (N_16842,N_16548,N_16623);
nor U16843 (N_16843,N_16629,N_16523);
and U16844 (N_16844,N_16610,N_16569);
xnor U16845 (N_16845,N_16709,N_16780);
and U16846 (N_16846,N_16517,N_16598);
xor U16847 (N_16847,N_16677,N_16591);
nor U16848 (N_16848,N_16525,N_16778);
or U16849 (N_16849,N_16699,N_16582);
or U16850 (N_16850,N_16735,N_16536);
nor U16851 (N_16851,N_16730,N_16753);
and U16852 (N_16852,N_16724,N_16762);
and U16853 (N_16853,N_16606,N_16529);
and U16854 (N_16854,N_16580,N_16706);
and U16855 (N_16855,N_16658,N_16726);
and U16856 (N_16856,N_16793,N_16759);
or U16857 (N_16857,N_16603,N_16685);
and U16858 (N_16858,N_16710,N_16664);
or U16859 (N_16859,N_16559,N_16567);
nor U16860 (N_16860,N_16560,N_16776);
nand U16861 (N_16861,N_16502,N_16576);
xor U16862 (N_16862,N_16770,N_16763);
and U16863 (N_16863,N_16785,N_16652);
nand U16864 (N_16864,N_16501,N_16671);
or U16865 (N_16865,N_16689,N_16777);
nand U16866 (N_16866,N_16504,N_16734);
nand U16867 (N_16867,N_16693,N_16614);
xor U16868 (N_16868,N_16708,N_16632);
nor U16869 (N_16869,N_16786,N_16722);
or U16870 (N_16870,N_16712,N_16788);
nor U16871 (N_16871,N_16605,N_16518);
nand U16872 (N_16872,N_16604,N_16748);
xnor U16873 (N_16873,N_16578,N_16783);
xnor U16874 (N_16874,N_16799,N_16661);
nor U16875 (N_16875,N_16571,N_16557);
xor U16876 (N_16876,N_16789,N_16769);
nand U16877 (N_16877,N_16774,N_16544);
and U16878 (N_16878,N_16630,N_16541);
or U16879 (N_16879,N_16725,N_16634);
nor U16880 (N_16880,N_16535,N_16794);
xor U16881 (N_16881,N_16641,N_16597);
and U16882 (N_16882,N_16626,N_16672);
nor U16883 (N_16883,N_16552,N_16756);
nor U16884 (N_16884,N_16733,N_16515);
nand U16885 (N_16885,N_16587,N_16624);
or U16886 (N_16886,N_16647,N_16679);
and U16887 (N_16887,N_16585,N_16507);
nand U16888 (N_16888,N_16625,N_16736);
xnor U16889 (N_16889,N_16524,N_16715);
xnor U16890 (N_16890,N_16595,N_16566);
xor U16891 (N_16891,N_16586,N_16649);
nor U16892 (N_16892,N_16521,N_16564);
or U16893 (N_16893,N_16768,N_16695);
nand U16894 (N_16894,N_16773,N_16620);
and U16895 (N_16895,N_16665,N_16781);
and U16896 (N_16896,N_16775,N_16717);
xor U16897 (N_16897,N_16660,N_16654);
or U16898 (N_16898,N_16754,N_16751);
nor U16899 (N_16899,N_16508,N_16532);
nand U16900 (N_16900,N_16551,N_16615);
xor U16901 (N_16901,N_16749,N_16573);
nand U16902 (N_16902,N_16616,N_16510);
and U16903 (N_16903,N_16530,N_16666);
nand U16904 (N_16904,N_16675,N_16565);
nand U16905 (N_16905,N_16764,N_16738);
nor U16906 (N_16906,N_16700,N_16577);
nor U16907 (N_16907,N_16540,N_16790);
xnor U16908 (N_16908,N_16526,N_16668);
xnor U16909 (N_16909,N_16500,N_16728);
and U16910 (N_16910,N_16602,N_16771);
xnor U16911 (N_16911,N_16750,N_16678);
nor U16912 (N_16912,N_16737,N_16583);
and U16913 (N_16913,N_16687,N_16682);
nand U16914 (N_16914,N_16797,N_16648);
and U16915 (N_16915,N_16601,N_16703);
nor U16916 (N_16916,N_16511,N_16698);
and U16917 (N_16917,N_16627,N_16688);
xnor U16918 (N_16918,N_16527,N_16554);
or U16919 (N_16919,N_16505,N_16638);
and U16920 (N_16920,N_16659,N_16558);
nand U16921 (N_16921,N_16727,N_16684);
or U16922 (N_16922,N_16704,N_16745);
or U16923 (N_16923,N_16599,N_16637);
nor U16924 (N_16924,N_16663,N_16721);
xnor U16925 (N_16925,N_16669,N_16697);
xor U16926 (N_16926,N_16765,N_16643);
nand U16927 (N_16927,N_16711,N_16714);
and U16928 (N_16928,N_16572,N_16716);
xor U16929 (N_16929,N_16760,N_16752);
and U16930 (N_16930,N_16718,N_16608);
or U16931 (N_16931,N_16683,N_16686);
and U16932 (N_16932,N_16787,N_16758);
or U16933 (N_16933,N_16690,N_16772);
and U16934 (N_16934,N_16563,N_16542);
nand U16935 (N_16935,N_16691,N_16676);
nand U16936 (N_16936,N_16639,N_16555);
nor U16937 (N_16937,N_16549,N_16696);
or U16938 (N_16938,N_16791,N_16766);
nor U16939 (N_16939,N_16570,N_16670);
and U16940 (N_16940,N_16594,N_16538);
nand U16941 (N_16941,N_16662,N_16692);
or U16942 (N_16942,N_16611,N_16506);
nor U16943 (N_16943,N_16579,N_16612);
or U16944 (N_16944,N_16702,N_16533);
nand U16945 (N_16945,N_16509,N_16743);
xnor U16946 (N_16946,N_16516,N_16528);
nor U16947 (N_16947,N_16744,N_16646);
nand U16948 (N_16948,N_16681,N_16694);
nor U16949 (N_16949,N_16645,N_16732);
nor U16950 (N_16950,N_16541,N_16597);
xnor U16951 (N_16951,N_16642,N_16729);
xor U16952 (N_16952,N_16684,N_16510);
nand U16953 (N_16953,N_16512,N_16588);
nand U16954 (N_16954,N_16544,N_16719);
nor U16955 (N_16955,N_16688,N_16510);
or U16956 (N_16956,N_16701,N_16772);
or U16957 (N_16957,N_16717,N_16715);
or U16958 (N_16958,N_16589,N_16756);
nand U16959 (N_16959,N_16575,N_16665);
nor U16960 (N_16960,N_16641,N_16672);
and U16961 (N_16961,N_16547,N_16695);
and U16962 (N_16962,N_16657,N_16646);
nand U16963 (N_16963,N_16649,N_16704);
or U16964 (N_16964,N_16723,N_16689);
or U16965 (N_16965,N_16739,N_16629);
or U16966 (N_16966,N_16754,N_16698);
xnor U16967 (N_16967,N_16514,N_16615);
nand U16968 (N_16968,N_16714,N_16684);
nand U16969 (N_16969,N_16520,N_16616);
and U16970 (N_16970,N_16522,N_16626);
nand U16971 (N_16971,N_16547,N_16598);
or U16972 (N_16972,N_16708,N_16727);
xor U16973 (N_16973,N_16560,N_16587);
nor U16974 (N_16974,N_16637,N_16667);
and U16975 (N_16975,N_16746,N_16749);
xnor U16976 (N_16976,N_16765,N_16722);
or U16977 (N_16977,N_16540,N_16564);
xor U16978 (N_16978,N_16750,N_16545);
and U16979 (N_16979,N_16791,N_16626);
nand U16980 (N_16980,N_16586,N_16694);
nand U16981 (N_16981,N_16658,N_16750);
or U16982 (N_16982,N_16647,N_16660);
nand U16983 (N_16983,N_16556,N_16739);
xor U16984 (N_16984,N_16535,N_16719);
and U16985 (N_16985,N_16747,N_16782);
nor U16986 (N_16986,N_16648,N_16573);
nor U16987 (N_16987,N_16638,N_16757);
or U16988 (N_16988,N_16634,N_16619);
nor U16989 (N_16989,N_16534,N_16529);
or U16990 (N_16990,N_16577,N_16753);
nor U16991 (N_16991,N_16596,N_16744);
and U16992 (N_16992,N_16631,N_16510);
nor U16993 (N_16993,N_16772,N_16508);
xor U16994 (N_16994,N_16654,N_16607);
or U16995 (N_16995,N_16792,N_16591);
xor U16996 (N_16996,N_16780,N_16645);
nor U16997 (N_16997,N_16512,N_16749);
and U16998 (N_16998,N_16677,N_16532);
and U16999 (N_16999,N_16501,N_16792);
nand U17000 (N_17000,N_16774,N_16501);
or U17001 (N_17001,N_16761,N_16520);
and U17002 (N_17002,N_16548,N_16553);
and U17003 (N_17003,N_16639,N_16695);
nand U17004 (N_17004,N_16598,N_16796);
or U17005 (N_17005,N_16620,N_16763);
or U17006 (N_17006,N_16597,N_16590);
nor U17007 (N_17007,N_16735,N_16690);
or U17008 (N_17008,N_16790,N_16502);
nor U17009 (N_17009,N_16742,N_16703);
nor U17010 (N_17010,N_16711,N_16541);
xor U17011 (N_17011,N_16789,N_16552);
nor U17012 (N_17012,N_16606,N_16552);
and U17013 (N_17013,N_16513,N_16516);
or U17014 (N_17014,N_16587,N_16755);
nand U17015 (N_17015,N_16795,N_16699);
nand U17016 (N_17016,N_16596,N_16620);
and U17017 (N_17017,N_16630,N_16631);
xnor U17018 (N_17018,N_16594,N_16708);
nand U17019 (N_17019,N_16703,N_16683);
or U17020 (N_17020,N_16612,N_16528);
nor U17021 (N_17021,N_16789,N_16716);
xnor U17022 (N_17022,N_16676,N_16748);
nand U17023 (N_17023,N_16604,N_16761);
nor U17024 (N_17024,N_16785,N_16792);
nor U17025 (N_17025,N_16673,N_16766);
or U17026 (N_17026,N_16644,N_16669);
xnor U17027 (N_17027,N_16565,N_16634);
nand U17028 (N_17028,N_16542,N_16516);
and U17029 (N_17029,N_16737,N_16665);
xnor U17030 (N_17030,N_16586,N_16595);
nor U17031 (N_17031,N_16662,N_16789);
nor U17032 (N_17032,N_16555,N_16582);
and U17033 (N_17033,N_16601,N_16513);
or U17034 (N_17034,N_16602,N_16620);
or U17035 (N_17035,N_16636,N_16772);
nand U17036 (N_17036,N_16524,N_16788);
and U17037 (N_17037,N_16796,N_16767);
nor U17038 (N_17038,N_16686,N_16520);
nand U17039 (N_17039,N_16588,N_16761);
nand U17040 (N_17040,N_16527,N_16539);
nand U17041 (N_17041,N_16628,N_16506);
nand U17042 (N_17042,N_16560,N_16791);
or U17043 (N_17043,N_16794,N_16578);
and U17044 (N_17044,N_16649,N_16569);
xor U17045 (N_17045,N_16727,N_16618);
and U17046 (N_17046,N_16679,N_16550);
nand U17047 (N_17047,N_16697,N_16771);
nand U17048 (N_17048,N_16636,N_16727);
nor U17049 (N_17049,N_16532,N_16640);
xnor U17050 (N_17050,N_16745,N_16536);
nand U17051 (N_17051,N_16583,N_16523);
nand U17052 (N_17052,N_16703,N_16784);
nand U17053 (N_17053,N_16594,N_16726);
nand U17054 (N_17054,N_16587,N_16663);
xnor U17055 (N_17055,N_16768,N_16621);
xnor U17056 (N_17056,N_16767,N_16505);
nor U17057 (N_17057,N_16520,N_16775);
and U17058 (N_17058,N_16765,N_16578);
xnor U17059 (N_17059,N_16671,N_16596);
nand U17060 (N_17060,N_16503,N_16672);
or U17061 (N_17061,N_16732,N_16668);
and U17062 (N_17062,N_16535,N_16652);
and U17063 (N_17063,N_16559,N_16560);
nand U17064 (N_17064,N_16758,N_16796);
and U17065 (N_17065,N_16727,N_16629);
nand U17066 (N_17066,N_16684,N_16732);
nor U17067 (N_17067,N_16536,N_16527);
and U17068 (N_17068,N_16721,N_16537);
or U17069 (N_17069,N_16667,N_16563);
xnor U17070 (N_17070,N_16744,N_16686);
or U17071 (N_17071,N_16787,N_16696);
nor U17072 (N_17072,N_16534,N_16795);
and U17073 (N_17073,N_16614,N_16604);
xnor U17074 (N_17074,N_16715,N_16727);
nor U17075 (N_17075,N_16644,N_16607);
and U17076 (N_17076,N_16631,N_16550);
nor U17077 (N_17077,N_16503,N_16521);
nor U17078 (N_17078,N_16736,N_16563);
or U17079 (N_17079,N_16656,N_16684);
and U17080 (N_17080,N_16777,N_16539);
nand U17081 (N_17081,N_16637,N_16715);
nor U17082 (N_17082,N_16721,N_16529);
nand U17083 (N_17083,N_16599,N_16685);
nand U17084 (N_17084,N_16788,N_16537);
or U17085 (N_17085,N_16721,N_16540);
nor U17086 (N_17086,N_16605,N_16790);
and U17087 (N_17087,N_16762,N_16528);
and U17088 (N_17088,N_16553,N_16584);
nand U17089 (N_17089,N_16563,N_16555);
or U17090 (N_17090,N_16576,N_16690);
and U17091 (N_17091,N_16565,N_16756);
xnor U17092 (N_17092,N_16573,N_16632);
nand U17093 (N_17093,N_16682,N_16560);
nor U17094 (N_17094,N_16631,N_16642);
xnor U17095 (N_17095,N_16768,N_16718);
xnor U17096 (N_17096,N_16792,N_16684);
or U17097 (N_17097,N_16763,N_16704);
or U17098 (N_17098,N_16582,N_16579);
or U17099 (N_17099,N_16779,N_16521);
nor U17100 (N_17100,N_17073,N_17098);
or U17101 (N_17101,N_16880,N_17092);
nor U17102 (N_17102,N_17026,N_17057);
nor U17103 (N_17103,N_17095,N_16899);
and U17104 (N_17104,N_17055,N_17011);
and U17105 (N_17105,N_17076,N_17012);
or U17106 (N_17106,N_17041,N_16868);
nor U17107 (N_17107,N_17020,N_16925);
or U17108 (N_17108,N_17069,N_17049);
or U17109 (N_17109,N_16985,N_17010);
or U17110 (N_17110,N_16916,N_16898);
nand U17111 (N_17111,N_17090,N_16941);
nor U17112 (N_17112,N_16836,N_16883);
xor U17113 (N_17113,N_17022,N_16972);
nor U17114 (N_17114,N_16834,N_17050);
nand U17115 (N_17115,N_16931,N_17039);
or U17116 (N_17116,N_16831,N_16853);
nand U17117 (N_17117,N_17052,N_16966);
nor U17118 (N_17118,N_17056,N_16989);
and U17119 (N_17119,N_17001,N_17006);
xnor U17120 (N_17120,N_16873,N_16818);
nand U17121 (N_17121,N_17034,N_16806);
nor U17122 (N_17122,N_16903,N_16864);
xor U17123 (N_17123,N_17042,N_17091);
and U17124 (N_17124,N_17047,N_16970);
nor U17125 (N_17125,N_16805,N_16803);
xnor U17126 (N_17126,N_16832,N_16847);
nor U17127 (N_17127,N_16852,N_16808);
xor U17128 (N_17128,N_16924,N_16862);
nand U17129 (N_17129,N_16889,N_16912);
or U17130 (N_17130,N_16804,N_16987);
and U17131 (N_17131,N_16894,N_17004);
or U17132 (N_17132,N_16997,N_16950);
nand U17133 (N_17133,N_16877,N_16990);
nor U17134 (N_17134,N_16943,N_17027);
xor U17135 (N_17135,N_16963,N_16977);
xor U17136 (N_17136,N_16967,N_16917);
nor U17137 (N_17137,N_16910,N_17099);
or U17138 (N_17138,N_16976,N_16892);
or U17139 (N_17139,N_16998,N_16962);
and U17140 (N_17140,N_16927,N_16813);
and U17141 (N_17141,N_17059,N_16945);
nor U17142 (N_17142,N_17051,N_16965);
xnor U17143 (N_17143,N_16872,N_16914);
or U17144 (N_17144,N_17077,N_16956);
or U17145 (N_17145,N_16890,N_17023);
xor U17146 (N_17146,N_17066,N_16913);
xnor U17147 (N_17147,N_16844,N_16978);
xnor U17148 (N_17148,N_16930,N_17003);
or U17149 (N_17149,N_16871,N_17053);
xnor U17150 (N_17150,N_17037,N_17044);
xnor U17151 (N_17151,N_16902,N_16909);
nor U17152 (N_17152,N_16802,N_16935);
nand U17153 (N_17153,N_16863,N_16811);
nand U17154 (N_17154,N_16983,N_17009);
nand U17155 (N_17155,N_16933,N_16878);
xor U17156 (N_17156,N_16869,N_16827);
nor U17157 (N_17157,N_16820,N_16879);
and U17158 (N_17158,N_16837,N_16887);
nand U17159 (N_17159,N_16954,N_16857);
and U17160 (N_17160,N_16969,N_17007);
nand U17161 (N_17161,N_16961,N_16891);
or U17162 (N_17162,N_16815,N_16951);
xnor U17163 (N_17163,N_16822,N_16839);
nor U17164 (N_17164,N_17078,N_16854);
xnor U17165 (N_17165,N_16843,N_16896);
and U17166 (N_17166,N_16932,N_17029);
xnor U17167 (N_17167,N_16905,N_16842);
xnor U17168 (N_17168,N_17064,N_17079);
xor U17169 (N_17169,N_16856,N_17030);
and U17170 (N_17170,N_17016,N_16944);
xor U17171 (N_17171,N_16876,N_16981);
and U17172 (N_17172,N_16807,N_16937);
xor U17173 (N_17173,N_17074,N_16870);
or U17174 (N_17174,N_17005,N_17083);
nor U17175 (N_17175,N_17065,N_16838);
nand U17176 (N_17176,N_16800,N_16865);
xnor U17177 (N_17177,N_16918,N_16886);
nand U17178 (N_17178,N_16849,N_16810);
nor U17179 (N_17179,N_16960,N_16904);
nand U17180 (N_17180,N_16875,N_16845);
or U17181 (N_17181,N_16971,N_16915);
or U17182 (N_17182,N_16982,N_16835);
and U17183 (N_17183,N_16957,N_16988);
and U17184 (N_17184,N_16897,N_16929);
or U17185 (N_17185,N_17032,N_16814);
or U17186 (N_17186,N_16801,N_16851);
and U17187 (N_17187,N_17062,N_16816);
or U17188 (N_17188,N_17000,N_17058);
and U17189 (N_17189,N_16858,N_16991);
xor U17190 (N_17190,N_17002,N_16867);
and U17191 (N_17191,N_16830,N_16833);
or U17192 (N_17192,N_16848,N_16934);
xor U17193 (N_17193,N_17013,N_17082);
and U17194 (N_17194,N_16947,N_17017);
or U17195 (N_17195,N_16992,N_17085);
nand U17196 (N_17196,N_17072,N_17094);
xnor U17197 (N_17197,N_16979,N_16828);
or U17198 (N_17198,N_17087,N_17070);
and U17199 (N_17199,N_16819,N_17035);
nor U17200 (N_17200,N_16884,N_16911);
xnor U17201 (N_17201,N_16826,N_17019);
xnor U17202 (N_17202,N_17021,N_16938);
or U17203 (N_17203,N_16999,N_16885);
nor U17204 (N_17204,N_16986,N_16953);
and U17205 (N_17205,N_17067,N_16824);
and U17206 (N_17206,N_17097,N_16975);
xor U17207 (N_17207,N_16959,N_17018);
and U17208 (N_17208,N_16859,N_16952);
nor U17209 (N_17209,N_17048,N_17043);
nand U17210 (N_17210,N_16923,N_17038);
and U17211 (N_17211,N_16996,N_16895);
xnor U17212 (N_17212,N_16829,N_16906);
xor U17213 (N_17213,N_16920,N_17088);
nand U17214 (N_17214,N_16948,N_16955);
and U17215 (N_17215,N_17046,N_17045);
or U17216 (N_17216,N_16949,N_16939);
nand U17217 (N_17217,N_17089,N_16821);
nor U17218 (N_17218,N_16900,N_17093);
nand U17219 (N_17219,N_17084,N_16881);
nor U17220 (N_17220,N_16942,N_16882);
nor U17221 (N_17221,N_17014,N_17096);
and U17222 (N_17222,N_16888,N_16893);
and U17223 (N_17223,N_16861,N_16901);
and U17224 (N_17224,N_17080,N_17075);
xor U17225 (N_17225,N_17036,N_17025);
nand U17226 (N_17226,N_17033,N_16980);
and U17227 (N_17227,N_16840,N_16926);
xor U17228 (N_17228,N_17024,N_16994);
xor U17229 (N_17229,N_17060,N_17028);
nor U17230 (N_17230,N_16866,N_17015);
nand U17231 (N_17231,N_16823,N_16921);
nand U17232 (N_17232,N_16958,N_17063);
or U17233 (N_17233,N_16964,N_16812);
or U17234 (N_17234,N_17071,N_17031);
nor U17235 (N_17235,N_16936,N_16940);
or U17236 (N_17236,N_17040,N_16860);
nand U17237 (N_17237,N_16850,N_16973);
nor U17238 (N_17238,N_17008,N_16825);
xor U17239 (N_17239,N_17054,N_16907);
and U17240 (N_17240,N_16817,N_16993);
xnor U17241 (N_17241,N_17086,N_17068);
xor U17242 (N_17242,N_16995,N_16908);
and U17243 (N_17243,N_16974,N_16841);
or U17244 (N_17244,N_17061,N_16922);
xnor U17245 (N_17245,N_16984,N_16968);
nand U17246 (N_17246,N_17081,N_16928);
xnor U17247 (N_17247,N_16946,N_16855);
xnor U17248 (N_17248,N_16874,N_16919);
and U17249 (N_17249,N_16846,N_16809);
and U17250 (N_17250,N_16872,N_17047);
nand U17251 (N_17251,N_16872,N_16899);
or U17252 (N_17252,N_16988,N_16872);
xnor U17253 (N_17253,N_16959,N_17016);
or U17254 (N_17254,N_16860,N_16919);
xnor U17255 (N_17255,N_16855,N_16962);
nor U17256 (N_17256,N_17015,N_17075);
xnor U17257 (N_17257,N_16933,N_16934);
and U17258 (N_17258,N_16823,N_17060);
and U17259 (N_17259,N_16881,N_17026);
nand U17260 (N_17260,N_17039,N_17096);
or U17261 (N_17261,N_17059,N_17085);
and U17262 (N_17262,N_16970,N_17038);
nor U17263 (N_17263,N_16964,N_16957);
nor U17264 (N_17264,N_17028,N_16902);
xor U17265 (N_17265,N_16846,N_16865);
nand U17266 (N_17266,N_16849,N_16939);
nand U17267 (N_17267,N_17088,N_17058);
nand U17268 (N_17268,N_16986,N_17030);
xnor U17269 (N_17269,N_17034,N_16802);
or U17270 (N_17270,N_16983,N_16897);
xor U17271 (N_17271,N_16827,N_16851);
xnor U17272 (N_17272,N_17049,N_16972);
xnor U17273 (N_17273,N_17095,N_16919);
and U17274 (N_17274,N_16882,N_16937);
nand U17275 (N_17275,N_16986,N_17046);
or U17276 (N_17276,N_16876,N_16804);
and U17277 (N_17277,N_16861,N_16818);
or U17278 (N_17278,N_16888,N_16854);
and U17279 (N_17279,N_16807,N_16811);
nor U17280 (N_17280,N_17028,N_16914);
and U17281 (N_17281,N_16874,N_16817);
or U17282 (N_17282,N_16918,N_16919);
nor U17283 (N_17283,N_16819,N_16977);
xor U17284 (N_17284,N_16902,N_16833);
xor U17285 (N_17285,N_16959,N_16893);
xor U17286 (N_17286,N_16883,N_17074);
or U17287 (N_17287,N_16979,N_16876);
nand U17288 (N_17288,N_17008,N_16816);
and U17289 (N_17289,N_16937,N_16933);
and U17290 (N_17290,N_16926,N_17036);
xor U17291 (N_17291,N_16809,N_16898);
or U17292 (N_17292,N_17039,N_16980);
or U17293 (N_17293,N_16942,N_16832);
xnor U17294 (N_17294,N_16812,N_16864);
nor U17295 (N_17295,N_16997,N_17002);
or U17296 (N_17296,N_17090,N_16885);
nand U17297 (N_17297,N_17099,N_17085);
or U17298 (N_17298,N_16818,N_17042);
and U17299 (N_17299,N_16811,N_16805);
and U17300 (N_17300,N_16919,N_17005);
nand U17301 (N_17301,N_17099,N_17070);
and U17302 (N_17302,N_16815,N_17025);
xor U17303 (N_17303,N_17066,N_16837);
nor U17304 (N_17304,N_16881,N_16802);
and U17305 (N_17305,N_17011,N_16907);
nor U17306 (N_17306,N_16888,N_17081);
xnor U17307 (N_17307,N_17064,N_16981);
or U17308 (N_17308,N_16872,N_16977);
xnor U17309 (N_17309,N_16932,N_17063);
and U17310 (N_17310,N_16837,N_16931);
or U17311 (N_17311,N_16833,N_16922);
nor U17312 (N_17312,N_17006,N_16801);
nor U17313 (N_17313,N_16822,N_17000);
and U17314 (N_17314,N_16983,N_16821);
nor U17315 (N_17315,N_16866,N_16825);
and U17316 (N_17316,N_17063,N_16827);
nor U17317 (N_17317,N_17065,N_17028);
nor U17318 (N_17318,N_17015,N_16878);
and U17319 (N_17319,N_17072,N_17040);
or U17320 (N_17320,N_16853,N_17063);
nor U17321 (N_17321,N_16955,N_16965);
xor U17322 (N_17322,N_16842,N_17001);
nor U17323 (N_17323,N_16928,N_17029);
nand U17324 (N_17324,N_16824,N_16872);
and U17325 (N_17325,N_16922,N_16899);
nor U17326 (N_17326,N_17096,N_17027);
or U17327 (N_17327,N_16917,N_17014);
xnor U17328 (N_17328,N_16815,N_17063);
or U17329 (N_17329,N_16952,N_16979);
nor U17330 (N_17330,N_16935,N_16912);
xnor U17331 (N_17331,N_16831,N_16905);
nand U17332 (N_17332,N_17098,N_16858);
nand U17333 (N_17333,N_16896,N_16913);
xor U17334 (N_17334,N_17090,N_16862);
and U17335 (N_17335,N_16842,N_16884);
and U17336 (N_17336,N_16801,N_17019);
xor U17337 (N_17337,N_17050,N_16891);
nor U17338 (N_17338,N_16821,N_17038);
nor U17339 (N_17339,N_16802,N_16991);
nor U17340 (N_17340,N_16841,N_16943);
xnor U17341 (N_17341,N_17011,N_16903);
and U17342 (N_17342,N_16999,N_16953);
nand U17343 (N_17343,N_17093,N_16833);
or U17344 (N_17344,N_16972,N_16991);
or U17345 (N_17345,N_17030,N_17045);
nand U17346 (N_17346,N_17093,N_16807);
and U17347 (N_17347,N_17023,N_16817);
and U17348 (N_17348,N_17058,N_16853);
nor U17349 (N_17349,N_16865,N_16878);
nand U17350 (N_17350,N_16873,N_17042);
nor U17351 (N_17351,N_16839,N_16913);
and U17352 (N_17352,N_16891,N_17089);
xor U17353 (N_17353,N_16960,N_16989);
xor U17354 (N_17354,N_17050,N_16830);
xor U17355 (N_17355,N_17062,N_17037);
nand U17356 (N_17356,N_16837,N_16936);
xor U17357 (N_17357,N_16876,N_16862);
xnor U17358 (N_17358,N_16975,N_16840);
nand U17359 (N_17359,N_16908,N_16925);
nand U17360 (N_17360,N_16836,N_16894);
or U17361 (N_17361,N_16818,N_16966);
and U17362 (N_17362,N_16950,N_17098);
and U17363 (N_17363,N_16895,N_17084);
xor U17364 (N_17364,N_16994,N_16856);
xor U17365 (N_17365,N_16926,N_17001);
or U17366 (N_17366,N_16921,N_16973);
nor U17367 (N_17367,N_17014,N_17053);
nor U17368 (N_17368,N_16945,N_16948);
and U17369 (N_17369,N_16965,N_17039);
or U17370 (N_17370,N_17007,N_16841);
or U17371 (N_17371,N_16992,N_17036);
nor U17372 (N_17372,N_16868,N_16960);
nand U17373 (N_17373,N_16950,N_16923);
xor U17374 (N_17374,N_16845,N_16807);
nand U17375 (N_17375,N_17016,N_17048);
nand U17376 (N_17376,N_16893,N_16943);
nand U17377 (N_17377,N_16899,N_17023);
and U17378 (N_17378,N_16958,N_17069);
nand U17379 (N_17379,N_16919,N_17033);
xnor U17380 (N_17380,N_16875,N_16842);
nand U17381 (N_17381,N_17099,N_16962);
nor U17382 (N_17382,N_16912,N_16871);
or U17383 (N_17383,N_16998,N_16881);
xor U17384 (N_17384,N_16893,N_16934);
xnor U17385 (N_17385,N_16810,N_17004);
nand U17386 (N_17386,N_16816,N_17056);
nor U17387 (N_17387,N_16834,N_17099);
and U17388 (N_17388,N_17069,N_17056);
xnor U17389 (N_17389,N_16843,N_16928);
and U17390 (N_17390,N_16970,N_16853);
xor U17391 (N_17391,N_16935,N_16818);
nand U17392 (N_17392,N_17033,N_16900);
nor U17393 (N_17393,N_16820,N_16954);
nor U17394 (N_17394,N_17077,N_16818);
or U17395 (N_17395,N_17088,N_17099);
nor U17396 (N_17396,N_17096,N_16812);
nor U17397 (N_17397,N_16812,N_17013);
and U17398 (N_17398,N_16832,N_16908);
and U17399 (N_17399,N_16879,N_17031);
and U17400 (N_17400,N_17162,N_17142);
nor U17401 (N_17401,N_17361,N_17319);
xnor U17402 (N_17402,N_17278,N_17299);
and U17403 (N_17403,N_17171,N_17233);
or U17404 (N_17404,N_17148,N_17131);
nand U17405 (N_17405,N_17213,N_17260);
or U17406 (N_17406,N_17207,N_17373);
nor U17407 (N_17407,N_17225,N_17367);
nor U17408 (N_17408,N_17308,N_17310);
or U17409 (N_17409,N_17335,N_17270);
nor U17410 (N_17410,N_17371,N_17293);
xor U17411 (N_17411,N_17164,N_17140);
xor U17412 (N_17412,N_17156,N_17298);
nor U17413 (N_17413,N_17261,N_17221);
nor U17414 (N_17414,N_17248,N_17258);
and U17415 (N_17415,N_17129,N_17190);
and U17416 (N_17416,N_17269,N_17355);
and U17417 (N_17417,N_17337,N_17117);
nand U17418 (N_17418,N_17352,N_17363);
xor U17419 (N_17419,N_17132,N_17102);
nor U17420 (N_17420,N_17219,N_17262);
nor U17421 (N_17421,N_17229,N_17328);
or U17422 (N_17422,N_17120,N_17377);
nand U17423 (N_17423,N_17118,N_17399);
nand U17424 (N_17424,N_17271,N_17141);
nand U17425 (N_17425,N_17161,N_17397);
nor U17426 (N_17426,N_17199,N_17228);
nand U17427 (N_17427,N_17307,N_17292);
or U17428 (N_17428,N_17101,N_17323);
or U17429 (N_17429,N_17197,N_17191);
or U17430 (N_17430,N_17104,N_17253);
nor U17431 (N_17431,N_17332,N_17163);
nand U17432 (N_17432,N_17303,N_17185);
xnor U17433 (N_17433,N_17110,N_17180);
xnor U17434 (N_17434,N_17344,N_17134);
or U17435 (N_17435,N_17259,N_17317);
nor U17436 (N_17436,N_17331,N_17390);
xor U17437 (N_17437,N_17242,N_17126);
nand U17438 (N_17438,N_17297,N_17247);
xnor U17439 (N_17439,N_17284,N_17144);
or U17440 (N_17440,N_17217,N_17394);
nor U17441 (N_17441,N_17324,N_17153);
xor U17442 (N_17442,N_17179,N_17281);
xnor U17443 (N_17443,N_17183,N_17318);
nand U17444 (N_17444,N_17327,N_17112);
or U17445 (N_17445,N_17158,N_17305);
xor U17446 (N_17446,N_17300,N_17252);
or U17447 (N_17447,N_17325,N_17215);
xor U17448 (N_17448,N_17193,N_17218);
or U17449 (N_17449,N_17379,N_17157);
nand U17450 (N_17450,N_17339,N_17178);
nor U17451 (N_17451,N_17329,N_17301);
nor U17452 (N_17452,N_17238,N_17345);
nand U17453 (N_17453,N_17108,N_17240);
nand U17454 (N_17454,N_17200,N_17314);
nor U17455 (N_17455,N_17145,N_17383);
xnor U17456 (N_17456,N_17338,N_17273);
or U17457 (N_17457,N_17111,N_17257);
nor U17458 (N_17458,N_17155,N_17277);
xnor U17459 (N_17459,N_17234,N_17174);
xor U17460 (N_17460,N_17268,N_17266);
nor U17461 (N_17461,N_17378,N_17280);
or U17462 (N_17462,N_17276,N_17149);
nand U17463 (N_17463,N_17226,N_17232);
xnor U17464 (N_17464,N_17398,N_17351);
nor U17465 (N_17465,N_17154,N_17243);
nor U17466 (N_17466,N_17205,N_17194);
nor U17467 (N_17467,N_17249,N_17166);
xor U17468 (N_17468,N_17302,N_17267);
and U17469 (N_17469,N_17182,N_17103);
xor U17470 (N_17470,N_17186,N_17357);
or U17471 (N_17471,N_17152,N_17105);
nor U17472 (N_17472,N_17336,N_17125);
nor U17473 (N_17473,N_17356,N_17244);
xnor U17474 (N_17474,N_17384,N_17211);
nor U17475 (N_17475,N_17136,N_17347);
nand U17476 (N_17476,N_17151,N_17306);
nor U17477 (N_17477,N_17388,N_17181);
nand U17478 (N_17478,N_17294,N_17195);
nor U17479 (N_17479,N_17313,N_17263);
nor U17480 (N_17480,N_17382,N_17359);
nand U17481 (N_17481,N_17321,N_17150);
and U17482 (N_17482,N_17184,N_17121);
and U17483 (N_17483,N_17177,N_17208);
and U17484 (N_17484,N_17288,N_17212);
nor U17485 (N_17485,N_17380,N_17170);
or U17486 (N_17486,N_17393,N_17167);
nor U17487 (N_17487,N_17372,N_17204);
xor U17488 (N_17488,N_17387,N_17113);
nor U17489 (N_17489,N_17265,N_17311);
xor U17490 (N_17490,N_17330,N_17349);
and U17491 (N_17491,N_17369,N_17312);
and U17492 (N_17492,N_17346,N_17202);
nand U17493 (N_17493,N_17236,N_17285);
and U17494 (N_17494,N_17275,N_17139);
or U17495 (N_17495,N_17322,N_17224);
and U17496 (N_17496,N_17289,N_17395);
or U17497 (N_17497,N_17287,N_17386);
nand U17498 (N_17498,N_17159,N_17235);
or U17499 (N_17499,N_17348,N_17165);
nor U17500 (N_17500,N_17138,N_17214);
nor U17501 (N_17501,N_17133,N_17206);
nor U17502 (N_17502,N_17123,N_17175);
nor U17503 (N_17503,N_17230,N_17209);
or U17504 (N_17504,N_17256,N_17231);
nor U17505 (N_17505,N_17137,N_17295);
nor U17506 (N_17506,N_17146,N_17135);
and U17507 (N_17507,N_17147,N_17210);
nor U17508 (N_17508,N_17222,N_17362);
and U17509 (N_17509,N_17188,N_17143);
nor U17510 (N_17510,N_17114,N_17391);
xnor U17511 (N_17511,N_17350,N_17360);
nand U17512 (N_17512,N_17169,N_17189);
xor U17513 (N_17513,N_17353,N_17196);
nand U17514 (N_17514,N_17333,N_17246);
or U17515 (N_17515,N_17315,N_17291);
and U17516 (N_17516,N_17341,N_17130);
nor U17517 (N_17517,N_17389,N_17245);
xor U17518 (N_17518,N_17176,N_17366);
and U17519 (N_17519,N_17396,N_17122);
xor U17520 (N_17520,N_17320,N_17115);
or U17521 (N_17521,N_17250,N_17296);
and U17522 (N_17522,N_17201,N_17376);
xor U17523 (N_17523,N_17239,N_17342);
nand U17524 (N_17524,N_17223,N_17286);
nand U17525 (N_17525,N_17116,N_17283);
or U17526 (N_17526,N_17375,N_17368);
xnor U17527 (N_17527,N_17290,N_17264);
nand U17528 (N_17528,N_17392,N_17124);
or U17529 (N_17529,N_17119,N_17279);
or U17530 (N_17530,N_17237,N_17340);
nor U17531 (N_17531,N_17127,N_17187);
xnor U17532 (N_17532,N_17326,N_17251);
or U17533 (N_17533,N_17160,N_17216);
or U17534 (N_17534,N_17316,N_17227);
or U17535 (N_17535,N_17128,N_17109);
or U17536 (N_17536,N_17173,N_17106);
nor U17537 (N_17537,N_17255,N_17172);
xnor U17538 (N_17538,N_17358,N_17100);
nand U17539 (N_17539,N_17274,N_17364);
or U17540 (N_17540,N_17365,N_17203);
or U17541 (N_17541,N_17304,N_17220);
xnor U17542 (N_17542,N_17354,N_17370);
nand U17543 (N_17543,N_17107,N_17198);
nand U17544 (N_17544,N_17272,N_17241);
xor U17545 (N_17545,N_17282,N_17381);
and U17546 (N_17546,N_17254,N_17309);
nand U17547 (N_17547,N_17385,N_17343);
and U17548 (N_17548,N_17374,N_17168);
and U17549 (N_17549,N_17334,N_17192);
or U17550 (N_17550,N_17354,N_17116);
xor U17551 (N_17551,N_17265,N_17185);
or U17552 (N_17552,N_17237,N_17281);
xnor U17553 (N_17553,N_17380,N_17319);
xnor U17554 (N_17554,N_17399,N_17276);
xnor U17555 (N_17555,N_17214,N_17285);
xor U17556 (N_17556,N_17310,N_17106);
nor U17557 (N_17557,N_17331,N_17254);
nand U17558 (N_17558,N_17231,N_17226);
xor U17559 (N_17559,N_17232,N_17204);
nand U17560 (N_17560,N_17368,N_17290);
nor U17561 (N_17561,N_17299,N_17340);
nand U17562 (N_17562,N_17212,N_17250);
nor U17563 (N_17563,N_17181,N_17209);
and U17564 (N_17564,N_17122,N_17235);
nor U17565 (N_17565,N_17298,N_17182);
nand U17566 (N_17566,N_17339,N_17283);
nor U17567 (N_17567,N_17155,N_17330);
xnor U17568 (N_17568,N_17243,N_17168);
and U17569 (N_17569,N_17322,N_17368);
xor U17570 (N_17570,N_17238,N_17148);
or U17571 (N_17571,N_17160,N_17297);
and U17572 (N_17572,N_17299,N_17362);
nor U17573 (N_17573,N_17267,N_17132);
or U17574 (N_17574,N_17267,N_17339);
and U17575 (N_17575,N_17254,N_17278);
and U17576 (N_17576,N_17252,N_17222);
and U17577 (N_17577,N_17126,N_17220);
nand U17578 (N_17578,N_17365,N_17191);
or U17579 (N_17579,N_17292,N_17393);
or U17580 (N_17580,N_17127,N_17344);
and U17581 (N_17581,N_17186,N_17132);
and U17582 (N_17582,N_17225,N_17200);
or U17583 (N_17583,N_17262,N_17147);
and U17584 (N_17584,N_17347,N_17329);
or U17585 (N_17585,N_17274,N_17114);
or U17586 (N_17586,N_17318,N_17278);
or U17587 (N_17587,N_17380,N_17205);
nor U17588 (N_17588,N_17300,N_17253);
nand U17589 (N_17589,N_17354,N_17350);
nand U17590 (N_17590,N_17136,N_17339);
nand U17591 (N_17591,N_17202,N_17242);
xnor U17592 (N_17592,N_17322,N_17124);
nor U17593 (N_17593,N_17290,N_17394);
nor U17594 (N_17594,N_17344,N_17398);
and U17595 (N_17595,N_17101,N_17151);
or U17596 (N_17596,N_17365,N_17128);
nand U17597 (N_17597,N_17195,N_17392);
and U17598 (N_17598,N_17236,N_17359);
or U17599 (N_17599,N_17243,N_17257);
or U17600 (N_17600,N_17228,N_17246);
xor U17601 (N_17601,N_17288,N_17230);
and U17602 (N_17602,N_17371,N_17308);
or U17603 (N_17603,N_17142,N_17285);
xnor U17604 (N_17604,N_17331,N_17248);
nand U17605 (N_17605,N_17261,N_17243);
nand U17606 (N_17606,N_17200,N_17343);
or U17607 (N_17607,N_17347,N_17233);
or U17608 (N_17608,N_17119,N_17312);
or U17609 (N_17609,N_17295,N_17167);
nor U17610 (N_17610,N_17346,N_17273);
nor U17611 (N_17611,N_17344,N_17140);
xor U17612 (N_17612,N_17213,N_17358);
and U17613 (N_17613,N_17340,N_17234);
xor U17614 (N_17614,N_17231,N_17128);
xnor U17615 (N_17615,N_17175,N_17267);
and U17616 (N_17616,N_17161,N_17356);
nor U17617 (N_17617,N_17398,N_17192);
xor U17618 (N_17618,N_17219,N_17396);
and U17619 (N_17619,N_17285,N_17140);
xor U17620 (N_17620,N_17109,N_17222);
nand U17621 (N_17621,N_17221,N_17208);
nand U17622 (N_17622,N_17366,N_17378);
and U17623 (N_17623,N_17236,N_17299);
xor U17624 (N_17624,N_17136,N_17157);
xnor U17625 (N_17625,N_17365,N_17236);
and U17626 (N_17626,N_17375,N_17372);
xor U17627 (N_17627,N_17345,N_17350);
and U17628 (N_17628,N_17241,N_17137);
and U17629 (N_17629,N_17147,N_17180);
xor U17630 (N_17630,N_17302,N_17102);
nand U17631 (N_17631,N_17285,N_17237);
and U17632 (N_17632,N_17148,N_17145);
xnor U17633 (N_17633,N_17321,N_17362);
xnor U17634 (N_17634,N_17257,N_17135);
and U17635 (N_17635,N_17328,N_17365);
nor U17636 (N_17636,N_17399,N_17203);
and U17637 (N_17637,N_17341,N_17203);
nor U17638 (N_17638,N_17163,N_17191);
nor U17639 (N_17639,N_17158,N_17224);
nand U17640 (N_17640,N_17167,N_17365);
nor U17641 (N_17641,N_17149,N_17367);
and U17642 (N_17642,N_17184,N_17226);
xnor U17643 (N_17643,N_17276,N_17304);
and U17644 (N_17644,N_17123,N_17191);
and U17645 (N_17645,N_17100,N_17365);
and U17646 (N_17646,N_17208,N_17175);
or U17647 (N_17647,N_17219,N_17291);
xor U17648 (N_17648,N_17313,N_17234);
or U17649 (N_17649,N_17297,N_17116);
or U17650 (N_17650,N_17334,N_17347);
nor U17651 (N_17651,N_17130,N_17336);
and U17652 (N_17652,N_17258,N_17374);
and U17653 (N_17653,N_17340,N_17354);
nand U17654 (N_17654,N_17354,N_17115);
nand U17655 (N_17655,N_17166,N_17185);
nand U17656 (N_17656,N_17377,N_17262);
xor U17657 (N_17657,N_17319,N_17306);
nand U17658 (N_17658,N_17232,N_17181);
xnor U17659 (N_17659,N_17280,N_17239);
nor U17660 (N_17660,N_17140,N_17245);
xor U17661 (N_17661,N_17109,N_17190);
nor U17662 (N_17662,N_17253,N_17206);
and U17663 (N_17663,N_17191,N_17193);
nor U17664 (N_17664,N_17253,N_17317);
or U17665 (N_17665,N_17388,N_17197);
and U17666 (N_17666,N_17237,N_17273);
xnor U17667 (N_17667,N_17168,N_17190);
nor U17668 (N_17668,N_17261,N_17367);
nor U17669 (N_17669,N_17165,N_17355);
xor U17670 (N_17670,N_17260,N_17182);
or U17671 (N_17671,N_17192,N_17102);
nand U17672 (N_17672,N_17399,N_17263);
xor U17673 (N_17673,N_17121,N_17197);
and U17674 (N_17674,N_17160,N_17279);
or U17675 (N_17675,N_17107,N_17105);
xor U17676 (N_17676,N_17345,N_17229);
xor U17677 (N_17677,N_17324,N_17304);
nand U17678 (N_17678,N_17152,N_17262);
nand U17679 (N_17679,N_17324,N_17336);
nand U17680 (N_17680,N_17149,N_17369);
xor U17681 (N_17681,N_17196,N_17262);
and U17682 (N_17682,N_17357,N_17240);
nor U17683 (N_17683,N_17131,N_17241);
xnor U17684 (N_17684,N_17310,N_17131);
xnor U17685 (N_17685,N_17184,N_17369);
nor U17686 (N_17686,N_17105,N_17306);
nand U17687 (N_17687,N_17284,N_17321);
nand U17688 (N_17688,N_17338,N_17248);
xnor U17689 (N_17689,N_17261,N_17215);
nand U17690 (N_17690,N_17371,N_17381);
nand U17691 (N_17691,N_17148,N_17384);
nor U17692 (N_17692,N_17234,N_17316);
xnor U17693 (N_17693,N_17263,N_17245);
or U17694 (N_17694,N_17141,N_17138);
and U17695 (N_17695,N_17361,N_17283);
and U17696 (N_17696,N_17283,N_17323);
nand U17697 (N_17697,N_17374,N_17352);
nand U17698 (N_17698,N_17207,N_17240);
nand U17699 (N_17699,N_17167,N_17284);
nor U17700 (N_17700,N_17472,N_17494);
nor U17701 (N_17701,N_17541,N_17603);
or U17702 (N_17702,N_17584,N_17500);
nor U17703 (N_17703,N_17688,N_17487);
nor U17704 (N_17704,N_17548,N_17662);
or U17705 (N_17705,N_17474,N_17427);
nand U17706 (N_17706,N_17609,N_17608);
or U17707 (N_17707,N_17539,N_17461);
xnor U17708 (N_17708,N_17645,N_17590);
and U17709 (N_17709,N_17522,N_17643);
and U17710 (N_17710,N_17621,N_17518);
nand U17711 (N_17711,N_17563,N_17479);
xor U17712 (N_17712,N_17591,N_17554);
or U17713 (N_17713,N_17656,N_17660);
xnor U17714 (N_17714,N_17477,N_17686);
and U17715 (N_17715,N_17549,N_17690);
or U17716 (N_17716,N_17445,N_17529);
and U17717 (N_17717,N_17490,N_17484);
nand U17718 (N_17718,N_17499,N_17544);
nand U17719 (N_17719,N_17501,N_17587);
xor U17720 (N_17720,N_17543,N_17476);
and U17721 (N_17721,N_17663,N_17633);
or U17722 (N_17722,N_17630,N_17446);
or U17723 (N_17723,N_17460,N_17534);
xor U17724 (N_17724,N_17683,N_17561);
nand U17725 (N_17725,N_17449,N_17689);
and U17726 (N_17726,N_17575,N_17433);
and U17727 (N_17727,N_17564,N_17546);
nand U17728 (N_17728,N_17435,N_17647);
and U17729 (N_17729,N_17611,N_17443);
and U17730 (N_17730,N_17448,N_17637);
or U17731 (N_17731,N_17417,N_17439);
or U17732 (N_17732,N_17592,N_17400);
nor U17733 (N_17733,N_17558,N_17502);
and U17734 (N_17734,N_17426,N_17698);
nor U17735 (N_17735,N_17526,N_17465);
xnor U17736 (N_17736,N_17516,N_17676);
nor U17737 (N_17737,N_17491,N_17600);
xor U17738 (N_17738,N_17455,N_17551);
nor U17739 (N_17739,N_17595,N_17458);
and U17740 (N_17740,N_17638,N_17519);
and U17741 (N_17741,N_17412,N_17692);
nand U17742 (N_17742,N_17453,N_17661);
and U17743 (N_17743,N_17654,N_17614);
xnor U17744 (N_17744,N_17685,N_17639);
xor U17745 (N_17745,N_17571,N_17536);
xnor U17746 (N_17746,N_17635,N_17644);
or U17747 (N_17747,N_17521,N_17623);
xor U17748 (N_17748,N_17425,N_17576);
xnor U17749 (N_17749,N_17406,N_17462);
or U17750 (N_17750,N_17679,N_17678);
xnor U17751 (N_17751,N_17613,N_17489);
and U17752 (N_17752,N_17624,N_17533);
and U17753 (N_17753,N_17415,N_17673);
or U17754 (N_17754,N_17601,N_17572);
or U17755 (N_17755,N_17511,N_17599);
nor U17756 (N_17756,N_17681,N_17566);
xor U17757 (N_17757,N_17636,N_17421);
and U17758 (N_17758,N_17514,N_17675);
and U17759 (N_17759,N_17646,N_17506);
nor U17760 (N_17760,N_17431,N_17414);
nand U17761 (N_17761,N_17403,N_17481);
nand U17762 (N_17762,N_17666,N_17618);
or U17763 (N_17763,N_17694,N_17402);
nor U17764 (N_17764,N_17582,N_17670);
xor U17765 (N_17765,N_17416,N_17664);
xor U17766 (N_17766,N_17653,N_17610);
or U17767 (N_17767,N_17419,N_17615);
xnor U17768 (N_17768,N_17562,N_17648);
and U17769 (N_17769,N_17424,N_17578);
nor U17770 (N_17770,N_17464,N_17550);
and U17771 (N_17771,N_17510,N_17454);
nor U17772 (N_17772,N_17493,N_17565);
nor U17773 (N_17773,N_17428,N_17588);
nand U17774 (N_17774,N_17413,N_17629);
xor U17775 (N_17775,N_17408,N_17674);
nand U17776 (N_17776,N_17441,N_17482);
xnor U17777 (N_17777,N_17655,N_17513);
nand U17778 (N_17778,N_17530,N_17496);
and U17779 (N_17779,N_17498,N_17657);
xor U17780 (N_17780,N_17569,N_17467);
xnor U17781 (N_17781,N_17488,N_17555);
and U17782 (N_17782,N_17440,N_17557);
nand U17783 (N_17783,N_17410,N_17696);
or U17784 (N_17784,N_17581,N_17617);
nor U17785 (N_17785,N_17560,N_17520);
xnor U17786 (N_17786,N_17527,N_17622);
nor U17787 (N_17787,N_17537,N_17671);
nand U17788 (N_17788,N_17407,N_17602);
or U17789 (N_17789,N_17612,N_17432);
or U17790 (N_17790,N_17475,N_17650);
xnor U17791 (N_17791,N_17568,N_17628);
xor U17792 (N_17792,N_17471,N_17447);
nor U17793 (N_17793,N_17509,N_17409);
nor U17794 (N_17794,N_17525,N_17437);
xnor U17795 (N_17795,N_17631,N_17695);
and U17796 (N_17796,N_17463,N_17556);
nor U17797 (N_17797,N_17606,N_17697);
and U17798 (N_17798,N_17684,N_17542);
xor U17799 (N_17799,N_17559,N_17497);
or U17800 (N_17800,N_17570,N_17418);
and U17801 (N_17801,N_17658,N_17665);
nand U17802 (N_17802,N_17545,N_17423);
nand U17803 (N_17803,N_17405,N_17579);
nor U17804 (N_17804,N_17589,N_17508);
nor U17805 (N_17805,N_17597,N_17436);
or U17806 (N_17806,N_17457,N_17620);
nand U17807 (N_17807,N_17401,N_17507);
xor U17808 (N_17808,N_17450,N_17486);
or U17809 (N_17809,N_17430,N_17524);
xnor U17810 (N_17810,N_17640,N_17668);
xnor U17811 (N_17811,N_17625,N_17538);
xor U17812 (N_17812,N_17585,N_17649);
and U17813 (N_17813,N_17693,N_17573);
nand U17814 (N_17814,N_17485,N_17677);
xor U17815 (N_17815,N_17626,N_17429);
xor U17816 (N_17816,N_17619,N_17528);
xnor U17817 (N_17817,N_17480,N_17456);
and U17818 (N_17818,N_17605,N_17532);
nand U17819 (N_17819,N_17604,N_17552);
nand U17820 (N_17820,N_17452,N_17669);
and U17821 (N_17821,N_17607,N_17680);
or U17822 (N_17822,N_17478,N_17687);
and U17823 (N_17823,N_17632,N_17451);
xnor U17824 (N_17824,N_17652,N_17512);
and U17825 (N_17825,N_17503,N_17699);
nor U17826 (N_17826,N_17517,N_17438);
and U17827 (N_17827,N_17470,N_17627);
or U17828 (N_17828,N_17483,N_17442);
or U17829 (N_17829,N_17667,N_17553);
or U17830 (N_17830,N_17598,N_17492);
and U17831 (N_17831,N_17580,N_17682);
xnor U17832 (N_17832,N_17523,N_17444);
nor U17833 (N_17833,N_17616,N_17641);
nand U17834 (N_17834,N_17473,N_17586);
nor U17835 (N_17835,N_17567,N_17547);
nor U17836 (N_17836,N_17411,N_17642);
and U17837 (N_17837,N_17531,N_17466);
nand U17838 (N_17838,N_17594,N_17634);
and U17839 (N_17839,N_17596,N_17434);
or U17840 (N_17840,N_17593,N_17574);
xor U17841 (N_17841,N_17404,N_17420);
nor U17842 (N_17842,N_17659,N_17468);
xnor U17843 (N_17843,N_17459,N_17515);
or U17844 (N_17844,N_17469,N_17535);
nand U17845 (N_17845,N_17691,N_17577);
xnor U17846 (N_17846,N_17672,N_17651);
nand U17847 (N_17847,N_17505,N_17422);
nand U17848 (N_17848,N_17495,N_17540);
and U17849 (N_17849,N_17583,N_17504);
and U17850 (N_17850,N_17662,N_17554);
or U17851 (N_17851,N_17685,N_17567);
and U17852 (N_17852,N_17607,N_17550);
xnor U17853 (N_17853,N_17578,N_17420);
and U17854 (N_17854,N_17522,N_17667);
nor U17855 (N_17855,N_17675,N_17698);
xor U17856 (N_17856,N_17472,N_17550);
nand U17857 (N_17857,N_17419,N_17625);
or U17858 (N_17858,N_17491,N_17630);
nand U17859 (N_17859,N_17585,N_17582);
nand U17860 (N_17860,N_17606,N_17560);
nor U17861 (N_17861,N_17589,N_17646);
nor U17862 (N_17862,N_17544,N_17579);
nand U17863 (N_17863,N_17594,N_17649);
nor U17864 (N_17864,N_17462,N_17648);
and U17865 (N_17865,N_17645,N_17518);
and U17866 (N_17866,N_17588,N_17689);
xor U17867 (N_17867,N_17580,N_17571);
nand U17868 (N_17868,N_17421,N_17412);
nor U17869 (N_17869,N_17574,N_17591);
or U17870 (N_17870,N_17467,N_17576);
xor U17871 (N_17871,N_17693,N_17641);
or U17872 (N_17872,N_17608,N_17644);
and U17873 (N_17873,N_17627,N_17469);
and U17874 (N_17874,N_17644,N_17589);
xnor U17875 (N_17875,N_17596,N_17548);
nand U17876 (N_17876,N_17590,N_17545);
nor U17877 (N_17877,N_17484,N_17500);
or U17878 (N_17878,N_17563,N_17458);
or U17879 (N_17879,N_17605,N_17488);
nor U17880 (N_17880,N_17512,N_17491);
or U17881 (N_17881,N_17658,N_17549);
and U17882 (N_17882,N_17549,N_17694);
nand U17883 (N_17883,N_17510,N_17488);
nor U17884 (N_17884,N_17582,N_17519);
nor U17885 (N_17885,N_17506,N_17487);
xor U17886 (N_17886,N_17595,N_17484);
xnor U17887 (N_17887,N_17441,N_17519);
nor U17888 (N_17888,N_17500,N_17452);
or U17889 (N_17889,N_17693,N_17530);
nand U17890 (N_17890,N_17598,N_17639);
or U17891 (N_17891,N_17647,N_17481);
nor U17892 (N_17892,N_17568,N_17596);
or U17893 (N_17893,N_17431,N_17481);
nand U17894 (N_17894,N_17500,N_17421);
nand U17895 (N_17895,N_17448,N_17682);
nor U17896 (N_17896,N_17548,N_17496);
and U17897 (N_17897,N_17549,N_17418);
nor U17898 (N_17898,N_17464,N_17543);
nand U17899 (N_17899,N_17482,N_17551);
and U17900 (N_17900,N_17410,N_17471);
and U17901 (N_17901,N_17630,N_17440);
nor U17902 (N_17902,N_17547,N_17552);
and U17903 (N_17903,N_17691,N_17588);
and U17904 (N_17904,N_17684,N_17685);
xnor U17905 (N_17905,N_17468,N_17408);
nor U17906 (N_17906,N_17440,N_17616);
or U17907 (N_17907,N_17694,N_17677);
nand U17908 (N_17908,N_17672,N_17428);
nand U17909 (N_17909,N_17533,N_17457);
nand U17910 (N_17910,N_17534,N_17512);
xnor U17911 (N_17911,N_17566,N_17639);
or U17912 (N_17912,N_17456,N_17524);
or U17913 (N_17913,N_17559,N_17463);
or U17914 (N_17914,N_17431,N_17493);
nand U17915 (N_17915,N_17666,N_17574);
or U17916 (N_17916,N_17638,N_17600);
xnor U17917 (N_17917,N_17528,N_17681);
nand U17918 (N_17918,N_17677,N_17665);
xnor U17919 (N_17919,N_17690,N_17402);
nand U17920 (N_17920,N_17497,N_17465);
and U17921 (N_17921,N_17641,N_17613);
nand U17922 (N_17922,N_17618,N_17480);
nor U17923 (N_17923,N_17614,N_17426);
and U17924 (N_17924,N_17442,N_17433);
nand U17925 (N_17925,N_17665,N_17645);
nor U17926 (N_17926,N_17589,N_17431);
nor U17927 (N_17927,N_17546,N_17571);
and U17928 (N_17928,N_17494,N_17537);
xnor U17929 (N_17929,N_17468,N_17562);
or U17930 (N_17930,N_17684,N_17601);
nand U17931 (N_17931,N_17555,N_17685);
xnor U17932 (N_17932,N_17626,N_17413);
nand U17933 (N_17933,N_17512,N_17660);
nor U17934 (N_17934,N_17481,N_17428);
xnor U17935 (N_17935,N_17671,N_17491);
nor U17936 (N_17936,N_17681,N_17569);
and U17937 (N_17937,N_17609,N_17475);
nor U17938 (N_17938,N_17455,N_17468);
or U17939 (N_17939,N_17484,N_17521);
or U17940 (N_17940,N_17660,N_17506);
nor U17941 (N_17941,N_17446,N_17530);
xnor U17942 (N_17942,N_17548,N_17435);
nor U17943 (N_17943,N_17493,N_17509);
and U17944 (N_17944,N_17471,N_17408);
nand U17945 (N_17945,N_17505,N_17517);
xor U17946 (N_17946,N_17588,N_17590);
nand U17947 (N_17947,N_17447,N_17681);
or U17948 (N_17948,N_17558,N_17455);
nand U17949 (N_17949,N_17434,N_17454);
and U17950 (N_17950,N_17642,N_17477);
xnor U17951 (N_17951,N_17515,N_17517);
nand U17952 (N_17952,N_17417,N_17512);
nor U17953 (N_17953,N_17641,N_17588);
xor U17954 (N_17954,N_17674,N_17629);
or U17955 (N_17955,N_17625,N_17597);
or U17956 (N_17956,N_17674,N_17532);
or U17957 (N_17957,N_17668,N_17559);
xor U17958 (N_17958,N_17629,N_17627);
xnor U17959 (N_17959,N_17469,N_17441);
or U17960 (N_17960,N_17458,N_17648);
nor U17961 (N_17961,N_17443,N_17693);
nand U17962 (N_17962,N_17401,N_17438);
and U17963 (N_17963,N_17612,N_17686);
nand U17964 (N_17964,N_17640,N_17597);
nor U17965 (N_17965,N_17560,N_17676);
xnor U17966 (N_17966,N_17476,N_17579);
or U17967 (N_17967,N_17469,N_17540);
or U17968 (N_17968,N_17507,N_17568);
xnor U17969 (N_17969,N_17446,N_17546);
nand U17970 (N_17970,N_17655,N_17413);
nand U17971 (N_17971,N_17423,N_17465);
nor U17972 (N_17972,N_17484,N_17526);
nor U17973 (N_17973,N_17417,N_17596);
xor U17974 (N_17974,N_17401,N_17640);
xnor U17975 (N_17975,N_17570,N_17446);
or U17976 (N_17976,N_17478,N_17694);
nand U17977 (N_17977,N_17625,N_17589);
and U17978 (N_17978,N_17460,N_17553);
nor U17979 (N_17979,N_17421,N_17609);
xor U17980 (N_17980,N_17577,N_17455);
xor U17981 (N_17981,N_17536,N_17407);
nand U17982 (N_17982,N_17559,N_17606);
xor U17983 (N_17983,N_17673,N_17605);
xnor U17984 (N_17984,N_17520,N_17667);
nand U17985 (N_17985,N_17624,N_17475);
and U17986 (N_17986,N_17693,N_17456);
nand U17987 (N_17987,N_17463,N_17694);
nand U17988 (N_17988,N_17540,N_17673);
xnor U17989 (N_17989,N_17549,N_17685);
or U17990 (N_17990,N_17678,N_17419);
nor U17991 (N_17991,N_17452,N_17512);
and U17992 (N_17992,N_17477,N_17671);
nand U17993 (N_17993,N_17472,N_17536);
or U17994 (N_17994,N_17435,N_17599);
nand U17995 (N_17995,N_17475,N_17552);
xnor U17996 (N_17996,N_17553,N_17566);
nor U17997 (N_17997,N_17453,N_17553);
and U17998 (N_17998,N_17515,N_17649);
or U17999 (N_17999,N_17582,N_17501);
nor U18000 (N_18000,N_17911,N_17969);
or U18001 (N_18001,N_17816,N_17734);
or U18002 (N_18002,N_17772,N_17893);
or U18003 (N_18003,N_17704,N_17950);
nand U18004 (N_18004,N_17818,N_17812);
or U18005 (N_18005,N_17973,N_17897);
xnor U18006 (N_18006,N_17861,N_17762);
xnor U18007 (N_18007,N_17865,N_17882);
nand U18008 (N_18008,N_17930,N_17739);
nand U18009 (N_18009,N_17872,N_17994);
xor U18010 (N_18010,N_17776,N_17933);
nor U18011 (N_18011,N_17802,N_17714);
nor U18012 (N_18012,N_17877,N_17741);
xnor U18013 (N_18013,N_17706,N_17868);
and U18014 (N_18014,N_17754,N_17811);
xnor U18015 (N_18015,N_17743,N_17917);
or U18016 (N_18016,N_17855,N_17797);
and U18017 (N_18017,N_17889,N_17819);
nand U18018 (N_18018,N_17932,N_17923);
nand U18019 (N_18019,N_17867,N_17852);
or U18020 (N_18020,N_17866,N_17990);
and U18021 (N_18021,N_17744,N_17738);
and U18022 (N_18022,N_17759,N_17935);
or U18023 (N_18023,N_17902,N_17977);
nor U18024 (N_18024,N_17948,N_17783);
nor U18025 (N_18025,N_17792,N_17862);
xor U18026 (N_18026,N_17901,N_17824);
xnor U18027 (N_18027,N_17860,N_17922);
nor U18028 (N_18028,N_17947,N_17735);
nand U18029 (N_18029,N_17848,N_17747);
xnor U18030 (N_18030,N_17899,N_17884);
nand U18031 (N_18031,N_17849,N_17840);
nor U18032 (N_18032,N_17908,N_17844);
or U18033 (N_18033,N_17954,N_17795);
xor U18034 (N_18034,N_17980,N_17761);
or U18035 (N_18035,N_17916,N_17906);
or U18036 (N_18036,N_17707,N_17767);
xor U18037 (N_18037,N_17719,N_17913);
nor U18038 (N_18038,N_17712,N_17898);
nand U18039 (N_18039,N_17853,N_17752);
nand U18040 (N_18040,N_17750,N_17883);
nor U18041 (N_18041,N_17952,N_17838);
and U18042 (N_18042,N_17846,N_17753);
nor U18043 (N_18043,N_17927,N_17833);
and U18044 (N_18044,N_17788,N_17953);
nor U18045 (N_18045,N_17904,N_17956);
nand U18046 (N_18046,N_17859,N_17920);
nand U18047 (N_18047,N_17907,N_17723);
nand U18048 (N_18048,N_17803,N_17784);
nand U18049 (N_18049,N_17857,N_17722);
and U18050 (N_18050,N_17729,N_17715);
or U18051 (N_18051,N_17988,N_17779);
and U18052 (N_18052,N_17737,N_17800);
and U18053 (N_18053,N_17949,N_17945);
or U18054 (N_18054,N_17894,N_17934);
or U18055 (N_18055,N_17924,N_17998);
and U18056 (N_18056,N_17863,N_17778);
nor U18057 (N_18057,N_17847,N_17881);
xor U18058 (N_18058,N_17957,N_17966);
and U18059 (N_18059,N_17955,N_17826);
xnor U18060 (N_18060,N_17983,N_17978);
nand U18061 (N_18061,N_17773,N_17756);
xnor U18062 (N_18062,N_17742,N_17976);
or U18063 (N_18063,N_17909,N_17926);
and U18064 (N_18064,N_17946,N_17919);
nor U18065 (N_18065,N_17798,N_17769);
and U18066 (N_18066,N_17814,N_17968);
xor U18067 (N_18067,N_17777,N_17905);
or U18068 (N_18068,N_17999,N_17727);
or U18069 (N_18069,N_17710,N_17799);
nor U18070 (N_18070,N_17900,N_17944);
and U18071 (N_18071,N_17912,N_17869);
or U18072 (N_18072,N_17708,N_17961);
nor U18073 (N_18073,N_17965,N_17962);
nand U18074 (N_18074,N_17770,N_17749);
nand U18075 (N_18075,N_17937,N_17891);
nor U18076 (N_18076,N_17748,N_17982);
and U18077 (N_18077,N_17890,N_17972);
and U18078 (N_18078,N_17823,N_17871);
xor U18079 (N_18079,N_17931,N_17989);
xnor U18080 (N_18080,N_17886,N_17760);
and U18081 (N_18081,N_17959,N_17813);
nand U18082 (N_18082,N_17873,N_17766);
nor U18083 (N_18083,N_17718,N_17960);
xor U18084 (N_18084,N_17829,N_17717);
nand U18085 (N_18085,N_17815,N_17929);
and U18086 (N_18086,N_17987,N_17888);
nand U18087 (N_18087,N_17830,N_17786);
xor U18088 (N_18088,N_17822,N_17732);
and U18089 (N_18089,N_17915,N_17997);
or U18090 (N_18090,N_17880,N_17843);
xnor U18091 (N_18091,N_17796,N_17992);
nor U18092 (N_18092,N_17985,N_17771);
nand U18093 (N_18093,N_17974,N_17728);
nor U18094 (N_18094,N_17825,N_17809);
nor U18095 (N_18095,N_17763,N_17791);
and U18096 (N_18096,N_17765,N_17751);
nand U18097 (N_18097,N_17828,N_17836);
nor U18098 (N_18098,N_17793,N_17764);
and U18099 (N_18099,N_17851,N_17993);
and U18100 (N_18100,N_17970,N_17963);
or U18101 (N_18101,N_17746,N_17789);
and U18102 (N_18102,N_17757,N_17910);
or U18103 (N_18103,N_17925,N_17850);
or U18104 (N_18104,N_17892,N_17713);
nor U18105 (N_18105,N_17721,N_17805);
and U18106 (N_18106,N_17781,N_17940);
and U18107 (N_18107,N_17839,N_17858);
nor U18108 (N_18108,N_17705,N_17951);
xor U18109 (N_18109,N_17964,N_17856);
nand U18110 (N_18110,N_17984,N_17967);
or U18111 (N_18111,N_17981,N_17854);
nand U18112 (N_18112,N_17733,N_17979);
nand U18113 (N_18113,N_17870,N_17876);
or U18114 (N_18114,N_17831,N_17755);
nor U18115 (N_18115,N_17995,N_17842);
or U18116 (N_18116,N_17875,N_17817);
or U18117 (N_18117,N_17827,N_17736);
nor U18118 (N_18118,N_17730,N_17936);
nor U18119 (N_18119,N_17832,N_17941);
nor U18120 (N_18120,N_17938,N_17787);
and U18121 (N_18121,N_17971,N_17740);
nor U18122 (N_18122,N_17928,N_17794);
nand U18123 (N_18123,N_17702,N_17986);
nor U18124 (N_18124,N_17975,N_17806);
nor U18125 (N_18125,N_17775,N_17745);
nand U18126 (N_18126,N_17991,N_17808);
nor U18127 (N_18127,N_17921,N_17716);
nor U18128 (N_18128,N_17996,N_17725);
nor U18129 (N_18129,N_17810,N_17701);
and U18130 (N_18130,N_17782,N_17943);
and U18131 (N_18131,N_17731,N_17804);
nor U18132 (N_18132,N_17820,N_17720);
nand U18133 (N_18133,N_17780,N_17834);
or U18134 (N_18134,N_17864,N_17711);
xnor U18135 (N_18135,N_17958,N_17879);
nand U18136 (N_18136,N_17724,N_17807);
or U18137 (N_18137,N_17835,N_17758);
or U18138 (N_18138,N_17841,N_17709);
xnor U18139 (N_18139,N_17874,N_17885);
nor U18140 (N_18140,N_17914,N_17939);
nand U18141 (N_18141,N_17896,N_17918);
and U18142 (N_18142,N_17703,N_17942);
xor U18143 (N_18143,N_17790,N_17768);
xor U18144 (N_18144,N_17726,N_17878);
and U18145 (N_18145,N_17785,N_17774);
xnor U18146 (N_18146,N_17887,N_17821);
xor U18147 (N_18147,N_17837,N_17801);
or U18148 (N_18148,N_17700,N_17845);
and U18149 (N_18149,N_17903,N_17895);
nor U18150 (N_18150,N_17837,N_17978);
nand U18151 (N_18151,N_17781,N_17999);
or U18152 (N_18152,N_17873,N_17986);
or U18153 (N_18153,N_17823,N_17897);
xor U18154 (N_18154,N_17887,N_17969);
or U18155 (N_18155,N_17931,N_17828);
nor U18156 (N_18156,N_17732,N_17853);
and U18157 (N_18157,N_17817,N_17732);
or U18158 (N_18158,N_17905,N_17779);
nand U18159 (N_18159,N_17704,N_17727);
and U18160 (N_18160,N_17732,N_17920);
and U18161 (N_18161,N_17798,N_17998);
xor U18162 (N_18162,N_17700,N_17816);
xor U18163 (N_18163,N_17770,N_17904);
nand U18164 (N_18164,N_17928,N_17863);
xnor U18165 (N_18165,N_17931,N_17962);
nand U18166 (N_18166,N_17796,N_17832);
nand U18167 (N_18167,N_17957,N_17962);
and U18168 (N_18168,N_17730,N_17997);
nand U18169 (N_18169,N_17813,N_17949);
and U18170 (N_18170,N_17854,N_17937);
nor U18171 (N_18171,N_17721,N_17763);
and U18172 (N_18172,N_17898,N_17921);
nor U18173 (N_18173,N_17763,N_17989);
xnor U18174 (N_18174,N_17774,N_17960);
or U18175 (N_18175,N_17763,N_17761);
xnor U18176 (N_18176,N_17841,N_17768);
or U18177 (N_18177,N_17946,N_17930);
and U18178 (N_18178,N_17722,N_17977);
xnor U18179 (N_18179,N_17875,N_17785);
nand U18180 (N_18180,N_17879,N_17700);
xnor U18181 (N_18181,N_17870,N_17843);
nor U18182 (N_18182,N_17969,N_17710);
and U18183 (N_18183,N_17739,N_17873);
nor U18184 (N_18184,N_17754,N_17759);
nand U18185 (N_18185,N_17808,N_17834);
nand U18186 (N_18186,N_17745,N_17930);
nand U18187 (N_18187,N_17971,N_17771);
and U18188 (N_18188,N_17858,N_17707);
or U18189 (N_18189,N_17928,N_17912);
nor U18190 (N_18190,N_17941,N_17786);
xor U18191 (N_18191,N_17936,N_17868);
xnor U18192 (N_18192,N_17750,N_17904);
or U18193 (N_18193,N_17725,N_17913);
nor U18194 (N_18194,N_17759,N_17918);
or U18195 (N_18195,N_17830,N_17783);
nand U18196 (N_18196,N_17721,N_17788);
or U18197 (N_18197,N_17904,N_17763);
xor U18198 (N_18198,N_17700,N_17843);
and U18199 (N_18199,N_17990,N_17984);
nand U18200 (N_18200,N_17859,N_17990);
nand U18201 (N_18201,N_17921,N_17703);
nor U18202 (N_18202,N_17925,N_17800);
nand U18203 (N_18203,N_17735,N_17770);
xnor U18204 (N_18204,N_17848,N_17818);
xnor U18205 (N_18205,N_17857,N_17898);
and U18206 (N_18206,N_17953,N_17837);
xor U18207 (N_18207,N_17880,N_17703);
nand U18208 (N_18208,N_17956,N_17724);
xor U18209 (N_18209,N_17957,N_17843);
or U18210 (N_18210,N_17895,N_17995);
xnor U18211 (N_18211,N_17835,N_17851);
nand U18212 (N_18212,N_17734,N_17898);
xnor U18213 (N_18213,N_17868,N_17738);
xnor U18214 (N_18214,N_17769,N_17706);
nor U18215 (N_18215,N_17770,N_17986);
and U18216 (N_18216,N_17892,N_17949);
xor U18217 (N_18217,N_17770,N_17964);
nor U18218 (N_18218,N_17779,N_17897);
or U18219 (N_18219,N_17786,N_17867);
xnor U18220 (N_18220,N_17976,N_17817);
or U18221 (N_18221,N_17941,N_17988);
nand U18222 (N_18222,N_17747,N_17862);
nor U18223 (N_18223,N_17833,N_17925);
and U18224 (N_18224,N_17983,N_17901);
xnor U18225 (N_18225,N_17826,N_17820);
nor U18226 (N_18226,N_17983,N_17784);
or U18227 (N_18227,N_17938,N_17835);
or U18228 (N_18228,N_17732,N_17892);
nor U18229 (N_18229,N_17972,N_17814);
nand U18230 (N_18230,N_17757,N_17879);
or U18231 (N_18231,N_17812,N_17825);
nor U18232 (N_18232,N_17766,N_17969);
or U18233 (N_18233,N_17975,N_17934);
xnor U18234 (N_18234,N_17744,N_17790);
or U18235 (N_18235,N_17995,N_17790);
or U18236 (N_18236,N_17748,N_17995);
xor U18237 (N_18237,N_17769,N_17753);
nand U18238 (N_18238,N_17730,N_17906);
nor U18239 (N_18239,N_17790,N_17978);
nand U18240 (N_18240,N_17972,N_17924);
nor U18241 (N_18241,N_17779,N_17783);
xnor U18242 (N_18242,N_17854,N_17983);
or U18243 (N_18243,N_17790,N_17786);
nand U18244 (N_18244,N_17756,N_17788);
nor U18245 (N_18245,N_17872,N_17751);
or U18246 (N_18246,N_17786,N_17953);
xnor U18247 (N_18247,N_17814,N_17712);
nand U18248 (N_18248,N_17890,N_17721);
nor U18249 (N_18249,N_17874,N_17893);
nor U18250 (N_18250,N_17727,N_17757);
xnor U18251 (N_18251,N_17916,N_17860);
and U18252 (N_18252,N_17947,N_17893);
or U18253 (N_18253,N_17722,N_17856);
nor U18254 (N_18254,N_17960,N_17971);
nor U18255 (N_18255,N_17908,N_17876);
nand U18256 (N_18256,N_17919,N_17948);
and U18257 (N_18257,N_17945,N_17883);
xnor U18258 (N_18258,N_17997,N_17743);
xnor U18259 (N_18259,N_17923,N_17802);
nand U18260 (N_18260,N_17993,N_17867);
nor U18261 (N_18261,N_17885,N_17878);
nor U18262 (N_18262,N_17802,N_17871);
nand U18263 (N_18263,N_17932,N_17847);
nor U18264 (N_18264,N_17744,N_17785);
and U18265 (N_18265,N_17803,N_17970);
and U18266 (N_18266,N_17947,N_17734);
nor U18267 (N_18267,N_17883,N_17772);
xnor U18268 (N_18268,N_17883,N_17779);
nand U18269 (N_18269,N_17992,N_17710);
and U18270 (N_18270,N_17760,N_17813);
xor U18271 (N_18271,N_17749,N_17863);
nand U18272 (N_18272,N_17830,N_17968);
or U18273 (N_18273,N_17788,N_17819);
or U18274 (N_18274,N_17734,N_17919);
or U18275 (N_18275,N_17723,N_17867);
nand U18276 (N_18276,N_17780,N_17808);
or U18277 (N_18277,N_17819,N_17811);
or U18278 (N_18278,N_17793,N_17827);
nor U18279 (N_18279,N_17964,N_17897);
and U18280 (N_18280,N_17931,N_17745);
xor U18281 (N_18281,N_17759,N_17837);
and U18282 (N_18282,N_17772,N_17715);
and U18283 (N_18283,N_17761,N_17806);
nor U18284 (N_18284,N_17803,N_17799);
or U18285 (N_18285,N_17785,N_17953);
and U18286 (N_18286,N_17877,N_17842);
or U18287 (N_18287,N_17745,N_17860);
or U18288 (N_18288,N_17878,N_17806);
nand U18289 (N_18289,N_17754,N_17800);
xor U18290 (N_18290,N_17709,N_17795);
xor U18291 (N_18291,N_17820,N_17973);
xnor U18292 (N_18292,N_17876,N_17849);
or U18293 (N_18293,N_17707,N_17762);
or U18294 (N_18294,N_17793,N_17953);
nand U18295 (N_18295,N_17713,N_17844);
and U18296 (N_18296,N_17919,N_17868);
xor U18297 (N_18297,N_17945,N_17753);
xnor U18298 (N_18298,N_17874,N_17737);
nor U18299 (N_18299,N_17723,N_17738);
xnor U18300 (N_18300,N_18169,N_18112);
and U18301 (N_18301,N_18058,N_18289);
nand U18302 (N_18302,N_18168,N_18023);
nor U18303 (N_18303,N_18283,N_18294);
and U18304 (N_18304,N_18115,N_18074);
nand U18305 (N_18305,N_18253,N_18025);
or U18306 (N_18306,N_18237,N_18203);
nand U18307 (N_18307,N_18089,N_18245);
and U18308 (N_18308,N_18222,N_18062);
nand U18309 (N_18309,N_18265,N_18093);
or U18310 (N_18310,N_18045,N_18269);
nand U18311 (N_18311,N_18220,N_18207);
and U18312 (N_18312,N_18039,N_18102);
nand U18313 (N_18313,N_18216,N_18208);
xnor U18314 (N_18314,N_18183,N_18202);
nor U18315 (N_18315,N_18179,N_18196);
nor U18316 (N_18316,N_18091,N_18204);
xnor U18317 (N_18317,N_18211,N_18221);
and U18318 (N_18318,N_18188,N_18037);
and U18319 (N_18319,N_18078,N_18248);
nand U18320 (N_18320,N_18227,N_18218);
and U18321 (N_18321,N_18012,N_18212);
nor U18322 (N_18322,N_18247,N_18228);
nor U18323 (N_18323,N_18288,N_18138);
and U18324 (N_18324,N_18159,N_18182);
nand U18325 (N_18325,N_18139,N_18027);
and U18326 (N_18326,N_18140,N_18034);
or U18327 (N_18327,N_18243,N_18256);
nor U18328 (N_18328,N_18297,N_18080);
nor U18329 (N_18329,N_18121,N_18290);
nand U18330 (N_18330,N_18123,N_18257);
or U18331 (N_18331,N_18061,N_18068);
or U18332 (N_18332,N_18184,N_18049);
nand U18333 (N_18333,N_18164,N_18242);
xnor U18334 (N_18334,N_18051,N_18010);
and U18335 (N_18335,N_18065,N_18109);
or U18336 (N_18336,N_18022,N_18153);
xnor U18337 (N_18337,N_18124,N_18266);
and U18338 (N_18338,N_18152,N_18235);
or U18339 (N_18339,N_18285,N_18090);
or U18340 (N_18340,N_18261,N_18254);
or U18341 (N_18341,N_18021,N_18007);
nor U18342 (N_18342,N_18190,N_18251);
and U18343 (N_18343,N_18125,N_18267);
xor U18344 (N_18344,N_18018,N_18055);
and U18345 (N_18345,N_18250,N_18126);
xnor U18346 (N_18346,N_18154,N_18157);
nor U18347 (N_18347,N_18214,N_18099);
nor U18348 (N_18348,N_18083,N_18128);
or U18349 (N_18349,N_18239,N_18009);
nor U18350 (N_18350,N_18244,N_18024);
nand U18351 (N_18351,N_18141,N_18086);
xnor U18352 (N_18352,N_18110,N_18199);
and U18353 (N_18353,N_18017,N_18031);
nor U18354 (N_18354,N_18277,N_18134);
or U18355 (N_18355,N_18287,N_18286);
nor U18356 (N_18356,N_18100,N_18142);
nor U18357 (N_18357,N_18193,N_18106);
nand U18358 (N_18358,N_18215,N_18172);
xnor U18359 (N_18359,N_18019,N_18231);
nor U18360 (N_18360,N_18206,N_18298);
nand U18361 (N_18361,N_18054,N_18129);
nor U18362 (N_18362,N_18132,N_18013);
and U18363 (N_18363,N_18276,N_18291);
nor U18364 (N_18364,N_18205,N_18226);
or U18365 (N_18365,N_18005,N_18028);
and U18366 (N_18366,N_18175,N_18263);
and U18367 (N_18367,N_18252,N_18071);
nor U18368 (N_18368,N_18150,N_18198);
or U18369 (N_18369,N_18158,N_18066);
nand U18370 (N_18370,N_18120,N_18292);
nand U18371 (N_18371,N_18281,N_18200);
nand U18372 (N_18372,N_18060,N_18044);
nor U18373 (N_18373,N_18056,N_18187);
nor U18374 (N_18374,N_18166,N_18082);
nor U18375 (N_18375,N_18149,N_18156);
and U18376 (N_18376,N_18032,N_18059);
xnor U18377 (N_18377,N_18095,N_18224);
and U18378 (N_18378,N_18186,N_18042);
xnor U18379 (N_18379,N_18050,N_18163);
nand U18380 (N_18380,N_18268,N_18053);
or U18381 (N_18381,N_18209,N_18127);
nor U18382 (N_18382,N_18085,N_18043);
or U18383 (N_18383,N_18113,N_18104);
and U18384 (N_18384,N_18195,N_18006);
nand U18385 (N_18385,N_18219,N_18170);
or U18386 (N_18386,N_18236,N_18026);
xor U18387 (N_18387,N_18016,N_18255);
or U18388 (N_18388,N_18197,N_18264);
xnor U18389 (N_18389,N_18008,N_18155);
nand U18390 (N_18390,N_18259,N_18035);
nor U18391 (N_18391,N_18114,N_18118);
or U18392 (N_18392,N_18029,N_18246);
or U18393 (N_18393,N_18020,N_18223);
nand U18394 (N_18394,N_18122,N_18015);
or U18395 (N_18395,N_18213,N_18096);
xor U18396 (N_18396,N_18030,N_18052);
xnor U18397 (N_18397,N_18238,N_18194);
xnor U18398 (N_18398,N_18135,N_18084);
nor U18399 (N_18399,N_18041,N_18143);
xor U18400 (N_18400,N_18262,N_18145);
nand U18401 (N_18401,N_18040,N_18076);
xnor U18402 (N_18402,N_18271,N_18144);
and U18403 (N_18403,N_18240,N_18185);
nor U18404 (N_18404,N_18160,N_18148);
nor U18405 (N_18405,N_18210,N_18282);
xor U18406 (N_18406,N_18070,N_18130);
or U18407 (N_18407,N_18072,N_18270);
nor U18408 (N_18408,N_18284,N_18087);
xnor U18409 (N_18409,N_18181,N_18036);
xnor U18410 (N_18410,N_18094,N_18162);
xnor U18411 (N_18411,N_18098,N_18002);
nand U18412 (N_18412,N_18161,N_18146);
and U18413 (N_18413,N_18000,N_18151);
and U18414 (N_18414,N_18137,N_18105);
nor U18415 (N_18415,N_18003,N_18225);
and U18416 (N_18416,N_18189,N_18001);
nand U18417 (N_18417,N_18230,N_18064);
xnor U18418 (N_18418,N_18275,N_18131);
or U18419 (N_18419,N_18295,N_18077);
and U18420 (N_18420,N_18278,N_18279);
xnor U18421 (N_18421,N_18101,N_18191);
nor U18422 (N_18422,N_18046,N_18119);
nand U18423 (N_18423,N_18073,N_18232);
nand U18424 (N_18424,N_18047,N_18063);
nand U18425 (N_18425,N_18081,N_18011);
nand U18426 (N_18426,N_18293,N_18079);
xnor U18427 (N_18427,N_18241,N_18177);
xor U18428 (N_18428,N_18116,N_18180);
and U18429 (N_18429,N_18108,N_18249);
nand U18430 (N_18430,N_18107,N_18069);
nor U18431 (N_18431,N_18103,N_18234);
and U18432 (N_18432,N_18057,N_18097);
nand U18433 (N_18433,N_18038,N_18192);
and U18434 (N_18434,N_18174,N_18167);
nand U18435 (N_18435,N_18147,N_18260);
nor U18436 (N_18436,N_18173,N_18176);
xor U18437 (N_18437,N_18296,N_18299);
and U18438 (N_18438,N_18033,N_18067);
or U18439 (N_18439,N_18178,N_18092);
xnor U18440 (N_18440,N_18111,N_18075);
nor U18441 (N_18441,N_18117,N_18014);
nand U18442 (N_18442,N_18273,N_18136);
nor U18443 (N_18443,N_18274,N_18217);
nor U18444 (N_18444,N_18004,N_18280);
xnor U18445 (N_18445,N_18171,N_18229);
or U18446 (N_18446,N_18048,N_18201);
and U18447 (N_18447,N_18165,N_18088);
and U18448 (N_18448,N_18258,N_18233);
nor U18449 (N_18449,N_18133,N_18272);
and U18450 (N_18450,N_18070,N_18255);
nor U18451 (N_18451,N_18097,N_18068);
nor U18452 (N_18452,N_18223,N_18236);
and U18453 (N_18453,N_18157,N_18071);
xnor U18454 (N_18454,N_18105,N_18016);
or U18455 (N_18455,N_18171,N_18210);
and U18456 (N_18456,N_18285,N_18200);
nand U18457 (N_18457,N_18163,N_18237);
nor U18458 (N_18458,N_18252,N_18029);
or U18459 (N_18459,N_18297,N_18251);
xnor U18460 (N_18460,N_18092,N_18132);
or U18461 (N_18461,N_18290,N_18265);
and U18462 (N_18462,N_18001,N_18019);
nand U18463 (N_18463,N_18011,N_18217);
or U18464 (N_18464,N_18103,N_18106);
or U18465 (N_18465,N_18280,N_18178);
xor U18466 (N_18466,N_18292,N_18280);
xnor U18467 (N_18467,N_18133,N_18176);
nor U18468 (N_18468,N_18159,N_18110);
or U18469 (N_18469,N_18261,N_18207);
or U18470 (N_18470,N_18061,N_18197);
xor U18471 (N_18471,N_18030,N_18017);
or U18472 (N_18472,N_18235,N_18144);
or U18473 (N_18473,N_18063,N_18169);
nand U18474 (N_18474,N_18013,N_18019);
nor U18475 (N_18475,N_18159,N_18262);
and U18476 (N_18476,N_18188,N_18002);
and U18477 (N_18477,N_18223,N_18047);
and U18478 (N_18478,N_18173,N_18219);
or U18479 (N_18479,N_18073,N_18122);
nor U18480 (N_18480,N_18004,N_18283);
and U18481 (N_18481,N_18165,N_18286);
or U18482 (N_18482,N_18036,N_18250);
nand U18483 (N_18483,N_18149,N_18069);
or U18484 (N_18484,N_18293,N_18286);
and U18485 (N_18485,N_18151,N_18207);
and U18486 (N_18486,N_18008,N_18276);
or U18487 (N_18487,N_18167,N_18020);
and U18488 (N_18488,N_18069,N_18158);
nor U18489 (N_18489,N_18069,N_18265);
or U18490 (N_18490,N_18190,N_18116);
and U18491 (N_18491,N_18236,N_18158);
xor U18492 (N_18492,N_18073,N_18224);
nor U18493 (N_18493,N_18036,N_18234);
nor U18494 (N_18494,N_18191,N_18161);
or U18495 (N_18495,N_18010,N_18216);
and U18496 (N_18496,N_18017,N_18033);
nand U18497 (N_18497,N_18264,N_18093);
and U18498 (N_18498,N_18279,N_18079);
or U18499 (N_18499,N_18086,N_18053);
nor U18500 (N_18500,N_18188,N_18166);
nor U18501 (N_18501,N_18187,N_18118);
or U18502 (N_18502,N_18137,N_18214);
xor U18503 (N_18503,N_18219,N_18186);
or U18504 (N_18504,N_18026,N_18232);
xor U18505 (N_18505,N_18141,N_18171);
or U18506 (N_18506,N_18213,N_18199);
nand U18507 (N_18507,N_18079,N_18221);
and U18508 (N_18508,N_18247,N_18192);
or U18509 (N_18509,N_18285,N_18150);
xor U18510 (N_18510,N_18285,N_18058);
nand U18511 (N_18511,N_18211,N_18184);
or U18512 (N_18512,N_18047,N_18236);
xor U18513 (N_18513,N_18103,N_18054);
nor U18514 (N_18514,N_18066,N_18027);
xnor U18515 (N_18515,N_18169,N_18082);
nand U18516 (N_18516,N_18171,N_18218);
or U18517 (N_18517,N_18132,N_18024);
and U18518 (N_18518,N_18298,N_18264);
nor U18519 (N_18519,N_18163,N_18055);
and U18520 (N_18520,N_18105,N_18172);
or U18521 (N_18521,N_18139,N_18273);
or U18522 (N_18522,N_18108,N_18232);
or U18523 (N_18523,N_18176,N_18036);
and U18524 (N_18524,N_18124,N_18200);
and U18525 (N_18525,N_18136,N_18214);
nor U18526 (N_18526,N_18038,N_18240);
xor U18527 (N_18527,N_18255,N_18116);
nand U18528 (N_18528,N_18191,N_18026);
xor U18529 (N_18529,N_18065,N_18112);
xor U18530 (N_18530,N_18263,N_18183);
nand U18531 (N_18531,N_18121,N_18062);
nor U18532 (N_18532,N_18121,N_18131);
nor U18533 (N_18533,N_18181,N_18179);
or U18534 (N_18534,N_18215,N_18273);
nor U18535 (N_18535,N_18038,N_18207);
or U18536 (N_18536,N_18239,N_18187);
nor U18537 (N_18537,N_18108,N_18088);
or U18538 (N_18538,N_18283,N_18081);
nor U18539 (N_18539,N_18159,N_18065);
xnor U18540 (N_18540,N_18067,N_18000);
xnor U18541 (N_18541,N_18126,N_18056);
and U18542 (N_18542,N_18293,N_18172);
and U18543 (N_18543,N_18129,N_18137);
or U18544 (N_18544,N_18108,N_18125);
or U18545 (N_18545,N_18157,N_18198);
or U18546 (N_18546,N_18287,N_18102);
nand U18547 (N_18547,N_18124,N_18226);
and U18548 (N_18548,N_18029,N_18121);
nand U18549 (N_18549,N_18212,N_18245);
nand U18550 (N_18550,N_18052,N_18210);
nor U18551 (N_18551,N_18143,N_18193);
nor U18552 (N_18552,N_18078,N_18175);
and U18553 (N_18553,N_18041,N_18168);
xor U18554 (N_18554,N_18265,N_18116);
or U18555 (N_18555,N_18051,N_18050);
nor U18556 (N_18556,N_18224,N_18067);
and U18557 (N_18557,N_18025,N_18281);
nor U18558 (N_18558,N_18124,N_18167);
xnor U18559 (N_18559,N_18253,N_18143);
nor U18560 (N_18560,N_18059,N_18049);
or U18561 (N_18561,N_18075,N_18190);
and U18562 (N_18562,N_18105,N_18194);
and U18563 (N_18563,N_18002,N_18199);
nand U18564 (N_18564,N_18012,N_18188);
nand U18565 (N_18565,N_18136,N_18244);
and U18566 (N_18566,N_18299,N_18059);
xor U18567 (N_18567,N_18024,N_18124);
nor U18568 (N_18568,N_18205,N_18220);
nor U18569 (N_18569,N_18297,N_18126);
xor U18570 (N_18570,N_18072,N_18207);
or U18571 (N_18571,N_18147,N_18005);
nand U18572 (N_18572,N_18140,N_18132);
and U18573 (N_18573,N_18047,N_18278);
or U18574 (N_18574,N_18014,N_18277);
xnor U18575 (N_18575,N_18159,N_18149);
and U18576 (N_18576,N_18235,N_18243);
xnor U18577 (N_18577,N_18061,N_18111);
nor U18578 (N_18578,N_18162,N_18000);
xor U18579 (N_18579,N_18011,N_18098);
xor U18580 (N_18580,N_18189,N_18261);
or U18581 (N_18581,N_18233,N_18031);
and U18582 (N_18582,N_18092,N_18056);
xor U18583 (N_18583,N_18153,N_18267);
and U18584 (N_18584,N_18135,N_18059);
and U18585 (N_18585,N_18166,N_18251);
and U18586 (N_18586,N_18238,N_18089);
xnor U18587 (N_18587,N_18070,N_18031);
nor U18588 (N_18588,N_18150,N_18033);
and U18589 (N_18589,N_18119,N_18203);
xnor U18590 (N_18590,N_18116,N_18097);
or U18591 (N_18591,N_18047,N_18064);
and U18592 (N_18592,N_18295,N_18059);
or U18593 (N_18593,N_18048,N_18234);
xor U18594 (N_18594,N_18040,N_18057);
and U18595 (N_18595,N_18249,N_18005);
xnor U18596 (N_18596,N_18282,N_18114);
xor U18597 (N_18597,N_18166,N_18299);
nand U18598 (N_18598,N_18008,N_18270);
xor U18599 (N_18599,N_18238,N_18003);
or U18600 (N_18600,N_18516,N_18495);
nor U18601 (N_18601,N_18552,N_18592);
and U18602 (N_18602,N_18341,N_18308);
or U18603 (N_18603,N_18486,N_18527);
and U18604 (N_18604,N_18358,N_18304);
and U18605 (N_18605,N_18500,N_18441);
nand U18606 (N_18606,N_18593,N_18589);
or U18607 (N_18607,N_18459,N_18565);
nand U18608 (N_18608,N_18581,N_18555);
xor U18609 (N_18609,N_18519,N_18368);
and U18610 (N_18610,N_18361,N_18594);
or U18611 (N_18611,N_18417,N_18549);
nor U18612 (N_18612,N_18513,N_18332);
and U18613 (N_18613,N_18445,N_18585);
or U18614 (N_18614,N_18406,N_18442);
xnor U18615 (N_18615,N_18437,N_18520);
and U18616 (N_18616,N_18376,N_18498);
nor U18617 (N_18617,N_18384,N_18321);
xnor U18618 (N_18618,N_18313,N_18398);
and U18619 (N_18619,N_18464,N_18562);
and U18620 (N_18620,N_18378,N_18590);
and U18621 (N_18621,N_18392,N_18523);
xnor U18622 (N_18622,N_18506,N_18472);
nor U18623 (N_18623,N_18456,N_18521);
xor U18624 (N_18624,N_18305,N_18533);
nor U18625 (N_18625,N_18360,N_18333);
and U18626 (N_18626,N_18372,N_18393);
and U18627 (N_18627,N_18318,N_18310);
and U18628 (N_18628,N_18543,N_18388);
xnor U18629 (N_18629,N_18435,N_18327);
nor U18630 (N_18630,N_18535,N_18390);
nor U18631 (N_18631,N_18400,N_18381);
or U18632 (N_18632,N_18503,N_18575);
and U18633 (N_18633,N_18402,N_18343);
and U18634 (N_18634,N_18307,N_18349);
or U18635 (N_18635,N_18496,N_18499);
nand U18636 (N_18636,N_18342,N_18509);
and U18637 (N_18637,N_18493,N_18426);
nor U18638 (N_18638,N_18556,N_18409);
xnor U18639 (N_18639,N_18473,N_18316);
or U18640 (N_18640,N_18576,N_18548);
nor U18641 (N_18641,N_18557,N_18454);
nor U18642 (N_18642,N_18553,N_18383);
nor U18643 (N_18643,N_18465,N_18466);
and U18644 (N_18644,N_18369,N_18540);
and U18645 (N_18645,N_18325,N_18320);
nor U18646 (N_18646,N_18571,N_18559);
nand U18647 (N_18647,N_18582,N_18515);
or U18648 (N_18648,N_18474,N_18362);
nand U18649 (N_18649,N_18319,N_18531);
nand U18650 (N_18650,N_18444,N_18455);
nor U18651 (N_18651,N_18309,N_18588);
xor U18652 (N_18652,N_18526,N_18580);
nand U18653 (N_18653,N_18522,N_18447);
nand U18654 (N_18654,N_18364,N_18414);
xor U18655 (N_18655,N_18431,N_18355);
nand U18656 (N_18656,N_18598,N_18487);
xnor U18657 (N_18657,N_18363,N_18468);
xor U18658 (N_18658,N_18301,N_18488);
xor U18659 (N_18659,N_18425,N_18389);
nor U18660 (N_18660,N_18380,N_18353);
or U18661 (N_18661,N_18429,N_18405);
xor U18662 (N_18662,N_18373,N_18587);
xnor U18663 (N_18663,N_18412,N_18475);
nor U18664 (N_18664,N_18415,N_18458);
nor U18665 (N_18665,N_18323,N_18401);
or U18666 (N_18666,N_18558,N_18334);
nor U18667 (N_18667,N_18314,N_18397);
or U18668 (N_18668,N_18322,N_18326);
nand U18669 (N_18669,N_18542,N_18583);
xor U18670 (N_18670,N_18422,N_18508);
or U18671 (N_18671,N_18534,N_18382);
xor U18672 (N_18672,N_18324,N_18416);
and U18673 (N_18673,N_18505,N_18430);
nor U18674 (N_18674,N_18492,N_18586);
or U18675 (N_18675,N_18504,N_18350);
xor U18676 (N_18676,N_18428,N_18410);
or U18677 (N_18677,N_18329,N_18331);
nand U18678 (N_18678,N_18566,N_18423);
or U18679 (N_18679,N_18467,N_18420);
or U18680 (N_18680,N_18524,N_18356);
nor U18681 (N_18681,N_18525,N_18352);
and U18682 (N_18682,N_18469,N_18407);
nor U18683 (N_18683,N_18339,N_18532);
and U18684 (N_18684,N_18462,N_18501);
and U18685 (N_18685,N_18411,N_18460);
nor U18686 (N_18686,N_18560,N_18510);
nor U18687 (N_18687,N_18529,N_18507);
or U18688 (N_18688,N_18391,N_18591);
nand U18689 (N_18689,N_18317,N_18367);
nand U18690 (N_18690,N_18537,N_18547);
or U18691 (N_18691,N_18545,N_18370);
xnor U18692 (N_18692,N_18551,N_18311);
and U18693 (N_18693,N_18306,N_18427);
and U18694 (N_18694,N_18491,N_18479);
xor U18695 (N_18695,N_18345,N_18359);
nand U18696 (N_18696,N_18568,N_18517);
nand U18697 (N_18697,N_18448,N_18315);
nor U18698 (N_18698,N_18578,N_18434);
nor U18699 (N_18699,N_18512,N_18481);
xnor U18700 (N_18700,N_18336,N_18574);
xor U18701 (N_18701,N_18340,N_18569);
or U18702 (N_18702,N_18584,N_18404);
and U18703 (N_18703,N_18597,N_18436);
and U18704 (N_18704,N_18312,N_18482);
xor U18705 (N_18705,N_18302,N_18446);
nor U18706 (N_18706,N_18335,N_18375);
nor U18707 (N_18707,N_18573,N_18348);
nand U18708 (N_18708,N_18449,N_18502);
and U18709 (N_18709,N_18403,N_18344);
xnor U18710 (N_18710,N_18300,N_18563);
and U18711 (N_18711,N_18366,N_18528);
nor U18712 (N_18712,N_18541,N_18419);
and U18713 (N_18713,N_18424,N_18470);
and U18714 (N_18714,N_18579,N_18347);
xnor U18715 (N_18715,N_18377,N_18386);
and U18716 (N_18716,N_18371,N_18354);
nand U18717 (N_18717,N_18440,N_18554);
nand U18718 (N_18718,N_18599,N_18478);
nor U18719 (N_18719,N_18439,N_18570);
nand U18720 (N_18720,N_18489,N_18539);
or U18721 (N_18721,N_18453,N_18595);
xor U18722 (N_18722,N_18561,N_18572);
nand U18723 (N_18723,N_18408,N_18418);
xnor U18724 (N_18724,N_18538,N_18577);
and U18725 (N_18725,N_18374,N_18365);
xor U18726 (N_18726,N_18399,N_18596);
nor U18727 (N_18727,N_18484,N_18396);
nand U18728 (N_18728,N_18536,N_18338);
xor U18729 (N_18729,N_18511,N_18346);
xnor U18730 (N_18730,N_18357,N_18483);
nand U18731 (N_18731,N_18463,N_18413);
xnor U18732 (N_18732,N_18546,N_18450);
nor U18733 (N_18733,N_18451,N_18485);
nor U18734 (N_18734,N_18476,N_18457);
or U18735 (N_18735,N_18550,N_18395);
nand U18736 (N_18736,N_18452,N_18494);
or U18737 (N_18737,N_18303,N_18330);
xor U18738 (N_18738,N_18544,N_18564);
xnor U18739 (N_18739,N_18394,N_18461);
nor U18740 (N_18740,N_18328,N_18490);
and U18741 (N_18741,N_18432,N_18518);
nand U18742 (N_18742,N_18567,N_18337);
nor U18743 (N_18743,N_18443,N_18433);
xor U18744 (N_18744,N_18385,N_18438);
xor U18745 (N_18745,N_18471,N_18421);
xor U18746 (N_18746,N_18477,N_18530);
or U18747 (N_18747,N_18480,N_18379);
and U18748 (N_18748,N_18497,N_18387);
and U18749 (N_18749,N_18351,N_18514);
nor U18750 (N_18750,N_18333,N_18436);
nor U18751 (N_18751,N_18466,N_18412);
nor U18752 (N_18752,N_18587,N_18337);
nor U18753 (N_18753,N_18355,N_18554);
or U18754 (N_18754,N_18346,N_18556);
nand U18755 (N_18755,N_18457,N_18430);
xnor U18756 (N_18756,N_18437,N_18339);
or U18757 (N_18757,N_18536,N_18589);
and U18758 (N_18758,N_18388,N_18441);
and U18759 (N_18759,N_18576,N_18368);
and U18760 (N_18760,N_18372,N_18530);
or U18761 (N_18761,N_18556,N_18306);
xor U18762 (N_18762,N_18589,N_18594);
and U18763 (N_18763,N_18517,N_18562);
nand U18764 (N_18764,N_18327,N_18306);
nand U18765 (N_18765,N_18411,N_18347);
xor U18766 (N_18766,N_18434,N_18320);
or U18767 (N_18767,N_18411,N_18378);
nand U18768 (N_18768,N_18350,N_18576);
and U18769 (N_18769,N_18407,N_18565);
nand U18770 (N_18770,N_18544,N_18301);
nand U18771 (N_18771,N_18316,N_18529);
and U18772 (N_18772,N_18535,N_18588);
xor U18773 (N_18773,N_18494,N_18425);
xnor U18774 (N_18774,N_18423,N_18526);
and U18775 (N_18775,N_18350,N_18359);
or U18776 (N_18776,N_18545,N_18382);
nor U18777 (N_18777,N_18459,N_18474);
nand U18778 (N_18778,N_18336,N_18463);
nand U18779 (N_18779,N_18563,N_18475);
or U18780 (N_18780,N_18457,N_18586);
xnor U18781 (N_18781,N_18313,N_18339);
or U18782 (N_18782,N_18546,N_18421);
or U18783 (N_18783,N_18469,N_18321);
xnor U18784 (N_18784,N_18598,N_18512);
or U18785 (N_18785,N_18366,N_18468);
nor U18786 (N_18786,N_18369,N_18451);
nand U18787 (N_18787,N_18399,N_18473);
xor U18788 (N_18788,N_18428,N_18324);
or U18789 (N_18789,N_18582,N_18398);
nand U18790 (N_18790,N_18336,N_18537);
or U18791 (N_18791,N_18372,N_18361);
nand U18792 (N_18792,N_18388,N_18529);
and U18793 (N_18793,N_18399,N_18594);
and U18794 (N_18794,N_18450,N_18309);
or U18795 (N_18795,N_18365,N_18521);
and U18796 (N_18796,N_18554,N_18514);
xnor U18797 (N_18797,N_18563,N_18516);
or U18798 (N_18798,N_18446,N_18445);
xnor U18799 (N_18799,N_18347,N_18374);
nand U18800 (N_18800,N_18529,N_18555);
nor U18801 (N_18801,N_18597,N_18416);
or U18802 (N_18802,N_18429,N_18574);
nor U18803 (N_18803,N_18363,N_18460);
or U18804 (N_18804,N_18336,N_18307);
nor U18805 (N_18805,N_18446,N_18591);
nor U18806 (N_18806,N_18512,N_18421);
and U18807 (N_18807,N_18470,N_18441);
nor U18808 (N_18808,N_18419,N_18568);
or U18809 (N_18809,N_18594,N_18301);
nor U18810 (N_18810,N_18576,N_18412);
xor U18811 (N_18811,N_18478,N_18431);
nand U18812 (N_18812,N_18447,N_18431);
nor U18813 (N_18813,N_18408,N_18395);
xor U18814 (N_18814,N_18389,N_18443);
nor U18815 (N_18815,N_18392,N_18573);
xnor U18816 (N_18816,N_18566,N_18550);
nor U18817 (N_18817,N_18477,N_18408);
or U18818 (N_18818,N_18344,N_18380);
nand U18819 (N_18819,N_18599,N_18431);
and U18820 (N_18820,N_18514,N_18556);
and U18821 (N_18821,N_18578,N_18584);
or U18822 (N_18822,N_18358,N_18329);
nand U18823 (N_18823,N_18598,N_18559);
xor U18824 (N_18824,N_18426,N_18328);
or U18825 (N_18825,N_18492,N_18479);
and U18826 (N_18826,N_18553,N_18535);
and U18827 (N_18827,N_18598,N_18531);
or U18828 (N_18828,N_18329,N_18412);
and U18829 (N_18829,N_18478,N_18319);
nand U18830 (N_18830,N_18594,N_18471);
nand U18831 (N_18831,N_18506,N_18560);
or U18832 (N_18832,N_18537,N_18530);
or U18833 (N_18833,N_18452,N_18417);
nand U18834 (N_18834,N_18555,N_18340);
xor U18835 (N_18835,N_18543,N_18486);
or U18836 (N_18836,N_18381,N_18593);
or U18837 (N_18837,N_18305,N_18350);
and U18838 (N_18838,N_18500,N_18439);
nor U18839 (N_18839,N_18434,N_18319);
and U18840 (N_18840,N_18542,N_18469);
or U18841 (N_18841,N_18399,N_18560);
nand U18842 (N_18842,N_18494,N_18348);
nand U18843 (N_18843,N_18599,N_18400);
nand U18844 (N_18844,N_18336,N_18354);
nand U18845 (N_18845,N_18392,N_18452);
or U18846 (N_18846,N_18479,N_18455);
nor U18847 (N_18847,N_18493,N_18327);
and U18848 (N_18848,N_18414,N_18431);
xor U18849 (N_18849,N_18499,N_18434);
nand U18850 (N_18850,N_18392,N_18463);
nor U18851 (N_18851,N_18426,N_18507);
nand U18852 (N_18852,N_18524,N_18519);
xor U18853 (N_18853,N_18522,N_18353);
and U18854 (N_18854,N_18380,N_18524);
nor U18855 (N_18855,N_18564,N_18458);
and U18856 (N_18856,N_18409,N_18413);
and U18857 (N_18857,N_18328,N_18553);
nand U18858 (N_18858,N_18526,N_18309);
nor U18859 (N_18859,N_18321,N_18421);
or U18860 (N_18860,N_18302,N_18414);
nor U18861 (N_18861,N_18376,N_18494);
or U18862 (N_18862,N_18483,N_18428);
xor U18863 (N_18863,N_18393,N_18503);
xor U18864 (N_18864,N_18565,N_18306);
nand U18865 (N_18865,N_18554,N_18380);
or U18866 (N_18866,N_18568,N_18324);
nand U18867 (N_18867,N_18379,N_18559);
and U18868 (N_18868,N_18496,N_18436);
xor U18869 (N_18869,N_18490,N_18408);
nor U18870 (N_18870,N_18517,N_18309);
xor U18871 (N_18871,N_18351,N_18520);
xor U18872 (N_18872,N_18441,N_18565);
nand U18873 (N_18873,N_18454,N_18401);
and U18874 (N_18874,N_18522,N_18529);
and U18875 (N_18875,N_18397,N_18596);
nand U18876 (N_18876,N_18534,N_18414);
and U18877 (N_18877,N_18385,N_18509);
xnor U18878 (N_18878,N_18381,N_18453);
xor U18879 (N_18879,N_18504,N_18471);
nor U18880 (N_18880,N_18324,N_18453);
nor U18881 (N_18881,N_18398,N_18532);
and U18882 (N_18882,N_18312,N_18501);
nand U18883 (N_18883,N_18551,N_18512);
and U18884 (N_18884,N_18308,N_18481);
or U18885 (N_18885,N_18319,N_18442);
and U18886 (N_18886,N_18534,N_18545);
nor U18887 (N_18887,N_18579,N_18355);
and U18888 (N_18888,N_18475,N_18496);
xor U18889 (N_18889,N_18430,N_18321);
and U18890 (N_18890,N_18457,N_18596);
nor U18891 (N_18891,N_18481,N_18492);
or U18892 (N_18892,N_18337,N_18305);
xnor U18893 (N_18893,N_18405,N_18448);
nand U18894 (N_18894,N_18358,N_18453);
or U18895 (N_18895,N_18416,N_18303);
nand U18896 (N_18896,N_18317,N_18486);
or U18897 (N_18897,N_18391,N_18447);
or U18898 (N_18898,N_18585,N_18554);
nor U18899 (N_18899,N_18491,N_18437);
or U18900 (N_18900,N_18775,N_18727);
nand U18901 (N_18901,N_18711,N_18875);
xnor U18902 (N_18902,N_18826,N_18676);
and U18903 (N_18903,N_18600,N_18822);
nand U18904 (N_18904,N_18809,N_18800);
nor U18905 (N_18905,N_18625,N_18607);
nand U18906 (N_18906,N_18665,N_18740);
xnor U18907 (N_18907,N_18698,N_18797);
or U18908 (N_18908,N_18758,N_18679);
nand U18909 (N_18909,N_18692,N_18861);
xnor U18910 (N_18910,N_18680,N_18833);
nor U18911 (N_18911,N_18793,N_18883);
xnor U18912 (N_18912,N_18851,N_18701);
nor U18913 (N_18913,N_18706,N_18648);
and U18914 (N_18914,N_18777,N_18848);
or U18915 (N_18915,N_18629,N_18613);
nor U18916 (N_18916,N_18622,N_18685);
xor U18917 (N_18917,N_18879,N_18788);
and U18918 (N_18918,N_18650,N_18745);
nand U18919 (N_18919,N_18694,N_18762);
nand U18920 (N_18920,N_18636,N_18877);
xnor U18921 (N_18921,N_18691,N_18749);
nor U18922 (N_18922,N_18730,N_18836);
nand U18923 (N_18923,N_18683,N_18859);
xor U18924 (N_18924,N_18881,N_18667);
and U18925 (N_18925,N_18601,N_18811);
and U18926 (N_18926,N_18778,N_18824);
nand U18927 (N_18927,N_18717,N_18670);
nor U18928 (N_18928,N_18675,N_18885);
nand U18929 (N_18929,N_18684,N_18845);
or U18930 (N_18930,N_18755,N_18729);
nand U18931 (N_18931,N_18723,N_18897);
or U18932 (N_18932,N_18810,N_18825);
and U18933 (N_18933,N_18779,N_18733);
xnor U18934 (N_18934,N_18750,N_18737);
and U18935 (N_18935,N_18724,N_18721);
nand U18936 (N_18936,N_18772,N_18757);
nor U18937 (N_18937,N_18806,N_18850);
and U18938 (N_18938,N_18678,N_18681);
xnor U18939 (N_18939,N_18886,N_18889);
nand U18940 (N_18940,N_18817,N_18686);
xor U18941 (N_18941,N_18774,N_18651);
or U18942 (N_18942,N_18744,N_18865);
xor U18943 (N_18943,N_18888,N_18756);
nand U18944 (N_18944,N_18846,N_18771);
and U18945 (N_18945,N_18635,N_18718);
nand U18946 (N_18946,N_18766,N_18839);
nand U18947 (N_18947,N_18621,N_18747);
or U18948 (N_18948,N_18821,N_18827);
or U18949 (N_18949,N_18633,N_18695);
nand U18950 (N_18950,N_18884,N_18764);
nand U18951 (N_18951,N_18643,N_18853);
xnor U18952 (N_18952,N_18611,N_18672);
and U18953 (N_18953,N_18792,N_18693);
nand U18954 (N_18954,N_18869,N_18807);
or U18955 (N_18955,N_18830,N_18715);
xor U18956 (N_18956,N_18608,N_18834);
nor U18957 (N_18957,N_18702,N_18671);
and U18958 (N_18958,N_18798,N_18838);
nor U18959 (N_18959,N_18871,N_18882);
and U18960 (N_18960,N_18872,N_18713);
and U18961 (N_18961,N_18896,N_18832);
or U18962 (N_18962,N_18634,N_18697);
nand U18963 (N_18963,N_18722,N_18751);
xor U18964 (N_18964,N_18819,N_18725);
nand U18965 (N_18965,N_18782,N_18894);
nand U18966 (N_18966,N_18829,N_18734);
xor U18967 (N_18967,N_18644,N_18786);
xnor U18968 (N_18968,N_18812,N_18780);
nor U18969 (N_18969,N_18761,N_18759);
xnor U18970 (N_18970,N_18743,N_18794);
or U18971 (N_18971,N_18799,N_18620);
nor U18972 (N_18972,N_18820,N_18831);
xor U18973 (N_18973,N_18639,N_18688);
nor U18974 (N_18974,N_18705,N_18791);
and U18975 (N_18975,N_18768,N_18789);
or U18976 (N_18976,N_18752,N_18769);
and U18977 (N_18977,N_18874,N_18728);
and U18978 (N_18978,N_18606,N_18626);
or U18979 (N_18979,N_18887,N_18867);
xor U18980 (N_18980,N_18741,N_18638);
xnor U18981 (N_18981,N_18703,N_18652);
nor U18982 (N_18982,N_18708,N_18632);
or U18983 (N_18983,N_18687,N_18720);
xnor U18984 (N_18984,N_18842,N_18785);
xor U18985 (N_18985,N_18890,N_18815);
and U18986 (N_18986,N_18802,N_18689);
or U18987 (N_18987,N_18712,N_18707);
xor U18988 (N_18988,N_18658,N_18677);
xnor U18989 (N_18989,N_18862,N_18645);
nand U18990 (N_18990,N_18816,N_18619);
nand U18991 (N_18991,N_18837,N_18852);
xnor U18992 (N_18992,N_18790,N_18617);
and U18993 (N_18993,N_18849,N_18637);
nand U18994 (N_18994,N_18795,N_18742);
nand U18995 (N_18995,N_18623,N_18784);
nand U18996 (N_18996,N_18763,N_18714);
and U18997 (N_18997,N_18855,N_18630);
or U18998 (N_18998,N_18628,N_18835);
and U18999 (N_18999,N_18640,N_18893);
xnor U19000 (N_19000,N_18880,N_18863);
xor U19001 (N_19001,N_18878,N_18682);
and U19002 (N_19002,N_18899,N_18719);
and U19003 (N_19003,N_18736,N_18655);
nand U19004 (N_19004,N_18661,N_18843);
xnor U19005 (N_19005,N_18754,N_18814);
or U19006 (N_19006,N_18647,N_18609);
and U19007 (N_19007,N_18716,N_18746);
and U19008 (N_19008,N_18663,N_18892);
and U19009 (N_19009,N_18773,N_18783);
xor U19010 (N_19010,N_18602,N_18760);
nor U19011 (N_19011,N_18840,N_18805);
nand U19012 (N_19012,N_18732,N_18669);
and U19013 (N_19013,N_18738,N_18641);
and U19014 (N_19014,N_18603,N_18656);
xnor U19015 (N_19015,N_18854,N_18646);
or U19016 (N_19016,N_18776,N_18616);
xnor U19017 (N_19017,N_18631,N_18654);
xor U19018 (N_19018,N_18666,N_18624);
xnor U19019 (N_19019,N_18604,N_18813);
nand U19020 (N_19020,N_18748,N_18649);
nor U19021 (N_19021,N_18739,N_18781);
or U19022 (N_19022,N_18858,N_18664);
nand U19023 (N_19023,N_18726,N_18873);
and U19024 (N_19024,N_18808,N_18856);
xnor U19025 (N_19025,N_18699,N_18642);
or U19026 (N_19026,N_18866,N_18731);
nand U19027 (N_19027,N_18767,N_18674);
or U19028 (N_19028,N_18605,N_18787);
nor U19029 (N_19029,N_18660,N_18857);
xnor U19030 (N_19030,N_18659,N_18704);
nand U19031 (N_19031,N_18823,N_18895);
and U19032 (N_19032,N_18898,N_18804);
and U19033 (N_19033,N_18841,N_18735);
nand U19034 (N_19034,N_18627,N_18828);
nand U19035 (N_19035,N_18864,N_18657);
and U19036 (N_19036,N_18868,N_18770);
xor U19037 (N_19037,N_18700,N_18653);
nor U19038 (N_19038,N_18891,N_18673);
or U19039 (N_19039,N_18818,N_18765);
nand U19040 (N_19040,N_18690,N_18615);
nor U19041 (N_19041,N_18610,N_18876);
or U19042 (N_19042,N_18614,N_18612);
or U19043 (N_19043,N_18710,N_18860);
and U19044 (N_19044,N_18668,N_18753);
nor U19045 (N_19045,N_18796,N_18844);
or U19046 (N_19046,N_18696,N_18618);
nand U19047 (N_19047,N_18801,N_18847);
xor U19048 (N_19048,N_18709,N_18803);
nor U19049 (N_19049,N_18662,N_18870);
nand U19050 (N_19050,N_18635,N_18677);
nor U19051 (N_19051,N_18686,N_18816);
xnor U19052 (N_19052,N_18740,N_18660);
nand U19053 (N_19053,N_18617,N_18650);
and U19054 (N_19054,N_18639,N_18883);
nand U19055 (N_19055,N_18766,N_18892);
nor U19056 (N_19056,N_18702,N_18615);
nand U19057 (N_19057,N_18812,N_18795);
or U19058 (N_19058,N_18864,N_18850);
and U19059 (N_19059,N_18679,N_18686);
and U19060 (N_19060,N_18767,N_18707);
or U19061 (N_19061,N_18629,N_18713);
nor U19062 (N_19062,N_18852,N_18788);
nor U19063 (N_19063,N_18797,N_18860);
nor U19064 (N_19064,N_18797,N_18829);
nand U19065 (N_19065,N_18609,N_18855);
xnor U19066 (N_19066,N_18875,N_18715);
xor U19067 (N_19067,N_18680,N_18777);
nor U19068 (N_19068,N_18888,N_18858);
and U19069 (N_19069,N_18746,N_18604);
xor U19070 (N_19070,N_18719,N_18727);
or U19071 (N_19071,N_18831,N_18830);
xor U19072 (N_19072,N_18831,N_18823);
or U19073 (N_19073,N_18693,N_18861);
or U19074 (N_19074,N_18855,N_18683);
or U19075 (N_19075,N_18774,N_18653);
or U19076 (N_19076,N_18646,N_18636);
nand U19077 (N_19077,N_18872,N_18844);
xor U19078 (N_19078,N_18700,N_18736);
xnor U19079 (N_19079,N_18821,N_18822);
and U19080 (N_19080,N_18612,N_18857);
nor U19081 (N_19081,N_18854,N_18813);
nor U19082 (N_19082,N_18757,N_18650);
nand U19083 (N_19083,N_18721,N_18653);
nor U19084 (N_19084,N_18641,N_18880);
or U19085 (N_19085,N_18830,N_18871);
nand U19086 (N_19086,N_18761,N_18631);
xor U19087 (N_19087,N_18729,N_18833);
and U19088 (N_19088,N_18810,N_18830);
or U19089 (N_19089,N_18898,N_18722);
nand U19090 (N_19090,N_18705,N_18793);
xor U19091 (N_19091,N_18761,N_18663);
xor U19092 (N_19092,N_18628,N_18747);
nand U19093 (N_19093,N_18764,N_18640);
nor U19094 (N_19094,N_18762,N_18846);
xnor U19095 (N_19095,N_18741,N_18851);
xnor U19096 (N_19096,N_18642,N_18674);
and U19097 (N_19097,N_18864,N_18645);
nor U19098 (N_19098,N_18704,N_18848);
and U19099 (N_19099,N_18887,N_18831);
and U19100 (N_19100,N_18717,N_18768);
nand U19101 (N_19101,N_18857,N_18627);
nor U19102 (N_19102,N_18633,N_18868);
and U19103 (N_19103,N_18870,N_18777);
xnor U19104 (N_19104,N_18614,N_18867);
or U19105 (N_19105,N_18641,N_18865);
or U19106 (N_19106,N_18678,N_18646);
or U19107 (N_19107,N_18855,N_18835);
and U19108 (N_19108,N_18857,N_18607);
xor U19109 (N_19109,N_18612,N_18604);
and U19110 (N_19110,N_18794,N_18689);
nor U19111 (N_19111,N_18622,N_18795);
nand U19112 (N_19112,N_18613,N_18746);
or U19113 (N_19113,N_18655,N_18663);
nand U19114 (N_19114,N_18729,N_18872);
and U19115 (N_19115,N_18798,N_18617);
nor U19116 (N_19116,N_18644,N_18685);
or U19117 (N_19117,N_18754,N_18735);
xor U19118 (N_19118,N_18844,N_18897);
nor U19119 (N_19119,N_18820,N_18769);
nand U19120 (N_19120,N_18672,N_18629);
nor U19121 (N_19121,N_18888,N_18876);
xnor U19122 (N_19122,N_18629,N_18732);
nand U19123 (N_19123,N_18604,N_18608);
and U19124 (N_19124,N_18880,N_18836);
xor U19125 (N_19125,N_18705,N_18874);
and U19126 (N_19126,N_18753,N_18743);
or U19127 (N_19127,N_18630,N_18754);
and U19128 (N_19128,N_18799,N_18885);
and U19129 (N_19129,N_18802,N_18746);
and U19130 (N_19130,N_18876,N_18808);
xnor U19131 (N_19131,N_18649,N_18615);
and U19132 (N_19132,N_18889,N_18684);
or U19133 (N_19133,N_18833,N_18612);
nand U19134 (N_19134,N_18714,N_18841);
xnor U19135 (N_19135,N_18877,N_18619);
xnor U19136 (N_19136,N_18602,N_18625);
and U19137 (N_19137,N_18864,N_18720);
nor U19138 (N_19138,N_18647,N_18619);
or U19139 (N_19139,N_18611,N_18651);
nand U19140 (N_19140,N_18849,N_18658);
nand U19141 (N_19141,N_18603,N_18880);
and U19142 (N_19142,N_18686,N_18786);
or U19143 (N_19143,N_18808,N_18870);
and U19144 (N_19144,N_18790,N_18719);
xor U19145 (N_19145,N_18826,N_18778);
and U19146 (N_19146,N_18794,N_18710);
and U19147 (N_19147,N_18806,N_18838);
or U19148 (N_19148,N_18766,N_18793);
xnor U19149 (N_19149,N_18827,N_18793);
and U19150 (N_19150,N_18732,N_18821);
xnor U19151 (N_19151,N_18752,N_18826);
or U19152 (N_19152,N_18659,N_18683);
xnor U19153 (N_19153,N_18602,N_18885);
xor U19154 (N_19154,N_18622,N_18687);
and U19155 (N_19155,N_18787,N_18805);
xor U19156 (N_19156,N_18748,N_18795);
and U19157 (N_19157,N_18658,N_18683);
nand U19158 (N_19158,N_18804,N_18698);
nor U19159 (N_19159,N_18848,N_18822);
nand U19160 (N_19160,N_18772,N_18661);
or U19161 (N_19161,N_18701,N_18704);
nand U19162 (N_19162,N_18637,N_18664);
nor U19163 (N_19163,N_18622,N_18866);
and U19164 (N_19164,N_18652,N_18744);
xnor U19165 (N_19165,N_18784,N_18703);
xnor U19166 (N_19166,N_18846,N_18674);
xnor U19167 (N_19167,N_18671,N_18867);
nor U19168 (N_19168,N_18696,N_18610);
xnor U19169 (N_19169,N_18831,N_18622);
and U19170 (N_19170,N_18679,N_18761);
nor U19171 (N_19171,N_18742,N_18876);
and U19172 (N_19172,N_18796,N_18679);
nor U19173 (N_19173,N_18826,N_18812);
nand U19174 (N_19174,N_18876,N_18616);
and U19175 (N_19175,N_18756,N_18636);
nor U19176 (N_19176,N_18639,N_18719);
nor U19177 (N_19177,N_18858,N_18864);
xnor U19178 (N_19178,N_18647,N_18760);
xor U19179 (N_19179,N_18610,N_18808);
xnor U19180 (N_19180,N_18637,N_18654);
nor U19181 (N_19181,N_18757,N_18769);
nand U19182 (N_19182,N_18834,N_18712);
or U19183 (N_19183,N_18607,N_18696);
or U19184 (N_19184,N_18605,N_18730);
xor U19185 (N_19185,N_18664,N_18793);
nand U19186 (N_19186,N_18747,N_18746);
and U19187 (N_19187,N_18714,N_18744);
nor U19188 (N_19188,N_18739,N_18808);
nor U19189 (N_19189,N_18712,N_18782);
nand U19190 (N_19190,N_18876,N_18730);
or U19191 (N_19191,N_18707,N_18661);
xor U19192 (N_19192,N_18790,N_18621);
and U19193 (N_19193,N_18897,N_18804);
nand U19194 (N_19194,N_18776,N_18804);
or U19195 (N_19195,N_18658,N_18639);
and U19196 (N_19196,N_18604,N_18709);
or U19197 (N_19197,N_18764,N_18890);
nand U19198 (N_19198,N_18675,N_18727);
nand U19199 (N_19199,N_18698,N_18829);
nor U19200 (N_19200,N_18991,N_18952);
nor U19201 (N_19201,N_19032,N_18922);
and U19202 (N_19202,N_19087,N_19033);
and U19203 (N_19203,N_19026,N_18974);
and U19204 (N_19204,N_19127,N_19159);
nor U19205 (N_19205,N_19175,N_18975);
nor U19206 (N_19206,N_18933,N_19054);
nor U19207 (N_19207,N_18988,N_18941);
nor U19208 (N_19208,N_18967,N_18971);
or U19209 (N_19209,N_19156,N_19160);
xor U19210 (N_19210,N_19099,N_18924);
and U19211 (N_19211,N_19186,N_19094);
nand U19212 (N_19212,N_19072,N_18927);
or U19213 (N_19213,N_18955,N_18990);
xor U19214 (N_19214,N_19077,N_19133);
nor U19215 (N_19215,N_18936,N_19092);
or U19216 (N_19216,N_19070,N_19171);
or U19217 (N_19217,N_19045,N_19042);
and U19218 (N_19218,N_18931,N_19086);
nand U19219 (N_19219,N_19095,N_18934);
or U19220 (N_19220,N_19153,N_18997);
nor U19221 (N_19221,N_19108,N_19091);
nand U19222 (N_19222,N_18946,N_18930);
or U19223 (N_19223,N_18949,N_19164);
nor U19224 (N_19224,N_19125,N_19036);
xnor U19225 (N_19225,N_19196,N_19059);
or U19226 (N_19226,N_18903,N_19063);
nor U19227 (N_19227,N_18956,N_19199);
nor U19228 (N_19228,N_19101,N_19115);
nor U19229 (N_19229,N_19193,N_19058);
nand U19230 (N_19230,N_19148,N_18948);
or U19231 (N_19231,N_19006,N_19128);
and U19232 (N_19232,N_19126,N_19073);
and U19233 (N_19233,N_19177,N_18994);
and U19234 (N_19234,N_18915,N_19060);
nor U19235 (N_19235,N_19085,N_19136);
xor U19236 (N_19236,N_19104,N_19080);
nand U19237 (N_19237,N_18964,N_19114);
or U19238 (N_19238,N_19027,N_19075);
and U19239 (N_19239,N_19144,N_19025);
nor U19240 (N_19240,N_18937,N_18984);
nand U19241 (N_19241,N_18917,N_18965);
and U19242 (N_19242,N_19123,N_18995);
or U19243 (N_19243,N_18978,N_19020);
and U19244 (N_19244,N_19028,N_19037);
and U19245 (N_19245,N_18943,N_19141);
or U19246 (N_19246,N_19157,N_19056);
and U19247 (N_19247,N_19180,N_19001);
xor U19248 (N_19248,N_19170,N_18951);
nand U19249 (N_19249,N_19078,N_19000);
or U19250 (N_19250,N_19137,N_19035);
nor U19251 (N_19251,N_18916,N_19188);
or U19252 (N_19252,N_19038,N_19190);
xnor U19253 (N_19253,N_19161,N_18976);
nor U19254 (N_19254,N_18999,N_19043);
or U19255 (N_19255,N_19181,N_18985);
nand U19256 (N_19256,N_19079,N_19197);
nand U19257 (N_19257,N_19183,N_19098);
nand U19258 (N_19258,N_19097,N_19174);
or U19259 (N_19259,N_19018,N_19015);
and U19260 (N_19260,N_19021,N_19184);
nand U19261 (N_19261,N_19010,N_18972);
or U19262 (N_19262,N_19017,N_18908);
nor U19263 (N_19263,N_19191,N_19076);
and U19264 (N_19264,N_19048,N_19185);
nand U19265 (N_19265,N_19150,N_19074);
or U19266 (N_19266,N_18947,N_19049);
nand U19267 (N_19267,N_18981,N_19081);
and U19268 (N_19268,N_19132,N_19145);
and U19269 (N_19269,N_19192,N_19154);
and U19270 (N_19270,N_18977,N_19083);
xor U19271 (N_19271,N_18923,N_18904);
nor U19272 (N_19272,N_18954,N_18932);
and U19273 (N_19273,N_18959,N_19012);
or U19274 (N_19274,N_18986,N_18963);
nand U19275 (N_19275,N_18935,N_19142);
or U19276 (N_19276,N_19167,N_19189);
nor U19277 (N_19277,N_18913,N_19195);
and U19278 (N_19278,N_19050,N_18905);
nor U19279 (N_19279,N_19121,N_19014);
nand U19280 (N_19280,N_19030,N_18960);
or U19281 (N_19281,N_19082,N_19112);
and U19282 (N_19282,N_18912,N_19068);
and U19283 (N_19283,N_19007,N_19002);
xnor U19284 (N_19284,N_18966,N_19147);
nand U19285 (N_19285,N_18911,N_19120);
or U19286 (N_19286,N_19069,N_18907);
nand U19287 (N_19287,N_19071,N_19039);
nor U19288 (N_19288,N_18979,N_18902);
or U19289 (N_19289,N_19096,N_18944);
xnor U19290 (N_19290,N_19084,N_18939);
nor U19291 (N_19291,N_19117,N_19003);
and U19292 (N_19292,N_18970,N_18901);
and U19293 (N_19293,N_18914,N_19089);
xnor U19294 (N_19294,N_18980,N_18938);
or U19295 (N_19295,N_19198,N_18969);
and U19296 (N_19296,N_19152,N_19111);
nor U19297 (N_19297,N_19122,N_19165);
xor U19298 (N_19298,N_19105,N_18983);
or U19299 (N_19299,N_19149,N_19146);
or U19300 (N_19300,N_19051,N_19040);
nor U19301 (N_19301,N_19100,N_18968);
or U19302 (N_19302,N_19135,N_18998);
or U19303 (N_19303,N_19119,N_18945);
nand U19304 (N_19304,N_19151,N_19009);
nor U19305 (N_19305,N_19065,N_19046);
nor U19306 (N_19306,N_19052,N_19162);
nand U19307 (N_19307,N_19047,N_19102);
and U19308 (N_19308,N_19139,N_18961);
and U19309 (N_19309,N_19062,N_18900);
nor U19310 (N_19310,N_18919,N_18953);
nand U19311 (N_19311,N_19041,N_18958);
or U19312 (N_19312,N_19155,N_19031);
xnor U19313 (N_19313,N_18957,N_19194);
or U19314 (N_19314,N_19024,N_19163);
xnor U19315 (N_19315,N_19124,N_19113);
and U19316 (N_19316,N_19057,N_18918);
and U19317 (N_19317,N_18926,N_18996);
or U19318 (N_19318,N_19011,N_19131);
nor U19319 (N_19319,N_18910,N_19103);
nand U19320 (N_19320,N_19179,N_19143);
and U19321 (N_19321,N_19029,N_19053);
or U19322 (N_19322,N_19172,N_19173);
or U19323 (N_19323,N_19022,N_19187);
nand U19324 (N_19324,N_18921,N_19138);
nor U19325 (N_19325,N_18940,N_19019);
or U19326 (N_19326,N_18929,N_19129);
or U19327 (N_19327,N_18987,N_19178);
nand U19328 (N_19328,N_19166,N_18993);
and U19329 (N_19329,N_19064,N_19134);
nor U19330 (N_19330,N_19008,N_18906);
xnor U19331 (N_19331,N_19169,N_19116);
and U19332 (N_19332,N_19118,N_19023);
xnor U19333 (N_19333,N_18942,N_18925);
and U19334 (N_19334,N_19168,N_19093);
nand U19335 (N_19335,N_19140,N_18992);
nor U19336 (N_19336,N_19130,N_18989);
or U19337 (N_19337,N_19088,N_19016);
nand U19338 (N_19338,N_19176,N_19066);
or U19339 (N_19339,N_18962,N_19004);
or U19340 (N_19340,N_19110,N_19090);
nand U19341 (N_19341,N_19034,N_19044);
xor U19342 (N_19342,N_19109,N_18928);
nor U19343 (N_19343,N_19107,N_19061);
nand U19344 (N_19344,N_18973,N_19106);
nor U19345 (N_19345,N_19158,N_19055);
nand U19346 (N_19346,N_19067,N_18920);
nor U19347 (N_19347,N_19005,N_19013);
xnor U19348 (N_19348,N_18909,N_19182);
or U19349 (N_19349,N_18982,N_18950);
nand U19350 (N_19350,N_19023,N_19065);
and U19351 (N_19351,N_19076,N_19199);
nor U19352 (N_19352,N_19161,N_19035);
nand U19353 (N_19353,N_19021,N_19024);
nor U19354 (N_19354,N_19135,N_19026);
nor U19355 (N_19355,N_19052,N_19104);
and U19356 (N_19356,N_19022,N_19017);
nand U19357 (N_19357,N_18979,N_19051);
nor U19358 (N_19358,N_19163,N_19107);
nand U19359 (N_19359,N_19112,N_19063);
and U19360 (N_19360,N_19049,N_18953);
nand U19361 (N_19361,N_19054,N_18953);
and U19362 (N_19362,N_18994,N_19067);
xor U19363 (N_19363,N_18961,N_18977);
nand U19364 (N_19364,N_19109,N_19114);
nor U19365 (N_19365,N_19035,N_18902);
xor U19366 (N_19366,N_19039,N_18988);
nor U19367 (N_19367,N_18928,N_18931);
or U19368 (N_19368,N_18922,N_19135);
nand U19369 (N_19369,N_18901,N_18993);
nor U19370 (N_19370,N_18997,N_19115);
or U19371 (N_19371,N_18946,N_19097);
xnor U19372 (N_19372,N_19011,N_19107);
nor U19373 (N_19373,N_19096,N_18974);
nor U19374 (N_19374,N_19148,N_19119);
or U19375 (N_19375,N_19162,N_19196);
and U19376 (N_19376,N_18943,N_19166);
nor U19377 (N_19377,N_19030,N_18909);
nand U19378 (N_19378,N_19034,N_18973);
and U19379 (N_19379,N_19039,N_19040);
xor U19380 (N_19380,N_19189,N_19154);
nand U19381 (N_19381,N_19026,N_18915);
xor U19382 (N_19382,N_18981,N_19040);
or U19383 (N_19383,N_18947,N_19124);
xor U19384 (N_19384,N_19024,N_19110);
and U19385 (N_19385,N_19070,N_18962);
nand U19386 (N_19386,N_19195,N_18923);
nor U19387 (N_19387,N_18923,N_19009);
xnor U19388 (N_19388,N_19171,N_19144);
xor U19389 (N_19389,N_19169,N_18990);
nor U19390 (N_19390,N_19028,N_18979);
and U19391 (N_19391,N_18976,N_18997);
or U19392 (N_19392,N_19038,N_19188);
nand U19393 (N_19393,N_18967,N_18985);
xnor U19394 (N_19394,N_19106,N_18920);
xnor U19395 (N_19395,N_19120,N_18940);
xor U19396 (N_19396,N_19168,N_19059);
xnor U19397 (N_19397,N_19146,N_19108);
and U19398 (N_19398,N_19113,N_18903);
nor U19399 (N_19399,N_18978,N_18986);
nor U19400 (N_19400,N_18986,N_19053);
nand U19401 (N_19401,N_19144,N_19053);
nor U19402 (N_19402,N_19026,N_18903);
xnor U19403 (N_19403,N_18912,N_18991);
and U19404 (N_19404,N_19188,N_19161);
or U19405 (N_19405,N_19059,N_19166);
xnor U19406 (N_19406,N_19136,N_18964);
nand U19407 (N_19407,N_19150,N_18916);
nand U19408 (N_19408,N_18929,N_18965);
xor U19409 (N_19409,N_19020,N_19055);
nand U19410 (N_19410,N_19114,N_19171);
nor U19411 (N_19411,N_18979,N_18987);
nand U19412 (N_19412,N_18997,N_18985);
nand U19413 (N_19413,N_19027,N_18938);
nor U19414 (N_19414,N_19070,N_19032);
or U19415 (N_19415,N_19084,N_19114);
nand U19416 (N_19416,N_18950,N_18929);
nand U19417 (N_19417,N_18944,N_19161);
nand U19418 (N_19418,N_19127,N_18991);
nand U19419 (N_19419,N_19077,N_19186);
or U19420 (N_19420,N_18986,N_19047);
nor U19421 (N_19421,N_18988,N_19069);
or U19422 (N_19422,N_19156,N_18907);
and U19423 (N_19423,N_19194,N_18998);
and U19424 (N_19424,N_19063,N_18938);
or U19425 (N_19425,N_19189,N_19009);
and U19426 (N_19426,N_19046,N_18966);
xor U19427 (N_19427,N_19151,N_18938);
or U19428 (N_19428,N_18953,N_18978);
and U19429 (N_19429,N_19153,N_19055);
nor U19430 (N_19430,N_18959,N_19177);
and U19431 (N_19431,N_19120,N_18961);
or U19432 (N_19432,N_18963,N_18907);
nor U19433 (N_19433,N_19143,N_19019);
xnor U19434 (N_19434,N_18903,N_18965);
or U19435 (N_19435,N_18997,N_19061);
or U19436 (N_19436,N_18936,N_19069);
or U19437 (N_19437,N_18999,N_19109);
nor U19438 (N_19438,N_19170,N_19194);
xor U19439 (N_19439,N_18908,N_19058);
or U19440 (N_19440,N_19021,N_19084);
nand U19441 (N_19441,N_19188,N_18966);
and U19442 (N_19442,N_19001,N_19022);
or U19443 (N_19443,N_19139,N_18947);
or U19444 (N_19444,N_19105,N_19169);
nand U19445 (N_19445,N_18984,N_18943);
and U19446 (N_19446,N_19074,N_18910);
or U19447 (N_19447,N_19088,N_19005);
nand U19448 (N_19448,N_19179,N_19109);
xor U19449 (N_19449,N_19055,N_19109);
nand U19450 (N_19450,N_19167,N_19079);
xor U19451 (N_19451,N_18959,N_18966);
nor U19452 (N_19452,N_19049,N_18982);
nor U19453 (N_19453,N_19031,N_18914);
nor U19454 (N_19454,N_19005,N_18982);
and U19455 (N_19455,N_19111,N_19163);
nor U19456 (N_19456,N_18975,N_19079);
nand U19457 (N_19457,N_19039,N_19144);
nor U19458 (N_19458,N_18940,N_19000);
nor U19459 (N_19459,N_19059,N_18905);
nand U19460 (N_19460,N_18999,N_18998);
nand U19461 (N_19461,N_19128,N_19044);
nand U19462 (N_19462,N_19195,N_19162);
or U19463 (N_19463,N_19007,N_18955);
xnor U19464 (N_19464,N_18904,N_18903);
nand U19465 (N_19465,N_19152,N_18908);
or U19466 (N_19466,N_18943,N_19044);
nand U19467 (N_19467,N_19153,N_19175);
and U19468 (N_19468,N_19161,N_19128);
nor U19469 (N_19469,N_19046,N_19027);
nand U19470 (N_19470,N_19142,N_18936);
nand U19471 (N_19471,N_19176,N_19003);
nor U19472 (N_19472,N_19167,N_18904);
xor U19473 (N_19473,N_18916,N_19017);
or U19474 (N_19474,N_19025,N_19044);
nor U19475 (N_19475,N_19045,N_19164);
and U19476 (N_19476,N_19193,N_18949);
and U19477 (N_19477,N_19098,N_19101);
and U19478 (N_19478,N_19054,N_19078);
xnor U19479 (N_19479,N_19198,N_19074);
and U19480 (N_19480,N_19143,N_18906);
and U19481 (N_19481,N_19103,N_18985);
nand U19482 (N_19482,N_19097,N_18912);
xor U19483 (N_19483,N_19005,N_19067);
nor U19484 (N_19484,N_18932,N_18958);
nor U19485 (N_19485,N_19038,N_19117);
xor U19486 (N_19486,N_18991,N_19115);
or U19487 (N_19487,N_19001,N_19116);
nand U19488 (N_19488,N_19119,N_19018);
nor U19489 (N_19489,N_18951,N_18991);
nand U19490 (N_19490,N_19135,N_18985);
or U19491 (N_19491,N_18913,N_18927);
or U19492 (N_19492,N_19068,N_18922);
nand U19493 (N_19493,N_18928,N_19052);
or U19494 (N_19494,N_18930,N_19158);
nand U19495 (N_19495,N_19047,N_19142);
and U19496 (N_19496,N_19015,N_18927);
or U19497 (N_19497,N_19137,N_18926);
nand U19498 (N_19498,N_18952,N_18981);
nor U19499 (N_19499,N_19111,N_19054);
xor U19500 (N_19500,N_19318,N_19450);
nor U19501 (N_19501,N_19307,N_19471);
or U19502 (N_19502,N_19235,N_19456);
nand U19503 (N_19503,N_19209,N_19332);
xnor U19504 (N_19504,N_19345,N_19322);
and U19505 (N_19505,N_19395,N_19316);
or U19506 (N_19506,N_19373,N_19296);
and U19507 (N_19507,N_19300,N_19449);
nand U19508 (N_19508,N_19444,N_19493);
nand U19509 (N_19509,N_19398,N_19394);
nand U19510 (N_19510,N_19371,N_19416);
nor U19511 (N_19511,N_19245,N_19366);
or U19512 (N_19512,N_19341,N_19432);
nand U19513 (N_19513,N_19491,N_19213);
or U19514 (N_19514,N_19429,N_19272);
or U19515 (N_19515,N_19314,N_19287);
nand U19516 (N_19516,N_19333,N_19409);
xor U19517 (N_19517,N_19443,N_19362);
or U19518 (N_19518,N_19397,N_19410);
or U19519 (N_19519,N_19315,N_19472);
nand U19520 (N_19520,N_19492,N_19223);
nor U19521 (N_19521,N_19216,N_19446);
and U19522 (N_19522,N_19305,N_19474);
or U19523 (N_19523,N_19434,N_19384);
or U19524 (N_19524,N_19447,N_19352);
nor U19525 (N_19525,N_19377,N_19445);
and U19526 (N_19526,N_19228,N_19336);
nand U19527 (N_19527,N_19415,N_19263);
or U19528 (N_19528,N_19337,N_19277);
or U19529 (N_19529,N_19481,N_19278);
and U19530 (N_19530,N_19258,N_19479);
or U19531 (N_19531,N_19282,N_19460);
nand U19532 (N_19532,N_19291,N_19424);
and U19533 (N_19533,N_19349,N_19358);
nand U19534 (N_19534,N_19407,N_19422);
or U19535 (N_19535,N_19306,N_19311);
nor U19536 (N_19536,N_19390,N_19323);
xor U19537 (N_19537,N_19490,N_19431);
nand U19538 (N_19538,N_19230,N_19378);
or U19539 (N_19539,N_19265,N_19370);
and U19540 (N_19540,N_19383,N_19468);
nor U19541 (N_19541,N_19310,N_19374);
or U19542 (N_19542,N_19303,N_19484);
nand U19543 (N_19543,N_19357,N_19262);
nor U19544 (N_19544,N_19299,N_19498);
xnor U19545 (N_19545,N_19252,N_19388);
xor U19546 (N_19546,N_19288,N_19203);
xor U19547 (N_19547,N_19313,N_19381);
nand U19548 (N_19548,N_19419,N_19331);
nand U19549 (N_19549,N_19246,N_19380);
or U19550 (N_19550,N_19253,N_19321);
nor U19551 (N_19551,N_19236,N_19408);
nor U19552 (N_19552,N_19206,N_19465);
and U19553 (N_19553,N_19375,N_19273);
nor U19554 (N_19554,N_19309,N_19355);
and U19555 (N_19555,N_19241,N_19454);
nand U19556 (N_19556,N_19297,N_19229);
nand U19557 (N_19557,N_19205,N_19420);
xnor U19558 (N_19558,N_19342,N_19351);
or U19559 (N_19559,N_19275,N_19488);
and U19560 (N_19560,N_19254,N_19217);
xor U19561 (N_19561,N_19266,N_19347);
and U19562 (N_19562,N_19452,N_19391);
nand U19563 (N_19563,N_19251,N_19400);
nand U19564 (N_19564,N_19364,N_19274);
nor U19565 (N_19565,N_19289,N_19376);
nor U19566 (N_19566,N_19497,N_19346);
nor U19567 (N_19567,N_19379,N_19448);
and U19568 (N_19568,N_19312,N_19354);
nand U19569 (N_19569,N_19330,N_19234);
and U19570 (N_19570,N_19267,N_19319);
and U19571 (N_19571,N_19259,N_19283);
or U19572 (N_19572,N_19451,N_19269);
nor U19573 (N_19573,N_19353,N_19215);
xor U19574 (N_19574,N_19204,N_19393);
nand U19575 (N_19575,N_19281,N_19435);
or U19576 (N_19576,N_19290,N_19255);
xnor U19577 (N_19577,N_19276,N_19338);
nand U19578 (N_19578,N_19369,N_19461);
or U19579 (N_19579,N_19404,N_19495);
xor U19580 (N_19580,N_19427,N_19417);
and U19581 (N_19581,N_19208,N_19477);
xor U19582 (N_19582,N_19367,N_19414);
or U19583 (N_19583,N_19402,N_19486);
nor U19584 (N_19584,N_19457,N_19339);
or U19585 (N_19585,N_19441,N_19286);
or U19586 (N_19586,N_19250,N_19348);
or U19587 (N_19587,N_19294,N_19436);
or U19588 (N_19588,N_19324,N_19334);
or U19589 (N_19589,N_19210,N_19499);
and U19590 (N_19590,N_19264,N_19361);
nand U19591 (N_19591,N_19405,N_19249);
or U19592 (N_19592,N_19438,N_19200);
nor U19593 (N_19593,N_19487,N_19219);
xnor U19594 (N_19594,N_19257,N_19317);
or U19595 (N_19595,N_19463,N_19421);
or U19596 (N_19596,N_19406,N_19244);
xnor U19597 (N_19597,N_19225,N_19350);
nor U19598 (N_19598,N_19399,N_19295);
and U19599 (N_19599,N_19478,N_19320);
or U19600 (N_19600,N_19280,N_19248);
xor U19601 (N_19601,N_19308,N_19428);
or U19602 (N_19602,N_19467,N_19413);
or U19603 (N_19603,N_19401,N_19425);
or U19604 (N_19604,N_19279,N_19476);
nand U19605 (N_19605,N_19494,N_19458);
nor U19606 (N_19606,N_19207,N_19260);
nor U19607 (N_19607,N_19335,N_19242);
and U19608 (N_19608,N_19455,N_19247);
nand U19609 (N_19609,N_19464,N_19327);
and U19610 (N_19610,N_19466,N_19271);
and U19611 (N_19611,N_19411,N_19224);
nand U19612 (N_19612,N_19453,N_19270);
and U19613 (N_19613,N_19256,N_19233);
xor U19614 (N_19614,N_19365,N_19359);
and U19615 (N_19615,N_19485,N_19221);
or U19616 (N_19616,N_19469,N_19372);
xor U19617 (N_19617,N_19363,N_19238);
and U19618 (N_19618,N_19344,N_19268);
nor U19619 (N_19619,N_19387,N_19218);
or U19620 (N_19620,N_19433,N_19475);
or U19621 (N_19621,N_19462,N_19304);
nor U19622 (N_19622,N_19480,N_19392);
and U19623 (N_19623,N_19222,N_19227);
nor U19624 (N_19624,N_19423,N_19340);
xnor U19625 (N_19625,N_19496,N_19360);
xor U19626 (N_19626,N_19439,N_19326);
xor U19627 (N_19627,N_19261,N_19403);
nor U19628 (N_19628,N_19356,N_19489);
nand U19629 (N_19629,N_19243,N_19442);
nand U19630 (N_19630,N_19239,N_19343);
xnor U19631 (N_19631,N_19459,N_19293);
or U19632 (N_19632,N_19382,N_19214);
or U19633 (N_19633,N_19240,N_19418);
and U19634 (N_19634,N_19211,N_19220);
or U19635 (N_19635,N_19440,N_19482);
xnor U19636 (N_19636,N_19396,N_19301);
xor U19637 (N_19637,N_19385,N_19328);
and U19638 (N_19638,N_19226,N_19302);
xor U19639 (N_19639,N_19298,N_19412);
and U19640 (N_19640,N_19386,N_19325);
nor U19641 (N_19641,N_19237,N_19483);
and U19642 (N_19642,N_19231,N_19426);
nor U19643 (N_19643,N_19437,N_19284);
or U19644 (N_19644,N_19212,N_19430);
nor U19645 (N_19645,N_19473,N_19201);
nor U19646 (N_19646,N_19389,N_19368);
and U19647 (N_19647,N_19470,N_19232);
or U19648 (N_19648,N_19285,N_19292);
and U19649 (N_19649,N_19202,N_19329);
nor U19650 (N_19650,N_19452,N_19395);
or U19651 (N_19651,N_19321,N_19496);
and U19652 (N_19652,N_19371,N_19232);
nor U19653 (N_19653,N_19480,N_19289);
or U19654 (N_19654,N_19287,N_19438);
xor U19655 (N_19655,N_19290,N_19436);
xnor U19656 (N_19656,N_19468,N_19219);
or U19657 (N_19657,N_19317,N_19460);
nor U19658 (N_19658,N_19235,N_19299);
or U19659 (N_19659,N_19234,N_19305);
nand U19660 (N_19660,N_19275,N_19377);
or U19661 (N_19661,N_19443,N_19453);
and U19662 (N_19662,N_19445,N_19287);
and U19663 (N_19663,N_19483,N_19352);
nor U19664 (N_19664,N_19212,N_19215);
nor U19665 (N_19665,N_19414,N_19274);
nor U19666 (N_19666,N_19378,N_19228);
xor U19667 (N_19667,N_19492,N_19317);
nor U19668 (N_19668,N_19384,N_19228);
nor U19669 (N_19669,N_19276,N_19340);
or U19670 (N_19670,N_19369,N_19344);
and U19671 (N_19671,N_19332,N_19258);
and U19672 (N_19672,N_19354,N_19311);
nor U19673 (N_19673,N_19330,N_19443);
nand U19674 (N_19674,N_19262,N_19481);
or U19675 (N_19675,N_19217,N_19339);
xor U19676 (N_19676,N_19476,N_19328);
or U19677 (N_19677,N_19233,N_19413);
nand U19678 (N_19678,N_19329,N_19395);
and U19679 (N_19679,N_19247,N_19407);
nand U19680 (N_19680,N_19360,N_19275);
xor U19681 (N_19681,N_19331,N_19346);
or U19682 (N_19682,N_19300,N_19442);
and U19683 (N_19683,N_19222,N_19489);
and U19684 (N_19684,N_19356,N_19387);
nand U19685 (N_19685,N_19322,N_19326);
xnor U19686 (N_19686,N_19216,N_19301);
nand U19687 (N_19687,N_19260,N_19277);
xnor U19688 (N_19688,N_19243,N_19467);
nor U19689 (N_19689,N_19346,N_19244);
or U19690 (N_19690,N_19237,N_19318);
nor U19691 (N_19691,N_19403,N_19288);
and U19692 (N_19692,N_19250,N_19311);
xnor U19693 (N_19693,N_19306,N_19287);
or U19694 (N_19694,N_19443,N_19294);
nor U19695 (N_19695,N_19341,N_19329);
nor U19696 (N_19696,N_19219,N_19218);
xor U19697 (N_19697,N_19202,N_19413);
xnor U19698 (N_19698,N_19244,N_19338);
or U19699 (N_19699,N_19483,N_19489);
xnor U19700 (N_19700,N_19292,N_19342);
and U19701 (N_19701,N_19297,N_19438);
nor U19702 (N_19702,N_19273,N_19252);
nor U19703 (N_19703,N_19246,N_19465);
and U19704 (N_19704,N_19492,N_19318);
nand U19705 (N_19705,N_19467,N_19479);
nor U19706 (N_19706,N_19313,N_19387);
nor U19707 (N_19707,N_19496,N_19422);
xor U19708 (N_19708,N_19249,N_19473);
nor U19709 (N_19709,N_19365,N_19244);
and U19710 (N_19710,N_19482,N_19369);
xor U19711 (N_19711,N_19447,N_19353);
or U19712 (N_19712,N_19472,N_19474);
or U19713 (N_19713,N_19406,N_19227);
xnor U19714 (N_19714,N_19219,N_19245);
and U19715 (N_19715,N_19379,N_19466);
nand U19716 (N_19716,N_19304,N_19301);
and U19717 (N_19717,N_19336,N_19409);
nand U19718 (N_19718,N_19231,N_19332);
or U19719 (N_19719,N_19271,N_19279);
nor U19720 (N_19720,N_19426,N_19247);
or U19721 (N_19721,N_19221,N_19455);
nor U19722 (N_19722,N_19252,N_19357);
and U19723 (N_19723,N_19396,N_19308);
xor U19724 (N_19724,N_19424,N_19399);
or U19725 (N_19725,N_19450,N_19238);
and U19726 (N_19726,N_19441,N_19410);
xnor U19727 (N_19727,N_19239,N_19451);
nor U19728 (N_19728,N_19317,N_19203);
nand U19729 (N_19729,N_19226,N_19362);
nor U19730 (N_19730,N_19487,N_19393);
or U19731 (N_19731,N_19232,N_19499);
nor U19732 (N_19732,N_19391,N_19212);
xnor U19733 (N_19733,N_19276,N_19274);
nor U19734 (N_19734,N_19220,N_19345);
and U19735 (N_19735,N_19280,N_19218);
nor U19736 (N_19736,N_19381,N_19213);
nand U19737 (N_19737,N_19251,N_19478);
nand U19738 (N_19738,N_19202,N_19214);
xnor U19739 (N_19739,N_19411,N_19473);
and U19740 (N_19740,N_19355,N_19271);
and U19741 (N_19741,N_19362,N_19378);
and U19742 (N_19742,N_19496,N_19340);
xnor U19743 (N_19743,N_19433,N_19435);
and U19744 (N_19744,N_19287,N_19299);
nand U19745 (N_19745,N_19219,N_19485);
or U19746 (N_19746,N_19253,N_19254);
xnor U19747 (N_19747,N_19337,N_19253);
nand U19748 (N_19748,N_19444,N_19246);
xor U19749 (N_19749,N_19220,N_19245);
or U19750 (N_19750,N_19424,N_19347);
nand U19751 (N_19751,N_19227,N_19211);
nand U19752 (N_19752,N_19420,N_19294);
nand U19753 (N_19753,N_19259,N_19408);
and U19754 (N_19754,N_19219,N_19470);
nor U19755 (N_19755,N_19297,N_19264);
nor U19756 (N_19756,N_19395,N_19244);
and U19757 (N_19757,N_19443,N_19376);
nand U19758 (N_19758,N_19290,N_19499);
and U19759 (N_19759,N_19267,N_19459);
or U19760 (N_19760,N_19491,N_19350);
nor U19761 (N_19761,N_19456,N_19372);
nor U19762 (N_19762,N_19221,N_19384);
nand U19763 (N_19763,N_19417,N_19480);
or U19764 (N_19764,N_19213,N_19303);
nand U19765 (N_19765,N_19334,N_19476);
or U19766 (N_19766,N_19382,N_19462);
nor U19767 (N_19767,N_19413,N_19248);
and U19768 (N_19768,N_19209,N_19291);
nor U19769 (N_19769,N_19279,N_19322);
xor U19770 (N_19770,N_19355,N_19320);
nor U19771 (N_19771,N_19406,N_19417);
nand U19772 (N_19772,N_19410,N_19273);
and U19773 (N_19773,N_19262,N_19356);
xor U19774 (N_19774,N_19262,N_19382);
and U19775 (N_19775,N_19273,N_19285);
and U19776 (N_19776,N_19461,N_19301);
and U19777 (N_19777,N_19300,N_19343);
xnor U19778 (N_19778,N_19378,N_19335);
nand U19779 (N_19779,N_19262,N_19411);
and U19780 (N_19780,N_19280,N_19234);
xor U19781 (N_19781,N_19314,N_19368);
and U19782 (N_19782,N_19280,N_19315);
and U19783 (N_19783,N_19227,N_19487);
xor U19784 (N_19784,N_19401,N_19343);
nor U19785 (N_19785,N_19281,N_19254);
nand U19786 (N_19786,N_19430,N_19481);
xnor U19787 (N_19787,N_19263,N_19324);
or U19788 (N_19788,N_19477,N_19270);
or U19789 (N_19789,N_19219,N_19339);
nand U19790 (N_19790,N_19427,N_19389);
or U19791 (N_19791,N_19211,N_19304);
nor U19792 (N_19792,N_19496,N_19395);
or U19793 (N_19793,N_19308,N_19345);
or U19794 (N_19794,N_19400,N_19316);
nor U19795 (N_19795,N_19310,N_19262);
or U19796 (N_19796,N_19222,N_19387);
xnor U19797 (N_19797,N_19229,N_19261);
and U19798 (N_19798,N_19484,N_19394);
nor U19799 (N_19799,N_19332,N_19423);
nor U19800 (N_19800,N_19528,N_19512);
or U19801 (N_19801,N_19725,N_19754);
xor U19802 (N_19802,N_19755,N_19589);
and U19803 (N_19803,N_19652,N_19794);
xor U19804 (N_19804,N_19592,N_19553);
nor U19805 (N_19805,N_19764,N_19714);
nand U19806 (N_19806,N_19762,N_19639);
nor U19807 (N_19807,N_19751,N_19686);
xor U19808 (N_19808,N_19554,N_19692);
or U19809 (N_19809,N_19786,N_19783);
xor U19810 (N_19810,N_19775,N_19596);
xor U19811 (N_19811,N_19769,N_19524);
or U19812 (N_19812,N_19698,N_19758);
nand U19813 (N_19813,N_19649,N_19727);
xnor U19814 (N_19814,N_19689,N_19590);
nor U19815 (N_19815,N_19556,N_19543);
xnor U19816 (N_19816,N_19676,N_19618);
nor U19817 (N_19817,N_19566,N_19761);
or U19818 (N_19818,N_19748,N_19609);
nand U19819 (N_19819,N_19646,N_19627);
and U19820 (N_19820,N_19675,N_19508);
xnor U19821 (N_19821,N_19561,N_19572);
nor U19822 (N_19822,N_19626,N_19506);
nand U19823 (N_19823,N_19551,N_19549);
or U19824 (N_19824,N_19778,N_19700);
nor U19825 (N_19825,N_19611,N_19647);
and U19826 (N_19826,N_19516,N_19637);
or U19827 (N_19827,N_19580,N_19658);
nand U19828 (N_19828,N_19741,N_19671);
and U19829 (N_19829,N_19745,N_19530);
nor U19830 (N_19830,N_19797,N_19788);
nor U19831 (N_19831,N_19653,N_19708);
and U19832 (N_19832,N_19687,N_19739);
and U19833 (N_19833,N_19537,N_19756);
xnor U19834 (N_19834,N_19621,N_19677);
xor U19835 (N_19835,N_19520,N_19777);
and U19836 (N_19836,N_19555,N_19563);
nor U19837 (N_19837,N_19505,N_19548);
and U19838 (N_19838,N_19565,N_19685);
nand U19839 (N_19839,N_19582,N_19503);
or U19840 (N_19840,N_19730,N_19773);
xor U19841 (N_19841,N_19644,N_19594);
nor U19842 (N_19842,N_19791,N_19767);
nand U19843 (N_19843,N_19583,N_19624);
xor U19844 (N_19844,N_19720,N_19546);
and U19845 (N_19845,N_19779,N_19722);
and U19846 (N_19846,N_19604,N_19735);
and U19847 (N_19847,N_19796,N_19531);
or U19848 (N_19848,N_19705,N_19681);
xor U19849 (N_19849,N_19747,N_19519);
or U19850 (N_19850,N_19606,N_19614);
nand U19851 (N_19851,N_19655,N_19753);
and U19852 (N_19852,N_19544,N_19682);
or U19853 (N_19853,N_19518,N_19608);
xnor U19854 (N_19854,N_19522,N_19579);
xor U19855 (N_19855,N_19736,N_19645);
and U19856 (N_19856,N_19684,N_19776);
xor U19857 (N_19857,N_19673,N_19709);
nand U19858 (N_19858,N_19679,N_19691);
nand U19859 (N_19859,N_19651,N_19662);
nand U19860 (N_19860,N_19672,N_19517);
or U19861 (N_19861,N_19694,N_19663);
or U19862 (N_19862,N_19781,N_19703);
nand U19863 (N_19863,N_19719,N_19780);
xor U19864 (N_19864,N_19670,N_19630);
nand U19865 (N_19865,N_19772,N_19619);
or U19866 (N_19866,N_19558,N_19539);
nand U19867 (N_19867,N_19620,N_19667);
nand U19868 (N_19868,N_19657,N_19710);
and U19869 (N_19869,N_19527,N_19634);
nor U19870 (N_19870,N_19640,N_19521);
nor U19871 (N_19871,N_19731,N_19654);
nand U19872 (N_19872,N_19602,N_19633);
or U19873 (N_19873,N_19510,N_19711);
xnor U19874 (N_19874,N_19744,N_19540);
and U19875 (N_19875,N_19605,N_19501);
xor U19876 (N_19876,N_19683,N_19661);
nand U19877 (N_19877,N_19784,N_19623);
xnor U19878 (N_19878,N_19766,N_19538);
or U19879 (N_19879,N_19598,N_19502);
and U19880 (N_19880,N_19575,N_19523);
xnor U19881 (N_19881,N_19536,N_19511);
and U19882 (N_19882,N_19638,N_19770);
nand U19883 (N_19883,N_19718,N_19729);
or U19884 (N_19884,N_19631,N_19595);
nand U19885 (N_19885,N_19706,N_19799);
nand U19886 (N_19886,N_19678,N_19574);
nand U19887 (N_19887,N_19693,N_19577);
nor U19888 (N_19888,N_19534,N_19768);
and U19889 (N_19889,N_19750,N_19541);
or U19890 (N_19890,N_19588,N_19790);
and U19891 (N_19891,N_19732,N_19584);
xnor U19892 (N_19892,N_19532,N_19547);
nand U19893 (N_19893,N_19734,N_19571);
xor U19894 (N_19894,N_19615,N_19746);
nand U19895 (N_19895,N_19696,N_19629);
nand U19896 (N_19896,N_19642,N_19564);
nor U19897 (N_19897,N_19712,N_19789);
and U19898 (N_19898,N_19716,N_19576);
and U19899 (N_19899,N_19733,N_19636);
xor U19900 (N_19900,N_19635,N_19593);
nor U19901 (N_19901,N_19798,N_19728);
xnor U19902 (N_19902,N_19607,N_19585);
and U19903 (N_19903,N_19591,N_19717);
nand U19904 (N_19904,N_19697,N_19795);
and U19905 (N_19905,N_19507,N_19599);
nand U19906 (N_19906,N_19601,N_19567);
nor U19907 (N_19907,N_19550,N_19569);
nand U19908 (N_19908,N_19763,N_19526);
xnor U19909 (N_19909,N_19559,N_19665);
nor U19910 (N_19910,N_19664,N_19765);
and U19911 (N_19911,N_19740,N_19578);
or U19912 (N_19912,N_19560,N_19704);
nand U19913 (N_19913,N_19743,N_19656);
xnor U19914 (N_19914,N_19688,N_19785);
and U19915 (N_19915,N_19641,N_19724);
nor U19916 (N_19916,N_19525,N_19695);
xor U19917 (N_19917,N_19632,N_19668);
or U19918 (N_19918,N_19513,N_19557);
nand U19919 (N_19919,N_19699,N_19573);
nor U19920 (N_19920,N_19628,N_19622);
and U19921 (N_19921,N_19600,N_19792);
nand U19922 (N_19922,N_19648,N_19603);
nand U19923 (N_19923,N_19562,N_19509);
nor U19924 (N_19924,N_19535,N_19721);
xnor U19925 (N_19925,N_19581,N_19737);
or U19926 (N_19926,N_19597,N_19533);
and U19927 (N_19927,N_19723,N_19666);
xor U19928 (N_19928,N_19587,N_19782);
nand U19929 (N_19929,N_19542,N_19514);
or U19930 (N_19930,N_19616,N_19545);
nand U19931 (N_19931,N_19586,N_19669);
xor U19932 (N_19932,N_19759,N_19529);
nor U19933 (N_19933,N_19612,N_19701);
nor U19934 (N_19934,N_19674,N_19504);
nand U19935 (N_19935,N_19643,N_19713);
nand U19936 (N_19936,N_19726,N_19570);
or U19937 (N_19937,N_19707,N_19715);
xor U19938 (N_19938,N_19650,N_19568);
nor U19939 (N_19939,N_19690,N_19774);
or U19940 (N_19940,N_19617,N_19742);
or U19941 (N_19941,N_19660,N_19610);
nor U19942 (N_19942,N_19793,N_19659);
nand U19943 (N_19943,N_19771,N_19702);
and U19944 (N_19944,N_19613,N_19749);
nor U19945 (N_19945,N_19500,N_19760);
nand U19946 (N_19946,N_19680,N_19752);
nand U19947 (N_19947,N_19787,N_19757);
or U19948 (N_19948,N_19552,N_19738);
and U19949 (N_19949,N_19625,N_19515);
nand U19950 (N_19950,N_19676,N_19587);
nand U19951 (N_19951,N_19674,N_19508);
or U19952 (N_19952,N_19556,N_19521);
xnor U19953 (N_19953,N_19616,N_19742);
and U19954 (N_19954,N_19726,N_19602);
nor U19955 (N_19955,N_19767,N_19749);
nand U19956 (N_19956,N_19764,N_19758);
and U19957 (N_19957,N_19558,N_19691);
xor U19958 (N_19958,N_19686,N_19549);
xnor U19959 (N_19959,N_19590,N_19743);
xnor U19960 (N_19960,N_19689,N_19701);
nand U19961 (N_19961,N_19705,N_19696);
xnor U19962 (N_19962,N_19578,N_19661);
nor U19963 (N_19963,N_19780,N_19610);
or U19964 (N_19964,N_19702,N_19533);
nor U19965 (N_19965,N_19599,N_19577);
nor U19966 (N_19966,N_19654,N_19501);
nand U19967 (N_19967,N_19503,N_19558);
and U19968 (N_19968,N_19514,N_19633);
and U19969 (N_19969,N_19588,N_19640);
nor U19970 (N_19970,N_19651,N_19622);
nor U19971 (N_19971,N_19683,N_19744);
and U19972 (N_19972,N_19765,N_19501);
or U19973 (N_19973,N_19652,N_19519);
or U19974 (N_19974,N_19787,N_19732);
and U19975 (N_19975,N_19685,N_19688);
nor U19976 (N_19976,N_19653,N_19554);
nand U19977 (N_19977,N_19651,N_19781);
xnor U19978 (N_19978,N_19701,N_19733);
nand U19979 (N_19979,N_19759,N_19752);
xnor U19980 (N_19980,N_19535,N_19667);
and U19981 (N_19981,N_19679,N_19564);
nand U19982 (N_19982,N_19739,N_19656);
xor U19983 (N_19983,N_19713,N_19638);
nor U19984 (N_19984,N_19693,N_19518);
and U19985 (N_19985,N_19725,N_19534);
nor U19986 (N_19986,N_19543,N_19586);
or U19987 (N_19987,N_19685,N_19566);
nand U19988 (N_19988,N_19701,N_19725);
nand U19989 (N_19989,N_19666,N_19684);
xor U19990 (N_19990,N_19621,N_19565);
nand U19991 (N_19991,N_19680,N_19551);
nor U19992 (N_19992,N_19505,N_19568);
xnor U19993 (N_19993,N_19796,N_19518);
and U19994 (N_19994,N_19579,N_19791);
nand U19995 (N_19995,N_19587,N_19740);
and U19996 (N_19996,N_19580,N_19784);
and U19997 (N_19997,N_19716,N_19744);
and U19998 (N_19998,N_19549,N_19544);
and U19999 (N_19999,N_19516,N_19640);
nor U20000 (N_20000,N_19698,N_19793);
and U20001 (N_20001,N_19793,N_19674);
and U20002 (N_20002,N_19691,N_19710);
or U20003 (N_20003,N_19639,N_19582);
nand U20004 (N_20004,N_19510,N_19649);
xnor U20005 (N_20005,N_19620,N_19679);
nand U20006 (N_20006,N_19703,N_19771);
xor U20007 (N_20007,N_19627,N_19683);
xor U20008 (N_20008,N_19603,N_19725);
and U20009 (N_20009,N_19785,N_19588);
nand U20010 (N_20010,N_19662,N_19618);
nor U20011 (N_20011,N_19757,N_19551);
nand U20012 (N_20012,N_19551,N_19707);
nand U20013 (N_20013,N_19508,N_19687);
xnor U20014 (N_20014,N_19502,N_19668);
and U20015 (N_20015,N_19746,N_19511);
xor U20016 (N_20016,N_19629,N_19600);
nand U20017 (N_20017,N_19637,N_19758);
xor U20018 (N_20018,N_19514,N_19599);
xnor U20019 (N_20019,N_19606,N_19654);
xor U20020 (N_20020,N_19619,N_19618);
nor U20021 (N_20021,N_19764,N_19793);
nor U20022 (N_20022,N_19762,N_19600);
xnor U20023 (N_20023,N_19535,N_19767);
and U20024 (N_20024,N_19538,N_19687);
or U20025 (N_20025,N_19722,N_19759);
xor U20026 (N_20026,N_19654,N_19623);
nor U20027 (N_20027,N_19670,N_19529);
nor U20028 (N_20028,N_19552,N_19786);
nor U20029 (N_20029,N_19523,N_19701);
or U20030 (N_20030,N_19783,N_19564);
xor U20031 (N_20031,N_19541,N_19570);
nor U20032 (N_20032,N_19596,N_19600);
and U20033 (N_20033,N_19713,N_19712);
or U20034 (N_20034,N_19581,N_19771);
nor U20035 (N_20035,N_19608,N_19602);
nor U20036 (N_20036,N_19762,N_19793);
and U20037 (N_20037,N_19593,N_19721);
or U20038 (N_20038,N_19501,N_19794);
or U20039 (N_20039,N_19670,N_19608);
nand U20040 (N_20040,N_19708,N_19607);
or U20041 (N_20041,N_19599,N_19527);
xor U20042 (N_20042,N_19698,N_19554);
xnor U20043 (N_20043,N_19610,N_19701);
xnor U20044 (N_20044,N_19783,N_19793);
nor U20045 (N_20045,N_19663,N_19678);
and U20046 (N_20046,N_19605,N_19731);
nor U20047 (N_20047,N_19651,N_19524);
nand U20048 (N_20048,N_19700,N_19510);
or U20049 (N_20049,N_19603,N_19772);
nand U20050 (N_20050,N_19698,N_19590);
or U20051 (N_20051,N_19775,N_19753);
and U20052 (N_20052,N_19686,N_19735);
and U20053 (N_20053,N_19558,N_19759);
nor U20054 (N_20054,N_19632,N_19528);
nand U20055 (N_20055,N_19793,N_19630);
nor U20056 (N_20056,N_19526,N_19687);
nor U20057 (N_20057,N_19631,N_19514);
xor U20058 (N_20058,N_19574,N_19718);
or U20059 (N_20059,N_19686,N_19527);
nor U20060 (N_20060,N_19770,N_19573);
or U20061 (N_20061,N_19534,N_19509);
and U20062 (N_20062,N_19545,N_19695);
xnor U20063 (N_20063,N_19669,N_19752);
xnor U20064 (N_20064,N_19601,N_19586);
or U20065 (N_20065,N_19629,N_19618);
xnor U20066 (N_20066,N_19670,N_19646);
and U20067 (N_20067,N_19717,N_19629);
nand U20068 (N_20068,N_19623,N_19548);
nor U20069 (N_20069,N_19608,N_19586);
nand U20070 (N_20070,N_19798,N_19508);
nand U20071 (N_20071,N_19588,N_19674);
or U20072 (N_20072,N_19640,N_19548);
nand U20073 (N_20073,N_19502,N_19554);
or U20074 (N_20074,N_19599,N_19690);
or U20075 (N_20075,N_19660,N_19547);
nand U20076 (N_20076,N_19667,N_19655);
xnor U20077 (N_20077,N_19730,N_19614);
nand U20078 (N_20078,N_19699,N_19638);
nand U20079 (N_20079,N_19719,N_19507);
xnor U20080 (N_20080,N_19670,N_19749);
nand U20081 (N_20081,N_19770,N_19650);
xor U20082 (N_20082,N_19770,N_19772);
xor U20083 (N_20083,N_19641,N_19537);
xor U20084 (N_20084,N_19577,N_19610);
nand U20085 (N_20085,N_19787,N_19516);
xor U20086 (N_20086,N_19711,N_19629);
and U20087 (N_20087,N_19572,N_19674);
nor U20088 (N_20088,N_19715,N_19614);
or U20089 (N_20089,N_19675,N_19543);
or U20090 (N_20090,N_19714,N_19614);
nand U20091 (N_20091,N_19576,N_19669);
xnor U20092 (N_20092,N_19783,N_19688);
xor U20093 (N_20093,N_19617,N_19772);
or U20094 (N_20094,N_19747,N_19682);
or U20095 (N_20095,N_19717,N_19675);
xnor U20096 (N_20096,N_19747,N_19678);
xor U20097 (N_20097,N_19783,N_19610);
or U20098 (N_20098,N_19661,N_19534);
nand U20099 (N_20099,N_19703,N_19648);
nand U20100 (N_20100,N_19953,N_19980);
nor U20101 (N_20101,N_19960,N_19868);
nand U20102 (N_20102,N_20030,N_20058);
nand U20103 (N_20103,N_19928,N_19869);
or U20104 (N_20104,N_20070,N_19992);
nand U20105 (N_20105,N_19825,N_19888);
and U20106 (N_20106,N_20063,N_19937);
nand U20107 (N_20107,N_19801,N_20002);
or U20108 (N_20108,N_19856,N_19899);
nor U20109 (N_20109,N_19912,N_19995);
xor U20110 (N_20110,N_20007,N_20031);
and U20111 (N_20111,N_19982,N_20016);
or U20112 (N_20112,N_19839,N_19941);
nor U20113 (N_20113,N_19966,N_20073);
and U20114 (N_20114,N_20066,N_19885);
or U20115 (N_20115,N_19977,N_19927);
xnor U20116 (N_20116,N_20088,N_20005);
nand U20117 (N_20117,N_19851,N_19858);
xor U20118 (N_20118,N_19942,N_20082);
xor U20119 (N_20119,N_20013,N_19866);
xnor U20120 (N_20120,N_19891,N_19906);
and U20121 (N_20121,N_20068,N_19974);
nand U20122 (N_20122,N_19932,N_20062);
and U20123 (N_20123,N_19901,N_19809);
nand U20124 (N_20124,N_20095,N_19848);
xor U20125 (N_20125,N_20094,N_20035);
xor U20126 (N_20126,N_19894,N_19917);
nand U20127 (N_20127,N_19857,N_20099);
nand U20128 (N_20128,N_19827,N_19926);
and U20129 (N_20129,N_19908,N_19859);
and U20130 (N_20130,N_20026,N_19838);
nor U20131 (N_20131,N_19998,N_19824);
or U20132 (N_20132,N_19930,N_19812);
nor U20133 (N_20133,N_19915,N_19996);
nand U20134 (N_20134,N_19940,N_20050);
xor U20135 (N_20135,N_20064,N_20004);
nand U20136 (N_20136,N_19831,N_20049);
or U20137 (N_20137,N_20053,N_19979);
or U20138 (N_20138,N_19889,N_20020);
or U20139 (N_20139,N_19890,N_19882);
xnor U20140 (N_20140,N_19842,N_19808);
or U20141 (N_20141,N_20047,N_20079);
and U20142 (N_20142,N_20028,N_19962);
nand U20143 (N_20143,N_19922,N_19989);
nand U20144 (N_20144,N_19870,N_20033);
or U20145 (N_20145,N_20039,N_19903);
nand U20146 (N_20146,N_20097,N_19957);
nor U20147 (N_20147,N_20011,N_19850);
and U20148 (N_20148,N_20086,N_19916);
nand U20149 (N_20149,N_19909,N_19833);
or U20150 (N_20150,N_19892,N_19884);
nand U20151 (N_20151,N_19990,N_20021);
or U20152 (N_20152,N_20077,N_19847);
and U20153 (N_20153,N_19821,N_20076);
and U20154 (N_20154,N_19984,N_20008);
and U20155 (N_20155,N_19958,N_19867);
nor U20156 (N_20156,N_19835,N_19871);
xnor U20157 (N_20157,N_19967,N_19810);
and U20158 (N_20158,N_20009,N_20080);
nor U20159 (N_20159,N_19836,N_19852);
xnor U20160 (N_20160,N_19849,N_19804);
nand U20161 (N_20161,N_19945,N_19846);
nor U20162 (N_20162,N_19970,N_19834);
nand U20163 (N_20163,N_19875,N_20018);
nand U20164 (N_20164,N_19929,N_20074);
nand U20165 (N_20165,N_20041,N_19923);
nor U20166 (N_20166,N_19806,N_20061);
and U20167 (N_20167,N_19904,N_19818);
nand U20168 (N_20168,N_19947,N_19861);
and U20169 (N_20169,N_20036,N_19931);
xnor U20170 (N_20170,N_19817,N_19919);
and U20171 (N_20171,N_20022,N_19955);
or U20172 (N_20172,N_19981,N_19803);
nand U20173 (N_20173,N_19883,N_19999);
nor U20174 (N_20174,N_20089,N_19972);
nand U20175 (N_20175,N_19952,N_20081);
or U20176 (N_20176,N_19820,N_19959);
or U20177 (N_20177,N_20083,N_20059);
or U20178 (N_20178,N_19815,N_20046);
or U20179 (N_20179,N_19860,N_20045);
and U20180 (N_20180,N_19880,N_19874);
xnor U20181 (N_20181,N_19965,N_20037);
or U20182 (N_20182,N_19898,N_20014);
and U20183 (N_20183,N_19865,N_19934);
nand U20184 (N_20184,N_19924,N_19936);
nand U20185 (N_20185,N_19921,N_19954);
nand U20186 (N_20186,N_19956,N_19897);
and U20187 (N_20187,N_20017,N_20051);
and U20188 (N_20188,N_19991,N_20092);
or U20189 (N_20189,N_20048,N_19879);
nand U20190 (N_20190,N_19983,N_20024);
nand U20191 (N_20191,N_20091,N_19939);
nand U20192 (N_20192,N_20042,N_20010);
or U20193 (N_20193,N_19807,N_19948);
nand U20194 (N_20194,N_19905,N_20025);
nand U20195 (N_20195,N_19819,N_20096);
and U20196 (N_20196,N_19896,N_19895);
xor U20197 (N_20197,N_19853,N_19822);
or U20198 (N_20198,N_19826,N_19800);
nand U20199 (N_20199,N_19968,N_19855);
nor U20200 (N_20200,N_20075,N_19976);
nand U20201 (N_20201,N_20056,N_20090);
xnor U20202 (N_20202,N_20078,N_19878);
and U20203 (N_20203,N_19811,N_19832);
or U20204 (N_20204,N_19925,N_19914);
or U20205 (N_20205,N_19910,N_19862);
and U20206 (N_20206,N_20060,N_19872);
nand U20207 (N_20207,N_19877,N_19950);
and U20208 (N_20208,N_20044,N_19802);
and U20209 (N_20209,N_20003,N_19814);
nand U20210 (N_20210,N_19828,N_19913);
nand U20211 (N_20211,N_20043,N_19902);
or U20212 (N_20212,N_19837,N_19911);
or U20213 (N_20213,N_20055,N_19844);
or U20214 (N_20214,N_19951,N_19943);
nand U20215 (N_20215,N_20006,N_20071);
or U20216 (N_20216,N_20023,N_20069);
or U20217 (N_20217,N_20065,N_19907);
and U20218 (N_20218,N_20038,N_19971);
and U20219 (N_20219,N_19944,N_20072);
nor U20220 (N_20220,N_20012,N_19816);
and U20221 (N_20221,N_19978,N_20067);
or U20222 (N_20222,N_19994,N_19863);
or U20223 (N_20223,N_20052,N_20087);
xor U20224 (N_20224,N_19841,N_19938);
xnor U20225 (N_20225,N_20029,N_19993);
or U20226 (N_20226,N_19986,N_20040);
nand U20227 (N_20227,N_19918,N_19840);
xor U20228 (N_20228,N_19975,N_19933);
and U20229 (N_20229,N_19997,N_19829);
nor U20230 (N_20230,N_19876,N_19946);
nand U20231 (N_20231,N_19813,N_19881);
nor U20232 (N_20232,N_19854,N_20001);
nand U20233 (N_20233,N_19920,N_20034);
or U20234 (N_20234,N_19987,N_19843);
xnor U20235 (N_20235,N_19988,N_19823);
nor U20236 (N_20236,N_19961,N_20098);
nand U20237 (N_20237,N_20019,N_19893);
xnor U20238 (N_20238,N_20057,N_19864);
and U20239 (N_20239,N_19964,N_20027);
nand U20240 (N_20240,N_19886,N_20032);
or U20241 (N_20241,N_20015,N_19935);
or U20242 (N_20242,N_20054,N_19963);
and U20243 (N_20243,N_19969,N_19900);
nand U20244 (N_20244,N_19973,N_19845);
nor U20245 (N_20245,N_20000,N_19985);
and U20246 (N_20246,N_19805,N_20093);
and U20247 (N_20247,N_20085,N_19887);
xor U20248 (N_20248,N_19949,N_20084);
or U20249 (N_20249,N_19830,N_19873);
nor U20250 (N_20250,N_19975,N_19831);
or U20251 (N_20251,N_20010,N_20064);
nand U20252 (N_20252,N_20016,N_20079);
nand U20253 (N_20253,N_19880,N_19868);
and U20254 (N_20254,N_19927,N_19961);
and U20255 (N_20255,N_19990,N_19841);
and U20256 (N_20256,N_19967,N_20077);
or U20257 (N_20257,N_19983,N_20069);
nor U20258 (N_20258,N_20066,N_19887);
or U20259 (N_20259,N_19912,N_19833);
xnor U20260 (N_20260,N_19821,N_20020);
and U20261 (N_20261,N_20096,N_20016);
nand U20262 (N_20262,N_19865,N_20077);
or U20263 (N_20263,N_19817,N_20068);
xor U20264 (N_20264,N_20085,N_20098);
nor U20265 (N_20265,N_20031,N_20013);
xor U20266 (N_20266,N_20047,N_20061);
xnor U20267 (N_20267,N_19905,N_19836);
nand U20268 (N_20268,N_19825,N_19949);
xor U20269 (N_20269,N_20079,N_20004);
and U20270 (N_20270,N_19806,N_20001);
xor U20271 (N_20271,N_20043,N_20022);
xor U20272 (N_20272,N_19997,N_19962);
nand U20273 (N_20273,N_19947,N_19851);
nor U20274 (N_20274,N_19952,N_20034);
and U20275 (N_20275,N_20072,N_19876);
xnor U20276 (N_20276,N_19913,N_19997);
or U20277 (N_20277,N_20098,N_19998);
nand U20278 (N_20278,N_20089,N_19963);
nor U20279 (N_20279,N_20081,N_19883);
or U20280 (N_20280,N_20066,N_20064);
or U20281 (N_20281,N_19833,N_19928);
nand U20282 (N_20282,N_19953,N_19899);
and U20283 (N_20283,N_19896,N_19930);
and U20284 (N_20284,N_19851,N_19822);
nor U20285 (N_20285,N_19995,N_19872);
or U20286 (N_20286,N_19906,N_19876);
nand U20287 (N_20287,N_19891,N_19920);
xor U20288 (N_20288,N_19946,N_20075);
nor U20289 (N_20289,N_19851,N_20004);
xnor U20290 (N_20290,N_20027,N_20049);
nor U20291 (N_20291,N_19823,N_19989);
nor U20292 (N_20292,N_19858,N_19952);
and U20293 (N_20293,N_19876,N_20021);
xnor U20294 (N_20294,N_19917,N_19912);
nor U20295 (N_20295,N_20035,N_19944);
nor U20296 (N_20296,N_19963,N_20063);
and U20297 (N_20297,N_19834,N_20065);
nor U20298 (N_20298,N_20077,N_20024);
or U20299 (N_20299,N_20080,N_20096);
or U20300 (N_20300,N_19806,N_19970);
and U20301 (N_20301,N_19880,N_19948);
xnor U20302 (N_20302,N_19813,N_19849);
nand U20303 (N_20303,N_19900,N_19822);
nand U20304 (N_20304,N_20067,N_20003);
nand U20305 (N_20305,N_19892,N_19857);
or U20306 (N_20306,N_20013,N_19836);
or U20307 (N_20307,N_19921,N_19937);
or U20308 (N_20308,N_19976,N_19895);
nand U20309 (N_20309,N_19880,N_20033);
xor U20310 (N_20310,N_20030,N_19980);
or U20311 (N_20311,N_20091,N_20039);
nand U20312 (N_20312,N_19832,N_19813);
and U20313 (N_20313,N_20046,N_19889);
or U20314 (N_20314,N_20055,N_20058);
and U20315 (N_20315,N_20081,N_19829);
nor U20316 (N_20316,N_19860,N_20070);
or U20317 (N_20317,N_19987,N_19982);
and U20318 (N_20318,N_20024,N_19948);
xor U20319 (N_20319,N_19834,N_19924);
nor U20320 (N_20320,N_19814,N_19968);
and U20321 (N_20321,N_19922,N_19881);
xnor U20322 (N_20322,N_19831,N_19880);
and U20323 (N_20323,N_19832,N_19937);
and U20324 (N_20324,N_19991,N_19985);
and U20325 (N_20325,N_20099,N_19825);
or U20326 (N_20326,N_19906,N_19815);
and U20327 (N_20327,N_19975,N_19941);
xnor U20328 (N_20328,N_19909,N_19889);
nor U20329 (N_20329,N_19944,N_19837);
nor U20330 (N_20330,N_19960,N_19880);
or U20331 (N_20331,N_20014,N_20089);
nand U20332 (N_20332,N_20036,N_19948);
nand U20333 (N_20333,N_20047,N_19839);
and U20334 (N_20334,N_19919,N_20061);
xnor U20335 (N_20335,N_19836,N_19829);
nor U20336 (N_20336,N_19848,N_19936);
nor U20337 (N_20337,N_19946,N_19994);
or U20338 (N_20338,N_19920,N_19868);
and U20339 (N_20339,N_19890,N_19825);
xor U20340 (N_20340,N_19859,N_19846);
nand U20341 (N_20341,N_19882,N_20048);
and U20342 (N_20342,N_20081,N_19812);
xnor U20343 (N_20343,N_19889,N_19975);
and U20344 (N_20344,N_19823,N_19882);
nor U20345 (N_20345,N_19845,N_19827);
and U20346 (N_20346,N_19811,N_19840);
and U20347 (N_20347,N_20086,N_20058);
and U20348 (N_20348,N_19817,N_20037);
xnor U20349 (N_20349,N_19954,N_20009);
or U20350 (N_20350,N_19943,N_19835);
nand U20351 (N_20351,N_20079,N_19862);
xor U20352 (N_20352,N_19825,N_19942);
nand U20353 (N_20353,N_19967,N_19871);
and U20354 (N_20354,N_20010,N_19947);
and U20355 (N_20355,N_19996,N_19894);
and U20356 (N_20356,N_20083,N_19847);
nand U20357 (N_20357,N_20067,N_19866);
or U20358 (N_20358,N_19984,N_20055);
nor U20359 (N_20359,N_19856,N_20038);
nand U20360 (N_20360,N_20085,N_20065);
and U20361 (N_20361,N_19848,N_20045);
or U20362 (N_20362,N_19986,N_19936);
nor U20363 (N_20363,N_20045,N_19976);
xnor U20364 (N_20364,N_19824,N_19884);
nor U20365 (N_20365,N_19807,N_20017);
and U20366 (N_20366,N_19848,N_19829);
nand U20367 (N_20367,N_19824,N_19962);
or U20368 (N_20368,N_20093,N_20084);
xnor U20369 (N_20369,N_19981,N_20067);
or U20370 (N_20370,N_19876,N_19886);
nor U20371 (N_20371,N_19893,N_19802);
and U20372 (N_20372,N_19838,N_20054);
xnor U20373 (N_20373,N_19841,N_19828);
xnor U20374 (N_20374,N_19952,N_20063);
or U20375 (N_20375,N_19875,N_20044);
xor U20376 (N_20376,N_19875,N_19962);
xor U20377 (N_20377,N_19842,N_20099);
xnor U20378 (N_20378,N_19903,N_19846);
or U20379 (N_20379,N_19828,N_19877);
and U20380 (N_20380,N_19966,N_19823);
xnor U20381 (N_20381,N_20003,N_19906);
nand U20382 (N_20382,N_19990,N_19994);
nand U20383 (N_20383,N_19961,N_19910);
nor U20384 (N_20384,N_20010,N_19945);
and U20385 (N_20385,N_19954,N_19878);
or U20386 (N_20386,N_20093,N_19906);
nand U20387 (N_20387,N_20090,N_19941);
xnor U20388 (N_20388,N_19800,N_20010);
or U20389 (N_20389,N_19843,N_20036);
and U20390 (N_20390,N_19934,N_20098);
xor U20391 (N_20391,N_19990,N_20042);
xnor U20392 (N_20392,N_19906,N_19836);
nand U20393 (N_20393,N_19967,N_20074);
and U20394 (N_20394,N_19924,N_19896);
and U20395 (N_20395,N_19812,N_20019);
nor U20396 (N_20396,N_19810,N_19902);
and U20397 (N_20397,N_20072,N_19969);
nor U20398 (N_20398,N_19843,N_19809);
nand U20399 (N_20399,N_20094,N_19855);
nor U20400 (N_20400,N_20108,N_20321);
or U20401 (N_20401,N_20247,N_20398);
nand U20402 (N_20402,N_20155,N_20323);
nand U20403 (N_20403,N_20234,N_20113);
nor U20404 (N_20404,N_20236,N_20370);
nor U20405 (N_20405,N_20230,N_20166);
or U20406 (N_20406,N_20156,N_20190);
nor U20407 (N_20407,N_20202,N_20293);
nand U20408 (N_20408,N_20272,N_20248);
nor U20409 (N_20409,N_20197,N_20298);
nand U20410 (N_20410,N_20267,N_20210);
and U20411 (N_20411,N_20384,N_20393);
and U20412 (N_20412,N_20391,N_20180);
and U20413 (N_20413,N_20387,N_20324);
nand U20414 (N_20414,N_20304,N_20149);
or U20415 (N_20415,N_20366,N_20131);
or U20416 (N_20416,N_20227,N_20303);
xnor U20417 (N_20417,N_20151,N_20306);
nor U20418 (N_20418,N_20317,N_20237);
or U20419 (N_20419,N_20318,N_20231);
xor U20420 (N_20420,N_20390,N_20169);
and U20421 (N_20421,N_20283,N_20235);
nor U20422 (N_20422,N_20107,N_20146);
and U20423 (N_20423,N_20159,N_20208);
and U20424 (N_20424,N_20117,N_20338);
and U20425 (N_20425,N_20364,N_20171);
nand U20426 (N_20426,N_20377,N_20212);
or U20427 (N_20427,N_20359,N_20320);
xor U20428 (N_20428,N_20194,N_20204);
xnor U20429 (N_20429,N_20290,N_20136);
xor U20430 (N_20430,N_20285,N_20106);
and U20431 (N_20431,N_20329,N_20191);
xor U20432 (N_20432,N_20144,N_20174);
and U20433 (N_20433,N_20183,N_20223);
nand U20434 (N_20434,N_20240,N_20369);
nor U20435 (N_20435,N_20116,N_20375);
xnor U20436 (N_20436,N_20340,N_20343);
nand U20437 (N_20437,N_20326,N_20265);
or U20438 (N_20438,N_20309,N_20362);
xnor U20439 (N_20439,N_20308,N_20284);
and U20440 (N_20440,N_20262,N_20104);
xnor U20441 (N_20441,N_20275,N_20258);
nand U20442 (N_20442,N_20256,N_20115);
nor U20443 (N_20443,N_20335,N_20311);
xnor U20444 (N_20444,N_20389,N_20316);
nand U20445 (N_20445,N_20198,N_20216);
and U20446 (N_20446,N_20342,N_20182);
xnor U20447 (N_20447,N_20280,N_20121);
nand U20448 (N_20448,N_20167,N_20192);
xor U20449 (N_20449,N_20297,N_20196);
xor U20450 (N_20450,N_20336,N_20181);
or U20451 (N_20451,N_20118,N_20372);
or U20452 (N_20452,N_20138,N_20382);
nor U20453 (N_20453,N_20360,N_20385);
nor U20454 (N_20454,N_20242,N_20367);
or U20455 (N_20455,N_20341,N_20352);
or U20456 (N_20456,N_20220,N_20246);
nand U20457 (N_20457,N_20112,N_20257);
or U20458 (N_20458,N_20140,N_20289);
or U20459 (N_20459,N_20111,N_20282);
nand U20460 (N_20460,N_20383,N_20379);
and U20461 (N_20461,N_20261,N_20250);
and U20462 (N_20462,N_20253,N_20310);
or U20463 (N_20463,N_20294,N_20357);
or U20464 (N_20464,N_20354,N_20137);
nor U20465 (N_20465,N_20243,N_20126);
nand U20466 (N_20466,N_20207,N_20133);
xnor U20467 (N_20467,N_20187,N_20193);
nor U20468 (N_20468,N_20160,N_20353);
nand U20469 (N_20469,N_20244,N_20346);
or U20470 (N_20470,N_20270,N_20120);
or U20471 (N_20471,N_20328,N_20268);
nand U20472 (N_20472,N_20313,N_20214);
nand U20473 (N_20473,N_20200,N_20170);
xnor U20474 (N_20474,N_20228,N_20276);
nand U20475 (N_20475,N_20148,N_20176);
nor U20476 (N_20476,N_20172,N_20373);
and U20477 (N_20477,N_20397,N_20251);
xnor U20478 (N_20478,N_20396,N_20333);
xnor U20479 (N_20479,N_20150,N_20239);
nor U20480 (N_20480,N_20299,N_20100);
nand U20481 (N_20481,N_20245,N_20332);
nand U20482 (N_20482,N_20269,N_20205);
nand U20483 (N_20483,N_20296,N_20361);
and U20484 (N_20484,N_20273,N_20386);
xnor U20485 (N_20485,N_20162,N_20399);
or U20486 (N_20486,N_20134,N_20222);
nor U20487 (N_20487,N_20163,N_20233);
and U20488 (N_20488,N_20209,N_20254);
and U20489 (N_20489,N_20288,N_20186);
nor U20490 (N_20490,N_20266,N_20132);
and U20491 (N_20491,N_20103,N_20219);
xor U20492 (N_20492,N_20154,N_20394);
or U20493 (N_20493,N_20314,N_20221);
or U20494 (N_20494,N_20334,N_20135);
nor U20495 (N_20495,N_20215,N_20392);
nor U20496 (N_20496,N_20125,N_20277);
nand U20497 (N_20497,N_20128,N_20179);
xor U20498 (N_20498,N_20381,N_20337);
nor U20499 (N_20499,N_20229,N_20292);
or U20500 (N_20500,N_20119,N_20129);
and U20501 (N_20501,N_20226,N_20143);
and U20502 (N_20502,N_20175,N_20201);
or U20503 (N_20503,N_20165,N_20300);
xor U20504 (N_20504,N_20114,N_20139);
nand U20505 (N_20505,N_20152,N_20278);
xnor U20506 (N_20506,N_20161,N_20315);
nand U20507 (N_20507,N_20350,N_20213);
nand U20508 (N_20508,N_20274,N_20358);
or U20509 (N_20509,N_20348,N_20339);
or U20510 (N_20510,N_20302,N_20218);
xnor U20511 (N_20511,N_20264,N_20141);
nand U20512 (N_20512,N_20349,N_20363);
or U20513 (N_20513,N_20286,N_20355);
or U20514 (N_20514,N_20388,N_20206);
and U20515 (N_20515,N_20241,N_20351);
nor U20516 (N_20516,N_20344,N_20177);
and U20517 (N_20517,N_20153,N_20158);
xor U20518 (N_20518,N_20287,N_20380);
or U20519 (N_20519,N_20189,N_20305);
nand U20520 (N_20520,N_20249,N_20188);
and U20521 (N_20521,N_20295,N_20356);
nor U20522 (N_20522,N_20259,N_20238);
and U20523 (N_20523,N_20371,N_20203);
nor U20524 (N_20524,N_20365,N_20279);
nor U20525 (N_20525,N_20211,N_20173);
xnor U20526 (N_20526,N_20368,N_20345);
nand U20527 (N_20527,N_20327,N_20127);
nor U20528 (N_20528,N_20145,N_20232);
and U20529 (N_20529,N_20124,N_20281);
nor U20530 (N_20530,N_20319,N_20185);
or U20531 (N_20531,N_20252,N_20378);
nand U20532 (N_20532,N_20168,N_20110);
xnor U20533 (N_20533,N_20347,N_20178);
nor U20534 (N_20534,N_20184,N_20331);
nand U20535 (N_20535,N_20142,N_20109);
nor U20536 (N_20536,N_20105,N_20224);
nor U20537 (N_20537,N_20102,N_20157);
nor U20538 (N_20538,N_20199,N_20307);
nor U20539 (N_20539,N_20164,N_20330);
nand U20540 (N_20540,N_20395,N_20147);
xor U20541 (N_20541,N_20130,N_20195);
nor U20542 (N_20542,N_20263,N_20271);
nand U20543 (N_20543,N_20225,N_20322);
or U20544 (N_20544,N_20122,N_20101);
nand U20545 (N_20545,N_20255,N_20376);
xor U20546 (N_20546,N_20325,N_20123);
and U20547 (N_20547,N_20291,N_20374);
or U20548 (N_20548,N_20312,N_20260);
nor U20549 (N_20549,N_20301,N_20217);
nand U20550 (N_20550,N_20170,N_20224);
and U20551 (N_20551,N_20239,N_20381);
nor U20552 (N_20552,N_20362,N_20213);
nand U20553 (N_20553,N_20144,N_20365);
or U20554 (N_20554,N_20370,N_20142);
nand U20555 (N_20555,N_20305,N_20244);
xor U20556 (N_20556,N_20168,N_20104);
xor U20557 (N_20557,N_20214,N_20126);
or U20558 (N_20558,N_20103,N_20291);
or U20559 (N_20559,N_20156,N_20376);
xor U20560 (N_20560,N_20221,N_20156);
and U20561 (N_20561,N_20297,N_20240);
and U20562 (N_20562,N_20135,N_20227);
nand U20563 (N_20563,N_20156,N_20148);
xnor U20564 (N_20564,N_20166,N_20125);
nor U20565 (N_20565,N_20164,N_20204);
or U20566 (N_20566,N_20102,N_20120);
nor U20567 (N_20567,N_20242,N_20347);
or U20568 (N_20568,N_20322,N_20184);
nand U20569 (N_20569,N_20389,N_20358);
nand U20570 (N_20570,N_20159,N_20363);
nand U20571 (N_20571,N_20225,N_20154);
or U20572 (N_20572,N_20130,N_20274);
or U20573 (N_20573,N_20371,N_20218);
nand U20574 (N_20574,N_20111,N_20380);
nor U20575 (N_20575,N_20315,N_20391);
or U20576 (N_20576,N_20273,N_20345);
nor U20577 (N_20577,N_20182,N_20339);
and U20578 (N_20578,N_20295,N_20360);
nor U20579 (N_20579,N_20281,N_20295);
nor U20580 (N_20580,N_20217,N_20102);
nand U20581 (N_20581,N_20398,N_20228);
and U20582 (N_20582,N_20307,N_20156);
nand U20583 (N_20583,N_20226,N_20377);
or U20584 (N_20584,N_20385,N_20128);
xnor U20585 (N_20585,N_20115,N_20370);
nor U20586 (N_20586,N_20354,N_20304);
xor U20587 (N_20587,N_20151,N_20335);
and U20588 (N_20588,N_20226,N_20246);
xor U20589 (N_20589,N_20199,N_20244);
nor U20590 (N_20590,N_20168,N_20131);
xor U20591 (N_20591,N_20275,N_20336);
nor U20592 (N_20592,N_20161,N_20203);
or U20593 (N_20593,N_20113,N_20191);
or U20594 (N_20594,N_20301,N_20318);
and U20595 (N_20595,N_20158,N_20125);
or U20596 (N_20596,N_20291,N_20394);
and U20597 (N_20597,N_20383,N_20211);
nand U20598 (N_20598,N_20127,N_20215);
and U20599 (N_20599,N_20270,N_20362);
or U20600 (N_20600,N_20220,N_20335);
nand U20601 (N_20601,N_20253,N_20271);
xnor U20602 (N_20602,N_20208,N_20101);
nand U20603 (N_20603,N_20348,N_20296);
xor U20604 (N_20604,N_20233,N_20360);
xor U20605 (N_20605,N_20205,N_20153);
or U20606 (N_20606,N_20113,N_20186);
xnor U20607 (N_20607,N_20109,N_20128);
or U20608 (N_20608,N_20293,N_20299);
nor U20609 (N_20609,N_20383,N_20199);
nand U20610 (N_20610,N_20260,N_20378);
xor U20611 (N_20611,N_20175,N_20144);
xor U20612 (N_20612,N_20125,N_20317);
nor U20613 (N_20613,N_20345,N_20130);
and U20614 (N_20614,N_20338,N_20106);
or U20615 (N_20615,N_20139,N_20240);
nor U20616 (N_20616,N_20109,N_20310);
xnor U20617 (N_20617,N_20363,N_20395);
nor U20618 (N_20618,N_20173,N_20342);
and U20619 (N_20619,N_20158,N_20135);
nand U20620 (N_20620,N_20210,N_20234);
nand U20621 (N_20621,N_20343,N_20146);
nor U20622 (N_20622,N_20297,N_20336);
xor U20623 (N_20623,N_20131,N_20248);
xnor U20624 (N_20624,N_20128,N_20309);
nand U20625 (N_20625,N_20244,N_20184);
nand U20626 (N_20626,N_20176,N_20336);
or U20627 (N_20627,N_20120,N_20244);
and U20628 (N_20628,N_20355,N_20102);
and U20629 (N_20629,N_20308,N_20288);
or U20630 (N_20630,N_20210,N_20336);
or U20631 (N_20631,N_20242,N_20231);
nor U20632 (N_20632,N_20130,N_20369);
and U20633 (N_20633,N_20191,N_20310);
nand U20634 (N_20634,N_20144,N_20351);
or U20635 (N_20635,N_20374,N_20367);
nor U20636 (N_20636,N_20284,N_20187);
nor U20637 (N_20637,N_20295,N_20365);
nor U20638 (N_20638,N_20348,N_20160);
nor U20639 (N_20639,N_20108,N_20132);
and U20640 (N_20640,N_20369,N_20206);
or U20641 (N_20641,N_20254,N_20155);
and U20642 (N_20642,N_20308,N_20344);
xnor U20643 (N_20643,N_20137,N_20286);
nand U20644 (N_20644,N_20216,N_20153);
and U20645 (N_20645,N_20234,N_20275);
or U20646 (N_20646,N_20322,N_20146);
nand U20647 (N_20647,N_20215,N_20160);
and U20648 (N_20648,N_20128,N_20237);
and U20649 (N_20649,N_20122,N_20321);
nand U20650 (N_20650,N_20219,N_20194);
and U20651 (N_20651,N_20364,N_20296);
and U20652 (N_20652,N_20358,N_20345);
and U20653 (N_20653,N_20258,N_20169);
and U20654 (N_20654,N_20129,N_20182);
nor U20655 (N_20655,N_20291,N_20181);
nor U20656 (N_20656,N_20257,N_20247);
or U20657 (N_20657,N_20183,N_20276);
nand U20658 (N_20658,N_20341,N_20201);
xnor U20659 (N_20659,N_20285,N_20333);
or U20660 (N_20660,N_20106,N_20365);
and U20661 (N_20661,N_20201,N_20120);
and U20662 (N_20662,N_20191,N_20352);
and U20663 (N_20663,N_20254,N_20359);
nand U20664 (N_20664,N_20356,N_20339);
xor U20665 (N_20665,N_20211,N_20282);
and U20666 (N_20666,N_20343,N_20176);
xor U20667 (N_20667,N_20306,N_20209);
nand U20668 (N_20668,N_20388,N_20284);
nand U20669 (N_20669,N_20361,N_20271);
xor U20670 (N_20670,N_20146,N_20171);
nor U20671 (N_20671,N_20354,N_20188);
and U20672 (N_20672,N_20351,N_20290);
xnor U20673 (N_20673,N_20113,N_20397);
nand U20674 (N_20674,N_20369,N_20132);
xor U20675 (N_20675,N_20333,N_20292);
nand U20676 (N_20676,N_20308,N_20121);
xor U20677 (N_20677,N_20225,N_20274);
xnor U20678 (N_20678,N_20299,N_20186);
nor U20679 (N_20679,N_20326,N_20249);
and U20680 (N_20680,N_20379,N_20317);
and U20681 (N_20681,N_20121,N_20109);
and U20682 (N_20682,N_20183,N_20279);
nand U20683 (N_20683,N_20141,N_20391);
nand U20684 (N_20684,N_20137,N_20133);
nor U20685 (N_20685,N_20326,N_20321);
xnor U20686 (N_20686,N_20179,N_20193);
xnor U20687 (N_20687,N_20355,N_20179);
xor U20688 (N_20688,N_20158,N_20106);
nor U20689 (N_20689,N_20138,N_20245);
nand U20690 (N_20690,N_20188,N_20181);
nor U20691 (N_20691,N_20356,N_20212);
nand U20692 (N_20692,N_20127,N_20214);
and U20693 (N_20693,N_20102,N_20267);
nor U20694 (N_20694,N_20369,N_20189);
xor U20695 (N_20695,N_20140,N_20399);
and U20696 (N_20696,N_20363,N_20117);
and U20697 (N_20697,N_20288,N_20336);
xor U20698 (N_20698,N_20356,N_20221);
and U20699 (N_20699,N_20176,N_20333);
nor U20700 (N_20700,N_20477,N_20506);
and U20701 (N_20701,N_20510,N_20433);
nor U20702 (N_20702,N_20613,N_20482);
nor U20703 (N_20703,N_20499,N_20413);
and U20704 (N_20704,N_20550,N_20484);
xor U20705 (N_20705,N_20622,N_20443);
nand U20706 (N_20706,N_20574,N_20528);
nand U20707 (N_20707,N_20578,N_20672);
and U20708 (N_20708,N_20480,N_20615);
nor U20709 (N_20709,N_20436,N_20617);
xnor U20710 (N_20710,N_20448,N_20524);
nand U20711 (N_20711,N_20669,N_20555);
nor U20712 (N_20712,N_20680,N_20463);
nand U20713 (N_20713,N_20556,N_20474);
nor U20714 (N_20714,N_20554,N_20415);
and U20715 (N_20715,N_20453,N_20561);
and U20716 (N_20716,N_20646,N_20469);
nor U20717 (N_20717,N_20599,N_20620);
nand U20718 (N_20718,N_20426,N_20640);
or U20719 (N_20719,N_20569,N_20481);
and U20720 (N_20720,N_20589,N_20546);
and U20721 (N_20721,N_20668,N_20661);
nand U20722 (N_20722,N_20438,N_20663);
nand U20723 (N_20723,N_20697,N_20414);
nand U20724 (N_20724,N_20494,N_20424);
xor U20725 (N_20725,N_20431,N_20648);
xor U20726 (N_20726,N_20532,N_20459);
or U20727 (N_20727,N_20408,N_20501);
or U20728 (N_20728,N_20434,N_20639);
nor U20729 (N_20729,N_20526,N_20525);
and U20730 (N_20730,N_20597,N_20608);
nor U20731 (N_20731,N_20652,N_20460);
and U20732 (N_20732,N_20507,N_20437);
nand U20733 (N_20733,N_20551,N_20473);
xor U20734 (N_20734,N_20432,N_20479);
or U20735 (N_20735,N_20455,N_20403);
and U20736 (N_20736,N_20618,N_20591);
nand U20737 (N_20737,N_20637,N_20512);
nor U20738 (N_20738,N_20660,N_20564);
and U20739 (N_20739,N_20496,N_20505);
nor U20740 (N_20740,N_20435,N_20404);
xor U20741 (N_20741,N_20575,N_20504);
and U20742 (N_20742,N_20596,N_20445);
nand U20743 (N_20743,N_20584,N_20544);
nand U20744 (N_20744,N_20513,N_20470);
or U20745 (N_20745,N_20425,N_20645);
xnor U20746 (N_20746,N_20486,N_20405);
and U20747 (N_20747,N_20664,N_20605);
nor U20748 (N_20748,N_20684,N_20542);
and U20749 (N_20749,N_20458,N_20671);
xor U20750 (N_20750,N_20489,N_20698);
nor U20751 (N_20751,N_20562,N_20503);
nor U20752 (N_20752,N_20412,N_20641);
nand U20753 (N_20753,N_20402,N_20603);
or U20754 (N_20754,N_20446,N_20611);
and U20755 (N_20755,N_20511,N_20590);
or U20756 (N_20756,N_20449,N_20457);
nor U20757 (N_20757,N_20647,N_20471);
nor U20758 (N_20758,N_20444,N_20509);
and U20759 (N_20759,N_20441,N_20665);
nor U20760 (N_20760,N_20515,N_20587);
nor U20761 (N_20761,N_20523,N_20682);
xnor U20762 (N_20762,N_20655,N_20518);
nor U20763 (N_20763,N_20514,N_20442);
nand U20764 (N_20764,N_20450,N_20558);
or U20765 (N_20765,N_20520,N_20440);
nor U20766 (N_20766,N_20519,N_20421);
nand U20767 (N_20767,N_20643,N_20585);
nand U20768 (N_20768,N_20530,N_20699);
or U20769 (N_20769,N_20418,N_20543);
nand U20770 (N_20770,N_20649,N_20577);
nor U20771 (N_20771,N_20540,N_20670);
nand U20772 (N_20772,N_20678,N_20635);
xor U20773 (N_20773,N_20686,N_20651);
nor U20774 (N_20774,N_20619,N_20553);
or U20775 (N_20775,N_20644,N_20508);
and U20776 (N_20776,N_20560,N_20409);
and U20777 (N_20777,N_20485,N_20656);
nor U20778 (N_20778,N_20488,N_20498);
xnor U20779 (N_20779,N_20439,N_20472);
and U20780 (N_20780,N_20552,N_20570);
nor U20781 (N_20781,N_20527,N_20493);
or U20782 (N_20782,N_20679,N_20583);
nor U20783 (N_20783,N_20634,N_20571);
xor U20784 (N_20784,N_20566,N_20568);
and U20785 (N_20785,N_20447,N_20567);
or U20786 (N_20786,N_20588,N_20491);
or U20787 (N_20787,N_20632,N_20423);
nand U20788 (N_20788,N_20522,N_20411);
and U20789 (N_20789,N_20630,N_20419);
nor U20790 (N_20790,N_20610,N_20676);
or U20791 (N_20791,N_20538,N_20406);
nor U20792 (N_20792,N_20629,N_20666);
or U20793 (N_20793,N_20606,N_20475);
and U20794 (N_20794,N_20691,N_20462);
xor U20795 (N_20795,N_20696,N_20539);
and U20796 (N_20796,N_20685,N_20690);
or U20797 (N_20797,N_20502,N_20549);
nand U20798 (N_20798,N_20427,N_20401);
xnor U20799 (N_20799,N_20616,N_20536);
or U20800 (N_20800,N_20674,N_20417);
and U20801 (N_20801,N_20683,N_20614);
nand U20802 (N_20802,N_20521,N_20428);
nor U20803 (N_20803,N_20478,N_20633);
or U20804 (N_20804,N_20600,N_20658);
and U20805 (N_20805,N_20500,N_20464);
nand U20806 (N_20806,N_20430,N_20429);
nor U20807 (N_20807,N_20592,N_20563);
nand U20808 (N_20808,N_20586,N_20454);
xor U20809 (N_20809,N_20534,N_20642);
xnor U20810 (N_20810,N_20681,N_20689);
xor U20811 (N_20811,N_20529,N_20497);
and U20812 (N_20812,N_20541,N_20487);
or U20813 (N_20813,N_20692,N_20595);
nand U20814 (N_20814,N_20545,N_20667);
nand U20815 (N_20815,N_20559,N_20609);
and U20816 (N_20816,N_20580,N_20407);
nand U20817 (N_20817,N_20516,N_20483);
nor U20818 (N_20818,N_20626,N_20531);
and U20819 (N_20819,N_20631,N_20422);
or U20820 (N_20820,N_20593,N_20657);
xnor U20821 (N_20821,N_20492,N_20625);
nand U20822 (N_20822,N_20579,N_20582);
xor U20823 (N_20823,N_20688,N_20604);
xor U20824 (N_20824,N_20565,N_20467);
nand U20825 (N_20825,N_20602,N_20420);
and U20826 (N_20826,N_20612,N_20410);
nor U20827 (N_20827,N_20400,N_20628);
or U20828 (N_20828,N_20621,N_20659);
xnor U20829 (N_20829,N_20476,N_20624);
nand U20830 (N_20830,N_20693,N_20572);
nor U20831 (N_20831,N_20677,N_20662);
nand U20832 (N_20832,N_20451,N_20638);
or U20833 (N_20833,N_20607,N_20694);
xor U20834 (N_20834,N_20495,N_20576);
and U20835 (N_20835,N_20653,N_20650);
xor U20836 (N_20836,N_20623,N_20675);
or U20837 (N_20837,N_20465,N_20695);
or U20838 (N_20838,N_20557,N_20627);
and U20839 (N_20839,N_20547,N_20573);
and U20840 (N_20840,N_20673,N_20452);
nor U20841 (N_20841,N_20466,N_20461);
nand U20842 (N_20842,N_20456,N_20636);
and U20843 (N_20843,N_20598,N_20416);
xnor U20844 (N_20844,N_20594,N_20490);
nand U20845 (N_20845,N_20581,N_20468);
nand U20846 (N_20846,N_20535,N_20654);
nor U20847 (N_20847,N_20687,N_20548);
nor U20848 (N_20848,N_20533,N_20601);
and U20849 (N_20849,N_20537,N_20517);
and U20850 (N_20850,N_20433,N_20644);
nor U20851 (N_20851,N_20461,N_20631);
xnor U20852 (N_20852,N_20643,N_20436);
xor U20853 (N_20853,N_20648,N_20592);
and U20854 (N_20854,N_20577,N_20483);
nand U20855 (N_20855,N_20408,N_20519);
xor U20856 (N_20856,N_20431,N_20485);
xnor U20857 (N_20857,N_20549,N_20626);
xnor U20858 (N_20858,N_20472,N_20512);
nor U20859 (N_20859,N_20437,N_20438);
and U20860 (N_20860,N_20541,N_20551);
nor U20861 (N_20861,N_20604,N_20487);
nand U20862 (N_20862,N_20468,N_20505);
nor U20863 (N_20863,N_20462,N_20432);
and U20864 (N_20864,N_20544,N_20551);
nor U20865 (N_20865,N_20560,N_20680);
and U20866 (N_20866,N_20611,N_20597);
nor U20867 (N_20867,N_20666,N_20578);
xor U20868 (N_20868,N_20416,N_20518);
nand U20869 (N_20869,N_20573,N_20500);
nand U20870 (N_20870,N_20607,N_20664);
nor U20871 (N_20871,N_20519,N_20676);
and U20872 (N_20872,N_20619,N_20511);
nor U20873 (N_20873,N_20512,N_20449);
and U20874 (N_20874,N_20677,N_20522);
nand U20875 (N_20875,N_20676,N_20564);
and U20876 (N_20876,N_20441,N_20444);
nor U20877 (N_20877,N_20680,N_20618);
and U20878 (N_20878,N_20556,N_20445);
nor U20879 (N_20879,N_20632,N_20655);
nor U20880 (N_20880,N_20427,N_20423);
nor U20881 (N_20881,N_20622,N_20570);
xnor U20882 (N_20882,N_20545,N_20482);
or U20883 (N_20883,N_20441,N_20427);
xor U20884 (N_20884,N_20673,N_20559);
nand U20885 (N_20885,N_20448,N_20539);
and U20886 (N_20886,N_20621,N_20634);
or U20887 (N_20887,N_20547,N_20565);
xnor U20888 (N_20888,N_20495,N_20554);
nor U20889 (N_20889,N_20631,N_20645);
nand U20890 (N_20890,N_20490,N_20652);
and U20891 (N_20891,N_20682,N_20580);
nor U20892 (N_20892,N_20590,N_20545);
and U20893 (N_20893,N_20524,N_20420);
or U20894 (N_20894,N_20467,N_20609);
nor U20895 (N_20895,N_20455,N_20665);
xor U20896 (N_20896,N_20621,N_20497);
nand U20897 (N_20897,N_20680,N_20454);
xor U20898 (N_20898,N_20409,N_20555);
xnor U20899 (N_20899,N_20494,N_20671);
and U20900 (N_20900,N_20414,N_20595);
and U20901 (N_20901,N_20468,N_20512);
or U20902 (N_20902,N_20510,N_20693);
nand U20903 (N_20903,N_20516,N_20502);
xor U20904 (N_20904,N_20593,N_20556);
and U20905 (N_20905,N_20616,N_20619);
and U20906 (N_20906,N_20635,N_20625);
and U20907 (N_20907,N_20605,N_20663);
nor U20908 (N_20908,N_20602,N_20514);
or U20909 (N_20909,N_20616,N_20548);
or U20910 (N_20910,N_20501,N_20637);
xnor U20911 (N_20911,N_20463,N_20557);
nor U20912 (N_20912,N_20510,N_20664);
nor U20913 (N_20913,N_20659,N_20488);
xor U20914 (N_20914,N_20647,N_20539);
nor U20915 (N_20915,N_20661,N_20629);
nand U20916 (N_20916,N_20467,N_20450);
xnor U20917 (N_20917,N_20619,N_20445);
nor U20918 (N_20918,N_20450,N_20486);
nor U20919 (N_20919,N_20639,N_20643);
nor U20920 (N_20920,N_20575,N_20472);
xnor U20921 (N_20921,N_20451,N_20403);
or U20922 (N_20922,N_20454,N_20611);
xnor U20923 (N_20923,N_20528,N_20579);
xor U20924 (N_20924,N_20447,N_20549);
nand U20925 (N_20925,N_20600,N_20626);
or U20926 (N_20926,N_20655,N_20606);
nand U20927 (N_20927,N_20500,N_20424);
nand U20928 (N_20928,N_20655,N_20625);
nand U20929 (N_20929,N_20410,N_20694);
and U20930 (N_20930,N_20603,N_20404);
and U20931 (N_20931,N_20600,N_20411);
nor U20932 (N_20932,N_20616,N_20620);
xor U20933 (N_20933,N_20490,N_20534);
nor U20934 (N_20934,N_20626,N_20680);
and U20935 (N_20935,N_20591,N_20622);
nor U20936 (N_20936,N_20482,N_20572);
and U20937 (N_20937,N_20567,N_20446);
nand U20938 (N_20938,N_20484,N_20410);
or U20939 (N_20939,N_20541,N_20500);
or U20940 (N_20940,N_20675,N_20426);
or U20941 (N_20941,N_20649,N_20501);
or U20942 (N_20942,N_20620,N_20631);
and U20943 (N_20943,N_20630,N_20589);
nor U20944 (N_20944,N_20699,N_20437);
or U20945 (N_20945,N_20584,N_20457);
nand U20946 (N_20946,N_20697,N_20638);
or U20947 (N_20947,N_20592,N_20486);
nor U20948 (N_20948,N_20548,N_20489);
nand U20949 (N_20949,N_20570,N_20563);
xnor U20950 (N_20950,N_20620,N_20649);
xor U20951 (N_20951,N_20549,N_20529);
nor U20952 (N_20952,N_20521,N_20652);
nor U20953 (N_20953,N_20523,N_20665);
or U20954 (N_20954,N_20520,N_20424);
and U20955 (N_20955,N_20530,N_20509);
xor U20956 (N_20956,N_20505,N_20669);
xor U20957 (N_20957,N_20540,N_20638);
or U20958 (N_20958,N_20594,N_20653);
nand U20959 (N_20959,N_20637,N_20655);
or U20960 (N_20960,N_20435,N_20553);
xnor U20961 (N_20961,N_20495,N_20521);
and U20962 (N_20962,N_20692,N_20680);
and U20963 (N_20963,N_20451,N_20491);
nand U20964 (N_20964,N_20501,N_20551);
nand U20965 (N_20965,N_20682,N_20495);
and U20966 (N_20966,N_20633,N_20695);
xor U20967 (N_20967,N_20697,N_20618);
nand U20968 (N_20968,N_20524,N_20687);
and U20969 (N_20969,N_20531,N_20616);
xor U20970 (N_20970,N_20429,N_20558);
xnor U20971 (N_20971,N_20403,N_20635);
xnor U20972 (N_20972,N_20572,N_20655);
nand U20973 (N_20973,N_20504,N_20506);
nor U20974 (N_20974,N_20423,N_20594);
nor U20975 (N_20975,N_20533,N_20490);
nor U20976 (N_20976,N_20562,N_20514);
nor U20977 (N_20977,N_20422,N_20455);
nor U20978 (N_20978,N_20464,N_20661);
xnor U20979 (N_20979,N_20497,N_20481);
xor U20980 (N_20980,N_20475,N_20476);
xnor U20981 (N_20981,N_20584,N_20496);
and U20982 (N_20982,N_20426,N_20462);
and U20983 (N_20983,N_20531,N_20534);
xor U20984 (N_20984,N_20656,N_20666);
nor U20985 (N_20985,N_20625,N_20557);
or U20986 (N_20986,N_20467,N_20695);
or U20987 (N_20987,N_20698,N_20446);
nand U20988 (N_20988,N_20629,N_20571);
or U20989 (N_20989,N_20534,N_20591);
nor U20990 (N_20990,N_20419,N_20542);
or U20991 (N_20991,N_20448,N_20621);
nand U20992 (N_20992,N_20414,N_20601);
or U20993 (N_20993,N_20550,N_20524);
nor U20994 (N_20994,N_20506,N_20415);
nor U20995 (N_20995,N_20439,N_20444);
or U20996 (N_20996,N_20690,N_20668);
and U20997 (N_20997,N_20677,N_20434);
nor U20998 (N_20998,N_20562,N_20507);
xnor U20999 (N_20999,N_20436,N_20608);
nand U21000 (N_21000,N_20851,N_20933);
and U21001 (N_21001,N_20808,N_20870);
and U21002 (N_21002,N_20771,N_20833);
xor U21003 (N_21003,N_20999,N_20957);
xor U21004 (N_21004,N_20799,N_20845);
xnor U21005 (N_21005,N_20816,N_20832);
xor U21006 (N_21006,N_20947,N_20981);
or U21007 (N_21007,N_20891,N_20977);
xnor U21008 (N_21008,N_20922,N_20732);
xor U21009 (N_21009,N_20785,N_20759);
nand U21010 (N_21010,N_20804,N_20826);
or U21011 (N_21011,N_20730,N_20788);
and U21012 (N_21012,N_20797,N_20863);
and U21013 (N_21013,N_20745,N_20767);
or U21014 (N_21014,N_20979,N_20795);
nor U21015 (N_21015,N_20992,N_20841);
or U21016 (N_21016,N_20882,N_20945);
xor U21017 (N_21017,N_20813,N_20838);
or U21018 (N_21018,N_20938,N_20723);
nor U21019 (N_21019,N_20872,N_20777);
and U21020 (N_21020,N_20984,N_20878);
and U21021 (N_21021,N_20753,N_20954);
and U21022 (N_21022,N_20706,N_20887);
nor U21023 (N_21023,N_20839,N_20919);
nand U21024 (N_21024,N_20814,N_20748);
xnor U21025 (N_21025,N_20766,N_20873);
nor U21026 (N_21026,N_20798,N_20840);
nor U21027 (N_21027,N_20900,N_20969);
and U21028 (N_21028,N_20749,N_20881);
or U21029 (N_21029,N_20726,N_20711);
xor U21030 (N_21030,N_20800,N_20927);
nor U21031 (N_21031,N_20989,N_20725);
nand U21032 (N_21032,N_20850,N_20834);
xnor U21033 (N_21033,N_20971,N_20944);
and U21034 (N_21034,N_20751,N_20948);
xnor U21035 (N_21035,N_20964,N_20958);
nand U21036 (N_21036,N_20857,N_20915);
xor U21037 (N_21037,N_20731,N_20959);
and U21038 (N_21038,N_20994,N_20993);
or U21039 (N_21039,N_20868,N_20937);
or U21040 (N_21040,N_20862,N_20756);
nor U21041 (N_21041,N_20917,N_20936);
or U21042 (N_21042,N_20807,N_20941);
nor U21043 (N_21043,N_20859,N_20712);
and U21044 (N_21044,N_20960,N_20737);
or U21045 (N_21045,N_20794,N_20763);
xnor U21046 (N_21046,N_20988,N_20829);
and U21047 (N_21047,N_20860,N_20717);
xnor U21048 (N_21048,N_20889,N_20775);
nor U21049 (N_21049,N_20883,N_20893);
or U21050 (N_21050,N_20760,N_20789);
nand U21051 (N_21051,N_20827,N_20913);
xor U21052 (N_21052,N_20735,N_20925);
nor U21053 (N_21053,N_20768,N_20902);
or U21054 (N_21054,N_20781,N_20996);
nand U21055 (N_21055,N_20995,N_20973);
nor U21056 (N_21056,N_20783,N_20837);
and U21057 (N_21057,N_20871,N_20967);
nor U21058 (N_21058,N_20818,N_20740);
or U21059 (N_21059,N_20812,N_20793);
and U21060 (N_21060,N_20911,N_20802);
nand U21061 (N_21061,N_20907,N_20820);
or U21062 (N_21062,N_20714,N_20764);
and U21063 (N_21063,N_20782,N_20848);
or U21064 (N_21064,N_20719,N_20779);
nor U21065 (N_21065,N_20842,N_20806);
nor U21066 (N_21066,N_20910,N_20955);
and U21067 (N_21067,N_20940,N_20784);
and U21068 (N_21068,N_20817,N_20861);
xor U21069 (N_21069,N_20708,N_20985);
xor U21070 (N_21070,N_20769,N_20926);
and U21071 (N_21071,N_20978,N_20904);
nand U21072 (N_21072,N_20741,N_20884);
or U21073 (N_21073,N_20701,N_20895);
nor U21074 (N_21074,N_20931,N_20786);
xnor U21075 (N_21075,N_20844,N_20879);
and U21076 (N_21076,N_20700,N_20867);
or U21077 (N_21077,N_20787,N_20966);
or U21078 (N_21078,N_20847,N_20875);
nand U21079 (N_21079,N_20946,N_20976);
or U21080 (N_21080,N_20761,N_20953);
and U21081 (N_21081,N_20715,N_20974);
nand U21082 (N_21082,N_20803,N_20705);
nand U21083 (N_21083,N_20923,N_20928);
xnor U21084 (N_21084,N_20830,N_20930);
nand U21085 (N_21085,N_20890,N_20934);
nor U21086 (N_21086,N_20924,N_20939);
nand U21087 (N_21087,N_20811,N_20831);
xor U21088 (N_21088,N_20752,N_20754);
nand U21089 (N_21089,N_20724,N_20770);
and U21090 (N_21090,N_20986,N_20908);
or U21091 (N_21091,N_20773,N_20886);
xor U21092 (N_21092,N_20744,N_20949);
nand U21093 (N_21093,N_20774,N_20702);
or U21094 (N_21094,N_20896,N_20869);
nand U21095 (N_21095,N_20997,N_20982);
xnor U21096 (N_21096,N_20963,N_20746);
nand U21097 (N_21097,N_20961,N_20972);
xor U21098 (N_21098,N_20821,N_20728);
nor U21099 (N_21099,N_20738,N_20823);
and U21100 (N_21100,N_20858,N_20901);
and U21101 (N_21101,N_20885,N_20776);
xor U21102 (N_21102,N_20899,N_20935);
and U21103 (N_21103,N_20864,N_20758);
nor U21104 (N_21104,N_20718,N_20765);
or U21105 (N_21105,N_20897,N_20734);
xnor U21106 (N_21106,N_20877,N_20778);
nor U21107 (N_21107,N_20918,N_20727);
nand U21108 (N_21108,N_20750,N_20865);
and U21109 (N_21109,N_20920,N_20796);
nor U21110 (N_21110,N_20849,N_20757);
and U21111 (N_21111,N_20942,N_20828);
or U21112 (N_21112,N_20822,N_20853);
or U21113 (N_21113,N_20888,N_20790);
or U21114 (N_21114,N_20916,N_20835);
or U21115 (N_21115,N_20780,N_20703);
and U21116 (N_21116,N_20836,N_20716);
xnor U21117 (N_21117,N_20952,N_20713);
nor U21118 (N_21118,N_20747,N_20854);
nor U21119 (N_21119,N_20709,N_20707);
and U21120 (N_21120,N_20710,N_20729);
or U21121 (N_21121,N_20965,N_20892);
and U21122 (N_21122,N_20968,N_20898);
and U21123 (N_21123,N_20991,N_20912);
nand U21124 (N_21124,N_20903,N_20739);
xnor U21125 (N_21125,N_20801,N_20733);
nor U21126 (N_21126,N_20874,N_20894);
and U21127 (N_21127,N_20943,N_20805);
nor U21128 (N_21128,N_20736,N_20855);
xor U21129 (N_21129,N_20914,N_20720);
or U21130 (N_21130,N_20909,N_20852);
nand U21131 (N_21131,N_20843,N_20792);
nor U21132 (N_21132,N_20846,N_20762);
or U21133 (N_21133,N_20866,N_20921);
nand U21134 (N_21134,N_20951,N_20983);
and U21135 (N_21135,N_20704,N_20990);
nand U21136 (N_21136,N_20950,N_20905);
or U21137 (N_21137,N_20956,N_20742);
or U21138 (N_21138,N_20856,N_20721);
nor U21139 (N_21139,N_20906,N_20743);
nor U21140 (N_21140,N_20810,N_20815);
xnor U21141 (N_21141,N_20825,N_20824);
xnor U21142 (N_21142,N_20819,N_20722);
nand U21143 (N_21143,N_20791,N_20987);
and U21144 (N_21144,N_20929,N_20876);
nand U21145 (N_21145,N_20932,N_20970);
xor U21146 (N_21146,N_20755,N_20975);
nor U21147 (N_21147,N_20980,N_20962);
nand U21148 (N_21148,N_20998,N_20880);
xor U21149 (N_21149,N_20809,N_20772);
xor U21150 (N_21150,N_20831,N_20867);
and U21151 (N_21151,N_20722,N_20766);
xnor U21152 (N_21152,N_20972,N_20963);
nor U21153 (N_21153,N_20867,N_20788);
and U21154 (N_21154,N_20762,N_20968);
nor U21155 (N_21155,N_20972,N_20870);
and U21156 (N_21156,N_20882,N_20948);
and U21157 (N_21157,N_20817,N_20828);
or U21158 (N_21158,N_20837,N_20916);
or U21159 (N_21159,N_20862,N_20740);
and U21160 (N_21160,N_20727,N_20800);
and U21161 (N_21161,N_20844,N_20980);
or U21162 (N_21162,N_20941,N_20707);
or U21163 (N_21163,N_20878,N_20723);
nor U21164 (N_21164,N_20922,N_20733);
or U21165 (N_21165,N_20803,N_20938);
xnor U21166 (N_21166,N_20789,N_20763);
and U21167 (N_21167,N_20784,N_20736);
or U21168 (N_21168,N_20991,N_20846);
xor U21169 (N_21169,N_20768,N_20709);
and U21170 (N_21170,N_20802,N_20986);
xnor U21171 (N_21171,N_20762,N_20888);
nor U21172 (N_21172,N_20806,N_20742);
and U21173 (N_21173,N_20837,N_20872);
xnor U21174 (N_21174,N_20949,N_20803);
or U21175 (N_21175,N_20784,N_20762);
xor U21176 (N_21176,N_20769,N_20972);
nand U21177 (N_21177,N_20819,N_20923);
or U21178 (N_21178,N_20989,N_20863);
xnor U21179 (N_21179,N_20792,N_20882);
nor U21180 (N_21180,N_20796,N_20801);
nand U21181 (N_21181,N_20812,N_20778);
and U21182 (N_21182,N_20846,N_20852);
or U21183 (N_21183,N_20791,N_20811);
nor U21184 (N_21184,N_20998,N_20892);
nor U21185 (N_21185,N_20962,N_20781);
or U21186 (N_21186,N_20736,N_20884);
and U21187 (N_21187,N_20845,N_20896);
xor U21188 (N_21188,N_20903,N_20995);
and U21189 (N_21189,N_20839,N_20757);
and U21190 (N_21190,N_20762,N_20836);
xor U21191 (N_21191,N_20909,N_20785);
or U21192 (N_21192,N_20947,N_20802);
nand U21193 (N_21193,N_20910,N_20877);
or U21194 (N_21194,N_20980,N_20906);
or U21195 (N_21195,N_20736,N_20728);
nand U21196 (N_21196,N_20790,N_20998);
nand U21197 (N_21197,N_20780,N_20826);
or U21198 (N_21198,N_20995,N_20820);
xnor U21199 (N_21199,N_20842,N_20702);
nor U21200 (N_21200,N_20759,N_20886);
or U21201 (N_21201,N_20731,N_20982);
xnor U21202 (N_21202,N_20818,N_20876);
and U21203 (N_21203,N_20722,N_20815);
nand U21204 (N_21204,N_20781,N_20807);
xnor U21205 (N_21205,N_20720,N_20998);
xor U21206 (N_21206,N_20941,N_20800);
nand U21207 (N_21207,N_20781,N_20748);
nand U21208 (N_21208,N_20906,N_20876);
nand U21209 (N_21209,N_20820,N_20808);
xor U21210 (N_21210,N_20789,N_20888);
or U21211 (N_21211,N_20995,N_20949);
xnor U21212 (N_21212,N_20758,N_20928);
or U21213 (N_21213,N_20975,N_20736);
or U21214 (N_21214,N_20838,N_20750);
nor U21215 (N_21215,N_20984,N_20884);
and U21216 (N_21216,N_20984,N_20776);
xor U21217 (N_21217,N_20822,N_20722);
nor U21218 (N_21218,N_20861,N_20997);
and U21219 (N_21219,N_20930,N_20881);
nand U21220 (N_21220,N_20881,N_20849);
nor U21221 (N_21221,N_20706,N_20898);
xor U21222 (N_21222,N_20979,N_20895);
nor U21223 (N_21223,N_20711,N_20878);
or U21224 (N_21224,N_20791,N_20906);
nor U21225 (N_21225,N_20929,N_20914);
xor U21226 (N_21226,N_20956,N_20923);
xor U21227 (N_21227,N_20802,N_20787);
xnor U21228 (N_21228,N_20889,N_20959);
xnor U21229 (N_21229,N_20823,N_20890);
and U21230 (N_21230,N_20712,N_20981);
or U21231 (N_21231,N_20877,N_20978);
nor U21232 (N_21232,N_20752,N_20932);
or U21233 (N_21233,N_20772,N_20994);
and U21234 (N_21234,N_20864,N_20813);
and U21235 (N_21235,N_20735,N_20879);
xor U21236 (N_21236,N_20724,N_20789);
xnor U21237 (N_21237,N_20854,N_20716);
nor U21238 (N_21238,N_20976,N_20701);
or U21239 (N_21239,N_20990,N_20894);
nor U21240 (N_21240,N_20996,N_20997);
and U21241 (N_21241,N_20738,N_20984);
or U21242 (N_21242,N_20807,N_20820);
nand U21243 (N_21243,N_20944,N_20798);
or U21244 (N_21244,N_20869,N_20993);
nor U21245 (N_21245,N_20832,N_20958);
nor U21246 (N_21246,N_20779,N_20893);
xor U21247 (N_21247,N_20874,N_20773);
nand U21248 (N_21248,N_20866,N_20802);
or U21249 (N_21249,N_20891,N_20716);
nor U21250 (N_21250,N_20924,N_20713);
nand U21251 (N_21251,N_20737,N_20966);
nand U21252 (N_21252,N_20937,N_20712);
xor U21253 (N_21253,N_20727,N_20734);
and U21254 (N_21254,N_20796,N_20849);
xor U21255 (N_21255,N_20936,N_20834);
nand U21256 (N_21256,N_20991,N_20825);
and U21257 (N_21257,N_20715,N_20773);
xnor U21258 (N_21258,N_20800,N_20744);
nand U21259 (N_21259,N_20992,N_20963);
nor U21260 (N_21260,N_20762,N_20877);
nand U21261 (N_21261,N_20903,N_20836);
nor U21262 (N_21262,N_20992,N_20955);
and U21263 (N_21263,N_20920,N_20847);
nor U21264 (N_21264,N_20834,N_20759);
and U21265 (N_21265,N_20700,N_20901);
or U21266 (N_21266,N_20741,N_20894);
nand U21267 (N_21267,N_20722,N_20973);
and U21268 (N_21268,N_20765,N_20807);
nor U21269 (N_21269,N_20985,N_20909);
or U21270 (N_21270,N_20966,N_20830);
and U21271 (N_21271,N_20974,N_20777);
nor U21272 (N_21272,N_20935,N_20873);
nor U21273 (N_21273,N_20786,N_20751);
or U21274 (N_21274,N_20827,N_20915);
xnor U21275 (N_21275,N_20926,N_20932);
and U21276 (N_21276,N_20960,N_20827);
nor U21277 (N_21277,N_20940,N_20872);
nand U21278 (N_21278,N_20741,N_20972);
nor U21279 (N_21279,N_20908,N_20738);
and U21280 (N_21280,N_20769,N_20789);
and U21281 (N_21281,N_20766,N_20831);
or U21282 (N_21282,N_20868,N_20838);
or U21283 (N_21283,N_20739,N_20797);
nand U21284 (N_21284,N_20862,N_20874);
nor U21285 (N_21285,N_20895,N_20809);
and U21286 (N_21286,N_20772,N_20719);
nand U21287 (N_21287,N_20786,N_20905);
nand U21288 (N_21288,N_20777,N_20752);
nand U21289 (N_21289,N_20814,N_20823);
or U21290 (N_21290,N_20822,N_20820);
and U21291 (N_21291,N_20909,N_20870);
nor U21292 (N_21292,N_20783,N_20720);
xor U21293 (N_21293,N_20943,N_20911);
or U21294 (N_21294,N_20746,N_20998);
nand U21295 (N_21295,N_20886,N_20813);
nor U21296 (N_21296,N_20771,N_20949);
nor U21297 (N_21297,N_20700,N_20733);
xnor U21298 (N_21298,N_20748,N_20932);
xnor U21299 (N_21299,N_20780,N_20785);
and U21300 (N_21300,N_21154,N_21226);
nand U21301 (N_21301,N_21105,N_21031);
nor U21302 (N_21302,N_21066,N_21098);
or U21303 (N_21303,N_21288,N_21016);
nand U21304 (N_21304,N_21216,N_21296);
and U21305 (N_21305,N_21179,N_21027);
nor U21306 (N_21306,N_21071,N_21019);
and U21307 (N_21307,N_21135,N_21091);
nor U21308 (N_21308,N_21205,N_21033);
and U21309 (N_21309,N_21141,N_21078);
or U21310 (N_21310,N_21262,N_21238);
xor U21311 (N_21311,N_21284,N_21011);
or U21312 (N_21312,N_21042,N_21192);
or U21313 (N_21313,N_21291,N_21024);
xor U21314 (N_21314,N_21151,N_21047);
xor U21315 (N_21315,N_21058,N_21239);
nand U21316 (N_21316,N_21074,N_21169);
nor U21317 (N_21317,N_21144,N_21265);
and U21318 (N_21318,N_21231,N_21053);
nor U21319 (N_21319,N_21089,N_21211);
xnor U21320 (N_21320,N_21229,N_21132);
or U21321 (N_21321,N_21076,N_21250);
nor U21322 (N_21322,N_21195,N_21166);
nand U21323 (N_21323,N_21234,N_21094);
and U21324 (N_21324,N_21189,N_21110);
nand U21325 (N_21325,N_21082,N_21228);
xor U21326 (N_21326,N_21181,N_21059);
and U21327 (N_21327,N_21218,N_21023);
and U21328 (N_21328,N_21186,N_21138);
xor U21329 (N_21329,N_21115,N_21057);
nand U21330 (N_21330,N_21258,N_21128);
xor U21331 (N_21331,N_21209,N_21064);
and U21332 (N_21332,N_21001,N_21259);
nor U21333 (N_21333,N_21173,N_21029);
and U21334 (N_21334,N_21095,N_21269);
nand U21335 (N_21335,N_21271,N_21097);
nand U21336 (N_21336,N_21129,N_21009);
nor U21337 (N_21337,N_21180,N_21148);
xnor U21338 (N_21338,N_21063,N_21175);
nor U21339 (N_21339,N_21039,N_21103);
and U21340 (N_21340,N_21207,N_21213);
and U21341 (N_21341,N_21206,N_21150);
nor U21342 (N_21342,N_21187,N_21010);
and U21343 (N_21343,N_21070,N_21146);
nand U21344 (N_21344,N_21235,N_21194);
and U21345 (N_21345,N_21220,N_21037);
nand U21346 (N_21346,N_21117,N_21061);
or U21347 (N_21347,N_21268,N_21287);
and U21348 (N_21348,N_21118,N_21116);
nand U21349 (N_21349,N_21253,N_21130);
or U21350 (N_21350,N_21062,N_21090);
nand U21351 (N_21351,N_21295,N_21275);
nor U21352 (N_21352,N_21190,N_21297);
nor U21353 (N_21353,N_21005,N_21018);
xor U21354 (N_21354,N_21026,N_21096);
and U21355 (N_21355,N_21045,N_21160);
xnor U21356 (N_21356,N_21188,N_21164);
xnor U21357 (N_21357,N_21281,N_21157);
or U21358 (N_21358,N_21134,N_21083);
nor U21359 (N_21359,N_21214,N_21267);
nand U21360 (N_21360,N_21067,N_21102);
or U21361 (N_21361,N_21131,N_21075);
nand U21362 (N_21362,N_21012,N_21198);
and U21363 (N_21363,N_21167,N_21208);
or U21364 (N_21364,N_21145,N_21282);
xor U21365 (N_21365,N_21123,N_21152);
xor U21366 (N_21366,N_21125,N_21252);
xnor U21367 (N_21367,N_21162,N_21200);
or U21368 (N_21368,N_21017,N_21104);
nor U21369 (N_21369,N_21000,N_21093);
and U21370 (N_21370,N_21038,N_21004);
or U21371 (N_21371,N_21034,N_21197);
and U21372 (N_21372,N_21283,N_21286);
nand U21373 (N_21373,N_21032,N_21114);
nor U21374 (N_21374,N_21112,N_21247);
xor U21375 (N_21375,N_21241,N_21086);
and U21376 (N_21376,N_21273,N_21041);
xnor U21377 (N_21377,N_21035,N_21266);
or U21378 (N_21378,N_21278,N_21165);
nand U21379 (N_21379,N_21279,N_21088);
or U21380 (N_21380,N_21227,N_21084);
xor U21381 (N_21381,N_21137,N_21025);
and U21382 (N_21382,N_21100,N_21274);
nand U21383 (N_21383,N_21108,N_21133);
nor U21384 (N_21384,N_21008,N_21264);
nand U21385 (N_21385,N_21055,N_21174);
and U21386 (N_21386,N_21002,N_21290);
xor U21387 (N_21387,N_21245,N_21219);
or U21388 (N_21388,N_21298,N_21223);
and U21389 (N_21389,N_21246,N_21178);
and U21390 (N_21390,N_21243,N_21201);
nand U21391 (N_21391,N_21212,N_21251);
and U21392 (N_21392,N_21242,N_21050);
nand U21393 (N_21393,N_21109,N_21196);
or U21394 (N_21394,N_21036,N_21003);
xnor U21395 (N_21395,N_21254,N_21299);
nand U21396 (N_21396,N_21046,N_21065);
xnor U21397 (N_21397,N_21040,N_21007);
or U21398 (N_21398,N_21049,N_21043);
xor U21399 (N_21399,N_21289,N_21263);
and U21400 (N_21400,N_21244,N_21225);
or U21401 (N_21401,N_21028,N_21052);
nor U21402 (N_21402,N_21260,N_21221);
xnor U21403 (N_21403,N_21156,N_21230);
or U21404 (N_21404,N_21185,N_21294);
or U21405 (N_21405,N_21124,N_21222);
and U21406 (N_21406,N_21120,N_21060);
nor U21407 (N_21407,N_21199,N_21277);
xor U21408 (N_21408,N_21248,N_21056);
and U21409 (N_21409,N_21073,N_21285);
and U21410 (N_21410,N_21210,N_21163);
and U21411 (N_21411,N_21111,N_21072);
nand U21412 (N_21412,N_21183,N_21155);
xor U21413 (N_21413,N_21147,N_21069);
and U21414 (N_21414,N_21153,N_21126);
or U21415 (N_21415,N_21237,N_21044);
or U21416 (N_21416,N_21292,N_21014);
xor U21417 (N_21417,N_21092,N_21079);
nand U21418 (N_21418,N_21006,N_21232);
xnor U21419 (N_21419,N_21113,N_21149);
nand U21420 (N_21420,N_21280,N_21215);
and U21421 (N_21421,N_21139,N_21101);
and U21422 (N_21422,N_21158,N_21077);
nand U21423 (N_21423,N_21081,N_21127);
nand U21424 (N_21424,N_21020,N_21172);
or U21425 (N_21425,N_21143,N_21256);
or U21426 (N_21426,N_21048,N_21236);
or U21427 (N_21427,N_21119,N_21270);
and U21428 (N_21428,N_21217,N_21184);
nand U21429 (N_21429,N_21272,N_21257);
nand U21430 (N_21430,N_21099,N_21171);
nand U21431 (N_21431,N_21168,N_21054);
and U21432 (N_21432,N_21191,N_21177);
nor U21433 (N_21433,N_21170,N_21015);
or U21434 (N_21434,N_21085,N_21107);
nand U21435 (N_21435,N_21261,N_21249);
or U21436 (N_21436,N_21051,N_21022);
xor U21437 (N_21437,N_21142,N_21240);
nor U21438 (N_21438,N_21021,N_21140);
nand U21439 (N_21439,N_21122,N_21013);
nor U21440 (N_21440,N_21202,N_21106);
nand U21441 (N_21441,N_21193,N_21182);
and U21442 (N_21442,N_21224,N_21276);
and U21443 (N_21443,N_21121,N_21136);
nor U21444 (N_21444,N_21068,N_21233);
nor U21445 (N_21445,N_21204,N_21255);
and U21446 (N_21446,N_21087,N_21159);
nor U21447 (N_21447,N_21293,N_21080);
and U21448 (N_21448,N_21176,N_21030);
and U21449 (N_21449,N_21203,N_21161);
nand U21450 (N_21450,N_21192,N_21203);
nand U21451 (N_21451,N_21269,N_21092);
nand U21452 (N_21452,N_21090,N_21237);
nand U21453 (N_21453,N_21015,N_21100);
or U21454 (N_21454,N_21019,N_21130);
or U21455 (N_21455,N_21006,N_21157);
nor U21456 (N_21456,N_21243,N_21239);
xor U21457 (N_21457,N_21155,N_21238);
xor U21458 (N_21458,N_21040,N_21244);
or U21459 (N_21459,N_21073,N_21264);
xor U21460 (N_21460,N_21097,N_21185);
or U21461 (N_21461,N_21037,N_21072);
nor U21462 (N_21462,N_21182,N_21196);
nand U21463 (N_21463,N_21066,N_21076);
xnor U21464 (N_21464,N_21208,N_21040);
xnor U21465 (N_21465,N_21168,N_21291);
nor U21466 (N_21466,N_21009,N_21130);
nand U21467 (N_21467,N_21054,N_21209);
xor U21468 (N_21468,N_21201,N_21143);
nand U21469 (N_21469,N_21142,N_21182);
and U21470 (N_21470,N_21091,N_21025);
nor U21471 (N_21471,N_21221,N_21071);
nand U21472 (N_21472,N_21147,N_21016);
xnor U21473 (N_21473,N_21166,N_21032);
or U21474 (N_21474,N_21263,N_21083);
and U21475 (N_21475,N_21252,N_21064);
nand U21476 (N_21476,N_21202,N_21294);
and U21477 (N_21477,N_21096,N_21179);
xnor U21478 (N_21478,N_21267,N_21188);
xor U21479 (N_21479,N_21007,N_21080);
or U21480 (N_21480,N_21049,N_21205);
nand U21481 (N_21481,N_21266,N_21218);
nand U21482 (N_21482,N_21044,N_21151);
and U21483 (N_21483,N_21238,N_21221);
nor U21484 (N_21484,N_21143,N_21285);
or U21485 (N_21485,N_21213,N_21010);
and U21486 (N_21486,N_21179,N_21086);
and U21487 (N_21487,N_21238,N_21188);
or U21488 (N_21488,N_21027,N_21068);
nor U21489 (N_21489,N_21085,N_21290);
xor U21490 (N_21490,N_21218,N_21128);
xor U21491 (N_21491,N_21228,N_21017);
or U21492 (N_21492,N_21253,N_21044);
xor U21493 (N_21493,N_21101,N_21124);
and U21494 (N_21494,N_21124,N_21023);
xor U21495 (N_21495,N_21130,N_21170);
or U21496 (N_21496,N_21235,N_21085);
xor U21497 (N_21497,N_21087,N_21221);
nand U21498 (N_21498,N_21114,N_21119);
nand U21499 (N_21499,N_21183,N_21255);
xnor U21500 (N_21500,N_21151,N_21150);
nand U21501 (N_21501,N_21225,N_21235);
or U21502 (N_21502,N_21039,N_21206);
and U21503 (N_21503,N_21080,N_21075);
nand U21504 (N_21504,N_21041,N_21164);
xnor U21505 (N_21505,N_21110,N_21221);
xor U21506 (N_21506,N_21061,N_21029);
nor U21507 (N_21507,N_21110,N_21244);
xor U21508 (N_21508,N_21271,N_21174);
or U21509 (N_21509,N_21231,N_21171);
or U21510 (N_21510,N_21187,N_21101);
nor U21511 (N_21511,N_21001,N_21083);
and U21512 (N_21512,N_21196,N_21261);
xnor U21513 (N_21513,N_21046,N_21276);
nand U21514 (N_21514,N_21144,N_21058);
or U21515 (N_21515,N_21245,N_21161);
xnor U21516 (N_21516,N_21107,N_21168);
nand U21517 (N_21517,N_21107,N_21263);
or U21518 (N_21518,N_21186,N_21233);
xor U21519 (N_21519,N_21145,N_21284);
and U21520 (N_21520,N_21217,N_21182);
or U21521 (N_21521,N_21074,N_21265);
nor U21522 (N_21522,N_21113,N_21129);
and U21523 (N_21523,N_21288,N_21049);
nand U21524 (N_21524,N_21176,N_21129);
nor U21525 (N_21525,N_21111,N_21149);
nor U21526 (N_21526,N_21055,N_21054);
nor U21527 (N_21527,N_21157,N_21231);
nor U21528 (N_21528,N_21265,N_21193);
xor U21529 (N_21529,N_21225,N_21063);
or U21530 (N_21530,N_21103,N_21031);
or U21531 (N_21531,N_21076,N_21117);
nand U21532 (N_21532,N_21201,N_21133);
nand U21533 (N_21533,N_21102,N_21226);
or U21534 (N_21534,N_21070,N_21245);
or U21535 (N_21535,N_21145,N_21287);
nand U21536 (N_21536,N_21215,N_21060);
nor U21537 (N_21537,N_21031,N_21195);
nor U21538 (N_21538,N_21000,N_21259);
nor U21539 (N_21539,N_21268,N_21157);
nor U21540 (N_21540,N_21224,N_21263);
nor U21541 (N_21541,N_21071,N_21002);
xnor U21542 (N_21542,N_21199,N_21015);
nand U21543 (N_21543,N_21178,N_21140);
xnor U21544 (N_21544,N_21035,N_21211);
xnor U21545 (N_21545,N_21157,N_21192);
or U21546 (N_21546,N_21174,N_21159);
and U21547 (N_21547,N_21008,N_21035);
nor U21548 (N_21548,N_21251,N_21241);
nand U21549 (N_21549,N_21044,N_21004);
and U21550 (N_21550,N_21241,N_21122);
and U21551 (N_21551,N_21023,N_21264);
xor U21552 (N_21552,N_21278,N_21233);
nand U21553 (N_21553,N_21109,N_21076);
nor U21554 (N_21554,N_21135,N_21009);
xor U21555 (N_21555,N_21079,N_21272);
or U21556 (N_21556,N_21208,N_21235);
nor U21557 (N_21557,N_21019,N_21252);
xor U21558 (N_21558,N_21047,N_21189);
or U21559 (N_21559,N_21245,N_21281);
nand U21560 (N_21560,N_21246,N_21297);
nand U21561 (N_21561,N_21088,N_21079);
nand U21562 (N_21562,N_21118,N_21260);
nor U21563 (N_21563,N_21035,N_21131);
nand U21564 (N_21564,N_21131,N_21211);
xor U21565 (N_21565,N_21176,N_21175);
nand U21566 (N_21566,N_21042,N_21187);
and U21567 (N_21567,N_21053,N_21012);
xnor U21568 (N_21568,N_21258,N_21107);
or U21569 (N_21569,N_21052,N_21017);
nor U21570 (N_21570,N_21274,N_21087);
nor U21571 (N_21571,N_21087,N_21239);
nand U21572 (N_21572,N_21092,N_21031);
xnor U21573 (N_21573,N_21292,N_21205);
and U21574 (N_21574,N_21044,N_21145);
xnor U21575 (N_21575,N_21112,N_21208);
and U21576 (N_21576,N_21262,N_21260);
nor U21577 (N_21577,N_21000,N_21257);
nor U21578 (N_21578,N_21262,N_21226);
nand U21579 (N_21579,N_21117,N_21251);
or U21580 (N_21580,N_21034,N_21168);
xnor U21581 (N_21581,N_21295,N_21039);
and U21582 (N_21582,N_21293,N_21060);
nand U21583 (N_21583,N_21197,N_21132);
and U21584 (N_21584,N_21015,N_21120);
or U21585 (N_21585,N_21067,N_21047);
nand U21586 (N_21586,N_21122,N_21158);
and U21587 (N_21587,N_21286,N_21082);
or U21588 (N_21588,N_21200,N_21286);
nor U21589 (N_21589,N_21127,N_21193);
or U21590 (N_21590,N_21110,N_21297);
xor U21591 (N_21591,N_21151,N_21020);
nor U21592 (N_21592,N_21184,N_21135);
xnor U21593 (N_21593,N_21070,N_21006);
nand U21594 (N_21594,N_21096,N_21222);
nand U21595 (N_21595,N_21270,N_21268);
or U21596 (N_21596,N_21155,N_21172);
or U21597 (N_21597,N_21234,N_21210);
xor U21598 (N_21598,N_21150,N_21228);
and U21599 (N_21599,N_21028,N_21039);
nand U21600 (N_21600,N_21413,N_21448);
nor U21601 (N_21601,N_21542,N_21355);
nand U21602 (N_21602,N_21533,N_21528);
nor U21603 (N_21603,N_21302,N_21536);
xor U21604 (N_21604,N_21568,N_21336);
and U21605 (N_21605,N_21304,N_21566);
nand U21606 (N_21606,N_21353,N_21541);
nor U21607 (N_21607,N_21396,N_21330);
and U21608 (N_21608,N_21492,N_21548);
nor U21609 (N_21609,N_21476,N_21424);
and U21610 (N_21610,N_21497,N_21598);
xnor U21611 (N_21611,N_21459,N_21391);
and U21612 (N_21612,N_21559,N_21378);
xnor U21613 (N_21613,N_21417,N_21442);
or U21614 (N_21614,N_21576,N_21452);
xnor U21615 (N_21615,N_21578,N_21407);
nor U21616 (N_21616,N_21467,N_21496);
xnor U21617 (N_21617,N_21303,N_21591);
or U21618 (N_21618,N_21432,N_21325);
nand U21619 (N_21619,N_21509,N_21431);
nor U21620 (N_21620,N_21483,N_21338);
nor U21621 (N_21621,N_21398,N_21488);
or U21622 (N_21622,N_21331,N_21594);
or U21623 (N_21623,N_21346,N_21505);
nand U21624 (N_21624,N_21446,N_21337);
nand U21625 (N_21625,N_21320,N_21478);
xnor U21626 (N_21626,N_21361,N_21557);
xor U21627 (N_21627,N_21412,N_21313);
nand U21628 (N_21628,N_21362,N_21474);
and U21629 (N_21629,N_21575,N_21414);
nor U21630 (N_21630,N_21455,N_21597);
nor U21631 (N_21631,N_21399,N_21363);
or U21632 (N_21632,N_21444,N_21360);
nor U21633 (N_21633,N_21377,N_21502);
xnor U21634 (N_21634,N_21365,N_21599);
and U21635 (N_21635,N_21486,N_21352);
or U21636 (N_21636,N_21401,N_21529);
nor U21637 (N_21637,N_21511,N_21480);
xor U21638 (N_21638,N_21309,N_21384);
xor U21639 (N_21639,N_21383,N_21418);
xor U21640 (N_21640,N_21435,N_21580);
nor U21641 (N_21641,N_21489,N_21461);
or U21642 (N_21642,N_21341,N_21411);
xnor U21643 (N_21643,N_21322,N_21425);
or U21644 (N_21644,N_21538,N_21439);
or U21645 (N_21645,N_21312,N_21386);
and U21646 (N_21646,N_21571,N_21403);
and U21647 (N_21647,N_21438,N_21427);
nor U21648 (N_21648,N_21589,N_21545);
and U21649 (N_21649,N_21395,N_21404);
nand U21650 (N_21650,N_21370,N_21582);
nor U21651 (N_21651,N_21437,N_21326);
nor U21652 (N_21652,N_21526,N_21596);
xnor U21653 (N_21653,N_21408,N_21344);
or U21654 (N_21654,N_21410,N_21453);
and U21655 (N_21655,N_21462,N_21584);
and U21656 (N_21656,N_21433,N_21556);
nor U21657 (N_21657,N_21560,N_21314);
or U21658 (N_21658,N_21562,N_21315);
or U21659 (N_21659,N_21416,N_21306);
nor U21660 (N_21660,N_21570,N_21481);
nand U21661 (N_21661,N_21328,N_21555);
nor U21662 (N_21662,N_21521,N_21321);
nand U21663 (N_21663,N_21310,N_21517);
nand U21664 (N_21664,N_21450,N_21350);
nor U21665 (N_21665,N_21436,N_21340);
and U21666 (N_21666,N_21558,N_21587);
xnor U21667 (N_21667,N_21379,N_21335);
or U21668 (N_21668,N_21593,N_21485);
nor U21669 (N_21669,N_21394,N_21451);
xnor U21670 (N_21670,N_21458,N_21371);
nand U21671 (N_21671,N_21549,N_21380);
xnor U21672 (N_21672,N_21588,N_21323);
nand U21673 (N_21673,N_21551,N_21531);
nand U21674 (N_21674,N_21347,N_21527);
xnor U21675 (N_21675,N_21504,N_21506);
xnor U21676 (N_21676,N_21577,N_21369);
or U21677 (N_21677,N_21372,N_21420);
or U21678 (N_21678,N_21457,N_21507);
and U21679 (N_21679,N_21547,N_21388);
and U21680 (N_21680,N_21333,N_21554);
xor U21681 (N_21681,N_21469,N_21465);
and U21682 (N_21682,N_21464,N_21585);
xnor U21683 (N_21683,N_21454,N_21499);
and U21684 (N_21684,N_21430,N_21510);
and U21685 (N_21685,N_21482,N_21405);
and U21686 (N_21686,N_21423,N_21519);
xor U21687 (N_21687,N_21543,N_21429);
nor U21688 (N_21688,N_21441,N_21351);
xor U21689 (N_21689,N_21463,N_21493);
nor U21690 (N_21690,N_21305,N_21339);
or U21691 (N_21691,N_21516,N_21477);
nor U21692 (N_21692,N_21409,N_21348);
or U21693 (N_21693,N_21532,N_21534);
nor U21694 (N_21694,N_21358,N_21422);
xor U21695 (N_21695,N_21475,N_21523);
xnor U21696 (N_21696,N_21544,N_21579);
or U21697 (N_21697,N_21392,N_21468);
nand U21698 (N_21698,N_21592,N_21581);
or U21699 (N_21699,N_21316,N_21434);
nand U21700 (N_21700,N_21513,N_21368);
nand U21701 (N_21701,N_21397,N_21373);
nor U21702 (N_21702,N_21546,N_21428);
nand U21703 (N_21703,N_21415,N_21334);
xnor U21704 (N_21704,N_21550,N_21300);
xor U21705 (N_21705,N_21484,N_21381);
xor U21706 (N_21706,N_21524,N_21382);
xor U21707 (N_21707,N_21318,N_21374);
xor U21708 (N_21708,N_21552,N_21518);
and U21709 (N_21709,N_21343,N_21494);
nand U21710 (N_21710,N_21466,N_21421);
and U21711 (N_21711,N_21332,N_21574);
nor U21712 (N_21712,N_21500,N_21456);
and U21713 (N_21713,N_21349,N_21573);
and U21714 (N_21714,N_21449,N_21586);
nand U21715 (N_21715,N_21402,N_21512);
and U21716 (N_21716,N_21530,N_21356);
xor U21717 (N_21717,N_21359,N_21515);
or U21718 (N_21718,N_21501,N_21387);
nand U21719 (N_21719,N_21307,N_21471);
nand U21720 (N_21720,N_21525,N_21445);
or U21721 (N_21721,N_21508,N_21367);
or U21722 (N_21722,N_21472,N_21522);
or U21723 (N_21723,N_21537,N_21572);
nor U21724 (N_21724,N_21389,N_21495);
nand U21725 (N_21725,N_21440,N_21590);
and U21726 (N_21726,N_21375,N_21479);
nor U21727 (N_21727,N_21470,N_21535);
xor U21728 (N_21728,N_21406,N_21491);
nor U21729 (N_21729,N_21390,N_21498);
and U21730 (N_21730,N_21364,N_21376);
nor U21731 (N_21731,N_21443,N_21385);
xnor U21732 (N_21732,N_21393,N_21327);
and U21733 (N_21733,N_21311,N_21460);
nand U21734 (N_21734,N_21564,N_21319);
and U21735 (N_21735,N_21563,N_21565);
nor U21736 (N_21736,N_21317,N_21487);
and U21737 (N_21737,N_21324,N_21400);
xor U21738 (N_21738,N_21354,N_21419);
xor U21739 (N_21739,N_21345,N_21569);
nor U21740 (N_21740,N_21357,N_21342);
and U21741 (N_21741,N_21426,N_21540);
nand U21742 (N_21742,N_21514,N_21561);
nand U21743 (N_21743,N_21473,N_21520);
and U21744 (N_21744,N_21366,N_21503);
and U21745 (N_21745,N_21539,N_21490);
or U21746 (N_21746,N_21553,N_21567);
xnor U21747 (N_21747,N_21447,N_21301);
xnor U21748 (N_21748,N_21595,N_21583);
or U21749 (N_21749,N_21329,N_21308);
or U21750 (N_21750,N_21593,N_21374);
or U21751 (N_21751,N_21596,N_21331);
xor U21752 (N_21752,N_21309,N_21402);
or U21753 (N_21753,N_21538,N_21526);
xnor U21754 (N_21754,N_21562,N_21571);
xor U21755 (N_21755,N_21418,N_21497);
or U21756 (N_21756,N_21438,N_21476);
and U21757 (N_21757,N_21434,N_21545);
xnor U21758 (N_21758,N_21410,N_21387);
nor U21759 (N_21759,N_21599,N_21534);
nor U21760 (N_21760,N_21437,N_21584);
nor U21761 (N_21761,N_21536,N_21347);
and U21762 (N_21762,N_21338,N_21599);
or U21763 (N_21763,N_21471,N_21351);
xnor U21764 (N_21764,N_21350,N_21455);
nor U21765 (N_21765,N_21480,N_21389);
or U21766 (N_21766,N_21402,N_21409);
and U21767 (N_21767,N_21585,N_21353);
nand U21768 (N_21768,N_21433,N_21419);
nor U21769 (N_21769,N_21337,N_21300);
xnor U21770 (N_21770,N_21314,N_21587);
nand U21771 (N_21771,N_21307,N_21391);
and U21772 (N_21772,N_21327,N_21328);
or U21773 (N_21773,N_21372,N_21395);
nand U21774 (N_21774,N_21489,N_21587);
xnor U21775 (N_21775,N_21556,N_21336);
xor U21776 (N_21776,N_21471,N_21599);
nor U21777 (N_21777,N_21441,N_21377);
nor U21778 (N_21778,N_21556,N_21321);
nor U21779 (N_21779,N_21347,N_21314);
xor U21780 (N_21780,N_21511,N_21452);
xor U21781 (N_21781,N_21357,N_21458);
nand U21782 (N_21782,N_21514,N_21357);
and U21783 (N_21783,N_21547,N_21554);
nand U21784 (N_21784,N_21364,N_21475);
xor U21785 (N_21785,N_21493,N_21395);
or U21786 (N_21786,N_21467,N_21570);
nand U21787 (N_21787,N_21554,N_21431);
nor U21788 (N_21788,N_21450,N_21591);
and U21789 (N_21789,N_21503,N_21301);
nor U21790 (N_21790,N_21331,N_21383);
or U21791 (N_21791,N_21347,N_21498);
xor U21792 (N_21792,N_21548,N_21416);
or U21793 (N_21793,N_21504,N_21576);
nor U21794 (N_21794,N_21365,N_21460);
xor U21795 (N_21795,N_21371,N_21585);
nor U21796 (N_21796,N_21569,N_21332);
nand U21797 (N_21797,N_21497,N_21540);
nor U21798 (N_21798,N_21575,N_21409);
or U21799 (N_21799,N_21402,N_21324);
and U21800 (N_21800,N_21471,N_21404);
nand U21801 (N_21801,N_21391,N_21343);
and U21802 (N_21802,N_21420,N_21502);
xnor U21803 (N_21803,N_21590,N_21317);
or U21804 (N_21804,N_21322,N_21386);
and U21805 (N_21805,N_21495,N_21316);
nand U21806 (N_21806,N_21556,N_21499);
xor U21807 (N_21807,N_21422,N_21597);
and U21808 (N_21808,N_21427,N_21519);
and U21809 (N_21809,N_21342,N_21460);
or U21810 (N_21810,N_21509,N_21391);
xnor U21811 (N_21811,N_21360,N_21513);
nand U21812 (N_21812,N_21510,N_21501);
nand U21813 (N_21813,N_21340,N_21528);
xor U21814 (N_21814,N_21477,N_21568);
nor U21815 (N_21815,N_21459,N_21525);
xnor U21816 (N_21816,N_21386,N_21367);
and U21817 (N_21817,N_21419,N_21445);
nor U21818 (N_21818,N_21329,N_21417);
or U21819 (N_21819,N_21495,N_21377);
or U21820 (N_21820,N_21302,N_21423);
nor U21821 (N_21821,N_21546,N_21389);
and U21822 (N_21822,N_21318,N_21414);
xor U21823 (N_21823,N_21409,N_21437);
xor U21824 (N_21824,N_21423,N_21533);
nor U21825 (N_21825,N_21426,N_21433);
nor U21826 (N_21826,N_21574,N_21360);
nor U21827 (N_21827,N_21436,N_21433);
and U21828 (N_21828,N_21397,N_21552);
nand U21829 (N_21829,N_21473,N_21551);
and U21830 (N_21830,N_21473,N_21352);
and U21831 (N_21831,N_21350,N_21403);
or U21832 (N_21832,N_21357,N_21494);
or U21833 (N_21833,N_21308,N_21540);
nand U21834 (N_21834,N_21541,N_21302);
or U21835 (N_21835,N_21392,N_21472);
nand U21836 (N_21836,N_21399,N_21589);
and U21837 (N_21837,N_21392,N_21359);
xnor U21838 (N_21838,N_21310,N_21537);
and U21839 (N_21839,N_21380,N_21485);
and U21840 (N_21840,N_21494,N_21487);
nand U21841 (N_21841,N_21512,N_21580);
and U21842 (N_21842,N_21506,N_21342);
nor U21843 (N_21843,N_21508,N_21312);
nand U21844 (N_21844,N_21520,N_21551);
xnor U21845 (N_21845,N_21364,N_21451);
or U21846 (N_21846,N_21319,N_21395);
nand U21847 (N_21847,N_21426,N_21533);
xor U21848 (N_21848,N_21439,N_21337);
or U21849 (N_21849,N_21455,N_21335);
or U21850 (N_21850,N_21419,N_21535);
nor U21851 (N_21851,N_21331,N_21314);
nor U21852 (N_21852,N_21562,N_21444);
nand U21853 (N_21853,N_21443,N_21463);
xnor U21854 (N_21854,N_21427,N_21588);
xnor U21855 (N_21855,N_21389,N_21517);
nand U21856 (N_21856,N_21456,N_21447);
and U21857 (N_21857,N_21319,N_21313);
xor U21858 (N_21858,N_21369,N_21560);
xor U21859 (N_21859,N_21312,N_21422);
xor U21860 (N_21860,N_21321,N_21429);
or U21861 (N_21861,N_21353,N_21402);
nor U21862 (N_21862,N_21357,N_21543);
xnor U21863 (N_21863,N_21490,N_21378);
or U21864 (N_21864,N_21596,N_21407);
xnor U21865 (N_21865,N_21456,N_21377);
nand U21866 (N_21866,N_21407,N_21562);
or U21867 (N_21867,N_21462,N_21320);
or U21868 (N_21868,N_21352,N_21418);
nand U21869 (N_21869,N_21366,N_21364);
or U21870 (N_21870,N_21304,N_21344);
nor U21871 (N_21871,N_21433,N_21348);
and U21872 (N_21872,N_21404,N_21422);
nand U21873 (N_21873,N_21548,N_21343);
and U21874 (N_21874,N_21431,N_21396);
nand U21875 (N_21875,N_21349,N_21501);
or U21876 (N_21876,N_21356,N_21340);
or U21877 (N_21877,N_21557,N_21553);
nor U21878 (N_21878,N_21303,N_21467);
xor U21879 (N_21879,N_21504,N_21456);
or U21880 (N_21880,N_21378,N_21563);
xnor U21881 (N_21881,N_21509,N_21401);
nand U21882 (N_21882,N_21533,N_21501);
nor U21883 (N_21883,N_21596,N_21519);
nand U21884 (N_21884,N_21405,N_21490);
nand U21885 (N_21885,N_21455,N_21438);
and U21886 (N_21886,N_21455,N_21531);
or U21887 (N_21887,N_21446,N_21564);
nand U21888 (N_21888,N_21304,N_21461);
xor U21889 (N_21889,N_21512,N_21363);
or U21890 (N_21890,N_21524,N_21351);
nor U21891 (N_21891,N_21506,N_21519);
xor U21892 (N_21892,N_21594,N_21301);
xor U21893 (N_21893,N_21495,N_21373);
xor U21894 (N_21894,N_21461,N_21513);
or U21895 (N_21895,N_21537,N_21575);
nand U21896 (N_21896,N_21358,N_21369);
nand U21897 (N_21897,N_21578,N_21436);
xor U21898 (N_21898,N_21453,N_21342);
and U21899 (N_21899,N_21453,N_21463);
nor U21900 (N_21900,N_21877,N_21687);
nand U21901 (N_21901,N_21754,N_21624);
xnor U21902 (N_21902,N_21628,N_21758);
nor U21903 (N_21903,N_21619,N_21642);
nand U21904 (N_21904,N_21644,N_21615);
xnor U21905 (N_21905,N_21785,N_21647);
nor U21906 (N_21906,N_21717,N_21856);
nand U21907 (N_21907,N_21636,N_21750);
or U21908 (N_21908,N_21838,N_21732);
nor U21909 (N_21909,N_21871,N_21844);
and U21910 (N_21910,N_21777,N_21834);
and U21911 (N_21911,N_21799,N_21783);
xor U21912 (N_21912,N_21688,N_21842);
nand U21913 (N_21913,N_21665,N_21709);
xnor U21914 (N_21914,N_21755,N_21780);
xnor U21915 (N_21915,N_21649,N_21814);
and U21916 (N_21916,N_21663,N_21859);
or U21917 (N_21917,N_21802,N_21801);
or U21918 (N_21918,N_21828,N_21762);
nand U21919 (N_21919,N_21708,N_21811);
nand U21920 (N_21920,N_21635,N_21696);
nor U21921 (N_21921,N_21741,N_21793);
and U21922 (N_21922,N_21872,N_21770);
and U21923 (N_21923,N_21684,N_21716);
or U21924 (N_21924,N_21723,N_21671);
xnor U21925 (N_21925,N_21623,N_21662);
nand U21926 (N_21926,N_21724,N_21705);
or U21927 (N_21927,N_21867,N_21721);
xor U21928 (N_21928,N_21894,N_21769);
or U21929 (N_21929,N_21712,N_21673);
xor U21930 (N_21930,N_21809,N_21704);
xnor U21931 (N_21931,N_21786,N_21690);
nor U21932 (N_21932,N_21808,N_21691);
and U21933 (N_21933,N_21610,N_21693);
nand U21934 (N_21934,N_21831,N_21845);
xnor U21935 (N_21935,N_21676,N_21703);
nand U21936 (N_21936,N_21600,N_21745);
nand U21937 (N_21937,N_21678,N_21638);
xor U21938 (N_21938,N_21620,N_21836);
nor U21939 (N_21939,N_21847,N_21820);
or U21940 (N_21940,N_21781,N_21746);
nand U21941 (N_21941,N_21878,N_21775);
nor U21942 (N_21942,N_21860,N_21810);
nand U21943 (N_21943,N_21829,N_21759);
nor U21944 (N_21944,N_21627,N_21764);
or U21945 (N_21945,N_21695,N_21824);
xor U21946 (N_21946,N_21700,N_21886);
and U21947 (N_21947,N_21631,N_21885);
nor U21948 (N_21948,N_21617,N_21800);
and U21949 (N_21949,N_21643,N_21841);
xnor U21950 (N_21950,N_21735,N_21849);
nor U21951 (N_21951,N_21794,N_21651);
or U21952 (N_21952,N_21817,N_21654);
or U21953 (N_21953,N_21887,N_21603);
nor U21954 (N_21954,N_21602,N_21726);
and U21955 (N_21955,N_21792,N_21822);
and U21956 (N_21956,N_21702,N_21641);
or U21957 (N_21957,N_21694,N_21893);
nand U21958 (N_21958,N_21748,N_21753);
nor U21959 (N_21959,N_21664,N_21659);
or U21960 (N_21960,N_21742,N_21682);
xor U21961 (N_21961,N_21632,N_21895);
nand U21962 (N_21962,N_21701,N_21614);
nor U21963 (N_21963,N_21813,N_21760);
nor U21964 (N_21964,N_21692,N_21655);
and U21965 (N_21965,N_21848,N_21681);
nor U21966 (N_21966,N_21736,N_21622);
and U21967 (N_21967,N_21774,N_21605);
xor U21968 (N_21968,N_21881,N_21850);
xnor U21969 (N_21969,N_21680,N_21621);
or U21970 (N_21970,N_21675,N_21660);
nor U21971 (N_21971,N_21714,N_21639);
xor U21972 (N_21972,N_21719,N_21720);
nor U21973 (N_21973,N_21821,N_21648);
nand U21974 (N_21974,N_21843,N_21883);
nand U21975 (N_21975,N_21803,N_21782);
nand U21976 (N_21976,N_21618,N_21728);
nor U21977 (N_21977,N_21747,N_21870);
or U21978 (N_21978,N_21854,N_21862);
nor U21979 (N_21979,N_21882,N_21778);
nor U21980 (N_21980,N_21707,N_21879);
nand U21981 (N_21981,N_21890,N_21827);
nor U21982 (N_21982,N_21761,N_21865);
or U21983 (N_21983,N_21667,N_21805);
nor U21984 (N_21984,N_21731,N_21697);
nor U21985 (N_21985,N_21787,N_21630);
nor U21986 (N_21986,N_21689,N_21674);
xor U21987 (N_21987,N_21738,N_21767);
or U21988 (N_21988,N_21670,N_21823);
or U21989 (N_21989,N_21613,N_21896);
xor U21990 (N_21990,N_21863,N_21768);
xor U21991 (N_21991,N_21668,N_21725);
and U21992 (N_21992,N_21771,N_21650);
or U21993 (N_21993,N_21866,N_21818);
nor U21994 (N_21994,N_21629,N_21729);
or U21995 (N_21995,N_21727,N_21686);
or U21996 (N_21996,N_21640,N_21825);
and U21997 (N_21997,N_21855,N_21601);
nor U21998 (N_21998,N_21606,N_21791);
nand U21999 (N_21999,N_21772,N_21740);
nand U22000 (N_22000,N_21661,N_21652);
xnor U22001 (N_22001,N_21840,N_21857);
xor U22002 (N_22002,N_21889,N_21698);
xor U22003 (N_22003,N_21752,N_21611);
xor U22004 (N_22004,N_21658,N_21830);
nor U22005 (N_22005,N_21898,N_21853);
xnor U22006 (N_22006,N_21864,N_21733);
xnor U22007 (N_22007,N_21710,N_21739);
nor U22008 (N_22008,N_21626,N_21796);
and U22009 (N_22009,N_21656,N_21888);
and U22010 (N_22010,N_21784,N_21608);
or U22011 (N_22011,N_21730,N_21633);
nand U22012 (N_22012,N_21645,N_21666);
or U22013 (N_22013,N_21788,N_21763);
or U22014 (N_22014,N_21625,N_21815);
nand U22015 (N_22015,N_21826,N_21756);
xor U22016 (N_22016,N_21646,N_21892);
nor U22017 (N_22017,N_21743,N_21837);
and U22018 (N_22018,N_21711,N_21779);
or U22019 (N_22019,N_21683,N_21832);
nand U22020 (N_22020,N_21806,N_21751);
or U22021 (N_22021,N_21819,N_21873);
and U22022 (N_22022,N_21765,N_21861);
nor U22023 (N_22023,N_21713,N_21776);
nand U22024 (N_22024,N_21897,N_21876);
nand U22025 (N_22025,N_21744,N_21757);
and U22026 (N_22026,N_21699,N_21672);
and U22027 (N_22027,N_21609,N_21749);
and U22028 (N_22028,N_21715,N_21869);
or U22029 (N_22029,N_21891,N_21737);
nand U22030 (N_22030,N_21607,N_21653);
xor U22031 (N_22031,N_21734,N_21718);
or U22032 (N_22032,N_21685,N_21846);
and U22033 (N_22033,N_21851,N_21804);
and U22034 (N_22034,N_21839,N_21816);
nand U22035 (N_22035,N_21669,N_21795);
nor U22036 (N_22036,N_21899,N_21706);
nor U22037 (N_22037,N_21835,N_21790);
xnor U22038 (N_22038,N_21874,N_21833);
nor U22039 (N_22039,N_21858,N_21612);
and U22040 (N_22040,N_21868,N_21884);
and U22041 (N_22041,N_21789,N_21722);
and U22042 (N_22042,N_21852,N_21812);
xnor U22043 (N_22043,N_21679,N_21773);
nand U22044 (N_22044,N_21634,N_21880);
nor U22045 (N_22045,N_21766,N_21604);
nand U22046 (N_22046,N_21797,N_21616);
nand U22047 (N_22047,N_21807,N_21637);
nor U22048 (N_22048,N_21798,N_21677);
and U22049 (N_22049,N_21875,N_21657);
and U22050 (N_22050,N_21653,N_21665);
nand U22051 (N_22051,N_21793,N_21811);
xnor U22052 (N_22052,N_21639,N_21880);
xnor U22053 (N_22053,N_21631,N_21764);
or U22054 (N_22054,N_21889,N_21820);
and U22055 (N_22055,N_21622,N_21731);
xnor U22056 (N_22056,N_21792,N_21740);
xnor U22057 (N_22057,N_21751,N_21789);
xor U22058 (N_22058,N_21845,N_21846);
or U22059 (N_22059,N_21645,N_21772);
or U22060 (N_22060,N_21878,N_21720);
nor U22061 (N_22061,N_21728,N_21741);
nand U22062 (N_22062,N_21827,N_21777);
xor U22063 (N_22063,N_21864,N_21862);
or U22064 (N_22064,N_21881,N_21871);
nand U22065 (N_22065,N_21796,N_21660);
or U22066 (N_22066,N_21844,N_21755);
nor U22067 (N_22067,N_21829,N_21845);
or U22068 (N_22068,N_21728,N_21754);
or U22069 (N_22069,N_21785,N_21747);
and U22070 (N_22070,N_21723,N_21660);
nand U22071 (N_22071,N_21727,N_21875);
and U22072 (N_22072,N_21723,N_21632);
nor U22073 (N_22073,N_21770,N_21726);
xor U22074 (N_22074,N_21711,N_21765);
or U22075 (N_22075,N_21698,N_21632);
and U22076 (N_22076,N_21831,N_21868);
and U22077 (N_22077,N_21622,N_21805);
nor U22078 (N_22078,N_21700,N_21835);
nand U22079 (N_22079,N_21728,N_21840);
and U22080 (N_22080,N_21709,N_21842);
nor U22081 (N_22081,N_21863,N_21711);
nand U22082 (N_22082,N_21664,N_21830);
and U22083 (N_22083,N_21613,N_21702);
nor U22084 (N_22084,N_21764,N_21893);
and U22085 (N_22085,N_21611,N_21651);
nand U22086 (N_22086,N_21737,N_21659);
xnor U22087 (N_22087,N_21699,N_21869);
xnor U22088 (N_22088,N_21648,N_21780);
or U22089 (N_22089,N_21716,N_21803);
nand U22090 (N_22090,N_21604,N_21624);
nand U22091 (N_22091,N_21892,N_21855);
and U22092 (N_22092,N_21749,N_21857);
xor U22093 (N_22093,N_21660,N_21694);
xnor U22094 (N_22094,N_21793,N_21786);
or U22095 (N_22095,N_21813,N_21781);
or U22096 (N_22096,N_21822,N_21633);
nor U22097 (N_22097,N_21877,N_21789);
nor U22098 (N_22098,N_21766,N_21809);
xnor U22099 (N_22099,N_21878,N_21651);
nor U22100 (N_22100,N_21656,N_21678);
nand U22101 (N_22101,N_21850,N_21725);
nor U22102 (N_22102,N_21816,N_21614);
nand U22103 (N_22103,N_21755,N_21857);
or U22104 (N_22104,N_21689,N_21614);
nand U22105 (N_22105,N_21817,N_21695);
or U22106 (N_22106,N_21650,N_21699);
nand U22107 (N_22107,N_21845,N_21882);
or U22108 (N_22108,N_21876,N_21838);
or U22109 (N_22109,N_21754,N_21627);
nand U22110 (N_22110,N_21644,N_21726);
xor U22111 (N_22111,N_21686,N_21870);
nor U22112 (N_22112,N_21752,N_21871);
and U22113 (N_22113,N_21613,N_21852);
or U22114 (N_22114,N_21633,N_21816);
nor U22115 (N_22115,N_21689,N_21816);
xnor U22116 (N_22116,N_21768,N_21652);
and U22117 (N_22117,N_21793,N_21721);
and U22118 (N_22118,N_21616,N_21827);
nor U22119 (N_22119,N_21805,N_21850);
nor U22120 (N_22120,N_21892,N_21757);
or U22121 (N_22121,N_21713,N_21675);
nand U22122 (N_22122,N_21895,N_21713);
or U22123 (N_22123,N_21623,N_21838);
or U22124 (N_22124,N_21697,N_21890);
and U22125 (N_22125,N_21794,N_21893);
or U22126 (N_22126,N_21693,N_21765);
nor U22127 (N_22127,N_21769,N_21883);
nor U22128 (N_22128,N_21879,N_21648);
and U22129 (N_22129,N_21858,N_21834);
or U22130 (N_22130,N_21758,N_21763);
and U22131 (N_22131,N_21711,N_21667);
nand U22132 (N_22132,N_21780,N_21657);
nand U22133 (N_22133,N_21723,N_21826);
xnor U22134 (N_22134,N_21815,N_21805);
or U22135 (N_22135,N_21865,N_21735);
or U22136 (N_22136,N_21884,N_21708);
nand U22137 (N_22137,N_21760,N_21630);
and U22138 (N_22138,N_21650,N_21830);
and U22139 (N_22139,N_21638,N_21774);
nor U22140 (N_22140,N_21821,N_21624);
nor U22141 (N_22141,N_21785,N_21878);
nor U22142 (N_22142,N_21688,N_21708);
nand U22143 (N_22143,N_21670,N_21795);
and U22144 (N_22144,N_21898,N_21642);
xor U22145 (N_22145,N_21606,N_21854);
xor U22146 (N_22146,N_21650,N_21703);
xor U22147 (N_22147,N_21837,N_21793);
nand U22148 (N_22148,N_21682,N_21781);
nand U22149 (N_22149,N_21663,N_21806);
and U22150 (N_22150,N_21818,N_21797);
or U22151 (N_22151,N_21652,N_21891);
nand U22152 (N_22152,N_21789,N_21661);
nand U22153 (N_22153,N_21871,N_21650);
nand U22154 (N_22154,N_21611,N_21704);
and U22155 (N_22155,N_21627,N_21770);
nor U22156 (N_22156,N_21819,N_21874);
xor U22157 (N_22157,N_21725,N_21797);
nand U22158 (N_22158,N_21808,N_21881);
nand U22159 (N_22159,N_21861,N_21615);
xor U22160 (N_22160,N_21723,N_21815);
nand U22161 (N_22161,N_21656,N_21720);
nand U22162 (N_22162,N_21690,N_21613);
nor U22163 (N_22163,N_21879,N_21765);
and U22164 (N_22164,N_21625,N_21630);
nand U22165 (N_22165,N_21647,N_21666);
xnor U22166 (N_22166,N_21666,N_21732);
and U22167 (N_22167,N_21669,N_21616);
or U22168 (N_22168,N_21701,N_21721);
xor U22169 (N_22169,N_21754,N_21720);
xnor U22170 (N_22170,N_21860,N_21850);
nand U22171 (N_22171,N_21728,N_21810);
xor U22172 (N_22172,N_21635,N_21847);
and U22173 (N_22173,N_21848,N_21601);
nor U22174 (N_22174,N_21717,N_21865);
nor U22175 (N_22175,N_21849,N_21856);
nor U22176 (N_22176,N_21822,N_21855);
or U22177 (N_22177,N_21701,N_21600);
nor U22178 (N_22178,N_21684,N_21713);
or U22179 (N_22179,N_21666,N_21854);
or U22180 (N_22180,N_21885,N_21828);
xor U22181 (N_22181,N_21718,N_21739);
and U22182 (N_22182,N_21693,N_21752);
xnor U22183 (N_22183,N_21719,N_21881);
xnor U22184 (N_22184,N_21698,N_21620);
or U22185 (N_22185,N_21824,N_21604);
nand U22186 (N_22186,N_21874,N_21640);
and U22187 (N_22187,N_21816,N_21809);
and U22188 (N_22188,N_21863,N_21885);
xor U22189 (N_22189,N_21612,N_21776);
nand U22190 (N_22190,N_21859,N_21611);
or U22191 (N_22191,N_21640,N_21663);
xnor U22192 (N_22192,N_21814,N_21760);
nor U22193 (N_22193,N_21728,N_21702);
nor U22194 (N_22194,N_21888,N_21822);
or U22195 (N_22195,N_21738,N_21635);
nand U22196 (N_22196,N_21879,N_21818);
or U22197 (N_22197,N_21678,N_21850);
and U22198 (N_22198,N_21848,N_21711);
or U22199 (N_22199,N_21701,N_21772);
xnor U22200 (N_22200,N_22160,N_22155);
xor U22201 (N_22201,N_22020,N_21970);
and U22202 (N_22202,N_21954,N_22152);
or U22203 (N_22203,N_21992,N_22034);
nand U22204 (N_22204,N_22029,N_21936);
and U22205 (N_22205,N_21988,N_22134);
or U22206 (N_22206,N_22195,N_21985);
nor U22207 (N_22207,N_21913,N_22005);
or U22208 (N_22208,N_22122,N_21958);
nor U22209 (N_22209,N_22197,N_22085);
xnor U22210 (N_22210,N_22135,N_21937);
nor U22211 (N_22211,N_21959,N_21961);
xor U22212 (N_22212,N_22076,N_22073);
and U22213 (N_22213,N_22196,N_22113);
nand U22214 (N_22214,N_21938,N_22080);
nor U22215 (N_22215,N_21950,N_21953);
nor U22216 (N_22216,N_22012,N_22043);
xor U22217 (N_22217,N_21928,N_22088);
and U22218 (N_22218,N_22054,N_22000);
nand U22219 (N_22219,N_22041,N_22006);
nor U22220 (N_22220,N_22079,N_22099);
or U22221 (N_22221,N_22101,N_22042);
nor U22222 (N_22222,N_22180,N_22121);
xor U22223 (N_22223,N_22014,N_21956);
nand U22224 (N_22224,N_22100,N_22116);
or U22225 (N_22225,N_21907,N_22036);
xor U22226 (N_22226,N_21947,N_22127);
xnor U22227 (N_22227,N_22071,N_21997);
and U22228 (N_22228,N_21952,N_22106);
nor U22229 (N_22229,N_22037,N_22138);
or U22230 (N_22230,N_21911,N_22115);
xor U22231 (N_22231,N_21978,N_21935);
nor U22232 (N_22232,N_22078,N_22188);
nor U22233 (N_22233,N_22062,N_21948);
xor U22234 (N_22234,N_22170,N_22181);
nor U22235 (N_22235,N_22091,N_21968);
or U22236 (N_22236,N_22064,N_21920);
and U22237 (N_22237,N_22132,N_22087);
xor U22238 (N_22238,N_22068,N_21957);
xnor U22239 (N_22239,N_22129,N_22137);
nor U22240 (N_22240,N_22175,N_22019);
nor U22241 (N_22241,N_22198,N_22163);
and U22242 (N_22242,N_22161,N_22103);
nor U22243 (N_22243,N_22090,N_22186);
and U22244 (N_22244,N_21990,N_22112);
and U22245 (N_22245,N_21965,N_22108);
nand U22246 (N_22246,N_22104,N_22011);
nand U22247 (N_22247,N_21998,N_22060);
xor U22248 (N_22248,N_21902,N_21991);
nor U22249 (N_22249,N_22070,N_21945);
and U22250 (N_22250,N_22040,N_22063);
and U22251 (N_22251,N_21946,N_22072);
nor U22252 (N_22252,N_21966,N_22086);
xnor U22253 (N_22253,N_21964,N_22109);
xnor U22254 (N_22254,N_22118,N_21942);
and U22255 (N_22255,N_21924,N_22117);
nor U22256 (N_22256,N_21923,N_22102);
nor U22257 (N_22257,N_22153,N_21934);
nand U22258 (N_22258,N_22001,N_21908);
and U22259 (N_22259,N_22199,N_22089);
and U22260 (N_22260,N_22147,N_22150);
and U22261 (N_22261,N_22067,N_22139);
or U22262 (N_22262,N_21962,N_22105);
xor U22263 (N_22263,N_22096,N_22059);
nand U22264 (N_22264,N_21915,N_22171);
and U22265 (N_22265,N_22003,N_21967);
and U22266 (N_22266,N_21993,N_21951);
and U22267 (N_22267,N_22154,N_21901);
xnor U22268 (N_22268,N_22023,N_22049);
xor U22269 (N_22269,N_22074,N_22050);
or U22270 (N_22270,N_22039,N_22182);
xor U22271 (N_22271,N_22002,N_21989);
nand U22272 (N_22272,N_21944,N_21999);
or U22273 (N_22273,N_21983,N_22094);
xor U22274 (N_22274,N_21939,N_22051);
xnor U22275 (N_22275,N_22008,N_22111);
xnor U22276 (N_22276,N_22107,N_22169);
or U22277 (N_22277,N_22084,N_21941);
and U22278 (N_22278,N_21917,N_21903);
xnor U22279 (N_22279,N_22095,N_21919);
nor U22280 (N_22280,N_21984,N_21974);
or U22281 (N_22281,N_22056,N_21931);
nand U22282 (N_22282,N_22128,N_22114);
or U22283 (N_22283,N_21976,N_21979);
xor U22284 (N_22284,N_22066,N_22031);
nor U22285 (N_22285,N_22032,N_21927);
and U22286 (N_22286,N_21996,N_22048);
and U22287 (N_22287,N_22166,N_21973);
nor U22288 (N_22288,N_22173,N_22053);
nand U22289 (N_22289,N_21986,N_21921);
and U22290 (N_22290,N_22168,N_21930);
or U22291 (N_22291,N_22082,N_22017);
or U22292 (N_22292,N_21982,N_21949);
or U22293 (N_22293,N_22184,N_22027);
and U22294 (N_22294,N_21960,N_22052);
nand U22295 (N_22295,N_22044,N_22013);
and U22296 (N_22296,N_22035,N_21943);
and U22297 (N_22297,N_21918,N_22024);
and U22298 (N_22298,N_22026,N_22022);
and U22299 (N_22299,N_22081,N_22176);
nand U22300 (N_22300,N_22038,N_22172);
nand U22301 (N_22301,N_21929,N_22016);
nor U22302 (N_22302,N_22021,N_22004);
xor U22303 (N_22303,N_22164,N_21916);
or U22304 (N_22304,N_22030,N_22045);
and U22305 (N_22305,N_22140,N_22185);
and U22306 (N_22306,N_22069,N_22167);
or U22307 (N_22307,N_22046,N_22162);
and U22308 (N_22308,N_22110,N_22025);
nand U22309 (N_22309,N_21971,N_22065);
or U22310 (N_22310,N_21963,N_22083);
and U22311 (N_22311,N_22028,N_22018);
nor U22312 (N_22312,N_22131,N_22192);
nand U22313 (N_22313,N_22077,N_22179);
nor U22314 (N_22314,N_21904,N_21925);
and U22315 (N_22315,N_21975,N_22119);
nand U22316 (N_22316,N_22149,N_22047);
or U22317 (N_22317,N_21995,N_22061);
nand U22318 (N_22318,N_22151,N_22143);
and U22319 (N_22319,N_21977,N_22177);
nand U22320 (N_22320,N_21955,N_22133);
and U22321 (N_22321,N_22165,N_22092);
or U22322 (N_22322,N_22194,N_22189);
and U22323 (N_22323,N_22057,N_21969);
or U22324 (N_22324,N_22075,N_21906);
and U22325 (N_22325,N_21980,N_21994);
nor U22326 (N_22326,N_22033,N_22130);
xor U22327 (N_22327,N_22142,N_22055);
nor U22328 (N_22328,N_21940,N_22136);
or U22329 (N_22329,N_22126,N_21932);
nor U22330 (N_22330,N_22146,N_22193);
nor U22331 (N_22331,N_21981,N_21933);
nor U22332 (N_22332,N_22125,N_22156);
xnor U22333 (N_22333,N_22098,N_21972);
nand U22334 (N_22334,N_22124,N_21912);
or U22335 (N_22335,N_22174,N_21922);
nor U22336 (N_22336,N_21909,N_22148);
or U22337 (N_22337,N_22159,N_21987);
xnor U22338 (N_22338,N_22010,N_21914);
nor U22339 (N_22339,N_22190,N_22144);
and U22340 (N_22340,N_22178,N_22093);
xor U22341 (N_22341,N_22123,N_22141);
and U22342 (N_22342,N_22015,N_22058);
xnor U22343 (N_22343,N_22187,N_21905);
nor U22344 (N_22344,N_22183,N_22158);
xnor U22345 (N_22345,N_22009,N_21926);
xnor U22346 (N_22346,N_22120,N_22007);
nor U22347 (N_22347,N_22157,N_22191);
nand U22348 (N_22348,N_21910,N_22145);
or U22349 (N_22349,N_21900,N_22097);
and U22350 (N_22350,N_22079,N_22017);
and U22351 (N_22351,N_21955,N_21974);
or U22352 (N_22352,N_22122,N_22001);
xnor U22353 (N_22353,N_21933,N_21958);
and U22354 (N_22354,N_22125,N_21944);
xor U22355 (N_22355,N_21949,N_21965);
xor U22356 (N_22356,N_22092,N_22041);
xnor U22357 (N_22357,N_22155,N_21989);
xnor U22358 (N_22358,N_21960,N_22188);
xnor U22359 (N_22359,N_21972,N_22115);
and U22360 (N_22360,N_22152,N_22078);
nor U22361 (N_22361,N_21997,N_21934);
or U22362 (N_22362,N_22179,N_22121);
and U22363 (N_22363,N_22034,N_22089);
or U22364 (N_22364,N_22048,N_21901);
nor U22365 (N_22365,N_21962,N_21948);
nand U22366 (N_22366,N_21975,N_22195);
nand U22367 (N_22367,N_21951,N_21985);
and U22368 (N_22368,N_22025,N_21934);
and U22369 (N_22369,N_22052,N_21972);
nor U22370 (N_22370,N_22023,N_21909);
xor U22371 (N_22371,N_22193,N_22107);
xor U22372 (N_22372,N_22094,N_21939);
and U22373 (N_22373,N_21949,N_22110);
xnor U22374 (N_22374,N_22018,N_21963);
or U22375 (N_22375,N_22186,N_21904);
nor U22376 (N_22376,N_21991,N_21901);
nor U22377 (N_22377,N_22124,N_21937);
nor U22378 (N_22378,N_22173,N_21952);
and U22379 (N_22379,N_21913,N_21936);
nand U22380 (N_22380,N_22181,N_22048);
nor U22381 (N_22381,N_22060,N_22084);
nor U22382 (N_22382,N_22111,N_22102);
and U22383 (N_22383,N_21989,N_22030);
xor U22384 (N_22384,N_22144,N_22142);
and U22385 (N_22385,N_21948,N_22116);
nor U22386 (N_22386,N_21978,N_22147);
xnor U22387 (N_22387,N_22159,N_21980);
nand U22388 (N_22388,N_22141,N_22039);
nand U22389 (N_22389,N_21912,N_21999);
or U22390 (N_22390,N_21939,N_21971);
nand U22391 (N_22391,N_22007,N_22054);
and U22392 (N_22392,N_21914,N_22189);
and U22393 (N_22393,N_22038,N_22076);
or U22394 (N_22394,N_22143,N_22071);
nor U22395 (N_22395,N_21950,N_22064);
and U22396 (N_22396,N_22176,N_21942);
nand U22397 (N_22397,N_22116,N_22039);
xnor U22398 (N_22398,N_22161,N_22122);
xnor U22399 (N_22399,N_21974,N_22048);
nand U22400 (N_22400,N_21909,N_22047);
and U22401 (N_22401,N_22155,N_21991);
xnor U22402 (N_22402,N_22053,N_22141);
nand U22403 (N_22403,N_21914,N_22065);
or U22404 (N_22404,N_21920,N_21952);
nand U22405 (N_22405,N_22097,N_22100);
and U22406 (N_22406,N_21907,N_21926);
or U22407 (N_22407,N_22049,N_22073);
nor U22408 (N_22408,N_22082,N_21921);
and U22409 (N_22409,N_22153,N_22061);
nand U22410 (N_22410,N_22138,N_22192);
nand U22411 (N_22411,N_22168,N_21975);
or U22412 (N_22412,N_22149,N_21960);
or U22413 (N_22413,N_22093,N_22047);
xor U22414 (N_22414,N_22028,N_21905);
nand U22415 (N_22415,N_22041,N_22085);
xnor U22416 (N_22416,N_21910,N_21935);
xnor U22417 (N_22417,N_21937,N_22100);
or U22418 (N_22418,N_22110,N_21967);
xnor U22419 (N_22419,N_21938,N_22108);
nor U22420 (N_22420,N_21996,N_22037);
and U22421 (N_22421,N_22050,N_21912);
and U22422 (N_22422,N_22120,N_22186);
xnor U22423 (N_22423,N_22008,N_21995);
and U22424 (N_22424,N_22102,N_22107);
and U22425 (N_22425,N_21983,N_22174);
nor U22426 (N_22426,N_22171,N_22121);
and U22427 (N_22427,N_22040,N_22014);
and U22428 (N_22428,N_22101,N_22178);
xnor U22429 (N_22429,N_21945,N_22170);
nand U22430 (N_22430,N_22044,N_22065);
or U22431 (N_22431,N_22049,N_22074);
nor U22432 (N_22432,N_22008,N_22178);
xnor U22433 (N_22433,N_22022,N_21965);
nand U22434 (N_22434,N_22005,N_21945);
nand U22435 (N_22435,N_22193,N_22159);
nor U22436 (N_22436,N_22198,N_22098);
nor U22437 (N_22437,N_22152,N_22132);
nand U22438 (N_22438,N_21912,N_22041);
and U22439 (N_22439,N_22068,N_22077);
xor U22440 (N_22440,N_22106,N_22011);
nor U22441 (N_22441,N_21982,N_22110);
xnor U22442 (N_22442,N_22055,N_22124);
and U22443 (N_22443,N_22172,N_22077);
nor U22444 (N_22444,N_21993,N_22137);
xor U22445 (N_22445,N_21909,N_22042);
and U22446 (N_22446,N_22036,N_22065);
and U22447 (N_22447,N_22117,N_21908);
and U22448 (N_22448,N_22141,N_21993);
xor U22449 (N_22449,N_21913,N_22061);
nor U22450 (N_22450,N_22057,N_21919);
or U22451 (N_22451,N_21953,N_21910);
nor U22452 (N_22452,N_21962,N_22056);
nand U22453 (N_22453,N_21980,N_22037);
xnor U22454 (N_22454,N_22061,N_22093);
nand U22455 (N_22455,N_22024,N_22168);
and U22456 (N_22456,N_22008,N_21953);
nand U22457 (N_22457,N_21984,N_22150);
or U22458 (N_22458,N_21903,N_22014);
nor U22459 (N_22459,N_22139,N_22152);
nand U22460 (N_22460,N_22146,N_21978);
nor U22461 (N_22461,N_21947,N_22143);
nor U22462 (N_22462,N_22115,N_21964);
nor U22463 (N_22463,N_22002,N_22011);
and U22464 (N_22464,N_21980,N_22174);
and U22465 (N_22465,N_22099,N_21997);
nand U22466 (N_22466,N_22013,N_21963);
and U22467 (N_22467,N_22016,N_22091);
and U22468 (N_22468,N_21915,N_22077);
nand U22469 (N_22469,N_22029,N_22040);
or U22470 (N_22470,N_22155,N_21918);
and U22471 (N_22471,N_22000,N_21931);
nor U22472 (N_22472,N_21907,N_22145);
or U22473 (N_22473,N_22118,N_22015);
xnor U22474 (N_22474,N_21961,N_21932);
nand U22475 (N_22475,N_21960,N_21963);
or U22476 (N_22476,N_22135,N_22007);
xnor U22477 (N_22477,N_22072,N_22147);
or U22478 (N_22478,N_22087,N_21982);
xnor U22479 (N_22479,N_21957,N_21900);
nor U22480 (N_22480,N_22087,N_22117);
xor U22481 (N_22481,N_21948,N_21976);
or U22482 (N_22482,N_22069,N_22184);
nand U22483 (N_22483,N_21918,N_22110);
nor U22484 (N_22484,N_21928,N_22127);
or U22485 (N_22485,N_22107,N_22160);
or U22486 (N_22486,N_21933,N_21996);
or U22487 (N_22487,N_22011,N_22122);
nor U22488 (N_22488,N_22143,N_22173);
xor U22489 (N_22489,N_21960,N_21916);
and U22490 (N_22490,N_22138,N_21977);
nor U22491 (N_22491,N_21970,N_22193);
and U22492 (N_22492,N_21943,N_21940);
xnor U22493 (N_22493,N_22169,N_22002);
or U22494 (N_22494,N_21946,N_22125);
nor U22495 (N_22495,N_22111,N_22147);
or U22496 (N_22496,N_21986,N_22141);
nor U22497 (N_22497,N_22075,N_21960);
nand U22498 (N_22498,N_21952,N_21955);
or U22499 (N_22499,N_22101,N_21983);
nor U22500 (N_22500,N_22237,N_22436);
or U22501 (N_22501,N_22415,N_22404);
nor U22502 (N_22502,N_22482,N_22323);
nand U22503 (N_22503,N_22213,N_22255);
and U22504 (N_22504,N_22467,N_22478);
nor U22505 (N_22505,N_22310,N_22325);
or U22506 (N_22506,N_22433,N_22201);
or U22507 (N_22507,N_22494,N_22422);
nand U22508 (N_22508,N_22267,N_22400);
or U22509 (N_22509,N_22202,N_22474);
nand U22510 (N_22510,N_22289,N_22245);
nor U22511 (N_22511,N_22394,N_22428);
or U22512 (N_22512,N_22445,N_22456);
and U22513 (N_22513,N_22446,N_22409);
nor U22514 (N_22514,N_22278,N_22439);
nor U22515 (N_22515,N_22320,N_22357);
and U22516 (N_22516,N_22455,N_22443);
or U22517 (N_22517,N_22218,N_22485);
or U22518 (N_22518,N_22497,N_22376);
nor U22519 (N_22519,N_22227,N_22204);
nor U22520 (N_22520,N_22339,N_22381);
or U22521 (N_22521,N_22366,N_22312);
or U22522 (N_22522,N_22252,N_22346);
nand U22523 (N_22523,N_22276,N_22374);
and U22524 (N_22524,N_22210,N_22209);
nand U22525 (N_22525,N_22380,N_22224);
or U22526 (N_22526,N_22242,N_22230);
or U22527 (N_22527,N_22345,N_22269);
or U22528 (N_22528,N_22353,N_22338);
nor U22529 (N_22529,N_22238,N_22387);
nand U22530 (N_22530,N_22483,N_22321);
xnor U22531 (N_22531,N_22491,N_22362);
xnor U22532 (N_22532,N_22484,N_22275);
or U22533 (N_22533,N_22368,N_22486);
nand U22534 (N_22534,N_22263,N_22231);
or U22535 (N_22535,N_22383,N_22492);
xor U22536 (N_22536,N_22498,N_22305);
and U22537 (N_22537,N_22216,N_22359);
nand U22538 (N_22538,N_22264,N_22298);
and U22539 (N_22539,N_22297,N_22369);
or U22540 (N_22540,N_22435,N_22370);
and U22541 (N_22541,N_22342,N_22473);
and U22542 (N_22542,N_22408,N_22225);
and U22543 (N_22543,N_22287,N_22453);
nor U22544 (N_22544,N_22322,N_22277);
nor U22545 (N_22545,N_22481,N_22270);
nor U22546 (N_22546,N_22244,N_22337);
nor U22547 (N_22547,N_22349,N_22308);
nand U22548 (N_22548,N_22416,N_22313);
nand U22549 (N_22549,N_22347,N_22295);
or U22550 (N_22550,N_22356,N_22226);
or U22551 (N_22551,N_22360,N_22442);
xnor U22552 (N_22552,N_22214,N_22296);
xnor U22553 (N_22553,N_22493,N_22253);
nor U22554 (N_22554,N_22476,N_22273);
nor U22555 (N_22555,N_22251,N_22215);
nor U22556 (N_22556,N_22450,N_22274);
nor U22557 (N_22557,N_22340,N_22365);
and U22558 (N_22558,N_22470,N_22327);
xnor U22559 (N_22559,N_22306,N_22315);
and U22560 (N_22560,N_22441,N_22240);
xnor U22561 (N_22561,N_22316,N_22303);
nand U22562 (N_22562,N_22487,N_22311);
and U22563 (N_22563,N_22413,N_22351);
nand U22564 (N_22564,N_22336,N_22421);
and U22565 (N_22565,N_22375,N_22432);
and U22566 (N_22566,N_22265,N_22477);
nor U22567 (N_22567,N_22454,N_22222);
nand U22568 (N_22568,N_22283,N_22488);
xnor U22569 (N_22569,N_22377,N_22348);
and U22570 (N_22570,N_22268,N_22250);
or U22571 (N_22571,N_22479,N_22290);
or U22572 (N_22572,N_22334,N_22248);
nor U22573 (N_22573,N_22466,N_22367);
nand U22574 (N_22574,N_22355,N_22458);
nor U22575 (N_22575,N_22341,N_22233);
xor U22576 (N_22576,N_22438,N_22480);
nand U22577 (N_22577,N_22364,N_22472);
nand U22578 (N_22578,N_22257,N_22460);
nor U22579 (N_22579,N_22330,N_22280);
and U22580 (N_22580,N_22241,N_22372);
nand U22581 (N_22581,N_22399,N_22329);
and U22582 (N_22582,N_22457,N_22302);
nand U22583 (N_22583,N_22489,N_22284);
or U22584 (N_22584,N_22314,N_22464);
or U22585 (N_22585,N_22324,N_22221);
and U22586 (N_22586,N_22282,N_22319);
nand U22587 (N_22587,N_22254,N_22392);
xnor U22588 (N_22588,N_22462,N_22328);
nor U22589 (N_22589,N_22206,N_22326);
or U22590 (N_22590,N_22468,N_22279);
or U22591 (N_22591,N_22304,N_22220);
xor U22592 (N_22592,N_22317,N_22403);
xnor U22593 (N_22593,N_22299,N_22223);
nor U22594 (N_22594,N_22256,N_22475);
or U22595 (N_22595,N_22379,N_22496);
and U22596 (N_22596,N_22291,N_22207);
nor U22597 (N_22597,N_22499,N_22373);
or U22598 (N_22598,N_22262,N_22208);
nor U22599 (N_22599,N_22333,N_22294);
and U22600 (N_22600,N_22437,N_22419);
xor U22601 (N_22601,N_22463,N_22412);
nor U22602 (N_22602,N_22350,N_22212);
or U22603 (N_22603,N_22200,N_22363);
and U22604 (N_22604,N_22471,N_22246);
and U22605 (N_22605,N_22239,N_22449);
nor U22606 (N_22606,N_22229,N_22247);
nand U22607 (N_22607,N_22461,N_22281);
or U22608 (N_22608,N_22424,N_22411);
and U22609 (N_22609,N_22258,N_22249);
or U22610 (N_22610,N_22417,N_22234);
nor U22611 (N_22611,N_22371,N_22382);
nand U22612 (N_22612,N_22228,N_22384);
and U22613 (N_22613,N_22398,N_22318);
xor U22614 (N_22614,N_22393,N_22406);
xor U22615 (N_22615,N_22459,N_22465);
or U22616 (N_22616,N_22358,N_22451);
nor U22617 (N_22617,N_22469,N_22378);
nor U22618 (N_22618,N_22288,N_22495);
nor U22619 (N_22619,N_22236,N_22331);
or U22620 (N_22620,N_22452,N_22388);
nor U22621 (N_22621,N_22397,N_22401);
and U22622 (N_22622,N_22448,N_22285);
or U22623 (N_22623,N_22211,N_22447);
nand U22624 (N_22624,N_22418,N_22391);
nand U22625 (N_22625,N_22490,N_22420);
nor U22626 (N_22626,N_22430,N_22405);
or U22627 (N_22627,N_22260,N_22243);
nor U22628 (N_22628,N_22352,N_22232);
nand U22629 (N_22629,N_22292,N_22335);
and U22630 (N_22630,N_22385,N_22414);
and U22631 (N_22631,N_22390,N_22444);
or U22632 (N_22632,N_22272,N_22361);
or U22633 (N_22633,N_22389,N_22344);
nor U22634 (N_22634,N_22407,N_22425);
or U22635 (N_22635,N_22219,N_22266);
and U22636 (N_22636,N_22307,N_22300);
and U22637 (N_22637,N_22259,N_22235);
nor U22638 (N_22638,N_22271,N_22217);
nand U22639 (N_22639,N_22431,N_22354);
nor U22640 (N_22640,N_22286,N_22434);
xor U22641 (N_22641,N_22309,N_22426);
nand U22642 (N_22642,N_22427,N_22293);
and U22643 (N_22643,N_22440,N_22402);
and U22644 (N_22644,N_22429,N_22205);
nor U22645 (N_22645,N_22423,N_22301);
nor U22646 (N_22646,N_22261,N_22386);
and U22647 (N_22647,N_22343,N_22332);
nand U22648 (N_22648,N_22203,N_22395);
nand U22649 (N_22649,N_22410,N_22396);
xnor U22650 (N_22650,N_22313,N_22304);
or U22651 (N_22651,N_22392,N_22454);
or U22652 (N_22652,N_22348,N_22400);
or U22653 (N_22653,N_22367,N_22372);
xnor U22654 (N_22654,N_22468,N_22434);
nor U22655 (N_22655,N_22499,N_22223);
and U22656 (N_22656,N_22375,N_22457);
xor U22657 (N_22657,N_22480,N_22496);
nor U22658 (N_22658,N_22222,N_22435);
and U22659 (N_22659,N_22366,N_22249);
nor U22660 (N_22660,N_22266,N_22338);
nor U22661 (N_22661,N_22265,N_22388);
nand U22662 (N_22662,N_22447,N_22262);
xor U22663 (N_22663,N_22254,N_22350);
nor U22664 (N_22664,N_22491,N_22492);
and U22665 (N_22665,N_22447,N_22202);
or U22666 (N_22666,N_22302,N_22470);
xor U22667 (N_22667,N_22446,N_22495);
nand U22668 (N_22668,N_22363,N_22485);
or U22669 (N_22669,N_22435,N_22229);
nand U22670 (N_22670,N_22432,N_22494);
and U22671 (N_22671,N_22394,N_22304);
and U22672 (N_22672,N_22274,N_22458);
and U22673 (N_22673,N_22474,N_22250);
nand U22674 (N_22674,N_22362,N_22495);
nor U22675 (N_22675,N_22428,N_22446);
nor U22676 (N_22676,N_22480,N_22331);
nand U22677 (N_22677,N_22460,N_22314);
nand U22678 (N_22678,N_22417,N_22393);
xnor U22679 (N_22679,N_22405,N_22454);
nor U22680 (N_22680,N_22324,N_22435);
and U22681 (N_22681,N_22352,N_22462);
nor U22682 (N_22682,N_22239,N_22226);
nand U22683 (N_22683,N_22222,N_22215);
xor U22684 (N_22684,N_22326,N_22424);
xor U22685 (N_22685,N_22321,N_22412);
or U22686 (N_22686,N_22334,N_22373);
or U22687 (N_22687,N_22312,N_22259);
xnor U22688 (N_22688,N_22343,N_22291);
nor U22689 (N_22689,N_22246,N_22450);
and U22690 (N_22690,N_22410,N_22479);
and U22691 (N_22691,N_22468,N_22426);
nand U22692 (N_22692,N_22429,N_22329);
xnor U22693 (N_22693,N_22366,N_22258);
and U22694 (N_22694,N_22262,N_22215);
and U22695 (N_22695,N_22381,N_22438);
nand U22696 (N_22696,N_22229,N_22238);
or U22697 (N_22697,N_22384,N_22269);
and U22698 (N_22698,N_22386,N_22401);
and U22699 (N_22699,N_22215,N_22322);
and U22700 (N_22700,N_22253,N_22331);
nor U22701 (N_22701,N_22284,N_22281);
nand U22702 (N_22702,N_22438,N_22495);
and U22703 (N_22703,N_22230,N_22269);
xor U22704 (N_22704,N_22234,N_22290);
and U22705 (N_22705,N_22265,N_22323);
nor U22706 (N_22706,N_22491,N_22468);
nand U22707 (N_22707,N_22436,N_22281);
and U22708 (N_22708,N_22478,N_22392);
and U22709 (N_22709,N_22303,N_22407);
or U22710 (N_22710,N_22394,N_22268);
and U22711 (N_22711,N_22434,N_22463);
nand U22712 (N_22712,N_22293,N_22444);
and U22713 (N_22713,N_22348,N_22204);
or U22714 (N_22714,N_22341,N_22223);
and U22715 (N_22715,N_22266,N_22337);
nand U22716 (N_22716,N_22234,N_22464);
nand U22717 (N_22717,N_22428,N_22212);
xnor U22718 (N_22718,N_22440,N_22317);
nand U22719 (N_22719,N_22230,N_22379);
xnor U22720 (N_22720,N_22437,N_22314);
xor U22721 (N_22721,N_22285,N_22396);
nor U22722 (N_22722,N_22497,N_22384);
nand U22723 (N_22723,N_22412,N_22358);
xnor U22724 (N_22724,N_22262,N_22368);
nand U22725 (N_22725,N_22432,N_22290);
nor U22726 (N_22726,N_22216,N_22269);
nor U22727 (N_22727,N_22248,N_22263);
xor U22728 (N_22728,N_22491,N_22411);
or U22729 (N_22729,N_22461,N_22326);
and U22730 (N_22730,N_22376,N_22209);
nand U22731 (N_22731,N_22418,N_22379);
or U22732 (N_22732,N_22218,N_22403);
nor U22733 (N_22733,N_22226,N_22306);
or U22734 (N_22734,N_22407,N_22285);
or U22735 (N_22735,N_22241,N_22205);
and U22736 (N_22736,N_22436,N_22358);
or U22737 (N_22737,N_22331,N_22465);
and U22738 (N_22738,N_22495,N_22207);
xor U22739 (N_22739,N_22492,N_22318);
nor U22740 (N_22740,N_22397,N_22301);
nand U22741 (N_22741,N_22467,N_22443);
nor U22742 (N_22742,N_22454,N_22200);
nand U22743 (N_22743,N_22390,N_22357);
nand U22744 (N_22744,N_22362,N_22368);
or U22745 (N_22745,N_22300,N_22390);
xnor U22746 (N_22746,N_22369,N_22437);
or U22747 (N_22747,N_22242,N_22385);
nor U22748 (N_22748,N_22401,N_22312);
nor U22749 (N_22749,N_22444,N_22372);
nand U22750 (N_22750,N_22378,N_22457);
nand U22751 (N_22751,N_22265,N_22382);
or U22752 (N_22752,N_22440,N_22280);
and U22753 (N_22753,N_22415,N_22475);
nor U22754 (N_22754,N_22496,N_22393);
nor U22755 (N_22755,N_22238,N_22291);
or U22756 (N_22756,N_22269,N_22427);
and U22757 (N_22757,N_22321,N_22332);
or U22758 (N_22758,N_22271,N_22398);
or U22759 (N_22759,N_22463,N_22252);
nand U22760 (N_22760,N_22490,N_22450);
and U22761 (N_22761,N_22272,N_22494);
nand U22762 (N_22762,N_22331,N_22358);
or U22763 (N_22763,N_22230,N_22393);
or U22764 (N_22764,N_22209,N_22401);
nor U22765 (N_22765,N_22316,N_22310);
xor U22766 (N_22766,N_22484,N_22237);
nand U22767 (N_22767,N_22303,N_22406);
nand U22768 (N_22768,N_22372,N_22249);
nor U22769 (N_22769,N_22298,N_22430);
xnor U22770 (N_22770,N_22291,N_22372);
nand U22771 (N_22771,N_22255,N_22346);
nand U22772 (N_22772,N_22335,N_22408);
xor U22773 (N_22773,N_22497,N_22404);
or U22774 (N_22774,N_22317,N_22427);
nor U22775 (N_22775,N_22411,N_22225);
and U22776 (N_22776,N_22288,N_22398);
xnor U22777 (N_22777,N_22250,N_22224);
and U22778 (N_22778,N_22351,N_22436);
or U22779 (N_22779,N_22483,N_22201);
or U22780 (N_22780,N_22383,N_22234);
and U22781 (N_22781,N_22481,N_22475);
nor U22782 (N_22782,N_22417,N_22281);
nor U22783 (N_22783,N_22305,N_22206);
nand U22784 (N_22784,N_22278,N_22402);
or U22785 (N_22785,N_22430,N_22297);
nand U22786 (N_22786,N_22456,N_22291);
xor U22787 (N_22787,N_22413,N_22421);
or U22788 (N_22788,N_22273,N_22247);
and U22789 (N_22789,N_22307,N_22352);
or U22790 (N_22790,N_22288,N_22486);
and U22791 (N_22791,N_22202,N_22445);
nand U22792 (N_22792,N_22314,N_22408);
xor U22793 (N_22793,N_22479,N_22241);
or U22794 (N_22794,N_22267,N_22201);
nand U22795 (N_22795,N_22361,N_22248);
xnor U22796 (N_22796,N_22373,N_22473);
xor U22797 (N_22797,N_22263,N_22423);
xor U22798 (N_22798,N_22460,N_22471);
or U22799 (N_22799,N_22431,N_22424);
or U22800 (N_22800,N_22675,N_22643);
xnor U22801 (N_22801,N_22780,N_22599);
or U22802 (N_22802,N_22687,N_22559);
or U22803 (N_22803,N_22594,N_22688);
nand U22804 (N_22804,N_22770,N_22558);
nor U22805 (N_22805,N_22690,N_22564);
xor U22806 (N_22806,N_22792,N_22700);
and U22807 (N_22807,N_22680,N_22771);
xor U22808 (N_22808,N_22501,N_22672);
or U22809 (N_22809,N_22600,N_22767);
or U22810 (N_22810,N_22537,N_22717);
nor U22811 (N_22811,N_22679,N_22797);
or U22812 (N_22812,N_22569,N_22713);
xnor U22813 (N_22813,N_22755,N_22540);
and U22814 (N_22814,N_22794,N_22693);
and U22815 (N_22815,N_22533,N_22519);
and U22816 (N_22816,N_22644,N_22779);
xor U22817 (N_22817,N_22622,N_22646);
or U22818 (N_22818,N_22798,N_22743);
nand U22819 (N_22819,N_22510,N_22671);
nand U22820 (N_22820,N_22793,N_22545);
nand U22821 (N_22821,N_22721,N_22546);
xor U22822 (N_22822,N_22746,N_22560);
or U22823 (N_22823,N_22758,N_22511);
or U22824 (N_22824,N_22528,N_22682);
or U22825 (N_22825,N_22623,N_22653);
nor U22826 (N_22826,N_22584,N_22661);
and U22827 (N_22827,N_22503,N_22650);
nor U22828 (N_22828,N_22681,N_22762);
nor U22829 (N_22829,N_22570,N_22520);
nand U22830 (N_22830,N_22553,N_22589);
xor U22831 (N_22831,N_22765,N_22749);
xnor U22832 (N_22832,N_22581,N_22575);
xor U22833 (N_22833,N_22506,N_22522);
or U22834 (N_22834,N_22524,N_22636);
and U22835 (N_22835,N_22566,N_22605);
xor U22836 (N_22836,N_22773,N_22544);
or U22837 (N_22837,N_22696,N_22515);
and U22838 (N_22838,N_22538,N_22527);
nor U22839 (N_22839,N_22631,N_22722);
or U22840 (N_22840,N_22763,N_22744);
nand U22841 (N_22841,N_22638,N_22645);
and U22842 (N_22842,N_22610,N_22627);
xnor U22843 (N_22843,N_22572,N_22730);
xnor U22844 (N_22844,N_22669,N_22548);
and U22845 (N_22845,N_22521,N_22709);
nand U22846 (N_22846,N_22543,N_22563);
and U22847 (N_22847,N_22766,N_22505);
xnor U22848 (N_22848,N_22657,N_22651);
or U22849 (N_22849,N_22656,N_22635);
xor U22850 (N_22850,N_22789,N_22714);
and U22851 (N_22851,N_22590,N_22711);
xor U22852 (N_22852,N_22726,N_22745);
or U22853 (N_22853,N_22788,N_22565);
xor U22854 (N_22854,N_22684,N_22772);
or U22855 (N_22855,N_22579,N_22629);
and U22856 (N_22856,N_22534,N_22642);
xnor U22857 (N_22857,N_22753,N_22740);
xnor U22858 (N_22858,N_22757,N_22598);
or U22859 (N_22859,N_22787,N_22786);
nor U22860 (N_22860,N_22582,N_22585);
xnor U22861 (N_22861,N_22702,N_22776);
nor U22862 (N_22862,N_22677,N_22561);
and U22863 (N_22863,N_22716,N_22775);
and U22864 (N_22864,N_22507,N_22768);
xnor U22865 (N_22865,N_22574,N_22531);
nand U22866 (N_22866,N_22514,N_22735);
nor U22867 (N_22867,N_22576,N_22715);
and U22868 (N_22868,N_22781,N_22573);
or U22869 (N_22869,N_22760,N_22718);
nand U22870 (N_22870,N_22790,N_22603);
nand U22871 (N_22871,N_22625,N_22504);
nor U22872 (N_22872,N_22759,N_22748);
nand U22873 (N_22873,N_22778,N_22648);
xnor U22874 (N_22874,N_22796,N_22554);
nor U22875 (N_22875,N_22652,N_22706);
xor U22876 (N_22876,N_22666,N_22583);
xnor U22877 (N_22877,N_22799,N_22615);
or U22878 (N_22878,N_22526,N_22783);
nand U22879 (N_22879,N_22604,N_22791);
xor U22880 (N_22880,N_22729,N_22611);
and U22881 (N_22881,N_22731,N_22725);
nand U22882 (N_22882,N_22723,N_22707);
xnor U22883 (N_22883,N_22633,N_22597);
nand U22884 (N_22884,N_22676,N_22703);
xnor U22885 (N_22885,N_22624,N_22734);
or U22886 (N_22886,N_22609,N_22660);
xnor U22887 (N_22887,N_22732,N_22769);
or U22888 (N_22888,N_22518,N_22742);
xor U22889 (N_22889,N_22606,N_22513);
nor U22890 (N_22890,N_22712,N_22694);
nor U22891 (N_22891,N_22664,N_22630);
and U22892 (N_22892,N_22761,N_22542);
or U22893 (N_22893,N_22502,N_22632);
nand U22894 (N_22894,N_22752,N_22557);
nand U22895 (N_22895,N_22555,N_22512);
and U22896 (N_22896,N_22620,N_22591);
or U22897 (N_22897,N_22782,N_22785);
nand U22898 (N_22898,N_22649,N_22739);
nand U22899 (N_22899,N_22530,N_22626);
or U22900 (N_22900,N_22509,N_22754);
or U22901 (N_22901,N_22710,N_22549);
nand U22902 (N_22902,N_22568,N_22724);
nand U22903 (N_22903,N_22665,N_22601);
xor U22904 (N_22904,N_22613,N_22634);
or U22905 (N_22905,N_22750,N_22689);
and U22906 (N_22906,N_22580,N_22532);
and U22907 (N_22907,N_22741,N_22697);
nor U22908 (N_22908,N_22727,N_22567);
or U22909 (N_22909,N_22662,N_22678);
nand U22910 (N_22910,N_22593,N_22500);
nor U22911 (N_22911,N_22618,N_22547);
nor U22912 (N_22912,N_22562,N_22586);
and U22913 (N_22913,N_22704,N_22578);
or U22914 (N_22914,N_22673,N_22535);
nor U22915 (N_22915,N_22736,N_22602);
or U22916 (N_22916,N_22508,N_22747);
and U22917 (N_22917,N_22667,N_22708);
nor U22918 (N_22918,N_22616,N_22647);
nand U22919 (N_22919,N_22637,N_22571);
nand U22920 (N_22920,N_22516,N_22720);
or U22921 (N_22921,N_22751,N_22621);
and U22922 (N_22922,N_22738,N_22592);
or U22923 (N_22923,N_22517,N_22784);
nor U22924 (N_22924,N_22686,N_22663);
and U22925 (N_22925,N_22777,N_22588);
or U22926 (N_22926,N_22541,N_22698);
nand U22927 (N_22927,N_22655,N_22685);
nand U22928 (N_22928,N_22699,N_22639);
and U22929 (N_22929,N_22536,N_22701);
xnor U22930 (N_22930,N_22587,N_22692);
xnor U22931 (N_22931,N_22595,N_22577);
and U22932 (N_22932,N_22764,N_22525);
and U22933 (N_22933,N_22691,N_22719);
and U22934 (N_22934,N_22756,N_22539);
and U22935 (N_22935,N_22640,N_22658);
and U22936 (N_22936,N_22733,N_22552);
nand U22937 (N_22937,N_22617,N_22556);
or U22938 (N_22938,N_22607,N_22654);
xnor U22939 (N_22939,N_22612,N_22529);
nand U22940 (N_22940,N_22737,N_22619);
nor U22941 (N_22941,N_22596,N_22705);
xor U22942 (N_22942,N_22668,N_22608);
nor U22943 (N_22943,N_22674,N_22695);
nand U22944 (N_22944,N_22614,N_22550);
or U22945 (N_22945,N_22670,N_22683);
nand U22946 (N_22946,N_22551,N_22795);
nor U22947 (N_22947,N_22523,N_22728);
nor U22948 (N_22948,N_22659,N_22641);
nand U22949 (N_22949,N_22774,N_22628);
or U22950 (N_22950,N_22712,N_22600);
nand U22951 (N_22951,N_22599,N_22616);
xor U22952 (N_22952,N_22710,N_22584);
nor U22953 (N_22953,N_22549,N_22599);
and U22954 (N_22954,N_22697,N_22735);
xnor U22955 (N_22955,N_22694,N_22579);
nand U22956 (N_22956,N_22605,N_22670);
xnor U22957 (N_22957,N_22658,N_22788);
and U22958 (N_22958,N_22730,N_22775);
and U22959 (N_22959,N_22742,N_22758);
nand U22960 (N_22960,N_22533,N_22602);
nor U22961 (N_22961,N_22727,N_22646);
nor U22962 (N_22962,N_22607,N_22538);
nand U22963 (N_22963,N_22575,N_22548);
xnor U22964 (N_22964,N_22788,N_22762);
nor U22965 (N_22965,N_22606,N_22753);
nand U22966 (N_22966,N_22760,N_22714);
nand U22967 (N_22967,N_22700,N_22603);
and U22968 (N_22968,N_22578,N_22799);
xnor U22969 (N_22969,N_22583,N_22710);
nand U22970 (N_22970,N_22533,N_22663);
nand U22971 (N_22971,N_22679,N_22657);
nor U22972 (N_22972,N_22785,N_22717);
or U22973 (N_22973,N_22775,N_22635);
and U22974 (N_22974,N_22505,N_22521);
and U22975 (N_22975,N_22675,N_22736);
or U22976 (N_22976,N_22644,N_22652);
nor U22977 (N_22977,N_22667,N_22555);
or U22978 (N_22978,N_22651,N_22511);
or U22979 (N_22979,N_22600,N_22565);
or U22980 (N_22980,N_22730,N_22644);
and U22981 (N_22981,N_22578,N_22627);
xor U22982 (N_22982,N_22506,N_22618);
nor U22983 (N_22983,N_22587,N_22791);
nor U22984 (N_22984,N_22649,N_22517);
and U22985 (N_22985,N_22606,N_22507);
xor U22986 (N_22986,N_22521,N_22684);
xnor U22987 (N_22987,N_22595,N_22611);
and U22988 (N_22988,N_22550,N_22798);
or U22989 (N_22989,N_22639,N_22759);
or U22990 (N_22990,N_22797,N_22571);
nor U22991 (N_22991,N_22599,N_22598);
and U22992 (N_22992,N_22584,N_22509);
or U22993 (N_22993,N_22614,N_22764);
or U22994 (N_22994,N_22776,N_22696);
or U22995 (N_22995,N_22571,N_22607);
nor U22996 (N_22996,N_22772,N_22661);
or U22997 (N_22997,N_22505,N_22681);
xnor U22998 (N_22998,N_22627,N_22539);
and U22999 (N_22999,N_22718,N_22750);
nand U23000 (N_23000,N_22772,N_22627);
nand U23001 (N_23001,N_22720,N_22789);
xnor U23002 (N_23002,N_22585,N_22633);
nor U23003 (N_23003,N_22558,N_22753);
or U23004 (N_23004,N_22570,N_22771);
xor U23005 (N_23005,N_22614,N_22684);
nor U23006 (N_23006,N_22662,N_22742);
nand U23007 (N_23007,N_22683,N_22779);
nor U23008 (N_23008,N_22660,N_22576);
nor U23009 (N_23009,N_22507,N_22661);
nor U23010 (N_23010,N_22797,N_22705);
or U23011 (N_23011,N_22783,N_22540);
nand U23012 (N_23012,N_22741,N_22575);
xor U23013 (N_23013,N_22620,N_22711);
and U23014 (N_23014,N_22670,N_22797);
xnor U23015 (N_23015,N_22651,N_22701);
and U23016 (N_23016,N_22574,N_22647);
xor U23017 (N_23017,N_22619,N_22647);
and U23018 (N_23018,N_22768,N_22650);
xor U23019 (N_23019,N_22701,N_22569);
and U23020 (N_23020,N_22558,N_22700);
and U23021 (N_23021,N_22711,N_22591);
nor U23022 (N_23022,N_22798,N_22547);
or U23023 (N_23023,N_22682,N_22513);
xnor U23024 (N_23024,N_22606,N_22677);
xnor U23025 (N_23025,N_22627,N_22702);
and U23026 (N_23026,N_22604,N_22634);
and U23027 (N_23027,N_22519,N_22585);
xnor U23028 (N_23028,N_22724,N_22779);
xor U23029 (N_23029,N_22782,N_22713);
nor U23030 (N_23030,N_22757,N_22754);
nand U23031 (N_23031,N_22554,N_22672);
nor U23032 (N_23032,N_22633,N_22564);
or U23033 (N_23033,N_22725,N_22682);
nand U23034 (N_23034,N_22526,N_22650);
and U23035 (N_23035,N_22760,N_22665);
xnor U23036 (N_23036,N_22740,N_22503);
and U23037 (N_23037,N_22711,N_22743);
xor U23038 (N_23038,N_22673,N_22648);
xnor U23039 (N_23039,N_22778,N_22693);
or U23040 (N_23040,N_22599,N_22762);
nand U23041 (N_23041,N_22631,N_22657);
nor U23042 (N_23042,N_22638,N_22707);
nand U23043 (N_23043,N_22656,N_22648);
and U23044 (N_23044,N_22500,N_22530);
or U23045 (N_23045,N_22571,N_22548);
xnor U23046 (N_23046,N_22564,N_22691);
nand U23047 (N_23047,N_22680,N_22514);
or U23048 (N_23048,N_22543,N_22635);
xor U23049 (N_23049,N_22541,N_22758);
nand U23050 (N_23050,N_22729,N_22641);
nand U23051 (N_23051,N_22599,N_22760);
or U23052 (N_23052,N_22504,N_22741);
nand U23053 (N_23053,N_22508,N_22588);
or U23054 (N_23054,N_22579,N_22770);
nor U23055 (N_23055,N_22782,N_22754);
nor U23056 (N_23056,N_22752,N_22709);
nand U23057 (N_23057,N_22677,N_22664);
and U23058 (N_23058,N_22535,N_22681);
or U23059 (N_23059,N_22661,N_22601);
and U23060 (N_23060,N_22586,N_22773);
nor U23061 (N_23061,N_22766,N_22642);
xnor U23062 (N_23062,N_22550,N_22735);
or U23063 (N_23063,N_22509,N_22529);
and U23064 (N_23064,N_22560,N_22519);
or U23065 (N_23065,N_22501,N_22640);
nor U23066 (N_23066,N_22561,N_22678);
xnor U23067 (N_23067,N_22724,N_22795);
xor U23068 (N_23068,N_22665,N_22581);
or U23069 (N_23069,N_22758,N_22664);
nor U23070 (N_23070,N_22781,N_22700);
and U23071 (N_23071,N_22629,N_22631);
or U23072 (N_23072,N_22502,N_22755);
xnor U23073 (N_23073,N_22743,N_22748);
nand U23074 (N_23074,N_22771,N_22573);
nor U23075 (N_23075,N_22536,N_22553);
nor U23076 (N_23076,N_22674,N_22772);
xor U23077 (N_23077,N_22760,N_22788);
nor U23078 (N_23078,N_22677,N_22635);
xnor U23079 (N_23079,N_22518,N_22658);
xor U23080 (N_23080,N_22659,N_22509);
and U23081 (N_23081,N_22710,N_22524);
and U23082 (N_23082,N_22546,N_22727);
or U23083 (N_23083,N_22741,N_22701);
xor U23084 (N_23084,N_22514,N_22533);
xnor U23085 (N_23085,N_22508,N_22580);
nand U23086 (N_23086,N_22514,N_22513);
xnor U23087 (N_23087,N_22797,N_22648);
xor U23088 (N_23088,N_22659,N_22580);
xor U23089 (N_23089,N_22712,N_22785);
nand U23090 (N_23090,N_22596,N_22664);
nor U23091 (N_23091,N_22796,N_22701);
and U23092 (N_23092,N_22763,N_22643);
or U23093 (N_23093,N_22642,N_22797);
nand U23094 (N_23094,N_22726,N_22514);
nor U23095 (N_23095,N_22712,N_22749);
nand U23096 (N_23096,N_22510,N_22772);
nand U23097 (N_23097,N_22705,N_22601);
or U23098 (N_23098,N_22601,N_22739);
xor U23099 (N_23099,N_22513,N_22763);
nand U23100 (N_23100,N_22903,N_23069);
and U23101 (N_23101,N_23037,N_22891);
xnor U23102 (N_23102,N_23033,N_22922);
nand U23103 (N_23103,N_22875,N_22999);
or U23104 (N_23104,N_22805,N_22950);
nor U23105 (N_23105,N_22898,N_22860);
and U23106 (N_23106,N_23035,N_22929);
nand U23107 (N_23107,N_22850,N_22863);
and U23108 (N_23108,N_23073,N_22956);
xor U23109 (N_23109,N_22995,N_23020);
nor U23110 (N_23110,N_22955,N_22815);
or U23111 (N_23111,N_23021,N_22983);
and U23112 (N_23112,N_23050,N_22902);
xor U23113 (N_23113,N_22952,N_23002);
xor U23114 (N_23114,N_23023,N_22835);
xnor U23115 (N_23115,N_23083,N_22967);
xor U23116 (N_23116,N_22817,N_22802);
or U23117 (N_23117,N_22871,N_22880);
and U23118 (N_23118,N_22866,N_23057);
nand U23119 (N_23119,N_22869,N_23026);
nand U23120 (N_23120,N_22960,N_22979);
and U23121 (N_23121,N_22978,N_23079);
and U23122 (N_23122,N_22966,N_22827);
nand U23123 (N_23123,N_22806,N_23067);
nor U23124 (N_23124,N_22857,N_23001);
nor U23125 (N_23125,N_23097,N_23095);
nand U23126 (N_23126,N_23015,N_22911);
or U23127 (N_23127,N_23017,N_22877);
or U23128 (N_23128,N_22941,N_23005);
nor U23129 (N_23129,N_22972,N_22804);
nor U23130 (N_23130,N_22887,N_23091);
or U23131 (N_23131,N_22836,N_22886);
xor U23132 (N_23132,N_22820,N_22907);
xnor U23133 (N_23133,N_23077,N_22818);
nand U23134 (N_23134,N_22948,N_23041);
and U23135 (N_23135,N_22816,N_23009);
and U23136 (N_23136,N_22964,N_22943);
nand U23137 (N_23137,N_23031,N_22923);
and U23138 (N_23138,N_23048,N_22984);
or U23139 (N_23139,N_23036,N_22969);
nand U23140 (N_23140,N_22930,N_23089);
or U23141 (N_23141,N_23051,N_22945);
nand U23142 (N_23142,N_23049,N_22993);
or U23143 (N_23143,N_22822,N_22914);
xnor U23144 (N_23144,N_22940,N_22883);
or U23145 (N_23145,N_22986,N_23000);
and U23146 (N_23146,N_22974,N_22897);
nor U23147 (N_23147,N_22894,N_23012);
and U23148 (N_23148,N_22991,N_22998);
and U23149 (N_23149,N_23082,N_23078);
nand U23150 (N_23150,N_22989,N_22918);
nor U23151 (N_23151,N_22992,N_22849);
and U23152 (N_23152,N_22946,N_22888);
and U23153 (N_23153,N_22878,N_22977);
or U23154 (N_23154,N_22884,N_22861);
nand U23155 (N_23155,N_23081,N_23003);
nor U23156 (N_23156,N_22890,N_22963);
or U23157 (N_23157,N_23008,N_22851);
and U23158 (N_23158,N_22821,N_22809);
xnor U23159 (N_23159,N_22812,N_22811);
nand U23160 (N_23160,N_22831,N_23004);
and U23161 (N_23161,N_22900,N_22959);
and U23162 (N_23162,N_22868,N_23094);
or U23163 (N_23163,N_23087,N_22926);
nand U23164 (N_23164,N_22833,N_22919);
or U23165 (N_23165,N_23063,N_22932);
nor U23166 (N_23166,N_22867,N_23076);
nand U23167 (N_23167,N_22909,N_22843);
nor U23168 (N_23168,N_22913,N_23090);
and U23169 (N_23169,N_23092,N_23075);
nor U23170 (N_23170,N_23028,N_22904);
xor U23171 (N_23171,N_22881,N_23086);
nand U23172 (N_23172,N_23060,N_23061);
nand U23173 (N_23173,N_22801,N_22874);
or U23174 (N_23174,N_22864,N_23053);
nor U23175 (N_23175,N_22813,N_22839);
and U23176 (N_23176,N_22858,N_23047);
or U23177 (N_23177,N_23093,N_22824);
nor U23178 (N_23178,N_23016,N_23024);
or U23179 (N_23179,N_22934,N_22954);
or U23180 (N_23180,N_22915,N_22971);
nand U23181 (N_23181,N_23052,N_23022);
xnor U23182 (N_23182,N_23039,N_23088);
or U23183 (N_23183,N_22828,N_22951);
or U23184 (N_23184,N_22896,N_22873);
and U23185 (N_23185,N_23072,N_22845);
nor U23186 (N_23186,N_22825,N_22865);
nor U23187 (N_23187,N_22924,N_22962);
nand U23188 (N_23188,N_22917,N_22834);
nand U23189 (N_23189,N_23014,N_22856);
nor U23190 (N_23190,N_22800,N_22910);
and U23191 (N_23191,N_22852,N_23068);
or U23192 (N_23192,N_22838,N_23084);
nand U23193 (N_23193,N_22997,N_23058);
or U23194 (N_23194,N_23025,N_22939);
or U23195 (N_23195,N_22958,N_22942);
or U23196 (N_23196,N_22899,N_22920);
and U23197 (N_23197,N_22925,N_23040);
and U23198 (N_23198,N_22933,N_23027);
nor U23199 (N_23199,N_22814,N_22837);
xnor U23200 (N_23200,N_22844,N_22981);
nor U23201 (N_23201,N_22807,N_22853);
nand U23202 (N_23202,N_22990,N_23018);
and U23203 (N_23203,N_23045,N_22882);
or U23204 (N_23204,N_23007,N_23034);
xnor U23205 (N_23205,N_22808,N_22935);
nor U23206 (N_23206,N_23030,N_22889);
nand U23207 (N_23207,N_22829,N_22872);
nor U23208 (N_23208,N_22803,N_23046);
and U23209 (N_23209,N_23013,N_22819);
nor U23210 (N_23210,N_23042,N_22975);
or U23211 (N_23211,N_22988,N_23019);
xor U23212 (N_23212,N_23099,N_22893);
nor U23213 (N_23213,N_23043,N_22876);
xnor U23214 (N_23214,N_22859,N_23032);
nand U23215 (N_23215,N_22879,N_22862);
xor U23216 (N_23216,N_22996,N_22987);
nor U23217 (N_23217,N_22840,N_22976);
or U23218 (N_23218,N_23070,N_22846);
nor U23219 (N_23219,N_22994,N_22927);
xnor U23220 (N_23220,N_22944,N_22854);
and U23221 (N_23221,N_23062,N_22830);
and U23222 (N_23222,N_22985,N_23098);
xnor U23223 (N_23223,N_22982,N_23059);
nor U23224 (N_23224,N_22855,N_22892);
or U23225 (N_23225,N_22823,N_22965);
nand U23226 (N_23226,N_22947,N_23044);
and U23227 (N_23227,N_23038,N_22905);
nor U23228 (N_23228,N_22848,N_22949);
nand U23229 (N_23229,N_22870,N_22847);
nand U23230 (N_23230,N_23054,N_23065);
and U23231 (N_23231,N_22980,N_22937);
nor U23232 (N_23232,N_22936,N_23056);
nor U23233 (N_23233,N_22906,N_22885);
xnor U23234 (N_23234,N_23080,N_23085);
nand U23235 (N_23235,N_22973,N_22895);
and U23236 (N_23236,N_22961,N_22938);
or U23237 (N_23237,N_22928,N_22968);
nor U23238 (N_23238,N_23096,N_22832);
xnor U23239 (N_23239,N_22931,N_23066);
nand U23240 (N_23240,N_23055,N_23006);
or U23241 (N_23241,N_22953,N_22916);
nor U23242 (N_23242,N_22841,N_23011);
nor U23243 (N_23243,N_22957,N_23074);
nor U23244 (N_23244,N_23064,N_23010);
and U23245 (N_23245,N_23029,N_22842);
and U23246 (N_23246,N_22810,N_23071);
xnor U23247 (N_23247,N_22912,N_22921);
nor U23248 (N_23248,N_22901,N_22908);
nor U23249 (N_23249,N_22970,N_22826);
xor U23250 (N_23250,N_23090,N_22840);
or U23251 (N_23251,N_23039,N_22887);
and U23252 (N_23252,N_23093,N_22936);
nor U23253 (N_23253,N_22911,N_23097);
or U23254 (N_23254,N_23077,N_23048);
nor U23255 (N_23255,N_22881,N_22910);
nand U23256 (N_23256,N_22888,N_22953);
or U23257 (N_23257,N_22969,N_22842);
nand U23258 (N_23258,N_23041,N_22955);
xor U23259 (N_23259,N_22928,N_22988);
or U23260 (N_23260,N_22854,N_23051);
and U23261 (N_23261,N_23063,N_22926);
nor U23262 (N_23262,N_23005,N_23065);
or U23263 (N_23263,N_23007,N_22816);
xor U23264 (N_23264,N_22867,N_22938);
nor U23265 (N_23265,N_22954,N_22961);
or U23266 (N_23266,N_23090,N_22855);
xnor U23267 (N_23267,N_23046,N_22900);
xor U23268 (N_23268,N_22987,N_22804);
xnor U23269 (N_23269,N_23031,N_22851);
and U23270 (N_23270,N_23072,N_22802);
nor U23271 (N_23271,N_22829,N_22898);
or U23272 (N_23272,N_23036,N_22818);
and U23273 (N_23273,N_22822,N_22883);
xnor U23274 (N_23274,N_23055,N_23053);
nor U23275 (N_23275,N_23006,N_23005);
nand U23276 (N_23276,N_22975,N_23073);
xnor U23277 (N_23277,N_22946,N_23061);
and U23278 (N_23278,N_22910,N_22920);
xor U23279 (N_23279,N_22861,N_22834);
nor U23280 (N_23280,N_22912,N_23000);
xor U23281 (N_23281,N_22910,N_23021);
and U23282 (N_23282,N_23000,N_22879);
nand U23283 (N_23283,N_22820,N_22964);
and U23284 (N_23284,N_23037,N_22812);
nand U23285 (N_23285,N_22837,N_22924);
nand U23286 (N_23286,N_22875,N_22813);
and U23287 (N_23287,N_22958,N_22945);
or U23288 (N_23288,N_22813,N_22838);
xor U23289 (N_23289,N_22992,N_22848);
or U23290 (N_23290,N_23023,N_23039);
or U23291 (N_23291,N_22969,N_22957);
and U23292 (N_23292,N_22967,N_22813);
or U23293 (N_23293,N_23069,N_22888);
nor U23294 (N_23294,N_22936,N_23004);
xor U23295 (N_23295,N_22802,N_22895);
and U23296 (N_23296,N_23065,N_22988);
or U23297 (N_23297,N_22911,N_23031);
nand U23298 (N_23298,N_22818,N_22996);
and U23299 (N_23299,N_22885,N_22913);
or U23300 (N_23300,N_23042,N_23061);
and U23301 (N_23301,N_23010,N_22887);
xnor U23302 (N_23302,N_23063,N_22985);
and U23303 (N_23303,N_23008,N_23032);
and U23304 (N_23304,N_23082,N_23087);
xnor U23305 (N_23305,N_23044,N_22960);
nor U23306 (N_23306,N_22879,N_23022);
or U23307 (N_23307,N_22806,N_22810);
nor U23308 (N_23308,N_22817,N_22967);
xor U23309 (N_23309,N_22827,N_22971);
and U23310 (N_23310,N_23059,N_22905);
nand U23311 (N_23311,N_22934,N_23035);
and U23312 (N_23312,N_22962,N_22810);
or U23313 (N_23313,N_23078,N_22903);
xor U23314 (N_23314,N_22962,N_22974);
nand U23315 (N_23315,N_22827,N_22884);
xor U23316 (N_23316,N_23090,N_22864);
nor U23317 (N_23317,N_22907,N_23042);
xnor U23318 (N_23318,N_23090,N_22809);
nor U23319 (N_23319,N_23040,N_22828);
and U23320 (N_23320,N_23061,N_22950);
xor U23321 (N_23321,N_23065,N_22940);
and U23322 (N_23322,N_23040,N_22827);
and U23323 (N_23323,N_22808,N_22933);
and U23324 (N_23324,N_22874,N_22867);
nand U23325 (N_23325,N_23085,N_23054);
or U23326 (N_23326,N_22944,N_22997);
nand U23327 (N_23327,N_23051,N_22915);
or U23328 (N_23328,N_22822,N_22918);
or U23329 (N_23329,N_23087,N_22813);
nor U23330 (N_23330,N_22879,N_23092);
and U23331 (N_23331,N_23048,N_22840);
or U23332 (N_23332,N_22979,N_22931);
nand U23333 (N_23333,N_22916,N_22850);
nand U23334 (N_23334,N_22865,N_22883);
nor U23335 (N_23335,N_22845,N_23093);
nand U23336 (N_23336,N_22966,N_22811);
nand U23337 (N_23337,N_23018,N_22946);
or U23338 (N_23338,N_23009,N_22991);
nand U23339 (N_23339,N_22910,N_22803);
nor U23340 (N_23340,N_23049,N_23008);
nand U23341 (N_23341,N_22902,N_23020);
xor U23342 (N_23342,N_22819,N_22923);
xnor U23343 (N_23343,N_22928,N_22957);
nand U23344 (N_23344,N_22976,N_23084);
or U23345 (N_23345,N_22802,N_22844);
nand U23346 (N_23346,N_22970,N_22991);
and U23347 (N_23347,N_22968,N_22897);
nand U23348 (N_23348,N_22810,N_22871);
nand U23349 (N_23349,N_22918,N_22867);
or U23350 (N_23350,N_23019,N_22895);
xor U23351 (N_23351,N_22853,N_22979);
xor U23352 (N_23352,N_22984,N_22829);
or U23353 (N_23353,N_22957,N_22812);
nor U23354 (N_23354,N_23033,N_23068);
nand U23355 (N_23355,N_23000,N_22825);
or U23356 (N_23356,N_23012,N_22980);
or U23357 (N_23357,N_22846,N_23031);
nor U23358 (N_23358,N_22947,N_22892);
nand U23359 (N_23359,N_22963,N_23021);
nor U23360 (N_23360,N_22965,N_22974);
xor U23361 (N_23361,N_23059,N_22825);
or U23362 (N_23362,N_22986,N_22928);
or U23363 (N_23363,N_22974,N_22925);
or U23364 (N_23364,N_22877,N_22915);
xnor U23365 (N_23365,N_22897,N_22827);
nor U23366 (N_23366,N_22883,N_22948);
xor U23367 (N_23367,N_22807,N_22827);
or U23368 (N_23368,N_22954,N_22814);
nand U23369 (N_23369,N_22961,N_23037);
xor U23370 (N_23370,N_23004,N_23060);
and U23371 (N_23371,N_22886,N_22831);
nor U23372 (N_23372,N_23052,N_22883);
and U23373 (N_23373,N_22975,N_22835);
nand U23374 (N_23374,N_22973,N_23095);
nand U23375 (N_23375,N_22866,N_23005);
xor U23376 (N_23376,N_22943,N_22939);
or U23377 (N_23377,N_22851,N_22819);
nor U23378 (N_23378,N_22971,N_23057);
nor U23379 (N_23379,N_22947,N_22911);
or U23380 (N_23380,N_22854,N_22911);
xor U23381 (N_23381,N_22982,N_23034);
nand U23382 (N_23382,N_22935,N_23048);
or U23383 (N_23383,N_23031,N_22944);
and U23384 (N_23384,N_23089,N_22890);
nand U23385 (N_23385,N_22825,N_23064);
or U23386 (N_23386,N_23034,N_22983);
nor U23387 (N_23387,N_23026,N_23092);
or U23388 (N_23388,N_22806,N_22861);
nor U23389 (N_23389,N_22802,N_22906);
or U23390 (N_23390,N_22877,N_23088);
and U23391 (N_23391,N_22841,N_22989);
xnor U23392 (N_23392,N_22891,N_22882);
xor U23393 (N_23393,N_22811,N_22945);
or U23394 (N_23394,N_22904,N_22976);
nand U23395 (N_23395,N_22881,N_22955);
or U23396 (N_23396,N_23095,N_22956);
and U23397 (N_23397,N_22824,N_22977);
nand U23398 (N_23398,N_22872,N_22936);
or U23399 (N_23399,N_22996,N_22978);
or U23400 (N_23400,N_23329,N_23284);
nor U23401 (N_23401,N_23190,N_23232);
and U23402 (N_23402,N_23230,N_23367);
or U23403 (N_23403,N_23368,N_23266);
xor U23404 (N_23404,N_23293,N_23122);
or U23405 (N_23405,N_23247,N_23208);
nor U23406 (N_23406,N_23352,N_23276);
or U23407 (N_23407,N_23181,N_23334);
nand U23408 (N_23408,N_23177,N_23186);
or U23409 (N_23409,N_23174,N_23298);
nor U23410 (N_23410,N_23264,N_23341);
xor U23411 (N_23411,N_23254,N_23219);
or U23412 (N_23412,N_23101,N_23176);
xor U23413 (N_23413,N_23178,N_23320);
nand U23414 (N_23414,N_23381,N_23103);
or U23415 (N_23415,N_23241,N_23288);
xnor U23416 (N_23416,N_23185,N_23315);
xnor U23417 (N_23417,N_23119,N_23326);
nand U23418 (N_23418,N_23160,N_23244);
or U23419 (N_23419,N_23162,N_23117);
xnor U23420 (N_23420,N_23283,N_23307);
and U23421 (N_23421,N_23205,N_23248);
nand U23422 (N_23422,N_23173,N_23280);
and U23423 (N_23423,N_23379,N_23384);
or U23424 (N_23424,N_23207,N_23359);
xor U23425 (N_23425,N_23339,N_23242);
nand U23426 (N_23426,N_23279,N_23191);
and U23427 (N_23427,N_23135,N_23277);
or U23428 (N_23428,N_23378,N_23150);
nor U23429 (N_23429,N_23209,N_23121);
nand U23430 (N_23430,N_23151,N_23102);
or U23431 (N_23431,N_23202,N_23172);
or U23432 (N_23432,N_23217,N_23371);
and U23433 (N_23433,N_23147,N_23170);
nor U23434 (N_23434,N_23336,N_23218);
nand U23435 (N_23435,N_23356,N_23155);
or U23436 (N_23436,N_23297,N_23164);
nand U23437 (N_23437,N_23152,N_23364);
nor U23438 (N_23438,N_23107,N_23196);
nand U23439 (N_23439,N_23259,N_23304);
and U23440 (N_23440,N_23385,N_23161);
nor U23441 (N_23441,N_23255,N_23233);
and U23442 (N_23442,N_23245,N_23347);
nand U23443 (N_23443,N_23204,N_23260);
and U23444 (N_23444,N_23194,N_23169);
nand U23445 (N_23445,N_23372,N_23394);
and U23446 (N_23446,N_23136,N_23396);
and U23447 (N_23447,N_23370,N_23183);
nand U23448 (N_23448,N_23104,N_23335);
or U23449 (N_23449,N_23234,N_23321);
nand U23450 (N_23450,N_23295,N_23322);
and U23451 (N_23451,N_23327,N_23148);
or U23452 (N_23452,N_23342,N_23109);
or U23453 (N_23453,N_23210,N_23100);
nor U23454 (N_23454,N_23224,N_23332);
or U23455 (N_23455,N_23115,N_23249);
or U23456 (N_23456,N_23363,N_23392);
or U23457 (N_23457,N_23262,N_23299);
xor U23458 (N_23458,N_23243,N_23310);
nor U23459 (N_23459,N_23200,N_23128);
nand U23460 (N_23460,N_23362,N_23201);
or U23461 (N_23461,N_23383,N_23361);
or U23462 (N_23462,N_23349,N_23149);
nand U23463 (N_23463,N_23134,N_23229);
xor U23464 (N_23464,N_23206,N_23132);
xor U23465 (N_23465,N_23274,N_23153);
and U23466 (N_23466,N_23373,N_23388);
xor U23467 (N_23467,N_23195,N_23308);
nand U23468 (N_23468,N_23222,N_23171);
or U23469 (N_23469,N_23389,N_23289);
nand U23470 (N_23470,N_23272,N_23351);
or U23471 (N_23471,N_23286,N_23225);
xnor U23472 (N_23472,N_23330,N_23125);
and U23473 (N_23473,N_23211,N_23301);
nand U23474 (N_23474,N_23126,N_23246);
and U23475 (N_23475,N_23138,N_23139);
and U23476 (N_23476,N_23393,N_23311);
and U23477 (N_23477,N_23313,N_23358);
or U23478 (N_23478,N_23236,N_23131);
xnor U23479 (N_23479,N_23380,N_23340);
xor U23480 (N_23480,N_23346,N_23338);
and U23481 (N_23481,N_23157,N_23158);
nand U23482 (N_23482,N_23213,N_23220);
or U23483 (N_23483,N_23319,N_23163);
or U23484 (N_23484,N_23268,N_23116);
nand U23485 (N_23485,N_23110,N_23198);
nor U23486 (N_23486,N_23386,N_23300);
and U23487 (N_23487,N_23221,N_23154);
or U23488 (N_23488,N_23325,N_23285);
or U23489 (N_23489,N_23303,N_23273);
nor U23490 (N_23490,N_23212,N_23318);
xnor U23491 (N_23491,N_23261,N_23124);
and U23492 (N_23492,N_23253,N_23267);
or U23493 (N_23493,N_23193,N_23216);
nor U23494 (N_23494,N_23294,N_23187);
nand U23495 (N_23495,N_23398,N_23108);
or U23496 (N_23496,N_23270,N_23395);
or U23497 (N_23497,N_23214,N_23203);
nor U23498 (N_23498,N_23156,N_23146);
xnor U23499 (N_23499,N_23377,N_23328);
nand U23500 (N_23500,N_23235,N_23348);
or U23501 (N_23501,N_23112,N_23227);
nor U23502 (N_23502,N_23312,N_23281);
or U23503 (N_23503,N_23344,N_23114);
nor U23504 (N_23504,N_23337,N_23137);
xor U23505 (N_23505,N_23179,N_23106);
nor U23506 (N_23506,N_23275,N_23350);
nor U23507 (N_23507,N_23166,N_23240);
nor U23508 (N_23508,N_23357,N_23366);
or U23509 (N_23509,N_23111,N_23228);
xor U23510 (N_23510,N_23355,N_23399);
or U23511 (N_23511,N_23159,N_23215);
xor U23512 (N_23512,N_23323,N_23353);
nand U23513 (N_23513,N_23309,N_23271);
and U23514 (N_23514,N_23113,N_23127);
nand U23515 (N_23515,N_23291,N_23197);
xnor U23516 (N_23516,N_23316,N_23129);
xnor U23517 (N_23517,N_23278,N_23369);
xnor U23518 (N_23518,N_23123,N_23302);
nor U23519 (N_23519,N_23331,N_23250);
nand U23520 (N_23520,N_23292,N_23251);
xor U23521 (N_23521,N_23182,N_23118);
and U23522 (N_23522,N_23333,N_23226);
nor U23523 (N_23523,N_23391,N_23189);
and U23524 (N_23524,N_23237,N_23144);
xor U23525 (N_23525,N_23263,N_23376);
nand U23526 (N_23526,N_23343,N_23296);
nand U23527 (N_23527,N_23175,N_23238);
nor U23528 (N_23528,N_23239,N_23375);
and U23529 (N_23529,N_23165,N_23305);
nand U23530 (N_23530,N_23390,N_23354);
nor U23531 (N_23531,N_23252,N_23143);
nor U23532 (N_23532,N_23282,N_23192);
xor U23533 (N_23533,N_23167,N_23133);
or U23534 (N_23534,N_23120,N_23374);
and U23535 (N_23535,N_23314,N_23324);
nand U23536 (N_23536,N_23269,N_23256);
and U23537 (N_23537,N_23141,N_23360);
or U23538 (N_23538,N_23142,N_23317);
nor U23539 (N_23539,N_23180,N_23257);
nand U23540 (N_23540,N_23105,N_23231);
nand U23541 (N_23541,N_23130,N_23223);
nand U23542 (N_23542,N_23265,N_23397);
or U23543 (N_23543,N_23365,N_23145);
xor U23544 (N_23544,N_23168,N_23382);
nor U23545 (N_23545,N_23258,N_23387);
xor U23546 (N_23546,N_23188,N_23290);
and U23547 (N_23547,N_23140,N_23306);
or U23548 (N_23548,N_23287,N_23199);
and U23549 (N_23549,N_23345,N_23184);
or U23550 (N_23550,N_23236,N_23285);
nor U23551 (N_23551,N_23323,N_23176);
nand U23552 (N_23552,N_23324,N_23139);
nor U23553 (N_23553,N_23102,N_23338);
xor U23554 (N_23554,N_23339,N_23381);
nor U23555 (N_23555,N_23261,N_23151);
and U23556 (N_23556,N_23322,N_23381);
nor U23557 (N_23557,N_23285,N_23346);
or U23558 (N_23558,N_23178,N_23328);
nor U23559 (N_23559,N_23247,N_23314);
xnor U23560 (N_23560,N_23332,N_23166);
and U23561 (N_23561,N_23110,N_23341);
or U23562 (N_23562,N_23195,N_23365);
and U23563 (N_23563,N_23377,N_23252);
or U23564 (N_23564,N_23120,N_23203);
xnor U23565 (N_23565,N_23399,N_23152);
nor U23566 (N_23566,N_23140,N_23189);
nor U23567 (N_23567,N_23135,N_23148);
and U23568 (N_23568,N_23196,N_23187);
and U23569 (N_23569,N_23257,N_23243);
or U23570 (N_23570,N_23200,N_23201);
xnor U23571 (N_23571,N_23103,N_23158);
nand U23572 (N_23572,N_23179,N_23184);
xnor U23573 (N_23573,N_23327,N_23254);
or U23574 (N_23574,N_23375,N_23115);
xnor U23575 (N_23575,N_23384,N_23232);
nor U23576 (N_23576,N_23278,N_23207);
and U23577 (N_23577,N_23179,N_23109);
nand U23578 (N_23578,N_23221,N_23284);
xor U23579 (N_23579,N_23274,N_23176);
xnor U23580 (N_23580,N_23375,N_23303);
nand U23581 (N_23581,N_23287,N_23309);
nor U23582 (N_23582,N_23335,N_23216);
nand U23583 (N_23583,N_23101,N_23378);
nand U23584 (N_23584,N_23235,N_23369);
xnor U23585 (N_23585,N_23268,N_23216);
or U23586 (N_23586,N_23301,N_23186);
nor U23587 (N_23587,N_23361,N_23121);
xnor U23588 (N_23588,N_23380,N_23320);
nor U23589 (N_23589,N_23361,N_23313);
nor U23590 (N_23590,N_23194,N_23148);
nor U23591 (N_23591,N_23363,N_23186);
nand U23592 (N_23592,N_23399,N_23339);
or U23593 (N_23593,N_23368,N_23329);
nand U23594 (N_23594,N_23106,N_23383);
or U23595 (N_23595,N_23223,N_23238);
xor U23596 (N_23596,N_23353,N_23280);
xnor U23597 (N_23597,N_23380,N_23177);
and U23598 (N_23598,N_23268,N_23237);
and U23599 (N_23599,N_23341,N_23167);
and U23600 (N_23600,N_23155,N_23115);
xor U23601 (N_23601,N_23322,N_23168);
nand U23602 (N_23602,N_23198,N_23252);
and U23603 (N_23603,N_23173,N_23197);
xnor U23604 (N_23604,N_23184,N_23172);
or U23605 (N_23605,N_23250,N_23337);
and U23606 (N_23606,N_23317,N_23347);
xnor U23607 (N_23607,N_23327,N_23265);
xor U23608 (N_23608,N_23315,N_23241);
or U23609 (N_23609,N_23127,N_23391);
or U23610 (N_23610,N_23285,N_23349);
nor U23611 (N_23611,N_23361,N_23315);
xnor U23612 (N_23612,N_23224,N_23352);
nand U23613 (N_23613,N_23190,N_23259);
nand U23614 (N_23614,N_23240,N_23296);
or U23615 (N_23615,N_23158,N_23194);
nor U23616 (N_23616,N_23171,N_23177);
nand U23617 (N_23617,N_23355,N_23214);
nor U23618 (N_23618,N_23151,N_23291);
xor U23619 (N_23619,N_23242,N_23353);
xor U23620 (N_23620,N_23188,N_23201);
nor U23621 (N_23621,N_23378,N_23256);
xor U23622 (N_23622,N_23102,N_23286);
xor U23623 (N_23623,N_23144,N_23142);
and U23624 (N_23624,N_23338,N_23127);
or U23625 (N_23625,N_23309,N_23150);
and U23626 (N_23626,N_23276,N_23120);
xnor U23627 (N_23627,N_23145,N_23217);
or U23628 (N_23628,N_23376,N_23125);
xor U23629 (N_23629,N_23396,N_23370);
and U23630 (N_23630,N_23252,N_23177);
and U23631 (N_23631,N_23173,N_23269);
and U23632 (N_23632,N_23316,N_23190);
or U23633 (N_23633,N_23340,N_23374);
and U23634 (N_23634,N_23134,N_23120);
xor U23635 (N_23635,N_23359,N_23234);
or U23636 (N_23636,N_23197,N_23375);
nand U23637 (N_23637,N_23277,N_23262);
nand U23638 (N_23638,N_23260,N_23280);
xnor U23639 (N_23639,N_23388,N_23164);
nand U23640 (N_23640,N_23265,N_23264);
nand U23641 (N_23641,N_23127,N_23200);
and U23642 (N_23642,N_23250,N_23349);
xnor U23643 (N_23643,N_23290,N_23147);
and U23644 (N_23644,N_23393,N_23277);
xor U23645 (N_23645,N_23185,N_23302);
nand U23646 (N_23646,N_23357,N_23116);
or U23647 (N_23647,N_23247,N_23375);
nand U23648 (N_23648,N_23363,N_23252);
and U23649 (N_23649,N_23252,N_23294);
xnor U23650 (N_23650,N_23391,N_23209);
and U23651 (N_23651,N_23388,N_23285);
or U23652 (N_23652,N_23353,N_23287);
nor U23653 (N_23653,N_23308,N_23282);
nand U23654 (N_23654,N_23320,N_23399);
and U23655 (N_23655,N_23332,N_23168);
or U23656 (N_23656,N_23334,N_23309);
nor U23657 (N_23657,N_23382,N_23361);
or U23658 (N_23658,N_23339,N_23201);
and U23659 (N_23659,N_23390,N_23158);
xor U23660 (N_23660,N_23278,N_23212);
or U23661 (N_23661,N_23198,N_23171);
and U23662 (N_23662,N_23318,N_23242);
or U23663 (N_23663,N_23234,N_23328);
xor U23664 (N_23664,N_23382,N_23267);
nand U23665 (N_23665,N_23326,N_23168);
nand U23666 (N_23666,N_23268,N_23395);
and U23667 (N_23667,N_23194,N_23196);
and U23668 (N_23668,N_23313,N_23246);
xor U23669 (N_23669,N_23347,N_23188);
xnor U23670 (N_23670,N_23173,N_23393);
nand U23671 (N_23671,N_23376,N_23149);
or U23672 (N_23672,N_23287,N_23182);
and U23673 (N_23673,N_23274,N_23123);
and U23674 (N_23674,N_23117,N_23327);
xor U23675 (N_23675,N_23297,N_23221);
nand U23676 (N_23676,N_23127,N_23399);
nor U23677 (N_23677,N_23295,N_23245);
nand U23678 (N_23678,N_23305,N_23106);
and U23679 (N_23679,N_23186,N_23283);
nand U23680 (N_23680,N_23192,N_23161);
nor U23681 (N_23681,N_23175,N_23283);
and U23682 (N_23682,N_23222,N_23218);
and U23683 (N_23683,N_23283,N_23342);
nand U23684 (N_23684,N_23278,N_23224);
xor U23685 (N_23685,N_23160,N_23203);
nand U23686 (N_23686,N_23133,N_23163);
or U23687 (N_23687,N_23399,N_23380);
or U23688 (N_23688,N_23215,N_23338);
nor U23689 (N_23689,N_23122,N_23287);
xnor U23690 (N_23690,N_23311,N_23394);
nand U23691 (N_23691,N_23314,N_23329);
or U23692 (N_23692,N_23350,N_23221);
and U23693 (N_23693,N_23333,N_23216);
or U23694 (N_23694,N_23244,N_23190);
xnor U23695 (N_23695,N_23190,N_23182);
xnor U23696 (N_23696,N_23194,N_23352);
and U23697 (N_23697,N_23369,N_23331);
xor U23698 (N_23698,N_23245,N_23133);
or U23699 (N_23699,N_23260,N_23347);
xnor U23700 (N_23700,N_23536,N_23522);
and U23701 (N_23701,N_23681,N_23544);
nor U23702 (N_23702,N_23644,N_23577);
nand U23703 (N_23703,N_23525,N_23584);
and U23704 (N_23704,N_23563,N_23501);
nor U23705 (N_23705,N_23404,N_23573);
xor U23706 (N_23706,N_23658,N_23618);
nand U23707 (N_23707,N_23461,N_23580);
xnor U23708 (N_23708,N_23492,N_23433);
or U23709 (N_23709,N_23636,N_23490);
xor U23710 (N_23710,N_23402,N_23635);
or U23711 (N_23711,N_23499,N_23669);
and U23712 (N_23712,N_23534,N_23429);
xor U23713 (N_23713,N_23532,N_23460);
xnor U23714 (N_23714,N_23511,N_23673);
nand U23715 (N_23715,N_23697,N_23611);
xor U23716 (N_23716,N_23470,N_23489);
and U23717 (N_23717,N_23675,N_23473);
xnor U23718 (N_23718,N_23684,N_23406);
or U23719 (N_23719,N_23463,N_23449);
nand U23720 (N_23720,N_23556,N_23453);
and U23721 (N_23721,N_23459,N_23469);
or U23722 (N_23722,N_23553,N_23477);
nand U23723 (N_23723,N_23615,N_23550);
or U23724 (N_23724,N_23543,N_23627);
nand U23725 (N_23725,N_23415,N_23476);
and U23726 (N_23726,N_23509,N_23652);
xnor U23727 (N_23727,N_23515,N_23457);
nand U23728 (N_23728,N_23612,N_23602);
or U23729 (N_23729,N_23554,N_23596);
nor U23730 (N_23730,N_23471,N_23408);
xor U23731 (N_23731,N_23436,N_23451);
nor U23732 (N_23732,N_23467,N_23437);
and U23733 (N_23733,N_23672,N_23628);
or U23734 (N_23734,N_23416,N_23533);
xnor U23735 (N_23735,N_23633,N_23486);
and U23736 (N_23736,N_23680,N_23606);
or U23737 (N_23737,N_23514,N_23592);
or U23738 (N_23738,N_23435,N_23425);
nor U23739 (N_23739,N_23480,N_23495);
and U23740 (N_23740,N_23447,N_23430);
or U23741 (N_23741,N_23518,N_23665);
nor U23742 (N_23742,N_23696,N_23616);
and U23743 (N_23743,N_23448,N_23693);
or U23744 (N_23744,N_23513,N_23656);
xor U23745 (N_23745,N_23411,N_23421);
xnor U23746 (N_23746,N_23605,N_23657);
and U23747 (N_23747,N_23601,N_23519);
or U23748 (N_23748,N_23527,N_23564);
or U23749 (N_23749,N_23438,N_23503);
and U23750 (N_23750,N_23427,N_23566);
or U23751 (N_23751,N_23547,N_23642);
and U23752 (N_23752,N_23502,N_23688);
or U23753 (N_23753,N_23649,N_23560);
or U23754 (N_23754,N_23524,N_23428);
xor U23755 (N_23755,N_23588,N_23569);
or U23756 (N_23756,N_23521,N_23494);
nand U23757 (N_23757,N_23426,N_23419);
or U23758 (N_23758,N_23455,N_23695);
nor U23759 (N_23759,N_23510,N_23660);
xor U23760 (N_23760,N_23674,N_23617);
nand U23761 (N_23761,N_23487,N_23526);
nor U23762 (N_23762,N_23557,N_23529);
xor U23763 (N_23763,N_23434,N_23497);
and U23764 (N_23764,N_23456,N_23450);
or U23765 (N_23765,N_23661,N_23587);
or U23766 (N_23766,N_23694,N_23539);
and U23767 (N_23767,N_23454,N_23632);
and U23768 (N_23768,N_23662,N_23488);
and U23769 (N_23769,N_23578,N_23698);
nor U23770 (N_23770,N_23639,N_23679);
nor U23771 (N_23771,N_23687,N_23599);
or U23772 (N_23772,N_23498,N_23608);
and U23773 (N_23773,N_23496,N_23574);
and U23774 (N_23774,N_23607,N_23548);
nor U23775 (N_23775,N_23481,N_23439);
nor U23776 (N_23776,N_23546,N_23555);
nor U23777 (N_23777,N_23572,N_23655);
nand U23778 (N_23778,N_23575,N_23619);
xnor U23779 (N_23779,N_23666,N_23541);
or U23780 (N_23780,N_23683,N_23598);
xnor U23781 (N_23781,N_23603,N_23690);
or U23782 (N_23782,N_23646,N_23508);
and U23783 (N_23783,N_23412,N_23462);
xnor U23784 (N_23784,N_23631,N_23610);
and U23785 (N_23785,N_23540,N_23422);
xnor U23786 (N_23786,N_23483,N_23582);
or U23787 (N_23787,N_23468,N_23484);
xor U23788 (N_23788,N_23401,N_23663);
nand U23789 (N_23789,N_23620,N_23609);
xor U23790 (N_23790,N_23600,N_23579);
nor U23791 (N_23791,N_23651,N_23441);
nand U23792 (N_23792,N_23593,N_23668);
nand U23793 (N_23793,N_23581,N_23670);
nor U23794 (N_23794,N_23559,N_23407);
or U23795 (N_23795,N_23570,N_23400);
nand U23796 (N_23796,N_23645,N_23640);
or U23797 (N_23797,N_23568,N_23589);
or U23798 (N_23798,N_23423,N_23659);
xnor U23799 (N_23799,N_23590,N_23478);
and U23800 (N_23800,N_23637,N_23479);
nor U23801 (N_23801,N_23594,N_23552);
nor U23802 (N_23802,N_23613,N_23561);
nand U23803 (N_23803,N_23597,N_23586);
nand U23804 (N_23804,N_23537,N_23623);
xnor U23805 (N_23805,N_23418,N_23630);
or U23806 (N_23806,N_23409,N_23530);
nand U23807 (N_23807,N_23551,N_23466);
nor U23808 (N_23808,N_23410,N_23405);
and U23809 (N_23809,N_23622,N_23604);
xnor U23810 (N_23810,N_23624,N_23482);
nor U23811 (N_23811,N_23691,N_23689);
or U23812 (N_23812,N_23629,N_23558);
and U23813 (N_23813,N_23676,N_23507);
xor U23814 (N_23814,N_23504,N_23491);
nand U23815 (N_23815,N_23535,N_23440);
nand U23816 (N_23816,N_23614,N_23464);
or U23817 (N_23817,N_23638,N_23699);
nand U23818 (N_23818,N_23692,N_23505);
nor U23819 (N_23819,N_23667,N_23452);
nor U23820 (N_23820,N_23542,N_23567);
nand U23821 (N_23821,N_23565,N_23403);
xor U23822 (N_23822,N_23664,N_23445);
xnor U23823 (N_23823,N_23643,N_23549);
or U23824 (N_23824,N_23528,N_23648);
or U23825 (N_23825,N_23621,N_23654);
xor U23826 (N_23826,N_23576,N_23431);
xnor U23827 (N_23827,N_23677,N_23458);
nand U23828 (N_23828,N_23516,N_23685);
nand U23829 (N_23829,N_23538,N_23653);
and U23830 (N_23830,N_23446,N_23432);
and U23831 (N_23831,N_23531,N_23625);
xnor U23832 (N_23832,N_23506,N_23472);
nand U23833 (N_23833,N_23512,N_23650);
nor U23834 (N_23834,N_23591,N_23583);
nor U23835 (N_23835,N_23443,N_23465);
xor U23836 (N_23836,N_23414,N_23647);
xor U23837 (N_23837,N_23523,N_23686);
or U23838 (N_23838,N_23413,N_23493);
or U23839 (N_23839,N_23485,N_23442);
and U23840 (N_23840,N_23500,N_23682);
xnor U23841 (N_23841,N_23444,N_23571);
nor U23842 (N_23842,N_23585,N_23424);
and U23843 (N_23843,N_23520,N_23626);
and U23844 (N_23844,N_23420,N_23474);
xnor U23845 (N_23845,N_23545,N_23517);
nor U23846 (N_23846,N_23562,N_23671);
nand U23847 (N_23847,N_23634,N_23475);
xnor U23848 (N_23848,N_23641,N_23417);
or U23849 (N_23849,N_23595,N_23678);
or U23850 (N_23850,N_23544,N_23537);
nand U23851 (N_23851,N_23649,N_23679);
and U23852 (N_23852,N_23514,N_23644);
nor U23853 (N_23853,N_23528,N_23516);
or U23854 (N_23854,N_23664,N_23463);
nor U23855 (N_23855,N_23529,N_23674);
xnor U23856 (N_23856,N_23452,N_23597);
nand U23857 (N_23857,N_23665,N_23540);
nor U23858 (N_23858,N_23442,N_23571);
or U23859 (N_23859,N_23533,N_23439);
and U23860 (N_23860,N_23421,N_23586);
or U23861 (N_23861,N_23684,N_23622);
or U23862 (N_23862,N_23468,N_23633);
and U23863 (N_23863,N_23486,N_23666);
nor U23864 (N_23864,N_23589,N_23573);
or U23865 (N_23865,N_23622,N_23639);
nor U23866 (N_23866,N_23573,N_23587);
or U23867 (N_23867,N_23535,N_23515);
and U23868 (N_23868,N_23675,N_23448);
or U23869 (N_23869,N_23513,N_23509);
nand U23870 (N_23870,N_23538,N_23536);
nand U23871 (N_23871,N_23686,N_23440);
or U23872 (N_23872,N_23531,N_23416);
xor U23873 (N_23873,N_23403,N_23423);
xnor U23874 (N_23874,N_23472,N_23512);
xor U23875 (N_23875,N_23627,N_23653);
xor U23876 (N_23876,N_23418,N_23596);
nor U23877 (N_23877,N_23472,N_23561);
or U23878 (N_23878,N_23440,N_23536);
nor U23879 (N_23879,N_23663,N_23615);
nor U23880 (N_23880,N_23510,N_23482);
nand U23881 (N_23881,N_23585,N_23566);
nor U23882 (N_23882,N_23569,N_23410);
xor U23883 (N_23883,N_23661,N_23542);
nor U23884 (N_23884,N_23588,N_23480);
nor U23885 (N_23885,N_23461,N_23603);
nand U23886 (N_23886,N_23645,N_23520);
nand U23887 (N_23887,N_23653,N_23579);
or U23888 (N_23888,N_23406,N_23654);
nor U23889 (N_23889,N_23475,N_23536);
xnor U23890 (N_23890,N_23566,N_23589);
nand U23891 (N_23891,N_23560,N_23531);
and U23892 (N_23892,N_23680,N_23421);
and U23893 (N_23893,N_23612,N_23402);
or U23894 (N_23894,N_23628,N_23640);
nand U23895 (N_23895,N_23600,N_23679);
nor U23896 (N_23896,N_23562,N_23637);
nor U23897 (N_23897,N_23560,N_23611);
or U23898 (N_23898,N_23598,N_23435);
or U23899 (N_23899,N_23481,N_23679);
nor U23900 (N_23900,N_23591,N_23557);
nand U23901 (N_23901,N_23612,N_23647);
and U23902 (N_23902,N_23605,N_23680);
and U23903 (N_23903,N_23610,N_23499);
nand U23904 (N_23904,N_23596,N_23678);
and U23905 (N_23905,N_23503,N_23432);
nand U23906 (N_23906,N_23465,N_23454);
and U23907 (N_23907,N_23488,N_23483);
or U23908 (N_23908,N_23660,N_23630);
nor U23909 (N_23909,N_23532,N_23685);
or U23910 (N_23910,N_23614,N_23620);
and U23911 (N_23911,N_23427,N_23617);
nor U23912 (N_23912,N_23626,N_23627);
or U23913 (N_23913,N_23565,N_23626);
nor U23914 (N_23914,N_23686,N_23659);
and U23915 (N_23915,N_23538,N_23662);
nor U23916 (N_23916,N_23591,N_23553);
or U23917 (N_23917,N_23648,N_23698);
xor U23918 (N_23918,N_23535,N_23610);
nor U23919 (N_23919,N_23624,N_23635);
xnor U23920 (N_23920,N_23423,N_23641);
and U23921 (N_23921,N_23439,N_23493);
nor U23922 (N_23922,N_23565,N_23528);
nor U23923 (N_23923,N_23626,N_23504);
nor U23924 (N_23924,N_23669,N_23430);
and U23925 (N_23925,N_23621,N_23570);
xnor U23926 (N_23926,N_23585,N_23561);
nor U23927 (N_23927,N_23654,N_23674);
nand U23928 (N_23928,N_23620,N_23540);
nand U23929 (N_23929,N_23526,N_23625);
and U23930 (N_23930,N_23401,N_23595);
xnor U23931 (N_23931,N_23499,N_23695);
or U23932 (N_23932,N_23663,N_23641);
xnor U23933 (N_23933,N_23674,N_23533);
nand U23934 (N_23934,N_23516,N_23417);
or U23935 (N_23935,N_23519,N_23687);
nand U23936 (N_23936,N_23449,N_23583);
nor U23937 (N_23937,N_23541,N_23600);
and U23938 (N_23938,N_23430,N_23592);
nor U23939 (N_23939,N_23629,N_23433);
xnor U23940 (N_23940,N_23687,N_23503);
nand U23941 (N_23941,N_23449,N_23557);
nand U23942 (N_23942,N_23583,N_23684);
xnor U23943 (N_23943,N_23456,N_23637);
nand U23944 (N_23944,N_23689,N_23646);
or U23945 (N_23945,N_23465,N_23433);
nand U23946 (N_23946,N_23549,N_23511);
nor U23947 (N_23947,N_23646,N_23492);
nand U23948 (N_23948,N_23523,N_23574);
xnor U23949 (N_23949,N_23654,N_23466);
nand U23950 (N_23950,N_23665,N_23478);
xnor U23951 (N_23951,N_23687,N_23427);
and U23952 (N_23952,N_23699,N_23463);
xor U23953 (N_23953,N_23425,N_23480);
nor U23954 (N_23954,N_23566,N_23647);
nand U23955 (N_23955,N_23482,N_23672);
nor U23956 (N_23956,N_23506,N_23547);
xnor U23957 (N_23957,N_23515,N_23659);
nor U23958 (N_23958,N_23500,N_23557);
and U23959 (N_23959,N_23429,N_23699);
or U23960 (N_23960,N_23520,N_23681);
and U23961 (N_23961,N_23622,N_23403);
and U23962 (N_23962,N_23495,N_23410);
or U23963 (N_23963,N_23676,N_23682);
or U23964 (N_23964,N_23590,N_23544);
nand U23965 (N_23965,N_23544,N_23530);
nor U23966 (N_23966,N_23481,N_23479);
and U23967 (N_23967,N_23614,N_23538);
or U23968 (N_23968,N_23645,N_23546);
nor U23969 (N_23969,N_23548,N_23498);
nor U23970 (N_23970,N_23613,N_23429);
nor U23971 (N_23971,N_23475,N_23483);
nor U23972 (N_23972,N_23416,N_23489);
nor U23973 (N_23973,N_23595,N_23641);
or U23974 (N_23974,N_23551,N_23587);
or U23975 (N_23975,N_23411,N_23548);
nor U23976 (N_23976,N_23619,N_23543);
and U23977 (N_23977,N_23636,N_23498);
nor U23978 (N_23978,N_23605,N_23577);
nor U23979 (N_23979,N_23441,N_23661);
nor U23980 (N_23980,N_23439,N_23634);
xnor U23981 (N_23981,N_23568,N_23601);
nand U23982 (N_23982,N_23495,N_23423);
xor U23983 (N_23983,N_23659,N_23561);
nor U23984 (N_23984,N_23436,N_23607);
nand U23985 (N_23985,N_23547,N_23609);
nor U23986 (N_23986,N_23523,N_23695);
and U23987 (N_23987,N_23424,N_23605);
and U23988 (N_23988,N_23627,N_23660);
or U23989 (N_23989,N_23676,N_23536);
xor U23990 (N_23990,N_23484,N_23541);
nand U23991 (N_23991,N_23524,N_23533);
and U23992 (N_23992,N_23485,N_23599);
nand U23993 (N_23993,N_23599,N_23486);
nor U23994 (N_23994,N_23483,N_23424);
or U23995 (N_23995,N_23643,N_23563);
and U23996 (N_23996,N_23630,N_23515);
or U23997 (N_23997,N_23545,N_23536);
xnor U23998 (N_23998,N_23544,N_23414);
xor U23999 (N_23999,N_23503,N_23558);
nor U24000 (N_24000,N_23724,N_23734);
nand U24001 (N_24001,N_23886,N_23969);
nand U24002 (N_24002,N_23779,N_23878);
and U24003 (N_24003,N_23850,N_23730);
nor U24004 (N_24004,N_23804,N_23813);
nand U24005 (N_24005,N_23739,N_23719);
nand U24006 (N_24006,N_23748,N_23713);
xnor U24007 (N_24007,N_23950,N_23865);
and U24008 (N_24008,N_23907,N_23841);
or U24009 (N_24009,N_23728,N_23760);
xnor U24010 (N_24010,N_23992,N_23765);
nand U24011 (N_24011,N_23960,N_23857);
xnor U24012 (N_24012,N_23717,N_23711);
nor U24013 (N_24013,N_23993,N_23921);
nand U24014 (N_24014,N_23922,N_23811);
and U24015 (N_24015,N_23831,N_23877);
or U24016 (N_24016,N_23936,N_23819);
xor U24017 (N_24017,N_23957,N_23727);
and U24018 (N_24018,N_23823,N_23942);
nor U24019 (N_24019,N_23762,N_23836);
xor U24020 (N_24020,N_23966,N_23832);
and U24021 (N_24021,N_23704,N_23733);
nand U24022 (N_24022,N_23741,N_23926);
or U24023 (N_24023,N_23833,N_23732);
or U24024 (N_24024,N_23737,N_23964);
and U24025 (N_24025,N_23754,N_23888);
nand U24026 (N_24026,N_23934,N_23860);
and U24027 (N_24027,N_23961,N_23837);
nor U24028 (N_24028,N_23978,N_23894);
and U24029 (N_24029,N_23736,N_23712);
xor U24030 (N_24030,N_23847,N_23856);
nand U24031 (N_24031,N_23842,N_23979);
nand U24032 (N_24032,N_23740,N_23801);
nor U24033 (N_24033,N_23987,N_23786);
xor U24034 (N_24034,N_23884,N_23827);
and U24035 (N_24035,N_23773,N_23974);
and U24036 (N_24036,N_23889,N_23759);
and U24037 (N_24037,N_23803,N_23795);
and U24038 (N_24038,N_23800,N_23753);
xnor U24039 (N_24039,N_23797,N_23814);
and U24040 (N_24040,N_23875,N_23780);
nand U24041 (N_24041,N_23913,N_23710);
and U24042 (N_24042,N_23862,N_23903);
nand U24043 (N_24043,N_23977,N_23720);
or U24044 (N_24044,N_23876,N_23943);
nor U24045 (N_24045,N_23777,N_23920);
nor U24046 (N_24046,N_23703,N_23802);
or U24047 (N_24047,N_23916,N_23988);
xor U24048 (N_24048,N_23822,N_23905);
nor U24049 (N_24049,N_23805,N_23817);
or U24050 (N_24050,N_23815,N_23967);
or U24051 (N_24051,N_23947,N_23812);
xnor U24052 (N_24052,N_23887,N_23818);
or U24053 (N_24053,N_23873,N_23744);
nand U24054 (N_24054,N_23756,N_23839);
nand U24055 (N_24055,N_23864,N_23882);
nand U24056 (N_24056,N_23866,N_23830);
xor U24057 (N_24057,N_23743,N_23859);
or U24058 (N_24058,N_23941,N_23844);
xor U24059 (N_24059,N_23828,N_23932);
and U24060 (N_24060,N_23789,N_23949);
xor U24061 (N_24061,N_23925,N_23787);
or U24062 (N_24062,N_23790,N_23799);
nand U24063 (N_24063,N_23846,N_23915);
or U24064 (N_24064,N_23928,N_23778);
nor U24065 (N_24065,N_23810,N_23820);
nor U24066 (N_24066,N_23930,N_23821);
or U24067 (N_24067,N_23870,N_23763);
xor U24068 (N_24068,N_23924,N_23793);
or U24069 (N_24069,N_23955,N_23749);
nand U24070 (N_24070,N_23874,N_23718);
nand U24071 (N_24071,N_23808,N_23959);
and U24072 (N_24072,N_23895,N_23852);
xor U24073 (N_24073,N_23791,N_23963);
nand U24074 (N_24074,N_23906,N_23902);
and U24075 (N_24075,N_23958,N_23854);
and U24076 (N_24076,N_23707,N_23742);
nor U24077 (N_24077,N_23807,N_23745);
and U24078 (N_24078,N_23776,N_23824);
or U24079 (N_24079,N_23984,N_23723);
and U24080 (N_24080,N_23702,N_23935);
nor U24081 (N_24081,N_23994,N_23785);
or U24082 (N_24082,N_23904,N_23953);
xor U24083 (N_24083,N_23829,N_23881);
nor U24084 (N_24084,N_23918,N_23991);
or U24085 (N_24085,N_23701,N_23998);
xor U24086 (N_24086,N_23982,N_23772);
xnor U24087 (N_24087,N_23910,N_23806);
nand U24088 (N_24088,N_23757,N_23900);
nor U24089 (N_24089,N_23954,N_23867);
nand U24090 (N_24090,N_23851,N_23911);
nand U24091 (N_24091,N_23968,N_23775);
xor U24092 (N_24092,N_23892,N_23764);
nor U24093 (N_24093,N_23809,N_23970);
and U24094 (N_24094,N_23869,N_23845);
nor U24095 (N_24095,N_23986,N_23995);
or U24096 (N_24096,N_23834,N_23835);
nand U24097 (N_24097,N_23853,N_23996);
xnor U24098 (N_24098,N_23972,N_23825);
xnor U24099 (N_24099,N_23976,N_23898);
xor U24100 (N_24100,N_23956,N_23783);
xor U24101 (N_24101,N_23938,N_23927);
nand U24102 (N_24102,N_23937,N_23971);
xor U24103 (N_24103,N_23784,N_23879);
nand U24104 (N_24104,N_23989,N_23990);
nor U24105 (N_24105,N_23899,N_23973);
xnor U24106 (N_24106,N_23735,N_23939);
nand U24107 (N_24107,N_23826,N_23917);
and U24108 (N_24108,N_23774,N_23933);
nor U24109 (N_24109,N_23883,N_23891);
nand U24110 (N_24110,N_23893,N_23944);
nor U24111 (N_24111,N_23999,N_23709);
and U24112 (N_24112,N_23729,N_23750);
xor U24113 (N_24113,N_23716,N_23722);
and U24114 (N_24114,N_23975,N_23962);
xnor U24115 (N_24115,N_23731,N_23767);
nand U24116 (N_24116,N_23738,N_23769);
nor U24117 (N_24117,N_23983,N_23768);
and U24118 (N_24118,N_23940,N_23700);
and U24119 (N_24119,N_23848,N_23912);
and U24120 (N_24120,N_23923,N_23946);
and U24121 (N_24121,N_23725,N_23872);
and U24122 (N_24122,N_23751,N_23914);
or U24123 (N_24123,N_23840,N_23794);
and U24124 (N_24124,N_23746,N_23788);
or U24125 (N_24125,N_23755,N_23965);
or U24126 (N_24126,N_23909,N_23766);
xor U24127 (N_24127,N_23792,N_23985);
nand U24128 (N_24128,N_23816,N_23849);
xor U24129 (N_24129,N_23715,N_23908);
xor U24130 (N_24130,N_23901,N_23747);
nand U24131 (N_24131,N_23770,N_23885);
xnor U24132 (N_24132,N_23796,N_23863);
or U24133 (N_24133,N_23897,N_23952);
or U24134 (N_24134,N_23714,N_23896);
nor U24135 (N_24135,N_23855,N_23708);
and U24136 (N_24136,N_23706,N_23880);
xnor U24137 (N_24137,N_23843,N_23761);
xnor U24138 (N_24138,N_23771,N_23948);
xnor U24139 (N_24139,N_23798,N_23929);
xnor U24140 (N_24140,N_23981,N_23890);
nand U24141 (N_24141,N_23871,N_23861);
and U24142 (N_24142,N_23781,N_23919);
or U24143 (N_24143,N_23705,N_23758);
and U24144 (N_24144,N_23951,N_23752);
nor U24145 (N_24145,N_23726,N_23721);
xor U24146 (N_24146,N_23868,N_23997);
and U24147 (N_24147,N_23931,N_23838);
nand U24148 (N_24148,N_23945,N_23858);
nand U24149 (N_24149,N_23980,N_23782);
or U24150 (N_24150,N_23883,N_23949);
nand U24151 (N_24151,N_23810,N_23840);
xnor U24152 (N_24152,N_23868,N_23740);
nand U24153 (N_24153,N_23720,N_23737);
or U24154 (N_24154,N_23933,N_23892);
and U24155 (N_24155,N_23975,N_23979);
nand U24156 (N_24156,N_23959,N_23922);
nand U24157 (N_24157,N_23792,N_23946);
nor U24158 (N_24158,N_23843,N_23939);
and U24159 (N_24159,N_23834,N_23800);
or U24160 (N_24160,N_23748,N_23940);
nor U24161 (N_24161,N_23948,N_23934);
xnor U24162 (N_24162,N_23709,N_23974);
nand U24163 (N_24163,N_23851,N_23983);
nand U24164 (N_24164,N_23929,N_23890);
and U24165 (N_24165,N_23701,N_23719);
nand U24166 (N_24166,N_23704,N_23764);
nor U24167 (N_24167,N_23976,N_23795);
xnor U24168 (N_24168,N_23712,N_23759);
and U24169 (N_24169,N_23755,N_23851);
or U24170 (N_24170,N_23819,N_23757);
nor U24171 (N_24171,N_23763,N_23983);
nand U24172 (N_24172,N_23719,N_23778);
nand U24173 (N_24173,N_23844,N_23956);
or U24174 (N_24174,N_23972,N_23798);
and U24175 (N_24175,N_23755,N_23961);
or U24176 (N_24176,N_23840,N_23959);
xnor U24177 (N_24177,N_23924,N_23960);
nand U24178 (N_24178,N_23720,N_23925);
or U24179 (N_24179,N_23796,N_23730);
or U24180 (N_24180,N_23796,N_23789);
or U24181 (N_24181,N_23775,N_23724);
nor U24182 (N_24182,N_23984,N_23718);
xnor U24183 (N_24183,N_23798,N_23747);
nor U24184 (N_24184,N_23736,N_23871);
xnor U24185 (N_24185,N_23842,N_23860);
nand U24186 (N_24186,N_23848,N_23858);
and U24187 (N_24187,N_23705,N_23910);
xnor U24188 (N_24188,N_23932,N_23968);
or U24189 (N_24189,N_23719,N_23981);
nand U24190 (N_24190,N_23861,N_23842);
nor U24191 (N_24191,N_23987,N_23799);
nor U24192 (N_24192,N_23945,N_23760);
and U24193 (N_24193,N_23884,N_23879);
nor U24194 (N_24194,N_23803,N_23948);
and U24195 (N_24195,N_23939,N_23807);
xnor U24196 (N_24196,N_23935,N_23896);
nor U24197 (N_24197,N_23817,N_23787);
nor U24198 (N_24198,N_23953,N_23869);
or U24199 (N_24199,N_23956,N_23937);
and U24200 (N_24200,N_23856,N_23876);
nor U24201 (N_24201,N_23857,N_23930);
xnor U24202 (N_24202,N_23946,N_23882);
nor U24203 (N_24203,N_23947,N_23798);
nor U24204 (N_24204,N_23875,N_23808);
nor U24205 (N_24205,N_23899,N_23827);
nand U24206 (N_24206,N_23828,N_23772);
nor U24207 (N_24207,N_23980,N_23848);
and U24208 (N_24208,N_23842,N_23933);
nor U24209 (N_24209,N_23970,N_23960);
or U24210 (N_24210,N_23744,N_23752);
and U24211 (N_24211,N_23951,N_23812);
xnor U24212 (N_24212,N_23907,N_23735);
and U24213 (N_24213,N_23981,N_23933);
and U24214 (N_24214,N_23788,N_23775);
nand U24215 (N_24215,N_23879,N_23757);
xor U24216 (N_24216,N_23987,N_23726);
and U24217 (N_24217,N_23945,N_23824);
or U24218 (N_24218,N_23728,N_23995);
xnor U24219 (N_24219,N_23925,N_23851);
nand U24220 (N_24220,N_23873,N_23733);
and U24221 (N_24221,N_23915,N_23966);
xor U24222 (N_24222,N_23940,N_23934);
and U24223 (N_24223,N_23796,N_23775);
xnor U24224 (N_24224,N_23722,N_23749);
xor U24225 (N_24225,N_23761,N_23890);
and U24226 (N_24226,N_23996,N_23744);
nand U24227 (N_24227,N_23874,N_23818);
and U24228 (N_24228,N_23804,N_23743);
nor U24229 (N_24229,N_23991,N_23994);
xor U24230 (N_24230,N_23774,N_23883);
nor U24231 (N_24231,N_23970,N_23997);
nor U24232 (N_24232,N_23711,N_23896);
nor U24233 (N_24233,N_23876,N_23900);
nand U24234 (N_24234,N_23800,N_23879);
nor U24235 (N_24235,N_23918,N_23741);
nand U24236 (N_24236,N_23728,N_23787);
xor U24237 (N_24237,N_23826,N_23725);
nand U24238 (N_24238,N_23989,N_23851);
xnor U24239 (N_24239,N_23828,N_23906);
xnor U24240 (N_24240,N_23824,N_23802);
xnor U24241 (N_24241,N_23795,N_23804);
nand U24242 (N_24242,N_23792,N_23842);
xor U24243 (N_24243,N_23875,N_23705);
and U24244 (N_24244,N_23800,N_23881);
and U24245 (N_24245,N_23992,N_23858);
xnor U24246 (N_24246,N_23919,N_23949);
or U24247 (N_24247,N_23987,N_23877);
or U24248 (N_24248,N_23765,N_23858);
or U24249 (N_24249,N_23782,N_23865);
nor U24250 (N_24250,N_23795,N_23841);
xor U24251 (N_24251,N_23796,N_23779);
nor U24252 (N_24252,N_23819,N_23761);
and U24253 (N_24253,N_23991,N_23721);
or U24254 (N_24254,N_23931,N_23730);
nand U24255 (N_24255,N_23866,N_23732);
nor U24256 (N_24256,N_23708,N_23838);
xnor U24257 (N_24257,N_23865,N_23766);
or U24258 (N_24258,N_23905,N_23925);
nor U24259 (N_24259,N_23878,N_23883);
nor U24260 (N_24260,N_23919,N_23864);
nand U24261 (N_24261,N_23944,N_23788);
nand U24262 (N_24262,N_23857,N_23962);
nand U24263 (N_24263,N_23992,N_23844);
nor U24264 (N_24264,N_23814,N_23958);
nor U24265 (N_24265,N_23806,N_23907);
xnor U24266 (N_24266,N_23888,N_23968);
nand U24267 (N_24267,N_23917,N_23974);
nand U24268 (N_24268,N_23909,N_23920);
nand U24269 (N_24269,N_23985,N_23946);
nand U24270 (N_24270,N_23786,N_23758);
nand U24271 (N_24271,N_23761,N_23771);
xor U24272 (N_24272,N_23794,N_23810);
or U24273 (N_24273,N_23741,N_23996);
and U24274 (N_24274,N_23877,N_23922);
nand U24275 (N_24275,N_23987,N_23750);
xor U24276 (N_24276,N_23955,N_23885);
nor U24277 (N_24277,N_23811,N_23832);
nand U24278 (N_24278,N_23863,N_23947);
or U24279 (N_24279,N_23974,N_23761);
or U24280 (N_24280,N_23754,N_23886);
nor U24281 (N_24281,N_23824,N_23816);
nor U24282 (N_24282,N_23783,N_23954);
nand U24283 (N_24283,N_23827,N_23881);
or U24284 (N_24284,N_23975,N_23745);
nor U24285 (N_24285,N_23944,N_23860);
and U24286 (N_24286,N_23798,N_23979);
or U24287 (N_24287,N_23811,N_23876);
or U24288 (N_24288,N_23852,N_23762);
or U24289 (N_24289,N_23751,N_23929);
nor U24290 (N_24290,N_23707,N_23810);
nor U24291 (N_24291,N_23701,N_23771);
nand U24292 (N_24292,N_23928,N_23932);
xnor U24293 (N_24293,N_23821,N_23814);
nor U24294 (N_24294,N_23937,N_23831);
and U24295 (N_24295,N_23821,N_23954);
xor U24296 (N_24296,N_23773,N_23754);
nor U24297 (N_24297,N_23912,N_23855);
and U24298 (N_24298,N_23883,N_23791);
nand U24299 (N_24299,N_23895,N_23921);
or U24300 (N_24300,N_24107,N_24075);
or U24301 (N_24301,N_24015,N_24116);
nor U24302 (N_24302,N_24241,N_24064);
and U24303 (N_24303,N_24145,N_24211);
xor U24304 (N_24304,N_24005,N_24087);
or U24305 (N_24305,N_24168,N_24082);
or U24306 (N_24306,N_24181,N_24163);
xor U24307 (N_24307,N_24101,N_24115);
or U24308 (N_24308,N_24249,N_24024);
xnor U24309 (N_24309,N_24261,N_24166);
nand U24310 (N_24310,N_24222,N_24191);
and U24311 (N_24311,N_24004,N_24045);
nor U24312 (N_24312,N_24276,N_24006);
xor U24313 (N_24313,N_24210,N_24277);
nand U24314 (N_24314,N_24054,N_24170);
nand U24315 (N_24315,N_24028,N_24287);
nand U24316 (N_24316,N_24259,N_24032);
and U24317 (N_24317,N_24150,N_24144);
and U24318 (N_24318,N_24068,N_24072);
xnor U24319 (N_24319,N_24117,N_24043);
or U24320 (N_24320,N_24111,N_24256);
nor U24321 (N_24321,N_24027,N_24169);
and U24322 (N_24322,N_24238,N_24047);
nor U24323 (N_24323,N_24153,N_24281);
xor U24324 (N_24324,N_24013,N_24127);
nor U24325 (N_24325,N_24297,N_24227);
xnor U24326 (N_24326,N_24177,N_24262);
nor U24327 (N_24327,N_24193,N_24001);
and U24328 (N_24328,N_24282,N_24011);
and U24329 (N_24329,N_24129,N_24212);
nor U24330 (N_24330,N_24288,N_24190);
xnor U24331 (N_24331,N_24050,N_24201);
xor U24332 (N_24332,N_24065,N_24076);
xor U24333 (N_24333,N_24188,N_24199);
and U24334 (N_24334,N_24203,N_24074);
or U24335 (N_24335,N_24073,N_24096);
xnor U24336 (N_24336,N_24205,N_24062);
xor U24337 (N_24337,N_24292,N_24112);
or U24338 (N_24338,N_24114,N_24067);
xnor U24339 (N_24339,N_24186,N_24198);
or U24340 (N_24340,N_24136,N_24159);
nand U24341 (N_24341,N_24274,N_24160);
nor U24342 (N_24342,N_24118,N_24021);
nand U24343 (N_24343,N_24202,N_24183);
and U24344 (N_24344,N_24030,N_24132);
xor U24345 (N_24345,N_24046,N_24023);
nor U24346 (N_24346,N_24290,N_24229);
nand U24347 (N_24347,N_24059,N_24156);
and U24348 (N_24348,N_24128,N_24206);
and U24349 (N_24349,N_24061,N_24296);
or U24350 (N_24350,N_24138,N_24265);
nand U24351 (N_24351,N_24099,N_24167);
nor U24352 (N_24352,N_24063,N_24134);
and U24353 (N_24353,N_24095,N_24180);
and U24354 (N_24354,N_24230,N_24234);
nand U24355 (N_24355,N_24052,N_24187);
xor U24356 (N_24356,N_24056,N_24279);
nand U24357 (N_24357,N_24143,N_24051);
or U24358 (N_24358,N_24091,N_24025);
nand U24359 (N_24359,N_24247,N_24041);
nor U24360 (N_24360,N_24066,N_24228);
xor U24361 (N_24361,N_24020,N_24236);
nand U24362 (N_24362,N_24079,N_24235);
and U24363 (N_24363,N_24295,N_24184);
xor U24364 (N_24364,N_24103,N_24185);
xor U24365 (N_24365,N_24218,N_24273);
nand U24366 (N_24366,N_24192,N_24098);
or U24367 (N_24367,N_24215,N_24240);
xor U24368 (N_24368,N_24033,N_24171);
xnor U24369 (N_24369,N_24182,N_24008);
xor U24370 (N_24370,N_24179,N_24034);
and U24371 (N_24371,N_24083,N_24239);
xnor U24372 (N_24372,N_24044,N_24258);
nor U24373 (N_24373,N_24016,N_24286);
nand U24374 (N_24374,N_24175,N_24264);
nand U24375 (N_24375,N_24246,N_24263);
xnor U24376 (N_24376,N_24251,N_24130);
or U24377 (N_24377,N_24086,N_24084);
nand U24378 (N_24378,N_24208,N_24070);
xor U24379 (N_24379,N_24283,N_24142);
nor U24380 (N_24380,N_24233,N_24197);
xor U24381 (N_24381,N_24172,N_24154);
xor U24382 (N_24382,N_24140,N_24007);
and U24383 (N_24383,N_24060,N_24146);
nor U24384 (N_24384,N_24161,N_24289);
or U24385 (N_24385,N_24100,N_24176);
xnor U24386 (N_24386,N_24120,N_24037);
nor U24387 (N_24387,N_24189,N_24242);
nor U24388 (N_24388,N_24194,N_24105);
nor U24389 (N_24389,N_24058,N_24108);
xnor U24390 (N_24390,N_24124,N_24085);
nor U24391 (N_24391,N_24260,N_24029);
xnor U24392 (N_24392,N_24255,N_24254);
nand U24393 (N_24393,N_24121,N_24225);
nor U24394 (N_24394,N_24017,N_24071);
and U24395 (N_24395,N_24040,N_24269);
and U24396 (N_24396,N_24223,N_24137);
nand U24397 (N_24397,N_24152,N_24147);
xor U24398 (N_24398,N_24113,N_24135);
xor U24399 (N_24399,N_24026,N_24131);
nor U24400 (N_24400,N_24220,N_24231);
xnor U24401 (N_24401,N_24195,N_24055);
and U24402 (N_24402,N_24110,N_24275);
or U24403 (N_24403,N_24093,N_24232);
xor U24404 (N_24404,N_24216,N_24092);
nor U24405 (N_24405,N_24155,N_24217);
xor U24406 (N_24406,N_24294,N_24162);
nand U24407 (N_24407,N_24009,N_24019);
xnor U24408 (N_24408,N_24226,N_24042);
and U24409 (N_24409,N_24158,N_24053);
nor U24410 (N_24410,N_24012,N_24039);
xnor U24411 (N_24411,N_24250,N_24278);
nand U24412 (N_24412,N_24209,N_24003);
nand U24413 (N_24413,N_24245,N_24031);
and U24414 (N_24414,N_24224,N_24077);
xor U24415 (N_24415,N_24293,N_24257);
and U24416 (N_24416,N_24204,N_24038);
xnor U24417 (N_24417,N_24000,N_24097);
nor U24418 (N_24418,N_24069,N_24139);
or U24419 (N_24419,N_24022,N_24078);
xnor U24420 (N_24420,N_24148,N_24106);
and U24421 (N_24421,N_24164,N_24048);
nand U24422 (N_24422,N_24243,N_24119);
nand U24423 (N_24423,N_24291,N_24094);
and U24424 (N_24424,N_24213,N_24080);
nor U24425 (N_24425,N_24244,N_24125);
or U24426 (N_24426,N_24122,N_24266);
and U24427 (N_24427,N_24252,N_24272);
nor U24428 (N_24428,N_24271,N_24149);
nand U24429 (N_24429,N_24270,N_24104);
xor U24430 (N_24430,N_24298,N_24268);
nor U24431 (N_24431,N_24126,N_24299);
nor U24432 (N_24432,N_24173,N_24102);
nand U24433 (N_24433,N_24141,N_24133);
nand U24434 (N_24434,N_24090,N_24221);
nand U24435 (N_24435,N_24165,N_24151);
nand U24436 (N_24436,N_24280,N_24267);
nand U24437 (N_24437,N_24174,N_24178);
nor U24438 (N_24438,N_24002,N_24248);
nand U24439 (N_24439,N_24109,N_24088);
and U24440 (N_24440,N_24200,N_24157);
nor U24441 (N_24441,N_24036,N_24219);
and U24442 (N_24442,N_24081,N_24237);
nand U24443 (N_24443,N_24035,N_24207);
nand U24444 (N_24444,N_24089,N_24010);
nand U24445 (N_24445,N_24285,N_24284);
or U24446 (N_24446,N_24014,N_24123);
nand U24447 (N_24447,N_24196,N_24214);
and U24448 (N_24448,N_24253,N_24049);
or U24449 (N_24449,N_24057,N_24018);
xor U24450 (N_24450,N_24051,N_24287);
nor U24451 (N_24451,N_24053,N_24169);
and U24452 (N_24452,N_24079,N_24053);
nand U24453 (N_24453,N_24154,N_24285);
nand U24454 (N_24454,N_24128,N_24117);
and U24455 (N_24455,N_24040,N_24012);
or U24456 (N_24456,N_24011,N_24290);
nor U24457 (N_24457,N_24243,N_24251);
and U24458 (N_24458,N_24296,N_24224);
or U24459 (N_24459,N_24262,N_24092);
xnor U24460 (N_24460,N_24031,N_24123);
or U24461 (N_24461,N_24044,N_24108);
or U24462 (N_24462,N_24239,N_24159);
or U24463 (N_24463,N_24132,N_24189);
and U24464 (N_24464,N_24130,N_24253);
and U24465 (N_24465,N_24000,N_24295);
nor U24466 (N_24466,N_24175,N_24195);
nor U24467 (N_24467,N_24282,N_24008);
nand U24468 (N_24468,N_24282,N_24170);
xor U24469 (N_24469,N_24089,N_24082);
xnor U24470 (N_24470,N_24299,N_24024);
xnor U24471 (N_24471,N_24044,N_24122);
xnor U24472 (N_24472,N_24030,N_24104);
nand U24473 (N_24473,N_24067,N_24093);
xnor U24474 (N_24474,N_24107,N_24081);
or U24475 (N_24475,N_24002,N_24211);
and U24476 (N_24476,N_24090,N_24087);
or U24477 (N_24477,N_24239,N_24090);
and U24478 (N_24478,N_24273,N_24176);
nor U24479 (N_24479,N_24147,N_24265);
xor U24480 (N_24480,N_24191,N_24167);
or U24481 (N_24481,N_24067,N_24286);
or U24482 (N_24482,N_24093,N_24019);
nand U24483 (N_24483,N_24049,N_24047);
nand U24484 (N_24484,N_24218,N_24193);
nor U24485 (N_24485,N_24249,N_24151);
xnor U24486 (N_24486,N_24135,N_24221);
nand U24487 (N_24487,N_24121,N_24029);
nor U24488 (N_24488,N_24082,N_24190);
or U24489 (N_24489,N_24103,N_24013);
nor U24490 (N_24490,N_24152,N_24011);
nand U24491 (N_24491,N_24287,N_24211);
nor U24492 (N_24492,N_24066,N_24123);
xnor U24493 (N_24493,N_24212,N_24047);
nand U24494 (N_24494,N_24236,N_24291);
nor U24495 (N_24495,N_24159,N_24180);
nand U24496 (N_24496,N_24106,N_24260);
nand U24497 (N_24497,N_24183,N_24082);
nand U24498 (N_24498,N_24028,N_24071);
and U24499 (N_24499,N_24244,N_24036);
nand U24500 (N_24500,N_24215,N_24110);
xnor U24501 (N_24501,N_24278,N_24094);
and U24502 (N_24502,N_24212,N_24249);
nor U24503 (N_24503,N_24202,N_24294);
xor U24504 (N_24504,N_24035,N_24032);
and U24505 (N_24505,N_24181,N_24148);
and U24506 (N_24506,N_24002,N_24278);
xnor U24507 (N_24507,N_24100,N_24227);
or U24508 (N_24508,N_24062,N_24266);
xor U24509 (N_24509,N_24224,N_24017);
nor U24510 (N_24510,N_24200,N_24021);
xor U24511 (N_24511,N_24219,N_24166);
nand U24512 (N_24512,N_24244,N_24052);
nor U24513 (N_24513,N_24053,N_24272);
or U24514 (N_24514,N_24227,N_24190);
nor U24515 (N_24515,N_24154,N_24234);
or U24516 (N_24516,N_24154,N_24248);
nand U24517 (N_24517,N_24154,N_24219);
nor U24518 (N_24518,N_24011,N_24141);
or U24519 (N_24519,N_24125,N_24033);
and U24520 (N_24520,N_24015,N_24265);
and U24521 (N_24521,N_24111,N_24060);
nor U24522 (N_24522,N_24042,N_24229);
nor U24523 (N_24523,N_24256,N_24048);
and U24524 (N_24524,N_24063,N_24193);
xnor U24525 (N_24525,N_24276,N_24161);
nand U24526 (N_24526,N_24174,N_24291);
nor U24527 (N_24527,N_24168,N_24297);
and U24528 (N_24528,N_24123,N_24225);
nand U24529 (N_24529,N_24116,N_24114);
nand U24530 (N_24530,N_24171,N_24012);
and U24531 (N_24531,N_24192,N_24091);
xnor U24532 (N_24532,N_24158,N_24160);
nor U24533 (N_24533,N_24014,N_24287);
nor U24534 (N_24534,N_24078,N_24142);
or U24535 (N_24535,N_24127,N_24184);
xor U24536 (N_24536,N_24149,N_24068);
or U24537 (N_24537,N_24230,N_24248);
xor U24538 (N_24538,N_24117,N_24269);
xnor U24539 (N_24539,N_24022,N_24203);
nand U24540 (N_24540,N_24025,N_24008);
xnor U24541 (N_24541,N_24004,N_24026);
nor U24542 (N_24542,N_24106,N_24011);
nor U24543 (N_24543,N_24099,N_24011);
nor U24544 (N_24544,N_24259,N_24104);
nand U24545 (N_24545,N_24206,N_24278);
or U24546 (N_24546,N_24267,N_24138);
nand U24547 (N_24547,N_24101,N_24131);
or U24548 (N_24548,N_24295,N_24153);
or U24549 (N_24549,N_24030,N_24138);
or U24550 (N_24550,N_24229,N_24018);
nor U24551 (N_24551,N_24058,N_24095);
nor U24552 (N_24552,N_24113,N_24184);
or U24553 (N_24553,N_24049,N_24252);
and U24554 (N_24554,N_24112,N_24065);
nand U24555 (N_24555,N_24177,N_24272);
or U24556 (N_24556,N_24251,N_24295);
nand U24557 (N_24557,N_24279,N_24016);
or U24558 (N_24558,N_24041,N_24092);
nor U24559 (N_24559,N_24089,N_24163);
nor U24560 (N_24560,N_24149,N_24016);
nor U24561 (N_24561,N_24106,N_24159);
and U24562 (N_24562,N_24284,N_24169);
xor U24563 (N_24563,N_24055,N_24057);
nor U24564 (N_24564,N_24005,N_24048);
nor U24565 (N_24565,N_24024,N_24032);
nor U24566 (N_24566,N_24084,N_24221);
or U24567 (N_24567,N_24001,N_24132);
and U24568 (N_24568,N_24137,N_24292);
nor U24569 (N_24569,N_24265,N_24150);
nand U24570 (N_24570,N_24202,N_24215);
xor U24571 (N_24571,N_24129,N_24254);
xnor U24572 (N_24572,N_24088,N_24171);
nand U24573 (N_24573,N_24077,N_24037);
nand U24574 (N_24574,N_24011,N_24053);
and U24575 (N_24575,N_24111,N_24020);
xor U24576 (N_24576,N_24179,N_24228);
or U24577 (N_24577,N_24023,N_24216);
and U24578 (N_24578,N_24265,N_24293);
nor U24579 (N_24579,N_24101,N_24221);
or U24580 (N_24580,N_24291,N_24145);
xnor U24581 (N_24581,N_24143,N_24182);
xor U24582 (N_24582,N_24038,N_24285);
xor U24583 (N_24583,N_24145,N_24237);
nand U24584 (N_24584,N_24205,N_24116);
or U24585 (N_24585,N_24189,N_24095);
xnor U24586 (N_24586,N_24194,N_24109);
nand U24587 (N_24587,N_24044,N_24101);
nand U24588 (N_24588,N_24176,N_24026);
xnor U24589 (N_24589,N_24231,N_24131);
xor U24590 (N_24590,N_24092,N_24274);
and U24591 (N_24591,N_24205,N_24165);
or U24592 (N_24592,N_24268,N_24062);
and U24593 (N_24593,N_24001,N_24122);
nand U24594 (N_24594,N_24063,N_24069);
nand U24595 (N_24595,N_24056,N_24224);
or U24596 (N_24596,N_24041,N_24031);
or U24597 (N_24597,N_24256,N_24015);
or U24598 (N_24598,N_24294,N_24257);
or U24599 (N_24599,N_24085,N_24206);
nor U24600 (N_24600,N_24572,N_24384);
nand U24601 (N_24601,N_24400,N_24588);
xnor U24602 (N_24602,N_24470,N_24399);
nor U24603 (N_24603,N_24359,N_24308);
or U24604 (N_24604,N_24348,N_24346);
and U24605 (N_24605,N_24430,N_24582);
nand U24606 (N_24606,N_24301,N_24403);
or U24607 (N_24607,N_24366,N_24448);
nor U24608 (N_24608,N_24445,N_24435);
or U24609 (N_24609,N_24369,N_24475);
and U24610 (N_24610,N_24482,N_24313);
or U24611 (N_24611,N_24554,N_24454);
or U24612 (N_24612,N_24500,N_24335);
nor U24613 (N_24613,N_24375,N_24570);
or U24614 (N_24614,N_24391,N_24559);
xnor U24615 (N_24615,N_24552,N_24450);
and U24616 (N_24616,N_24441,N_24349);
and U24617 (N_24617,N_24396,N_24537);
or U24618 (N_24618,N_24498,N_24446);
nand U24619 (N_24619,N_24584,N_24327);
and U24620 (N_24620,N_24342,N_24513);
or U24621 (N_24621,N_24465,N_24533);
or U24622 (N_24622,N_24434,N_24458);
xor U24623 (N_24623,N_24364,N_24317);
nand U24624 (N_24624,N_24426,N_24550);
nor U24625 (N_24625,N_24388,N_24480);
xor U24626 (N_24626,N_24367,N_24436);
or U24627 (N_24627,N_24468,N_24325);
nor U24628 (N_24628,N_24319,N_24438);
nand U24629 (N_24629,N_24521,N_24451);
or U24630 (N_24630,N_24376,N_24493);
or U24631 (N_24631,N_24423,N_24562);
and U24632 (N_24632,N_24352,N_24383);
xor U24633 (N_24633,N_24504,N_24495);
or U24634 (N_24634,N_24315,N_24431);
nand U24635 (N_24635,N_24569,N_24303);
and U24636 (N_24636,N_24525,N_24425);
nand U24637 (N_24637,N_24326,N_24336);
or U24638 (N_24638,N_24437,N_24380);
or U24639 (N_24639,N_24305,N_24517);
nand U24640 (N_24640,N_24402,N_24401);
or U24641 (N_24641,N_24474,N_24432);
and U24642 (N_24642,N_24372,N_24501);
xor U24643 (N_24643,N_24463,N_24549);
and U24644 (N_24644,N_24444,N_24574);
nor U24645 (N_24645,N_24338,N_24520);
nor U24646 (N_24646,N_24331,N_24389);
nand U24647 (N_24647,N_24515,N_24377);
or U24648 (N_24648,N_24339,N_24539);
nand U24649 (N_24649,N_24421,N_24528);
nor U24650 (N_24650,N_24427,N_24361);
or U24651 (N_24651,N_24412,N_24408);
and U24652 (N_24652,N_24439,N_24486);
or U24653 (N_24653,N_24394,N_24512);
xor U24654 (N_24654,N_24510,N_24589);
or U24655 (N_24655,N_24548,N_24507);
or U24656 (N_24656,N_24575,N_24362);
and U24657 (N_24657,N_24527,N_24485);
nand U24658 (N_24658,N_24419,N_24347);
and U24659 (N_24659,N_24344,N_24395);
nor U24660 (N_24660,N_24545,N_24566);
nand U24661 (N_24661,N_24576,N_24511);
xnor U24662 (N_24662,N_24534,N_24387);
nand U24663 (N_24663,N_24540,N_24573);
or U24664 (N_24664,N_24370,N_24553);
or U24665 (N_24665,N_24586,N_24557);
or U24666 (N_24666,N_24476,N_24373);
nor U24667 (N_24667,N_24538,N_24484);
and U24668 (N_24668,N_24343,N_24543);
nand U24669 (N_24669,N_24453,N_24508);
or U24670 (N_24670,N_24580,N_24378);
nand U24671 (N_24671,N_24505,N_24420);
nor U24672 (N_24672,N_24316,N_24332);
or U24673 (N_24673,N_24531,N_24466);
nor U24674 (N_24674,N_24302,N_24487);
and U24675 (N_24675,N_24320,N_24506);
xnor U24676 (N_24676,N_24304,N_24494);
nand U24677 (N_24677,N_24462,N_24565);
nor U24678 (N_24678,N_24481,N_24314);
nand U24679 (N_24679,N_24404,N_24499);
or U24680 (N_24680,N_24357,N_24488);
xor U24681 (N_24681,N_24595,N_24546);
or U24682 (N_24682,N_24447,N_24371);
nand U24683 (N_24683,N_24307,N_24321);
or U24684 (N_24684,N_24330,N_24312);
and U24685 (N_24685,N_24502,N_24392);
nor U24686 (N_24686,N_24567,N_24407);
xnor U24687 (N_24687,N_24583,N_24522);
or U24688 (N_24688,N_24405,N_24341);
nand U24689 (N_24689,N_24353,N_24577);
xor U24690 (N_24690,N_24382,N_24532);
and U24691 (N_24691,N_24328,N_24422);
nor U24692 (N_24692,N_24479,N_24418);
nand U24693 (N_24693,N_24443,N_24597);
or U24694 (N_24694,N_24509,N_24599);
and U24695 (N_24695,N_24491,N_24581);
or U24696 (N_24696,N_24542,N_24558);
nor U24697 (N_24697,N_24568,N_24490);
nand U24698 (N_24698,N_24306,N_24452);
nor U24699 (N_24699,N_24415,N_24593);
and U24700 (N_24700,N_24477,N_24417);
xnor U24701 (N_24701,N_24355,N_24469);
and U24702 (N_24702,N_24591,N_24428);
nand U24703 (N_24703,N_24345,N_24350);
nor U24704 (N_24704,N_24406,N_24547);
and U24705 (N_24705,N_24464,N_24414);
nand U24706 (N_24706,N_24351,N_24524);
xnor U24707 (N_24707,N_24544,N_24503);
nand U24708 (N_24708,N_24449,N_24478);
and U24709 (N_24709,N_24322,N_24529);
or U24710 (N_24710,N_24311,N_24472);
nor U24711 (N_24711,N_24492,N_24497);
and U24712 (N_24712,N_24598,N_24535);
nor U24713 (N_24713,N_24496,N_24440);
xor U24714 (N_24714,N_24358,N_24333);
nor U24715 (N_24715,N_24363,N_24354);
and U24716 (N_24716,N_24386,N_24587);
nor U24717 (N_24717,N_24471,N_24416);
nor U24718 (N_24718,N_24519,N_24526);
nor U24719 (N_24719,N_24556,N_24555);
or U24720 (N_24720,N_24393,N_24579);
and U24721 (N_24721,N_24560,N_24324);
or U24722 (N_24722,N_24518,N_24374);
nor U24723 (N_24723,N_24455,N_24483);
and U24724 (N_24724,N_24467,N_24442);
and U24725 (N_24725,N_24360,N_24596);
and U24726 (N_24726,N_24585,N_24429);
and U24727 (N_24727,N_24541,N_24424);
and U24728 (N_24728,N_24459,N_24337);
nor U24729 (N_24729,N_24318,N_24592);
xor U24730 (N_24730,N_24300,N_24516);
nor U24731 (N_24731,N_24571,N_24564);
and U24732 (N_24732,N_24340,N_24530);
or U24733 (N_24733,N_24561,N_24410);
xnor U24734 (N_24734,N_24594,N_24409);
nor U24735 (N_24735,N_24590,N_24489);
nand U24736 (N_24736,N_24385,N_24381);
and U24737 (N_24737,N_24398,N_24356);
or U24738 (N_24738,N_24473,N_24368);
nor U24739 (N_24739,N_24457,N_24411);
or U24740 (N_24740,N_24329,N_24323);
xor U24741 (N_24741,N_24413,N_24563);
and U24742 (N_24742,N_24460,N_24310);
nor U24743 (N_24743,N_24365,N_24433);
nand U24744 (N_24744,N_24578,N_24397);
and U24745 (N_24745,N_24334,N_24390);
or U24746 (N_24746,N_24379,N_24536);
nand U24747 (N_24747,N_24456,N_24461);
nor U24748 (N_24748,N_24514,N_24309);
nand U24749 (N_24749,N_24523,N_24551);
nor U24750 (N_24750,N_24364,N_24521);
xor U24751 (N_24751,N_24554,N_24356);
or U24752 (N_24752,N_24443,N_24337);
xor U24753 (N_24753,N_24552,N_24487);
xor U24754 (N_24754,N_24564,N_24595);
and U24755 (N_24755,N_24509,N_24533);
xor U24756 (N_24756,N_24551,N_24418);
and U24757 (N_24757,N_24515,N_24508);
xor U24758 (N_24758,N_24484,N_24524);
and U24759 (N_24759,N_24388,N_24406);
or U24760 (N_24760,N_24418,N_24382);
xnor U24761 (N_24761,N_24435,N_24366);
nand U24762 (N_24762,N_24415,N_24333);
xor U24763 (N_24763,N_24583,N_24461);
or U24764 (N_24764,N_24560,N_24334);
nand U24765 (N_24765,N_24541,N_24545);
and U24766 (N_24766,N_24582,N_24391);
xnor U24767 (N_24767,N_24544,N_24476);
or U24768 (N_24768,N_24490,N_24342);
nor U24769 (N_24769,N_24446,N_24402);
nand U24770 (N_24770,N_24557,N_24357);
xor U24771 (N_24771,N_24310,N_24578);
and U24772 (N_24772,N_24477,N_24469);
or U24773 (N_24773,N_24303,N_24349);
and U24774 (N_24774,N_24334,N_24332);
and U24775 (N_24775,N_24481,N_24460);
nand U24776 (N_24776,N_24368,N_24303);
and U24777 (N_24777,N_24589,N_24501);
nand U24778 (N_24778,N_24379,N_24463);
and U24779 (N_24779,N_24563,N_24426);
xor U24780 (N_24780,N_24484,N_24405);
and U24781 (N_24781,N_24316,N_24550);
or U24782 (N_24782,N_24443,N_24366);
or U24783 (N_24783,N_24309,N_24372);
nand U24784 (N_24784,N_24528,N_24334);
or U24785 (N_24785,N_24342,N_24480);
and U24786 (N_24786,N_24495,N_24370);
nand U24787 (N_24787,N_24470,N_24370);
or U24788 (N_24788,N_24512,N_24505);
nand U24789 (N_24789,N_24402,N_24489);
nor U24790 (N_24790,N_24470,N_24532);
or U24791 (N_24791,N_24333,N_24414);
nor U24792 (N_24792,N_24377,N_24576);
and U24793 (N_24793,N_24344,N_24331);
xnor U24794 (N_24794,N_24474,N_24334);
nor U24795 (N_24795,N_24395,N_24472);
nand U24796 (N_24796,N_24459,N_24406);
xnor U24797 (N_24797,N_24425,N_24435);
nand U24798 (N_24798,N_24342,N_24456);
nand U24799 (N_24799,N_24417,N_24507);
and U24800 (N_24800,N_24448,N_24576);
or U24801 (N_24801,N_24434,N_24372);
and U24802 (N_24802,N_24344,N_24343);
xor U24803 (N_24803,N_24487,N_24319);
or U24804 (N_24804,N_24314,N_24488);
xnor U24805 (N_24805,N_24483,N_24450);
xor U24806 (N_24806,N_24555,N_24401);
nand U24807 (N_24807,N_24413,N_24326);
nand U24808 (N_24808,N_24547,N_24364);
and U24809 (N_24809,N_24375,N_24558);
and U24810 (N_24810,N_24383,N_24359);
nand U24811 (N_24811,N_24374,N_24547);
and U24812 (N_24812,N_24552,N_24405);
nand U24813 (N_24813,N_24493,N_24373);
xor U24814 (N_24814,N_24578,N_24515);
nor U24815 (N_24815,N_24581,N_24467);
nor U24816 (N_24816,N_24366,N_24596);
nor U24817 (N_24817,N_24434,N_24320);
xor U24818 (N_24818,N_24489,N_24398);
and U24819 (N_24819,N_24425,N_24579);
and U24820 (N_24820,N_24333,N_24471);
and U24821 (N_24821,N_24449,N_24564);
xor U24822 (N_24822,N_24562,N_24348);
nand U24823 (N_24823,N_24509,N_24447);
nand U24824 (N_24824,N_24417,N_24483);
xnor U24825 (N_24825,N_24443,N_24406);
nand U24826 (N_24826,N_24516,N_24503);
and U24827 (N_24827,N_24361,N_24381);
nor U24828 (N_24828,N_24361,N_24476);
nand U24829 (N_24829,N_24406,N_24395);
and U24830 (N_24830,N_24542,N_24535);
or U24831 (N_24831,N_24497,N_24559);
or U24832 (N_24832,N_24407,N_24453);
or U24833 (N_24833,N_24554,N_24403);
xnor U24834 (N_24834,N_24309,N_24330);
and U24835 (N_24835,N_24324,N_24359);
nand U24836 (N_24836,N_24397,N_24554);
and U24837 (N_24837,N_24571,N_24566);
xor U24838 (N_24838,N_24306,N_24488);
or U24839 (N_24839,N_24560,N_24594);
and U24840 (N_24840,N_24538,N_24574);
nor U24841 (N_24841,N_24375,N_24468);
nor U24842 (N_24842,N_24565,N_24485);
xnor U24843 (N_24843,N_24480,N_24449);
or U24844 (N_24844,N_24568,N_24433);
or U24845 (N_24845,N_24475,N_24549);
nand U24846 (N_24846,N_24535,N_24578);
xor U24847 (N_24847,N_24478,N_24455);
nand U24848 (N_24848,N_24552,N_24390);
xor U24849 (N_24849,N_24348,N_24577);
xor U24850 (N_24850,N_24569,N_24475);
and U24851 (N_24851,N_24566,N_24363);
or U24852 (N_24852,N_24454,N_24426);
nand U24853 (N_24853,N_24310,N_24471);
nand U24854 (N_24854,N_24509,N_24569);
nor U24855 (N_24855,N_24437,N_24329);
nand U24856 (N_24856,N_24468,N_24388);
nand U24857 (N_24857,N_24345,N_24580);
or U24858 (N_24858,N_24330,N_24362);
xor U24859 (N_24859,N_24423,N_24465);
nor U24860 (N_24860,N_24312,N_24541);
xnor U24861 (N_24861,N_24345,N_24459);
nand U24862 (N_24862,N_24589,N_24548);
nor U24863 (N_24863,N_24360,N_24524);
xor U24864 (N_24864,N_24525,N_24554);
nor U24865 (N_24865,N_24390,N_24556);
or U24866 (N_24866,N_24547,N_24342);
xnor U24867 (N_24867,N_24471,N_24306);
nand U24868 (N_24868,N_24492,N_24366);
nand U24869 (N_24869,N_24422,N_24414);
or U24870 (N_24870,N_24423,N_24413);
and U24871 (N_24871,N_24394,N_24523);
or U24872 (N_24872,N_24520,N_24573);
xnor U24873 (N_24873,N_24395,N_24435);
or U24874 (N_24874,N_24572,N_24338);
and U24875 (N_24875,N_24498,N_24459);
or U24876 (N_24876,N_24359,N_24341);
or U24877 (N_24877,N_24302,N_24468);
or U24878 (N_24878,N_24461,N_24453);
nand U24879 (N_24879,N_24544,N_24534);
xor U24880 (N_24880,N_24567,N_24558);
nand U24881 (N_24881,N_24346,N_24410);
nand U24882 (N_24882,N_24340,N_24584);
and U24883 (N_24883,N_24454,N_24473);
xnor U24884 (N_24884,N_24311,N_24392);
nand U24885 (N_24885,N_24488,N_24523);
nand U24886 (N_24886,N_24410,N_24351);
and U24887 (N_24887,N_24560,N_24392);
xor U24888 (N_24888,N_24593,N_24426);
and U24889 (N_24889,N_24593,N_24598);
nor U24890 (N_24890,N_24445,N_24578);
nand U24891 (N_24891,N_24475,N_24491);
or U24892 (N_24892,N_24389,N_24362);
or U24893 (N_24893,N_24427,N_24552);
nor U24894 (N_24894,N_24578,N_24485);
nand U24895 (N_24895,N_24510,N_24536);
xor U24896 (N_24896,N_24550,N_24334);
nand U24897 (N_24897,N_24565,N_24498);
or U24898 (N_24898,N_24517,N_24542);
xnor U24899 (N_24899,N_24440,N_24374);
nand U24900 (N_24900,N_24773,N_24811);
and U24901 (N_24901,N_24642,N_24662);
and U24902 (N_24902,N_24776,N_24667);
nand U24903 (N_24903,N_24777,N_24756);
nand U24904 (N_24904,N_24890,N_24889);
and U24905 (N_24905,N_24767,N_24719);
and U24906 (N_24906,N_24800,N_24749);
nor U24907 (N_24907,N_24651,N_24782);
or U24908 (N_24908,N_24859,N_24857);
and U24909 (N_24909,N_24637,N_24673);
or U24910 (N_24910,N_24631,N_24623);
nand U24911 (N_24911,N_24609,N_24712);
xor U24912 (N_24912,N_24624,N_24751);
and U24913 (N_24913,N_24748,N_24701);
xor U24914 (N_24914,N_24725,N_24818);
or U24915 (N_24915,N_24675,N_24614);
nand U24916 (N_24916,N_24763,N_24718);
or U24917 (N_24917,N_24657,N_24850);
nand U24918 (N_24918,N_24722,N_24634);
and U24919 (N_24919,N_24611,N_24691);
and U24920 (N_24920,N_24689,N_24666);
and U24921 (N_24921,N_24787,N_24726);
and U24922 (N_24922,N_24703,N_24677);
or U24923 (N_24923,N_24600,N_24660);
nand U24924 (N_24924,N_24752,N_24664);
or U24925 (N_24925,N_24815,N_24622);
and U24926 (N_24926,N_24669,N_24710);
xnor U24927 (N_24927,N_24698,N_24647);
nor U24928 (N_24928,N_24661,N_24806);
nand U24929 (N_24929,N_24605,N_24682);
xor U24930 (N_24930,N_24692,N_24617);
xor U24931 (N_24931,N_24625,N_24741);
and U24932 (N_24932,N_24670,N_24835);
nand U24933 (N_24933,N_24855,N_24868);
or U24934 (N_24934,N_24744,N_24709);
nand U24935 (N_24935,N_24872,N_24863);
or U24936 (N_24936,N_24869,N_24804);
and U24937 (N_24937,N_24791,N_24728);
or U24938 (N_24938,N_24711,N_24615);
and U24939 (N_24939,N_24760,N_24616);
nor U24940 (N_24940,N_24650,N_24892);
and U24941 (N_24941,N_24653,N_24731);
and U24942 (N_24942,N_24607,N_24619);
nor U24943 (N_24943,N_24780,N_24796);
xnor U24944 (N_24944,N_24674,N_24739);
or U24945 (N_24945,N_24628,N_24789);
nand U24946 (N_24946,N_24747,N_24668);
or U24947 (N_24947,N_24658,N_24684);
xor U24948 (N_24948,N_24715,N_24795);
nand U24949 (N_24949,N_24817,N_24633);
or U24950 (N_24950,N_24785,N_24823);
nor U24951 (N_24951,N_24608,N_24851);
or U24952 (N_24952,N_24734,N_24706);
or U24953 (N_24953,N_24781,N_24893);
or U24954 (N_24954,N_24813,N_24758);
and U24955 (N_24955,N_24814,N_24862);
nor U24956 (N_24956,N_24672,N_24688);
nand U24957 (N_24957,N_24648,N_24694);
nand U24958 (N_24958,N_24879,N_24831);
nand U24959 (N_24959,N_24884,N_24833);
and U24960 (N_24960,N_24839,N_24696);
and U24961 (N_24961,N_24654,N_24630);
nand U24962 (N_24962,N_24699,N_24742);
or U24963 (N_24963,N_24641,N_24656);
nand U24964 (N_24964,N_24663,N_24700);
xnor U24965 (N_24965,N_24730,N_24613);
and U24966 (N_24966,N_24768,N_24881);
or U24967 (N_24967,N_24612,N_24603);
nor U24968 (N_24968,N_24895,N_24871);
nand U24969 (N_24969,N_24632,N_24860);
nand U24970 (N_24970,N_24717,N_24652);
xor U24971 (N_24971,N_24671,N_24626);
nor U24972 (N_24972,N_24878,N_24792);
nand U24973 (N_24973,N_24841,N_24784);
and U24974 (N_24974,N_24679,N_24897);
nor U24975 (N_24975,N_24894,N_24604);
or U24976 (N_24976,N_24783,N_24870);
nand U24977 (N_24977,N_24874,N_24723);
nor U24978 (N_24978,N_24610,N_24743);
xnor U24979 (N_24979,N_24707,N_24721);
xor U24980 (N_24980,N_24816,N_24759);
nand U24981 (N_24981,N_24853,N_24645);
nor U24982 (N_24982,N_24770,N_24812);
xor U24983 (N_24983,N_24713,N_24635);
or U24984 (N_24984,N_24690,N_24858);
nor U24985 (N_24985,N_24724,N_24888);
nor U24986 (N_24986,N_24819,N_24793);
and U24987 (N_24987,N_24809,N_24798);
nor U24988 (N_24988,N_24774,N_24882);
xnor U24989 (N_24989,N_24765,N_24627);
nor U24990 (N_24990,N_24824,N_24753);
xor U24991 (N_24991,N_24766,N_24886);
or U24992 (N_24992,N_24716,N_24877);
or U24993 (N_24993,N_24695,N_24738);
and U24994 (N_24994,N_24810,N_24762);
xor U24995 (N_24995,N_24643,N_24832);
nand U24996 (N_24996,N_24827,N_24891);
nand U24997 (N_24997,N_24786,N_24757);
nor U24998 (N_24998,N_24842,N_24705);
or U24999 (N_24999,N_24830,N_24720);
xnor U25000 (N_25000,N_24865,N_24733);
or U25001 (N_25001,N_24794,N_24704);
xnor U25002 (N_25002,N_24880,N_24828);
or U25003 (N_25003,N_24686,N_24807);
or U25004 (N_25004,N_24867,N_24856);
xnor U25005 (N_25005,N_24640,N_24649);
xnor U25006 (N_25006,N_24693,N_24746);
or U25007 (N_25007,N_24779,N_24834);
and U25008 (N_25008,N_24801,N_24829);
and U25009 (N_25009,N_24875,N_24646);
and U25010 (N_25010,N_24852,N_24771);
and U25011 (N_25011,N_24848,N_24764);
nand U25012 (N_25012,N_24638,N_24644);
nand U25013 (N_25013,N_24676,N_24639);
nand U25014 (N_25014,N_24896,N_24799);
nor U25015 (N_25015,N_24845,N_24846);
xor U25016 (N_25016,N_24772,N_24714);
xor U25017 (N_25017,N_24887,N_24737);
or U25018 (N_25018,N_24601,N_24797);
or U25019 (N_25019,N_24775,N_24826);
xor U25020 (N_25020,N_24864,N_24655);
or U25021 (N_25021,N_24750,N_24727);
and U25022 (N_25022,N_24697,N_24636);
or U25023 (N_25023,N_24849,N_24821);
nand U25024 (N_25024,N_24755,N_24876);
and U25025 (N_25025,N_24825,N_24899);
and U25026 (N_25026,N_24735,N_24803);
and U25027 (N_25027,N_24847,N_24732);
xnor U25028 (N_25028,N_24898,N_24620);
xor U25029 (N_25029,N_24822,N_24736);
nor U25030 (N_25030,N_24708,N_24618);
xnor U25031 (N_25031,N_24680,N_24836);
nor U25032 (N_25032,N_24740,N_24659);
or U25033 (N_25033,N_24602,N_24861);
and U25034 (N_25034,N_24883,N_24769);
xnor U25035 (N_25035,N_24843,N_24778);
nor U25036 (N_25036,N_24678,N_24702);
nor U25037 (N_25037,N_24844,N_24873);
nand U25038 (N_25038,N_24808,N_24621);
xnor U25039 (N_25039,N_24665,N_24790);
or U25040 (N_25040,N_24687,N_24840);
and U25041 (N_25041,N_24683,N_24761);
and U25042 (N_25042,N_24820,N_24837);
nand U25043 (N_25043,N_24681,N_24854);
nand U25044 (N_25044,N_24838,N_24788);
nand U25045 (N_25045,N_24629,N_24729);
and U25046 (N_25046,N_24685,N_24802);
xor U25047 (N_25047,N_24754,N_24745);
nand U25048 (N_25048,N_24606,N_24866);
or U25049 (N_25049,N_24885,N_24805);
or U25050 (N_25050,N_24836,N_24641);
or U25051 (N_25051,N_24773,N_24628);
or U25052 (N_25052,N_24779,N_24721);
nand U25053 (N_25053,N_24876,N_24816);
xor U25054 (N_25054,N_24692,N_24742);
nor U25055 (N_25055,N_24630,N_24807);
and U25056 (N_25056,N_24751,N_24621);
and U25057 (N_25057,N_24646,N_24755);
and U25058 (N_25058,N_24820,N_24605);
nand U25059 (N_25059,N_24774,N_24756);
and U25060 (N_25060,N_24601,N_24654);
and U25061 (N_25061,N_24625,N_24680);
nand U25062 (N_25062,N_24732,N_24810);
nor U25063 (N_25063,N_24778,N_24739);
xnor U25064 (N_25064,N_24619,N_24766);
or U25065 (N_25065,N_24851,N_24693);
xor U25066 (N_25066,N_24608,N_24894);
or U25067 (N_25067,N_24656,N_24816);
xor U25068 (N_25068,N_24749,N_24651);
and U25069 (N_25069,N_24602,N_24798);
nand U25070 (N_25070,N_24841,N_24831);
nand U25071 (N_25071,N_24607,N_24896);
xnor U25072 (N_25072,N_24852,N_24718);
nand U25073 (N_25073,N_24654,N_24755);
nor U25074 (N_25074,N_24792,N_24700);
and U25075 (N_25075,N_24718,N_24751);
nor U25076 (N_25076,N_24829,N_24775);
and U25077 (N_25077,N_24607,N_24824);
nand U25078 (N_25078,N_24637,N_24677);
nand U25079 (N_25079,N_24783,N_24779);
nor U25080 (N_25080,N_24712,N_24749);
and U25081 (N_25081,N_24684,N_24766);
nor U25082 (N_25082,N_24771,N_24640);
nand U25083 (N_25083,N_24802,N_24820);
nor U25084 (N_25084,N_24601,N_24812);
xor U25085 (N_25085,N_24723,N_24642);
and U25086 (N_25086,N_24858,N_24618);
nand U25087 (N_25087,N_24843,N_24672);
and U25088 (N_25088,N_24830,N_24721);
or U25089 (N_25089,N_24775,N_24649);
and U25090 (N_25090,N_24697,N_24796);
or U25091 (N_25091,N_24644,N_24837);
xor U25092 (N_25092,N_24835,N_24627);
xor U25093 (N_25093,N_24679,N_24850);
nor U25094 (N_25094,N_24658,N_24856);
nor U25095 (N_25095,N_24754,N_24721);
xnor U25096 (N_25096,N_24813,N_24783);
or U25097 (N_25097,N_24762,N_24896);
nand U25098 (N_25098,N_24722,N_24894);
nand U25099 (N_25099,N_24697,N_24802);
xnor U25100 (N_25100,N_24801,N_24838);
xnor U25101 (N_25101,N_24657,N_24890);
and U25102 (N_25102,N_24837,N_24813);
nor U25103 (N_25103,N_24719,N_24661);
xnor U25104 (N_25104,N_24671,N_24700);
nand U25105 (N_25105,N_24861,N_24843);
nand U25106 (N_25106,N_24716,N_24832);
xnor U25107 (N_25107,N_24739,N_24810);
nor U25108 (N_25108,N_24690,N_24660);
nor U25109 (N_25109,N_24636,N_24639);
and U25110 (N_25110,N_24836,N_24834);
nor U25111 (N_25111,N_24632,N_24633);
xor U25112 (N_25112,N_24650,N_24710);
and U25113 (N_25113,N_24887,N_24641);
and U25114 (N_25114,N_24883,N_24789);
nor U25115 (N_25115,N_24661,N_24805);
or U25116 (N_25116,N_24699,N_24801);
nand U25117 (N_25117,N_24791,N_24698);
xnor U25118 (N_25118,N_24700,N_24623);
xnor U25119 (N_25119,N_24714,N_24771);
xor U25120 (N_25120,N_24894,N_24771);
nor U25121 (N_25121,N_24890,N_24646);
or U25122 (N_25122,N_24899,N_24884);
xor U25123 (N_25123,N_24751,N_24899);
or U25124 (N_25124,N_24871,N_24767);
nand U25125 (N_25125,N_24803,N_24760);
and U25126 (N_25126,N_24744,N_24887);
nor U25127 (N_25127,N_24791,N_24628);
and U25128 (N_25128,N_24869,N_24768);
or U25129 (N_25129,N_24622,N_24828);
xor U25130 (N_25130,N_24731,N_24670);
xor U25131 (N_25131,N_24658,N_24743);
and U25132 (N_25132,N_24809,N_24860);
or U25133 (N_25133,N_24698,N_24649);
nor U25134 (N_25134,N_24738,N_24743);
xnor U25135 (N_25135,N_24684,N_24687);
or U25136 (N_25136,N_24735,N_24642);
nand U25137 (N_25137,N_24689,N_24749);
or U25138 (N_25138,N_24720,N_24776);
xnor U25139 (N_25139,N_24664,N_24796);
xnor U25140 (N_25140,N_24760,N_24770);
nor U25141 (N_25141,N_24838,N_24786);
and U25142 (N_25142,N_24762,N_24723);
xor U25143 (N_25143,N_24861,N_24827);
or U25144 (N_25144,N_24653,N_24675);
or U25145 (N_25145,N_24627,N_24739);
or U25146 (N_25146,N_24673,N_24609);
nor U25147 (N_25147,N_24784,N_24794);
xor U25148 (N_25148,N_24876,N_24812);
nor U25149 (N_25149,N_24770,N_24815);
and U25150 (N_25150,N_24672,N_24847);
xnor U25151 (N_25151,N_24890,N_24756);
or U25152 (N_25152,N_24733,N_24732);
xnor U25153 (N_25153,N_24711,N_24810);
and U25154 (N_25154,N_24899,N_24765);
xnor U25155 (N_25155,N_24749,N_24799);
or U25156 (N_25156,N_24781,N_24632);
or U25157 (N_25157,N_24727,N_24791);
nand U25158 (N_25158,N_24651,N_24653);
or U25159 (N_25159,N_24685,N_24753);
nand U25160 (N_25160,N_24834,N_24770);
or U25161 (N_25161,N_24710,N_24728);
or U25162 (N_25162,N_24814,N_24820);
and U25163 (N_25163,N_24778,N_24750);
or U25164 (N_25164,N_24724,N_24678);
or U25165 (N_25165,N_24646,N_24667);
or U25166 (N_25166,N_24717,N_24787);
xnor U25167 (N_25167,N_24843,N_24701);
xnor U25168 (N_25168,N_24805,N_24612);
nand U25169 (N_25169,N_24836,N_24654);
xnor U25170 (N_25170,N_24743,N_24698);
and U25171 (N_25171,N_24726,N_24653);
or U25172 (N_25172,N_24703,N_24811);
and U25173 (N_25173,N_24642,N_24853);
or U25174 (N_25174,N_24659,N_24601);
and U25175 (N_25175,N_24768,N_24631);
or U25176 (N_25176,N_24775,N_24638);
and U25177 (N_25177,N_24671,N_24869);
nand U25178 (N_25178,N_24789,N_24642);
nor U25179 (N_25179,N_24869,N_24623);
and U25180 (N_25180,N_24718,N_24684);
and U25181 (N_25181,N_24624,N_24791);
xnor U25182 (N_25182,N_24676,N_24613);
nand U25183 (N_25183,N_24617,N_24898);
or U25184 (N_25184,N_24838,N_24750);
xnor U25185 (N_25185,N_24648,N_24731);
or U25186 (N_25186,N_24834,N_24833);
xor U25187 (N_25187,N_24805,N_24722);
nor U25188 (N_25188,N_24661,N_24662);
or U25189 (N_25189,N_24889,N_24650);
xor U25190 (N_25190,N_24744,N_24817);
nor U25191 (N_25191,N_24663,N_24657);
nor U25192 (N_25192,N_24800,N_24777);
or U25193 (N_25193,N_24787,N_24772);
xnor U25194 (N_25194,N_24795,N_24663);
nand U25195 (N_25195,N_24892,N_24834);
or U25196 (N_25196,N_24886,N_24662);
and U25197 (N_25197,N_24720,N_24848);
nor U25198 (N_25198,N_24650,N_24660);
nand U25199 (N_25199,N_24734,N_24843);
or U25200 (N_25200,N_25130,N_24960);
and U25201 (N_25201,N_25138,N_25013);
or U25202 (N_25202,N_25051,N_24988);
or U25203 (N_25203,N_24979,N_25065);
xor U25204 (N_25204,N_25096,N_25137);
and U25205 (N_25205,N_25077,N_24962);
xnor U25206 (N_25206,N_25176,N_24903);
xnor U25207 (N_25207,N_24902,N_25018);
or U25208 (N_25208,N_25181,N_25122);
or U25209 (N_25209,N_25135,N_24920);
nor U25210 (N_25210,N_25136,N_25030);
nor U25211 (N_25211,N_25008,N_24906);
and U25212 (N_25212,N_25174,N_25159);
or U25213 (N_25213,N_25047,N_24956);
or U25214 (N_25214,N_24987,N_24997);
and U25215 (N_25215,N_25022,N_25190);
nand U25216 (N_25216,N_25192,N_25119);
nand U25217 (N_25217,N_25028,N_25070);
nand U25218 (N_25218,N_24952,N_24992);
nor U25219 (N_25219,N_24913,N_25066);
and U25220 (N_25220,N_25011,N_25058);
xnor U25221 (N_25221,N_24976,N_24951);
and U25222 (N_25222,N_24936,N_25179);
nand U25223 (N_25223,N_25154,N_25186);
xnor U25224 (N_25224,N_25015,N_25195);
and U25225 (N_25225,N_25064,N_24989);
xnor U25226 (N_25226,N_25095,N_25105);
and U25227 (N_25227,N_25081,N_25061);
nand U25228 (N_25228,N_25072,N_25032);
and U25229 (N_25229,N_25131,N_24901);
nand U25230 (N_25230,N_24995,N_24963);
and U25231 (N_25231,N_25099,N_24929);
xor U25232 (N_25232,N_25182,N_24925);
xnor U25233 (N_25233,N_25183,N_25053);
xor U25234 (N_25234,N_25000,N_25162);
and U25235 (N_25235,N_24941,N_25090);
or U25236 (N_25236,N_24953,N_25091);
or U25237 (N_25237,N_25088,N_24923);
nand U25238 (N_25238,N_25149,N_24994);
or U25239 (N_25239,N_25123,N_25073);
xor U25240 (N_25240,N_24933,N_25056);
nor U25241 (N_25241,N_25098,N_25161);
nand U25242 (N_25242,N_24955,N_24984);
and U25243 (N_25243,N_25129,N_25045);
nor U25244 (N_25244,N_25026,N_25168);
nand U25245 (N_25245,N_25194,N_25101);
or U25246 (N_25246,N_24990,N_24968);
nand U25247 (N_25247,N_25115,N_25148);
or U25248 (N_25248,N_25164,N_24912);
or U25249 (N_25249,N_25049,N_24939);
or U25250 (N_25250,N_25158,N_25092);
nand U25251 (N_25251,N_24981,N_25150);
nor U25252 (N_25252,N_25003,N_25116);
nor U25253 (N_25253,N_25083,N_25062);
or U25254 (N_25254,N_25126,N_25075);
nand U25255 (N_25255,N_25144,N_25178);
and U25256 (N_25256,N_24938,N_24977);
xnor U25257 (N_25257,N_25108,N_24904);
or U25258 (N_25258,N_24980,N_25020);
or U25259 (N_25259,N_25040,N_25127);
nor U25260 (N_25260,N_25031,N_24983);
nor U25261 (N_25261,N_25079,N_25198);
nor U25262 (N_25262,N_25078,N_24944);
xnor U25263 (N_25263,N_24986,N_24975);
nand U25264 (N_25264,N_24943,N_25102);
nand U25265 (N_25265,N_25025,N_24921);
xnor U25266 (N_25266,N_25069,N_24961);
and U25267 (N_25267,N_25107,N_24965);
and U25268 (N_25268,N_25184,N_24937);
or U25269 (N_25269,N_25089,N_24922);
xor U25270 (N_25270,N_25009,N_25187);
and U25271 (N_25271,N_25146,N_25109);
and U25272 (N_25272,N_24967,N_24926);
or U25273 (N_25273,N_25068,N_25166);
nand U25274 (N_25274,N_25125,N_25170);
nand U25275 (N_25275,N_25171,N_25004);
or U25276 (N_25276,N_25059,N_25063);
or U25277 (N_25277,N_25165,N_25140);
or U25278 (N_25278,N_25046,N_25044);
nor U25279 (N_25279,N_25177,N_24928);
nor U25280 (N_25280,N_24935,N_25001);
and U25281 (N_25281,N_25118,N_25087);
nand U25282 (N_25282,N_24993,N_25139);
nand U25283 (N_25283,N_25104,N_24918);
nor U25284 (N_25284,N_24910,N_25006);
nor U25285 (N_25285,N_25067,N_25050);
or U25286 (N_25286,N_24966,N_25120);
nand U25287 (N_25287,N_25021,N_24934);
xnor U25288 (N_25288,N_25114,N_25017);
nand U25289 (N_25289,N_25048,N_25097);
xnor U25290 (N_25290,N_25023,N_25103);
nand U25291 (N_25291,N_25193,N_25094);
nand U25292 (N_25292,N_25010,N_24964);
and U25293 (N_25293,N_24919,N_25106);
and U25294 (N_25294,N_25110,N_25113);
or U25295 (N_25295,N_24970,N_24957);
nand U25296 (N_25296,N_25111,N_24914);
and U25297 (N_25297,N_25042,N_24958);
and U25298 (N_25298,N_25086,N_25157);
nand U25299 (N_25299,N_25076,N_25145);
or U25300 (N_25300,N_24991,N_25036);
nand U25301 (N_25301,N_25147,N_24908);
xnor U25302 (N_25302,N_24959,N_24971);
or U25303 (N_25303,N_25160,N_25175);
and U25304 (N_25304,N_25156,N_25172);
nand U25305 (N_25305,N_24917,N_25043);
xnor U25306 (N_25306,N_24969,N_25054);
nand U25307 (N_25307,N_25124,N_24996);
nor U25308 (N_25308,N_25173,N_25167);
nor U25309 (N_25309,N_25117,N_25191);
and U25310 (N_25310,N_24974,N_24973);
xor U25311 (N_25311,N_25121,N_25112);
or U25312 (N_25312,N_25084,N_25038);
nand U25313 (N_25313,N_25012,N_25141);
nand U25314 (N_25314,N_25060,N_25163);
xnor U25315 (N_25315,N_24915,N_24948);
xor U25316 (N_25316,N_25037,N_24907);
xnor U25317 (N_25317,N_25153,N_25019);
xor U25318 (N_25318,N_24940,N_25071);
nand U25319 (N_25319,N_25080,N_24982);
and U25320 (N_25320,N_24932,N_25151);
nand U25321 (N_25321,N_25133,N_25197);
xor U25322 (N_25322,N_25093,N_25100);
and U25323 (N_25323,N_25188,N_25057);
nand U25324 (N_25324,N_24946,N_25029);
nand U25325 (N_25325,N_25134,N_25143);
xnor U25326 (N_25326,N_24972,N_25196);
xor U25327 (N_25327,N_25027,N_24931);
nor U25328 (N_25328,N_24911,N_24947);
xor U25329 (N_25329,N_25155,N_24985);
nand U25330 (N_25330,N_25199,N_24924);
xor U25331 (N_25331,N_24930,N_25014);
and U25332 (N_25332,N_25035,N_24916);
and U25333 (N_25333,N_24954,N_25007);
nor U25334 (N_25334,N_25033,N_24927);
nand U25335 (N_25335,N_25185,N_25055);
and U25336 (N_25336,N_25039,N_25034);
nand U25337 (N_25337,N_25189,N_25016);
nor U25338 (N_25338,N_25142,N_24999);
xnor U25339 (N_25339,N_25041,N_25082);
nand U25340 (N_25340,N_24998,N_25024);
or U25341 (N_25341,N_25074,N_24949);
nor U25342 (N_25342,N_25180,N_25132);
nor U25343 (N_25343,N_24945,N_25169);
and U25344 (N_25344,N_25085,N_24950);
nand U25345 (N_25345,N_25128,N_25052);
and U25346 (N_25346,N_24900,N_25002);
nand U25347 (N_25347,N_24905,N_24942);
or U25348 (N_25348,N_24978,N_25152);
nand U25349 (N_25349,N_24909,N_25005);
nor U25350 (N_25350,N_24972,N_24911);
and U25351 (N_25351,N_25129,N_24948);
or U25352 (N_25352,N_25106,N_24942);
nor U25353 (N_25353,N_25106,N_25044);
or U25354 (N_25354,N_24965,N_25155);
and U25355 (N_25355,N_25187,N_24986);
and U25356 (N_25356,N_25073,N_25069);
nand U25357 (N_25357,N_25062,N_25154);
nor U25358 (N_25358,N_25100,N_25169);
nand U25359 (N_25359,N_24989,N_25032);
nor U25360 (N_25360,N_25153,N_25011);
or U25361 (N_25361,N_24923,N_25183);
and U25362 (N_25362,N_25108,N_25016);
or U25363 (N_25363,N_25166,N_25037);
nand U25364 (N_25364,N_25036,N_25154);
nand U25365 (N_25365,N_25088,N_25067);
or U25366 (N_25366,N_24912,N_24951);
nand U25367 (N_25367,N_24961,N_25177);
xor U25368 (N_25368,N_25187,N_24917);
or U25369 (N_25369,N_25090,N_24946);
nor U25370 (N_25370,N_25028,N_25155);
xnor U25371 (N_25371,N_25145,N_24936);
and U25372 (N_25372,N_25086,N_25119);
nor U25373 (N_25373,N_24992,N_25005);
and U25374 (N_25374,N_25199,N_24984);
nor U25375 (N_25375,N_25060,N_25142);
nor U25376 (N_25376,N_24988,N_25178);
nand U25377 (N_25377,N_25069,N_25142);
or U25378 (N_25378,N_24995,N_25160);
and U25379 (N_25379,N_24933,N_24955);
xor U25380 (N_25380,N_25068,N_25062);
or U25381 (N_25381,N_24959,N_25021);
nor U25382 (N_25382,N_25187,N_25013);
nor U25383 (N_25383,N_25118,N_24969);
xnor U25384 (N_25384,N_25108,N_25132);
nor U25385 (N_25385,N_25095,N_25076);
and U25386 (N_25386,N_25052,N_25112);
and U25387 (N_25387,N_25153,N_25141);
nor U25388 (N_25388,N_25175,N_25104);
or U25389 (N_25389,N_24923,N_25120);
nand U25390 (N_25390,N_24961,N_25172);
and U25391 (N_25391,N_24973,N_25078);
nand U25392 (N_25392,N_25164,N_25146);
nand U25393 (N_25393,N_25033,N_24979);
or U25394 (N_25394,N_24910,N_25138);
and U25395 (N_25395,N_24978,N_24928);
nor U25396 (N_25396,N_25139,N_24945);
or U25397 (N_25397,N_25191,N_25182);
nand U25398 (N_25398,N_24923,N_24942);
or U25399 (N_25399,N_25184,N_25072);
nand U25400 (N_25400,N_24956,N_24947);
nor U25401 (N_25401,N_24958,N_24971);
nand U25402 (N_25402,N_25107,N_24923);
or U25403 (N_25403,N_25035,N_25182);
xor U25404 (N_25404,N_24919,N_25003);
nand U25405 (N_25405,N_24964,N_25007);
nor U25406 (N_25406,N_25077,N_25036);
and U25407 (N_25407,N_24956,N_24981);
nor U25408 (N_25408,N_25184,N_24917);
and U25409 (N_25409,N_24928,N_25070);
xnor U25410 (N_25410,N_24934,N_25007);
and U25411 (N_25411,N_25197,N_25114);
nor U25412 (N_25412,N_24985,N_25086);
or U25413 (N_25413,N_25101,N_25147);
and U25414 (N_25414,N_25075,N_25034);
xor U25415 (N_25415,N_25188,N_24946);
or U25416 (N_25416,N_25194,N_25001);
xor U25417 (N_25417,N_25083,N_24940);
xnor U25418 (N_25418,N_24924,N_25068);
and U25419 (N_25419,N_25014,N_25091);
xnor U25420 (N_25420,N_25056,N_25094);
nor U25421 (N_25421,N_25107,N_25082);
or U25422 (N_25422,N_25134,N_25178);
nand U25423 (N_25423,N_25063,N_25139);
nand U25424 (N_25424,N_25154,N_24995);
nor U25425 (N_25425,N_25098,N_25011);
or U25426 (N_25426,N_24907,N_25072);
and U25427 (N_25427,N_25032,N_24992);
nand U25428 (N_25428,N_25196,N_25178);
nand U25429 (N_25429,N_25111,N_25193);
xor U25430 (N_25430,N_24901,N_24921);
nand U25431 (N_25431,N_25138,N_24936);
or U25432 (N_25432,N_25110,N_24953);
or U25433 (N_25433,N_24976,N_25095);
and U25434 (N_25434,N_24932,N_24908);
xor U25435 (N_25435,N_24945,N_25031);
xor U25436 (N_25436,N_24904,N_25094);
nor U25437 (N_25437,N_25032,N_24909);
xor U25438 (N_25438,N_25153,N_24972);
xnor U25439 (N_25439,N_25022,N_24903);
or U25440 (N_25440,N_24997,N_25128);
nor U25441 (N_25441,N_25048,N_24960);
xor U25442 (N_25442,N_25142,N_25024);
and U25443 (N_25443,N_25141,N_25132);
xor U25444 (N_25444,N_25049,N_25115);
nor U25445 (N_25445,N_24926,N_25137);
or U25446 (N_25446,N_24900,N_25009);
xor U25447 (N_25447,N_25149,N_25186);
xnor U25448 (N_25448,N_25150,N_25028);
nor U25449 (N_25449,N_25092,N_25151);
or U25450 (N_25450,N_24914,N_25031);
or U25451 (N_25451,N_25176,N_24970);
xnor U25452 (N_25452,N_25154,N_25198);
nor U25453 (N_25453,N_25170,N_24988);
and U25454 (N_25454,N_24949,N_24997);
nand U25455 (N_25455,N_25107,N_25159);
and U25456 (N_25456,N_25083,N_25149);
nor U25457 (N_25457,N_25145,N_25053);
xnor U25458 (N_25458,N_25051,N_25161);
xor U25459 (N_25459,N_24903,N_25119);
or U25460 (N_25460,N_25148,N_24923);
or U25461 (N_25461,N_24970,N_25030);
nand U25462 (N_25462,N_25036,N_24905);
nand U25463 (N_25463,N_24968,N_24996);
xnor U25464 (N_25464,N_25066,N_25182);
nor U25465 (N_25465,N_25160,N_24920);
xnor U25466 (N_25466,N_25079,N_25162);
xnor U25467 (N_25467,N_25105,N_24948);
and U25468 (N_25468,N_25130,N_25185);
or U25469 (N_25469,N_24946,N_25023);
nor U25470 (N_25470,N_25056,N_25083);
nand U25471 (N_25471,N_24907,N_25124);
nand U25472 (N_25472,N_25057,N_25030);
nand U25473 (N_25473,N_25111,N_24920);
and U25474 (N_25474,N_25013,N_25008);
and U25475 (N_25475,N_24963,N_25187);
and U25476 (N_25476,N_25148,N_24982);
nand U25477 (N_25477,N_24954,N_24924);
and U25478 (N_25478,N_25007,N_25165);
or U25479 (N_25479,N_25147,N_25031);
nor U25480 (N_25480,N_24912,N_25001);
xnor U25481 (N_25481,N_25197,N_25126);
and U25482 (N_25482,N_25198,N_25047);
and U25483 (N_25483,N_25190,N_25096);
nand U25484 (N_25484,N_25064,N_25187);
and U25485 (N_25485,N_25111,N_25073);
or U25486 (N_25486,N_25178,N_25013);
xor U25487 (N_25487,N_25141,N_25020);
xor U25488 (N_25488,N_24992,N_25061);
and U25489 (N_25489,N_25062,N_25151);
nand U25490 (N_25490,N_25112,N_25120);
nand U25491 (N_25491,N_24973,N_25037);
nor U25492 (N_25492,N_25128,N_25132);
xor U25493 (N_25493,N_25105,N_24961);
and U25494 (N_25494,N_25036,N_25005);
and U25495 (N_25495,N_25127,N_25013);
and U25496 (N_25496,N_24973,N_25103);
nand U25497 (N_25497,N_25088,N_25176);
nand U25498 (N_25498,N_24981,N_25028);
and U25499 (N_25499,N_25161,N_24907);
and U25500 (N_25500,N_25261,N_25344);
nor U25501 (N_25501,N_25346,N_25356);
and U25502 (N_25502,N_25306,N_25370);
nor U25503 (N_25503,N_25294,N_25234);
and U25504 (N_25504,N_25366,N_25478);
or U25505 (N_25505,N_25242,N_25333);
and U25506 (N_25506,N_25412,N_25498);
and U25507 (N_25507,N_25372,N_25295);
nand U25508 (N_25508,N_25482,N_25380);
and U25509 (N_25509,N_25290,N_25390);
xor U25510 (N_25510,N_25238,N_25436);
xnor U25511 (N_25511,N_25212,N_25291);
nor U25512 (N_25512,N_25236,N_25287);
nand U25513 (N_25513,N_25387,N_25357);
and U25514 (N_25514,N_25223,N_25442);
nand U25515 (N_25515,N_25447,N_25309);
nor U25516 (N_25516,N_25209,N_25389);
and U25517 (N_25517,N_25484,N_25247);
and U25518 (N_25518,N_25258,N_25456);
nor U25519 (N_25519,N_25406,N_25487);
xnor U25520 (N_25520,N_25351,N_25324);
xnor U25521 (N_25521,N_25373,N_25367);
and U25522 (N_25522,N_25248,N_25493);
nor U25523 (N_25523,N_25336,N_25231);
nand U25524 (N_25524,N_25379,N_25299);
xnor U25525 (N_25525,N_25435,N_25345);
and U25526 (N_25526,N_25264,N_25489);
or U25527 (N_25527,N_25490,N_25250);
or U25528 (N_25528,N_25292,N_25217);
nand U25529 (N_25529,N_25363,N_25414);
nor U25530 (N_25530,N_25469,N_25448);
or U25531 (N_25531,N_25471,N_25419);
or U25532 (N_25532,N_25497,N_25218);
nand U25533 (N_25533,N_25265,N_25378);
or U25534 (N_25534,N_25381,N_25303);
nand U25535 (N_25535,N_25480,N_25492);
xor U25536 (N_25536,N_25206,N_25313);
nor U25537 (N_25537,N_25252,N_25385);
or U25538 (N_25538,N_25316,N_25279);
xor U25539 (N_25539,N_25369,N_25288);
nand U25540 (N_25540,N_25340,N_25483);
nand U25541 (N_25541,N_25254,N_25266);
and U25542 (N_25542,N_25360,N_25496);
and U25543 (N_25543,N_25437,N_25410);
nand U25544 (N_25544,N_25396,N_25273);
nor U25545 (N_25545,N_25349,N_25286);
nor U25546 (N_25546,N_25225,N_25458);
or U25547 (N_25547,N_25451,N_25411);
nor U25548 (N_25548,N_25241,N_25454);
and U25549 (N_25549,N_25255,N_25439);
nor U25550 (N_25550,N_25479,N_25429);
xnor U25551 (N_25551,N_25260,N_25401);
or U25552 (N_25552,N_25335,N_25404);
nand U25553 (N_25553,N_25251,N_25315);
nor U25554 (N_25554,N_25210,N_25278);
nor U25555 (N_25555,N_25359,N_25470);
nor U25556 (N_25556,N_25276,N_25337);
or U25557 (N_25557,N_25450,N_25308);
or U25558 (N_25558,N_25394,N_25358);
xor U25559 (N_25559,N_25220,N_25243);
nor U25560 (N_25560,N_25499,N_25213);
nor U25561 (N_25561,N_25204,N_25466);
nand U25562 (N_25562,N_25481,N_25417);
nand U25563 (N_25563,N_25233,N_25216);
nor U25564 (N_25564,N_25343,N_25226);
nor U25565 (N_25565,N_25472,N_25457);
nand U25566 (N_25566,N_25432,N_25219);
nand U25567 (N_25567,N_25418,N_25215);
or U25568 (N_25568,N_25441,N_25235);
nor U25569 (N_25569,N_25269,N_25208);
nand U25570 (N_25570,N_25323,N_25334);
xor U25571 (N_25571,N_25297,N_25444);
xnor U25572 (N_25572,N_25203,N_25443);
or U25573 (N_25573,N_25326,N_25293);
nor U25574 (N_25574,N_25267,N_25377);
nor U25575 (N_25575,N_25362,N_25465);
nand U25576 (N_25576,N_25416,N_25371);
nor U25577 (N_25577,N_25259,N_25227);
nand U25578 (N_25578,N_25473,N_25398);
or U25579 (N_25579,N_25352,N_25364);
nand U25580 (N_25580,N_25329,N_25240);
nor U25581 (N_25581,N_25317,N_25397);
nand U25582 (N_25582,N_25449,N_25455);
or U25583 (N_25583,N_25228,N_25459);
nor U25584 (N_25584,N_25232,N_25301);
nor U25585 (N_25585,N_25393,N_25495);
and U25586 (N_25586,N_25423,N_25452);
nand U25587 (N_25587,N_25305,N_25403);
and U25588 (N_25588,N_25244,N_25376);
and U25589 (N_25589,N_25282,N_25318);
or U25590 (N_25590,N_25491,N_25424);
nand U25591 (N_25591,N_25440,N_25339);
nand U25592 (N_25592,N_25427,N_25270);
and U25593 (N_25593,N_25304,N_25428);
and U25594 (N_25594,N_25311,N_25374);
and U25595 (N_25595,N_25302,N_25409);
and U25596 (N_25596,N_25271,N_25361);
or U25597 (N_25597,N_25272,N_25284);
and U25598 (N_25598,N_25486,N_25201);
or U25599 (N_25599,N_25395,N_25388);
nand U25600 (N_25600,N_25268,N_25342);
xnor U25601 (N_25601,N_25474,N_25433);
nor U25602 (N_25602,N_25280,N_25296);
or U25603 (N_25603,N_25327,N_25391);
xnor U25604 (N_25604,N_25224,N_25420);
nor U25605 (N_25605,N_25462,N_25485);
nand U25606 (N_25606,N_25307,N_25475);
xnor U25607 (N_25607,N_25330,N_25365);
and U25608 (N_25608,N_25331,N_25353);
or U25609 (N_25609,N_25230,N_25319);
nand U25610 (N_25610,N_25263,N_25467);
nor U25611 (N_25611,N_25275,N_25382);
or U25612 (N_25612,N_25328,N_25256);
nor U25613 (N_25613,N_25354,N_25375);
nand U25614 (N_25614,N_25430,N_25245);
xnor U25615 (N_25615,N_25214,N_25249);
nand U25616 (N_25616,N_25383,N_25408);
and U25617 (N_25617,N_25281,N_25431);
xnor U25618 (N_25618,N_25274,N_25283);
nor U25619 (N_25619,N_25445,N_25229);
and U25620 (N_25620,N_25341,N_25314);
and U25621 (N_25621,N_25253,N_25348);
xnor U25622 (N_25622,N_25325,N_25463);
xnor U25623 (N_25623,N_25277,N_25298);
nand U25624 (N_25624,N_25392,N_25321);
and U25625 (N_25625,N_25338,N_25453);
or U25626 (N_25626,N_25421,N_25322);
or U25627 (N_25627,N_25207,N_25257);
nand U25628 (N_25628,N_25320,N_25405);
and U25629 (N_25629,N_25476,N_25221);
xor U25630 (N_25630,N_25205,N_25350);
nand U25631 (N_25631,N_25426,N_25222);
nor U25632 (N_25632,N_25425,N_25211);
and U25633 (N_25633,N_25434,N_25347);
and U25634 (N_25634,N_25285,N_25464);
and U25635 (N_25635,N_25438,N_25332);
and U25636 (N_25636,N_25460,N_25312);
or U25637 (N_25637,N_25239,N_25477);
nor U25638 (N_25638,N_25399,N_25422);
xnor U25639 (N_25639,N_25446,N_25246);
xnor U25640 (N_25640,N_25461,N_25262);
xor U25641 (N_25641,N_25402,N_25468);
nand U25642 (N_25642,N_25386,N_25488);
nand U25643 (N_25643,N_25310,N_25400);
and U25644 (N_25644,N_25415,N_25237);
and U25645 (N_25645,N_25300,N_25413);
or U25646 (N_25646,N_25407,N_25200);
or U25647 (N_25647,N_25494,N_25355);
xnor U25648 (N_25648,N_25202,N_25384);
and U25649 (N_25649,N_25289,N_25368);
nand U25650 (N_25650,N_25279,N_25452);
nand U25651 (N_25651,N_25424,N_25347);
xor U25652 (N_25652,N_25490,N_25286);
xnor U25653 (N_25653,N_25204,N_25257);
or U25654 (N_25654,N_25264,N_25267);
nor U25655 (N_25655,N_25271,N_25318);
xor U25656 (N_25656,N_25232,N_25253);
xnor U25657 (N_25657,N_25205,N_25328);
and U25658 (N_25658,N_25302,N_25444);
nand U25659 (N_25659,N_25358,N_25279);
nor U25660 (N_25660,N_25279,N_25412);
nand U25661 (N_25661,N_25204,N_25406);
or U25662 (N_25662,N_25345,N_25321);
and U25663 (N_25663,N_25303,N_25292);
or U25664 (N_25664,N_25486,N_25424);
nor U25665 (N_25665,N_25319,N_25447);
or U25666 (N_25666,N_25424,N_25373);
or U25667 (N_25667,N_25438,N_25444);
nor U25668 (N_25668,N_25350,N_25289);
nand U25669 (N_25669,N_25253,N_25228);
xnor U25670 (N_25670,N_25237,N_25477);
nor U25671 (N_25671,N_25459,N_25307);
xnor U25672 (N_25672,N_25491,N_25293);
nor U25673 (N_25673,N_25432,N_25443);
nand U25674 (N_25674,N_25489,N_25413);
nor U25675 (N_25675,N_25446,N_25220);
or U25676 (N_25676,N_25431,N_25288);
and U25677 (N_25677,N_25248,N_25386);
and U25678 (N_25678,N_25293,N_25342);
nor U25679 (N_25679,N_25402,N_25318);
xor U25680 (N_25680,N_25451,N_25430);
xor U25681 (N_25681,N_25234,N_25413);
nor U25682 (N_25682,N_25289,N_25230);
and U25683 (N_25683,N_25214,N_25283);
and U25684 (N_25684,N_25307,N_25370);
nand U25685 (N_25685,N_25401,N_25460);
or U25686 (N_25686,N_25378,N_25417);
nor U25687 (N_25687,N_25458,N_25490);
xnor U25688 (N_25688,N_25216,N_25259);
or U25689 (N_25689,N_25331,N_25325);
and U25690 (N_25690,N_25430,N_25389);
or U25691 (N_25691,N_25246,N_25258);
and U25692 (N_25692,N_25205,N_25329);
xnor U25693 (N_25693,N_25385,N_25242);
xor U25694 (N_25694,N_25419,N_25285);
xnor U25695 (N_25695,N_25355,N_25275);
nor U25696 (N_25696,N_25336,N_25404);
and U25697 (N_25697,N_25486,N_25379);
nand U25698 (N_25698,N_25382,N_25473);
nand U25699 (N_25699,N_25330,N_25429);
nand U25700 (N_25700,N_25460,N_25382);
and U25701 (N_25701,N_25492,N_25389);
nor U25702 (N_25702,N_25259,N_25410);
nor U25703 (N_25703,N_25299,N_25235);
and U25704 (N_25704,N_25319,N_25208);
nand U25705 (N_25705,N_25344,N_25214);
xnor U25706 (N_25706,N_25389,N_25343);
nand U25707 (N_25707,N_25333,N_25327);
nor U25708 (N_25708,N_25381,N_25230);
and U25709 (N_25709,N_25370,N_25496);
or U25710 (N_25710,N_25446,N_25425);
xor U25711 (N_25711,N_25354,N_25470);
nor U25712 (N_25712,N_25340,N_25273);
nor U25713 (N_25713,N_25440,N_25389);
or U25714 (N_25714,N_25221,N_25317);
or U25715 (N_25715,N_25311,N_25285);
or U25716 (N_25716,N_25271,N_25460);
or U25717 (N_25717,N_25319,N_25222);
nor U25718 (N_25718,N_25467,N_25225);
or U25719 (N_25719,N_25231,N_25205);
xnor U25720 (N_25720,N_25276,N_25404);
nor U25721 (N_25721,N_25217,N_25257);
nor U25722 (N_25722,N_25488,N_25392);
or U25723 (N_25723,N_25211,N_25204);
or U25724 (N_25724,N_25242,N_25364);
and U25725 (N_25725,N_25469,N_25490);
nor U25726 (N_25726,N_25408,N_25274);
and U25727 (N_25727,N_25348,N_25219);
nor U25728 (N_25728,N_25212,N_25230);
xnor U25729 (N_25729,N_25499,N_25254);
nand U25730 (N_25730,N_25362,N_25278);
nor U25731 (N_25731,N_25206,N_25305);
nand U25732 (N_25732,N_25419,N_25274);
nor U25733 (N_25733,N_25493,N_25470);
xnor U25734 (N_25734,N_25487,N_25447);
or U25735 (N_25735,N_25483,N_25231);
or U25736 (N_25736,N_25492,N_25242);
xnor U25737 (N_25737,N_25333,N_25399);
or U25738 (N_25738,N_25201,N_25425);
nor U25739 (N_25739,N_25331,N_25382);
nor U25740 (N_25740,N_25413,N_25269);
nand U25741 (N_25741,N_25340,N_25234);
nor U25742 (N_25742,N_25385,N_25296);
nor U25743 (N_25743,N_25400,N_25365);
or U25744 (N_25744,N_25395,N_25442);
nor U25745 (N_25745,N_25377,N_25239);
nand U25746 (N_25746,N_25209,N_25246);
or U25747 (N_25747,N_25499,N_25230);
or U25748 (N_25748,N_25344,N_25404);
xor U25749 (N_25749,N_25376,N_25299);
or U25750 (N_25750,N_25334,N_25456);
xor U25751 (N_25751,N_25291,N_25294);
nor U25752 (N_25752,N_25432,N_25416);
and U25753 (N_25753,N_25495,N_25210);
nand U25754 (N_25754,N_25222,N_25457);
nor U25755 (N_25755,N_25300,N_25287);
nor U25756 (N_25756,N_25374,N_25394);
nor U25757 (N_25757,N_25444,N_25272);
and U25758 (N_25758,N_25423,N_25257);
or U25759 (N_25759,N_25388,N_25263);
and U25760 (N_25760,N_25345,N_25229);
or U25761 (N_25761,N_25477,N_25273);
nand U25762 (N_25762,N_25410,N_25221);
or U25763 (N_25763,N_25338,N_25476);
xnor U25764 (N_25764,N_25344,N_25237);
and U25765 (N_25765,N_25443,N_25370);
nor U25766 (N_25766,N_25474,N_25381);
xnor U25767 (N_25767,N_25243,N_25434);
or U25768 (N_25768,N_25426,N_25295);
nor U25769 (N_25769,N_25322,N_25382);
xnor U25770 (N_25770,N_25277,N_25444);
nand U25771 (N_25771,N_25263,N_25221);
nor U25772 (N_25772,N_25282,N_25293);
xnor U25773 (N_25773,N_25348,N_25262);
xnor U25774 (N_25774,N_25459,N_25331);
nor U25775 (N_25775,N_25401,N_25457);
and U25776 (N_25776,N_25449,N_25274);
xnor U25777 (N_25777,N_25422,N_25465);
xnor U25778 (N_25778,N_25264,N_25469);
xnor U25779 (N_25779,N_25325,N_25295);
xnor U25780 (N_25780,N_25407,N_25460);
xnor U25781 (N_25781,N_25458,N_25349);
xnor U25782 (N_25782,N_25231,N_25208);
xnor U25783 (N_25783,N_25354,N_25211);
or U25784 (N_25784,N_25437,N_25211);
or U25785 (N_25785,N_25242,N_25233);
xor U25786 (N_25786,N_25319,N_25436);
and U25787 (N_25787,N_25396,N_25320);
nand U25788 (N_25788,N_25404,N_25257);
and U25789 (N_25789,N_25329,N_25227);
xnor U25790 (N_25790,N_25441,N_25206);
nor U25791 (N_25791,N_25424,N_25270);
and U25792 (N_25792,N_25201,N_25342);
nor U25793 (N_25793,N_25218,N_25447);
xor U25794 (N_25794,N_25459,N_25317);
nor U25795 (N_25795,N_25491,N_25227);
xnor U25796 (N_25796,N_25359,N_25355);
nand U25797 (N_25797,N_25402,N_25276);
xnor U25798 (N_25798,N_25248,N_25255);
or U25799 (N_25799,N_25217,N_25436);
or U25800 (N_25800,N_25501,N_25606);
xnor U25801 (N_25801,N_25671,N_25558);
nand U25802 (N_25802,N_25712,N_25579);
nor U25803 (N_25803,N_25667,N_25670);
xor U25804 (N_25804,N_25698,N_25769);
nand U25805 (N_25805,N_25738,N_25687);
nor U25806 (N_25806,N_25770,N_25685);
and U25807 (N_25807,N_25677,N_25648);
nor U25808 (N_25808,N_25663,N_25504);
and U25809 (N_25809,N_25506,N_25608);
and U25810 (N_25810,N_25693,N_25537);
or U25811 (N_25811,N_25597,N_25748);
xnor U25812 (N_25812,N_25633,N_25603);
nor U25813 (N_25813,N_25795,N_25510);
nand U25814 (N_25814,N_25610,N_25666);
and U25815 (N_25815,N_25621,N_25650);
nand U25816 (N_25816,N_25699,N_25594);
nand U25817 (N_25817,N_25611,N_25562);
xnor U25818 (N_25818,N_25747,N_25785);
and U25819 (N_25819,N_25742,N_25532);
xnor U25820 (N_25820,N_25707,N_25762);
nor U25821 (N_25821,N_25741,N_25798);
nor U25822 (N_25822,N_25694,N_25549);
xnor U25823 (N_25823,N_25786,N_25651);
and U25824 (N_25824,N_25753,N_25706);
nand U25825 (N_25825,N_25616,N_25787);
and U25826 (N_25826,N_25635,N_25701);
or U25827 (N_25827,N_25729,N_25727);
or U25828 (N_25828,N_25530,N_25774);
and U25829 (N_25829,N_25561,N_25593);
xor U25830 (N_25830,N_25642,N_25613);
nand U25831 (N_25831,N_25732,N_25777);
xor U25832 (N_25832,N_25797,N_25540);
and U25833 (N_25833,N_25796,N_25527);
nand U25834 (N_25834,N_25662,N_25511);
or U25835 (N_25835,N_25581,N_25719);
nor U25836 (N_25836,N_25776,N_25578);
nor U25837 (N_25837,N_25631,N_25512);
and U25838 (N_25838,N_25546,N_25690);
and U25839 (N_25839,N_25580,N_25709);
or U25840 (N_25840,N_25682,N_25627);
xnor U25841 (N_25841,N_25730,N_25592);
and U25842 (N_25842,N_25585,N_25521);
nor U25843 (N_25843,N_25559,N_25684);
nor U25844 (N_25844,N_25531,N_25615);
nor U25845 (N_25845,N_25743,N_25724);
or U25846 (N_25846,N_25636,N_25586);
and U25847 (N_25847,N_25516,N_25656);
nor U25848 (N_25848,N_25704,N_25551);
or U25849 (N_25849,N_25710,N_25756);
nor U25850 (N_25850,N_25764,N_25723);
or U25851 (N_25851,N_25788,N_25639);
and U25852 (N_25852,N_25657,N_25605);
and U25853 (N_25853,N_25523,N_25573);
xnor U25854 (N_25854,N_25507,N_25643);
and U25855 (N_25855,N_25522,N_25519);
nand U25856 (N_25856,N_25628,N_25691);
and U25857 (N_25857,N_25721,N_25761);
xnor U25858 (N_25858,N_25675,N_25536);
nor U25859 (N_25859,N_25588,N_25751);
nand U25860 (N_25860,N_25728,N_25660);
and U25861 (N_25861,N_25789,N_25508);
nor U25862 (N_25862,N_25705,N_25619);
nor U25863 (N_25863,N_25618,N_25572);
xnor U25864 (N_25864,N_25574,N_25653);
and U25865 (N_25865,N_25525,N_25524);
and U25866 (N_25866,N_25544,N_25791);
nand U25867 (N_25867,N_25543,N_25654);
xnor U25868 (N_25868,N_25604,N_25553);
nand U25869 (N_25869,N_25731,N_25718);
xnor U25870 (N_25870,N_25576,N_25645);
or U25871 (N_25871,N_25552,N_25600);
xnor U25872 (N_25872,N_25768,N_25715);
nand U25873 (N_25873,N_25735,N_25595);
nand U25874 (N_25874,N_25548,N_25711);
xor U25875 (N_25875,N_25503,N_25649);
xnor U25876 (N_25876,N_25708,N_25526);
and U25877 (N_25877,N_25695,N_25745);
or U25878 (N_25878,N_25505,N_25517);
and U25879 (N_25879,N_25793,N_25584);
or U25880 (N_25880,N_25513,N_25757);
xor U25881 (N_25881,N_25655,N_25535);
xor U25882 (N_25882,N_25620,N_25775);
xnor U25883 (N_25883,N_25583,N_25779);
and U25884 (N_25884,N_25759,N_25717);
or U25885 (N_25885,N_25577,N_25547);
nor U25886 (N_25886,N_25734,N_25533);
or U25887 (N_25887,N_25782,N_25590);
and U25888 (N_25888,N_25612,N_25567);
nand U25889 (N_25889,N_25765,N_25744);
nand U25890 (N_25890,N_25689,N_25541);
xnor U25891 (N_25891,N_25601,N_25570);
xor U25892 (N_25892,N_25638,N_25569);
xnor U25893 (N_25893,N_25542,N_25652);
nand U25894 (N_25894,N_25672,N_25599);
nand U25895 (N_25895,N_25713,N_25538);
nand U25896 (N_25896,N_25629,N_25509);
xor U25897 (N_25897,N_25784,N_25529);
or U25898 (N_25898,N_25767,N_25754);
nor U25899 (N_25899,N_25587,N_25736);
or U25900 (N_25900,N_25725,N_25700);
nor U25901 (N_25901,N_25560,N_25726);
or U25902 (N_25902,N_25591,N_25557);
and U25903 (N_25903,N_25669,N_25534);
nand U25904 (N_25904,N_25678,N_25617);
or U25905 (N_25905,N_25683,N_25539);
nor U25906 (N_25906,N_25720,N_25598);
nand U25907 (N_25907,N_25799,N_25518);
xor U25908 (N_25908,N_25686,N_25783);
or U25909 (N_25909,N_25750,N_25630);
xnor U25910 (N_25910,N_25575,N_25668);
or U25911 (N_25911,N_25520,N_25568);
and U25912 (N_25912,N_25676,N_25515);
and U25913 (N_25913,N_25647,N_25688);
or U25914 (N_25914,N_25703,N_25607);
or U25915 (N_25915,N_25740,N_25555);
and U25916 (N_25916,N_25614,N_25755);
or U25917 (N_25917,N_25737,N_25664);
nor U25918 (N_25918,N_25766,N_25564);
and U25919 (N_25919,N_25609,N_25622);
nand U25920 (N_25920,N_25771,N_25658);
and U25921 (N_25921,N_25644,N_25596);
nor U25922 (N_25922,N_25571,N_25632);
or U25923 (N_25923,N_25545,N_25665);
nor U25924 (N_25924,N_25674,N_25714);
xor U25925 (N_25925,N_25589,N_25746);
or U25926 (N_25926,N_25692,N_25556);
xnor U25927 (N_25927,N_25528,N_25763);
xnor U25928 (N_25928,N_25772,N_25697);
or U25929 (N_25929,N_25624,N_25739);
or U25930 (N_25930,N_25566,N_25500);
nor U25931 (N_25931,N_25733,N_25563);
nand U25932 (N_25932,N_25623,N_25792);
or U25933 (N_25933,N_25696,N_25582);
xnor U25934 (N_25934,N_25749,N_25758);
xnor U25935 (N_25935,N_25625,N_25550);
or U25936 (N_25936,N_25565,N_25760);
nor U25937 (N_25937,N_25646,N_25502);
nor U25938 (N_25938,N_25702,N_25514);
xor U25939 (N_25939,N_25626,N_25602);
nor U25940 (N_25940,N_25640,N_25661);
nand U25941 (N_25941,N_25679,N_25778);
xnor U25942 (N_25942,N_25780,N_25773);
nand U25943 (N_25943,N_25641,N_25659);
and U25944 (N_25944,N_25781,N_25554);
nand U25945 (N_25945,N_25752,N_25673);
nor U25946 (N_25946,N_25680,N_25716);
nand U25947 (N_25947,N_25790,N_25634);
nand U25948 (N_25948,N_25637,N_25794);
nand U25949 (N_25949,N_25681,N_25722);
nor U25950 (N_25950,N_25543,N_25622);
nand U25951 (N_25951,N_25651,N_25638);
or U25952 (N_25952,N_25765,N_25771);
or U25953 (N_25953,N_25520,N_25709);
nand U25954 (N_25954,N_25690,N_25678);
xnor U25955 (N_25955,N_25681,N_25717);
nor U25956 (N_25956,N_25694,N_25702);
or U25957 (N_25957,N_25776,N_25765);
xor U25958 (N_25958,N_25747,N_25629);
nand U25959 (N_25959,N_25637,N_25537);
xnor U25960 (N_25960,N_25739,N_25545);
and U25961 (N_25961,N_25690,N_25697);
nor U25962 (N_25962,N_25572,N_25622);
xor U25963 (N_25963,N_25725,N_25624);
nor U25964 (N_25964,N_25771,N_25527);
xnor U25965 (N_25965,N_25776,N_25740);
or U25966 (N_25966,N_25563,N_25613);
nor U25967 (N_25967,N_25670,N_25785);
and U25968 (N_25968,N_25656,N_25562);
or U25969 (N_25969,N_25775,N_25709);
nand U25970 (N_25970,N_25593,N_25580);
or U25971 (N_25971,N_25634,N_25775);
nor U25972 (N_25972,N_25696,N_25712);
xor U25973 (N_25973,N_25615,N_25644);
or U25974 (N_25974,N_25664,N_25533);
nand U25975 (N_25975,N_25527,N_25659);
and U25976 (N_25976,N_25698,N_25743);
and U25977 (N_25977,N_25545,N_25590);
nand U25978 (N_25978,N_25608,N_25513);
nand U25979 (N_25979,N_25669,N_25678);
nand U25980 (N_25980,N_25627,N_25595);
xnor U25981 (N_25981,N_25732,N_25729);
xor U25982 (N_25982,N_25651,N_25655);
nor U25983 (N_25983,N_25511,N_25731);
or U25984 (N_25984,N_25517,N_25583);
nand U25985 (N_25985,N_25698,N_25565);
and U25986 (N_25986,N_25706,N_25574);
xor U25987 (N_25987,N_25703,N_25575);
xnor U25988 (N_25988,N_25544,N_25568);
nor U25989 (N_25989,N_25544,N_25669);
xor U25990 (N_25990,N_25761,N_25612);
nor U25991 (N_25991,N_25539,N_25740);
or U25992 (N_25992,N_25620,N_25662);
and U25993 (N_25993,N_25590,N_25768);
nor U25994 (N_25994,N_25623,N_25541);
nor U25995 (N_25995,N_25770,N_25797);
and U25996 (N_25996,N_25711,N_25597);
xor U25997 (N_25997,N_25551,N_25518);
and U25998 (N_25998,N_25544,N_25770);
nand U25999 (N_25999,N_25762,N_25663);
and U26000 (N_26000,N_25588,N_25698);
and U26001 (N_26001,N_25650,N_25512);
xnor U26002 (N_26002,N_25766,N_25554);
or U26003 (N_26003,N_25515,N_25647);
and U26004 (N_26004,N_25618,N_25763);
xnor U26005 (N_26005,N_25724,N_25587);
nor U26006 (N_26006,N_25735,N_25521);
nor U26007 (N_26007,N_25517,N_25572);
nand U26008 (N_26008,N_25751,N_25766);
and U26009 (N_26009,N_25558,N_25666);
xnor U26010 (N_26010,N_25550,N_25542);
or U26011 (N_26011,N_25512,N_25692);
nand U26012 (N_26012,N_25749,N_25597);
xor U26013 (N_26013,N_25756,N_25511);
xor U26014 (N_26014,N_25786,N_25576);
or U26015 (N_26015,N_25673,N_25503);
or U26016 (N_26016,N_25794,N_25658);
or U26017 (N_26017,N_25647,N_25772);
or U26018 (N_26018,N_25653,N_25551);
nor U26019 (N_26019,N_25613,N_25661);
and U26020 (N_26020,N_25688,N_25544);
and U26021 (N_26021,N_25506,N_25661);
xnor U26022 (N_26022,N_25561,N_25560);
xor U26023 (N_26023,N_25646,N_25597);
or U26024 (N_26024,N_25649,N_25610);
xor U26025 (N_26025,N_25698,N_25653);
nand U26026 (N_26026,N_25595,N_25711);
and U26027 (N_26027,N_25615,N_25541);
xor U26028 (N_26028,N_25627,N_25641);
or U26029 (N_26029,N_25625,N_25534);
nor U26030 (N_26030,N_25614,N_25622);
nor U26031 (N_26031,N_25717,N_25691);
or U26032 (N_26032,N_25624,N_25708);
and U26033 (N_26033,N_25529,N_25770);
or U26034 (N_26034,N_25643,N_25547);
or U26035 (N_26035,N_25502,N_25674);
or U26036 (N_26036,N_25642,N_25700);
and U26037 (N_26037,N_25532,N_25766);
nor U26038 (N_26038,N_25712,N_25531);
nor U26039 (N_26039,N_25712,N_25779);
or U26040 (N_26040,N_25502,N_25622);
and U26041 (N_26041,N_25527,N_25758);
nand U26042 (N_26042,N_25694,N_25573);
nor U26043 (N_26043,N_25501,N_25519);
and U26044 (N_26044,N_25613,N_25567);
nand U26045 (N_26045,N_25660,N_25698);
and U26046 (N_26046,N_25595,N_25688);
or U26047 (N_26047,N_25694,N_25778);
nand U26048 (N_26048,N_25694,N_25506);
nand U26049 (N_26049,N_25564,N_25736);
nor U26050 (N_26050,N_25728,N_25704);
xor U26051 (N_26051,N_25697,N_25658);
and U26052 (N_26052,N_25767,N_25540);
xnor U26053 (N_26053,N_25770,N_25649);
or U26054 (N_26054,N_25650,N_25559);
nor U26055 (N_26055,N_25681,N_25672);
xor U26056 (N_26056,N_25632,N_25797);
and U26057 (N_26057,N_25718,N_25704);
and U26058 (N_26058,N_25760,N_25799);
xor U26059 (N_26059,N_25790,N_25797);
or U26060 (N_26060,N_25681,N_25668);
and U26061 (N_26061,N_25548,N_25614);
xnor U26062 (N_26062,N_25507,N_25611);
or U26063 (N_26063,N_25577,N_25502);
nand U26064 (N_26064,N_25626,N_25786);
or U26065 (N_26065,N_25650,N_25611);
and U26066 (N_26066,N_25526,N_25604);
nor U26067 (N_26067,N_25509,N_25608);
xnor U26068 (N_26068,N_25622,N_25509);
xor U26069 (N_26069,N_25518,N_25735);
or U26070 (N_26070,N_25753,N_25740);
or U26071 (N_26071,N_25762,N_25513);
or U26072 (N_26072,N_25511,N_25724);
nand U26073 (N_26073,N_25579,N_25545);
nor U26074 (N_26074,N_25533,N_25526);
and U26075 (N_26075,N_25506,N_25500);
nand U26076 (N_26076,N_25571,N_25620);
and U26077 (N_26077,N_25758,N_25563);
and U26078 (N_26078,N_25732,N_25602);
or U26079 (N_26079,N_25723,N_25684);
and U26080 (N_26080,N_25574,N_25590);
and U26081 (N_26081,N_25556,N_25529);
nor U26082 (N_26082,N_25603,N_25589);
xor U26083 (N_26083,N_25782,N_25701);
nand U26084 (N_26084,N_25503,N_25538);
or U26085 (N_26085,N_25670,N_25514);
and U26086 (N_26086,N_25705,N_25587);
nor U26087 (N_26087,N_25554,N_25686);
and U26088 (N_26088,N_25714,N_25682);
or U26089 (N_26089,N_25548,N_25736);
nor U26090 (N_26090,N_25527,N_25767);
nand U26091 (N_26091,N_25792,N_25527);
nand U26092 (N_26092,N_25597,N_25531);
nor U26093 (N_26093,N_25528,N_25571);
or U26094 (N_26094,N_25683,N_25555);
nand U26095 (N_26095,N_25752,N_25713);
nand U26096 (N_26096,N_25617,N_25657);
nand U26097 (N_26097,N_25590,N_25510);
xnor U26098 (N_26098,N_25584,N_25586);
and U26099 (N_26099,N_25736,N_25531);
or U26100 (N_26100,N_25845,N_25859);
nand U26101 (N_26101,N_25950,N_25930);
xor U26102 (N_26102,N_25963,N_26042);
nor U26103 (N_26103,N_25972,N_25957);
and U26104 (N_26104,N_25800,N_25877);
xnor U26105 (N_26105,N_25976,N_25966);
and U26106 (N_26106,N_25994,N_25843);
nor U26107 (N_26107,N_26067,N_25992);
nor U26108 (N_26108,N_26036,N_25836);
nor U26109 (N_26109,N_26069,N_25909);
nand U26110 (N_26110,N_25929,N_26028);
nor U26111 (N_26111,N_25857,N_25915);
or U26112 (N_26112,N_25871,N_25946);
nand U26113 (N_26113,N_26090,N_25886);
nor U26114 (N_26114,N_26077,N_25967);
nor U26115 (N_26115,N_26003,N_25860);
nor U26116 (N_26116,N_25823,N_26046);
xor U26117 (N_26117,N_26099,N_26006);
or U26118 (N_26118,N_25889,N_25934);
and U26119 (N_26119,N_25893,N_26068);
or U26120 (N_26120,N_25986,N_25977);
and U26121 (N_26121,N_26092,N_26001);
nor U26122 (N_26122,N_25983,N_25898);
and U26123 (N_26123,N_26014,N_25818);
or U26124 (N_26124,N_26011,N_25942);
nor U26125 (N_26125,N_26039,N_26029);
nor U26126 (N_26126,N_26071,N_25858);
xnor U26127 (N_26127,N_25959,N_26026);
or U26128 (N_26128,N_26076,N_25892);
nand U26129 (N_26129,N_25861,N_25921);
nand U26130 (N_26130,N_25901,N_26048);
nand U26131 (N_26131,N_26016,N_26096);
or U26132 (N_26132,N_25896,N_26040);
or U26133 (N_26133,N_26051,N_26019);
and U26134 (N_26134,N_26088,N_26027);
nand U26135 (N_26135,N_25989,N_25903);
and U26136 (N_26136,N_25944,N_25820);
xor U26137 (N_26137,N_25815,N_25844);
xor U26138 (N_26138,N_25951,N_26023);
xor U26139 (N_26139,N_25811,N_25936);
and U26140 (N_26140,N_25827,N_25812);
xor U26141 (N_26141,N_25801,N_26091);
and U26142 (N_26142,N_25924,N_25872);
or U26143 (N_26143,N_25945,N_25852);
nand U26144 (N_26144,N_25848,N_25943);
nor U26145 (N_26145,N_25937,N_25810);
xor U26146 (N_26146,N_26047,N_25826);
xor U26147 (N_26147,N_25825,N_25952);
xor U26148 (N_26148,N_26020,N_26044);
nor U26149 (N_26149,N_25956,N_25895);
xor U26150 (N_26150,N_25922,N_25968);
and U26151 (N_26151,N_25833,N_26097);
nor U26152 (N_26152,N_25985,N_26082);
nor U26153 (N_26153,N_25862,N_25870);
nand U26154 (N_26154,N_25980,N_26045);
xor U26155 (N_26155,N_25802,N_26010);
or U26156 (N_26156,N_25918,N_25867);
or U26157 (N_26157,N_26075,N_25856);
or U26158 (N_26158,N_25923,N_25916);
nor U26159 (N_26159,N_26030,N_25840);
xor U26160 (N_26160,N_25806,N_26033);
or U26161 (N_26161,N_25958,N_25987);
or U26162 (N_26162,N_26087,N_26064);
nor U26163 (N_26163,N_26080,N_25873);
or U26164 (N_26164,N_26083,N_25891);
and U26165 (N_26165,N_25809,N_25878);
nor U26166 (N_26166,N_25814,N_25865);
nand U26167 (N_26167,N_25965,N_25875);
xor U26168 (N_26168,N_25947,N_26066);
xnor U26169 (N_26169,N_25949,N_25854);
and U26170 (N_26170,N_25869,N_26000);
xor U26171 (N_26171,N_26086,N_26085);
nand U26172 (N_26172,N_25926,N_25970);
xor U26173 (N_26173,N_26089,N_25824);
or U26174 (N_26174,N_25851,N_26095);
nor U26175 (N_26175,N_25998,N_25997);
and U26176 (N_26176,N_25808,N_25919);
xor U26177 (N_26177,N_25908,N_25881);
and U26178 (N_26178,N_25839,N_26049);
and U26179 (N_26179,N_25971,N_25821);
and U26180 (N_26180,N_26050,N_25961);
nand U26181 (N_26181,N_25962,N_26098);
nor U26182 (N_26182,N_25828,N_26084);
or U26183 (N_26183,N_25885,N_25981);
xnor U26184 (N_26184,N_25969,N_25931);
or U26185 (N_26185,N_25855,N_26070);
nand U26186 (N_26186,N_26041,N_25803);
or U26187 (N_26187,N_25834,N_25807);
or U26188 (N_26188,N_26038,N_25991);
and U26189 (N_26189,N_25884,N_26057);
and U26190 (N_26190,N_25832,N_26035);
nor U26191 (N_26191,N_25978,N_25876);
nor U26192 (N_26192,N_25954,N_25911);
and U26193 (N_26193,N_25847,N_26094);
nor U26194 (N_26194,N_25887,N_25928);
xnor U26195 (N_26195,N_25993,N_26002);
nand U26196 (N_26196,N_25964,N_25984);
and U26197 (N_26197,N_26081,N_25842);
nand U26198 (N_26198,N_25879,N_26054);
nand U26199 (N_26199,N_25804,N_26061);
nand U26200 (N_26200,N_25831,N_25912);
and U26201 (N_26201,N_25904,N_26004);
and U26202 (N_26202,N_25973,N_26024);
nor U26203 (N_26203,N_26093,N_26032);
nor U26204 (N_26204,N_25974,N_25938);
nor U26205 (N_26205,N_25932,N_26008);
nor U26206 (N_26206,N_25910,N_25866);
nand U26207 (N_26207,N_26052,N_26063);
nor U26208 (N_26208,N_25846,N_25899);
nand U26209 (N_26209,N_25917,N_25850);
and U26210 (N_26210,N_26079,N_26007);
xnor U26211 (N_26211,N_25925,N_25888);
xnor U26212 (N_26212,N_25868,N_25953);
xnor U26213 (N_26213,N_26009,N_25913);
nor U26214 (N_26214,N_26022,N_25894);
or U26215 (N_26215,N_26012,N_25822);
and U26216 (N_26216,N_25874,N_25907);
nand U26217 (N_26217,N_26078,N_26060);
nor U26218 (N_26218,N_25960,N_25941);
nor U26219 (N_26219,N_26053,N_25920);
or U26220 (N_26220,N_26005,N_25883);
and U26221 (N_26221,N_25835,N_25819);
nor U26222 (N_26222,N_25939,N_25805);
nand U26223 (N_26223,N_25990,N_25940);
nor U26224 (N_26224,N_25882,N_26073);
nor U26225 (N_26225,N_25890,N_26034);
xnor U26226 (N_26226,N_25933,N_25841);
and U26227 (N_26227,N_25813,N_25837);
xnor U26228 (N_26228,N_26018,N_26013);
or U26229 (N_26229,N_26062,N_26017);
or U26230 (N_26230,N_25955,N_25935);
or U26231 (N_26231,N_25829,N_26037);
nand U26232 (N_26232,N_25996,N_26056);
and U26233 (N_26233,N_25906,N_26055);
and U26234 (N_26234,N_25982,N_25927);
nand U26235 (N_26235,N_26015,N_25979);
xor U26236 (N_26236,N_25864,N_25995);
xnor U26237 (N_26237,N_25816,N_25863);
or U26238 (N_26238,N_25975,N_25838);
and U26239 (N_26239,N_26025,N_25999);
xor U26240 (N_26240,N_25905,N_25830);
or U26241 (N_26241,N_26058,N_26021);
xor U26242 (N_26242,N_26043,N_25849);
xnor U26243 (N_26243,N_25897,N_25817);
or U26244 (N_26244,N_25948,N_25902);
nand U26245 (N_26245,N_25900,N_25988);
or U26246 (N_26246,N_25880,N_26059);
and U26247 (N_26247,N_26065,N_25914);
or U26248 (N_26248,N_26072,N_25853);
or U26249 (N_26249,N_26031,N_26074);
nor U26250 (N_26250,N_26052,N_25800);
xor U26251 (N_26251,N_25838,N_25822);
and U26252 (N_26252,N_25803,N_25872);
or U26253 (N_26253,N_25995,N_25984);
xnor U26254 (N_26254,N_25906,N_25936);
xor U26255 (N_26255,N_25896,N_25955);
xor U26256 (N_26256,N_26002,N_25844);
nor U26257 (N_26257,N_25894,N_26026);
nand U26258 (N_26258,N_26043,N_25977);
nand U26259 (N_26259,N_25871,N_26058);
nor U26260 (N_26260,N_25975,N_26002);
and U26261 (N_26261,N_25826,N_25892);
or U26262 (N_26262,N_26019,N_25900);
or U26263 (N_26263,N_25988,N_25911);
or U26264 (N_26264,N_25805,N_26002);
nand U26265 (N_26265,N_25904,N_25937);
nor U26266 (N_26266,N_25913,N_25914);
nand U26267 (N_26267,N_25849,N_25978);
xnor U26268 (N_26268,N_25902,N_25975);
and U26269 (N_26269,N_26099,N_25918);
or U26270 (N_26270,N_25846,N_25914);
nor U26271 (N_26271,N_26039,N_25934);
nand U26272 (N_26272,N_25923,N_26053);
and U26273 (N_26273,N_25957,N_26013);
nand U26274 (N_26274,N_26059,N_26001);
or U26275 (N_26275,N_25853,N_26092);
nand U26276 (N_26276,N_26035,N_25924);
nor U26277 (N_26277,N_25831,N_25859);
or U26278 (N_26278,N_26054,N_25990);
nor U26279 (N_26279,N_26092,N_25885);
nand U26280 (N_26280,N_25876,N_26043);
nor U26281 (N_26281,N_25918,N_25802);
nor U26282 (N_26282,N_25904,N_26094);
and U26283 (N_26283,N_25992,N_26007);
nor U26284 (N_26284,N_26048,N_26033);
nand U26285 (N_26285,N_26056,N_25912);
and U26286 (N_26286,N_26031,N_25900);
nand U26287 (N_26287,N_25972,N_25806);
or U26288 (N_26288,N_25986,N_25861);
or U26289 (N_26289,N_25882,N_25966);
nand U26290 (N_26290,N_25945,N_25825);
nor U26291 (N_26291,N_25843,N_26062);
or U26292 (N_26292,N_25980,N_25846);
and U26293 (N_26293,N_25890,N_25895);
xnor U26294 (N_26294,N_25982,N_25884);
nor U26295 (N_26295,N_25981,N_25974);
nor U26296 (N_26296,N_25976,N_26055);
or U26297 (N_26297,N_26049,N_25827);
nand U26298 (N_26298,N_25998,N_25964);
nor U26299 (N_26299,N_25953,N_26055);
and U26300 (N_26300,N_25827,N_25841);
nor U26301 (N_26301,N_25934,N_25965);
nand U26302 (N_26302,N_25962,N_25837);
nand U26303 (N_26303,N_26025,N_26090);
or U26304 (N_26304,N_25873,N_26047);
nor U26305 (N_26305,N_25882,N_25875);
nor U26306 (N_26306,N_26069,N_25965);
and U26307 (N_26307,N_25885,N_26003);
nor U26308 (N_26308,N_25822,N_25850);
xnor U26309 (N_26309,N_26002,N_25894);
nor U26310 (N_26310,N_25956,N_26078);
and U26311 (N_26311,N_25898,N_25812);
nor U26312 (N_26312,N_25954,N_25968);
and U26313 (N_26313,N_25845,N_25825);
or U26314 (N_26314,N_25963,N_26031);
and U26315 (N_26315,N_25805,N_25991);
xor U26316 (N_26316,N_26029,N_25858);
and U26317 (N_26317,N_26004,N_25908);
or U26318 (N_26318,N_25832,N_26001);
nand U26319 (N_26319,N_25839,N_25913);
or U26320 (N_26320,N_25987,N_25971);
or U26321 (N_26321,N_25979,N_25949);
or U26322 (N_26322,N_25883,N_25821);
and U26323 (N_26323,N_25974,N_26088);
or U26324 (N_26324,N_25971,N_25985);
nand U26325 (N_26325,N_25827,N_26090);
xor U26326 (N_26326,N_25939,N_25908);
xor U26327 (N_26327,N_25994,N_25965);
xor U26328 (N_26328,N_26057,N_25857);
nand U26329 (N_26329,N_25859,N_26063);
nand U26330 (N_26330,N_25861,N_25962);
or U26331 (N_26331,N_25820,N_25934);
and U26332 (N_26332,N_26060,N_26031);
xor U26333 (N_26333,N_25947,N_25988);
nand U26334 (N_26334,N_25964,N_25981);
nor U26335 (N_26335,N_26069,N_25963);
and U26336 (N_26336,N_25986,N_25965);
and U26337 (N_26337,N_25803,N_25999);
nand U26338 (N_26338,N_26010,N_26009);
and U26339 (N_26339,N_26045,N_26010);
or U26340 (N_26340,N_25836,N_26021);
or U26341 (N_26341,N_25849,N_26069);
and U26342 (N_26342,N_25841,N_26004);
nand U26343 (N_26343,N_26072,N_25882);
and U26344 (N_26344,N_26011,N_25936);
and U26345 (N_26345,N_25886,N_26005);
nor U26346 (N_26346,N_26075,N_26096);
nand U26347 (N_26347,N_25967,N_25891);
nand U26348 (N_26348,N_25810,N_25833);
or U26349 (N_26349,N_26017,N_26074);
and U26350 (N_26350,N_26072,N_25938);
nor U26351 (N_26351,N_25888,N_25840);
nor U26352 (N_26352,N_25829,N_25819);
or U26353 (N_26353,N_26059,N_25898);
nand U26354 (N_26354,N_25881,N_26025);
nor U26355 (N_26355,N_25981,N_25980);
or U26356 (N_26356,N_25880,N_26077);
and U26357 (N_26357,N_25801,N_25828);
nand U26358 (N_26358,N_25814,N_25917);
nand U26359 (N_26359,N_25855,N_25991);
and U26360 (N_26360,N_26028,N_26084);
nor U26361 (N_26361,N_25909,N_25891);
nor U26362 (N_26362,N_25944,N_26051);
or U26363 (N_26363,N_26052,N_25858);
xor U26364 (N_26364,N_25936,N_25918);
xnor U26365 (N_26365,N_25824,N_25871);
and U26366 (N_26366,N_25833,N_25983);
nor U26367 (N_26367,N_25987,N_25917);
nor U26368 (N_26368,N_26030,N_25856);
nor U26369 (N_26369,N_25969,N_26051);
nand U26370 (N_26370,N_25980,N_25919);
nand U26371 (N_26371,N_26019,N_25884);
xnor U26372 (N_26372,N_25928,N_26085);
nor U26373 (N_26373,N_25831,N_26091);
or U26374 (N_26374,N_26077,N_25837);
and U26375 (N_26375,N_26011,N_26016);
and U26376 (N_26376,N_26091,N_25856);
nand U26377 (N_26377,N_25855,N_26074);
and U26378 (N_26378,N_25801,N_26056);
and U26379 (N_26379,N_26053,N_26037);
or U26380 (N_26380,N_26054,N_25871);
or U26381 (N_26381,N_26067,N_25839);
and U26382 (N_26382,N_26072,N_25866);
nor U26383 (N_26383,N_25840,N_26028);
xnor U26384 (N_26384,N_26052,N_25886);
or U26385 (N_26385,N_26071,N_25878);
xnor U26386 (N_26386,N_26008,N_25822);
nor U26387 (N_26387,N_26075,N_26046);
xnor U26388 (N_26388,N_26098,N_26000);
and U26389 (N_26389,N_25944,N_25813);
or U26390 (N_26390,N_25810,N_25938);
nor U26391 (N_26391,N_26033,N_26000);
and U26392 (N_26392,N_25832,N_25888);
xor U26393 (N_26393,N_26017,N_25859);
nor U26394 (N_26394,N_26080,N_25968);
and U26395 (N_26395,N_25883,N_26070);
or U26396 (N_26396,N_26071,N_26085);
xnor U26397 (N_26397,N_25894,N_26054);
xor U26398 (N_26398,N_25869,N_26070);
nand U26399 (N_26399,N_26056,N_25853);
nand U26400 (N_26400,N_26282,N_26185);
and U26401 (N_26401,N_26235,N_26184);
and U26402 (N_26402,N_26112,N_26110);
xor U26403 (N_26403,N_26256,N_26115);
nand U26404 (N_26404,N_26169,N_26118);
or U26405 (N_26405,N_26365,N_26198);
xnor U26406 (N_26406,N_26250,N_26124);
nor U26407 (N_26407,N_26190,N_26237);
nand U26408 (N_26408,N_26176,N_26214);
nor U26409 (N_26409,N_26108,N_26348);
and U26410 (N_26410,N_26297,N_26173);
or U26411 (N_26411,N_26161,N_26123);
and U26412 (N_26412,N_26224,N_26276);
xnor U26413 (N_26413,N_26195,N_26130);
or U26414 (N_26414,N_26245,N_26377);
and U26415 (N_26415,N_26272,N_26391);
nor U26416 (N_26416,N_26151,N_26189);
nand U26417 (N_26417,N_26232,N_26261);
and U26418 (N_26418,N_26278,N_26229);
or U26419 (N_26419,N_26144,N_26100);
nor U26420 (N_26420,N_26322,N_26305);
nor U26421 (N_26421,N_26179,N_26273);
and U26422 (N_26422,N_26353,N_26341);
nand U26423 (N_26423,N_26139,N_26363);
or U26424 (N_26424,N_26283,N_26317);
and U26425 (N_26425,N_26394,N_26172);
or U26426 (N_26426,N_26233,N_26113);
nor U26427 (N_26427,N_26208,N_26309);
xnor U26428 (N_26428,N_26323,N_26340);
or U26429 (N_26429,N_26145,N_26399);
nand U26430 (N_26430,N_26375,N_26180);
xor U26431 (N_26431,N_26152,N_26116);
and U26432 (N_26432,N_26385,N_26114);
xnor U26433 (N_26433,N_26201,N_26243);
xor U26434 (N_26434,N_26149,N_26398);
and U26435 (N_26435,N_26390,N_26136);
nand U26436 (N_26436,N_26102,N_26327);
xor U26437 (N_26437,N_26227,N_26117);
or U26438 (N_26438,N_26131,N_26264);
xor U26439 (N_26439,N_26147,N_26247);
nand U26440 (N_26440,N_26171,N_26226);
nor U26441 (N_26441,N_26133,N_26164);
nor U26442 (N_26442,N_26339,N_26174);
or U26443 (N_26443,N_26334,N_26343);
and U26444 (N_26444,N_26397,N_26350);
or U26445 (N_26445,N_26213,N_26137);
nand U26446 (N_26446,N_26292,N_26215);
and U26447 (N_26447,N_26351,N_26298);
nor U26448 (N_26448,N_26357,N_26295);
or U26449 (N_26449,N_26335,N_26143);
and U26450 (N_26450,N_26200,N_26105);
or U26451 (N_26451,N_26236,N_26158);
and U26452 (N_26452,N_26234,N_26203);
nor U26453 (N_26453,N_26396,N_26155);
nand U26454 (N_26454,N_26177,N_26393);
nand U26455 (N_26455,N_26209,N_26382);
nand U26456 (N_26456,N_26395,N_26331);
xor U26457 (N_26457,N_26303,N_26142);
xor U26458 (N_26458,N_26175,N_26205);
nand U26459 (N_26459,N_26374,N_26355);
nand U26460 (N_26460,N_26157,N_26358);
or U26461 (N_26461,N_26128,N_26300);
or U26462 (N_26462,N_26294,N_26329);
or U26463 (N_26463,N_26153,N_26103);
nor U26464 (N_26464,N_26249,N_26378);
xor U26465 (N_26465,N_26325,N_26244);
and U26466 (N_26466,N_26321,N_26275);
xor U26467 (N_26467,N_26356,N_26231);
or U26468 (N_26468,N_26299,N_26218);
or U26469 (N_26469,N_26310,N_26333);
nor U26470 (N_26470,N_26107,N_26207);
and U26471 (N_26471,N_26217,N_26212);
xor U26472 (N_26472,N_26274,N_26251);
nand U26473 (N_26473,N_26289,N_26269);
or U26474 (N_26474,N_26266,N_26277);
xor U26475 (N_26475,N_26312,N_26220);
and U26476 (N_26476,N_26337,N_26252);
nand U26477 (N_26477,N_26210,N_26186);
xnor U26478 (N_26478,N_26165,N_26387);
and U26479 (N_26479,N_26242,N_26359);
nor U26480 (N_26480,N_26285,N_26362);
and U26481 (N_26481,N_26293,N_26265);
nor U26482 (N_26482,N_26119,N_26346);
nor U26483 (N_26483,N_26379,N_26140);
nand U26484 (N_26484,N_26354,N_26257);
xnor U26485 (N_26485,N_26349,N_26336);
and U26486 (N_26486,N_26127,N_26125);
and U26487 (N_26487,N_26302,N_26286);
nand U26488 (N_26488,N_26255,N_26246);
nor U26489 (N_26489,N_26320,N_26221);
and U26490 (N_26490,N_26366,N_26120);
or U26491 (N_26491,N_26319,N_26156);
nor U26492 (N_26492,N_26187,N_26267);
nor U26493 (N_26493,N_26216,N_26141);
or U26494 (N_26494,N_26338,N_26192);
xnor U26495 (N_26495,N_26315,N_26202);
nor U26496 (N_26496,N_26368,N_26230);
or U26497 (N_26497,N_26370,N_26388);
xnor U26498 (N_26498,N_26318,N_26330);
and U26499 (N_26499,N_26160,N_26361);
xor U26500 (N_26500,N_26225,N_26238);
xnor U26501 (N_26501,N_26268,N_26270);
and U26502 (N_26502,N_26188,N_26376);
nor U26503 (N_26503,N_26240,N_26306);
and U26504 (N_26504,N_26248,N_26109);
or U26505 (N_26505,N_26367,N_26287);
nand U26506 (N_26506,N_26347,N_26260);
xnor U26507 (N_26507,N_26206,N_26219);
or U26508 (N_26508,N_26148,N_26223);
nor U26509 (N_26509,N_26284,N_26181);
nand U26510 (N_26510,N_26162,N_26360);
nor U26511 (N_26511,N_26288,N_26163);
or U26512 (N_26512,N_26134,N_26182);
nor U26513 (N_26513,N_26371,N_26352);
and U26514 (N_26514,N_26138,N_26191);
nand U26515 (N_26515,N_26121,N_26239);
nand U26516 (N_26516,N_26381,N_26183);
nor U26517 (N_26517,N_26369,N_26228);
xnor U26518 (N_26518,N_26263,N_26146);
nor U26519 (N_26519,N_26386,N_26222);
or U26520 (N_26520,N_26178,N_26258);
or U26521 (N_26521,N_26159,N_26328);
nor U26522 (N_26522,N_26332,N_26392);
xor U26523 (N_26523,N_26101,N_26106);
nor U26524 (N_26524,N_26129,N_26262);
and U26525 (N_26525,N_26167,N_26154);
xor U26526 (N_26526,N_26308,N_26166);
or U26527 (N_26527,N_26307,N_26104);
nand U26528 (N_26528,N_26345,N_26170);
nor U26529 (N_26529,N_26150,N_26326);
nor U26530 (N_26530,N_26314,N_26290);
and U26531 (N_26531,N_26193,N_26122);
and U26532 (N_26532,N_26241,N_26311);
and U26533 (N_26533,N_26279,N_26194);
or U26534 (N_26534,N_26111,N_26364);
xnor U26535 (N_26535,N_26126,N_26253);
nor U26536 (N_26536,N_26254,N_26296);
nand U26537 (N_26537,N_26384,N_26383);
or U26538 (N_26538,N_26304,N_26373);
and U26539 (N_26539,N_26316,N_26168);
xnor U26540 (N_26540,N_26281,N_26301);
nor U26541 (N_26541,N_26132,N_26380);
or U26542 (N_26542,N_26344,N_26259);
nor U26543 (N_26543,N_26372,N_26324);
nand U26544 (N_26544,N_26204,N_26389);
xnor U26545 (N_26545,N_26342,N_26280);
or U26546 (N_26546,N_26199,N_26313);
nor U26547 (N_26547,N_26291,N_26196);
or U26548 (N_26548,N_26211,N_26135);
or U26549 (N_26549,N_26271,N_26197);
nand U26550 (N_26550,N_26140,N_26221);
or U26551 (N_26551,N_26234,N_26102);
and U26552 (N_26552,N_26278,N_26163);
nand U26553 (N_26553,N_26165,N_26105);
and U26554 (N_26554,N_26280,N_26388);
xor U26555 (N_26555,N_26367,N_26319);
and U26556 (N_26556,N_26144,N_26102);
nand U26557 (N_26557,N_26132,N_26178);
and U26558 (N_26558,N_26241,N_26182);
nand U26559 (N_26559,N_26248,N_26133);
nor U26560 (N_26560,N_26395,N_26359);
and U26561 (N_26561,N_26398,N_26289);
nor U26562 (N_26562,N_26199,N_26393);
and U26563 (N_26563,N_26192,N_26335);
nor U26564 (N_26564,N_26121,N_26118);
and U26565 (N_26565,N_26266,N_26155);
or U26566 (N_26566,N_26160,N_26177);
xnor U26567 (N_26567,N_26198,N_26298);
nor U26568 (N_26568,N_26108,N_26174);
or U26569 (N_26569,N_26253,N_26233);
nand U26570 (N_26570,N_26105,N_26152);
nor U26571 (N_26571,N_26372,N_26329);
or U26572 (N_26572,N_26102,N_26389);
or U26573 (N_26573,N_26318,N_26345);
xnor U26574 (N_26574,N_26390,N_26361);
nand U26575 (N_26575,N_26173,N_26352);
xor U26576 (N_26576,N_26249,N_26365);
nor U26577 (N_26577,N_26314,N_26100);
xor U26578 (N_26578,N_26369,N_26336);
or U26579 (N_26579,N_26241,N_26396);
nor U26580 (N_26580,N_26261,N_26268);
or U26581 (N_26581,N_26356,N_26258);
nand U26582 (N_26582,N_26337,N_26393);
and U26583 (N_26583,N_26110,N_26239);
xnor U26584 (N_26584,N_26287,N_26185);
xor U26585 (N_26585,N_26155,N_26337);
nor U26586 (N_26586,N_26371,N_26222);
nor U26587 (N_26587,N_26316,N_26376);
nor U26588 (N_26588,N_26230,N_26388);
or U26589 (N_26589,N_26101,N_26228);
or U26590 (N_26590,N_26121,N_26360);
xnor U26591 (N_26591,N_26326,N_26169);
nor U26592 (N_26592,N_26286,N_26208);
or U26593 (N_26593,N_26269,N_26139);
nor U26594 (N_26594,N_26171,N_26222);
or U26595 (N_26595,N_26151,N_26341);
nor U26596 (N_26596,N_26144,N_26307);
nor U26597 (N_26597,N_26218,N_26267);
xor U26598 (N_26598,N_26173,N_26121);
nand U26599 (N_26599,N_26158,N_26126);
nor U26600 (N_26600,N_26317,N_26115);
or U26601 (N_26601,N_26383,N_26304);
and U26602 (N_26602,N_26116,N_26233);
nor U26603 (N_26603,N_26260,N_26382);
and U26604 (N_26604,N_26301,N_26119);
and U26605 (N_26605,N_26201,N_26306);
nor U26606 (N_26606,N_26170,N_26396);
xor U26607 (N_26607,N_26114,N_26164);
nor U26608 (N_26608,N_26370,N_26220);
xnor U26609 (N_26609,N_26278,N_26333);
nand U26610 (N_26610,N_26328,N_26129);
and U26611 (N_26611,N_26103,N_26213);
xnor U26612 (N_26612,N_26113,N_26267);
nand U26613 (N_26613,N_26246,N_26140);
nand U26614 (N_26614,N_26340,N_26261);
nand U26615 (N_26615,N_26169,N_26340);
xor U26616 (N_26616,N_26300,N_26117);
or U26617 (N_26617,N_26342,N_26320);
and U26618 (N_26618,N_26311,N_26320);
nand U26619 (N_26619,N_26339,N_26230);
and U26620 (N_26620,N_26339,N_26335);
nand U26621 (N_26621,N_26393,N_26249);
or U26622 (N_26622,N_26292,N_26157);
or U26623 (N_26623,N_26284,N_26354);
or U26624 (N_26624,N_26200,N_26248);
xor U26625 (N_26625,N_26223,N_26162);
and U26626 (N_26626,N_26365,N_26209);
nand U26627 (N_26627,N_26254,N_26115);
nand U26628 (N_26628,N_26367,N_26120);
or U26629 (N_26629,N_26154,N_26156);
xnor U26630 (N_26630,N_26291,N_26188);
or U26631 (N_26631,N_26365,N_26199);
and U26632 (N_26632,N_26177,N_26399);
nand U26633 (N_26633,N_26260,N_26231);
xnor U26634 (N_26634,N_26319,N_26295);
nand U26635 (N_26635,N_26151,N_26313);
nand U26636 (N_26636,N_26171,N_26284);
or U26637 (N_26637,N_26398,N_26272);
or U26638 (N_26638,N_26304,N_26347);
nand U26639 (N_26639,N_26134,N_26160);
and U26640 (N_26640,N_26231,N_26250);
nor U26641 (N_26641,N_26344,N_26151);
and U26642 (N_26642,N_26329,N_26269);
xnor U26643 (N_26643,N_26287,N_26330);
and U26644 (N_26644,N_26182,N_26323);
or U26645 (N_26645,N_26238,N_26273);
xor U26646 (N_26646,N_26195,N_26174);
xnor U26647 (N_26647,N_26199,N_26218);
nand U26648 (N_26648,N_26324,N_26178);
and U26649 (N_26649,N_26261,N_26285);
nand U26650 (N_26650,N_26202,N_26163);
xnor U26651 (N_26651,N_26388,N_26281);
xnor U26652 (N_26652,N_26283,N_26301);
nor U26653 (N_26653,N_26146,N_26347);
or U26654 (N_26654,N_26203,N_26312);
and U26655 (N_26655,N_26228,N_26207);
and U26656 (N_26656,N_26333,N_26350);
xnor U26657 (N_26657,N_26227,N_26310);
or U26658 (N_26658,N_26196,N_26241);
xnor U26659 (N_26659,N_26199,N_26175);
and U26660 (N_26660,N_26193,N_26221);
nor U26661 (N_26661,N_26182,N_26385);
xor U26662 (N_26662,N_26212,N_26353);
and U26663 (N_26663,N_26130,N_26206);
and U26664 (N_26664,N_26222,N_26370);
nor U26665 (N_26665,N_26322,N_26287);
xor U26666 (N_26666,N_26223,N_26164);
and U26667 (N_26667,N_26241,N_26294);
or U26668 (N_26668,N_26345,N_26218);
and U26669 (N_26669,N_26236,N_26205);
nor U26670 (N_26670,N_26138,N_26381);
xor U26671 (N_26671,N_26187,N_26116);
nand U26672 (N_26672,N_26355,N_26397);
nand U26673 (N_26673,N_26263,N_26355);
xnor U26674 (N_26674,N_26171,N_26325);
xor U26675 (N_26675,N_26261,N_26381);
and U26676 (N_26676,N_26319,N_26288);
or U26677 (N_26677,N_26320,N_26137);
nor U26678 (N_26678,N_26362,N_26327);
and U26679 (N_26679,N_26295,N_26190);
nand U26680 (N_26680,N_26210,N_26389);
nor U26681 (N_26681,N_26363,N_26275);
and U26682 (N_26682,N_26392,N_26139);
or U26683 (N_26683,N_26236,N_26263);
nor U26684 (N_26684,N_26156,N_26245);
nor U26685 (N_26685,N_26283,N_26219);
and U26686 (N_26686,N_26129,N_26161);
and U26687 (N_26687,N_26193,N_26130);
and U26688 (N_26688,N_26270,N_26224);
and U26689 (N_26689,N_26163,N_26256);
and U26690 (N_26690,N_26239,N_26267);
or U26691 (N_26691,N_26134,N_26179);
xnor U26692 (N_26692,N_26258,N_26260);
and U26693 (N_26693,N_26276,N_26304);
nand U26694 (N_26694,N_26372,N_26240);
nand U26695 (N_26695,N_26312,N_26211);
or U26696 (N_26696,N_26168,N_26195);
or U26697 (N_26697,N_26158,N_26293);
nand U26698 (N_26698,N_26105,N_26340);
and U26699 (N_26699,N_26377,N_26179);
nor U26700 (N_26700,N_26687,N_26523);
nand U26701 (N_26701,N_26453,N_26405);
xnor U26702 (N_26702,N_26494,N_26509);
and U26703 (N_26703,N_26467,N_26540);
or U26704 (N_26704,N_26518,N_26586);
and U26705 (N_26705,N_26526,N_26555);
nand U26706 (N_26706,N_26628,N_26525);
nor U26707 (N_26707,N_26570,N_26412);
nor U26708 (N_26708,N_26419,N_26591);
nor U26709 (N_26709,N_26432,N_26473);
nor U26710 (N_26710,N_26476,N_26444);
xor U26711 (N_26711,N_26692,N_26638);
or U26712 (N_26712,N_26534,N_26440);
nand U26713 (N_26713,N_26533,N_26679);
nand U26714 (N_26714,N_26451,N_26578);
xnor U26715 (N_26715,N_26513,N_26436);
nor U26716 (N_26716,N_26481,N_26546);
nor U26717 (N_26717,N_26668,N_26404);
and U26718 (N_26718,N_26437,N_26439);
xor U26719 (N_26719,N_26564,N_26684);
xor U26720 (N_26720,N_26625,N_26532);
and U26721 (N_26721,N_26423,N_26401);
nand U26722 (N_26722,N_26461,N_26593);
nand U26723 (N_26723,N_26511,N_26415);
or U26724 (N_26724,N_26561,N_26619);
nor U26725 (N_26725,N_26448,N_26601);
nand U26726 (N_26726,N_26411,N_26633);
xor U26727 (N_26727,N_26691,N_26568);
or U26728 (N_26728,N_26611,N_26403);
and U26729 (N_26729,N_26592,N_26636);
xnor U26730 (N_26730,N_26562,N_26400);
nor U26731 (N_26731,N_26535,N_26589);
xnor U26732 (N_26732,N_26531,N_26681);
xnor U26733 (N_26733,N_26567,N_26604);
nand U26734 (N_26734,N_26580,N_26699);
xnor U26735 (N_26735,N_26641,N_26514);
or U26736 (N_26736,N_26443,N_26522);
nand U26737 (N_26737,N_26563,N_26541);
nor U26738 (N_26738,N_26459,N_26651);
nand U26739 (N_26739,N_26414,N_26677);
xnor U26740 (N_26740,N_26682,N_26410);
xnor U26741 (N_26741,N_26585,N_26474);
nor U26742 (N_26742,N_26630,N_26462);
and U26743 (N_26743,N_26507,N_26635);
xor U26744 (N_26744,N_26445,N_26458);
and U26745 (N_26745,N_26502,N_26538);
xor U26746 (N_26746,N_26623,N_26571);
and U26747 (N_26747,N_26560,N_26676);
nor U26748 (N_26748,N_26551,N_26698);
and U26749 (N_26749,N_26663,N_26433);
nor U26750 (N_26750,N_26618,N_26613);
xor U26751 (N_26751,N_26552,N_26637);
and U26752 (N_26752,N_26504,N_26421);
or U26753 (N_26753,N_26470,N_26446);
or U26754 (N_26754,N_26420,N_26626);
and U26755 (N_26755,N_26598,N_26639);
or U26756 (N_26756,N_26424,N_26671);
nor U26757 (N_26757,N_26683,N_26644);
and U26758 (N_26758,N_26491,N_26457);
xnor U26759 (N_26759,N_26550,N_26498);
xor U26760 (N_26760,N_26631,N_26452);
nand U26761 (N_26761,N_26643,N_26442);
xor U26762 (N_26762,N_26553,N_26664);
or U26763 (N_26763,N_26670,N_26483);
and U26764 (N_26764,N_26480,N_26594);
nor U26765 (N_26765,N_26455,N_26587);
and U26766 (N_26766,N_26500,N_26646);
nand U26767 (N_26767,N_26603,N_26431);
nor U26768 (N_26768,N_26556,N_26475);
and U26769 (N_26769,N_26557,N_26621);
xnor U26770 (N_26770,N_26501,N_26554);
or U26771 (N_26771,N_26599,N_26487);
and U26772 (N_26772,N_26666,N_26524);
or U26773 (N_26773,N_26549,N_26482);
and U26774 (N_26774,N_26427,N_26669);
xor U26775 (N_26775,N_26607,N_26629);
xnor U26776 (N_26776,N_26672,N_26655);
nor U26777 (N_26777,N_26545,N_26409);
nand U26778 (N_26778,N_26581,N_26678);
or U26779 (N_26779,N_26417,N_26688);
nor U26780 (N_26780,N_26624,N_26649);
nand U26781 (N_26781,N_26584,N_26573);
or U26782 (N_26782,N_26430,N_26695);
xnor U26783 (N_26783,N_26460,N_26620);
nand U26784 (N_26784,N_26582,N_26579);
xor U26785 (N_26785,N_26503,N_26429);
or U26786 (N_26786,N_26450,N_26685);
or U26787 (N_26787,N_26558,N_26542);
nor U26788 (N_26788,N_26616,N_26686);
or U26789 (N_26789,N_26612,N_26539);
xor U26790 (N_26790,N_26577,N_26590);
nand U26791 (N_26791,N_26499,N_26661);
or U26792 (N_26792,N_26657,N_26529);
or U26793 (N_26793,N_26466,N_26426);
nand U26794 (N_26794,N_26527,N_26662);
and U26795 (N_26795,N_26454,N_26696);
xor U26796 (N_26796,N_26456,N_26548);
nor U26797 (N_26797,N_26674,N_26615);
nand U26798 (N_26798,N_26627,N_26441);
nand U26799 (N_26799,N_26510,N_26485);
xnor U26800 (N_26800,N_26469,N_26600);
nor U26801 (N_26801,N_26428,N_26537);
and U26802 (N_26802,N_26596,N_26413);
nand U26803 (N_26803,N_26640,N_26543);
xnor U26804 (N_26804,N_26647,N_26680);
or U26805 (N_26805,N_26508,N_26665);
and U26806 (N_26806,N_26516,N_26574);
xor U26807 (N_26807,N_26425,N_26667);
or U26808 (N_26808,N_26653,N_26402);
nand U26809 (N_26809,N_26536,N_26468);
or U26810 (N_26810,N_26505,N_26506);
nor U26811 (N_26811,N_26464,N_26634);
nor U26812 (N_26812,N_26658,N_26659);
xnor U26813 (N_26813,N_26471,N_26478);
or U26814 (N_26814,N_26654,N_26407);
and U26815 (N_26815,N_26608,N_26477);
and U26816 (N_26816,N_26694,N_26689);
nor U26817 (N_26817,N_26486,N_26521);
nor U26818 (N_26818,N_26673,N_26632);
xor U26819 (N_26819,N_26416,N_26463);
or U26820 (N_26820,N_26434,N_26675);
or U26821 (N_26821,N_26490,N_26575);
nand U26822 (N_26822,N_26496,N_26489);
or U26823 (N_26823,N_26544,N_26572);
nand U26824 (N_26824,N_26565,N_26530);
nor U26825 (N_26825,N_26614,N_26656);
nor U26826 (N_26826,N_26660,N_26610);
nor U26827 (N_26827,N_26418,N_26652);
or U26828 (N_26828,N_26488,N_26492);
xnor U26829 (N_26829,N_26472,N_26605);
and U26830 (N_26830,N_26449,N_26566);
nor U26831 (N_26831,N_26645,N_26497);
nor U26832 (N_26832,N_26609,N_26493);
nor U26833 (N_26833,N_26693,N_26447);
or U26834 (N_26834,N_26622,N_26406);
or U26835 (N_26835,N_26479,N_26648);
and U26836 (N_26836,N_26617,N_26602);
xnor U26837 (N_26837,N_26465,N_26595);
nand U26838 (N_26838,N_26512,N_26520);
nand U26839 (N_26839,N_26422,N_26408);
xnor U26840 (N_26840,N_26495,N_26519);
and U26841 (N_26841,N_26597,N_26547);
or U26842 (N_26842,N_26569,N_26697);
nand U26843 (N_26843,N_26642,N_26588);
nor U26844 (N_26844,N_26515,N_26606);
nor U26845 (N_26845,N_26559,N_26435);
and U26846 (N_26846,N_26690,N_26528);
nand U26847 (N_26847,N_26517,N_26484);
nor U26848 (N_26848,N_26576,N_26650);
xor U26849 (N_26849,N_26583,N_26438);
xor U26850 (N_26850,N_26586,N_26587);
and U26851 (N_26851,N_26480,N_26648);
or U26852 (N_26852,N_26562,N_26565);
nand U26853 (N_26853,N_26442,N_26530);
or U26854 (N_26854,N_26538,N_26677);
nand U26855 (N_26855,N_26693,N_26474);
nand U26856 (N_26856,N_26446,N_26488);
xnor U26857 (N_26857,N_26657,N_26568);
or U26858 (N_26858,N_26498,N_26438);
xnor U26859 (N_26859,N_26496,N_26531);
nand U26860 (N_26860,N_26539,N_26672);
nor U26861 (N_26861,N_26658,N_26687);
xnor U26862 (N_26862,N_26633,N_26475);
or U26863 (N_26863,N_26684,N_26438);
xnor U26864 (N_26864,N_26617,N_26595);
and U26865 (N_26865,N_26409,N_26668);
and U26866 (N_26866,N_26672,N_26586);
and U26867 (N_26867,N_26545,N_26445);
nor U26868 (N_26868,N_26539,N_26685);
and U26869 (N_26869,N_26530,N_26459);
and U26870 (N_26870,N_26404,N_26484);
or U26871 (N_26871,N_26550,N_26615);
xor U26872 (N_26872,N_26413,N_26517);
xnor U26873 (N_26873,N_26664,N_26411);
or U26874 (N_26874,N_26699,N_26483);
nor U26875 (N_26875,N_26630,N_26422);
xnor U26876 (N_26876,N_26473,N_26560);
or U26877 (N_26877,N_26536,N_26652);
or U26878 (N_26878,N_26643,N_26422);
xor U26879 (N_26879,N_26596,N_26564);
xor U26880 (N_26880,N_26568,N_26674);
nand U26881 (N_26881,N_26415,N_26612);
and U26882 (N_26882,N_26553,N_26691);
xor U26883 (N_26883,N_26480,N_26460);
nand U26884 (N_26884,N_26625,N_26527);
nand U26885 (N_26885,N_26500,N_26415);
xor U26886 (N_26886,N_26591,N_26663);
nand U26887 (N_26887,N_26565,N_26688);
xnor U26888 (N_26888,N_26699,N_26464);
nand U26889 (N_26889,N_26693,N_26642);
nor U26890 (N_26890,N_26600,N_26655);
xnor U26891 (N_26891,N_26442,N_26421);
or U26892 (N_26892,N_26636,N_26639);
nand U26893 (N_26893,N_26402,N_26622);
nand U26894 (N_26894,N_26685,N_26574);
xnor U26895 (N_26895,N_26500,N_26688);
or U26896 (N_26896,N_26563,N_26502);
xnor U26897 (N_26897,N_26451,N_26666);
nand U26898 (N_26898,N_26449,N_26593);
xor U26899 (N_26899,N_26534,N_26564);
nor U26900 (N_26900,N_26446,N_26468);
xnor U26901 (N_26901,N_26640,N_26686);
nand U26902 (N_26902,N_26512,N_26629);
nor U26903 (N_26903,N_26668,N_26511);
and U26904 (N_26904,N_26422,N_26567);
nand U26905 (N_26905,N_26595,N_26462);
nor U26906 (N_26906,N_26653,N_26515);
or U26907 (N_26907,N_26563,N_26509);
or U26908 (N_26908,N_26481,N_26530);
or U26909 (N_26909,N_26622,N_26573);
nand U26910 (N_26910,N_26463,N_26625);
nor U26911 (N_26911,N_26613,N_26611);
or U26912 (N_26912,N_26698,N_26565);
xnor U26913 (N_26913,N_26592,N_26447);
nand U26914 (N_26914,N_26421,N_26498);
nor U26915 (N_26915,N_26551,N_26457);
nand U26916 (N_26916,N_26449,N_26459);
or U26917 (N_26917,N_26457,N_26558);
nand U26918 (N_26918,N_26584,N_26592);
xnor U26919 (N_26919,N_26676,N_26413);
xnor U26920 (N_26920,N_26537,N_26440);
xnor U26921 (N_26921,N_26600,N_26610);
or U26922 (N_26922,N_26583,N_26656);
xor U26923 (N_26923,N_26695,N_26525);
xor U26924 (N_26924,N_26505,N_26504);
nand U26925 (N_26925,N_26576,N_26546);
nor U26926 (N_26926,N_26671,N_26594);
or U26927 (N_26927,N_26633,N_26689);
or U26928 (N_26928,N_26583,N_26681);
and U26929 (N_26929,N_26538,N_26601);
and U26930 (N_26930,N_26655,N_26563);
or U26931 (N_26931,N_26573,N_26668);
and U26932 (N_26932,N_26686,N_26552);
or U26933 (N_26933,N_26675,N_26628);
nor U26934 (N_26934,N_26597,N_26565);
or U26935 (N_26935,N_26490,N_26662);
xor U26936 (N_26936,N_26431,N_26672);
nand U26937 (N_26937,N_26574,N_26457);
nor U26938 (N_26938,N_26585,N_26557);
xnor U26939 (N_26939,N_26680,N_26697);
xnor U26940 (N_26940,N_26644,N_26565);
or U26941 (N_26941,N_26651,N_26656);
xnor U26942 (N_26942,N_26605,N_26449);
xor U26943 (N_26943,N_26625,N_26659);
nor U26944 (N_26944,N_26654,N_26589);
or U26945 (N_26945,N_26404,N_26595);
or U26946 (N_26946,N_26532,N_26432);
and U26947 (N_26947,N_26412,N_26441);
and U26948 (N_26948,N_26599,N_26449);
nor U26949 (N_26949,N_26683,N_26651);
nand U26950 (N_26950,N_26493,N_26555);
xor U26951 (N_26951,N_26572,N_26423);
xor U26952 (N_26952,N_26693,N_26640);
and U26953 (N_26953,N_26511,N_26418);
nor U26954 (N_26954,N_26500,N_26628);
xor U26955 (N_26955,N_26699,N_26472);
xnor U26956 (N_26956,N_26682,N_26673);
and U26957 (N_26957,N_26600,N_26677);
or U26958 (N_26958,N_26474,N_26609);
nor U26959 (N_26959,N_26452,N_26471);
and U26960 (N_26960,N_26672,N_26486);
nand U26961 (N_26961,N_26603,N_26467);
nor U26962 (N_26962,N_26616,N_26456);
nand U26963 (N_26963,N_26434,N_26478);
or U26964 (N_26964,N_26511,N_26429);
nand U26965 (N_26965,N_26685,N_26557);
xor U26966 (N_26966,N_26625,N_26456);
or U26967 (N_26967,N_26586,N_26670);
and U26968 (N_26968,N_26526,N_26672);
and U26969 (N_26969,N_26536,N_26519);
nor U26970 (N_26970,N_26663,N_26661);
xnor U26971 (N_26971,N_26427,N_26588);
xnor U26972 (N_26972,N_26427,N_26481);
xor U26973 (N_26973,N_26433,N_26694);
and U26974 (N_26974,N_26522,N_26450);
and U26975 (N_26975,N_26671,N_26437);
or U26976 (N_26976,N_26486,N_26400);
xnor U26977 (N_26977,N_26696,N_26474);
nor U26978 (N_26978,N_26528,N_26480);
nor U26979 (N_26979,N_26634,N_26538);
and U26980 (N_26980,N_26410,N_26674);
and U26981 (N_26981,N_26459,N_26647);
or U26982 (N_26982,N_26566,N_26565);
nand U26983 (N_26983,N_26653,N_26610);
nand U26984 (N_26984,N_26668,N_26419);
nor U26985 (N_26985,N_26539,N_26622);
or U26986 (N_26986,N_26521,N_26628);
or U26987 (N_26987,N_26569,N_26652);
xor U26988 (N_26988,N_26480,N_26441);
or U26989 (N_26989,N_26582,N_26547);
or U26990 (N_26990,N_26602,N_26475);
nor U26991 (N_26991,N_26555,N_26659);
xor U26992 (N_26992,N_26569,N_26458);
and U26993 (N_26993,N_26426,N_26409);
nor U26994 (N_26994,N_26454,N_26574);
xor U26995 (N_26995,N_26552,N_26572);
and U26996 (N_26996,N_26611,N_26669);
xnor U26997 (N_26997,N_26546,N_26586);
xnor U26998 (N_26998,N_26401,N_26626);
xor U26999 (N_26999,N_26581,N_26419);
or U27000 (N_27000,N_26851,N_26816);
xnor U27001 (N_27001,N_26882,N_26963);
nand U27002 (N_27002,N_26973,N_26869);
nor U27003 (N_27003,N_26974,N_26806);
nand U27004 (N_27004,N_26920,N_26790);
and U27005 (N_27005,N_26709,N_26717);
nand U27006 (N_27006,N_26912,N_26944);
nor U27007 (N_27007,N_26834,N_26906);
or U27008 (N_27008,N_26899,N_26821);
and U27009 (N_27009,N_26789,N_26833);
and U27010 (N_27010,N_26783,N_26889);
or U27011 (N_27011,N_26870,N_26757);
and U27012 (N_27012,N_26811,N_26896);
nor U27013 (N_27013,N_26951,N_26764);
and U27014 (N_27014,N_26738,N_26769);
xor U27015 (N_27015,N_26865,N_26726);
nor U27016 (N_27016,N_26961,N_26955);
nor U27017 (N_27017,N_26964,N_26942);
or U27018 (N_27018,N_26732,N_26954);
or U27019 (N_27019,N_26916,N_26838);
nor U27020 (N_27020,N_26873,N_26765);
and U27021 (N_27021,N_26980,N_26815);
nor U27022 (N_27022,N_26890,N_26760);
nor U27023 (N_27023,N_26958,N_26972);
and U27024 (N_27024,N_26736,N_26953);
nand U27025 (N_27025,N_26730,N_26842);
xor U27026 (N_27026,N_26703,N_26910);
nand U27027 (N_27027,N_26802,N_26772);
nor U27028 (N_27028,N_26818,N_26728);
nor U27029 (N_27029,N_26932,N_26948);
nand U27030 (N_27030,N_26830,N_26918);
and U27031 (N_27031,N_26798,N_26771);
and U27032 (N_27032,N_26983,N_26985);
nor U27033 (N_27033,N_26844,N_26823);
nor U27034 (N_27034,N_26747,N_26863);
xor U27035 (N_27035,N_26875,N_26817);
and U27036 (N_27036,N_26744,N_26923);
xnor U27037 (N_27037,N_26734,N_26911);
or U27038 (N_27038,N_26977,N_26861);
or U27039 (N_27039,N_26839,N_26814);
and U27040 (N_27040,N_26768,N_26917);
nor U27041 (N_27041,N_26722,N_26903);
nand U27042 (N_27042,N_26957,N_26803);
nor U27043 (N_27043,N_26895,N_26724);
or U27044 (N_27044,N_26746,N_26827);
nand U27045 (N_27045,N_26813,N_26856);
nand U27046 (N_27046,N_26743,N_26849);
or U27047 (N_27047,N_26805,N_26782);
or U27048 (N_27048,N_26721,N_26763);
nand U27049 (N_27049,N_26959,N_26926);
nor U27050 (N_27050,N_26930,N_26967);
nand U27051 (N_27051,N_26779,N_26737);
xnor U27052 (N_27052,N_26919,N_26902);
and U27053 (N_27053,N_26982,N_26727);
xnor U27054 (N_27054,N_26981,N_26725);
nor U27055 (N_27055,N_26710,N_26745);
and U27056 (N_27056,N_26829,N_26800);
nand U27057 (N_27057,N_26778,N_26824);
nand U27058 (N_27058,N_26759,N_26949);
and U27059 (N_27059,N_26794,N_26872);
nor U27060 (N_27060,N_26925,N_26787);
xor U27061 (N_27061,N_26960,N_26820);
xnor U27062 (N_27062,N_26795,N_26792);
nand U27063 (N_27063,N_26975,N_26888);
and U27064 (N_27064,N_26993,N_26828);
xor U27065 (N_27065,N_26868,N_26988);
nor U27066 (N_27066,N_26892,N_26719);
or U27067 (N_27067,N_26854,N_26705);
and U27068 (N_27068,N_26773,N_26715);
and U27069 (N_27069,N_26947,N_26898);
xnor U27070 (N_27070,N_26855,N_26884);
xnor U27071 (N_27071,N_26952,N_26943);
xor U27072 (N_27072,N_26840,N_26755);
and U27073 (N_27073,N_26785,N_26996);
or U27074 (N_27074,N_26822,N_26809);
or U27075 (N_27075,N_26804,N_26843);
and U27076 (N_27076,N_26825,N_26990);
or U27077 (N_27077,N_26893,N_26720);
nor U27078 (N_27078,N_26788,N_26819);
and U27079 (N_27079,N_26994,N_26812);
and U27080 (N_27080,N_26950,N_26801);
nand U27081 (N_27081,N_26940,N_26986);
xor U27082 (N_27082,N_26756,N_26716);
and U27083 (N_27083,N_26791,N_26879);
nor U27084 (N_27084,N_26739,N_26700);
or U27085 (N_27085,N_26946,N_26810);
and U27086 (N_27086,N_26968,N_26832);
xnor U27087 (N_27087,N_26797,N_26714);
nor U27088 (N_27088,N_26987,N_26992);
and U27089 (N_27089,N_26702,N_26876);
nor U27090 (N_27090,N_26859,N_26799);
xor U27091 (N_27091,N_26729,N_26965);
nor U27092 (N_27092,N_26999,N_26853);
or U27093 (N_27093,N_26826,N_26749);
nor U27094 (N_27094,N_26924,N_26897);
nand U27095 (N_27095,N_26885,N_26862);
nor U27096 (N_27096,N_26742,N_26713);
or U27097 (N_27097,N_26984,N_26939);
xnor U27098 (N_27098,N_26945,N_26708);
nor U27099 (N_27099,N_26740,N_26780);
nor U27100 (N_27100,N_26748,N_26887);
nor U27101 (N_27101,N_26786,N_26704);
or U27102 (N_27102,N_26864,N_26793);
or U27103 (N_27103,N_26808,N_26979);
and U27104 (N_27104,N_26883,N_26845);
xnor U27105 (N_27105,N_26937,N_26762);
nand U27106 (N_27106,N_26871,N_26796);
nor U27107 (N_27107,N_26886,N_26841);
xnor U27108 (N_27108,N_26835,N_26989);
nor U27109 (N_27109,N_26978,N_26881);
xnor U27110 (N_27110,N_26877,N_26933);
or U27111 (N_27111,N_26781,N_26904);
xnor U27112 (N_27112,N_26711,N_26901);
nand U27113 (N_27113,N_26770,N_26846);
nor U27114 (N_27114,N_26733,N_26878);
and U27115 (N_27115,N_26761,N_26894);
nor U27116 (N_27116,N_26866,N_26934);
and U27117 (N_27117,N_26741,N_26712);
nand U27118 (N_27118,N_26752,N_26936);
nand U27119 (N_27119,N_26701,N_26837);
or U27120 (N_27120,N_26751,N_26836);
xor U27121 (N_27121,N_26767,N_26928);
nand U27122 (N_27122,N_26922,N_26847);
nor U27123 (N_27123,N_26867,N_26758);
and U27124 (N_27124,N_26962,N_26766);
and U27125 (N_27125,N_26754,N_26857);
xor U27126 (N_27126,N_26706,N_26874);
and U27127 (N_27127,N_26707,N_26905);
or U27128 (N_27128,N_26900,N_26731);
nor U27129 (N_27129,N_26921,N_26907);
xnor U27130 (N_27130,N_26929,N_26880);
or U27131 (N_27131,N_26775,N_26753);
nand U27132 (N_27132,N_26831,N_26850);
nor U27133 (N_27133,N_26848,N_26718);
or U27134 (N_27134,N_26935,N_26941);
and U27135 (N_27135,N_26777,N_26969);
xnor U27136 (N_27136,N_26971,N_26860);
xor U27137 (N_27137,N_26852,N_26914);
or U27138 (N_27138,N_26909,N_26966);
and U27139 (N_27139,N_26998,N_26970);
and U27140 (N_27140,N_26997,N_26931);
nor U27141 (N_27141,N_26807,N_26891);
xnor U27142 (N_27142,N_26938,N_26995);
and U27143 (N_27143,N_26991,N_26913);
and U27144 (N_27144,N_26723,N_26976);
nand U27145 (N_27145,N_26908,N_26776);
nor U27146 (N_27146,N_26784,N_26735);
or U27147 (N_27147,N_26915,N_26956);
nor U27148 (N_27148,N_26858,N_26927);
or U27149 (N_27149,N_26750,N_26774);
nor U27150 (N_27150,N_26994,N_26711);
nand U27151 (N_27151,N_26824,N_26962);
or U27152 (N_27152,N_26959,N_26887);
and U27153 (N_27153,N_26990,N_26961);
nand U27154 (N_27154,N_26833,N_26830);
xnor U27155 (N_27155,N_26950,N_26848);
xor U27156 (N_27156,N_26932,N_26703);
or U27157 (N_27157,N_26726,N_26802);
or U27158 (N_27158,N_26972,N_26973);
nand U27159 (N_27159,N_26971,N_26881);
xnor U27160 (N_27160,N_26738,N_26984);
nor U27161 (N_27161,N_26797,N_26889);
nand U27162 (N_27162,N_26798,N_26961);
or U27163 (N_27163,N_26952,N_26868);
or U27164 (N_27164,N_26936,N_26946);
and U27165 (N_27165,N_26867,N_26791);
xor U27166 (N_27166,N_26937,N_26739);
nand U27167 (N_27167,N_26736,N_26847);
nor U27168 (N_27168,N_26869,N_26979);
or U27169 (N_27169,N_26934,N_26923);
xor U27170 (N_27170,N_26718,N_26808);
nand U27171 (N_27171,N_26885,N_26777);
nand U27172 (N_27172,N_26739,N_26864);
nand U27173 (N_27173,N_26946,N_26805);
or U27174 (N_27174,N_26720,N_26908);
and U27175 (N_27175,N_26924,N_26986);
or U27176 (N_27176,N_26986,N_26952);
or U27177 (N_27177,N_26792,N_26789);
nor U27178 (N_27178,N_26980,N_26782);
xor U27179 (N_27179,N_26706,N_26825);
or U27180 (N_27180,N_26703,N_26960);
xor U27181 (N_27181,N_26766,N_26740);
nor U27182 (N_27182,N_26725,N_26977);
and U27183 (N_27183,N_26950,N_26904);
nor U27184 (N_27184,N_26728,N_26891);
nor U27185 (N_27185,N_26786,N_26902);
xnor U27186 (N_27186,N_26809,N_26915);
xor U27187 (N_27187,N_26776,N_26809);
or U27188 (N_27188,N_26832,N_26900);
or U27189 (N_27189,N_26855,N_26999);
nand U27190 (N_27190,N_26807,N_26881);
nand U27191 (N_27191,N_26884,N_26804);
nand U27192 (N_27192,N_26952,N_26807);
and U27193 (N_27193,N_26931,N_26944);
nand U27194 (N_27194,N_26982,N_26767);
or U27195 (N_27195,N_26970,N_26935);
or U27196 (N_27196,N_26807,N_26862);
and U27197 (N_27197,N_26887,N_26738);
nor U27198 (N_27198,N_26992,N_26882);
nand U27199 (N_27199,N_26740,N_26890);
nand U27200 (N_27200,N_26911,N_26811);
and U27201 (N_27201,N_26806,N_26825);
and U27202 (N_27202,N_26718,N_26931);
nor U27203 (N_27203,N_26929,N_26735);
xor U27204 (N_27204,N_26998,N_26787);
nand U27205 (N_27205,N_26791,N_26892);
xnor U27206 (N_27206,N_26951,N_26964);
and U27207 (N_27207,N_26868,N_26700);
and U27208 (N_27208,N_26947,N_26866);
and U27209 (N_27209,N_26709,N_26981);
nor U27210 (N_27210,N_26904,N_26826);
and U27211 (N_27211,N_26739,N_26816);
nand U27212 (N_27212,N_26989,N_26840);
nand U27213 (N_27213,N_26707,N_26808);
nor U27214 (N_27214,N_26890,N_26850);
xnor U27215 (N_27215,N_26925,N_26956);
or U27216 (N_27216,N_26868,N_26955);
nor U27217 (N_27217,N_26742,N_26815);
or U27218 (N_27218,N_26769,N_26938);
xor U27219 (N_27219,N_26935,N_26902);
nand U27220 (N_27220,N_26940,N_26968);
xnor U27221 (N_27221,N_26923,N_26901);
nor U27222 (N_27222,N_26844,N_26963);
or U27223 (N_27223,N_26933,N_26860);
and U27224 (N_27224,N_26928,N_26830);
nor U27225 (N_27225,N_26717,N_26826);
nor U27226 (N_27226,N_26729,N_26720);
and U27227 (N_27227,N_26903,N_26732);
or U27228 (N_27228,N_26777,N_26762);
and U27229 (N_27229,N_26809,N_26804);
nor U27230 (N_27230,N_26767,N_26770);
nor U27231 (N_27231,N_26805,N_26944);
nand U27232 (N_27232,N_26989,N_26754);
nand U27233 (N_27233,N_26789,N_26806);
nor U27234 (N_27234,N_26797,N_26711);
nor U27235 (N_27235,N_26765,N_26912);
or U27236 (N_27236,N_26828,N_26997);
xnor U27237 (N_27237,N_26927,N_26897);
nand U27238 (N_27238,N_26900,N_26983);
or U27239 (N_27239,N_26856,N_26920);
or U27240 (N_27240,N_26952,N_26753);
nor U27241 (N_27241,N_26843,N_26759);
xnor U27242 (N_27242,N_26712,N_26840);
xnor U27243 (N_27243,N_26898,N_26887);
nor U27244 (N_27244,N_26994,N_26745);
nor U27245 (N_27245,N_26877,N_26863);
nand U27246 (N_27246,N_26846,N_26861);
xnor U27247 (N_27247,N_26789,N_26700);
xnor U27248 (N_27248,N_26895,N_26717);
nor U27249 (N_27249,N_26700,N_26860);
nand U27250 (N_27250,N_26923,N_26914);
nand U27251 (N_27251,N_26771,N_26945);
or U27252 (N_27252,N_26924,N_26741);
and U27253 (N_27253,N_26963,N_26990);
nor U27254 (N_27254,N_26822,N_26750);
xnor U27255 (N_27255,N_26723,N_26778);
xor U27256 (N_27256,N_26820,N_26746);
xnor U27257 (N_27257,N_26983,N_26998);
and U27258 (N_27258,N_26878,N_26746);
or U27259 (N_27259,N_26878,N_26831);
nor U27260 (N_27260,N_26985,N_26720);
or U27261 (N_27261,N_26809,N_26773);
nand U27262 (N_27262,N_26942,N_26977);
and U27263 (N_27263,N_26969,N_26860);
and U27264 (N_27264,N_26898,N_26865);
and U27265 (N_27265,N_26799,N_26870);
xnor U27266 (N_27266,N_26780,N_26926);
nor U27267 (N_27267,N_26826,N_26845);
nand U27268 (N_27268,N_26981,N_26914);
xor U27269 (N_27269,N_26792,N_26767);
xor U27270 (N_27270,N_26819,N_26984);
and U27271 (N_27271,N_26887,N_26726);
xor U27272 (N_27272,N_26981,N_26862);
nor U27273 (N_27273,N_26746,N_26976);
xnor U27274 (N_27274,N_26835,N_26759);
nand U27275 (N_27275,N_26710,N_26823);
nand U27276 (N_27276,N_26857,N_26895);
nor U27277 (N_27277,N_26727,N_26774);
and U27278 (N_27278,N_26750,N_26898);
xor U27279 (N_27279,N_26886,N_26772);
or U27280 (N_27280,N_26707,N_26765);
and U27281 (N_27281,N_26703,N_26734);
nor U27282 (N_27282,N_26960,N_26879);
and U27283 (N_27283,N_26880,N_26813);
nor U27284 (N_27284,N_26766,N_26782);
and U27285 (N_27285,N_26705,N_26910);
and U27286 (N_27286,N_26929,N_26886);
nor U27287 (N_27287,N_26947,N_26981);
and U27288 (N_27288,N_26767,N_26989);
or U27289 (N_27289,N_26826,N_26935);
nor U27290 (N_27290,N_26978,N_26817);
and U27291 (N_27291,N_26752,N_26868);
and U27292 (N_27292,N_26835,N_26701);
or U27293 (N_27293,N_26927,N_26875);
xor U27294 (N_27294,N_26874,N_26974);
and U27295 (N_27295,N_26771,N_26967);
nor U27296 (N_27296,N_26885,N_26926);
xor U27297 (N_27297,N_26970,N_26937);
and U27298 (N_27298,N_26862,N_26962);
xnor U27299 (N_27299,N_26760,N_26775);
and U27300 (N_27300,N_27039,N_27199);
or U27301 (N_27301,N_27181,N_27262);
nand U27302 (N_27302,N_27245,N_27286);
or U27303 (N_27303,N_27022,N_27281);
nand U27304 (N_27304,N_27004,N_27086);
nor U27305 (N_27305,N_27073,N_27047);
nand U27306 (N_27306,N_27146,N_27087);
or U27307 (N_27307,N_27111,N_27065);
or U27308 (N_27308,N_27099,N_27008);
and U27309 (N_27309,N_27154,N_27029);
or U27310 (N_27310,N_27200,N_27159);
nor U27311 (N_27311,N_27297,N_27057);
nand U27312 (N_27312,N_27062,N_27156);
or U27313 (N_27313,N_27220,N_27042);
xnor U27314 (N_27314,N_27189,N_27265);
xnor U27315 (N_27315,N_27107,N_27205);
and U27316 (N_27316,N_27048,N_27138);
and U27317 (N_27317,N_27270,N_27168);
nand U27318 (N_27318,N_27137,N_27150);
or U27319 (N_27319,N_27035,N_27158);
and U27320 (N_27320,N_27152,N_27006);
nor U27321 (N_27321,N_27292,N_27052);
or U27322 (N_27322,N_27080,N_27186);
nand U27323 (N_27323,N_27058,N_27216);
nand U27324 (N_27324,N_27295,N_27132);
and U27325 (N_27325,N_27142,N_27083);
or U27326 (N_27326,N_27256,N_27036);
xnor U27327 (N_27327,N_27275,N_27192);
or U27328 (N_27328,N_27153,N_27160);
xor U27329 (N_27329,N_27026,N_27155);
or U27330 (N_27330,N_27070,N_27112);
xor U27331 (N_27331,N_27088,N_27074);
and U27332 (N_27332,N_27278,N_27093);
nand U27333 (N_27333,N_27028,N_27121);
and U27334 (N_27334,N_27082,N_27248);
nand U27335 (N_27335,N_27236,N_27110);
nor U27336 (N_27336,N_27187,N_27257);
nand U27337 (N_27337,N_27225,N_27097);
nand U27338 (N_27338,N_27049,N_27218);
nor U27339 (N_27339,N_27059,N_27209);
nand U27340 (N_27340,N_27238,N_27179);
xnor U27341 (N_27341,N_27227,N_27113);
or U27342 (N_27342,N_27119,N_27207);
nor U27343 (N_27343,N_27217,N_27269);
nand U27344 (N_27344,N_27069,N_27233);
nand U27345 (N_27345,N_27244,N_27180);
xnor U27346 (N_27346,N_27274,N_27007);
or U27347 (N_27347,N_27147,N_27041);
and U27348 (N_27348,N_27287,N_27056);
xor U27349 (N_27349,N_27229,N_27260);
and U27350 (N_27350,N_27298,N_27151);
nand U27351 (N_27351,N_27118,N_27279);
nand U27352 (N_27352,N_27068,N_27096);
or U27353 (N_27353,N_27271,N_27226);
xnor U27354 (N_27354,N_27104,N_27081);
or U27355 (N_27355,N_27023,N_27296);
xnor U27356 (N_27356,N_27291,N_27050);
nor U27357 (N_27357,N_27264,N_27182);
or U27358 (N_27358,N_27173,N_27003);
and U27359 (N_27359,N_27195,N_27123);
xnor U27360 (N_27360,N_27067,N_27231);
and U27361 (N_27361,N_27024,N_27045);
xnor U27362 (N_27362,N_27253,N_27040);
or U27363 (N_27363,N_27166,N_27149);
and U27364 (N_27364,N_27183,N_27198);
xor U27365 (N_27365,N_27013,N_27066);
xnor U27366 (N_27366,N_27184,N_27239);
and U27367 (N_27367,N_27098,N_27230);
and U27368 (N_27368,N_27079,N_27090);
and U27369 (N_27369,N_27294,N_27289);
nor U27370 (N_27370,N_27208,N_27014);
nand U27371 (N_27371,N_27115,N_27011);
xnor U27372 (N_27372,N_27191,N_27176);
xor U27373 (N_27373,N_27285,N_27091);
or U27374 (N_27374,N_27135,N_27247);
nand U27375 (N_27375,N_27178,N_27078);
nor U27376 (N_27376,N_27143,N_27009);
or U27377 (N_27377,N_27054,N_27246);
or U27378 (N_27378,N_27272,N_27219);
xor U27379 (N_27379,N_27105,N_27197);
nor U27380 (N_27380,N_27202,N_27204);
nand U27381 (N_27381,N_27266,N_27157);
nand U27382 (N_27382,N_27017,N_27016);
nor U27383 (N_27383,N_27114,N_27046);
nand U27384 (N_27384,N_27134,N_27237);
nor U27385 (N_27385,N_27128,N_27224);
nand U27386 (N_27386,N_27201,N_27072);
nand U27387 (N_27387,N_27051,N_27221);
and U27388 (N_27388,N_27136,N_27234);
nand U27389 (N_27389,N_27268,N_27288);
nand U27390 (N_27390,N_27276,N_27196);
and U27391 (N_27391,N_27002,N_27232);
and U27392 (N_27392,N_27211,N_27133);
nor U27393 (N_27393,N_27139,N_27163);
or U27394 (N_27394,N_27077,N_27129);
and U27395 (N_27395,N_27188,N_27243);
nor U27396 (N_27396,N_27255,N_27190);
and U27397 (N_27397,N_27251,N_27206);
nand U27398 (N_27398,N_27053,N_27005);
or U27399 (N_27399,N_27030,N_27164);
nor U27400 (N_27400,N_27018,N_27215);
or U27401 (N_27401,N_27043,N_27259);
and U27402 (N_27402,N_27060,N_27012);
nand U27403 (N_27403,N_27092,N_27020);
or U27404 (N_27404,N_27071,N_27290);
and U27405 (N_27405,N_27293,N_27252);
nand U27406 (N_27406,N_27263,N_27027);
xor U27407 (N_27407,N_27064,N_27172);
or U27408 (N_27408,N_27075,N_27167);
nand U27409 (N_27409,N_27165,N_27241);
nor U27410 (N_27410,N_27210,N_27063);
and U27411 (N_27411,N_27015,N_27124);
xor U27412 (N_27412,N_27171,N_27108);
and U27413 (N_27413,N_27250,N_27019);
xor U27414 (N_27414,N_27001,N_27228);
xor U27415 (N_27415,N_27100,N_27185);
nand U27416 (N_27416,N_27240,N_27038);
nand U27417 (N_27417,N_27174,N_27125);
or U27418 (N_27418,N_27084,N_27130);
and U27419 (N_27419,N_27120,N_27273);
xnor U27420 (N_27420,N_27212,N_27122);
nor U27421 (N_27421,N_27094,N_27021);
or U27422 (N_27422,N_27169,N_27102);
or U27423 (N_27423,N_27076,N_27170);
or U27424 (N_27424,N_27106,N_27061);
nor U27425 (N_27425,N_27034,N_27126);
nor U27426 (N_27426,N_27235,N_27213);
nor U27427 (N_27427,N_27037,N_27280);
nor U27428 (N_27428,N_27109,N_27055);
nand U27429 (N_27429,N_27258,N_27010);
or U27430 (N_27430,N_27223,N_27161);
and U27431 (N_27431,N_27085,N_27141);
xor U27432 (N_27432,N_27162,N_27032);
or U27433 (N_27433,N_27214,N_27044);
xnor U27434 (N_27434,N_27117,N_27140);
nand U27435 (N_27435,N_27144,N_27283);
xor U27436 (N_27436,N_27175,N_27249);
nor U27437 (N_27437,N_27261,N_27131);
xor U27438 (N_27438,N_27267,N_27145);
nor U27439 (N_27439,N_27203,N_27193);
nand U27440 (N_27440,N_27222,N_27025);
and U27441 (N_27441,N_27116,N_27031);
nand U27442 (N_27442,N_27299,N_27194);
nor U27443 (N_27443,N_27127,N_27254);
or U27444 (N_27444,N_27282,N_27242);
and U27445 (N_27445,N_27148,N_27089);
or U27446 (N_27446,N_27177,N_27103);
nor U27447 (N_27447,N_27277,N_27033);
nand U27448 (N_27448,N_27284,N_27095);
nand U27449 (N_27449,N_27101,N_27000);
nor U27450 (N_27450,N_27079,N_27122);
nand U27451 (N_27451,N_27018,N_27087);
nand U27452 (N_27452,N_27188,N_27101);
and U27453 (N_27453,N_27171,N_27048);
or U27454 (N_27454,N_27032,N_27207);
and U27455 (N_27455,N_27019,N_27054);
and U27456 (N_27456,N_27151,N_27133);
and U27457 (N_27457,N_27226,N_27248);
nor U27458 (N_27458,N_27100,N_27200);
or U27459 (N_27459,N_27282,N_27287);
or U27460 (N_27460,N_27183,N_27081);
or U27461 (N_27461,N_27239,N_27188);
nand U27462 (N_27462,N_27041,N_27231);
nand U27463 (N_27463,N_27091,N_27144);
nor U27464 (N_27464,N_27252,N_27112);
nor U27465 (N_27465,N_27251,N_27266);
nor U27466 (N_27466,N_27227,N_27230);
nor U27467 (N_27467,N_27032,N_27258);
or U27468 (N_27468,N_27057,N_27081);
or U27469 (N_27469,N_27149,N_27041);
and U27470 (N_27470,N_27095,N_27078);
xnor U27471 (N_27471,N_27220,N_27069);
and U27472 (N_27472,N_27106,N_27160);
and U27473 (N_27473,N_27005,N_27160);
nor U27474 (N_27474,N_27015,N_27163);
nor U27475 (N_27475,N_27100,N_27043);
or U27476 (N_27476,N_27108,N_27097);
and U27477 (N_27477,N_27215,N_27223);
xor U27478 (N_27478,N_27209,N_27290);
or U27479 (N_27479,N_27173,N_27028);
nand U27480 (N_27480,N_27263,N_27161);
nand U27481 (N_27481,N_27036,N_27067);
xor U27482 (N_27482,N_27262,N_27194);
xnor U27483 (N_27483,N_27204,N_27034);
xnor U27484 (N_27484,N_27030,N_27026);
nand U27485 (N_27485,N_27146,N_27017);
or U27486 (N_27486,N_27293,N_27268);
nor U27487 (N_27487,N_27176,N_27056);
xnor U27488 (N_27488,N_27118,N_27188);
nand U27489 (N_27489,N_27041,N_27285);
nor U27490 (N_27490,N_27126,N_27163);
nor U27491 (N_27491,N_27156,N_27110);
xor U27492 (N_27492,N_27028,N_27073);
nor U27493 (N_27493,N_27029,N_27245);
nand U27494 (N_27494,N_27258,N_27084);
and U27495 (N_27495,N_27178,N_27140);
xnor U27496 (N_27496,N_27264,N_27252);
xor U27497 (N_27497,N_27008,N_27288);
and U27498 (N_27498,N_27299,N_27045);
or U27499 (N_27499,N_27162,N_27172);
xnor U27500 (N_27500,N_27111,N_27195);
nor U27501 (N_27501,N_27010,N_27164);
nor U27502 (N_27502,N_27009,N_27170);
nand U27503 (N_27503,N_27271,N_27160);
nor U27504 (N_27504,N_27151,N_27224);
or U27505 (N_27505,N_27024,N_27251);
xnor U27506 (N_27506,N_27285,N_27046);
nand U27507 (N_27507,N_27240,N_27277);
and U27508 (N_27508,N_27244,N_27246);
or U27509 (N_27509,N_27214,N_27049);
or U27510 (N_27510,N_27191,N_27144);
xnor U27511 (N_27511,N_27186,N_27115);
or U27512 (N_27512,N_27035,N_27032);
or U27513 (N_27513,N_27169,N_27297);
and U27514 (N_27514,N_27086,N_27299);
xnor U27515 (N_27515,N_27192,N_27014);
or U27516 (N_27516,N_27095,N_27163);
and U27517 (N_27517,N_27285,N_27267);
xnor U27518 (N_27518,N_27207,N_27227);
and U27519 (N_27519,N_27080,N_27047);
or U27520 (N_27520,N_27208,N_27159);
and U27521 (N_27521,N_27001,N_27054);
and U27522 (N_27522,N_27207,N_27298);
or U27523 (N_27523,N_27256,N_27179);
or U27524 (N_27524,N_27241,N_27283);
xor U27525 (N_27525,N_27003,N_27058);
and U27526 (N_27526,N_27030,N_27213);
xnor U27527 (N_27527,N_27129,N_27248);
nor U27528 (N_27528,N_27209,N_27198);
xor U27529 (N_27529,N_27223,N_27217);
or U27530 (N_27530,N_27096,N_27035);
or U27531 (N_27531,N_27116,N_27125);
or U27532 (N_27532,N_27264,N_27055);
xnor U27533 (N_27533,N_27153,N_27021);
or U27534 (N_27534,N_27119,N_27255);
nor U27535 (N_27535,N_27294,N_27273);
nand U27536 (N_27536,N_27200,N_27154);
nor U27537 (N_27537,N_27059,N_27290);
nand U27538 (N_27538,N_27040,N_27073);
nor U27539 (N_27539,N_27160,N_27236);
nand U27540 (N_27540,N_27189,N_27247);
nand U27541 (N_27541,N_27031,N_27135);
or U27542 (N_27542,N_27101,N_27017);
nor U27543 (N_27543,N_27017,N_27144);
nand U27544 (N_27544,N_27212,N_27255);
xor U27545 (N_27545,N_27235,N_27165);
nor U27546 (N_27546,N_27237,N_27017);
or U27547 (N_27547,N_27104,N_27254);
xor U27548 (N_27548,N_27122,N_27096);
or U27549 (N_27549,N_27254,N_27232);
or U27550 (N_27550,N_27292,N_27031);
nand U27551 (N_27551,N_27090,N_27038);
xnor U27552 (N_27552,N_27212,N_27227);
or U27553 (N_27553,N_27086,N_27239);
nor U27554 (N_27554,N_27165,N_27297);
nand U27555 (N_27555,N_27176,N_27062);
nand U27556 (N_27556,N_27120,N_27282);
xnor U27557 (N_27557,N_27269,N_27148);
nor U27558 (N_27558,N_27015,N_27056);
xor U27559 (N_27559,N_27002,N_27008);
nor U27560 (N_27560,N_27035,N_27083);
nand U27561 (N_27561,N_27210,N_27112);
nand U27562 (N_27562,N_27201,N_27222);
or U27563 (N_27563,N_27100,N_27045);
or U27564 (N_27564,N_27268,N_27285);
nand U27565 (N_27565,N_27129,N_27062);
xnor U27566 (N_27566,N_27009,N_27113);
and U27567 (N_27567,N_27119,N_27128);
nor U27568 (N_27568,N_27226,N_27096);
or U27569 (N_27569,N_27002,N_27009);
xor U27570 (N_27570,N_27190,N_27125);
nor U27571 (N_27571,N_27265,N_27218);
or U27572 (N_27572,N_27013,N_27194);
nand U27573 (N_27573,N_27091,N_27042);
and U27574 (N_27574,N_27254,N_27272);
nor U27575 (N_27575,N_27168,N_27035);
nand U27576 (N_27576,N_27112,N_27266);
nand U27577 (N_27577,N_27077,N_27248);
nand U27578 (N_27578,N_27071,N_27170);
nand U27579 (N_27579,N_27144,N_27260);
and U27580 (N_27580,N_27113,N_27280);
nor U27581 (N_27581,N_27034,N_27011);
nand U27582 (N_27582,N_27098,N_27200);
and U27583 (N_27583,N_27018,N_27013);
nor U27584 (N_27584,N_27126,N_27049);
or U27585 (N_27585,N_27186,N_27146);
nand U27586 (N_27586,N_27261,N_27094);
nand U27587 (N_27587,N_27115,N_27083);
or U27588 (N_27588,N_27176,N_27082);
and U27589 (N_27589,N_27194,N_27060);
nor U27590 (N_27590,N_27178,N_27281);
and U27591 (N_27591,N_27009,N_27036);
xnor U27592 (N_27592,N_27183,N_27194);
or U27593 (N_27593,N_27033,N_27224);
nor U27594 (N_27594,N_27076,N_27036);
or U27595 (N_27595,N_27105,N_27235);
or U27596 (N_27596,N_27247,N_27170);
nor U27597 (N_27597,N_27239,N_27253);
nor U27598 (N_27598,N_27265,N_27192);
nor U27599 (N_27599,N_27058,N_27203);
and U27600 (N_27600,N_27525,N_27397);
nor U27601 (N_27601,N_27438,N_27565);
xnor U27602 (N_27602,N_27328,N_27484);
nand U27603 (N_27603,N_27553,N_27408);
nor U27604 (N_27604,N_27335,N_27535);
or U27605 (N_27605,N_27352,N_27540);
xnor U27606 (N_27606,N_27378,N_27522);
or U27607 (N_27607,N_27470,N_27389);
xor U27608 (N_27608,N_27490,N_27430);
nand U27609 (N_27609,N_27375,N_27423);
xnor U27610 (N_27610,N_27353,N_27569);
xor U27611 (N_27611,N_27455,N_27336);
nor U27612 (N_27612,N_27555,N_27413);
or U27613 (N_27613,N_27447,N_27339);
xor U27614 (N_27614,N_27479,N_27394);
nand U27615 (N_27615,N_27581,N_27477);
xnor U27616 (N_27616,N_27518,N_27305);
and U27617 (N_27617,N_27530,N_27402);
nor U27618 (N_27618,N_27376,N_27452);
or U27619 (N_27619,N_27340,N_27363);
nor U27620 (N_27620,N_27310,N_27506);
xnor U27621 (N_27621,N_27431,N_27531);
or U27622 (N_27622,N_27457,N_27383);
nor U27623 (N_27623,N_27445,N_27496);
nand U27624 (N_27624,N_27332,N_27492);
or U27625 (N_27625,N_27349,N_27382);
nand U27626 (N_27626,N_27485,N_27466);
and U27627 (N_27627,N_27521,N_27460);
nand U27628 (N_27628,N_27356,N_27308);
xor U27629 (N_27629,N_27331,N_27415);
or U27630 (N_27630,N_27343,N_27410);
nor U27631 (N_27631,N_27468,N_27591);
xor U27632 (N_27632,N_27421,N_27385);
nor U27633 (N_27633,N_27598,N_27585);
or U27634 (N_27634,N_27437,N_27502);
and U27635 (N_27635,N_27347,N_27323);
and U27636 (N_27636,N_27509,N_27354);
nand U27637 (N_27637,N_27412,N_27481);
nor U27638 (N_27638,N_27568,N_27450);
xor U27639 (N_27639,N_27558,N_27360);
or U27640 (N_27640,N_27514,N_27393);
and U27641 (N_27641,N_27465,N_27440);
and U27642 (N_27642,N_27498,N_27384);
xnor U27643 (N_27643,N_27529,N_27510);
and U27644 (N_27644,N_27491,N_27566);
nor U27645 (N_27645,N_27417,N_27401);
nand U27646 (N_27646,N_27409,N_27419);
nand U27647 (N_27647,N_27507,N_27444);
nor U27648 (N_27648,N_27513,N_27346);
nor U27649 (N_27649,N_27420,N_27330);
nand U27650 (N_27650,N_27309,N_27588);
and U27651 (N_27651,N_27392,N_27592);
nand U27652 (N_27652,N_27511,N_27319);
and U27653 (N_27653,N_27501,N_27303);
and U27654 (N_27654,N_27435,N_27536);
nand U27655 (N_27655,N_27391,N_27441);
and U27656 (N_27656,N_27489,N_27398);
and U27657 (N_27657,N_27395,N_27472);
xnor U27658 (N_27658,N_27379,N_27453);
and U27659 (N_27659,N_27311,N_27541);
nor U27660 (N_27660,N_27414,N_27570);
nand U27661 (N_27661,N_27390,N_27517);
xor U27662 (N_27662,N_27315,N_27550);
nor U27663 (N_27663,N_27436,N_27579);
or U27664 (N_27664,N_27596,N_27373);
nor U27665 (N_27665,N_27345,N_27451);
nor U27666 (N_27666,N_27473,N_27334);
xor U27667 (N_27667,N_27351,N_27478);
and U27668 (N_27668,N_27377,N_27563);
or U27669 (N_27669,N_27371,N_27512);
nor U27670 (N_27670,N_27306,N_27543);
and U27671 (N_27671,N_27562,N_27590);
nand U27672 (N_27672,N_27316,N_27503);
and U27673 (N_27673,N_27442,N_27405);
nand U27674 (N_27674,N_27427,N_27554);
xnor U27675 (N_27675,N_27443,N_27552);
nand U27676 (N_27676,N_27344,N_27586);
nor U27677 (N_27677,N_27559,N_27547);
and U27678 (N_27678,N_27314,N_27333);
xor U27679 (N_27679,N_27464,N_27580);
nor U27680 (N_27680,N_27583,N_27462);
and U27681 (N_27681,N_27388,N_27483);
and U27682 (N_27682,N_27359,N_27534);
nand U27683 (N_27683,N_27320,N_27557);
and U27684 (N_27684,N_27533,N_27301);
or U27685 (N_27685,N_27422,N_27317);
nor U27686 (N_27686,N_27322,N_27572);
xnor U27687 (N_27687,N_27428,N_27575);
nand U27688 (N_27688,N_27399,N_27471);
and U27689 (N_27689,N_27571,N_27500);
or U27690 (N_27690,N_27355,N_27487);
or U27691 (N_27691,N_27404,N_27364);
xnor U27692 (N_27692,N_27499,N_27381);
or U27693 (N_27693,N_27561,N_27337);
and U27694 (N_27694,N_27476,N_27459);
and U27695 (N_27695,N_27454,N_27495);
and U27696 (N_27696,N_27577,N_27368);
and U27697 (N_27697,N_27300,N_27527);
or U27698 (N_27698,N_27474,N_27467);
or U27699 (N_27699,N_27325,N_27432);
and U27700 (N_27700,N_27307,N_27429);
nand U27701 (N_27701,N_27520,N_27519);
nand U27702 (N_27702,N_27505,N_27304);
nand U27703 (N_27703,N_27326,N_27488);
xnor U27704 (N_27704,N_27365,N_27573);
nand U27705 (N_27705,N_27313,N_27539);
and U27706 (N_27706,N_27387,N_27538);
xnor U27707 (N_27707,N_27551,N_27482);
nor U27708 (N_27708,N_27549,N_27584);
or U27709 (N_27709,N_27595,N_27458);
nor U27710 (N_27710,N_27537,N_27342);
and U27711 (N_27711,N_27348,N_27523);
or U27712 (N_27712,N_27528,N_27321);
xor U27713 (N_27713,N_27302,N_27480);
nand U27714 (N_27714,N_27526,N_27411);
or U27715 (N_27715,N_27407,N_27396);
nand U27716 (N_27716,N_27548,N_27456);
or U27717 (N_27717,N_27403,N_27357);
nand U27718 (N_27718,N_27369,N_27434);
nor U27719 (N_27719,N_27448,N_27329);
xor U27720 (N_27720,N_27416,N_27524);
xnor U27721 (N_27721,N_27564,N_27576);
or U27722 (N_27722,N_27424,N_27475);
nand U27723 (N_27723,N_27338,N_27469);
or U27724 (N_27724,N_27556,N_27589);
and U27725 (N_27725,N_27515,N_27560);
nor U27726 (N_27726,N_27532,N_27599);
or U27727 (N_27727,N_27461,N_27374);
or U27728 (N_27728,N_27358,N_27406);
nor U27729 (N_27729,N_27366,N_27362);
nor U27730 (N_27730,N_27544,N_27425);
or U27731 (N_27731,N_27312,N_27324);
or U27732 (N_27732,N_27593,N_27494);
or U27733 (N_27733,N_27361,N_27587);
nor U27734 (N_27734,N_27594,N_27341);
or U27735 (N_27735,N_27380,N_27400);
xnor U27736 (N_27736,N_27318,N_27350);
or U27737 (N_27737,N_27327,N_27486);
xor U27738 (N_27738,N_27546,N_27386);
nor U27739 (N_27739,N_27504,N_27426);
nor U27740 (N_27740,N_27463,N_27516);
and U27741 (N_27741,N_27449,N_27493);
or U27742 (N_27742,N_27439,N_27446);
and U27743 (N_27743,N_27497,N_27418);
or U27744 (N_27744,N_27372,N_27370);
nand U27745 (N_27745,N_27567,N_27545);
nor U27746 (N_27746,N_27578,N_27582);
nor U27747 (N_27747,N_27542,N_27433);
xor U27748 (N_27748,N_27574,N_27367);
and U27749 (N_27749,N_27508,N_27597);
nor U27750 (N_27750,N_27597,N_27444);
or U27751 (N_27751,N_27344,N_27559);
or U27752 (N_27752,N_27338,N_27592);
nor U27753 (N_27753,N_27452,N_27366);
and U27754 (N_27754,N_27344,N_27448);
nand U27755 (N_27755,N_27455,N_27426);
or U27756 (N_27756,N_27331,N_27396);
xnor U27757 (N_27757,N_27449,N_27334);
or U27758 (N_27758,N_27558,N_27585);
and U27759 (N_27759,N_27512,N_27518);
or U27760 (N_27760,N_27495,N_27354);
nand U27761 (N_27761,N_27353,N_27551);
nand U27762 (N_27762,N_27384,N_27572);
nor U27763 (N_27763,N_27306,N_27464);
nand U27764 (N_27764,N_27544,N_27373);
nand U27765 (N_27765,N_27523,N_27555);
nor U27766 (N_27766,N_27531,N_27474);
and U27767 (N_27767,N_27400,N_27455);
and U27768 (N_27768,N_27563,N_27511);
nor U27769 (N_27769,N_27511,N_27536);
nor U27770 (N_27770,N_27339,N_27442);
and U27771 (N_27771,N_27398,N_27518);
nor U27772 (N_27772,N_27595,N_27472);
nor U27773 (N_27773,N_27352,N_27340);
xor U27774 (N_27774,N_27497,N_27470);
nor U27775 (N_27775,N_27365,N_27597);
nand U27776 (N_27776,N_27511,N_27520);
or U27777 (N_27777,N_27515,N_27323);
nand U27778 (N_27778,N_27597,N_27473);
and U27779 (N_27779,N_27305,N_27369);
nand U27780 (N_27780,N_27327,N_27582);
and U27781 (N_27781,N_27450,N_27506);
xor U27782 (N_27782,N_27552,N_27579);
xor U27783 (N_27783,N_27388,N_27566);
or U27784 (N_27784,N_27376,N_27349);
or U27785 (N_27785,N_27417,N_27442);
xnor U27786 (N_27786,N_27411,N_27563);
nor U27787 (N_27787,N_27506,N_27424);
and U27788 (N_27788,N_27308,N_27435);
xnor U27789 (N_27789,N_27526,N_27542);
xor U27790 (N_27790,N_27405,N_27451);
nand U27791 (N_27791,N_27588,N_27389);
xnor U27792 (N_27792,N_27560,N_27364);
nor U27793 (N_27793,N_27321,N_27530);
xor U27794 (N_27794,N_27587,N_27563);
nand U27795 (N_27795,N_27488,N_27346);
nand U27796 (N_27796,N_27419,N_27400);
or U27797 (N_27797,N_27555,N_27565);
and U27798 (N_27798,N_27387,N_27522);
nor U27799 (N_27799,N_27399,N_27315);
or U27800 (N_27800,N_27530,N_27537);
nand U27801 (N_27801,N_27566,N_27372);
xnor U27802 (N_27802,N_27594,N_27475);
nand U27803 (N_27803,N_27440,N_27549);
nand U27804 (N_27804,N_27384,N_27449);
nor U27805 (N_27805,N_27536,N_27312);
xor U27806 (N_27806,N_27404,N_27546);
or U27807 (N_27807,N_27434,N_27449);
or U27808 (N_27808,N_27552,N_27404);
and U27809 (N_27809,N_27570,N_27318);
or U27810 (N_27810,N_27574,N_27572);
or U27811 (N_27811,N_27463,N_27549);
nand U27812 (N_27812,N_27328,N_27494);
nand U27813 (N_27813,N_27318,N_27508);
nor U27814 (N_27814,N_27386,N_27564);
nand U27815 (N_27815,N_27328,N_27385);
xnor U27816 (N_27816,N_27335,N_27553);
nor U27817 (N_27817,N_27509,N_27454);
or U27818 (N_27818,N_27422,N_27420);
nor U27819 (N_27819,N_27304,N_27431);
and U27820 (N_27820,N_27557,N_27469);
xnor U27821 (N_27821,N_27383,N_27576);
and U27822 (N_27822,N_27517,N_27569);
nor U27823 (N_27823,N_27444,N_27341);
or U27824 (N_27824,N_27400,N_27459);
nor U27825 (N_27825,N_27560,N_27530);
xnor U27826 (N_27826,N_27320,N_27531);
nand U27827 (N_27827,N_27533,N_27504);
nor U27828 (N_27828,N_27531,N_27592);
or U27829 (N_27829,N_27392,N_27427);
xor U27830 (N_27830,N_27442,N_27512);
xnor U27831 (N_27831,N_27487,N_27304);
xnor U27832 (N_27832,N_27568,N_27318);
nor U27833 (N_27833,N_27521,N_27405);
nand U27834 (N_27834,N_27424,N_27564);
and U27835 (N_27835,N_27375,N_27480);
nor U27836 (N_27836,N_27433,N_27567);
nor U27837 (N_27837,N_27530,N_27518);
or U27838 (N_27838,N_27353,N_27445);
xor U27839 (N_27839,N_27490,N_27314);
xor U27840 (N_27840,N_27372,N_27578);
or U27841 (N_27841,N_27396,N_27471);
and U27842 (N_27842,N_27598,N_27419);
nor U27843 (N_27843,N_27358,N_27553);
xor U27844 (N_27844,N_27513,N_27409);
xnor U27845 (N_27845,N_27416,N_27477);
nor U27846 (N_27846,N_27533,N_27399);
nand U27847 (N_27847,N_27463,N_27453);
nand U27848 (N_27848,N_27441,N_27459);
nand U27849 (N_27849,N_27535,N_27363);
xor U27850 (N_27850,N_27305,N_27443);
nor U27851 (N_27851,N_27518,N_27477);
or U27852 (N_27852,N_27538,N_27565);
and U27853 (N_27853,N_27308,N_27409);
and U27854 (N_27854,N_27590,N_27465);
and U27855 (N_27855,N_27504,N_27358);
nor U27856 (N_27856,N_27568,N_27345);
nand U27857 (N_27857,N_27352,N_27571);
and U27858 (N_27858,N_27375,N_27419);
xnor U27859 (N_27859,N_27576,N_27586);
or U27860 (N_27860,N_27516,N_27483);
nor U27861 (N_27861,N_27303,N_27466);
and U27862 (N_27862,N_27519,N_27333);
nand U27863 (N_27863,N_27379,N_27538);
nor U27864 (N_27864,N_27341,N_27532);
and U27865 (N_27865,N_27356,N_27431);
xor U27866 (N_27866,N_27350,N_27543);
and U27867 (N_27867,N_27435,N_27389);
nor U27868 (N_27868,N_27557,N_27395);
nor U27869 (N_27869,N_27483,N_27425);
nand U27870 (N_27870,N_27423,N_27574);
or U27871 (N_27871,N_27542,N_27440);
nor U27872 (N_27872,N_27345,N_27305);
nor U27873 (N_27873,N_27441,N_27574);
xnor U27874 (N_27874,N_27493,N_27315);
nor U27875 (N_27875,N_27367,N_27439);
nor U27876 (N_27876,N_27516,N_27519);
xor U27877 (N_27877,N_27431,N_27439);
and U27878 (N_27878,N_27339,N_27509);
and U27879 (N_27879,N_27311,N_27449);
xor U27880 (N_27880,N_27321,N_27444);
nand U27881 (N_27881,N_27491,N_27520);
or U27882 (N_27882,N_27370,N_27366);
nor U27883 (N_27883,N_27447,N_27543);
nor U27884 (N_27884,N_27397,N_27473);
and U27885 (N_27885,N_27342,N_27314);
xor U27886 (N_27886,N_27426,N_27596);
xor U27887 (N_27887,N_27329,N_27570);
and U27888 (N_27888,N_27510,N_27329);
and U27889 (N_27889,N_27329,N_27371);
or U27890 (N_27890,N_27501,N_27443);
nand U27891 (N_27891,N_27591,N_27400);
xnor U27892 (N_27892,N_27567,N_27495);
nand U27893 (N_27893,N_27438,N_27330);
xnor U27894 (N_27894,N_27526,N_27556);
nor U27895 (N_27895,N_27416,N_27340);
nand U27896 (N_27896,N_27510,N_27355);
and U27897 (N_27897,N_27490,N_27561);
or U27898 (N_27898,N_27340,N_27399);
and U27899 (N_27899,N_27368,N_27564);
nand U27900 (N_27900,N_27709,N_27815);
xor U27901 (N_27901,N_27670,N_27856);
and U27902 (N_27902,N_27819,N_27684);
or U27903 (N_27903,N_27801,N_27798);
nor U27904 (N_27904,N_27702,N_27778);
nand U27905 (N_27905,N_27857,N_27604);
nand U27906 (N_27906,N_27853,N_27727);
or U27907 (N_27907,N_27636,N_27607);
nand U27908 (N_27908,N_27791,N_27738);
nand U27909 (N_27909,N_27679,N_27692);
nor U27910 (N_27910,N_27848,N_27644);
xnor U27911 (N_27911,N_27659,N_27745);
and U27912 (N_27912,N_27790,N_27690);
and U27913 (N_27913,N_27601,N_27872);
xor U27914 (N_27914,N_27754,N_27897);
nor U27915 (N_27915,N_27775,N_27810);
or U27916 (N_27916,N_27715,N_27662);
nand U27917 (N_27917,N_27806,N_27732);
and U27918 (N_27918,N_27718,N_27839);
and U27919 (N_27919,N_27637,N_27752);
xnor U27920 (N_27920,N_27698,N_27657);
or U27921 (N_27921,N_27630,N_27640);
or U27922 (N_27922,N_27693,N_27681);
or U27923 (N_27923,N_27820,N_27749);
and U27924 (N_27924,N_27890,N_27844);
nor U27925 (N_27925,N_27629,N_27850);
or U27926 (N_27926,N_27833,N_27643);
nor U27927 (N_27927,N_27697,N_27700);
and U27928 (N_27928,N_27838,N_27765);
or U27929 (N_27929,N_27647,N_27612);
or U27930 (N_27930,N_27606,N_27770);
nor U27931 (N_27931,N_27882,N_27773);
nand U27932 (N_27932,N_27734,N_27739);
or U27933 (N_27933,N_27809,N_27748);
nor U27934 (N_27934,N_27879,N_27691);
xnor U27935 (N_27935,N_27795,N_27895);
nand U27936 (N_27936,N_27769,N_27781);
xor U27937 (N_27937,N_27812,N_27859);
and U27938 (N_27938,N_27652,N_27863);
xnor U27939 (N_27939,N_27631,N_27656);
or U27940 (N_27940,N_27864,N_27811);
and U27941 (N_27941,N_27704,N_27868);
nand U27942 (N_27942,N_27825,N_27733);
xor U27943 (N_27943,N_27837,N_27755);
nor U27944 (N_27944,N_27625,N_27663);
or U27945 (N_27945,N_27685,N_27766);
and U27946 (N_27946,N_27677,N_27741);
xnor U27947 (N_27947,N_27807,N_27880);
or U27948 (N_27948,N_27676,N_27768);
xnor U27949 (N_27949,N_27746,N_27878);
and U27950 (N_27950,N_27826,N_27683);
or U27951 (N_27951,N_27628,N_27874);
nand U27952 (N_27952,N_27642,N_27696);
nor U27953 (N_27953,N_27694,N_27830);
and U27954 (N_27954,N_27860,N_27666);
xnor U27955 (N_27955,N_27701,N_27831);
nor U27956 (N_27956,N_27731,N_27805);
and U27957 (N_27957,N_27892,N_27703);
or U27958 (N_27958,N_27852,N_27821);
nor U27959 (N_27959,N_27780,N_27808);
nor U27960 (N_27960,N_27846,N_27608);
nor U27961 (N_27961,N_27743,N_27651);
xor U27962 (N_27962,N_27641,N_27602);
nand U27963 (N_27963,N_27646,N_27623);
nand U27964 (N_27964,N_27744,N_27610);
nand U27965 (N_27965,N_27619,N_27638);
nand U27966 (N_27966,N_27621,N_27776);
nor U27967 (N_27967,N_27876,N_27842);
nand U27968 (N_27968,N_27869,N_27854);
and U27969 (N_27969,N_27764,N_27689);
xnor U27970 (N_27970,N_27843,N_27664);
nor U27971 (N_27971,N_27871,N_27841);
nor U27972 (N_27972,N_27803,N_27779);
nand U27973 (N_27973,N_27829,N_27726);
xor U27974 (N_27974,N_27672,N_27721);
and U27975 (N_27975,N_27740,N_27817);
xnor U27976 (N_27976,N_27688,N_27858);
and U27977 (N_27977,N_27639,N_27832);
nand U27978 (N_27978,N_27896,N_27712);
or U27979 (N_27979,N_27814,N_27802);
or U27980 (N_27980,N_27634,N_27759);
and U27981 (N_27981,N_27635,N_27706);
nand U27982 (N_27982,N_27788,N_27665);
xor U27983 (N_27983,N_27615,N_27785);
or U27984 (N_27984,N_27645,N_27671);
and U27985 (N_27985,N_27626,N_27816);
or U27986 (N_27986,N_27894,N_27855);
or U27987 (N_27987,N_27763,N_27678);
or U27988 (N_27988,N_27705,N_27654);
and U27989 (N_27989,N_27633,N_27742);
xor U27990 (N_27990,N_27865,N_27762);
or U27991 (N_27991,N_27613,N_27614);
nor U27992 (N_27992,N_27822,N_27714);
and U27993 (N_27993,N_27753,N_27772);
nor U27994 (N_27994,N_27632,N_27867);
nand U27995 (N_27995,N_27888,N_27877);
and U27996 (N_27996,N_27899,N_27669);
and U27997 (N_27997,N_27680,N_27827);
xor U27998 (N_27998,N_27710,N_27747);
and U27999 (N_27999,N_27787,N_27620);
nand U28000 (N_28000,N_27756,N_27618);
nor U28001 (N_28001,N_27616,N_27728);
xor U28002 (N_28002,N_27862,N_27883);
or U28003 (N_28003,N_27797,N_27760);
nor U28004 (N_28004,N_27722,N_27655);
and U28005 (N_28005,N_27717,N_27845);
nand U28006 (N_28006,N_27611,N_27761);
or U28007 (N_28007,N_27873,N_27716);
nor U28008 (N_28008,N_27751,N_27730);
xnor U28009 (N_28009,N_27886,N_27884);
or U28010 (N_28010,N_27675,N_27725);
and U28011 (N_28011,N_27835,N_27667);
xnor U28012 (N_28012,N_27875,N_27605);
nand U28013 (N_28013,N_27783,N_27881);
and U28014 (N_28014,N_27849,N_27794);
xnor U28015 (N_28015,N_27834,N_27673);
nand U28016 (N_28016,N_27840,N_27847);
xor U28017 (N_28017,N_27711,N_27650);
or U28018 (N_28018,N_27813,N_27889);
xnor U28019 (N_28019,N_27796,N_27818);
and U28020 (N_28020,N_27800,N_27600);
or U28021 (N_28021,N_27767,N_27782);
nand U28022 (N_28022,N_27686,N_27699);
and U28023 (N_28023,N_27866,N_27649);
nor U28024 (N_28024,N_27861,N_27624);
nor U28025 (N_28025,N_27828,N_27851);
nor U28026 (N_28026,N_27648,N_27789);
and U28027 (N_28027,N_27719,N_27713);
nor U28028 (N_28028,N_27898,N_27870);
xnor U28029 (N_28029,N_27758,N_27786);
or U28030 (N_28030,N_27799,N_27887);
nor U28031 (N_28031,N_27771,N_27658);
or U28032 (N_28032,N_27723,N_27777);
or U28033 (N_28033,N_27603,N_27707);
nor U28034 (N_28034,N_27668,N_27774);
xnor U28035 (N_28035,N_27784,N_27724);
nor U28036 (N_28036,N_27792,N_27891);
nor U28037 (N_28037,N_27729,N_27757);
or U28038 (N_28038,N_27823,N_27804);
nand U28039 (N_28039,N_27695,N_27674);
xor U28040 (N_28040,N_27661,N_27627);
nand U28041 (N_28041,N_27720,N_27737);
or U28042 (N_28042,N_27609,N_27893);
xnor U28043 (N_28043,N_27708,N_27617);
xnor U28044 (N_28044,N_27793,N_27622);
nand U28045 (N_28045,N_27736,N_27824);
nand U28046 (N_28046,N_27660,N_27682);
or U28047 (N_28047,N_27750,N_27653);
nand U28048 (N_28048,N_27885,N_27735);
nand U28049 (N_28049,N_27687,N_27836);
nand U28050 (N_28050,N_27769,N_27806);
or U28051 (N_28051,N_27767,N_27897);
and U28052 (N_28052,N_27891,N_27651);
nor U28053 (N_28053,N_27750,N_27765);
and U28054 (N_28054,N_27861,N_27799);
nor U28055 (N_28055,N_27825,N_27671);
or U28056 (N_28056,N_27773,N_27627);
and U28057 (N_28057,N_27699,N_27895);
and U28058 (N_28058,N_27786,N_27655);
or U28059 (N_28059,N_27795,N_27680);
nand U28060 (N_28060,N_27890,N_27762);
xor U28061 (N_28061,N_27755,N_27845);
and U28062 (N_28062,N_27747,N_27839);
or U28063 (N_28063,N_27824,N_27619);
and U28064 (N_28064,N_27738,N_27754);
nand U28065 (N_28065,N_27793,N_27665);
or U28066 (N_28066,N_27715,N_27607);
or U28067 (N_28067,N_27681,N_27770);
and U28068 (N_28068,N_27669,N_27729);
or U28069 (N_28069,N_27832,N_27732);
xor U28070 (N_28070,N_27811,N_27675);
nor U28071 (N_28071,N_27690,N_27604);
nand U28072 (N_28072,N_27803,N_27732);
xnor U28073 (N_28073,N_27674,N_27808);
or U28074 (N_28074,N_27697,N_27763);
or U28075 (N_28075,N_27886,N_27720);
nand U28076 (N_28076,N_27839,N_27709);
or U28077 (N_28077,N_27831,N_27722);
and U28078 (N_28078,N_27618,N_27753);
or U28079 (N_28079,N_27656,N_27883);
and U28080 (N_28080,N_27892,N_27756);
or U28081 (N_28081,N_27600,N_27612);
or U28082 (N_28082,N_27805,N_27817);
nor U28083 (N_28083,N_27612,N_27759);
and U28084 (N_28084,N_27610,N_27773);
nor U28085 (N_28085,N_27725,N_27716);
xor U28086 (N_28086,N_27715,N_27806);
and U28087 (N_28087,N_27874,N_27810);
nand U28088 (N_28088,N_27657,N_27639);
nand U28089 (N_28089,N_27898,N_27696);
xor U28090 (N_28090,N_27776,N_27777);
nand U28091 (N_28091,N_27784,N_27829);
xor U28092 (N_28092,N_27883,N_27865);
nor U28093 (N_28093,N_27874,N_27726);
xnor U28094 (N_28094,N_27706,N_27795);
xor U28095 (N_28095,N_27629,N_27805);
xnor U28096 (N_28096,N_27813,N_27714);
nand U28097 (N_28097,N_27724,N_27818);
or U28098 (N_28098,N_27746,N_27761);
xnor U28099 (N_28099,N_27823,N_27774);
xnor U28100 (N_28100,N_27795,N_27739);
or U28101 (N_28101,N_27675,N_27740);
nor U28102 (N_28102,N_27736,N_27619);
and U28103 (N_28103,N_27896,N_27702);
and U28104 (N_28104,N_27776,N_27833);
nor U28105 (N_28105,N_27672,N_27806);
or U28106 (N_28106,N_27890,N_27796);
or U28107 (N_28107,N_27851,N_27787);
and U28108 (N_28108,N_27744,N_27882);
nor U28109 (N_28109,N_27765,N_27605);
nor U28110 (N_28110,N_27747,N_27817);
nor U28111 (N_28111,N_27727,N_27713);
and U28112 (N_28112,N_27672,N_27665);
nand U28113 (N_28113,N_27735,N_27652);
nor U28114 (N_28114,N_27774,N_27830);
nor U28115 (N_28115,N_27721,N_27851);
xor U28116 (N_28116,N_27898,N_27666);
and U28117 (N_28117,N_27767,N_27776);
nand U28118 (N_28118,N_27785,N_27657);
nand U28119 (N_28119,N_27892,N_27730);
and U28120 (N_28120,N_27779,N_27655);
and U28121 (N_28121,N_27740,N_27668);
and U28122 (N_28122,N_27847,N_27829);
and U28123 (N_28123,N_27662,N_27869);
xnor U28124 (N_28124,N_27712,N_27675);
nor U28125 (N_28125,N_27835,N_27650);
nand U28126 (N_28126,N_27617,N_27738);
or U28127 (N_28127,N_27668,N_27743);
nand U28128 (N_28128,N_27661,N_27822);
xor U28129 (N_28129,N_27666,N_27855);
and U28130 (N_28130,N_27783,N_27676);
or U28131 (N_28131,N_27845,N_27732);
xor U28132 (N_28132,N_27809,N_27895);
and U28133 (N_28133,N_27603,N_27777);
and U28134 (N_28134,N_27888,N_27777);
nor U28135 (N_28135,N_27814,N_27707);
nand U28136 (N_28136,N_27693,N_27601);
nor U28137 (N_28137,N_27693,N_27766);
and U28138 (N_28138,N_27711,N_27831);
or U28139 (N_28139,N_27849,N_27702);
nor U28140 (N_28140,N_27806,N_27616);
and U28141 (N_28141,N_27827,N_27852);
nand U28142 (N_28142,N_27706,N_27602);
nand U28143 (N_28143,N_27779,N_27678);
nor U28144 (N_28144,N_27674,N_27778);
xnor U28145 (N_28145,N_27709,N_27618);
or U28146 (N_28146,N_27743,N_27700);
nor U28147 (N_28147,N_27837,N_27619);
nand U28148 (N_28148,N_27899,N_27808);
nand U28149 (N_28149,N_27673,N_27689);
nor U28150 (N_28150,N_27783,N_27795);
xor U28151 (N_28151,N_27898,N_27752);
nor U28152 (N_28152,N_27834,N_27799);
or U28153 (N_28153,N_27686,N_27784);
nand U28154 (N_28154,N_27748,N_27729);
or U28155 (N_28155,N_27761,N_27871);
and U28156 (N_28156,N_27683,N_27682);
nand U28157 (N_28157,N_27643,N_27736);
xnor U28158 (N_28158,N_27692,N_27889);
nor U28159 (N_28159,N_27663,N_27609);
xor U28160 (N_28160,N_27615,N_27744);
nor U28161 (N_28161,N_27860,N_27872);
or U28162 (N_28162,N_27747,N_27729);
nor U28163 (N_28163,N_27719,N_27763);
or U28164 (N_28164,N_27652,N_27849);
nand U28165 (N_28165,N_27618,N_27759);
xor U28166 (N_28166,N_27700,N_27736);
xnor U28167 (N_28167,N_27714,N_27613);
nand U28168 (N_28168,N_27614,N_27725);
nor U28169 (N_28169,N_27712,N_27679);
nor U28170 (N_28170,N_27670,N_27705);
xnor U28171 (N_28171,N_27859,N_27625);
or U28172 (N_28172,N_27601,N_27619);
nor U28173 (N_28173,N_27632,N_27734);
xnor U28174 (N_28174,N_27666,N_27868);
nand U28175 (N_28175,N_27692,N_27600);
xor U28176 (N_28176,N_27665,N_27654);
nand U28177 (N_28177,N_27805,N_27645);
nand U28178 (N_28178,N_27885,N_27743);
nand U28179 (N_28179,N_27834,N_27624);
nand U28180 (N_28180,N_27677,N_27743);
and U28181 (N_28181,N_27601,N_27689);
nor U28182 (N_28182,N_27681,N_27787);
and U28183 (N_28183,N_27841,N_27614);
nand U28184 (N_28184,N_27754,N_27893);
nor U28185 (N_28185,N_27835,N_27711);
nand U28186 (N_28186,N_27836,N_27752);
nand U28187 (N_28187,N_27801,N_27648);
or U28188 (N_28188,N_27796,N_27672);
and U28189 (N_28189,N_27709,N_27844);
nand U28190 (N_28190,N_27768,N_27846);
or U28191 (N_28191,N_27812,N_27629);
and U28192 (N_28192,N_27600,N_27648);
nand U28193 (N_28193,N_27774,N_27853);
or U28194 (N_28194,N_27892,N_27646);
nor U28195 (N_28195,N_27728,N_27898);
or U28196 (N_28196,N_27658,N_27847);
xnor U28197 (N_28197,N_27679,N_27619);
and U28198 (N_28198,N_27840,N_27800);
or U28199 (N_28199,N_27726,N_27773);
xnor U28200 (N_28200,N_28115,N_28124);
and U28201 (N_28201,N_28090,N_28184);
nand U28202 (N_28202,N_28154,N_28104);
and U28203 (N_28203,N_28082,N_27928);
nor U28204 (N_28204,N_27951,N_28084);
and U28205 (N_28205,N_28022,N_27975);
nand U28206 (N_28206,N_28064,N_28152);
nand U28207 (N_28207,N_28185,N_27913);
xor U28208 (N_28208,N_28103,N_28164);
or U28209 (N_28209,N_28187,N_27908);
and U28210 (N_28210,N_28063,N_28175);
and U28211 (N_28211,N_28140,N_28179);
nor U28212 (N_28212,N_28173,N_27930);
and U28213 (N_28213,N_28050,N_28067);
nand U28214 (N_28214,N_28027,N_28037);
nor U28215 (N_28215,N_27915,N_27956);
nor U28216 (N_28216,N_28125,N_28126);
nand U28217 (N_28217,N_28088,N_27921);
nor U28218 (N_28218,N_27950,N_27994);
nand U28219 (N_28219,N_27940,N_27963);
and U28220 (N_28220,N_27924,N_28052);
and U28221 (N_28221,N_28180,N_28135);
xor U28222 (N_28222,N_27984,N_27902);
nor U28223 (N_28223,N_28111,N_27979);
and U28224 (N_28224,N_27912,N_27926);
or U28225 (N_28225,N_28036,N_28095);
nor U28226 (N_28226,N_27969,N_28150);
nand U28227 (N_28227,N_28094,N_27953);
and U28228 (N_28228,N_28193,N_28003);
nand U28229 (N_28229,N_28109,N_28192);
and U28230 (N_28230,N_28174,N_27907);
xnor U28231 (N_28231,N_28081,N_28038);
or U28232 (N_28232,N_27996,N_28083);
nor U28233 (N_28233,N_27925,N_28007);
xnor U28234 (N_28234,N_28043,N_28048);
xnor U28235 (N_28235,N_28098,N_27932);
or U28236 (N_28236,N_28080,N_28089);
nor U28237 (N_28237,N_27977,N_27986);
nand U28238 (N_28238,N_27966,N_27946);
nor U28239 (N_28239,N_28128,N_28097);
or U28240 (N_28240,N_28156,N_28108);
and U28241 (N_28241,N_28051,N_28024);
nand U28242 (N_28242,N_27993,N_28077);
xnor U28243 (N_28243,N_27938,N_27937);
or U28244 (N_28244,N_27998,N_27962);
xnor U28245 (N_28245,N_27955,N_28114);
or U28246 (N_28246,N_27964,N_27904);
nor U28247 (N_28247,N_28112,N_28001);
xor U28248 (N_28248,N_28087,N_27933);
or U28249 (N_28249,N_28075,N_28079);
nand U28250 (N_28250,N_28054,N_28198);
or U28251 (N_28251,N_28162,N_28199);
nor U28252 (N_28252,N_28044,N_27910);
or U28253 (N_28253,N_28113,N_28107);
xor U28254 (N_28254,N_28056,N_28130);
nand U28255 (N_28255,N_28146,N_28129);
and U28256 (N_28256,N_27978,N_27991);
or U28257 (N_28257,N_28099,N_28190);
nor U28258 (N_28258,N_28117,N_28053);
nand U28259 (N_28259,N_27989,N_27918);
xor U28260 (N_28260,N_28055,N_28002);
nor U28261 (N_28261,N_28138,N_28158);
xor U28262 (N_28262,N_27922,N_27945);
xnor U28263 (N_28263,N_28172,N_28159);
nand U28264 (N_28264,N_28183,N_28049);
nand U28265 (N_28265,N_28131,N_28033);
xnor U28266 (N_28266,N_28071,N_28145);
xor U28267 (N_28267,N_28015,N_28119);
or U28268 (N_28268,N_27982,N_27959);
and U28269 (N_28269,N_28042,N_27916);
or U28270 (N_28270,N_28076,N_27941);
and U28271 (N_28271,N_28149,N_27968);
nor U28272 (N_28272,N_27943,N_28170);
nand U28273 (N_28273,N_28147,N_28134);
xor U28274 (N_28274,N_28045,N_28065);
and U28275 (N_28275,N_28100,N_27917);
and U28276 (N_28276,N_27948,N_28058);
xnor U28277 (N_28277,N_28072,N_27958);
nor U28278 (N_28278,N_28195,N_27944);
and U28279 (N_28279,N_28106,N_28165);
xor U28280 (N_28280,N_28060,N_28014);
or U28281 (N_28281,N_28029,N_28069);
nand U28282 (N_28282,N_28040,N_28030);
xnor U28283 (N_28283,N_27923,N_28035);
xnor U28284 (N_28284,N_27981,N_28144);
xnor U28285 (N_28285,N_28120,N_27949);
nor U28286 (N_28286,N_28078,N_28092);
xnor U28287 (N_28287,N_27987,N_28163);
nand U28288 (N_28288,N_28132,N_28110);
and U28289 (N_28289,N_28148,N_27900);
xnor U28290 (N_28290,N_28018,N_28013);
and U28291 (N_28291,N_28121,N_28116);
xnor U28292 (N_28292,N_28039,N_27967);
xor U28293 (N_28293,N_28068,N_28177);
nand U28294 (N_28294,N_28197,N_28186);
and U28295 (N_28295,N_28141,N_28182);
and U28296 (N_28296,N_28016,N_28086);
and U28297 (N_28297,N_28176,N_27970);
nand U28298 (N_28298,N_27920,N_28139);
and U28299 (N_28299,N_27965,N_28155);
and U28300 (N_28300,N_27960,N_27961);
nor U28301 (N_28301,N_28085,N_27909);
nor U28302 (N_28302,N_27997,N_28194);
or U28303 (N_28303,N_27985,N_28005);
nor U28304 (N_28304,N_27980,N_27983);
nor U28305 (N_28305,N_28021,N_28032);
nor U28306 (N_28306,N_28167,N_28178);
and U28307 (N_28307,N_27935,N_27972);
xnor U28308 (N_28308,N_28166,N_28153);
xnor U28309 (N_28309,N_28020,N_27939);
nand U28310 (N_28310,N_27999,N_28023);
xnor U28311 (N_28311,N_27988,N_28123);
xnor U28312 (N_28312,N_28091,N_28171);
or U28313 (N_28313,N_28031,N_28061);
nor U28314 (N_28314,N_28143,N_28006);
or U28315 (N_28315,N_28102,N_27934);
xnor U28316 (N_28316,N_27942,N_27901);
or U28317 (N_28317,N_28073,N_28074);
nand U28318 (N_28318,N_27957,N_28000);
or U28319 (N_28319,N_28168,N_28028);
xor U28320 (N_28320,N_28019,N_27992);
nor U28321 (N_28321,N_28012,N_27947);
nor U28322 (N_28322,N_28010,N_28136);
xor U28323 (N_28323,N_27974,N_28047);
xnor U28324 (N_28324,N_27954,N_28157);
and U28325 (N_28325,N_27936,N_28137);
xor U28326 (N_28326,N_28133,N_28189);
and U28327 (N_28327,N_28004,N_27927);
nand U28328 (N_28328,N_27914,N_27931);
nor U28329 (N_28329,N_27919,N_28057);
and U28330 (N_28330,N_28151,N_28062);
or U28331 (N_28331,N_27906,N_28011);
nor U28332 (N_28332,N_28161,N_28096);
nor U28333 (N_28333,N_28025,N_27995);
and U28334 (N_28334,N_28008,N_27911);
xnor U28335 (N_28335,N_27990,N_28196);
or U28336 (N_28336,N_27976,N_28127);
or U28337 (N_28337,N_28026,N_28093);
nor U28338 (N_28338,N_28191,N_28122);
and U28339 (N_28339,N_27971,N_28070);
xnor U28340 (N_28340,N_28160,N_28059);
and U28341 (N_28341,N_28034,N_28142);
and U28342 (N_28342,N_28017,N_27973);
and U28343 (N_28343,N_28188,N_28101);
nor U28344 (N_28344,N_27905,N_28118);
xnor U28345 (N_28345,N_28041,N_27903);
nor U28346 (N_28346,N_28105,N_28181);
xnor U28347 (N_28347,N_27929,N_28009);
and U28348 (N_28348,N_28066,N_28169);
xor U28349 (N_28349,N_27952,N_28046);
or U28350 (N_28350,N_28025,N_28191);
nand U28351 (N_28351,N_28087,N_28057);
and U28352 (N_28352,N_27962,N_28056);
nand U28353 (N_28353,N_28050,N_28143);
xnor U28354 (N_28354,N_27956,N_28186);
nor U28355 (N_28355,N_27928,N_27993);
xor U28356 (N_28356,N_28178,N_27976);
and U28357 (N_28357,N_28167,N_28083);
nand U28358 (N_28358,N_27961,N_28050);
nor U28359 (N_28359,N_28100,N_28119);
and U28360 (N_28360,N_27976,N_28193);
xor U28361 (N_28361,N_28040,N_28189);
and U28362 (N_28362,N_28195,N_28012);
nand U28363 (N_28363,N_28126,N_28159);
xnor U28364 (N_28364,N_27925,N_28072);
nand U28365 (N_28365,N_28069,N_28152);
nand U28366 (N_28366,N_28180,N_28086);
nand U28367 (N_28367,N_28098,N_28198);
xor U28368 (N_28368,N_28133,N_28062);
nor U28369 (N_28369,N_28013,N_28150);
or U28370 (N_28370,N_28130,N_28162);
nor U28371 (N_28371,N_28185,N_28126);
xor U28372 (N_28372,N_27917,N_28024);
nor U28373 (N_28373,N_27971,N_28109);
nor U28374 (N_28374,N_28110,N_27927);
nand U28375 (N_28375,N_28150,N_28176);
or U28376 (N_28376,N_28122,N_27996);
or U28377 (N_28377,N_27953,N_28072);
nand U28378 (N_28378,N_28034,N_27943);
and U28379 (N_28379,N_27913,N_28159);
nor U28380 (N_28380,N_28033,N_27928);
nand U28381 (N_28381,N_28140,N_28168);
nand U28382 (N_28382,N_28118,N_28058);
xnor U28383 (N_28383,N_27958,N_28176);
or U28384 (N_28384,N_28075,N_28197);
nand U28385 (N_28385,N_27927,N_27937);
nand U28386 (N_28386,N_27930,N_28115);
xor U28387 (N_28387,N_27993,N_28027);
xnor U28388 (N_28388,N_28086,N_28047);
and U28389 (N_28389,N_28039,N_27971);
xor U28390 (N_28390,N_28182,N_28120);
and U28391 (N_28391,N_28121,N_28006);
xnor U28392 (N_28392,N_27987,N_28106);
nor U28393 (N_28393,N_27946,N_28171);
and U28394 (N_28394,N_28078,N_28102);
nor U28395 (N_28395,N_28088,N_28071);
nand U28396 (N_28396,N_28144,N_28130);
and U28397 (N_28397,N_27913,N_28046);
or U28398 (N_28398,N_28055,N_28143);
xor U28399 (N_28399,N_28170,N_27981);
nand U28400 (N_28400,N_28024,N_28168);
nor U28401 (N_28401,N_28050,N_28069);
and U28402 (N_28402,N_28168,N_27953);
nor U28403 (N_28403,N_28021,N_28146);
and U28404 (N_28404,N_27952,N_27934);
or U28405 (N_28405,N_28195,N_27965);
nand U28406 (N_28406,N_28198,N_28159);
and U28407 (N_28407,N_27984,N_28147);
nor U28408 (N_28408,N_28046,N_28127);
or U28409 (N_28409,N_28153,N_27956);
or U28410 (N_28410,N_27995,N_28164);
xor U28411 (N_28411,N_27921,N_28067);
or U28412 (N_28412,N_28070,N_28074);
nand U28413 (N_28413,N_27927,N_28133);
or U28414 (N_28414,N_27986,N_28083);
or U28415 (N_28415,N_28046,N_27924);
nor U28416 (N_28416,N_28194,N_28103);
nor U28417 (N_28417,N_27978,N_28105);
or U28418 (N_28418,N_27920,N_28177);
nand U28419 (N_28419,N_27940,N_27990);
and U28420 (N_28420,N_28104,N_27981);
xnor U28421 (N_28421,N_28183,N_28050);
nand U28422 (N_28422,N_28111,N_27991);
and U28423 (N_28423,N_28048,N_27915);
and U28424 (N_28424,N_28173,N_28068);
nand U28425 (N_28425,N_28054,N_28189);
xor U28426 (N_28426,N_28016,N_27987);
xnor U28427 (N_28427,N_28170,N_27975);
and U28428 (N_28428,N_28083,N_28009);
or U28429 (N_28429,N_28058,N_28109);
or U28430 (N_28430,N_28151,N_27975);
or U28431 (N_28431,N_28115,N_28143);
nor U28432 (N_28432,N_27938,N_28111);
and U28433 (N_28433,N_28181,N_28051);
xnor U28434 (N_28434,N_28171,N_28152);
nor U28435 (N_28435,N_28004,N_28007);
nand U28436 (N_28436,N_28058,N_28056);
nor U28437 (N_28437,N_27963,N_28120);
or U28438 (N_28438,N_28085,N_27994);
nand U28439 (N_28439,N_28107,N_27910);
xor U28440 (N_28440,N_28034,N_28195);
nor U28441 (N_28441,N_28141,N_28052);
nor U28442 (N_28442,N_27992,N_28168);
nor U28443 (N_28443,N_27989,N_28090);
xnor U28444 (N_28444,N_28101,N_28087);
nor U28445 (N_28445,N_28198,N_28068);
xor U28446 (N_28446,N_28055,N_27952);
nand U28447 (N_28447,N_28114,N_28062);
or U28448 (N_28448,N_28062,N_28172);
xnor U28449 (N_28449,N_28153,N_28052);
nor U28450 (N_28450,N_28179,N_28103);
nor U28451 (N_28451,N_27904,N_28049);
xor U28452 (N_28452,N_28001,N_28044);
and U28453 (N_28453,N_28073,N_28130);
xnor U28454 (N_28454,N_28042,N_28144);
xnor U28455 (N_28455,N_27980,N_28011);
nor U28456 (N_28456,N_28176,N_28148);
nand U28457 (N_28457,N_27978,N_28005);
xnor U28458 (N_28458,N_27921,N_28161);
nor U28459 (N_28459,N_27916,N_28074);
nand U28460 (N_28460,N_28167,N_27999);
and U28461 (N_28461,N_28072,N_28108);
nor U28462 (N_28462,N_27940,N_28153);
nand U28463 (N_28463,N_28176,N_28130);
nor U28464 (N_28464,N_28136,N_28120);
nor U28465 (N_28465,N_28128,N_28147);
nor U28466 (N_28466,N_28156,N_28197);
nand U28467 (N_28467,N_27954,N_28009);
and U28468 (N_28468,N_28154,N_28086);
or U28469 (N_28469,N_28001,N_27973);
and U28470 (N_28470,N_28197,N_28138);
and U28471 (N_28471,N_28035,N_28165);
nor U28472 (N_28472,N_27935,N_27954);
nand U28473 (N_28473,N_28096,N_28071);
nor U28474 (N_28474,N_28149,N_27994);
xor U28475 (N_28475,N_28007,N_27961);
and U28476 (N_28476,N_28030,N_28044);
and U28477 (N_28477,N_28149,N_27915);
or U28478 (N_28478,N_27908,N_28017);
nand U28479 (N_28479,N_27990,N_27977);
and U28480 (N_28480,N_28185,N_28064);
xnor U28481 (N_28481,N_27913,N_28101);
and U28482 (N_28482,N_28085,N_27992);
nand U28483 (N_28483,N_28007,N_27941);
nor U28484 (N_28484,N_27949,N_28134);
and U28485 (N_28485,N_28194,N_28072);
nand U28486 (N_28486,N_28157,N_28060);
nand U28487 (N_28487,N_27939,N_28133);
nor U28488 (N_28488,N_28151,N_28032);
xnor U28489 (N_28489,N_28135,N_28187);
and U28490 (N_28490,N_28076,N_27968);
xnor U28491 (N_28491,N_27999,N_28064);
or U28492 (N_28492,N_27922,N_27915);
nor U28493 (N_28493,N_28166,N_28197);
nand U28494 (N_28494,N_28008,N_28087);
nand U28495 (N_28495,N_28029,N_28038);
nand U28496 (N_28496,N_27973,N_27904);
and U28497 (N_28497,N_27943,N_28093);
xor U28498 (N_28498,N_27994,N_27905);
or U28499 (N_28499,N_28012,N_27929);
and U28500 (N_28500,N_28450,N_28396);
or U28501 (N_28501,N_28244,N_28227);
xor U28502 (N_28502,N_28355,N_28214);
or U28503 (N_28503,N_28216,N_28342);
and U28504 (N_28504,N_28384,N_28424);
or U28505 (N_28505,N_28315,N_28204);
and U28506 (N_28506,N_28276,N_28377);
and U28507 (N_28507,N_28333,N_28291);
or U28508 (N_28508,N_28222,N_28220);
or U28509 (N_28509,N_28314,N_28295);
xor U28510 (N_28510,N_28260,N_28438);
xor U28511 (N_28511,N_28458,N_28452);
nand U28512 (N_28512,N_28322,N_28442);
nand U28513 (N_28513,N_28329,N_28358);
nand U28514 (N_28514,N_28336,N_28407);
xor U28515 (N_28515,N_28344,N_28369);
nand U28516 (N_28516,N_28376,N_28350);
nand U28517 (N_28517,N_28427,N_28460);
xor U28518 (N_28518,N_28219,N_28443);
xnor U28519 (N_28519,N_28262,N_28261);
nor U28520 (N_28520,N_28309,N_28236);
and U28521 (N_28521,N_28226,N_28257);
and U28522 (N_28522,N_28425,N_28400);
and U28523 (N_28523,N_28431,N_28280);
xor U28524 (N_28524,N_28312,N_28383);
nor U28525 (N_28525,N_28239,N_28439);
or U28526 (N_28526,N_28398,N_28284);
or U28527 (N_28527,N_28434,N_28489);
or U28528 (N_28528,N_28492,N_28463);
nand U28529 (N_28529,N_28328,N_28411);
or U28530 (N_28530,N_28391,N_28302);
nor U28531 (N_28531,N_28402,N_28343);
nor U28532 (N_28532,N_28325,N_28242);
nand U28533 (N_28533,N_28478,N_28475);
xor U28534 (N_28534,N_28285,N_28359);
nand U28535 (N_28535,N_28386,N_28483);
nand U28536 (N_28536,N_28298,N_28406);
and U28537 (N_28537,N_28320,N_28403);
nand U28538 (N_28538,N_28437,N_28297);
nor U28539 (N_28539,N_28332,N_28253);
nand U28540 (N_28540,N_28313,N_28490);
nand U28541 (N_28541,N_28341,N_28390);
xnor U28542 (N_28542,N_28331,N_28357);
and U28543 (N_28543,N_28299,N_28356);
xor U28544 (N_28544,N_28468,N_28401);
and U28545 (N_28545,N_28232,N_28334);
or U28546 (N_28546,N_28388,N_28347);
xor U28547 (N_28547,N_28353,N_28279);
and U28548 (N_28548,N_28224,N_28337);
xor U28549 (N_28549,N_28381,N_28399);
nor U28550 (N_28550,N_28282,N_28385);
or U28551 (N_28551,N_28428,N_28471);
xnor U28552 (N_28552,N_28250,N_28472);
or U28553 (N_28553,N_28362,N_28352);
nand U28554 (N_28554,N_28270,N_28354);
nand U28555 (N_28555,N_28497,N_28267);
nand U28556 (N_28556,N_28290,N_28271);
xor U28557 (N_28557,N_28293,N_28237);
or U28558 (N_28558,N_28202,N_28494);
nor U28559 (N_28559,N_28387,N_28209);
or U28560 (N_28560,N_28351,N_28374);
xor U28561 (N_28561,N_28349,N_28441);
xnor U28562 (N_28562,N_28397,N_28476);
xor U28563 (N_28563,N_28498,N_28340);
or U28564 (N_28564,N_28304,N_28382);
xor U28565 (N_28565,N_28311,N_28266);
or U28566 (N_28566,N_28462,N_28234);
nand U28567 (N_28567,N_28496,N_28417);
and U28568 (N_28568,N_28429,N_28335);
or U28569 (N_28569,N_28485,N_28433);
xor U28570 (N_28570,N_28466,N_28221);
xnor U28571 (N_28571,N_28208,N_28361);
and U28572 (N_28572,N_28430,N_28327);
nor U28573 (N_28573,N_28455,N_28269);
nand U28574 (N_28574,N_28435,N_28405);
and U28575 (N_28575,N_28287,N_28368);
or U28576 (N_28576,N_28464,N_28346);
nand U28577 (N_28577,N_28486,N_28206);
nand U28578 (N_28578,N_28372,N_28223);
nand U28579 (N_28579,N_28263,N_28414);
and U28580 (N_28580,N_28415,N_28409);
nor U28581 (N_28581,N_28495,N_28255);
and U28582 (N_28582,N_28445,N_28394);
and U28583 (N_28583,N_28413,N_28316);
and U28584 (N_28584,N_28319,N_28461);
xnor U28585 (N_28585,N_28278,N_28395);
xnor U28586 (N_28586,N_28225,N_28488);
and U28587 (N_28587,N_28310,N_28467);
xor U28588 (N_28588,N_28248,N_28373);
and U28589 (N_28589,N_28212,N_28251);
or U28590 (N_28590,N_28470,N_28229);
nor U28591 (N_28591,N_28419,N_28481);
xnor U28592 (N_28592,N_28249,N_28321);
and U28593 (N_28593,N_28203,N_28393);
or U28594 (N_28594,N_28281,N_28423);
xor U28595 (N_28595,N_28477,N_28348);
and U28596 (N_28596,N_28252,N_28367);
nand U28597 (N_28597,N_28453,N_28245);
and U28598 (N_28598,N_28338,N_28451);
or U28599 (N_28599,N_28231,N_28364);
xnor U28600 (N_28600,N_28449,N_28412);
or U28601 (N_28601,N_28200,N_28375);
nor U28602 (N_28602,N_28247,N_28294);
nand U28603 (N_28603,N_28233,N_28241);
xnor U28604 (N_28604,N_28421,N_28446);
xor U28605 (N_28605,N_28317,N_28389);
nor U28606 (N_28606,N_28459,N_28210);
or U28607 (N_28607,N_28201,N_28366);
xor U28608 (N_28608,N_28360,N_28286);
and U28609 (N_28609,N_28456,N_28418);
nand U28610 (N_28610,N_28379,N_28211);
and U28611 (N_28611,N_28215,N_28499);
or U28612 (N_28612,N_28303,N_28440);
nand U28613 (N_28613,N_28420,N_28432);
nor U28614 (N_28614,N_28392,N_28479);
nand U28615 (N_28615,N_28482,N_28305);
and U28616 (N_28616,N_28408,N_28330);
or U28617 (N_28617,N_28448,N_28491);
or U28618 (N_28618,N_28457,N_28288);
and U28619 (N_28619,N_28370,N_28217);
nor U28620 (N_28620,N_28275,N_28306);
xor U28621 (N_28621,N_28259,N_28426);
or U28622 (N_28622,N_28345,N_28363);
nand U28623 (N_28623,N_28487,N_28205);
nand U28624 (N_28624,N_28296,N_28289);
xnor U28625 (N_28625,N_28274,N_28235);
or U28626 (N_28626,N_28272,N_28465);
and U28627 (N_28627,N_28326,N_28243);
xnor U28628 (N_28628,N_28283,N_28277);
or U28629 (N_28629,N_28256,N_28473);
nor U28630 (N_28630,N_28240,N_28323);
and U28631 (N_28631,N_28246,N_28301);
and U28632 (N_28632,N_28469,N_28444);
nor U28633 (N_28633,N_28273,N_28218);
or U28634 (N_28634,N_28493,N_28238);
nand U28635 (N_28635,N_28339,N_28447);
nor U28636 (N_28636,N_28454,N_28416);
nand U28637 (N_28637,N_28371,N_28207);
and U28638 (N_28638,N_28480,N_28410);
nor U28639 (N_28639,N_28318,N_28365);
xnor U28640 (N_28640,N_28228,N_28307);
xnor U28641 (N_28641,N_28265,N_28300);
or U28642 (N_28642,N_28264,N_28254);
nor U28643 (N_28643,N_28378,N_28292);
and U28644 (N_28644,N_28436,N_28474);
nand U28645 (N_28645,N_28324,N_28258);
xnor U28646 (N_28646,N_28380,N_28484);
xor U28647 (N_28647,N_28308,N_28422);
nor U28648 (N_28648,N_28404,N_28268);
and U28649 (N_28649,N_28213,N_28230);
xnor U28650 (N_28650,N_28268,N_28393);
and U28651 (N_28651,N_28309,N_28456);
nor U28652 (N_28652,N_28384,N_28291);
nor U28653 (N_28653,N_28309,N_28337);
nor U28654 (N_28654,N_28369,N_28460);
nor U28655 (N_28655,N_28384,N_28487);
and U28656 (N_28656,N_28247,N_28234);
nor U28657 (N_28657,N_28320,N_28204);
and U28658 (N_28658,N_28334,N_28403);
nor U28659 (N_28659,N_28378,N_28453);
xor U28660 (N_28660,N_28206,N_28350);
nand U28661 (N_28661,N_28417,N_28430);
and U28662 (N_28662,N_28469,N_28334);
and U28663 (N_28663,N_28312,N_28489);
xnor U28664 (N_28664,N_28346,N_28285);
or U28665 (N_28665,N_28474,N_28287);
or U28666 (N_28666,N_28376,N_28341);
or U28667 (N_28667,N_28314,N_28285);
nand U28668 (N_28668,N_28343,N_28433);
nand U28669 (N_28669,N_28444,N_28277);
or U28670 (N_28670,N_28258,N_28297);
nand U28671 (N_28671,N_28374,N_28387);
and U28672 (N_28672,N_28237,N_28437);
or U28673 (N_28673,N_28354,N_28234);
and U28674 (N_28674,N_28348,N_28455);
xor U28675 (N_28675,N_28334,N_28227);
or U28676 (N_28676,N_28439,N_28351);
nand U28677 (N_28677,N_28450,N_28366);
and U28678 (N_28678,N_28281,N_28385);
nand U28679 (N_28679,N_28234,N_28298);
xor U28680 (N_28680,N_28448,N_28465);
nor U28681 (N_28681,N_28497,N_28276);
nor U28682 (N_28682,N_28282,N_28347);
nand U28683 (N_28683,N_28308,N_28262);
nand U28684 (N_28684,N_28267,N_28463);
nor U28685 (N_28685,N_28316,N_28298);
xor U28686 (N_28686,N_28437,N_28202);
nand U28687 (N_28687,N_28483,N_28332);
and U28688 (N_28688,N_28399,N_28282);
or U28689 (N_28689,N_28325,N_28453);
and U28690 (N_28690,N_28209,N_28358);
and U28691 (N_28691,N_28452,N_28498);
xnor U28692 (N_28692,N_28276,N_28220);
xnor U28693 (N_28693,N_28366,N_28213);
nor U28694 (N_28694,N_28421,N_28402);
nor U28695 (N_28695,N_28209,N_28364);
nor U28696 (N_28696,N_28460,N_28331);
or U28697 (N_28697,N_28477,N_28256);
xnor U28698 (N_28698,N_28467,N_28414);
nand U28699 (N_28699,N_28404,N_28295);
nand U28700 (N_28700,N_28211,N_28465);
xnor U28701 (N_28701,N_28332,N_28289);
and U28702 (N_28702,N_28246,N_28245);
nor U28703 (N_28703,N_28206,N_28405);
and U28704 (N_28704,N_28201,N_28417);
nor U28705 (N_28705,N_28303,N_28480);
nor U28706 (N_28706,N_28341,N_28377);
xor U28707 (N_28707,N_28353,N_28484);
nor U28708 (N_28708,N_28327,N_28356);
xnor U28709 (N_28709,N_28307,N_28391);
nor U28710 (N_28710,N_28328,N_28489);
xnor U28711 (N_28711,N_28313,N_28212);
nor U28712 (N_28712,N_28242,N_28419);
xor U28713 (N_28713,N_28343,N_28398);
nand U28714 (N_28714,N_28211,N_28200);
nand U28715 (N_28715,N_28420,N_28451);
xor U28716 (N_28716,N_28299,N_28261);
nor U28717 (N_28717,N_28381,N_28241);
and U28718 (N_28718,N_28231,N_28370);
nand U28719 (N_28719,N_28399,N_28341);
nor U28720 (N_28720,N_28301,N_28488);
xor U28721 (N_28721,N_28405,N_28342);
xor U28722 (N_28722,N_28311,N_28290);
xnor U28723 (N_28723,N_28361,N_28349);
and U28724 (N_28724,N_28434,N_28402);
nand U28725 (N_28725,N_28200,N_28330);
xnor U28726 (N_28726,N_28277,N_28248);
nand U28727 (N_28727,N_28333,N_28471);
nor U28728 (N_28728,N_28421,N_28431);
and U28729 (N_28729,N_28469,N_28459);
xor U28730 (N_28730,N_28452,N_28328);
nand U28731 (N_28731,N_28211,N_28375);
nor U28732 (N_28732,N_28343,N_28424);
nand U28733 (N_28733,N_28338,N_28226);
nor U28734 (N_28734,N_28215,N_28495);
nor U28735 (N_28735,N_28465,N_28431);
and U28736 (N_28736,N_28406,N_28274);
nor U28737 (N_28737,N_28464,N_28337);
or U28738 (N_28738,N_28489,N_28294);
or U28739 (N_28739,N_28234,N_28307);
xnor U28740 (N_28740,N_28424,N_28383);
nor U28741 (N_28741,N_28473,N_28246);
xor U28742 (N_28742,N_28471,N_28477);
nand U28743 (N_28743,N_28427,N_28336);
nand U28744 (N_28744,N_28433,N_28305);
nand U28745 (N_28745,N_28230,N_28243);
or U28746 (N_28746,N_28227,N_28408);
xnor U28747 (N_28747,N_28311,N_28471);
nor U28748 (N_28748,N_28247,N_28315);
xnor U28749 (N_28749,N_28364,N_28268);
nand U28750 (N_28750,N_28494,N_28388);
nor U28751 (N_28751,N_28460,N_28476);
nor U28752 (N_28752,N_28438,N_28437);
xor U28753 (N_28753,N_28233,N_28276);
nor U28754 (N_28754,N_28491,N_28265);
nor U28755 (N_28755,N_28333,N_28261);
nand U28756 (N_28756,N_28206,N_28290);
nand U28757 (N_28757,N_28405,N_28308);
or U28758 (N_28758,N_28342,N_28469);
or U28759 (N_28759,N_28455,N_28249);
and U28760 (N_28760,N_28214,N_28379);
xnor U28761 (N_28761,N_28204,N_28451);
nor U28762 (N_28762,N_28228,N_28403);
or U28763 (N_28763,N_28361,N_28252);
and U28764 (N_28764,N_28376,N_28301);
or U28765 (N_28765,N_28325,N_28330);
nor U28766 (N_28766,N_28205,N_28470);
nor U28767 (N_28767,N_28224,N_28454);
nor U28768 (N_28768,N_28381,N_28281);
xor U28769 (N_28769,N_28357,N_28299);
or U28770 (N_28770,N_28211,N_28346);
xnor U28771 (N_28771,N_28324,N_28226);
nor U28772 (N_28772,N_28439,N_28337);
nor U28773 (N_28773,N_28251,N_28450);
or U28774 (N_28774,N_28226,N_28355);
or U28775 (N_28775,N_28207,N_28271);
xnor U28776 (N_28776,N_28472,N_28476);
and U28777 (N_28777,N_28381,N_28322);
and U28778 (N_28778,N_28254,N_28205);
nor U28779 (N_28779,N_28464,N_28438);
or U28780 (N_28780,N_28257,N_28473);
nand U28781 (N_28781,N_28424,N_28378);
and U28782 (N_28782,N_28282,N_28455);
or U28783 (N_28783,N_28300,N_28399);
nand U28784 (N_28784,N_28353,N_28208);
or U28785 (N_28785,N_28346,N_28364);
nand U28786 (N_28786,N_28438,N_28311);
nor U28787 (N_28787,N_28394,N_28341);
and U28788 (N_28788,N_28473,N_28265);
and U28789 (N_28789,N_28310,N_28477);
xor U28790 (N_28790,N_28404,N_28209);
nand U28791 (N_28791,N_28342,N_28474);
nor U28792 (N_28792,N_28299,N_28479);
and U28793 (N_28793,N_28472,N_28314);
and U28794 (N_28794,N_28406,N_28212);
and U28795 (N_28795,N_28499,N_28306);
nor U28796 (N_28796,N_28280,N_28396);
and U28797 (N_28797,N_28485,N_28262);
and U28798 (N_28798,N_28312,N_28352);
xnor U28799 (N_28799,N_28383,N_28478);
nand U28800 (N_28800,N_28507,N_28621);
nor U28801 (N_28801,N_28768,N_28628);
nand U28802 (N_28802,N_28648,N_28765);
xor U28803 (N_28803,N_28744,N_28565);
xor U28804 (N_28804,N_28559,N_28572);
xnor U28805 (N_28805,N_28767,N_28764);
or U28806 (N_28806,N_28723,N_28635);
nor U28807 (N_28807,N_28755,N_28590);
nand U28808 (N_28808,N_28567,N_28583);
nor U28809 (N_28809,N_28550,N_28784);
and U28810 (N_28810,N_28694,N_28704);
xnor U28811 (N_28811,N_28541,N_28643);
or U28812 (N_28812,N_28525,N_28763);
xor U28813 (N_28813,N_28523,N_28734);
nand U28814 (N_28814,N_28515,N_28516);
nand U28815 (N_28815,N_28672,N_28595);
or U28816 (N_28816,N_28599,N_28699);
nand U28817 (N_28817,N_28759,N_28573);
nand U28818 (N_28818,N_28613,N_28529);
nand U28819 (N_28819,N_28540,N_28773);
xnor U28820 (N_28820,N_28714,N_28566);
nand U28821 (N_28821,N_28782,N_28616);
nand U28822 (N_28822,N_28524,N_28553);
nand U28823 (N_28823,N_28504,N_28710);
nor U28824 (N_28824,N_28546,N_28799);
nor U28825 (N_28825,N_28508,N_28600);
nand U28826 (N_28826,N_28568,N_28646);
nand U28827 (N_28827,N_28593,N_28551);
nand U28828 (N_28828,N_28754,N_28554);
xnor U28829 (N_28829,N_28794,N_28732);
nand U28830 (N_28830,N_28711,N_28667);
or U28831 (N_28831,N_28776,N_28601);
and U28832 (N_28832,N_28505,N_28531);
nand U28833 (N_28833,N_28629,N_28545);
nand U28834 (N_28834,N_28502,N_28522);
xnor U28835 (N_28835,N_28530,N_28611);
or U28836 (N_28836,N_28618,N_28577);
xnor U28837 (N_28837,N_28552,N_28663);
xor U28838 (N_28838,N_28771,N_28544);
xnor U28839 (N_28839,N_28693,N_28718);
and U28840 (N_28840,N_28514,N_28602);
nor U28841 (N_28841,N_28561,N_28675);
or U28842 (N_28842,N_28781,N_28509);
and U28843 (N_28843,N_28574,N_28517);
nand U28844 (N_28844,N_28708,N_28797);
nor U28845 (N_28845,N_28757,N_28780);
and U28846 (N_28846,N_28690,N_28564);
or U28847 (N_28847,N_28790,N_28549);
and U28848 (N_28848,N_28778,N_28625);
and U28849 (N_28849,N_28696,N_28659);
and U28850 (N_28850,N_28604,N_28580);
nand U28851 (N_28851,N_28735,N_28706);
nor U28852 (N_28852,N_28686,N_28584);
xor U28853 (N_28853,N_28518,N_28692);
nor U28854 (N_28854,N_28715,N_28679);
and U28855 (N_28855,N_28750,N_28656);
nand U28856 (N_28856,N_28683,N_28701);
nor U28857 (N_28857,N_28615,N_28520);
nand U28858 (N_28858,N_28664,N_28647);
nor U28859 (N_28859,N_28669,N_28747);
nor U28860 (N_28860,N_28680,N_28570);
or U28861 (N_28861,N_28649,N_28605);
xnor U28862 (N_28862,N_28527,N_28576);
or U28863 (N_28863,N_28607,N_28660);
nand U28864 (N_28864,N_28684,N_28737);
nor U28865 (N_28865,N_28758,N_28627);
or U28866 (N_28866,N_28637,N_28779);
xor U28867 (N_28867,N_28712,N_28740);
nand U28868 (N_28868,N_28724,N_28623);
xnor U28869 (N_28869,N_28519,N_28700);
or U28870 (N_28870,N_28741,N_28538);
nor U28871 (N_28871,N_28762,N_28796);
and U28872 (N_28872,N_28707,N_28521);
nor U28873 (N_28873,N_28671,N_28639);
xnor U28874 (N_28874,N_28719,N_28526);
nand U28875 (N_28875,N_28716,N_28681);
and U28876 (N_28876,N_28726,N_28555);
xnor U28877 (N_28877,N_28745,N_28752);
xor U28878 (N_28878,N_28528,N_28666);
or U28879 (N_28879,N_28636,N_28542);
nor U28880 (N_28880,N_28697,N_28589);
nand U28881 (N_28881,N_28506,N_28617);
or U28882 (N_28882,N_28575,N_28569);
nand U28883 (N_28883,N_28634,N_28563);
and U28884 (N_28884,N_28727,N_28748);
nand U28885 (N_28885,N_28620,N_28788);
nand U28886 (N_28886,N_28743,N_28560);
and U28887 (N_28887,N_28674,N_28582);
nand U28888 (N_28888,N_28720,N_28698);
or U28889 (N_28889,N_28775,N_28500);
and U28890 (N_28890,N_28537,N_28606);
nor U28891 (N_28891,N_28774,N_28614);
nor U28892 (N_28892,N_28597,N_28705);
and U28893 (N_28893,N_28792,N_28512);
or U28894 (N_28894,N_28543,N_28766);
or U28895 (N_28895,N_28688,N_28548);
and U28896 (N_28896,N_28731,N_28510);
or U28897 (N_28897,N_28562,N_28685);
or U28898 (N_28898,N_28655,N_28594);
and U28899 (N_28899,N_28725,N_28558);
nand U28900 (N_28900,N_28578,N_28678);
xor U28901 (N_28901,N_28676,N_28689);
xnor U28902 (N_28902,N_28603,N_28652);
nor U28903 (N_28903,N_28587,N_28702);
nand U28904 (N_28904,N_28749,N_28695);
xnor U28905 (N_28905,N_28626,N_28783);
xor U28906 (N_28906,N_28772,N_28592);
nand U28907 (N_28907,N_28795,N_28556);
nand U28908 (N_28908,N_28728,N_28619);
nor U28909 (N_28909,N_28662,N_28585);
nand U28910 (N_28910,N_28756,N_28703);
nor U28911 (N_28911,N_28588,N_28557);
xor U28912 (N_28912,N_28691,N_28612);
or U28913 (N_28913,N_28677,N_28532);
nand U28914 (N_28914,N_28746,N_28798);
nor U28915 (N_28915,N_28729,N_28769);
xnor U28916 (N_28916,N_28608,N_28730);
and U28917 (N_28917,N_28736,N_28630);
and U28918 (N_28918,N_28642,N_28591);
nand U28919 (N_28919,N_28709,N_28761);
xor U28920 (N_28920,N_28622,N_28624);
or U28921 (N_28921,N_28658,N_28596);
nand U28922 (N_28922,N_28610,N_28793);
nand U28923 (N_28923,N_28738,N_28581);
xnor U28924 (N_28924,N_28503,N_28534);
xor U28925 (N_28925,N_28770,N_28644);
and U28926 (N_28926,N_28598,N_28511);
xnor U28927 (N_28927,N_28722,N_28645);
nor U28928 (N_28928,N_28539,N_28791);
or U28929 (N_28929,N_28668,N_28641);
and U28930 (N_28930,N_28753,N_28651);
and U28931 (N_28931,N_28721,N_28682);
or U28932 (N_28932,N_28609,N_28787);
or U28933 (N_28933,N_28654,N_28535);
nor U28934 (N_28934,N_28751,N_28547);
nor U28935 (N_28935,N_28733,N_28777);
nand U28936 (N_28936,N_28742,N_28533);
and U28937 (N_28937,N_28501,N_28670);
nor U28938 (N_28938,N_28665,N_28571);
xnor U28939 (N_28939,N_28632,N_28717);
and U28940 (N_28940,N_28789,N_28786);
nand U28941 (N_28941,N_28653,N_28586);
and U28942 (N_28942,N_28513,N_28650);
and U28943 (N_28943,N_28760,N_28661);
nor U28944 (N_28944,N_28638,N_28536);
xnor U28945 (N_28945,N_28673,N_28631);
xnor U28946 (N_28946,N_28640,N_28633);
or U28947 (N_28947,N_28785,N_28739);
xnor U28948 (N_28948,N_28713,N_28687);
and U28949 (N_28949,N_28579,N_28657);
or U28950 (N_28950,N_28710,N_28535);
nor U28951 (N_28951,N_28796,N_28545);
nand U28952 (N_28952,N_28776,N_28567);
and U28953 (N_28953,N_28520,N_28677);
and U28954 (N_28954,N_28526,N_28718);
nand U28955 (N_28955,N_28695,N_28756);
or U28956 (N_28956,N_28679,N_28731);
xnor U28957 (N_28957,N_28562,N_28736);
xnor U28958 (N_28958,N_28688,N_28622);
nor U28959 (N_28959,N_28622,N_28754);
and U28960 (N_28960,N_28698,N_28651);
nor U28961 (N_28961,N_28506,N_28651);
xnor U28962 (N_28962,N_28576,N_28765);
or U28963 (N_28963,N_28525,N_28600);
nand U28964 (N_28964,N_28625,N_28665);
or U28965 (N_28965,N_28530,N_28569);
nand U28966 (N_28966,N_28560,N_28606);
or U28967 (N_28967,N_28760,N_28633);
or U28968 (N_28968,N_28547,N_28654);
nand U28969 (N_28969,N_28625,N_28717);
xor U28970 (N_28970,N_28502,N_28546);
or U28971 (N_28971,N_28764,N_28505);
nor U28972 (N_28972,N_28662,N_28716);
nand U28973 (N_28973,N_28583,N_28785);
and U28974 (N_28974,N_28673,N_28795);
and U28975 (N_28975,N_28508,N_28799);
xor U28976 (N_28976,N_28621,N_28755);
and U28977 (N_28977,N_28506,N_28639);
and U28978 (N_28978,N_28679,N_28699);
xor U28979 (N_28979,N_28702,N_28513);
or U28980 (N_28980,N_28677,N_28753);
or U28981 (N_28981,N_28676,N_28765);
or U28982 (N_28982,N_28735,N_28618);
or U28983 (N_28983,N_28688,N_28734);
xnor U28984 (N_28984,N_28625,N_28789);
xnor U28985 (N_28985,N_28694,N_28544);
or U28986 (N_28986,N_28510,N_28622);
or U28987 (N_28987,N_28662,N_28529);
nor U28988 (N_28988,N_28544,N_28700);
xor U28989 (N_28989,N_28735,N_28660);
and U28990 (N_28990,N_28563,N_28571);
nand U28991 (N_28991,N_28519,N_28778);
nor U28992 (N_28992,N_28754,N_28570);
nor U28993 (N_28993,N_28617,N_28736);
or U28994 (N_28994,N_28740,N_28714);
nor U28995 (N_28995,N_28570,N_28539);
xor U28996 (N_28996,N_28504,N_28601);
nor U28997 (N_28997,N_28759,N_28625);
and U28998 (N_28998,N_28706,N_28534);
nor U28999 (N_28999,N_28723,N_28586);
or U29000 (N_29000,N_28728,N_28532);
or U29001 (N_29001,N_28619,N_28755);
nand U29002 (N_29002,N_28696,N_28543);
nor U29003 (N_29003,N_28602,N_28636);
nand U29004 (N_29004,N_28727,N_28663);
or U29005 (N_29005,N_28524,N_28631);
or U29006 (N_29006,N_28535,N_28570);
xor U29007 (N_29007,N_28513,N_28780);
nand U29008 (N_29008,N_28578,N_28543);
and U29009 (N_29009,N_28586,N_28551);
nor U29010 (N_29010,N_28555,N_28581);
and U29011 (N_29011,N_28743,N_28605);
and U29012 (N_29012,N_28741,N_28630);
and U29013 (N_29013,N_28730,N_28653);
or U29014 (N_29014,N_28578,N_28709);
xnor U29015 (N_29015,N_28655,N_28699);
or U29016 (N_29016,N_28523,N_28780);
and U29017 (N_29017,N_28712,N_28512);
nor U29018 (N_29018,N_28629,N_28795);
or U29019 (N_29019,N_28540,N_28516);
and U29020 (N_29020,N_28550,N_28541);
xnor U29021 (N_29021,N_28670,N_28791);
and U29022 (N_29022,N_28637,N_28575);
or U29023 (N_29023,N_28773,N_28745);
nand U29024 (N_29024,N_28567,N_28634);
xor U29025 (N_29025,N_28690,N_28696);
and U29026 (N_29026,N_28548,N_28657);
xnor U29027 (N_29027,N_28735,N_28603);
and U29028 (N_29028,N_28704,N_28791);
nand U29029 (N_29029,N_28760,N_28766);
xnor U29030 (N_29030,N_28733,N_28501);
and U29031 (N_29031,N_28526,N_28695);
nor U29032 (N_29032,N_28669,N_28634);
xor U29033 (N_29033,N_28693,N_28647);
xnor U29034 (N_29034,N_28616,N_28501);
nor U29035 (N_29035,N_28719,N_28767);
and U29036 (N_29036,N_28793,N_28707);
nand U29037 (N_29037,N_28796,N_28651);
nor U29038 (N_29038,N_28767,N_28717);
nand U29039 (N_29039,N_28511,N_28602);
xnor U29040 (N_29040,N_28781,N_28744);
nor U29041 (N_29041,N_28692,N_28766);
nor U29042 (N_29042,N_28776,N_28572);
xor U29043 (N_29043,N_28607,N_28647);
xor U29044 (N_29044,N_28692,N_28519);
or U29045 (N_29045,N_28597,N_28661);
nand U29046 (N_29046,N_28625,N_28608);
nand U29047 (N_29047,N_28676,N_28519);
xnor U29048 (N_29048,N_28778,N_28557);
or U29049 (N_29049,N_28691,N_28748);
nand U29050 (N_29050,N_28617,N_28569);
nand U29051 (N_29051,N_28525,N_28548);
and U29052 (N_29052,N_28520,N_28735);
nor U29053 (N_29053,N_28502,N_28739);
nor U29054 (N_29054,N_28736,N_28769);
and U29055 (N_29055,N_28502,N_28763);
and U29056 (N_29056,N_28645,N_28697);
or U29057 (N_29057,N_28750,N_28652);
or U29058 (N_29058,N_28596,N_28705);
nor U29059 (N_29059,N_28778,N_28771);
or U29060 (N_29060,N_28675,N_28734);
nand U29061 (N_29061,N_28740,N_28577);
nand U29062 (N_29062,N_28524,N_28572);
or U29063 (N_29063,N_28591,N_28669);
or U29064 (N_29064,N_28641,N_28799);
nand U29065 (N_29065,N_28747,N_28686);
nor U29066 (N_29066,N_28502,N_28788);
nor U29067 (N_29067,N_28623,N_28525);
xor U29068 (N_29068,N_28534,N_28713);
and U29069 (N_29069,N_28778,N_28709);
or U29070 (N_29070,N_28640,N_28631);
and U29071 (N_29071,N_28566,N_28593);
or U29072 (N_29072,N_28652,N_28755);
xnor U29073 (N_29073,N_28527,N_28504);
xnor U29074 (N_29074,N_28613,N_28516);
nor U29075 (N_29075,N_28558,N_28749);
or U29076 (N_29076,N_28767,N_28600);
xor U29077 (N_29077,N_28744,N_28660);
or U29078 (N_29078,N_28681,N_28639);
or U29079 (N_29079,N_28502,N_28521);
xor U29080 (N_29080,N_28531,N_28547);
nand U29081 (N_29081,N_28628,N_28667);
and U29082 (N_29082,N_28676,N_28741);
and U29083 (N_29083,N_28723,N_28550);
nand U29084 (N_29084,N_28608,N_28562);
xnor U29085 (N_29085,N_28738,N_28698);
nor U29086 (N_29086,N_28741,N_28550);
nor U29087 (N_29087,N_28620,N_28658);
nor U29088 (N_29088,N_28696,N_28674);
nor U29089 (N_29089,N_28507,N_28663);
nand U29090 (N_29090,N_28564,N_28684);
or U29091 (N_29091,N_28659,N_28503);
nor U29092 (N_29092,N_28551,N_28626);
or U29093 (N_29093,N_28790,N_28748);
nor U29094 (N_29094,N_28774,N_28644);
or U29095 (N_29095,N_28683,N_28751);
or U29096 (N_29096,N_28728,N_28757);
nand U29097 (N_29097,N_28774,N_28590);
nand U29098 (N_29098,N_28673,N_28578);
nand U29099 (N_29099,N_28613,N_28603);
nand U29100 (N_29100,N_28963,N_28984);
and U29101 (N_29101,N_28856,N_28947);
nor U29102 (N_29102,N_29060,N_28944);
xor U29103 (N_29103,N_28999,N_29095);
xor U29104 (N_29104,N_29058,N_28970);
or U29105 (N_29105,N_28985,N_29065);
xor U29106 (N_29106,N_28954,N_28829);
nor U29107 (N_29107,N_28868,N_28859);
xor U29108 (N_29108,N_29082,N_28835);
and U29109 (N_29109,N_28851,N_28857);
nor U29110 (N_29110,N_29089,N_29024);
and U29111 (N_29111,N_28921,N_28839);
and U29112 (N_29112,N_29075,N_28909);
and U29113 (N_29113,N_28973,N_28917);
xor U29114 (N_29114,N_28802,N_28831);
and U29115 (N_29115,N_28866,N_29009);
and U29116 (N_29116,N_28879,N_28939);
or U29117 (N_29117,N_28867,N_28886);
nand U29118 (N_29118,N_28925,N_29015);
xnor U29119 (N_29119,N_29054,N_29079);
or U29120 (N_29120,N_29043,N_28942);
and U29121 (N_29121,N_28920,N_28957);
nor U29122 (N_29122,N_28924,N_28810);
xnor U29123 (N_29123,N_29038,N_29094);
xor U29124 (N_29124,N_28908,N_29007);
nor U29125 (N_29125,N_28896,N_29053);
or U29126 (N_29126,N_29077,N_28864);
nand U29127 (N_29127,N_28847,N_29088);
nor U29128 (N_29128,N_29031,N_28823);
nand U29129 (N_29129,N_29049,N_28885);
or U29130 (N_29130,N_29001,N_28865);
or U29131 (N_29131,N_29022,N_29018);
nand U29132 (N_29132,N_28949,N_28837);
xor U29133 (N_29133,N_28931,N_28993);
xnor U29134 (N_29134,N_28907,N_28982);
nor U29135 (N_29135,N_28858,N_28945);
nand U29136 (N_29136,N_29008,N_28998);
or U29137 (N_29137,N_28843,N_29037);
nor U29138 (N_29138,N_28912,N_29061);
or U29139 (N_29139,N_28995,N_28933);
xor U29140 (N_29140,N_28891,N_28961);
xor U29141 (N_29141,N_28978,N_28874);
nand U29142 (N_29142,N_29035,N_28911);
nor U29143 (N_29143,N_28811,N_28934);
nor U29144 (N_29144,N_29003,N_29011);
or U29145 (N_29145,N_29039,N_29067);
xor U29146 (N_29146,N_28930,N_28997);
xnor U29147 (N_29147,N_29002,N_28923);
nor U29148 (N_29148,N_28817,N_29032);
xnor U29149 (N_29149,N_28910,N_28878);
nand U29150 (N_29150,N_28992,N_28893);
nand U29151 (N_29151,N_28950,N_28850);
xor U29152 (N_29152,N_28832,N_29052);
and U29153 (N_29153,N_28935,N_29017);
and U29154 (N_29154,N_28914,N_28814);
nor U29155 (N_29155,N_29026,N_29096);
or U29156 (N_29156,N_28975,N_28894);
nor U29157 (N_29157,N_29041,N_28827);
or U29158 (N_29158,N_28861,N_28953);
nor U29159 (N_29159,N_29059,N_28981);
nor U29160 (N_29160,N_29062,N_28880);
or U29161 (N_29161,N_28951,N_28876);
or U29162 (N_29162,N_28972,N_28964);
nand U29163 (N_29163,N_29080,N_28956);
nand U29164 (N_29164,N_28889,N_28980);
or U29165 (N_29165,N_28820,N_28812);
xnor U29166 (N_29166,N_28884,N_28840);
nor U29167 (N_29167,N_28943,N_28853);
and U29168 (N_29168,N_28989,N_28826);
xor U29169 (N_29169,N_28875,N_28825);
or U29170 (N_29170,N_29005,N_28870);
and U29171 (N_29171,N_28929,N_28815);
nand U29172 (N_29172,N_29081,N_28994);
and U29173 (N_29173,N_28807,N_28897);
or U29174 (N_29174,N_28872,N_28960);
nand U29175 (N_29175,N_28854,N_28828);
and U29176 (N_29176,N_29021,N_29012);
and U29177 (N_29177,N_29093,N_28986);
xor U29178 (N_29178,N_28813,N_28955);
xor U29179 (N_29179,N_28983,N_29025);
nand U29180 (N_29180,N_28824,N_28969);
and U29181 (N_29181,N_28927,N_29090);
xnor U29182 (N_29182,N_29083,N_29070);
or U29183 (N_29183,N_29076,N_28821);
xnor U29184 (N_29184,N_28901,N_28882);
xor U29185 (N_29185,N_28845,N_29027);
nand U29186 (N_29186,N_29040,N_29056);
or U29187 (N_29187,N_29064,N_29014);
xnor U29188 (N_29188,N_29048,N_28852);
or U29189 (N_29189,N_28898,N_28869);
nand U29190 (N_29190,N_28948,N_28819);
nor U29191 (N_29191,N_28892,N_28838);
nor U29192 (N_29192,N_28979,N_29050);
xor U29193 (N_29193,N_28900,N_28836);
nand U29194 (N_29194,N_28906,N_28941);
nor U29195 (N_29195,N_28855,N_29084);
or U29196 (N_29196,N_29033,N_28881);
nor U29197 (N_29197,N_28806,N_28805);
and U29198 (N_29198,N_29029,N_28996);
nand U29199 (N_29199,N_29000,N_29087);
xnor U29200 (N_29200,N_29055,N_29023);
xor U29201 (N_29201,N_28818,N_28905);
xor U29202 (N_29202,N_29086,N_28940);
xnor U29203 (N_29203,N_28976,N_28959);
or U29204 (N_29204,N_28966,N_29028);
nor U29205 (N_29205,N_28863,N_29051);
nand U29206 (N_29206,N_28877,N_29044);
xnor U29207 (N_29207,N_29098,N_28903);
nor U29208 (N_29208,N_28977,N_28803);
nor U29209 (N_29209,N_28974,N_28873);
or U29210 (N_29210,N_28846,N_28860);
nor U29211 (N_29211,N_28958,N_29099);
nand U29212 (N_29212,N_28987,N_29057);
xor U29213 (N_29213,N_28990,N_28952);
or U29214 (N_29214,N_28988,N_29068);
nand U29215 (N_29215,N_28918,N_28926);
xnor U29216 (N_29216,N_29092,N_28965);
and U29217 (N_29217,N_29030,N_28919);
nand U29218 (N_29218,N_28871,N_29046);
xor U29219 (N_29219,N_29063,N_28895);
xor U29220 (N_29220,N_29071,N_28830);
or U29221 (N_29221,N_28841,N_29013);
xnor U29222 (N_29222,N_29045,N_28928);
or U29223 (N_29223,N_29034,N_29085);
or U29224 (N_29224,N_28915,N_28800);
or U29225 (N_29225,N_29010,N_29073);
and U29226 (N_29226,N_28904,N_28801);
nand U29227 (N_29227,N_28967,N_28833);
nand U29228 (N_29228,N_29042,N_28902);
xor U29229 (N_29229,N_28804,N_28968);
xor U29230 (N_29230,N_28913,N_29066);
and U29231 (N_29231,N_28842,N_28936);
xor U29232 (N_29232,N_28834,N_28932);
xnor U29233 (N_29233,N_29006,N_28991);
and U29234 (N_29234,N_28938,N_28848);
and U29235 (N_29235,N_28862,N_28887);
xnor U29236 (N_29236,N_28899,N_29047);
nand U29237 (N_29237,N_29016,N_28937);
and U29238 (N_29238,N_28971,N_29019);
and U29239 (N_29239,N_28916,N_29004);
and U29240 (N_29240,N_29020,N_28890);
xor U29241 (N_29241,N_29072,N_28922);
xor U29242 (N_29242,N_29074,N_29091);
nor U29243 (N_29243,N_29097,N_28962);
nor U29244 (N_29244,N_29069,N_28816);
or U29245 (N_29245,N_28888,N_29078);
xnor U29246 (N_29246,N_28808,N_28809);
and U29247 (N_29247,N_28844,N_29036);
and U29248 (N_29248,N_28849,N_28883);
xor U29249 (N_29249,N_28946,N_28822);
or U29250 (N_29250,N_28934,N_28886);
nand U29251 (N_29251,N_29061,N_29088);
and U29252 (N_29252,N_28833,N_28907);
or U29253 (N_29253,N_29084,N_28875);
nor U29254 (N_29254,N_29030,N_29006);
nand U29255 (N_29255,N_28811,N_28898);
xnor U29256 (N_29256,N_28959,N_28900);
nor U29257 (N_29257,N_29019,N_29036);
or U29258 (N_29258,N_28859,N_28834);
xor U29259 (N_29259,N_28919,N_28905);
and U29260 (N_29260,N_28962,N_28943);
nand U29261 (N_29261,N_28944,N_29048);
and U29262 (N_29262,N_29004,N_28831);
nor U29263 (N_29263,N_28800,N_29022);
or U29264 (N_29264,N_29049,N_28942);
xnor U29265 (N_29265,N_29053,N_29036);
nor U29266 (N_29266,N_28937,N_29071);
and U29267 (N_29267,N_28866,N_29002);
nor U29268 (N_29268,N_28964,N_28980);
or U29269 (N_29269,N_29043,N_28984);
or U29270 (N_29270,N_28990,N_28856);
and U29271 (N_29271,N_28890,N_28993);
and U29272 (N_29272,N_28854,N_28964);
or U29273 (N_29273,N_28930,N_28838);
nand U29274 (N_29274,N_29038,N_28852);
xnor U29275 (N_29275,N_28956,N_28859);
xor U29276 (N_29276,N_29029,N_28871);
and U29277 (N_29277,N_29012,N_29048);
or U29278 (N_29278,N_28819,N_28846);
nand U29279 (N_29279,N_28996,N_28938);
nand U29280 (N_29280,N_29084,N_28921);
nand U29281 (N_29281,N_28867,N_29075);
xnor U29282 (N_29282,N_28935,N_28938);
or U29283 (N_29283,N_29020,N_29081);
and U29284 (N_29284,N_28955,N_28867);
xor U29285 (N_29285,N_28826,N_29097);
or U29286 (N_29286,N_28925,N_28872);
and U29287 (N_29287,N_29046,N_29092);
or U29288 (N_29288,N_28923,N_28871);
nor U29289 (N_29289,N_28860,N_28865);
nand U29290 (N_29290,N_29028,N_28873);
nand U29291 (N_29291,N_28864,N_29013);
xor U29292 (N_29292,N_28840,N_28990);
nor U29293 (N_29293,N_28918,N_28982);
nor U29294 (N_29294,N_29055,N_28874);
nand U29295 (N_29295,N_28986,N_29061);
and U29296 (N_29296,N_28868,N_28838);
and U29297 (N_29297,N_28846,N_28997);
nor U29298 (N_29298,N_28934,N_28890);
xor U29299 (N_29299,N_29045,N_29008);
or U29300 (N_29300,N_28932,N_29005);
and U29301 (N_29301,N_29032,N_28843);
nor U29302 (N_29302,N_28924,N_28834);
nand U29303 (N_29303,N_28839,N_28846);
nor U29304 (N_29304,N_29045,N_28983);
nor U29305 (N_29305,N_28880,N_28928);
nand U29306 (N_29306,N_28983,N_28809);
nand U29307 (N_29307,N_28972,N_29086);
nand U29308 (N_29308,N_28837,N_28812);
nor U29309 (N_29309,N_29091,N_29018);
and U29310 (N_29310,N_29020,N_28875);
and U29311 (N_29311,N_28895,N_29059);
xor U29312 (N_29312,N_28998,N_28930);
nand U29313 (N_29313,N_28828,N_29066);
nor U29314 (N_29314,N_28970,N_29099);
nor U29315 (N_29315,N_28868,N_28883);
nor U29316 (N_29316,N_28904,N_28830);
xor U29317 (N_29317,N_28919,N_28920);
xnor U29318 (N_29318,N_28820,N_28979);
and U29319 (N_29319,N_28872,N_28890);
and U29320 (N_29320,N_29098,N_28817);
or U29321 (N_29321,N_28875,N_28942);
or U29322 (N_29322,N_29064,N_28902);
nor U29323 (N_29323,N_28967,N_28988);
or U29324 (N_29324,N_28909,N_29022);
nor U29325 (N_29325,N_28895,N_29039);
or U29326 (N_29326,N_29067,N_28834);
or U29327 (N_29327,N_28923,N_28999);
xnor U29328 (N_29328,N_29040,N_28861);
nand U29329 (N_29329,N_28936,N_28836);
nand U29330 (N_29330,N_28992,N_28996);
nor U29331 (N_29331,N_28880,N_28971);
nand U29332 (N_29332,N_29054,N_28981);
nand U29333 (N_29333,N_28882,N_28955);
nand U29334 (N_29334,N_29078,N_28910);
nand U29335 (N_29335,N_29048,N_28890);
nor U29336 (N_29336,N_29008,N_28971);
and U29337 (N_29337,N_29061,N_29059);
xnor U29338 (N_29338,N_28841,N_29016);
xor U29339 (N_29339,N_28905,N_28855);
nor U29340 (N_29340,N_28963,N_28940);
or U29341 (N_29341,N_29065,N_28838);
or U29342 (N_29342,N_28962,N_28927);
or U29343 (N_29343,N_29059,N_28919);
nor U29344 (N_29344,N_28947,N_28914);
xor U29345 (N_29345,N_28960,N_28832);
or U29346 (N_29346,N_28906,N_28922);
or U29347 (N_29347,N_28980,N_29021);
nand U29348 (N_29348,N_28969,N_28880);
xor U29349 (N_29349,N_28985,N_28905);
nor U29350 (N_29350,N_28993,N_29096);
and U29351 (N_29351,N_28969,N_28970);
or U29352 (N_29352,N_29081,N_28836);
or U29353 (N_29353,N_28999,N_28983);
nand U29354 (N_29354,N_29050,N_28841);
and U29355 (N_29355,N_28811,N_28808);
or U29356 (N_29356,N_28825,N_28899);
xor U29357 (N_29357,N_29008,N_28938);
xnor U29358 (N_29358,N_29081,N_29087);
or U29359 (N_29359,N_29023,N_28943);
nor U29360 (N_29360,N_28802,N_28922);
xnor U29361 (N_29361,N_28820,N_28953);
and U29362 (N_29362,N_29056,N_28970);
nand U29363 (N_29363,N_28913,N_28953);
xnor U29364 (N_29364,N_29091,N_28953);
and U29365 (N_29365,N_29019,N_29097);
nor U29366 (N_29366,N_29025,N_29034);
and U29367 (N_29367,N_29036,N_28804);
nand U29368 (N_29368,N_28845,N_29058);
nor U29369 (N_29369,N_29044,N_29053);
or U29370 (N_29370,N_29051,N_28920);
or U29371 (N_29371,N_29031,N_28862);
or U29372 (N_29372,N_29058,N_28841);
or U29373 (N_29373,N_28914,N_28928);
nor U29374 (N_29374,N_28817,N_28946);
xor U29375 (N_29375,N_28845,N_28849);
and U29376 (N_29376,N_28978,N_28963);
nand U29377 (N_29377,N_29094,N_28972);
xnor U29378 (N_29378,N_29069,N_29045);
and U29379 (N_29379,N_28861,N_28975);
and U29380 (N_29380,N_28888,N_28909);
xnor U29381 (N_29381,N_29037,N_28977);
or U29382 (N_29382,N_28879,N_28976);
or U29383 (N_29383,N_28890,N_29054);
nor U29384 (N_29384,N_28806,N_29040);
or U29385 (N_29385,N_28973,N_28807);
nor U29386 (N_29386,N_28850,N_28802);
nand U29387 (N_29387,N_28893,N_28967);
nand U29388 (N_29388,N_28815,N_28927);
nor U29389 (N_29389,N_28941,N_29048);
and U29390 (N_29390,N_29027,N_29055);
and U29391 (N_29391,N_29088,N_29044);
xnor U29392 (N_29392,N_28821,N_28831);
and U29393 (N_29393,N_29028,N_28902);
or U29394 (N_29394,N_28914,N_29062);
and U29395 (N_29395,N_28997,N_28957);
nor U29396 (N_29396,N_28844,N_28935);
nand U29397 (N_29397,N_29048,N_28848);
nand U29398 (N_29398,N_28875,N_28892);
and U29399 (N_29399,N_28855,N_29058);
nor U29400 (N_29400,N_29236,N_29183);
or U29401 (N_29401,N_29140,N_29277);
or U29402 (N_29402,N_29152,N_29393);
and U29403 (N_29403,N_29395,N_29282);
and U29404 (N_29404,N_29276,N_29122);
and U29405 (N_29405,N_29284,N_29392);
and U29406 (N_29406,N_29143,N_29255);
nand U29407 (N_29407,N_29220,N_29352);
and U29408 (N_29408,N_29253,N_29199);
or U29409 (N_29409,N_29307,N_29125);
xor U29410 (N_29410,N_29147,N_29138);
xnor U29411 (N_29411,N_29345,N_29113);
xnor U29412 (N_29412,N_29158,N_29268);
nor U29413 (N_29413,N_29322,N_29339);
nor U29414 (N_29414,N_29387,N_29356);
xnor U29415 (N_29415,N_29193,N_29161);
xor U29416 (N_29416,N_29285,N_29377);
or U29417 (N_29417,N_29132,N_29357);
nand U29418 (N_29418,N_29141,N_29351);
nand U29419 (N_29419,N_29270,N_29200);
nand U29420 (N_29420,N_29370,N_29226);
or U29421 (N_29421,N_29373,N_29251);
xor U29422 (N_29422,N_29330,N_29272);
nor U29423 (N_29423,N_29348,N_29361);
and U29424 (N_29424,N_29104,N_29308);
and U29425 (N_29425,N_29372,N_29157);
or U29426 (N_29426,N_29262,N_29365);
xnor U29427 (N_29427,N_29342,N_29165);
nand U29428 (N_29428,N_29368,N_29194);
and U29429 (N_29429,N_29114,N_29205);
nor U29430 (N_29430,N_29297,N_29190);
or U29431 (N_29431,N_29213,N_29232);
xor U29432 (N_29432,N_29206,N_29327);
nand U29433 (N_29433,N_29334,N_29210);
nor U29434 (N_29434,N_29292,N_29398);
nor U29435 (N_29435,N_29371,N_29310);
nand U29436 (N_29436,N_29128,N_29304);
xnor U29437 (N_29437,N_29344,N_29375);
nor U29438 (N_29438,N_29177,N_29159);
or U29439 (N_29439,N_29259,N_29329);
or U29440 (N_29440,N_29315,N_29328);
or U29441 (N_29441,N_29313,N_29211);
and U29442 (N_29442,N_29216,N_29376);
nor U29443 (N_29443,N_29135,N_29231);
or U29444 (N_29444,N_29233,N_29188);
or U29445 (N_29445,N_29399,N_29256);
or U29446 (N_29446,N_29127,N_29198);
and U29447 (N_29447,N_29353,N_29343);
or U29448 (N_29448,N_29337,N_29317);
nor U29449 (N_29449,N_29367,N_29303);
or U29450 (N_29450,N_29151,N_29153);
nand U29451 (N_29451,N_29112,N_29243);
and U29452 (N_29452,N_29212,N_29245);
and U29453 (N_29453,N_29316,N_29103);
nor U29454 (N_29454,N_29203,N_29336);
or U29455 (N_29455,N_29222,N_29111);
nand U29456 (N_29456,N_29115,N_29109);
xnor U29457 (N_29457,N_29293,N_29275);
nor U29458 (N_29458,N_29170,N_29230);
or U29459 (N_29459,N_29283,N_29228);
xor U29460 (N_29460,N_29129,N_29173);
or U29461 (N_29461,N_29287,N_29291);
nor U29462 (N_29462,N_29364,N_29269);
or U29463 (N_29463,N_29281,N_29130);
xor U29464 (N_29464,N_29207,N_29234);
nor U29465 (N_29465,N_29278,N_29389);
or U29466 (N_29466,N_29363,N_29145);
xnor U29467 (N_29467,N_29325,N_29358);
and U29468 (N_29468,N_29254,N_29175);
nor U29469 (N_29469,N_29182,N_29306);
xnor U29470 (N_29470,N_29340,N_29227);
xor U29471 (N_29471,N_29267,N_29362);
xor U29472 (N_29472,N_29390,N_29279);
nand U29473 (N_29473,N_29119,N_29181);
nor U29474 (N_29474,N_29369,N_29296);
nand U29475 (N_29475,N_29150,N_29397);
nand U29476 (N_29476,N_29381,N_29260);
nor U29477 (N_29477,N_29391,N_29106);
nor U29478 (N_29478,N_29101,N_29217);
or U29479 (N_29479,N_29380,N_29263);
and U29480 (N_29480,N_29202,N_29176);
nand U29481 (N_29481,N_29242,N_29289);
nor U29482 (N_29482,N_29108,N_29186);
nor U29483 (N_29483,N_29318,N_29288);
xor U29484 (N_29484,N_29335,N_29136);
and U29485 (N_29485,N_29218,N_29154);
xnor U29486 (N_29486,N_29331,N_29366);
xnor U29487 (N_29487,N_29346,N_29214);
xnor U29488 (N_29488,N_29384,N_29379);
xor U29489 (N_29489,N_29221,N_29238);
and U29490 (N_29490,N_29110,N_29219);
and U29491 (N_29491,N_29155,N_29169);
or U29492 (N_29492,N_29332,N_29144);
nor U29493 (N_29493,N_29388,N_29355);
nor U29494 (N_29494,N_29174,N_29160);
xor U29495 (N_29495,N_29225,N_29149);
or U29496 (N_29496,N_29298,N_29240);
xnor U29497 (N_29497,N_29142,N_29299);
and U29498 (N_29498,N_29187,N_29359);
xnor U29499 (N_29499,N_29273,N_29349);
or U29500 (N_29500,N_29264,N_29324);
and U29501 (N_29501,N_29396,N_29224);
or U29502 (N_29502,N_29146,N_29320);
xor U29503 (N_29503,N_29191,N_29178);
and U29504 (N_29504,N_29131,N_29139);
and U29505 (N_29505,N_29185,N_29168);
nand U29506 (N_29506,N_29350,N_29244);
nand U29507 (N_29507,N_29137,N_29148);
and U29508 (N_29508,N_29252,N_29166);
or U29509 (N_29509,N_29247,N_29126);
nor U29510 (N_29510,N_29338,N_29196);
nor U29511 (N_29511,N_29378,N_29265);
xnor U29512 (N_29512,N_29333,N_29167);
or U29513 (N_29513,N_29223,N_29347);
nand U29514 (N_29514,N_29123,N_29105);
and U29515 (N_29515,N_29360,N_29249);
nor U29516 (N_29516,N_29134,N_29250);
nor U29517 (N_29517,N_29102,N_29107);
and U29518 (N_29518,N_29208,N_29266);
and U29519 (N_29519,N_29302,N_29385);
xor U29520 (N_29520,N_29309,N_29189);
nand U29521 (N_29521,N_29323,N_29117);
nand U29522 (N_29522,N_29394,N_29305);
nand U29523 (N_29523,N_29118,N_29341);
nand U29524 (N_29524,N_29235,N_29156);
xnor U29525 (N_29525,N_29195,N_29172);
or U29526 (N_29526,N_29300,N_29257);
xnor U29527 (N_29527,N_29163,N_29274);
and U29528 (N_29528,N_29301,N_29180);
or U29529 (N_29529,N_29124,N_29171);
or U29530 (N_29530,N_29100,N_29164);
nand U29531 (N_29531,N_29201,N_29192);
xor U29532 (N_29532,N_29204,N_29383);
nand U29533 (N_29533,N_29248,N_29314);
nand U29534 (N_29534,N_29286,N_29116);
nand U29535 (N_29535,N_29162,N_29382);
xor U29536 (N_29536,N_29209,N_29239);
or U29537 (N_29537,N_29179,N_29290);
nand U29538 (N_29538,N_29241,N_29295);
nand U29539 (N_29539,N_29354,N_29374);
nand U29540 (N_29540,N_29280,N_29311);
xor U29541 (N_29541,N_29215,N_29197);
and U29542 (N_29542,N_29246,N_29258);
xor U29543 (N_29543,N_29271,N_29321);
or U29544 (N_29544,N_29386,N_29261);
or U29545 (N_29545,N_29120,N_29326);
or U29546 (N_29546,N_29237,N_29184);
xnor U29547 (N_29547,N_29133,N_29121);
and U29548 (N_29548,N_29229,N_29319);
nand U29549 (N_29549,N_29312,N_29294);
and U29550 (N_29550,N_29172,N_29284);
or U29551 (N_29551,N_29350,N_29268);
xor U29552 (N_29552,N_29353,N_29327);
xnor U29553 (N_29553,N_29317,N_29373);
xnor U29554 (N_29554,N_29368,N_29147);
nor U29555 (N_29555,N_29383,N_29159);
or U29556 (N_29556,N_29183,N_29357);
xor U29557 (N_29557,N_29304,N_29336);
xnor U29558 (N_29558,N_29178,N_29341);
xor U29559 (N_29559,N_29303,N_29199);
or U29560 (N_29560,N_29248,N_29365);
nand U29561 (N_29561,N_29273,N_29376);
nand U29562 (N_29562,N_29343,N_29357);
nand U29563 (N_29563,N_29168,N_29334);
nand U29564 (N_29564,N_29305,N_29229);
nor U29565 (N_29565,N_29398,N_29139);
nand U29566 (N_29566,N_29246,N_29272);
nor U29567 (N_29567,N_29392,N_29223);
and U29568 (N_29568,N_29252,N_29147);
xnor U29569 (N_29569,N_29180,N_29366);
or U29570 (N_29570,N_29131,N_29170);
xnor U29571 (N_29571,N_29263,N_29183);
and U29572 (N_29572,N_29344,N_29379);
nand U29573 (N_29573,N_29263,N_29348);
and U29574 (N_29574,N_29346,N_29302);
or U29575 (N_29575,N_29255,N_29284);
nand U29576 (N_29576,N_29361,N_29281);
nand U29577 (N_29577,N_29132,N_29173);
nand U29578 (N_29578,N_29383,N_29243);
or U29579 (N_29579,N_29186,N_29130);
nand U29580 (N_29580,N_29207,N_29206);
xor U29581 (N_29581,N_29209,N_29234);
nor U29582 (N_29582,N_29311,N_29316);
xor U29583 (N_29583,N_29299,N_29113);
nor U29584 (N_29584,N_29383,N_29207);
nand U29585 (N_29585,N_29108,N_29147);
or U29586 (N_29586,N_29276,N_29206);
or U29587 (N_29587,N_29151,N_29108);
nand U29588 (N_29588,N_29231,N_29338);
and U29589 (N_29589,N_29216,N_29359);
and U29590 (N_29590,N_29397,N_29148);
nand U29591 (N_29591,N_29346,N_29305);
nor U29592 (N_29592,N_29354,N_29365);
and U29593 (N_29593,N_29384,N_29195);
or U29594 (N_29594,N_29299,N_29153);
and U29595 (N_29595,N_29112,N_29183);
or U29596 (N_29596,N_29127,N_29267);
nand U29597 (N_29597,N_29236,N_29330);
and U29598 (N_29598,N_29131,N_29122);
and U29599 (N_29599,N_29163,N_29237);
or U29600 (N_29600,N_29320,N_29117);
or U29601 (N_29601,N_29244,N_29317);
nor U29602 (N_29602,N_29393,N_29353);
xnor U29603 (N_29603,N_29343,N_29283);
nor U29604 (N_29604,N_29246,N_29110);
nor U29605 (N_29605,N_29139,N_29243);
and U29606 (N_29606,N_29321,N_29152);
or U29607 (N_29607,N_29294,N_29120);
nor U29608 (N_29608,N_29365,N_29237);
xor U29609 (N_29609,N_29148,N_29322);
nand U29610 (N_29610,N_29387,N_29376);
or U29611 (N_29611,N_29224,N_29360);
or U29612 (N_29612,N_29271,N_29263);
or U29613 (N_29613,N_29244,N_29104);
and U29614 (N_29614,N_29312,N_29206);
xor U29615 (N_29615,N_29237,N_29203);
nor U29616 (N_29616,N_29183,N_29107);
or U29617 (N_29617,N_29213,N_29269);
or U29618 (N_29618,N_29174,N_29210);
nand U29619 (N_29619,N_29264,N_29272);
nor U29620 (N_29620,N_29317,N_29144);
nand U29621 (N_29621,N_29219,N_29250);
xor U29622 (N_29622,N_29207,N_29228);
and U29623 (N_29623,N_29104,N_29350);
xor U29624 (N_29624,N_29175,N_29248);
xnor U29625 (N_29625,N_29202,N_29157);
nand U29626 (N_29626,N_29202,N_29331);
and U29627 (N_29627,N_29266,N_29207);
xnor U29628 (N_29628,N_29332,N_29378);
nor U29629 (N_29629,N_29316,N_29363);
xor U29630 (N_29630,N_29185,N_29176);
and U29631 (N_29631,N_29211,N_29207);
and U29632 (N_29632,N_29195,N_29123);
nand U29633 (N_29633,N_29122,N_29325);
or U29634 (N_29634,N_29285,N_29383);
xor U29635 (N_29635,N_29335,N_29312);
xor U29636 (N_29636,N_29296,N_29329);
or U29637 (N_29637,N_29329,N_29295);
or U29638 (N_29638,N_29116,N_29239);
or U29639 (N_29639,N_29161,N_29329);
xor U29640 (N_29640,N_29219,N_29264);
xnor U29641 (N_29641,N_29296,N_29241);
xor U29642 (N_29642,N_29248,N_29194);
or U29643 (N_29643,N_29177,N_29143);
or U29644 (N_29644,N_29248,N_29359);
or U29645 (N_29645,N_29218,N_29202);
nor U29646 (N_29646,N_29395,N_29119);
nand U29647 (N_29647,N_29147,N_29382);
or U29648 (N_29648,N_29372,N_29177);
nor U29649 (N_29649,N_29309,N_29116);
nand U29650 (N_29650,N_29361,N_29298);
nand U29651 (N_29651,N_29203,N_29279);
xnor U29652 (N_29652,N_29241,N_29183);
and U29653 (N_29653,N_29197,N_29273);
nor U29654 (N_29654,N_29163,N_29166);
nand U29655 (N_29655,N_29161,N_29157);
and U29656 (N_29656,N_29359,N_29301);
nand U29657 (N_29657,N_29153,N_29277);
nand U29658 (N_29658,N_29223,N_29351);
and U29659 (N_29659,N_29152,N_29159);
xnor U29660 (N_29660,N_29129,N_29350);
nand U29661 (N_29661,N_29326,N_29253);
xnor U29662 (N_29662,N_29356,N_29365);
xor U29663 (N_29663,N_29150,N_29137);
nor U29664 (N_29664,N_29135,N_29198);
xor U29665 (N_29665,N_29293,N_29272);
and U29666 (N_29666,N_29366,N_29294);
xnor U29667 (N_29667,N_29177,N_29396);
nand U29668 (N_29668,N_29272,N_29311);
or U29669 (N_29669,N_29274,N_29167);
nand U29670 (N_29670,N_29338,N_29217);
and U29671 (N_29671,N_29187,N_29341);
and U29672 (N_29672,N_29304,N_29285);
nor U29673 (N_29673,N_29317,N_29187);
nand U29674 (N_29674,N_29295,N_29279);
nor U29675 (N_29675,N_29373,N_29312);
nor U29676 (N_29676,N_29353,N_29332);
and U29677 (N_29677,N_29300,N_29290);
nor U29678 (N_29678,N_29103,N_29169);
nand U29679 (N_29679,N_29306,N_29103);
nor U29680 (N_29680,N_29192,N_29344);
xor U29681 (N_29681,N_29169,N_29359);
xor U29682 (N_29682,N_29323,N_29310);
or U29683 (N_29683,N_29155,N_29371);
or U29684 (N_29684,N_29179,N_29133);
nor U29685 (N_29685,N_29332,N_29280);
nor U29686 (N_29686,N_29174,N_29374);
or U29687 (N_29687,N_29256,N_29397);
nor U29688 (N_29688,N_29146,N_29298);
nand U29689 (N_29689,N_29240,N_29244);
and U29690 (N_29690,N_29384,N_29377);
nand U29691 (N_29691,N_29293,N_29185);
nor U29692 (N_29692,N_29291,N_29304);
or U29693 (N_29693,N_29126,N_29370);
nor U29694 (N_29694,N_29234,N_29389);
xor U29695 (N_29695,N_29317,N_29326);
nor U29696 (N_29696,N_29304,N_29158);
xnor U29697 (N_29697,N_29107,N_29180);
nor U29698 (N_29698,N_29248,N_29368);
and U29699 (N_29699,N_29307,N_29347);
xnor U29700 (N_29700,N_29600,N_29511);
or U29701 (N_29701,N_29686,N_29625);
nand U29702 (N_29702,N_29678,N_29482);
nand U29703 (N_29703,N_29428,N_29501);
xor U29704 (N_29704,N_29486,N_29659);
xor U29705 (N_29705,N_29635,N_29680);
or U29706 (N_29706,N_29634,N_29427);
xor U29707 (N_29707,N_29568,N_29466);
nor U29708 (N_29708,N_29518,N_29582);
nor U29709 (N_29709,N_29467,N_29690);
or U29710 (N_29710,N_29664,N_29611);
nand U29711 (N_29711,N_29638,N_29505);
or U29712 (N_29712,N_29566,N_29603);
xnor U29713 (N_29713,N_29460,N_29410);
and U29714 (N_29714,N_29683,N_29435);
nand U29715 (N_29715,N_29617,N_29676);
xnor U29716 (N_29716,N_29451,N_29517);
nor U29717 (N_29717,N_29627,N_29503);
nor U29718 (N_29718,N_29510,N_29536);
and U29719 (N_29719,N_29576,N_29624);
and U29720 (N_29720,N_29669,N_29520);
xor U29721 (N_29721,N_29557,N_29577);
xnor U29722 (N_29722,N_29654,N_29637);
or U29723 (N_29723,N_29424,N_29684);
xor U29724 (N_29724,N_29549,N_29475);
nor U29725 (N_29725,N_29695,N_29551);
xor U29726 (N_29726,N_29402,N_29585);
xor U29727 (N_29727,N_29662,N_29552);
nand U29728 (N_29728,N_29494,N_29495);
xnor U29729 (N_29729,N_29693,N_29484);
or U29730 (N_29730,N_29647,N_29496);
xor U29731 (N_29731,N_29499,N_29526);
xnor U29732 (N_29732,N_29458,N_29653);
or U29733 (N_29733,N_29689,N_29614);
nor U29734 (N_29734,N_29504,N_29632);
xnor U29735 (N_29735,N_29480,N_29667);
nor U29736 (N_29736,N_29622,N_29457);
nor U29737 (N_29737,N_29436,N_29623);
or U29738 (N_29738,N_29408,N_29613);
xnor U29739 (N_29739,N_29607,N_29569);
and U29740 (N_29740,N_29497,N_29406);
xnor U29741 (N_29741,N_29485,N_29414);
xor U29742 (N_29742,N_29530,N_29651);
xnor U29743 (N_29743,N_29619,N_29469);
and U29744 (N_29744,N_29409,N_29419);
or U29745 (N_29745,N_29432,N_29620);
or U29746 (N_29746,N_29564,N_29612);
and U29747 (N_29747,N_29610,N_29567);
and U29748 (N_29748,N_29575,N_29593);
and U29749 (N_29749,N_29444,N_29668);
nor U29750 (N_29750,N_29509,N_29465);
and U29751 (N_29751,N_29594,N_29443);
or U29752 (N_29752,N_29642,N_29514);
and U29753 (N_29753,N_29697,N_29578);
xor U29754 (N_29754,N_29649,N_29473);
nor U29755 (N_29755,N_29455,N_29584);
nor U29756 (N_29756,N_29571,N_29452);
nor U29757 (N_29757,N_29687,N_29450);
and U29758 (N_29758,N_29655,N_29645);
nor U29759 (N_29759,N_29660,N_29437);
nor U29760 (N_29760,N_29539,N_29434);
nor U29761 (N_29761,N_29616,N_29556);
xnor U29762 (N_29762,N_29464,N_29438);
xor U29763 (N_29763,N_29646,N_29542);
xnor U29764 (N_29764,N_29404,N_29553);
nor U29765 (N_29765,N_29493,N_29533);
nor U29766 (N_29766,N_29519,N_29629);
or U29767 (N_29767,N_29604,N_29681);
or U29768 (N_29768,N_29691,N_29430);
and U29769 (N_29769,N_29512,N_29574);
nand U29770 (N_29770,N_29546,N_29413);
and U29771 (N_29771,N_29483,N_29601);
nand U29772 (N_29772,N_29538,N_29562);
or U29773 (N_29773,N_29488,N_29698);
nand U29774 (N_29774,N_29440,N_29605);
xnor U29775 (N_29775,N_29657,N_29420);
nor U29776 (N_29776,N_29589,N_29415);
nand U29777 (N_29777,N_29658,N_29547);
or U29778 (N_29778,N_29550,N_29426);
nor U29779 (N_29779,N_29588,N_29537);
or U29780 (N_29780,N_29648,N_29487);
nand U29781 (N_29781,N_29565,N_29447);
or U29782 (N_29782,N_29598,N_29468);
and U29783 (N_29783,N_29679,N_29591);
and U29784 (N_29784,N_29677,N_29532);
nand U29785 (N_29785,N_29491,N_29454);
and U29786 (N_29786,N_29639,N_29543);
and U29787 (N_29787,N_29506,N_29525);
or U29788 (N_29788,N_29489,N_29433);
and U29789 (N_29789,N_29448,N_29685);
nor U29790 (N_29790,N_29661,N_29423);
and U29791 (N_29791,N_29515,N_29560);
or U29792 (N_29792,N_29592,N_29643);
or U29793 (N_29793,N_29596,N_29522);
xnor U29794 (N_29794,N_29570,N_29573);
or U29795 (N_29795,N_29516,N_29682);
and U29796 (N_29796,N_29535,N_29597);
and U29797 (N_29797,N_29507,N_29548);
nor U29798 (N_29798,N_29405,N_29441);
nand U29799 (N_29799,N_29692,N_29595);
nor U29800 (N_29800,N_29583,N_29670);
and U29801 (N_29801,N_29545,N_29498);
nand U29802 (N_29802,N_29492,N_29508);
nand U29803 (N_29803,N_29500,N_29558);
xor U29804 (N_29804,N_29618,N_29666);
and U29805 (N_29805,N_29572,N_29416);
and U29806 (N_29806,N_29644,N_29445);
nor U29807 (N_29807,N_29580,N_29412);
xor U29808 (N_29808,N_29425,N_29431);
nand U29809 (N_29809,N_29609,N_29615);
or U29810 (N_29810,N_29674,N_29534);
xor U29811 (N_29811,N_29688,N_29403);
nand U29812 (N_29812,N_29401,N_29476);
xor U29813 (N_29813,N_29608,N_29665);
and U29814 (N_29814,N_29462,N_29672);
nand U29815 (N_29815,N_29671,N_29590);
nor U29816 (N_29816,N_29587,N_29449);
or U29817 (N_29817,N_29418,N_29477);
and U29818 (N_29818,N_29636,N_29650);
nor U29819 (N_29819,N_29478,N_29581);
or U29820 (N_29820,N_29439,N_29630);
or U29821 (N_29821,N_29579,N_29640);
and U29822 (N_29822,N_29400,N_29699);
or U29823 (N_29823,N_29559,N_29621);
nor U29824 (N_29824,N_29472,N_29694);
xnor U29825 (N_29825,N_29463,N_29554);
nor U29826 (N_29826,N_29474,N_29641);
nor U29827 (N_29827,N_29656,N_29540);
or U29828 (N_29828,N_29555,N_29599);
and U29829 (N_29829,N_29490,N_29631);
nand U29830 (N_29830,N_29529,N_29527);
or U29831 (N_29831,N_29675,N_29456);
nand U29832 (N_29832,N_29446,N_29663);
or U29833 (N_29833,N_29471,N_29470);
nand U29834 (N_29834,N_29502,N_29586);
xnor U29835 (N_29835,N_29633,N_29524);
nand U29836 (N_29836,N_29407,N_29561);
xnor U29837 (N_29837,N_29442,N_29417);
or U29838 (N_29838,N_29544,N_29673);
xor U29839 (N_29839,N_29523,N_29628);
or U29840 (N_29840,N_29606,N_29461);
and U29841 (N_29841,N_29429,N_29602);
xor U29842 (N_29842,N_29652,N_29696);
xor U29843 (N_29843,N_29411,N_29453);
nand U29844 (N_29844,N_29513,N_29563);
nand U29845 (N_29845,N_29528,N_29459);
and U29846 (N_29846,N_29421,N_29521);
xor U29847 (N_29847,N_29531,N_29541);
nor U29848 (N_29848,N_29479,N_29481);
or U29849 (N_29849,N_29626,N_29422);
xnor U29850 (N_29850,N_29421,N_29497);
or U29851 (N_29851,N_29480,N_29555);
and U29852 (N_29852,N_29572,N_29648);
and U29853 (N_29853,N_29533,N_29576);
xor U29854 (N_29854,N_29409,N_29616);
or U29855 (N_29855,N_29420,N_29529);
nand U29856 (N_29856,N_29452,N_29632);
or U29857 (N_29857,N_29467,N_29518);
nand U29858 (N_29858,N_29444,N_29652);
and U29859 (N_29859,N_29692,N_29602);
nand U29860 (N_29860,N_29484,N_29519);
or U29861 (N_29861,N_29677,N_29552);
xnor U29862 (N_29862,N_29504,N_29582);
or U29863 (N_29863,N_29697,N_29436);
nor U29864 (N_29864,N_29639,N_29686);
nor U29865 (N_29865,N_29535,N_29609);
xnor U29866 (N_29866,N_29595,N_29577);
and U29867 (N_29867,N_29520,N_29524);
nor U29868 (N_29868,N_29571,N_29404);
and U29869 (N_29869,N_29478,N_29584);
nand U29870 (N_29870,N_29516,N_29567);
xnor U29871 (N_29871,N_29587,N_29662);
and U29872 (N_29872,N_29657,N_29614);
or U29873 (N_29873,N_29492,N_29431);
nand U29874 (N_29874,N_29659,N_29663);
nor U29875 (N_29875,N_29505,N_29629);
nor U29876 (N_29876,N_29667,N_29645);
nand U29877 (N_29877,N_29548,N_29477);
or U29878 (N_29878,N_29451,N_29612);
and U29879 (N_29879,N_29497,N_29585);
nand U29880 (N_29880,N_29560,N_29453);
xor U29881 (N_29881,N_29500,N_29679);
and U29882 (N_29882,N_29576,N_29480);
and U29883 (N_29883,N_29445,N_29638);
or U29884 (N_29884,N_29645,N_29505);
and U29885 (N_29885,N_29653,N_29549);
nor U29886 (N_29886,N_29637,N_29699);
nand U29887 (N_29887,N_29528,N_29438);
and U29888 (N_29888,N_29606,N_29439);
xnor U29889 (N_29889,N_29464,N_29488);
or U29890 (N_29890,N_29684,N_29463);
xnor U29891 (N_29891,N_29403,N_29460);
nor U29892 (N_29892,N_29566,N_29560);
nand U29893 (N_29893,N_29678,N_29663);
xor U29894 (N_29894,N_29678,N_29695);
nor U29895 (N_29895,N_29482,N_29670);
and U29896 (N_29896,N_29540,N_29454);
nor U29897 (N_29897,N_29600,N_29666);
or U29898 (N_29898,N_29501,N_29510);
nor U29899 (N_29899,N_29504,N_29626);
nor U29900 (N_29900,N_29515,N_29430);
or U29901 (N_29901,N_29616,N_29506);
nand U29902 (N_29902,N_29654,N_29586);
and U29903 (N_29903,N_29635,N_29434);
nor U29904 (N_29904,N_29447,N_29534);
xnor U29905 (N_29905,N_29433,N_29446);
and U29906 (N_29906,N_29536,N_29589);
or U29907 (N_29907,N_29570,N_29692);
and U29908 (N_29908,N_29576,N_29488);
nor U29909 (N_29909,N_29617,N_29625);
nor U29910 (N_29910,N_29628,N_29504);
and U29911 (N_29911,N_29496,N_29598);
and U29912 (N_29912,N_29487,N_29697);
nor U29913 (N_29913,N_29636,N_29562);
or U29914 (N_29914,N_29520,N_29579);
and U29915 (N_29915,N_29539,N_29534);
and U29916 (N_29916,N_29438,N_29419);
nand U29917 (N_29917,N_29690,N_29444);
xnor U29918 (N_29918,N_29540,N_29400);
xor U29919 (N_29919,N_29563,N_29453);
or U29920 (N_29920,N_29636,N_29424);
xnor U29921 (N_29921,N_29670,N_29471);
nand U29922 (N_29922,N_29685,N_29646);
xnor U29923 (N_29923,N_29474,N_29580);
and U29924 (N_29924,N_29609,N_29633);
nand U29925 (N_29925,N_29659,N_29400);
or U29926 (N_29926,N_29680,N_29498);
xor U29927 (N_29927,N_29660,N_29478);
or U29928 (N_29928,N_29494,N_29507);
and U29929 (N_29929,N_29417,N_29558);
xor U29930 (N_29930,N_29549,N_29414);
nor U29931 (N_29931,N_29635,N_29595);
or U29932 (N_29932,N_29623,N_29470);
and U29933 (N_29933,N_29511,N_29403);
and U29934 (N_29934,N_29488,N_29525);
xor U29935 (N_29935,N_29581,N_29425);
and U29936 (N_29936,N_29630,N_29480);
nor U29937 (N_29937,N_29622,N_29535);
or U29938 (N_29938,N_29582,N_29603);
nor U29939 (N_29939,N_29490,N_29625);
and U29940 (N_29940,N_29503,N_29629);
and U29941 (N_29941,N_29643,N_29646);
nor U29942 (N_29942,N_29695,N_29624);
nand U29943 (N_29943,N_29650,N_29619);
nand U29944 (N_29944,N_29515,N_29662);
or U29945 (N_29945,N_29681,N_29533);
nand U29946 (N_29946,N_29451,N_29610);
xnor U29947 (N_29947,N_29581,N_29545);
nor U29948 (N_29948,N_29563,N_29667);
nand U29949 (N_29949,N_29698,N_29466);
or U29950 (N_29950,N_29404,N_29421);
nand U29951 (N_29951,N_29579,N_29646);
nor U29952 (N_29952,N_29427,N_29569);
nand U29953 (N_29953,N_29569,N_29691);
nor U29954 (N_29954,N_29453,N_29413);
or U29955 (N_29955,N_29661,N_29535);
nor U29956 (N_29956,N_29453,N_29468);
nor U29957 (N_29957,N_29549,N_29642);
xor U29958 (N_29958,N_29560,N_29667);
or U29959 (N_29959,N_29682,N_29559);
nand U29960 (N_29960,N_29570,N_29649);
xnor U29961 (N_29961,N_29461,N_29590);
xor U29962 (N_29962,N_29646,N_29680);
and U29963 (N_29963,N_29697,N_29572);
or U29964 (N_29964,N_29674,N_29629);
nor U29965 (N_29965,N_29694,N_29463);
or U29966 (N_29966,N_29478,N_29626);
and U29967 (N_29967,N_29679,N_29529);
or U29968 (N_29968,N_29452,N_29527);
nand U29969 (N_29969,N_29613,N_29568);
or U29970 (N_29970,N_29426,N_29402);
and U29971 (N_29971,N_29474,N_29573);
nor U29972 (N_29972,N_29553,N_29551);
nor U29973 (N_29973,N_29424,N_29503);
xnor U29974 (N_29974,N_29590,N_29523);
or U29975 (N_29975,N_29518,N_29501);
nor U29976 (N_29976,N_29491,N_29618);
and U29977 (N_29977,N_29625,N_29663);
nor U29978 (N_29978,N_29509,N_29489);
or U29979 (N_29979,N_29569,N_29484);
nand U29980 (N_29980,N_29673,N_29676);
nand U29981 (N_29981,N_29416,N_29519);
xnor U29982 (N_29982,N_29520,N_29529);
and U29983 (N_29983,N_29453,N_29573);
nand U29984 (N_29984,N_29502,N_29648);
nand U29985 (N_29985,N_29505,N_29401);
and U29986 (N_29986,N_29544,N_29621);
xnor U29987 (N_29987,N_29408,N_29478);
or U29988 (N_29988,N_29487,N_29519);
nor U29989 (N_29989,N_29448,N_29668);
xnor U29990 (N_29990,N_29636,N_29576);
nand U29991 (N_29991,N_29423,N_29624);
nand U29992 (N_29992,N_29654,N_29666);
xnor U29993 (N_29993,N_29620,N_29438);
and U29994 (N_29994,N_29635,N_29459);
or U29995 (N_29995,N_29412,N_29550);
xor U29996 (N_29996,N_29479,N_29648);
or U29997 (N_29997,N_29685,N_29557);
and U29998 (N_29998,N_29653,N_29627);
or U29999 (N_29999,N_29584,N_29443);
and UO_0 (O_0,N_29994,N_29713);
or UO_1 (O_1,N_29818,N_29938);
xor UO_2 (O_2,N_29944,N_29989);
xnor UO_3 (O_3,N_29720,N_29814);
and UO_4 (O_4,N_29942,N_29785);
and UO_5 (O_5,N_29904,N_29862);
and UO_6 (O_6,N_29748,N_29891);
or UO_7 (O_7,N_29963,N_29867);
xor UO_8 (O_8,N_29722,N_29831);
or UO_9 (O_9,N_29802,N_29875);
nand UO_10 (O_10,N_29728,N_29741);
nor UO_11 (O_11,N_29856,N_29917);
nor UO_12 (O_12,N_29727,N_29845);
xnor UO_13 (O_13,N_29988,N_29721);
nand UO_14 (O_14,N_29954,N_29786);
nand UO_15 (O_15,N_29704,N_29740);
or UO_16 (O_16,N_29842,N_29705);
nand UO_17 (O_17,N_29796,N_29811);
nor UO_18 (O_18,N_29913,N_29799);
or UO_19 (O_19,N_29821,N_29815);
nor UO_20 (O_20,N_29706,N_29798);
or UO_21 (O_21,N_29747,N_29810);
nand UO_22 (O_22,N_29742,N_29813);
nor UO_23 (O_23,N_29829,N_29969);
and UO_24 (O_24,N_29890,N_29937);
xnor UO_25 (O_25,N_29768,N_29964);
or UO_26 (O_26,N_29899,N_29883);
xnor UO_27 (O_27,N_29953,N_29962);
nand UO_28 (O_28,N_29877,N_29724);
xor UO_29 (O_29,N_29718,N_29983);
xor UO_30 (O_30,N_29987,N_29801);
nand UO_31 (O_31,N_29701,N_29966);
xnor UO_32 (O_32,N_29795,N_29971);
nor UO_33 (O_33,N_29751,N_29880);
nand UO_34 (O_34,N_29792,N_29844);
nand UO_35 (O_35,N_29873,N_29896);
or UO_36 (O_36,N_29931,N_29955);
nor UO_37 (O_37,N_29895,N_29929);
nand UO_38 (O_38,N_29783,N_29761);
nor UO_39 (O_39,N_29870,N_29947);
nor UO_40 (O_40,N_29835,N_29833);
nand UO_41 (O_41,N_29847,N_29744);
or UO_42 (O_42,N_29933,N_29843);
and UO_43 (O_43,N_29738,N_29996);
or UO_44 (O_44,N_29789,N_29960);
nor UO_45 (O_45,N_29952,N_29965);
nand UO_46 (O_46,N_29772,N_29733);
nand UO_47 (O_47,N_29916,N_29851);
and UO_48 (O_48,N_29709,N_29788);
xnor UO_49 (O_49,N_29872,N_29758);
nor UO_50 (O_50,N_29806,N_29759);
xor UO_51 (O_51,N_29878,N_29900);
and UO_52 (O_52,N_29812,N_29743);
nand UO_53 (O_53,N_29949,N_29848);
or UO_54 (O_54,N_29749,N_29779);
and UO_55 (O_55,N_29997,N_29825);
and UO_56 (O_56,N_29860,N_29961);
xnor UO_57 (O_57,N_29850,N_29755);
or UO_58 (O_58,N_29750,N_29946);
nand UO_59 (O_59,N_29972,N_29841);
and UO_60 (O_60,N_29708,N_29771);
xnor UO_61 (O_61,N_29995,N_29840);
xnor UO_62 (O_62,N_29817,N_29926);
nand UO_63 (O_63,N_29777,N_29927);
and UO_64 (O_64,N_29975,N_29828);
nor UO_65 (O_65,N_29957,N_29914);
xor UO_66 (O_66,N_29726,N_29716);
and UO_67 (O_67,N_29711,N_29893);
nand UO_68 (O_68,N_29981,N_29808);
nor UO_69 (O_69,N_29864,N_29930);
xor UO_70 (O_70,N_29869,N_29824);
xor UO_71 (O_71,N_29710,N_29924);
xnor UO_72 (O_72,N_29967,N_29909);
nand UO_73 (O_73,N_29919,N_29837);
or UO_74 (O_74,N_29736,N_29876);
nand UO_75 (O_75,N_29910,N_29908);
nor UO_76 (O_76,N_29888,N_29712);
nor UO_77 (O_77,N_29912,N_29948);
and UO_78 (O_78,N_29935,N_29719);
or UO_79 (O_79,N_29700,N_29836);
and UO_80 (O_80,N_29902,N_29868);
nor UO_81 (O_81,N_29846,N_29918);
xnor UO_82 (O_82,N_29739,N_29855);
or UO_83 (O_83,N_29839,N_29977);
nand UO_84 (O_84,N_29781,N_29974);
and UO_85 (O_85,N_29936,N_29764);
nand UO_86 (O_86,N_29999,N_29832);
nand UO_87 (O_87,N_29885,N_29773);
nor UO_88 (O_88,N_29959,N_29854);
and UO_89 (O_89,N_29940,N_29898);
nand UO_90 (O_90,N_29984,N_29730);
nor UO_91 (O_91,N_29906,N_29932);
nor UO_92 (O_92,N_29915,N_29787);
nor UO_93 (O_93,N_29760,N_29853);
nand UO_94 (O_94,N_29993,N_29830);
nor UO_95 (O_95,N_29889,N_29911);
xor UO_96 (O_96,N_29816,N_29901);
xnor UO_97 (O_97,N_29731,N_29746);
or UO_98 (O_98,N_29928,N_29702);
nor UO_99 (O_99,N_29894,N_29881);
and UO_100 (O_100,N_29945,N_29861);
nand UO_101 (O_101,N_29980,N_29852);
nor UO_102 (O_102,N_29715,N_29866);
and UO_103 (O_103,N_29794,N_29897);
nor UO_104 (O_104,N_29859,N_29790);
and UO_105 (O_105,N_29970,N_29703);
or UO_106 (O_106,N_29791,N_29769);
and UO_107 (O_107,N_29725,N_29822);
nand UO_108 (O_108,N_29905,N_29990);
or UO_109 (O_109,N_29784,N_29780);
nor UO_110 (O_110,N_29754,N_29797);
and UO_111 (O_111,N_29734,N_29778);
and UO_112 (O_112,N_29717,N_29732);
nand UO_113 (O_113,N_29770,N_29978);
xnor UO_114 (O_114,N_29737,N_29879);
nor UO_115 (O_115,N_29887,N_29958);
nand UO_116 (O_116,N_29762,N_29968);
nor UO_117 (O_117,N_29776,N_29807);
and UO_118 (O_118,N_29979,N_29809);
xor UO_119 (O_119,N_29823,N_29757);
nand UO_120 (O_120,N_29982,N_29941);
nand UO_121 (O_121,N_29775,N_29849);
nand UO_122 (O_122,N_29745,N_29903);
or UO_123 (O_123,N_29782,N_29943);
or UO_124 (O_124,N_29882,N_29907);
xor UO_125 (O_125,N_29863,N_29986);
nand UO_126 (O_126,N_29729,N_29774);
nand UO_127 (O_127,N_29923,N_29973);
nand UO_128 (O_128,N_29892,N_29874);
nor UO_129 (O_129,N_29921,N_29976);
nand UO_130 (O_130,N_29820,N_29950);
nor UO_131 (O_131,N_29838,N_29991);
or UO_132 (O_132,N_29707,N_29805);
and UO_133 (O_133,N_29992,N_29920);
nor UO_134 (O_134,N_29857,N_29804);
nand UO_135 (O_135,N_29827,N_29956);
xnor UO_136 (O_136,N_29884,N_29752);
or UO_137 (O_137,N_29998,N_29934);
or UO_138 (O_138,N_29763,N_29714);
and UO_139 (O_139,N_29767,N_29886);
or UO_140 (O_140,N_29756,N_29925);
and UO_141 (O_141,N_29922,N_29793);
xnor UO_142 (O_142,N_29753,N_29865);
or UO_143 (O_143,N_29723,N_29951);
nor UO_144 (O_144,N_29765,N_29858);
and UO_145 (O_145,N_29871,N_29766);
or UO_146 (O_146,N_29735,N_29803);
or UO_147 (O_147,N_29800,N_29834);
and UO_148 (O_148,N_29939,N_29826);
nor UO_149 (O_149,N_29985,N_29819);
or UO_150 (O_150,N_29740,N_29932);
nand UO_151 (O_151,N_29816,N_29971);
or UO_152 (O_152,N_29735,N_29824);
nor UO_153 (O_153,N_29756,N_29873);
nor UO_154 (O_154,N_29734,N_29933);
xor UO_155 (O_155,N_29828,N_29704);
nand UO_156 (O_156,N_29945,N_29717);
nor UO_157 (O_157,N_29898,N_29858);
nor UO_158 (O_158,N_29889,N_29737);
nand UO_159 (O_159,N_29898,N_29970);
or UO_160 (O_160,N_29777,N_29901);
nand UO_161 (O_161,N_29919,N_29970);
nand UO_162 (O_162,N_29744,N_29855);
or UO_163 (O_163,N_29765,N_29925);
nor UO_164 (O_164,N_29895,N_29833);
or UO_165 (O_165,N_29888,N_29819);
or UO_166 (O_166,N_29759,N_29799);
and UO_167 (O_167,N_29922,N_29906);
or UO_168 (O_168,N_29884,N_29742);
and UO_169 (O_169,N_29898,N_29831);
nand UO_170 (O_170,N_29926,N_29743);
nor UO_171 (O_171,N_29705,N_29923);
nand UO_172 (O_172,N_29932,N_29726);
nand UO_173 (O_173,N_29858,N_29817);
and UO_174 (O_174,N_29992,N_29965);
xor UO_175 (O_175,N_29721,N_29803);
and UO_176 (O_176,N_29976,N_29847);
nor UO_177 (O_177,N_29717,N_29986);
nor UO_178 (O_178,N_29973,N_29951);
xor UO_179 (O_179,N_29921,N_29993);
nor UO_180 (O_180,N_29989,N_29785);
and UO_181 (O_181,N_29706,N_29826);
nor UO_182 (O_182,N_29895,N_29896);
xnor UO_183 (O_183,N_29734,N_29891);
nand UO_184 (O_184,N_29902,N_29814);
or UO_185 (O_185,N_29775,N_29744);
nor UO_186 (O_186,N_29898,N_29988);
or UO_187 (O_187,N_29876,N_29859);
and UO_188 (O_188,N_29970,N_29945);
or UO_189 (O_189,N_29709,N_29860);
nand UO_190 (O_190,N_29941,N_29757);
nand UO_191 (O_191,N_29863,N_29778);
or UO_192 (O_192,N_29985,N_29737);
nand UO_193 (O_193,N_29968,N_29916);
nor UO_194 (O_194,N_29758,N_29856);
nand UO_195 (O_195,N_29908,N_29855);
nand UO_196 (O_196,N_29763,N_29856);
or UO_197 (O_197,N_29831,N_29838);
xor UO_198 (O_198,N_29925,N_29704);
xor UO_199 (O_199,N_29888,N_29922);
or UO_200 (O_200,N_29811,N_29881);
and UO_201 (O_201,N_29930,N_29951);
nor UO_202 (O_202,N_29980,N_29921);
nor UO_203 (O_203,N_29726,N_29842);
or UO_204 (O_204,N_29822,N_29772);
nand UO_205 (O_205,N_29993,N_29872);
and UO_206 (O_206,N_29787,N_29766);
xor UO_207 (O_207,N_29822,N_29976);
xnor UO_208 (O_208,N_29856,N_29836);
or UO_209 (O_209,N_29795,N_29937);
and UO_210 (O_210,N_29727,N_29742);
nand UO_211 (O_211,N_29904,N_29840);
nand UO_212 (O_212,N_29940,N_29929);
and UO_213 (O_213,N_29831,N_29767);
nand UO_214 (O_214,N_29745,N_29840);
or UO_215 (O_215,N_29990,N_29724);
xor UO_216 (O_216,N_29871,N_29884);
and UO_217 (O_217,N_29929,N_29848);
nand UO_218 (O_218,N_29725,N_29736);
nand UO_219 (O_219,N_29832,N_29888);
and UO_220 (O_220,N_29747,N_29927);
or UO_221 (O_221,N_29700,N_29831);
or UO_222 (O_222,N_29872,N_29998);
nor UO_223 (O_223,N_29920,N_29738);
or UO_224 (O_224,N_29803,N_29772);
nor UO_225 (O_225,N_29810,N_29748);
nand UO_226 (O_226,N_29752,N_29859);
nand UO_227 (O_227,N_29789,N_29749);
and UO_228 (O_228,N_29816,N_29942);
xor UO_229 (O_229,N_29869,N_29907);
nor UO_230 (O_230,N_29865,N_29708);
and UO_231 (O_231,N_29829,N_29997);
xor UO_232 (O_232,N_29734,N_29879);
nor UO_233 (O_233,N_29807,N_29830);
or UO_234 (O_234,N_29871,N_29867);
xnor UO_235 (O_235,N_29796,N_29908);
nand UO_236 (O_236,N_29829,N_29891);
nand UO_237 (O_237,N_29740,N_29822);
nand UO_238 (O_238,N_29927,N_29700);
or UO_239 (O_239,N_29770,N_29783);
nor UO_240 (O_240,N_29714,N_29740);
or UO_241 (O_241,N_29842,N_29984);
or UO_242 (O_242,N_29883,N_29826);
nand UO_243 (O_243,N_29742,N_29700);
or UO_244 (O_244,N_29721,N_29779);
and UO_245 (O_245,N_29735,N_29850);
xnor UO_246 (O_246,N_29795,N_29891);
xor UO_247 (O_247,N_29724,N_29927);
nand UO_248 (O_248,N_29715,N_29979);
xnor UO_249 (O_249,N_29901,N_29791);
nor UO_250 (O_250,N_29888,N_29769);
nand UO_251 (O_251,N_29792,N_29708);
or UO_252 (O_252,N_29874,N_29751);
nand UO_253 (O_253,N_29887,N_29869);
nor UO_254 (O_254,N_29935,N_29906);
xnor UO_255 (O_255,N_29732,N_29734);
and UO_256 (O_256,N_29751,N_29716);
nor UO_257 (O_257,N_29959,N_29749);
or UO_258 (O_258,N_29846,N_29882);
nor UO_259 (O_259,N_29925,N_29742);
xnor UO_260 (O_260,N_29970,N_29894);
nand UO_261 (O_261,N_29768,N_29729);
nor UO_262 (O_262,N_29823,N_29782);
and UO_263 (O_263,N_29818,N_29987);
nor UO_264 (O_264,N_29906,N_29875);
and UO_265 (O_265,N_29941,N_29976);
nand UO_266 (O_266,N_29974,N_29813);
nand UO_267 (O_267,N_29953,N_29871);
or UO_268 (O_268,N_29804,N_29839);
nand UO_269 (O_269,N_29700,N_29705);
xor UO_270 (O_270,N_29803,N_29773);
xnor UO_271 (O_271,N_29860,N_29778);
or UO_272 (O_272,N_29783,N_29763);
nand UO_273 (O_273,N_29718,N_29767);
nand UO_274 (O_274,N_29724,N_29827);
or UO_275 (O_275,N_29758,N_29893);
nand UO_276 (O_276,N_29993,N_29739);
xnor UO_277 (O_277,N_29941,N_29927);
or UO_278 (O_278,N_29783,N_29933);
nand UO_279 (O_279,N_29945,N_29768);
xor UO_280 (O_280,N_29911,N_29960);
or UO_281 (O_281,N_29856,N_29897);
xor UO_282 (O_282,N_29853,N_29791);
and UO_283 (O_283,N_29851,N_29830);
nand UO_284 (O_284,N_29894,N_29707);
and UO_285 (O_285,N_29877,N_29764);
or UO_286 (O_286,N_29991,N_29932);
xor UO_287 (O_287,N_29929,N_29765);
and UO_288 (O_288,N_29837,N_29854);
or UO_289 (O_289,N_29847,N_29989);
nand UO_290 (O_290,N_29814,N_29950);
nand UO_291 (O_291,N_29963,N_29844);
nor UO_292 (O_292,N_29946,N_29812);
or UO_293 (O_293,N_29882,N_29771);
or UO_294 (O_294,N_29943,N_29794);
nor UO_295 (O_295,N_29929,N_29867);
and UO_296 (O_296,N_29866,N_29703);
nand UO_297 (O_297,N_29847,N_29772);
and UO_298 (O_298,N_29805,N_29944);
nor UO_299 (O_299,N_29937,N_29705);
nand UO_300 (O_300,N_29998,N_29983);
and UO_301 (O_301,N_29918,N_29858);
xor UO_302 (O_302,N_29948,N_29851);
nor UO_303 (O_303,N_29773,N_29960);
or UO_304 (O_304,N_29834,N_29975);
xnor UO_305 (O_305,N_29832,N_29836);
xnor UO_306 (O_306,N_29951,N_29986);
nand UO_307 (O_307,N_29999,N_29803);
xnor UO_308 (O_308,N_29905,N_29999);
and UO_309 (O_309,N_29815,N_29887);
nor UO_310 (O_310,N_29715,N_29743);
or UO_311 (O_311,N_29961,N_29889);
xor UO_312 (O_312,N_29783,N_29704);
or UO_313 (O_313,N_29810,N_29811);
nor UO_314 (O_314,N_29991,N_29891);
nand UO_315 (O_315,N_29787,N_29867);
xnor UO_316 (O_316,N_29729,N_29728);
xor UO_317 (O_317,N_29910,N_29787);
nor UO_318 (O_318,N_29935,N_29916);
nor UO_319 (O_319,N_29998,N_29942);
nand UO_320 (O_320,N_29710,N_29892);
nor UO_321 (O_321,N_29962,N_29803);
or UO_322 (O_322,N_29944,N_29810);
nand UO_323 (O_323,N_29866,N_29863);
and UO_324 (O_324,N_29955,N_29759);
or UO_325 (O_325,N_29919,N_29998);
nor UO_326 (O_326,N_29860,N_29736);
or UO_327 (O_327,N_29796,N_29973);
or UO_328 (O_328,N_29910,N_29994);
nand UO_329 (O_329,N_29735,N_29952);
and UO_330 (O_330,N_29912,N_29724);
or UO_331 (O_331,N_29721,N_29990);
nor UO_332 (O_332,N_29993,N_29746);
or UO_333 (O_333,N_29956,N_29707);
nand UO_334 (O_334,N_29743,N_29947);
nor UO_335 (O_335,N_29753,N_29987);
nor UO_336 (O_336,N_29716,N_29761);
or UO_337 (O_337,N_29898,N_29960);
or UO_338 (O_338,N_29799,N_29854);
nor UO_339 (O_339,N_29961,N_29890);
nand UO_340 (O_340,N_29762,N_29800);
or UO_341 (O_341,N_29916,N_29909);
nor UO_342 (O_342,N_29927,N_29996);
nor UO_343 (O_343,N_29942,N_29813);
or UO_344 (O_344,N_29870,N_29920);
nand UO_345 (O_345,N_29968,N_29796);
nor UO_346 (O_346,N_29851,N_29710);
or UO_347 (O_347,N_29724,N_29991);
nand UO_348 (O_348,N_29839,N_29882);
or UO_349 (O_349,N_29937,N_29810);
or UO_350 (O_350,N_29975,N_29791);
or UO_351 (O_351,N_29715,N_29885);
xnor UO_352 (O_352,N_29938,N_29796);
or UO_353 (O_353,N_29911,N_29935);
nand UO_354 (O_354,N_29868,N_29762);
nor UO_355 (O_355,N_29758,N_29701);
and UO_356 (O_356,N_29916,N_29960);
xnor UO_357 (O_357,N_29870,N_29961);
xor UO_358 (O_358,N_29888,N_29887);
xor UO_359 (O_359,N_29871,N_29707);
and UO_360 (O_360,N_29843,N_29936);
nand UO_361 (O_361,N_29859,N_29845);
or UO_362 (O_362,N_29917,N_29951);
nand UO_363 (O_363,N_29862,N_29819);
nand UO_364 (O_364,N_29919,N_29757);
xnor UO_365 (O_365,N_29775,N_29734);
nand UO_366 (O_366,N_29999,N_29838);
and UO_367 (O_367,N_29965,N_29774);
xor UO_368 (O_368,N_29948,N_29703);
nor UO_369 (O_369,N_29830,N_29857);
nor UO_370 (O_370,N_29999,N_29783);
xor UO_371 (O_371,N_29702,N_29878);
or UO_372 (O_372,N_29711,N_29736);
nand UO_373 (O_373,N_29826,N_29728);
nand UO_374 (O_374,N_29778,N_29995);
or UO_375 (O_375,N_29993,N_29960);
or UO_376 (O_376,N_29845,N_29952);
nor UO_377 (O_377,N_29715,N_29837);
nor UO_378 (O_378,N_29711,N_29753);
xnor UO_379 (O_379,N_29991,N_29822);
xnor UO_380 (O_380,N_29757,N_29884);
nor UO_381 (O_381,N_29809,N_29769);
nor UO_382 (O_382,N_29929,N_29746);
or UO_383 (O_383,N_29899,N_29812);
nand UO_384 (O_384,N_29768,N_29887);
or UO_385 (O_385,N_29848,N_29702);
nor UO_386 (O_386,N_29715,N_29731);
xor UO_387 (O_387,N_29721,N_29759);
nand UO_388 (O_388,N_29709,N_29814);
or UO_389 (O_389,N_29723,N_29877);
and UO_390 (O_390,N_29892,N_29915);
and UO_391 (O_391,N_29992,N_29751);
and UO_392 (O_392,N_29756,N_29705);
nand UO_393 (O_393,N_29782,N_29785);
nor UO_394 (O_394,N_29762,N_29908);
nand UO_395 (O_395,N_29741,N_29856);
nor UO_396 (O_396,N_29717,N_29991);
xor UO_397 (O_397,N_29901,N_29936);
and UO_398 (O_398,N_29707,N_29952);
xor UO_399 (O_399,N_29735,N_29949);
nand UO_400 (O_400,N_29906,N_29736);
or UO_401 (O_401,N_29966,N_29837);
or UO_402 (O_402,N_29802,N_29795);
xor UO_403 (O_403,N_29816,N_29958);
and UO_404 (O_404,N_29871,N_29910);
and UO_405 (O_405,N_29835,N_29925);
and UO_406 (O_406,N_29925,N_29845);
and UO_407 (O_407,N_29895,N_29813);
and UO_408 (O_408,N_29782,N_29985);
xnor UO_409 (O_409,N_29778,N_29735);
nor UO_410 (O_410,N_29985,N_29998);
nand UO_411 (O_411,N_29966,N_29770);
nand UO_412 (O_412,N_29995,N_29753);
nor UO_413 (O_413,N_29968,N_29748);
nand UO_414 (O_414,N_29828,N_29918);
and UO_415 (O_415,N_29884,N_29828);
xor UO_416 (O_416,N_29826,N_29736);
nor UO_417 (O_417,N_29914,N_29723);
or UO_418 (O_418,N_29988,N_29834);
and UO_419 (O_419,N_29962,N_29892);
nor UO_420 (O_420,N_29881,N_29931);
and UO_421 (O_421,N_29716,N_29972);
xor UO_422 (O_422,N_29918,N_29766);
nor UO_423 (O_423,N_29722,N_29732);
or UO_424 (O_424,N_29775,N_29840);
and UO_425 (O_425,N_29886,N_29812);
nor UO_426 (O_426,N_29751,N_29899);
xor UO_427 (O_427,N_29850,N_29776);
and UO_428 (O_428,N_29715,N_29777);
or UO_429 (O_429,N_29751,N_29805);
xnor UO_430 (O_430,N_29819,N_29920);
or UO_431 (O_431,N_29806,N_29898);
or UO_432 (O_432,N_29722,N_29734);
or UO_433 (O_433,N_29774,N_29824);
nand UO_434 (O_434,N_29805,N_29997);
nand UO_435 (O_435,N_29932,N_29822);
nor UO_436 (O_436,N_29797,N_29744);
or UO_437 (O_437,N_29719,N_29928);
or UO_438 (O_438,N_29745,N_29935);
and UO_439 (O_439,N_29903,N_29841);
xor UO_440 (O_440,N_29835,N_29736);
and UO_441 (O_441,N_29749,N_29989);
xnor UO_442 (O_442,N_29928,N_29948);
nand UO_443 (O_443,N_29896,N_29768);
or UO_444 (O_444,N_29923,N_29948);
or UO_445 (O_445,N_29869,N_29863);
or UO_446 (O_446,N_29793,N_29831);
xnor UO_447 (O_447,N_29964,N_29720);
nand UO_448 (O_448,N_29779,N_29846);
xnor UO_449 (O_449,N_29870,N_29992);
nor UO_450 (O_450,N_29855,N_29793);
xnor UO_451 (O_451,N_29730,N_29924);
nor UO_452 (O_452,N_29936,N_29965);
and UO_453 (O_453,N_29860,N_29914);
nand UO_454 (O_454,N_29721,N_29702);
nor UO_455 (O_455,N_29717,N_29721);
xnor UO_456 (O_456,N_29800,N_29946);
and UO_457 (O_457,N_29967,N_29900);
and UO_458 (O_458,N_29909,N_29846);
nand UO_459 (O_459,N_29778,N_29979);
xnor UO_460 (O_460,N_29710,N_29805);
or UO_461 (O_461,N_29759,N_29957);
xnor UO_462 (O_462,N_29962,N_29734);
nand UO_463 (O_463,N_29882,N_29989);
nor UO_464 (O_464,N_29934,N_29831);
or UO_465 (O_465,N_29846,N_29905);
xor UO_466 (O_466,N_29810,N_29946);
nand UO_467 (O_467,N_29890,N_29944);
nor UO_468 (O_468,N_29879,N_29743);
and UO_469 (O_469,N_29738,N_29782);
or UO_470 (O_470,N_29780,N_29745);
and UO_471 (O_471,N_29955,N_29817);
xor UO_472 (O_472,N_29845,N_29804);
and UO_473 (O_473,N_29915,N_29757);
and UO_474 (O_474,N_29810,N_29870);
nand UO_475 (O_475,N_29856,N_29870);
and UO_476 (O_476,N_29903,N_29898);
xor UO_477 (O_477,N_29824,N_29844);
nand UO_478 (O_478,N_29725,N_29949);
nand UO_479 (O_479,N_29943,N_29770);
nor UO_480 (O_480,N_29827,N_29779);
and UO_481 (O_481,N_29991,N_29825);
nand UO_482 (O_482,N_29954,N_29899);
and UO_483 (O_483,N_29755,N_29872);
or UO_484 (O_484,N_29778,N_29994);
xnor UO_485 (O_485,N_29811,N_29725);
nand UO_486 (O_486,N_29786,N_29773);
nand UO_487 (O_487,N_29909,N_29969);
xnor UO_488 (O_488,N_29845,N_29700);
or UO_489 (O_489,N_29713,N_29963);
and UO_490 (O_490,N_29841,N_29937);
xor UO_491 (O_491,N_29829,N_29856);
or UO_492 (O_492,N_29725,N_29857);
or UO_493 (O_493,N_29906,N_29705);
and UO_494 (O_494,N_29864,N_29789);
or UO_495 (O_495,N_29841,N_29794);
xnor UO_496 (O_496,N_29727,N_29825);
and UO_497 (O_497,N_29841,N_29959);
nand UO_498 (O_498,N_29811,N_29736);
and UO_499 (O_499,N_29744,N_29848);
xnor UO_500 (O_500,N_29871,N_29727);
or UO_501 (O_501,N_29930,N_29767);
xor UO_502 (O_502,N_29973,N_29972);
nor UO_503 (O_503,N_29972,N_29987);
and UO_504 (O_504,N_29985,N_29786);
or UO_505 (O_505,N_29705,N_29874);
xor UO_506 (O_506,N_29822,N_29947);
xnor UO_507 (O_507,N_29969,N_29937);
nor UO_508 (O_508,N_29853,N_29866);
and UO_509 (O_509,N_29739,N_29895);
nand UO_510 (O_510,N_29963,N_29993);
or UO_511 (O_511,N_29721,N_29701);
or UO_512 (O_512,N_29742,N_29912);
nand UO_513 (O_513,N_29969,N_29852);
xnor UO_514 (O_514,N_29999,N_29771);
xor UO_515 (O_515,N_29925,N_29785);
or UO_516 (O_516,N_29701,N_29834);
nand UO_517 (O_517,N_29894,N_29932);
nor UO_518 (O_518,N_29848,N_29880);
xnor UO_519 (O_519,N_29787,N_29776);
nor UO_520 (O_520,N_29844,N_29839);
xnor UO_521 (O_521,N_29956,N_29703);
nand UO_522 (O_522,N_29840,N_29900);
nor UO_523 (O_523,N_29818,N_29931);
xor UO_524 (O_524,N_29800,N_29813);
xor UO_525 (O_525,N_29979,N_29806);
nand UO_526 (O_526,N_29916,N_29952);
and UO_527 (O_527,N_29811,N_29938);
xor UO_528 (O_528,N_29886,N_29797);
nor UO_529 (O_529,N_29941,N_29953);
nand UO_530 (O_530,N_29797,N_29840);
xor UO_531 (O_531,N_29917,N_29766);
or UO_532 (O_532,N_29903,N_29761);
nor UO_533 (O_533,N_29975,N_29718);
nor UO_534 (O_534,N_29723,N_29766);
and UO_535 (O_535,N_29887,N_29965);
and UO_536 (O_536,N_29891,N_29868);
xnor UO_537 (O_537,N_29859,N_29985);
nand UO_538 (O_538,N_29773,N_29976);
nor UO_539 (O_539,N_29948,N_29987);
nand UO_540 (O_540,N_29791,N_29704);
or UO_541 (O_541,N_29760,N_29732);
nand UO_542 (O_542,N_29876,N_29998);
or UO_543 (O_543,N_29837,N_29812);
xor UO_544 (O_544,N_29831,N_29816);
or UO_545 (O_545,N_29701,N_29840);
and UO_546 (O_546,N_29930,N_29725);
or UO_547 (O_547,N_29770,N_29805);
nand UO_548 (O_548,N_29914,N_29782);
nand UO_549 (O_549,N_29722,N_29769);
nor UO_550 (O_550,N_29916,N_29702);
and UO_551 (O_551,N_29861,N_29718);
nor UO_552 (O_552,N_29957,N_29911);
and UO_553 (O_553,N_29734,N_29744);
and UO_554 (O_554,N_29905,N_29813);
xnor UO_555 (O_555,N_29785,N_29914);
nor UO_556 (O_556,N_29880,N_29799);
nor UO_557 (O_557,N_29993,N_29977);
or UO_558 (O_558,N_29730,N_29942);
and UO_559 (O_559,N_29749,N_29914);
xor UO_560 (O_560,N_29946,N_29738);
nand UO_561 (O_561,N_29851,N_29725);
xnor UO_562 (O_562,N_29724,N_29804);
nor UO_563 (O_563,N_29784,N_29949);
and UO_564 (O_564,N_29957,N_29790);
nor UO_565 (O_565,N_29767,N_29837);
nor UO_566 (O_566,N_29731,N_29805);
xnor UO_567 (O_567,N_29712,N_29764);
or UO_568 (O_568,N_29800,N_29801);
xor UO_569 (O_569,N_29758,N_29889);
nor UO_570 (O_570,N_29740,N_29833);
or UO_571 (O_571,N_29957,N_29767);
and UO_572 (O_572,N_29758,N_29987);
and UO_573 (O_573,N_29710,N_29976);
nor UO_574 (O_574,N_29923,N_29922);
and UO_575 (O_575,N_29971,N_29861);
nand UO_576 (O_576,N_29982,N_29780);
xnor UO_577 (O_577,N_29852,N_29789);
xor UO_578 (O_578,N_29857,N_29721);
or UO_579 (O_579,N_29893,N_29960);
nor UO_580 (O_580,N_29973,N_29865);
nand UO_581 (O_581,N_29810,N_29749);
nand UO_582 (O_582,N_29756,N_29968);
and UO_583 (O_583,N_29961,N_29906);
and UO_584 (O_584,N_29877,N_29848);
xnor UO_585 (O_585,N_29965,N_29733);
nor UO_586 (O_586,N_29996,N_29895);
and UO_587 (O_587,N_29882,N_29920);
or UO_588 (O_588,N_29847,N_29927);
nand UO_589 (O_589,N_29762,N_29969);
or UO_590 (O_590,N_29751,N_29831);
nor UO_591 (O_591,N_29703,N_29833);
and UO_592 (O_592,N_29942,N_29721);
or UO_593 (O_593,N_29854,N_29943);
and UO_594 (O_594,N_29930,N_29738);
nand UO_595 (O_595,N_29793,N_29977);
nor UO_596 (O_596,N_29922,N_29790);
or UO_597 (O_597,N_29828,N_29994);
nor UO_598 (O_598,N_29943,N_29994);
nand UO_599 (O_599,N_29887,N_29909);
nor UO_600 (O_600,N_29791,N_29839);
xnor UO_601 (O_601,N_29716,N_29940);
nand UO_602 (O_602,N_29770,N_29922);
xor UO_603 (O_603,N_29979,N_29713);
or UO_604 (O_604,N_29860,N_29965);
or UO_605 (O_605,N_29948,N_29765);
and UO_606 (O_606,N_29820,N_29702);
nor UO_607 (O_607,N_29704,N_29920);
xor UO_608 (O_608,N_29836,N_29737);
nor UO_609 (O_609,N_29759,N_29867);
nor UO_610 (O_610,N_29828,N_29999);
xnor UO_611 (O_611,N_29997,N_29866);
or UO_612 (O_612,N_29729,N_29758);
nand UO_613 (O_613,N_29996,N_29828);
xor UO_614 (O_614,N_29784,N_29861);
xor UO_615 (O_615,N_29761,N_29908);
and UO_616 (O_616,N_29831,N_29901);
and UO_617 (O_617,N_29830,N_29913);
and UO_618 (O_618,N_29922,N_29904);
xor UO_619 (O_619,N_29957,N_29908);
and UO_620 (O_620,N_29721,N_29907);
or UO_621 (O_621,N_29948,N_29746);
nand UO_622 (O_622,N_29972,N_29860);
xor UO_623 (O_623,N_29999,N_29958);
nor UO_624 (O_624,N_29823,N_29960);
xor UO_625 (O_625,N_29708,N_29849);
xnor UO_626 (O_626,N_29822,N_29856);
xor UO_627 (O_627,N_29823,N_29809);
and UO_628 (O_628,N_29981,N_29824);
nand UO_629 (O_629,N_29809,N_29735);
nand UO_630 (O_630,N_29980,N_29969);
or UO_631 (O_631,N_29710,N_29848);
xnor UO_632 (O_632,N_29944,N_29716);
or UO_633 (O_633,N_29878,N_29713);
or UO_634 (O_634,N_29739,N_29880);
nor UO_635 (O_635,N_29781,N_29953);
or UO_636 (O_636,N_29762,N_29839);
and UO_637 (O_637,N_29734,N_29749);
nor UO_638 (O_638,N_29710,N_29883);
and UO_639 (O_639,N_29887,N_29825);
and UO_640 (O_640,N_29700,N_29731);
or UO_641 (O_641,N_29894,N_29964);
and UO_642 (O_642,N_29917,N_29978);
and UO_643 (O_643,N_29722,N_29948);
xnor UO_644 (O_644,N_29815,N_29891);
nand UO_645 (O_645,N_29830,N_29972);
and UO_646 (O_646,N_29980,N_29958);
xnor UO_647 (O_647,N_29839,N_29780);
xor UO_648 (O_648,N_29770,N_29931);
nor UO_649 (O_649,N_29899,N_29750);
xor UO_650 (O_650,N_29936,N_29983);
xor UO_651 (O_651,N_29734,N_29737);
nand UO_652 (O_652,N_29817,N_29913);
nand UO_653 (O_653,N_29710,N_29914);
xor UO_654 (O_654,N_29876,N_29878);
xor UO_655 (O_655,N_29928,N_29925);
xor UO_656 (O_656,N_29908,N_29921);
and UO_657 (O_657,N_29797,N_29936);
nand UO_658 (O_658,N_29713,N_29737);
nor UO_659 (O_659,N_29839,N_29773);
and UO_660 (O_660,N_29739,N_29784);
xor UO_661 (O_661,N_29831,N_29795);
or UO_662 (O_662,N_29728,N_29713);
nor UO_663 (O_663,N_29706,N_29795);
xnor UO_664 (O_664,N_29885,N_29844);
or UO_665 (O_665,N_29820,N_29794);
xnor UO_666 (O_666,N_29981,N_29762);
or UO_667 (O_667,N_29990,N_29973);
or UO_668 (O_668,N_29813,N_29793);
and UO_669 (O_669,N_29852,N_29963);
nand UO_670 (O_670,N_29817,N_29813);
nor UO_671 (O_671,N_29985,N_29979);
and UO_672 (O_672,N_29869,N_29882);
and UO_673 (O_673,N_29983,N_29761);
and UO_674 (O_674,N_29916,N_29752);
or UO_675 (O_675,N_29799,N_29999);
xnor UO_676 (O_676,N_29836,N_29701);
and UO_677 (O_677,N_29869,N_29879);
or UO_678 (O_678,N_29793,N_29723);
xor UO_679 (O_679,N_29908,N_29715);
and UO_680 (O_680,N_29903,N_29721);
xor UO_681 (O_681,N_29906,N_29848);
xor UO_682 (O_682,N_29758,N_29750);
nand UO_683 (O_683,N_29809,N_29779);
nand UO_684 (O_684,N_29908,N_29830);
nand UO_685 (O_685,N_29792,N_29776);
xor UO_686 (O_686,N_29955,N_29719);
xnor UO_687 (O_687,N_29930,N_29941);
or UO_688 (O_688,N_29817,N_29921);
or UO_689 (O_689,N_29744,N_29920);
and UO_690 (O_690,N_29864,N_29950);
or UO_691 (O_691,N_29834,N_29810);
xor UO_692 (O_692,N_29805,N_29861);
xor UO_693 (O_693,N_29914,N_29726);
nand UO_694 (O_694,N_29939,N_29902);
and UO_695 (O_695,N_29895,N_29733);
xnor UO_696 (O_696,N_29997,N_29838);
nor UO_697 (O_697,N_29950,N_29746);
nor UO_698 (O_698,N_29793,N_29715);
nand UO_699 (O_699,N_29825,N_29724);
nor UO_700 (O_700,N_29837,N_29766);
or UO_701 (O_701,N_29874,N_29993);
xor UO_702 (O_702,N_29962,N_29918);
nor UO_703 (O_703,N_29716,N_29779);
xor UO_704 (O_704,N_29829,N_29983);
nand UO_705 (O_705,N_29738,N_29860);
xnor UO_706 (O_706,N_29828,N_29886);
nor UO_707 (O_707,N_29856,N_29710);
nor UO_708 (O_708,N_29996,N_29854);
or UO_709 (O_709,N_29981,N_29742);
nand UO_710 (O_710,N_29922,N_29868);
nor UO_711 (O_711,N_29803,N_29924);
and UO_712 (O_712,N_29990,N_29725);
or UO_713 (O_713,N_29966,N_29707);
nor UO_714 (O_714,N_29706,N_29830);
nand UO_715 (O_715,N_29703,N_29836);
or UO_716 (O_716,N_29861,N_29992);
xnor UO_717 (O_717,N_29829,N_29801);
or UO_718 (O_718,N_29855,N_29715);
nand UO_719 (O_719,N_29940,N_29759);
xnor UO_720 (O_720,N_29897,N_29919);
nand UO_721 (O_721,N_29830,N_29914);
xnor UO_722 (O_722,N_29981,N_29720);
nand UO_723 (O_723,N_29753,N_29930);
nor UO_724 (O_724,N_29933,N_29703);
nor UO_725 (O_725,N_29926,N_29915);
nand UO_726 (O_726,N_29770,N_29955);
nand UO_727 (O_727,N_29732,N_29968);
or UO_728 (O_728,N_29760,N_29828);
or UO_729 (O_729,N_29781,N_29752);
nand UO_730 (O_730,N_29991,N_29755);
or UO_731 (O_731,N_29780,N_29820);
nor UO_732 (O_732,N_29805,N_29949);
nor UO_733 (O_733,N_29843,N_29785);
nor UO_734 (O_734,N_29996,N_29959);
xor UO_735 (O_735,N_29854,N_29902);
xor UO_736 (O_736,N_29775,N_29890);
xor UO_737 (O_737,N_29704,N_29883);
and UO_738 (O_738,N_29884,N_29803);
nor UO_739 (O_739,N_29829,N_29787);
or UO_740 (O_740,N_29993,N_29770);
xor UO_741 (O_741,N_29871,N_29713);
or UO_742 (O_742,N_29899,N_29895);
and UO_743 (O_743,N_29988,N_29860);
or UO_744 (O_744,N_29714,N_29873);
or UO_745 (O_745,N_29897,N_29741);
nor UO_746 (O_746,N_29999,N_29752);
nor UO_747 (O_747,N_29979,N_29899);
and UO_748 (O_748,N_29908,N_29818);
and UO_749 (O_749,N_29722,N_29938);
xor UO_750 (O_750,N_29726,N_29869);
xor UO_751 (O_751,N_29922,N_29794);
nor UO_752 (O_752,N_29898,N_29771);
or UO_753 (O_753,N_29970,N_29720);
and UO_754 (O_754,N_29807,N_29786);
and UO_755 (O_755,N_29787,N_29778);
nor UO_756 (O_756,N_29880,N_29864);
xnor UO_757 (O_757,N_29897,N_29716);
or UO_758 (O_758,N_29889,N_29844);
nand UO_759 (O_759,N_29938,N_29729);
xnor UO_760 (O_760,N_29733,N_29859);
nor UO_761 (O_761,N_29787,N_29855);
nand UO_762 (O_762,N_29814,N_29997);
or UO_763 (O_763,N_29991,N_29741);
or UO_764 (O_764,N_29788,N_29956);
nand UO_765 (O_765,N_29821,N_29768);
nand UO_766 (O_766,N_29862,N_29977);
nand UO_767 (O_767,N_29852,N_29939);
or UO_768 (O_768,N_29778,N_29943);
and UO_769 (O_769,N_29754,N_29876);
xnor UO_770 (O_770,N_29858,N_29795);
nand UO_771 (O_771,N_29708,N_29782);
nor UO_772 (O_772,N_29824,N_29739);
and UO_773 (O_773,N_29847,N_29889);
nor UO_774 (O_774,N_29704,N_29745);
nor UO_775 (O_775,N_29733,N_29728);
nor UO_776 (O_776,N_29745,N_29918);
or UO_777 (O_777,N_29926,N_29884);
or UO_778 (O_778,N_29984,N_29711);
or UO_779 (O_779,N_29968,N_29884);
xor UO_780 (O_780,N_29864,N_29839);
or UO_781 (O_781,N_29744,N_29743);
and UO_782 (O_782,N_29912,N_29879);
xnor UO_783 (O_783,N_29763,N_29864);
nand UO_784 (O_784,N_29759,N_29925);
nand UO_785 (O_785,N_29821,N_29851);
nand UO_786 (O_786,N_29930,N_29815);
and UO_787 (O_787,N_29935,N_29890);
or UO_788 (O_788,N_29845,N_29877);
xnor UO_789 (O_789,N_29754,N_29712);
or UO_790 (O_790,N_29797,N_29774);
nor UO_791 (O_791,N_29902,N_29866);
nand UO_792 (O_792,N_29924,N_29866);
and UO_793 (O_793,N_29993,N_29905);
and UO_794 (O_794,N_29919,N_29907);
or UO_795 (O_795,N_29952,N_29984);
xor UO_796 (O_796,N_29868,N_29831);
nand UO_797 (O_797,N_29903,N_29893);
and UO_798 (O_798,N_29742,N_29809);
xor UO_799 (O_799,N_29723,N_29929);
and UO_800 (O_800,N_29777,N_29760);
or UO_801 (O_801,N_29947,N_29786);
nand UO_802 (O_802,N_29815,N_29702);
nand UO_803 (O_803,N_29994,N_29992);
nor UO_804 (O_804,N_29731,N_29873);
nand UO_805 (O_805,N_29856,N_29898);
xor UO_806 (O_806,N_29772,N_29843);
nor UO_807 (O_807,N_29870,N_29929);
nor UO_808 (O_808,N_29827,N_29748);
nor UO_809 (O_809,N_29833,N_29813);
nand UO_810 (O_810,N_29854,N_29921);
xor UO_811 (O_811,N_29765,N_29957);
xor UO_812 (O_812,N_29829,N_29770);
nand UO_813 (O_813,N_29808,N_29740);
nor UO_814 (O_814,N_29874,N_29960);
nand UO_815 (O_815,N_29891,N_29823);
nor UO_816 (O_816,N_29854,N_29896);
xnor UO_817 (O_817,N_29818,N_29786);
nor UO_818 (O_818,N_29825,N_29780);
nand UO_819 (O_819,N_29921,N_29996);
nor UO_820 (O_820,N_29776,N_29966);
and UO_821 (O_821,N_29855,N_29920);
nand UO_822 (O_822,N_29861,N_29779);
or UO_823 (O_823,N_29998,N_29993);
nand UO_824 (O_824,N_29822,N_29866);
xor UO_825 (O_825,N_29946,N_29910);
nor UO_826 (O_826,N_29986,N_29875);
or UO_827 (O_827,N_29858,N_29867);
nor UO_828 (O_828,N_29835,N_29942);
nand UO_829 (O_829,N_29837,N_29969);
nor UO_830 (O_830,N_29779,N_29892);
xor UO_831 (O_831,N_29791,N_29899);
and UO_832 (O_832,N_29912,N_29927);
nand UO_833 (O_833,N_29924,N_29930);
nor UO_834 (O_834,N_29832,N_29821);
and UO_835 (O_835,N_29820,N_29960);
nor UO_836 (O_836,N_29874,N_29710);
nor UO_837 (O_837,N_29873,N_29704);
nand UO_838 (O_838,N_29802,N_29738);
and UO_839 (O_839,N_29713,N_29986);
or UO_840 (O_840,N_29925,N_29919);
and UO_841 (O_841,N_29799,N_29998);
nor UO_842 (O_842,N_29912,N_29738);
and UO_843 (O_843,N_29806,N_29810);
xnor UO_844 (O_844,N_29801,N_29784);
nand UO_845 (O_845,N_29718,N_29923);
or UO_846 (O_846,N_29998,N_29938);
or UO_847 (O_847,N_29874,N_29878);
xor UO_848 (O_848,N_29822,N_29883);
xnor UO_849 (O_849,N_29969,N_29961);
xor UO_850 (O_850,N_29769,N_29774);
nor UO_851 (O_851,N_29932,N_29970);
xor UO_852 (O_852,N_29708,N_29894);
or UO_853 (O_853,N_29767,N_29866);
and UO_854 (O_854,N_29818,N_29742);
nand UO_855 (O_855,N_29793,N_29843);
nand UO_856 (O_856,N_29992,N_29794);
and UO_857 (O_857,N_29709,N_29987);
xnor UO_858 (O_858,N_29978,N_29873);
nand UO_859 (O_859,N_29863,N_29882);
or UO_860 (O_860,N_29760,N_29978);
nand UO_861 (O_861,N_29999,N_29876);
and UO_862 (O_862,N_29971,N_29767);
nand UO_863 (O_863,N_29863,N_29819);
or UO_864 (O_864,N_29805,N_29980);
xor UO_865 (O_865,N_29829,N_29824);
or UO_866 (O_866,N_29929,N_29706);
or UO_867 (O_867,N_29916,N_29807);
and UO_868 (O_868,N_29729,N_29825);
or UO_869 (O_869,N_29905,N_29868);
or UO_870 (O_870,N_29755,N_29845);
and UO_871 (O_871,N_29838,N_29726);
nor UO_872 (O_872,N_29986,N_29906);
nand UO_873 (O_873,N_29879,N_29753);
and UO_874 (O_874,N_29993,N_29847);
nor UO_875 (O_875,N_29945,N_29822);
or UO_876 (O_876,N_29804,N_29984);
xnor UO_877 (O_877,N_29789,N_29824);
and UO_878 (O_878,N_29985,N_29980);
xor UO_879 (O_879,N_29931,N_29873);
and UO_880 (O_880,N_29767,N_29813);
nand UO_881 (O_881,N_29962,N_29738);
or UO_882 (O_882,N_29992,N_29895);
or UO_883 (O_883,N_29905,N_29764);
xnor UO_884 (O_884,N_29741,N_29799);
and UO_885 (O_885,N_29891,N_29717);
nor UO_886 (O_886,N_29923,N_29854);
or UO_887 (O_887,N_29864,N_29999);
xnor UO_888 (O_888,N_29999,N_29824);
nor UO_889 (O_889,N_29973,N_29984);
nor UO_890 (O_890,N_29945,N_29947);
and UO_891 (O_891,N_29859,N_29946);
xor UO_892 (O_892,N_29786,N_29906);
nand UO_893 (O_893,N_29775,N_29799);
or UO_894 (O_894,N_29820,N_29828);
or UO_895 (O_895,N_29858,N_29962);
and UO_896 (O_896,N_29917,N_29746);
nand UO_897 (O_897,N_29950,N_29785);
nand UO_898 (O_898,N_29859,N_29737);
or UO_899 (O_899,N_29884,N_29832);
or UO_900 (O_900,N_29908,N_29907);
or UO_901 (O_901,N_29840,N_29849);
xor UO_902 (O_902,N_29763,N_29707);
or UO_903 (O_903,N_29994,N_29918);
nand UO_904 (O_904,N_29969,N_29821);
nand UO_905 (O_905,N_29710,N_29739);
and UO_906 (O_906,N_29718,N_29713);
or UO_907 (O_907,N_29822,N_29724);
nor UO_908 (O_908,N_29719,N_29871);
and UO_909 (O_909,N_29779,N_29942);
nand UO_910 (O_910,N_29867,N_29725);
nand UO_911 (O_911,N_29778,N_29821);
nor UO_912 (O_912,N_29756,N_29837);
nand UO_913 (O_913,N_29991,N_29874);
or UO_914 (O_914,N_29816,N_29871);
xor UO_915 (O_915,N_29805,N_29752);
nand UO_916 (O_916,N_29960,N_29767);
and UO_917 (O_917,N_29889,N_29720);
xnor UO_918 (O_918,N_29853,N_29931);
nor UO_919 (O_919,N_29965,N_29911);
xnor UO_920 (O_920,N_29833,N_29831);
nor UO_921 (O_921,N_29918,N_29866);
or UO_922 (O_922,N_29936,N_29989);
xor UO_923 (O_923,N_29835,N_29824);
xor UO_924 (O_924,N_29856,N_29800);
nand UO_925 (O_925,N_29945,N_29810);
and UO_926 (O_926,N_29995,N_29797);
and UO_927 (O_927,N_29818,N_29878);
nand UO_928 (O_928,N_29782,N_29892);
xor UO_929 (O_929,N_29954,N_29966);
or UO_930 (O_930,N_29932,N_29765);
xor UO_931 (O_931,N_29990,N_29983);
or UO_932 (O_932,N_29784,N_29884);
nand UO_933 (O_933,N_29748,N_29773);
and UO_934 (O_934,N_29757,N_29728);
nor UO_935 (O_935,N_29712,N_29900);
nor UO_936 (O_936,N_29959,N_29793);
or UO_937 (O_937,N_29958,N_29779);
and UO_938 (O_938,N_29811,N_29898);
and UO_939 (O_939,N_29779,N_29765);
or UO_940 (O_940,N_29878,N_29717);
and UO_941 (O_941,N_29717,N_29748);
nor UO_942 (O_942,N_29754,N_29802);
xor UO_943 (O_943,N_29774,N_29707);
or UO_944 (O_944,N_29756,N_29946);
nor UO_945 (O_945,N_29705,N_29938);
nor UO_946 (O_946,N_29874,N_29864);
or UO_947 (O_947,N_29705,N_29777);
nor UO_948 (O_948,N_29998,N_29894);
or UO_949 (O_949,N_29757,N_29891);
nor UO_950 (O_950,N_29919,N_29830);
xor UO_951 (O_951,N_29765,N_29840);
xor UO_952 (O_952,N_29934,N_29839);
nor UO_953 (O_953,N_29835,N_29787);
nand UO_954 (O_954,N_29922,N_29914);
nand UO_955 (O_955,N_29872,N_29751);
and UO_956 (O_956,N_29837,N_29776);
or UO_957 (O_957,N_29902,N_29863);
and UO_958 (O_958,N_29775,N_29764);
or UO_959 (O_959,N_29700,N_29739);
nor UO_960 (O_960,N_29869,N_29733);
and UO_961 (O_961,N_29828,N_29924);
or UO_962 (O_962,N_29908,N_29773);
nand UO_963 (O_963,N_29791,N_29997);
or UO_964 (O_964,N_29892,N_29908);
or UO_965 (O_965,N_29937,N_29737);
or UO_966 (O_966,N_29935,N_29899);
or UO_967 (O_967,N_29949,N_29976);
xnor UO_968 (O_968,N_29954,N_29933);
xor UO_969 (O_969,N_29999,N_29815);
xnor UO_970 (O_970,N_29834,N_29796);
or UO_971 (O_971,N_29985,N_29902);
nand UO_972 (O_972,N_29828,N_29970);
and UO_973 (O_973,N_29971,N_29989);
xor UO_974 (O_974,N_29988,N_29811);
nand UO_975 (O_975,N_29726,N_29957);
nor UO_976 (O_976,N_29762,N_29877);
nand UO_977 (O_977,N_29891,N_29925);
nand UO_978 (O_978,N_29897,N_29709);
or UO_979 (O_979,N_29952,N_29824);
xnor UO_980 (O_980,N_29702,N_29907);
nor UO_981 (O_981,N_29807,N_29991);
nand UO_982 (O_982,N_29975,N_29783);
nand UO_983 (O_983,N_29768,N_29996);
nand UO_984 (O_984,N_29853,N_29948);
nor UO_985 (O_985,N_29817,N_29743);
nor UO_986 (O_986,N_29762,N_29892);
nor UO_987 (O_987,N_29811,N_29903);
xor UO_988 (O_988,N_29726,N_29892);
xor UO_989 (O_989,N_29890,N_29889);
or UO_990 (O_990,N_29719,N_29704);
and UO_991 (O_991,N_29757,N_29898);
or UO_992 (O_992,N_29740,N_29818);
nor UO_993 (O_993,N_29887,N_29980);
nand UO_994 (O_994,N_29862,N_29982);
nor UO_995 (O_995,N_29921,N_29841);
and UO_996 (O_996,N_29748,N_29909);
xnor UO_997 (O_997,N_29990,N_29931);
or UO_998 (O_998,N_29973,N_29726);
xor UO_999 (O_999,N_29841,N_29824);
xnor UO_1000 (O_1000,N_29833,N_29774);
nand UO_1001 (O_1001,N_29982,N_29819);
or UO_1002 (O_1002,N_29821,N_29806);
nand UO_1003 (O_1003,N_29928,N_29785);
nand UO_1004 (O_1004,N_29752,N_29838);
nor UO_1005 (O_1005,N_29805,N_29709);
and UO_1006 (O_1006,N_29950,N_29824);
xor UO_1007 (O_1007,N_29881,N_29916);
and UO_1008 (O_1008,N_29726,N_29747);
and UO_1009 (O_1009,N_29840,N_29753);
xnor UO_1010 (O_1010,N_29866,N_29812);
nor UO_1011 (O_1011,N_29897,N_29811);
nor UO_1012 (O_1012,N_29831,N_29905);
nor UO_1013 (O_1013,N_29902,N_29920);
nand UO_1014 (O_1014,N_29706,N_29956);
nand UO_1015 (O_1015,N_29985,N_29910);
nor UO_1016 (O_1016,N_29835,N_29972);
nor UO_1017 (O_1017,N_29846,N_29787);
and UO_1018 (O_1018,N_29962,N_29898);
xor UO_1019 (O_1019,N_29726,N_29878);
and UO_1020 (O_1020,N_29907,N_29856);
xor UO_1021 (O_1021,N_29992,N_29899);
nand UO_1022 (O_1022,N_29974,N_29905);
xor UO_1023 (O_1023,N_29857,N_29842);
or UO_1024 (O_1024,N_29820,N_29735);
nor UO_1025 (O_1025,N_29725,N_29792);
nor UO_1026 (O_1026,N_29817,N_29802);
xnor UO_1027 (O_1027,N_29713,N_29811);
xnor UO_1028 (O_1028,N_29706,N_29992);
nor UO_1029 (O_1029,N_29913,N_29954);
and UO_1030 (O_1030,N_29794,N_29972);
nor UO_1031 (O_1031,N_29791,N_29797);
or UO_1032 (O_1032,N_29713,N_29973);
or UO_1033 (O_1033,N_29898,N_29997);
or UO_1034 (O_1034,N_29867,N_29890);
xnor UO_1035 (O_1035,N_29930,N_29975);
nor UO_1036 (O_1036,N_29821,N_29731);
and UO_1037 (O_1037,N_29900,N_29780);
nor UO_1038 (O_1038,N_29796,N_29739);
xor UO_1039 (O_1039,N_29873,N_29890);
nand UO_1040 (O_1040,N_29976,N_29930);
or UO_1041 (O_1041,N_29789,N_29989);
and UO_1042 (O_1042,N_29928,N_29814);
xnor UO_1043 (O_1043,N_29922,N_29769);
xnor UO_1044 (O_1044,N_29934,N_29880);
xnor UO_1045 (O_1045,N_29757,N_29729);
xor UO_1046 (O_1046,N_29930,N_29887);
nor UO_1047 (O_1047,N_29859,N_29735);
xnor UO_1048 (O_1048,N_29707,N_29950);
nor UO_1049 (O_1049,N_29844,N_29955);
nand UO_1050 (O_1050,N_29848,N_29786);
nor UO_1051 (O_1051,N_29803,N_29853);
nand UO_1052 (O_1052,N_29838,N_29709);
or UO_1053 (O_1053,N_29971,N_29850);
and UO_1054 (O_1054,N_29912,N_29715);
nor UO_1055 (O_1055,N_29956,N_29948);
nand UO_1056 (O_1056,N_29966,N_29934);
nand UO_1057 (O_1057,N_29822,N_29746);
and UO_1058 (O_1058,N_29755,N_29948);
or UO_1059 (O_1059,N_29899,N_29957);
and UO_1060 (O_1060,N_29838,N_29887);
nand UO_1061 (O_1061,N_29747,N_29841);
or UO_1062 (O_1062,N_29737,N_29722);
or UO_1063 (O_1063,N_29761,N_29817);
nand UO_1064 (O_1064,N_29926,N_29858);
nand UO_1065 (O_1065,N_29968,N_29737);
or UO_1066 (O_1066,N_29863,N_29752);
nand UO_1067 (O_1067,N_29979,N_29705);
nor UO_1068 (O_1068,N_29916,N_29837);
nor UO_1069 (O_1069,N_29911,N_29764);
nand UO_1070 (O_1070,N_29750,N_29822);
or UO_1071 (O_1071,N_29848,N_29762);
and UO_1072 (O_1072,N_29715,N_29922);
or UO_1073 (O_1073,N_29948,N_29904);
or UO_1074 (O_1074,N_29731,N_29799);
nor UO_1075 (O_1075,N_29714,N_29827);
nand UO_1076 (O_1076,N_29972,N_29770);
nand UO_1077 (O_1077,N_29783,N_29824);
nand UO_1078 (O_1078,N_29864,N_29856);
and UO_1079 (O_1079,N_29853,N_29770);
nor UO_1080 (O_1080,N_29803,N_29896);
nor UO_1081 (O_1081,N_29833,N_29908);
nand UO_1082 (O_1082,N_29888,N_29837);
or UO_1083 (O_1083,N_29987,N_29756);
or UO_1084 (O_1084,N_29757,N_29809);
or UO_1085 (O_1085,N_29816,N_29969);
or UO_1086 (O_1086,N_29889,N_29912);
and UO_1087 (O_1087,N_29712,N_29880);
xnor UO_1088 (O_1088,N_29816,N_29954);
and UO_1089 (O_1089,N_29810,N_29919);
nor UO_1090 (O_1090,N_29806,N_29803);
nor UO_1091 (O_1091,N_29838,N_29916);
nor UO_1092 (O_1092,N_29810,N_29848);
or UO_1093 (O_1093,N_29928,N_29889);
nor UO_1094 (O_1094,N_29906,N_29719);
or UO_1095 (O_1095,N_29734,N_29884);
or UO_1096 (O_1096,N_29960,N_29826);
nand UO_1097 (O_1097,N_29740,N_29876);
xnor UO_1098 (O_1098,N_29737,N_29745);
nand UO_1099 (O_1099,N_29801,N_29872);
nor UO_1100 (O_1100,N_29829,N_29704);
nand UO_1101 (O_1101,N_29882,N_29779);
nand UO_1102 (O_1102,N_29718,N_29873);
or UO_1103 (O_1103,N_29763,N_29881);
xnor UO_1104 (O_1104,N_29855,N_29975);
xor UO_1105 (O_1105,N_29772,N_29748);
xnor UO_1106 (O_1106,N_29902,N_29869);
or UO_1107 (O_1107,N_29799,N_29934);
nand UO_1108 (O_1108,N_29976,N_29848);
and UO_1109 (O_1109,N_29989,N_29719);
xnor UO_1110 (O_1110,N_29788,N_29979);
or UO_1111 (O_1111,N_29869,N_29789);
or UO_1112 (O_1112,N_29889,N_29896);
nor UO_1113 (O_1113,N_29852,N_29967);
nor UO_1114 (O_1114,N_29909,N_29971);
xnor UO_1115 (O_1115,N_29909,N_29894);
and UO_1116 (O_1116,N_29880,N_29749);
or UO_1117 (O_1117,N_29983,N_29740);
nor UO_1118 (O_1118,N_29981,N_29876);
and UO_1119 (O_1119,N_29925,N_29714);
and UO_1120 (O_1120,N_29885,N_29713);
xnor UO_1121 (O_1121,N_29837,N_29786);
and UO_1122 (O_1122,N_29981,N_29875);
xor UO_1123 (O_1123,N_29962,N_29861);
nand UO_1124 (O_1124,N_29742,N_29920);
nor UO_1125 (O_1125,N_29745,N_29872);
and UO_1126 (O_1126,N_29836,N_29965);
nand UO_1127 (O_1127,N_29780,N_29705);
nor UO_1128 (O_1128,N_29968,N_29972);
and UO_1129 (O_1129,N_29990,N_29799);
or UO_1130 (O_1130,N_29744,N_29739);
nor UO_1131 (O_1131,N_29706,N_29854);
nand UO_1132 (O_1132,N_29709,N_29729);
or UO_1133 (O_1133,N_29905,N_29715);
nand UO_1134 (O_1134,N_29828,N_29764);
or UO_1135 (O_1135,N_29841,N_29729);
nor UO_1136 (O_1136,N_29930,N_29981);
nor UO_1137 (O_1137,N_29816,N_29789);
or UO_1138 (O_1138,N_29935,N_29920);
xor UO_1139 (O_1139,N_29916,N_29803);
nor UO_1140 (O_1140,N_29994,N_29907);
nand UO_1141 (O_1141,N_29788,N_29726);
and UO_1142 (O_1142,N_29921,N_29833);
nand UO_1143 (O_1143,N_29740,N_29797);
or UO_1144 (O_1144,N_29930,N_29804);
xnor UO_1145 (O_1145,N_29806,N_29981);
xnor UO_1146 (O_1146,N_29896,N_29918);
nand UO_1147 (O_1147,N_29704,N_29976);
or UO_1148 (O_1148,N_29878,N_29707);
and UO_1149 (O_1149,N_29701,N_29793);
or UO_1150 (O_1150,N_29980,N_29897);
xnor UO_1151 (O_1151,N_29808,N_29884);
and UO_1152 (O_1152,N_29858,N_29947);
nor UO_1153 (O_1153,N_29750,N_29917);
or UO_1154 (O_1154,N_29825,N_29912);
nor UO_1155 (O_1155,N_29839,N_29989);
nand UO_1156 (O_1156,N_29918,N_29776);
or UO_1157 (O_1157,N_29796,N_29872);
nor UO_1158 (O_1158,N_29956,N_29791);
and UO_1159 (O_1159,N_29913,N_29728);
nand UO_1160 (O_1160,N_29759,N_29854);
nand UO_1161 (O_1161,N_29888,N_29854);
or UO_1162 (O_1162,N_29990,N_29923);
nand UO_1163 (O_1163,N_29804,N_29810);
xor UO_1164 (O_1164,N_29772,N_29901);
or UO_1165 (O_1165,N_29905,N_29965);
or UO_1166 (O_1166,N_29811,N_29906);
nand UO_1167 (O_1167,N_29980,N_29716);
and UO_1168 (O_1168,N_29903,N_29785);
xnor UO_1169 (O_1169,N_29821,N_29792);
and UO_1170 (O_1170,N_29754,N_29752);
nand UO_1171 (O_1171,N_29963,N_29802);
and UO_1172 (O_1172,N_29992,N_29947);
or UO_1173 (O_1173,N_29837,N_29866);
nor UO_1174 (O_1174,N_29756,N_29986);
nand UO_1175 (O_1175,N_29733,N_29800);
nand UO_1176 (O_1176,N_29824,N_29758);
xor UO_1177 (O_1177,N_29920,N_29962);
nand UO_1178 (O_1178,N_29851,N_29700);
xnor UO_1179 (O_1179,N_29977,N_29804);
or UO_1180 (O_1180,N_29716,N_29755);
nor UO_1181 (O_1181,N_29779,N_29964);
and UO_1182 (O_1182,N_29838,N_29760);
nand UO_1183 (O_1183,N_29737,N_29775);
nand UO_1184 (O_1184,N_29704,N_29907);
xnor UO_1185 (O_1185,N_29806,N_29959);
nor UO_1186 (O_1186,N_29894,N_29781);
and UO_1187 (O_1187,N_29859,N_29777);
xor UO_1188 (O_1188,N_29969,N_29767);
and UO_1189 (O_1189,N_29851,N_29997);
nand UO_1190 (O_1190,N_29702,N_29936);
xnor UO_1191 (O_1191,N_29913,N_29761);
nor UO_1192 (O_1192,N_29971,N_29912);
xor UO_1193 (O_1193,N_29839,N_29921);
and UO_1194 (O_1194,N_29933,N_29939);
xnor UO_1195 (O_1195,N_29791,N_29822);
nor UO_1196 (O_1196,N_29885,N_29776);
nand UO_1197 (O_1197,N_29928,N_29825);
xor UO_1198 (O_1198,N_29781,N_29776);
nand UO_1199 (O_1199,N_29909,N_29921);
nand UO_1200 (O_1200,N_29842,N_29733);
xor UO_1201 (O_1201,N_29919,N_29767);
or UO_1202 (O_1202,N_29763,N_29721);
nand UO_1203 (O_1203,N_29783,N_29877);
nand UO_1204 (O_1204,N_29727,N_29931);
nand UO_1205 (O_1205,N_29801,N_29971);
or UO_1206 (O_1206,N_29999,N_29851);
and UO_1207 (O_1207,N_29933,N_29952);
nand UO_1208 (O_1208,N_29859,N_29883);
nand UO_1209 (O_1209,N_29933,N_29955);
nor UO_1210 (O_1210,N_29878,N_29778);
or UO_1211 (O_1211,N_29799,N_29961);
xnor UO_1212 (O_1212,N_29815,N_29943);
and UO_1213 (O_1213,N_29891,N_29947);
nand UO_1214 (O_1214,N_29855,N_29907);
or UO_1215 (O_1215,N_29872,N_29907);
xnor UO_1216 (O_1216,N_29755,N_29746);
nor UO_1217 (O_1217,N_29842,N_29751);
or UO_1218 (O_1218,N_29884,N_29865);
nor UO_1219 (O_1219,N_29713,N_29719);
nand UO_1220 (O_1220,N_29793,N_29818);
xnor UO_1221 (O_1221,N_29805,N_29824);
and UO_1222 (O_1222,N_29976,N_29876);
and UO_1223 (O_1223,N_29795,N_29710);
or UO_1224 (O_1224,N_29716,N_29949);
nor UO_1225 (O_1225,N_29987,N_29851);
xnor UO_1226 (O_1226,N_29765,N_29843);
and UO_1227 (O_1227,N_29952,N_29898);
and UO_1228 (O_1228,N_29775,N_29802);
xor UO_1229 (O_1229,N_29895,N_29964);
and UO_1230 (O_1230,N_29928,N_29963);
nor UO_1231 (O_1231,N_29711,N_29758);
and UO_1232 (O_1232,N_29752,N_29915);
and UO_1233 (O_1233,N_29894,N_29824);
nand UO_1234 (O_1234,N_29824,N_29840);
nand UO_1235 (O_1235,N_29906,N_29984);
and UO_1236 (O_1236,N_29705,N_29772);
or UO_1237 (O_1237,N_29882,N_29958);
or UO_1238 (O_1238,N_29983,N_29844);
xnor UO_1239 (O_1239,N_29863,N_29828);
and UO_1240 (O_1240,N_29788,N_29743);
nor UO_1241 (O_1241,N_29730,N_29717);
or UO_1242 (O_1242,N_29821,N_29910);
and UO_1243 (O_1243,N_29955,N_29764);
and UO_1244 (O_1244,N_29980,N_29945);
nor UO_1245 (O_1245,N_29877,N_29956);
nand UO_1246 (O_1246,N_29945,N_29770);
nor UO_1247 (O_1247,N_29862,N_29746);
nand UO_1248 (O_1248,N_29959,N_29962);
nor UO_1249 (O_1249,N_29886,N_29837);
or UO_1250 (O_1250,N_29716,N_29826);
xor UO_1251 (O_1251,N_29705,N_29860);
nand UO_1252 (O_1252,N_29838,N_29941);
and UO_1253 (O_1253,N_29724,N_29838);
nand UO_1254 (O_1254,N_29896,N_29898);
nor UO_1255 (O_1255,N_29730,N_29719);
nand UO_1256 (O_1256,N_29876,N_29857);
or UO_1257 (O_1257,N_29825,N_29952);
nand UO_1258 (O_1258,N_29970,N_29964);
xor UO_1259 (O_1259,N_29924,N_29863);
nand UO_1260 (O_1260,N_29846,N_29948);
xnor UO_1261 (O_1261,N_29818,N_29867);
or UO_1262 (O_1262,N_29864,N_29836);
nand UO_1263 (O_1263,N_29987,N_29976);
xor UO_1264 (O_1264,N_29932,N_29915);
nor UO_1265 (O_1265,N_29954,N_29712);
nand UO_1266 (O_1266,N_29988,N_29770);
nor UO_1267 (O_1267,N_29869,N_29940);
xor UO_1268 (O_1268,N_29727,N_29701);
nor UO_1269 (O_1269,N_29926,N_29901);
nand UO_1270 (O_1270,N_29854,N_29932);
nand UO_1271 (O_1271,N_29867,N_29798);
or UO_1272 (O_1272,N_29723,N_29924);
or UO_1273 (O_1273,N_29706,N_29792);
nand UO_1274 (O_1274,N_29790,N_29711);
nand UO_1275 (O_1275,N_29715,N_29851);
xor UO_1276 (O_1276,N_29764,N_29714);
nand UO_1277 (O_1277,N_29719,N_29876);
and UO_1278 (O_1278,N_29864,N_29786);
nor UO_1279 (O_1279,N_29725,N_29712);
nand UO_1280 (O_1280,N_29896,N_29932);
and UO_1281 (O_1281,N_29872,N_29858);
and UO_1282 (O_1282,N_29842,N_29759);
and UO_1283 (O_1283,N_29723,N_29973);
and UO_1284 (O_1284,N_29985,N_29862);
xnor UO_1285 (O_1285,N_29964,N_29969);
xor UO_1286 (O_1286,N_29841,N_29788);
nor UO_1287 (O_1287,N_29942,N_29919);
nor UO_1288 (O_1288,N_29817,N_29810);
nand UO_1289 (O_1289,N_29968,N_29985);
or UO_1290 (O_1290,N_29860,N_29784);
nor UO_1291 (O_1291,N_29904,N_29700);
and UO_1292 (O_1292,N_29851,N_29850);
and UO_1293 (O_1293,N_29999,N_29805);
or UO_1294 (O_1294,N_29943,N_29990);
xnor UO_1295 (O_1295,N_29876,N_29836);
nor UO_1296 (O_1296,N_29919,N_29852);
nand UO_1297 (O_1297,N_29747,N_29893);
xnor UO_1298 (O_1298,N_29876,N_29865);
and UO_1299 (O_1299,N_29842,N_29773);
xor UO_1300 (O_1300,N_29916,N_29845);
nor UO_1301 (O_1301,N_29767,N_29911);
nor UO_1302 (O_1302,N_29839,N_29991);
nand UO_1303 (O_1303,N_29865,N_29701);
nor UO_1304 (O_1304,N_29704,N_29736);
nor UO_1305 (O_1305,N_29992,N_29752);
or UO_1306 (O_1306,N_29953,N_29720);
or UO_1307 (O_1307,N_29848,N_29720);
xnor UO_1308 (O_1308,N_29929,N_29947);
or UO_1309 (O_1309,N_29998,N_29740);
nand UO_1310 (O_1310,N_29840,N_29959);
or UO_1311 (O_1311,N_29858,N_29838);
nor UO_1312 (O_1312,N_29827,N_29746);
nor UO_1313 (O_1313,N_29731,N_29824);
or UO_1314 (O_1314,N_29859,N_29814);
nand UO_1315 (O_1315,N_29780,N_29861);
xnor UO_1316 (O_1316,N_29864,N_29958);
nor UO_1317 (O_1317,N_29741,N_29994);
and UO_1318 (O_1318,N_29930,N_29791);
nor UO_1319 (O_1319,N_29926,N_29748);
nor UO_1320 (O_1320,N_29707,N_29889);
xnor UO_1321 (O_1321,N_29773,N_29910);
nor UO_1322 (O_1322,N_29892,N_29889);
nand UO_1323 (O_1323,N_29947,N_29843);
or UO_1324 (O_1324,N_29976,N_29724);
or UO_1325 (O_1325,N_29799,N_29931);
xnor UO_1326 (O_1326,N_29910,N_29923);
xnor UO_1327 (O_1327,N_29946,N_29841);
nor UO_1328 (O_1328,N_29760,N_29750);
or UO_1329 (O_1329,N_29929,N_29977);
and UO_1330 (O_1330,N_29782,N_29852);
or UO_1331 (O_1331,N_29976,N_29805);
nor UO_1332 (O_1332,N_29875,N_29998);
or UO_1333 (O_1333,N_29782,N_29974);
xor UO_1334 (O_1334,N_29709,N_29837);
xor UO_1335 (O_1335,N_29838,N_29889);
xnor UO_1336 (O_1336,N_29931,N_29747);
nor UO_1337 (O_1337,N_29843,N_29885);
nor UO_1338 (O_1338,N_29866,N_29868);
or UO_1339 (O_1339,N_29779,N_29906);
nor UO_1340 (O_1340,N_29941,N_29960);
xor UO_1341 (O_1341,N_29997,N_29715);
nand UO_1342 (O_1342,N_29851,N_29705);
nand UO_1343 (O_1343,N_29741,N_29915);
xor UO_1344 (O_1344,N_29999,N_29797);
nand UO_1345 (O_1345,N_29902,N_29992);
xor UO_1346 (O_1346,N_29778,N_29999);
nor UO_1347 (O_1347,N_29883,N_29795);
nor UO_1348 (O_1348,N_29835,N_29872);
xnor UO_1349 (O_1349,N_29755,N_29700);
nor UO_1350 (O_1350,N_29910,N_29825);
or UO_1351 (O_1351,N_29979,N_29776);
nand UO_1352 (O_1352,N_29903,N_29925);
xnor UO_1353 (O_1353,N_29819,N_29867);
and UO_1354 (O_1354,N_29717,N_29835);
xnor UO_1355 (O_1355,N_29821,N_29906);
and UO_1356 (O_1356,N_29755,N_29761);
or UO_1357 (O_1357,N_29740,N_29727);
xor UO_1358 (O_1358,N_29797,N_29966);
nor UO_1359 (O_1359,N_29736,N_29936);
or UO_1360 (O_1360,N_29863,N_29918);
nor UO_1361 (O_1361,N_29902,N_29935);
xor UO_1362 (O_1362,N_29925,N_29949);
nor UO_1363 (O_1363,N_29893,N_29771);
nor UO_1364 (O_1364,N_29988,N_29882);
or UO_1365 (O_1365,N_29782,N_29963);
and UO_1366 (O_1366,N_29926,N_29954);
nand UO_1367 (O_1367,N_29930,N_29826);
xnor UO_1368 (O_1368,N_29750,N_29744);
nand UO_1369 (O_1369,N_29798,N_29786);
xor UO_1370 (O_1370,N_29860,N_29902);
and UO_1371 (O_1371,N_29989,N_29896);
nand UO_1372 (O_1372,N_29844,N_29957);
or UO_1373 (O_1373,N_29962,N_29785);
and UO_1374 (O_1374,N_29792,N_29958);
or UO_1375 (O_1375,N_29842,N_29783);
xor UO_1376 (O_1376,N_29730,N_29963);
nor UO_1377 (O_1377,N_29992,N_29746);
xnor UO_1378 (O_1378,N_29791,N_29814);
nand UO_1379 (O_1379,N_29910,N_29860);
or UO_1380 (O_1380,N_29905,N_29893);
nand UO_1381 (O_1381,N_29720,N_29804);
xor UO_1382 (O_1382,N_29745,N_29708);
nand UO_1383 (O_1383,N_29854,N_29720);
and UO_1384 (O_1384,N_29707,N_29992);
nand UO_1385 (O_1385,N_29797,N_29856);
nor UO_1386 (O_1386,N_29900,N_29948);
and UO_1387 (O_1387,N_29870,N_29702);
xnor UO_1388 (O_1388,N_29965,N_29724);
nand UO_1389 (O_1389,N_29882,N_29979);
or UO_1390 (O_1390,N_29836,N_29742);
nand UO_1391 (O_1391,N_29943,N_29845);
nor UO_1392 (O_1392,N_29805,N_29706);
nand UO_1393 (O_1393,N_29701,N_29928);
and UO_1394 (O_1394,N_29812,N_29729);
and UO_1395 (O_1395,N_29848,N_29790);
nor UO_1396 (O_1396,N_29997,N_29771);
and UO_1397 (O_1397,N_29832,N_29962);
nand UO_1398 (O_1398,N_29792,N_29908);
nor UO_1399 (O_1399,N_29707,N_29969);
nor UO_1400 (O_1400,N_29827,N_29753);
or UO_1401 (O_1401,N_29928,N_29773);
or UO_1402 (O_1402,N_29968,N_29939);
xor UO_1403 (O_1403,N_29797,N_29824);
and UO_1404 (O_1404,N_29906,N_29725);
nor UO_1405 (O_1405,N_29737,N_29772);
and UO_1406 (O_1406,N_29966,N_29889);
nor UO_1407 (O_1407,N_29781,N_29741);
nor UO_1408 (O_1408,N_29831,N_29973);
and UO_1409 (O_1409,N_29724,N_29835);
nor UO_1410 (O_1410,N_29834,N_29811);
nand UO_1411 (O_1411,N_29891,N_29743);
or UO_1412 (O_1412,N_29841,N_29760);
xnor UO_1413 (O_1413,N_29897,N_29928);
xnor UO_1414 (O_1414,N_29709,N_29848);
nor UO_1415 (O_1415,N_29846,N_29874);
and UO_1416 (O_1416,N_29749,N_29745);
xnor UO_1417 (O_1417,N_29961,N_29769);
nor UO_1418 (O_1418,N_29860,N_29998);
nand UO_1419 (O_1419,N_29880,N_29968);
or UO_1420 (O_1420,N_29986,N_29757);
or UO_1421 (O_1421,N_29774,N_29882);
nor UO_1422 (O_1422,N_29964,N_29788);
nor UO_1423 (O_1423,N_29826,N_29866);
nor UO_1424 (O_1424,N_29955,N_29727);
or UO_1425 (O_1425,N_29852,N_29989);
and UO_1426 (O_1426,N_29781,N_29983);
xor UO_1427 (O_1427,N_29978,N_29777);
and UO_1428 (O_1428,N_29910,N_29705);
nor UO_1429 (O_1429,N_29962,N_29988);
nand UO_1430 (O_1430,N_29937,N_29824);
nor UO_1431 (O_1431,N_29714,N_29845);
or UO_1432 (O_1432,N_29730,N_29809);
or UO_1433 (O_1433,N_29709,N_29714);
xor UO_1434 (O_1434,N_29973,N_29721);
nand UO_1435 (O_1435,N_29798,N_29851);
xor UO_1436 (O_1436,N_29811,N_29973);
nor UO_1437 (O_1437,N_29862,N_29903);
xnor UO_1438 (O_1438,N_29935,N_29933);
or UO_1439 (O_1439,N_29959,N_29735);
or UO_1440 (O_1440,N_29950,N_29936);
nand UO_1441 (O_1441,N_29757,N_29737);
or UO_1442 (O_1442,N_29789,N_29978);
or UO_1443 (O_1443,N_29777,N_29808);
or UO_1444 (O_1444,N_29758,N_29845);
nand UO_1445 (O_1445,N_29707,N_29937);
xor UO_1446 (O_1446,N_29904,N_29838);
xnor UO_1447 (O_1447,N_29959,N_29855);
or UO_1448 (O_1448,N_29707,N_29970);
and UO_1449 (O_1449,N_29702,N_29771);
nor UO_1450 (O_1450,N_29958,N_29900);
and UO_1451 (O_1451,N_29724,N_29996);
and UO_1452 (O_1452,N_29844,N_29903);
or UO_1453 (O_1453,N_29852,N_29802);
and UO_1454 (O_1454,N_29962,N_29823);
nand UO_1455 (O_1455,N_29966,N_29743);
xor UO_1456 (O_1456,N_29934,N_29922);
xnor UO_1457 (O_1457,N_29777,N_29708);
nor UO_1458 (O_1458,N_29880,N_29894);
xor UO_1459 (O_1459,N_29812,N_29875);
xnor UO_1460 (O_1460,N_29782,N_29741);
nor UO_1461 (O_1461,N_29819,N_29840);
xor UO_1462 (O_1462,N_29962,N_29716);
nand UO_1463 (O_1463,N_29884,N_29728);
nor UO_1464 (O_1464,N_29830,N_29891);
xor UO_1465 (O_1465,N_29701,N_29825);
and UO_1466 (O_1466,N_29950,N_29817);
and UO_1467 (O_1467,N_29723,N_29857);
nand UO_1468 (O_1468,N_29844,N_29766);
or UO_1469 (O_1469,N_29709,N_29734);
xor UO_1470 (O_1470,N_29826,N_29993);
nor UO_1471 (O_1471,N_29912,N_29795);
and UO_1472 (O_1472,N_29802,N_29971);
and UO_1473 (O_1473,N_29824,N_29859);
xnor UO_1474 (O_1474,N_29802,N_29764);
nor UO_1475 (O_1475,N_29895,N_29723);
or UO_1476 (O_1476,N_29826,N_29789);
and UO_1477 (O_1477,N_29726,N_29704);
nand UO_1478 (O_1478,N_29767,N_29771);
xnor UO_1479 (O_1479,N_29904,N_29912);
and UO_1480 (O_1480,N_29737,N_29969);
and UO_1481 (O_1481,N_29719,N_29949);
nor UO_1482 (O_1482,N_29826,N_29957);
or UO_1483 (O_1483,N_29945,N_29712);
or UO_1484 (O_1484,N_29869,N_29916);
or UO_1485 (O_1485,N_29861,N_29952);
or UO_1486 (O_1486,N_29921,N_29765);
and UO_1487 (O_1487,N_29714,N_29966);
nand UO_1488 (O_1488,N_29932,N_29871);
nor UO_1489 (O_1489,N_29818,N_29768);
xor UO_1490 (O_1490,N_29902,N_29881);
nand UO_1491 (O_1491,N_29752,N_29832);
xor UO_1492 (O_1492,N_29742,N_29936);
nor UO_1493 (O_1493,N_29817,N_29714);
or UO_1494 (O_1494,N_29906,N_29754);
xor UO_1495 (O_1495,N_29959,N_29769);
or UO_1496 (O_1496,N_29959,N_29870);
or UO_1497 (O_1497,N_29903,N_29894);
xor UO_1498 (O_1498,N_29782,N_29954);
or UO_1499 (O_1499,N_29797,N_29708);
nor UO_1500 (O_1500,N_29750,N_29739);
nand UO_1501 (O_1501,N_29924,N_29998);
and UO_1502 (O_1502,N_29798,N_29795);
and UO_1503 (O_1503,N_29829,N_29807);
nand UO_1504 (O_1504,N_29812,N_29748);
nor UO_1505 (O_1505,N_29752,N_29700);
or UO_1506 (O_1506,N_29955,N_29816);
xnor UO_1507 (O_1507,N_29818,N_29952);
and UO_1508 (O_1508,N_29758,N_29720);
nand UO_1509 (O_1509,N_29854,N_29993);
xor UO_1510 (O_1510,N_29720,N_29956);
and UO_1511 (O_1511,N_29963,N_29913);
and UO_1512 (O_1512,N_29983,N_29931);
nand UO_1513 (O_1513,N_29769,N_29850);
nor UO_1514 (O_1514,N_29960,N_29863);
nand UO_1515 (O_1515,N_29890,N_29870);
xor UO_1516 (O_1516,N_29979,N_29861);
and UO_1517 (O_1517,N_29971,N_29919);
nor UO_1518 (O_1518,N_29773,N_29946);
nor UO_1519 (O_1519,N_29922,N_29802);
nor UO_1520 (O_1520,N_29896,N_29718);
and UO_1521 (O_1521,N_29860,N_29870);
nand UO_1522 (O_1522,N_29740,N_29726);
nand UO_1523 (O_1523,N_29999,N_29738);
and UO_1524 (O_1524,N_29775,N_29825);
xor UO_1525 (O_1525,N_29867,N_29713);
and UO_1526 (O_1526,N_29831,N_29822);
xnor UO_1527 (O_1527,N_29892,N_29738);
or UO_1528 (O_1528,N_29858,N_29837);
nor UO_1529 (O_1529,N_29918,N_29819);
or UO_1530 (O_1530,N_29754,N_29728);
nor UO_1531 (O_1531,N_29850,N_29714);
and UO_1532 (O_1532,N_29992,N_29831);
nand UO_1533 (O_1533,N_29739,N_29745);
nand UO_1534 (O_1534,N_29941,N_29794);
nand UO_1535 (O_1535,N_29850,N_29932);
nand UO_1536 (O_1536,N_29784,N_29707);
nand UO_1537 (O_1537,N_29961,N_29967);
xor UO_1538 (O_1538,N_29733,N_29952);
and UO_1539 (O_1539,N_29958,N_29896);
nand UO_1540 (O_1540,N_29785,N_29725);
or UO_1541 (O_1541,N_29977,N_29863);
nand UO_1542 (O_1542,N_29966,N_29962);
and UO_1543 (O_1543,N_29753,N_29981);
nor UO_1544 (O_1544,N_29941,N_29724);
nor UO_1545 (O_1545,N_29843,N_29951);
xnor UO_1546 (O_1546,N_29858,N_29806);
nand UO_1547 (O_1547,N_29700,N_29745);
nand UO_1548 (O_1548,N_29909,N_29838);
and UO_1549 (O_1549,N_29710,N_29912);
or UO_1550 (O_1550,N_29734,N_29716);
nor UO_1551 (O_1551,N_29847,N_29908);
or UO_1552 (O_1552,N_29779,N_29820);
nand UO_1553 (O_1553,N_29763,N_29933);
nand UO_1554 (O_1554,N_29703,N_29989);
xnor UO_1555 (O_1555,N_29974,N_29745);
or UO_1556 (O_1556,N_29882,N_29991);
nor UO_1557 (O_1557,N_29703,N_29890);
or UO_1558 (O_1558,N_29884,N_29858);
or UO_1559 (O_1559,N_29865,N_29871);
nor UO_1560 (O_1560,N_29845,N_29776);
xor UO_1561 (O_1561,N_29802,N_29910);
and UO_1562 (O_1562,N_29810,N_29989);
nand UO_1563 (O_1563,N_29896,N_29770);
nand UO_1564 (O_1564,N_29823,N_29815);
and UO_1565 (O_1565,N_29935,N_29723);
or UO_1566 (O_1566,N_29903,N_29730);
nand UO_1567 (O_1567,N_29932,N_29961);
nand UO_1568 (O_1568,N_29897,N_29983);
nor UO_1569 (O_1569,N_29768,N_29716);
nand UO_1570 (O_1570,N_29832,N_29997);
or UO_1571 (O_1571,N_29982,N_29736);
or UO_1572 (O_1572,N_29923,N_29702);
and UO_1573 (O_1573,N_29774,N_29905);
nor UO_1574 (O_1574,N_29778,N_29812);
or UO_1575 (O_1575,N_29892,N_29860);
nand UO_1576 (O_1576,N_29855,N_29711);
nor UO_1577 (O_1577,N_29716,N_29845);
nor UO_1578 (O_1578,N_29899,N_29719);
xor UO_1579 (O_1579,N_29771,N_29920);
or UO_1580 (O_1580,N_29897,N_29734);
nor UO_1581 (O_1581,N_29734,N_29812);
or UO_1582 (O_1582,N_29902,N_29993);
and UO_1583 (O_1583,N_29986,N_29894);
or UO_1584 (O_1584,N_29982,N_29990);
nor UO_1585 (O_1585,N_29740,N_29909);
and UO_1586 (O_1586,N_29798,N_29730);
xor UO_1587 (O_1587,N_29732,N_29924);
nor UO_1588 (O_1588,N_29783,N_29980);
and UO_1589 (O_1589,N_29735,N_29783);
or UO_1590 (O_1590,N_29777,N_29731);
or UO_1591 (O_1591,N_29871,N_29972);
xor UO_1592 (O_1592,N_29875,N_29900);
nor UO_1593 (O_1593,N_29770,N_29861);
xnor UO_1594 (O_1594,N_29716,N_29925);
and UO_1595 (O_1595,N_29844,N_29719);
nand UO_1596 (O_1596,N_29977,N_29992);
nor UO_1597 (O_1597,N_29857,N_29896);
nor UO_1598 (O_1598,N_29844,N_29833);
nor UO_1599 (O_1599,N_29816,N_29727);
nor UO_1600 (O_1600,N_29916,N_29890);
nand UO_1601 (O_1601,N_29983,N_29796);
nand UO_1602 (O_1602,N_29868,N_29876);
nand UO_1603 (O_1603,N_29746,N_29700);
xor UO_1604 (O_1604,N_29789,N_29724);
or UO_1605 (O_1605,N_29852,N_29769);
nand UO_1606 (O_1606,N_29921,N_29889);
and UO_1607 (O_1607,N_29919,N_29842);
nand UO_1608 (O_1608,N_29834,N_29915);
nor UO_1609 (O_1609,N_29841,N_29843);
xnor UO_1610 (O_1610,N_29858,N_29893);
and UO_1611 (O_1611,N_29737,N_29915);
nand UO_1612 (O_1612,N_29868,N_29904);
nand UO_1613 (O_1613,N_29793,N_29919);
or UO_1614 (O_1614,N_29932,N_29986);
and UO_1615 (O_1615,N_29984,N_29784);
nand UO_1616 (O_1616,N_29802,N_29895);
and UO_1617 (O_1617,N_29820,N_29757);
nand UO_1618 (O_1618,N_29911,N_29876);
xor UO_1619 (O_1619,N_29711,N_29779);
nand UO_1620 (O_1620,N_29979,N_29754);
and UO_1621 (O_1621,N_29875,N_29970);
xnor UO_1622 (O_1622,N_29888,N_29891);
or UO_1623 (O_1623,N_29903,N_29737);
xnor UO_1624 (O_1624,N_29791,N_29908);
or UO_1625 (O_1625,N_29961,N_29780);
and UO_1626 (O_1626,N_29918,N_29960);
and UO_1627 (O_1627,N_29862,N_29944);
and UO_1628 (O_1628,N_29905,N_29958);
nor UO_1629 (O_1629,N_29748,N_29863);
nor UO_1630 (O_1630,N_29721,N_29933);
nand UO_1631 (O_1631,N_29831,N_29792);
xnor UO_1632 (O_1632,N_29805,N_29853);
nand UO_1633 (O_1633,N_29765,N_29998);
and UO_1634 (O_1634,N_29713,N_29943);
and UO_1635 (O_1635,N_29965,N_29762);
or UO_1636 (O_1636,N_29847,N_29768);
nand UO_1637 (O_1637,N_29881,N_29999);
and UO_1638 (O_1638,N_29808,N_29956);
nor UO_1639 (O_1639,N_29884,N_29932);
or UO_1640 (O_1640,N_29912,N_29995);
nand UO_1641 (O_1641,N_29713,N_29980);
nand UO_1642 (O_1642,N_29972,N_29801);
nor UO_1643 (O_1643,N_29700,N_29850);
xor UO_1644 (O_1644,N_29829,N_29719);
or UO_1645 (O_1645,N_29856,N_29774);
nor UO_1646 (O_1646,N_29987,N_29925);
or UO_1647 (O_1647,N_29781,N_29952);
xor UO_1648 (O_1648,N_29789,N_29759);
and UO_1649 (O_1649,N_29866,N_29974);
or UO_1650 (O_1650,N_29757,N_29742);
and UO_1651 (O_1651,N_29708,N_29783);
nand UO_1652 (O_1652,N_29772,N_29791);
and UO_1653 (O_1653,N_29716,N_29813);
and UO_1654 (O_1654,N_29935,N_29974);
nand UO_1655 (O_1655,N_29857,N_29972);
xnor UO_1656 (O_1656,N_29854,N_29776);
xnor UO_1657 (O_1657,N_29709,N_29791);
or UO_1658 (O_1658,N_29807,N_29847);
nor UO_1659 (O_1659,N_29823,N_29822);
and UO_1660 (O_1660,N_29963,N_29926);
nand UO_1661 (O_1661,N_29893,N_29830);
nor UO_1662 (O_1662,N_29897,N_29802);
nor UO_1663 (O_1663,N_29803,N_29734);
nor UO_1664 (O_1664,N_29972,N_29804);
nor UO_1665 (O_1665,N_29823,N_29805);
or UO_1666 (O_1666,N_29734,N_29916);
or UO_1667 (O_1667,N_29845,N_29972);
and UO_1668 (O_1668,N_29951,N_29981);
and UO_1669 (O_1669,N_29986,N_29979);
or UO_1670 (O_1670,N_29767,N_29840);
nand UO_1671 (O_1671,N_29923,N_29714);
nor UO_1672 (O_1672,N_29935,N_29925);
and UO_1673 (O_1673,N_29931,N_29901);
nand UO_1674 (O_1674,N_29951,N_29945);
xor UO_1675 (O_1675,N_29910,N_29782);
nand UO_1676 (O_1676,N_29937,N_29977);
or UO_1677 (O_1677,N_29950,N_29804);
xor UO_1678 (O_1678,N_29705,N_29807);
nand UO_1679 (O_1679,N_29721,N_29791);
or UO_1680 (O_1680,N_29978,N_29895);
nand UO_1681 (O_1681,N_29852,N_29727);
nor UO_1682 (O_1682,N_29974,N_29920);
and UO_1683 (O_1683,N_29852,N_29706);
or UO_1684 (O_1684,N_29838,N_29750);
nand UO_1685 (O_1685,N_29937,N_29721);
and UO_1686 (O_1686,N_29723,N_29815);
and UO_1687 (O_1687,N_29966,N_29793);
nand UO_1688 (O_1688,N_29767,N_29871);
nor UO_1689 (O_1689,N_29723,N_29910);
and UO_1690 (O_1690,N_29785,N_29820);
or UO_1691 (O_1691,N_29968,N_29914);
or UO_1692 (O_1692,N_29952,N_29940);
nand UO_1693 (O_1693,N_29991,N_29883);
xor UO_1694 (O_1694,N_29992,N_29954);
xnor UO_1695 (O_1695,N_29931,N_29967);
xnor UO_1696 (O_1696,N_29885,N_29788);
and UO_1697 (O_1697,N_29725,N_29872);
and UO_1698 (O_1698,N_29953,N_29824);
xor UO_1699 (O_1699,N_29980,N_29933);
and UO_1700 (O_1700,N_29845,N_29865);
nand UO_1701 (O_1701,N_29964,N_29849);
and UO_1702 (O_1702,N_29925,N_29767);
nor UO_1703 (O_1703,N_29735,N_29806);
and UO_1704 (O_1704,N_29924,N_29936);
xor UO_1705 (O_1705,N_29847,N_29985);
xor UO_1706 (O_1706,N_29831,N_29746);
xnor UO_1707 (O_1707,N_29848,N_29923);
and UO_1708 (O_1708,N_29959,N_29940);
nor UO_1709 (O_1709,N_29705,N_29854);
nand UO_1710 (O_1710,N_29776,N_29819);
nand UO_1711 (O_1711,N_29755,N_29827);
or UO_1712 (O_1712,N_29807,N_29700);
xnor UO_1713 (O_1713,N_29747,N_29970);
xnor UO_1714 (O_1714,N_29848,N_29797);
or UO_1715 (O_1715,N_29871,N_29738);
and UO_1716 (O_1716,N_29961,N_29868);
xnor UO_1717 (O_1717,N_29952,N_29901);
xor UO_1718 (O_1718,N_29722,N_29840);
xor UO_1719 (O_1719,N_29997,N_29716);
nor UO_1720 (O_1720,N_29825,N_29713);
and UO_1721 (O_1721,N_29743,N_29728);
and UO_1722 (O_1722,N_29810,N_29724);
nand UO_1723 (O_1723,N_29805,N_29907);
and UO_1724 (O_1724,N_29821,N_29973);
and UO_1725 (O_1725,N_29942,N_29794);
nor UO_1726 (O_1726,N_29964,N_29772);
and UO_1727 (O_1727,N_29969,N_29742);
and UO_1728 (O_1728,N_29947,N_29939);
nand UO_1729 (O_1729,N_29811,N_29922);
xnor UO_1730 (O_1730,N_29708,N_29807);
nand UO_1731 (O_1731,N_29907,N_29780);
nand UO_1732 (O_1732,N_29809,N_29759);
or UO_1733 (O_1733,N_29774,N_29880);
and UO_1734 (O_1734,N_29865,N_29743);
nand UO_1735 (O_1735,N_29706,N_29891);
xnor UO_1736 (O_1736,N_29889,N_29948);
xor UO_1737 (O_1737,N_29731,N_29808);
or UO_1738 (O_1738,N_29988,N_29888);
nor UO_1739 (O_1739,N_29717,N_29808);
nand UO_1740 (O_1740,N_29901,N_29853);
and UO_1741 (O_1741,N_29780,N_29822);
and UO_1742 (O_1742,N_29829,N_29827);
or UO_1743 (O_1743,N_29842,N_29835);
nor UO_1744 (O_1744,N_29887,N_29845);
nor UO_1745 (O_1745,N_29921,N_29827);
and UO_1746 (O_1746,N_29830,N_29878);
xor UO_1747 (O_1747,N_29726,N_29969);
xnor UO_1748 (O_1748,N_29793,N_29819);
or UO_1749 (O_1749,N_29800,N_29920);
nor UO_1750 (O_1750,N_29732,N_29934);
nand UO_1751 (O_1751,N_29915,N_29924);
nand UO_1752 (O_1752,N_29929,N_29877);
nor UO_1753 (O_1753,N_29918,N_29928);
or UO_1754 (O_1754,N_29823,N_29909);
or UO_1755 (O_1755,N_29784,N_29938);
xor UO_1756 (O_1756,N_29913,N_29802);
or UO_1757 (O_1757,N_29873,N_29700);
nor UO_1758 (O_1758,N_29779,N_29710);
xor UO_1759 (O_1759,N_29915,N_29789);
xor UO_1760 (O_1760,N_29715,N_29921);
nand UO_1761 (O_1761,N_29789,N_29731);
or UO_1762 (O_1762,N_29798,N_29750);
xnor UO_1763 (O_1763,N_29981,N_29716);
nand UO_1764 (O_1764,N_29759,N_29742);
xor UO_1765 (O_1765,N_29861,N_29884);
nand UO_1766 (O_1766,N_29913,N_29839);
and UO_1767 (O_1767,N_29899,N_29702);
nor UO_1768 (O_1768,N_29728,N_29801);
and UO_1769 (O_1769,N_29900,N_29888);
or UO_1770 (O_1770,N_29991,N_29869);
or UO_1771 (O_1771,N_29899,N_29970);
and UO_1772 (O_1772,N_29850,N_29937);
or UO_1773 (O_1773,N_29780,N_29983);
nor UO_1774 (O_1774,N_29837,N_29994);
nand UO_1775 (O_1775,N_29885,N_29972);
nor UO_1776 (O_1776,N_29804,N_29758);
nor UO_1777 (O_1777,N_29946,N_29863);
nand UO_1778 (O_1778,N_29708,N_29789);
xor UO_1779 (O_1779,N_29920,N_29721);
and UO_1780 (O_1780,N_29946,N_29723);
and UO_1781 (O_1781,N_29701,N_29975);
xnor UO_1782 (O_1782,N_29934,N_29920);
xnor UO_1783 (O_1783,N_29903,N_29879);
xor UO_1784 (O_1784,N_29840,N_29795);
nand UO_1785 (O_1785,N_29866,N_29835);
nor UO_1786 (O_1786,N_29969,N_29794);
or UO_1787 (O_1787,N_29916,N_29809);
or UO_1788 (O_1788,N_29938,N_29826);
nor UO_1789 (O_1789,N_29844,N_29862);
and UO_1790 (O_1790,N_29899,N_29898);
xnor UO_1791 (O_1791,N_29943,N_29816);
xnor UO_1792 (O_1792,N_29925,N_29966);
nand UO_1793 (O_1793,N_29806,N_29972);
nor UO_1794 (O_1794,N_29858,N_29984);
xnor UO_1795 (O_1795,N_29878,N_29953);
nor UO_1796 (O_1796,N_29962,N_29755);
or UO_1797 (O_1797,N_29740,N_29750);
nor UO_1798 (O_1798,N_29788,N_29961);
nor UO_1799 (O_1799,N_29959,N_29819);
xnor UO_1800 (O_1800,N_29894,N_29863);
or UO_1801 (O_1801,N_29866,N_29746);
and UO_1802 (O_1802,N_29960,N_29785);
and UO_1803 (O_1803,N_29927,N_29856);
and UO_1804 (O_1804,N_29908,N_29845);
nor UO_1805 (O_1805,N_29907,N_29810);
nor UO_1806 (O_1806,N_29968,N_29931);
nand UO_1807 (O_1807,N_29760,N_29952);
and UO_1808 (O_1808,N_29920,N_29985);
or UO_1809 (O_1809,N_29866,N_29775);
nor UO_1810 (O_1810,N_29926,N_29856);
xnor UO_1811 (O_1811,N_29791,N_29883);
nand UO_1812 (O_1812,N_29807,N_29752);
or UO_1813 (O_1813,N_29753,N_29774);
xnor UO_1814 (O_1814,N_29983,N_29768);
xnor UO_1815 (O_1815,N_29875,N_29880);
xor UO_1816 (O_1816,N_29785,N_29792);
nor UO_1817 (O_1817,N_29812,N_29850);
xnor UO_1818 (O_1818,N_29806,N_29792);
xnor UO_1819 (O_1819,N_29857,N_29978);
xor UO_1820 (O_1820,N_29951,N_29838);
and UO_1821 (O_1821,N_29799,N_29896);
xnor UO_1822 (O_1822,N_29858,N_29736);
xor UO_1823 (O_1823,N_29917,N_29836);
and UO_1824 (O_1824,N_29720,N_29761);
nor UO_1825 (O_1825,N_29805,N_29708);
or UO_1826 (O_1826,N_29845,N_29870);
xor UO_1827 (O_1827,N_29801,N_29894);
or UO_1828 (O_1828,N_29934,N_29881);
xor UO_1829 (O_1829,N_29878,N_29827);
and UO_1830 (O_1830,N_29853,N_29762);
nor UO_1831 (O_1831,N_29934,N_29851);
and UO_1832 (O_1832,N_29861,N_29950);
or UO_1833 (O_1833,N_29776,N_29824);
or UO_1834 (O_1834,N_29894,N_29767);
or UO_1835 (O_1835,N_29777,N_29749);
nor UO_1836 (O_1836,N_29835,N_29768);
or UO_1837 (O_1837,N_29810,N_29880);
nor UO_1838 (O_1838,N_29713,N_29953);
nor UO_1839 (O_1839,N_29917,N_29974);
nor UO_1840 (O_1840,N_29877,N_29707);
nand UO_1841 (O_1841,N_29746,N_29868);
or UO_1842 (O_1842,N_29867,N_29986);
xor UO_1843 (O_1843,N_29934,N_29705);
xnor UO_1844 (O_1844,N_29952,N_29884);
xnor UO_1845 (O_1845,N_29851,N_29951);
xnor UO_1846 (O_1846,N_29876,N_29909);
or UO_1847 (O_1847,N_29978,N_29948);
and UO_1848 (O_1848,N_29864,N_29760);
xnor UO_1849 (O_1849,N_29736,N_29848);
nand UO_1850 (O_1850,N_29900,N_29981);
xnor UO_1851 (O_1851,N_29867,N_29843);
nor UO_1852 (O_1852,N_29738,N_29846);
nand UO_1853 (O_1853,N_29773,N_29975);
nand UO_1854 (O_1854,N_29946,N_29772);
xnor UO_1855 (O_1855,N_29711,N_29713);
nand UO_1856 (O_1856,N_29773,N_29728);
and UO_1857 (O_1857,N_29744,N_29836);
xnor UO_1858 (O_1858,N_29712,N_29784);
nand UO_1859 (O_1859,N_29717,N_29713);
nand UO_1860 (O_1860,N_29971,N_29810);
nand UO_1861 (O_1861,N_29967,N_29907);
nand UO_1862 (O_1862,N_29908,N_29834);
or UO_1863 (O_1863,N_29829,N_29921);
xnor UO_1864 (O_1864,N_29975,N_29996);
and UO_1865 (O_1865,N_29871,N_29791);
nor UO_1866 (O_1866,N_29769,N_29903);
xor UO_1867 (O_1867,N_29873,N_29994);
and UO_1868 (O_1868,N_29978,N_29892);
nor UO_1869 (O_1869,N_29852,N_29940);
and UO_1870 (O_1870,N_29806,N_29758);
or UO_1871 (O_1871,N_29930,N_29858);
xnor UO_1872 (O_1872,N_29793,N_29706);
xnor UO_1873 (O_1873,N_29721,N_29982);
and UO_1874 (O_1874,N_29939,N_29782);
nor UO_1875 (O_1875,N_29929,N_29965);
nor UO_1876 (O_1876,N_29917,N_29765);
xnor UO_1877 (O_1877,N_29955,N_29741);
or UO_1878 (O_1878,N_29811,N_29939);
nand UO_1879 (O_1879,N_29726,N_29873);
nor UO_1880 (O_1880,N_29952,N_29870);
xor UO_1881 (O_1881,N_29975,N_29881);
xor UO_1882 (O_1882,N_29921,N_29824);
nor UO_1883 (O_1883,N_29895,N_29747);
nor UO_1884 (O_1884,N_29764,N_29768);
nor UO_1885 (O_1885,N_29862,N_29719);
xnor UO_1886 (O_1886,N_29894,N_29755);
or UO_1887 (O_1887,N_29836,N_29996);
or UO_1888 (O_1888,N_29815,N_29811);
or UO_1889 (O_1889,N_29979,N_29940);
xnor UO_1890 (O_1890,N_29807,N_29714);
nand UO_1891 (O_1891,N_29775,N_29757);
or UO_1892 (O_1892,N_29925,N_29908);
nand UO_1893 (O_1893,N_29843,N_29800);
nand UO_1894 (O_1894,N_29981,N_29710);
nand UO_1895 (O_1895,N_29745,N_29991);
xnor UO_1896 (O_1896,N_29862,N_29920);
xor UO_1897 (O_1897,N_29713,N_29945);
xor UO_1898 (O_1898,N_29931,N_29724);
nand UO_1899 (O_1899,N_29867,N_29887);
nor UO_1900 (O_1900,N_29923,N_29775);
xnor UO_1901 (O_1901,N_29724,N_29725);
nand UO_1902 (O_1902,N_29777,N_29870);
nor UO_1903 (O_1903,N_29848,N_29776);
xor UO_1904 (O_1904,N_29753,N_29821);
and UO_1905 (O_1905,N_29779,N_29962);
nor UO_1906 (O_1906,N_29997,N_29885);
and UO_1907 (O_1907,N_29982,N_29771);
or UO_1908 (O_1908,N_29731,N_29787);
nor UO_1909 (O_1909,N_29870,N_29937);
xor UO_1910 (O_1910,N_29754,N_29707);
xor UO_1911 (O_1911,N_29825,N_29994);
nor UO_1912 (O_1912,N_29959,N_29788);
nand UO_1913 (O_1913,N_29930,N_29898);
nand UO_1914 (O_1914,N_29986,N_29984);
and UO_1915 (O_1915,N_29744,N_29903);
or UO_1916 (O_1916,N_29700,N_29960);
and UO_1917 (O_1917,N_29952,N_29817);
and UO_1918 (O_1918,N_29742,N_29962);
and UO_1919 (O_1919,N_29996,N_29776);
nor UO_1920 (O_1920,N_29916,N_29933);
and UO_1921 (O_1921,N_29762,N_29844);
or UO_1922 (O_1922,N_29852,N_29884);
nand UO_1923 (O_1923,N_29909,N_29834);
nor UO_1924 (O_1924,N_29989,N_29808);
nor UO_1925 (O_1925,N_29911,N_29860);
and UO_1926 (O_1926,N_29807,N_29846);
and UO_1927 (O_1927,N_29795,N_29778);
xor UO_1928 (O_1928,N_29988,N_29958);
and UO_1929 (O_1929,N_29762,N_29893);
or UO_1930 (O_1930,N_29949,N_29876);
nor UO_1931 (O_1931,N_29862,N_29801);
or UO_1932 (O_1932,N_29841,N_29990);
nor UO_1933 (O_1933,N_29843,N_29870);
xnor UO_1934 (O_1934,N_29702,N_29758);
xor UO_1935 (O_1935,N_29925,N_29849);
nor UO_1936 (O_1936,N_29813,N_29872);
xor UO_1937 (O_1937,N_29792,N_29929);
nand UO_1938 (O_1938,N_29761,N_29947);
xnor UO_1939 (O_1939,N_29762,N_29946);
and UO_1940 (O_1940,N_29782,N_29855);
nor UO_1941 (O_1941,N_29860,N_29720);
or UO_1942 (O_1942,N_29848,N_29983);
and UO_1943 (O_1943,N_29817,N_29736);
nand UO_1944 (O_1944,N_29831,N_29811);
and UO_1945 (O_1945,N_29834,N_29956);
nand UO_1946 (O_1946,N_29887,N_29884);
nor UO_1947 (O_1947,N_29767,N_29736);
xor UO_1948 (O_1948,N_29758,N_29876);
nand UO_1949 (O_1949,N_29888,N_29954);
nand UO_1950 (O_1950,N_29750,N_29957);
nand UO_1951 (O_1951,N_29964,N_29957);
and UO_1952 (O_1952,N_29871,N_29915);
nor UO_1953 (O_1953,N_29873,N_29925);
or UO_1954 (O_1954,N_29923,N_29760);
nor UO_1955 (O_1955,N_29733,N_29971);
xor UO_1956 (O_1956,N_29705,N_29790);
or UO_1957 (O_1957,N_29812,N_29760);
xor UO_1958 (O_1958,N_29799,N_29843);
or UO_1959 (O_1959,N_29717,N_29750);
and UO_1960 (O_1960,N_29719,N_29715);
nand UO_1961 (O_1961,N_29800,N_29794);
and UO_1962 (O_1962,N_29771,N_29836);
nand UO_1963 (O_1963,N_29918,N_29835);
nand UO_1964 (O_1964,N_29947,N_29742);
and UO_1965 (O_1965,N_29838,N_29942);
nand UO_1966 (O_1966,N_29989,N_29725);
and UO_1967 (O_1967,N_29702,N_29992);
nand UO_1968 (O_1968,N_29950,N_29970);
and UO_1969 (O_1969,N_29888,N_29701);
or UO_1970 (O_1970,N_29869,N_29777);
and UO_1971 (O_1971,N_29842,N_29951);
nor UO_1972 (O_1972,N_29869,N_29930);
xnor UO_1973 (O_1973,N_29934,N_29702);
and UO_1974 (O_1974,N_29872,N_29845);
or UO_1975 (O_1975,N_29760,N_29799);
or UO_1976 (O_1976,N_29856,N_29949);
or UO_1977 (O_1977,N_29932,N_29775);
or UO_1978 (O_1978,N_29877,N_29940);
and UO_1979 (O_1979,N_29928,N_29771);
nor UO_1980 (O_1980,N_29824,N_29811);
nand UO_1981 (O_1981,N_29950,N_29871);
or UO_1982 (O_1982,N_29844,N_29941);
and UO_1983 (O_1983,N_29927,N_29813);
nor UO_1984 (O_1984,N_29731,N_29971);
xnor UO_1985 (O_1985,N_29788,N_29746);
nand UO_1986 (O_1986,N_29980,N_29768);
or UO_1987 (O_1987,N_29893,N_29740);
nand UO_1988 (O_1988,N_29884,N_29919);
xnor UO_1989 (O_1989,N_29883,N_29948);
and UO_1990 (O_1990,N_29942,N_29978);
nand UO_1991 (O_1991,N_29915,N_29853);
and UO_1992 (O_1992,N_29790,N_29806);
xnor UO_1993 (O_1993,N_29843,N_29946);
or UO_1994 (O_1994,N_29900,N_29759);
nand UO_1995 (O_1995,N_29996,N_29748);
nor UO_1996 (O_1996,N_29940,N_29880);
or UO_1997 (O_1997,N_29747,N_29796);
nand UO_1998 (O_1998,N_29781,N_29944);
or UO_1999 (O_1999,N_29758,N_29981);
xnor UO_2000 (O_2000,N_29793,N_29797);
nand UO_2001 (O_2001,N_29736,N_29865);
nand UO_2002 (O_2002,N_29723,N_29940);
and UO_2003 (O_2003,N_29834,N_29965);
nand UO_2004 (O_2004,N_29924,N_29805);
nor UO_2005 (O_2005,N_29930,N_29813);
or UO_2006 (O_2006,N_29746,N_29879);
nor UO_2007 (O_2007,N_29996,N_29955);
xor UO_2008 (O_2008,N_29709,N_29924);
nor UO_2009 (O_2009,N_29737,N_29863);
nand UO_2010 (O_2010,N_29935,N_29758);
nor UO_2011 (O_2011,N_29934,N_29740);
nand UO_2012 (O_2012,N_29922,N_29733);
nor UO_2013 (O_2013,N_29759,N_29919);
xnor UO_2014 (O_2014,N_29849,N_29998);
or UO_2015 (O_2015,N_29763,N_29970);
nand UO_2016 (O_2016,N_29929,N_29810);
nor UO_2017 (O_2017,N_29755,N_29817);
nand UO_2018 (O_2018,N_29887,N_29911);
nor UO_2019 (O_2019,N_29881,N_29727);
xor UO_2020 (O_2020,N_29931,N_29781);
and UO_2021 (O_2021,N_29950,N_29806);
or UO_2022 (O_2022,N_29808,N_29848);
and UO_2023 (O_2023,N_29971,N_29857);
nor UO_2024 (O_2024,N_29736,N_29998);
nor UO_2025 (O_2025,N_29813,N_29721);
nand UO_2026 (O_2026,N_29790,N_29920);
nor UO_2027 (O_2027,N_29826,N_29927);
nor UO_2028 (O_2028,N_29727,N_29963);
or UO_2029 (O_2029,N_29734,N_29978);
nand UO_2030 (O_2030,N_29891,N_29912);
or UO_2031 (O_2031,N_29706,N_29867);
or UO_2032 (O_2032,N_29809,N_29749);
nand UO_2033 (O_2033,N_29957,N_29943);
and UO_2034 (O_2034,N_29704,N_29992);
xor UO_2035 (O_2035,N_29852,N_29962);
and UO_2036 (O_2036,N_29705,N_29745);
xor UO_2037 (O_2037,N_29820,N_29925);
or UO_2038 (O_2038,N_29806,N_29862);
nor UO_2039 (O_2039,N_29916,N_29720);
xnor UO_2040 (O_2040,N_29976,N_29786);
nand UO_2041 (O_2041,N_29991,N_29707);
xor UO_2042 (O_2042,N_29808,N_29736);
or UO_2043 (O_2043,N_29900,N_29824);
nor UO_2044 (O_2044,N_29811,N_29758);
nand UO_2045 (O_2045,N_29808,N_29751);
xnor UO_2046 (O_2046,N_29794,N_29952);
and UO_2047 (O_2047,N_29734,N_29713);
or UO_2048 (O_2048,N_29828,N_29767);
nand UO_2049 (O_2049,N_29970,N_29745);
xnor UO_2050 (O_2050,N_29896,N_29824);
and UO_2051 (O_2051,N_29785,N_29816);
xnor UO_2052 (O_2052,N_29705,N_29997);
xnor UO_2053 (O_2053,N_29962,N_29805);
nand UO_2054 (O_2054,N_29777,N_29790);
xnor UO_2055 (O_2055,N_29883,N_29876);
nand UO_2056 (O_2056,N_29778,N_29940);
and UO_2057 (O_2057,N_29862,N_29864);
nor UO_2058 (O_2058,N_29726,N_29850);
nor UO_2059 (O_2059,N_29814,N_29772);
or UO_2060 (O_2060,N_29947,N_29700);
or UO_2061 (O_2061,N_29708,N_29878);
or UO_2062 (O_2062,N_29828,N_29961);
nand UO_2063 (O_2063,N_29834,N_29871);
nor UO_2064 (O_2064,N_29952,N_29978);
nand UO_2065 (O_2065,N_29789,N_29752);
nand UO_2066 (O_2066,N_29958,N_29901);
nand UO_2067 (O_2067,N_29886,N_29722);
xor UO_2068 (O_2068,N_29771,N_29858);
nor UO_2069 (O_2069,N_29947,N_29918);
or UO_2070 (O_2070,N_29820,N_29905);
nand UO_2071 (O_2071,N_29862,N_29765);
nor UO_2072 (O_2072,N_29930,N_29783);
and UO_2073 (O_2073,N_29912,N_29933);
xnor UO_2074 (O_2074,N_29759,N_29796);
or UO_2075 (O_2075,N_29887,N_29725);
or UO_2076 (O_2076,N_29750,N_29988);
and UO_2077 (O_2077,N_29946,N_29811);
and UO_2078 (O_2078,N_29858,N_29917);
xor UO_2079 (O_2079,N_29765,N_29734);
nand UO_2080 (O_2080,N_29987,N_29890);
xor UO_2081 (O_2081,N_29976,N_29776);
and UO_2082 (O_2082,N_29979,N_29700);
or UO_2083 (O_2083,N_29744,N_29844);
nand UO_2084 (O_2084,N_29983,N_29830);
xnor UO_2085 (O_2085,N_29760,N_29969);
nand UO_2086 (O_2086,N_29744,N_29868);
and UO_2087 (O_2087,N_29789,N_29975);
or UO_2088 (O_2088,N_29955,N_29870);
and UO_2089 (O_2089,N_29788,N_29773);
nand UO_2090 (O_2090,N_29967,N_29733);
and UO_2091 (O_2091,N_29993,N_29966);
nor UO_2092 (O_2092,N_29843,N_29997);
or UO_2093 (O_2093,N_29926,N_29745);
and UO_2094 (O_2094,N_29763,N_29811);
nor UO_2095 (O_2095,N_29702,N_29967);
nor UO_2096 (O_2096,N_29871,N_29716);
xnor UO_2097 (O_2097,N_29903,N_29742);
xnor UO_2098 (O_2098,N_29847,N_29719);
nor UO_2099 (O_2099,N_29881,N_29945);
and UO_2100 (O_2100,N_29853,N_29959);
xnor UO_2101 (O_2101,N_29807,N_29837);
nor UO_2102 (O_2102,N_29951,N_29808);
nand UO_2103 (O_2103,N_29910,N_29865);
nand UO_2104 (O_2104,N_29891,N_29750);
nand UO_2105 (O_2105,N_29726,N_29984);
nor UO_2106 (O_2106,N_29866,N_29881);
nand UO_2107 (O_2107,N_29902,N_29721);
or UO_2108 (O_2108,N_29985,N_29854);
xor UO_2109 (O_2109,N_29795,N_29759);
or UO_2110 (O_2110,N_29848,N_29918);
nor UO_2111 (O_2111,N_29977,N_29755);
and UO_2112 (O_2112,N_29917,N_29894);
xnor UO_2113 (O_2113,N_29969,N_29861);
or UO_2114 (O_2114,N_29727,N_29870);
xor UO_2115 (O_2115,N_29799,N_29831);
xnor UO_2116 (O_2116,N_29941,N_29963);
or UO_2117 (O_2117,N_29954,N_29890);
nor UO_2118 (O_2118,N_29721,N_29896);
xnor UO_2119 (O_2119,N_29701,N_29827);
nand UO_2120 (O_2120,N_29899,N_29850);
or UO_2121 (O_2121,N_29926,N_29714);
nand UO_2122 (O_2122,N_29982,N_29921);
nand UO_2123 (O_2123,N_29937,N_29817);
xor UO_2124 (O_2124,N_29905,N_29943);
nand UO_2125 (O_2125,N_29988,N_29998);
xor UO_2126 (O_2126,N_29748,N_29943);
and UO_2127 (O_2127,N_29998,N_29908);
and UO_2128 (O_2128,N_29713,N_29702);
xor UO_2129 (O_2129,N_29840,N_29859);
nand UO_2130 (O_2130,N_29777,N_29922);
or UO_2131 (O_2131,N_29979,N_29945);
or UO_2132 (O_2132,N_29952,N_29701);
or UO_2133 (O_2133,N_29901,N_29963);
nand UO_2134 (O_2134,N_29867,N_29769);
nand UO_2135 (O_2135,N_29950,N_29893);
xor UO_2136 (O_2136,N_29886,N_29706);
xor UO_2137 (O_2137,N_29782,N_29759);
or UO_2138 (O_2138,N_29900,N_29765);
or UO_2139 (O_2139,N_29919,N_29892);
nor UO_2140 (O_2140,N_29806,N_29846);
and UO_2141 (O_2141,N_29752,N_29718);
nor UO_2142 (O_2142,N_29832,N_29759);
nand UO_2143 (O_2143,N_29745,N_29848);
nand UO_2144 (O_2144,N_29796,N_29798);
or UO_2145 (O_2145,N_29908,N_29760);
nor UO_2146 (O_2146,N_29769,N_29724);
xnor UO_2147 (O_2147,N_29922,N_29912);
nor UO_2148 (O_2148,N_29733,N_29963);
or UO_2149 (O_2149,N_29989,N_29805);
and UO_2150 (O_2150,N_29930,N_29982);
xnor UO_2151 (O_2151,N_29723,N_29986);
or UO_2152 (O_2152,N_29826,N_29747);
xor UO_2153 (O_2153,N_29942,N_29784);
xnor UO_2154 (O_2154,N_29819,N_29916);
xnor UO_2155 (O_2155,N_29855,N_29971);
nand UO_2156 (O_2156,N_29993,N_29720);
nor UO_2157 (O_2157,N_29963,N_29979);
or UO_2158 (O_2158,N_29729,N_29766);
and UO_2159 (O_2159,N_29791,N_29858);
or UO_2160 (O_2160,N_29729,N_29898);
or UO_2161 (O_2161,N_29955,N_29964);
xnor UO_2162 (O_2162,N_29921,N_29788);
nand UO_2163 (O_2163,N_29877,N_29846);
or UO_2164 (O_2164,N_29906,N_29965);
nand UO_2165 (O_2165,N_29874,N_29909);
or UO_2166 (O_2166,N_29737,N_29938);
xor UO_2167 (O_2167,N_29802,N_29906);
nand UO_2168 (O_2168,N_29706,N_29976);
nor UO_2169 (O_2169,N_29881,N_29745);
xnor UO_2170 (O_2170,N_29765,N_29735);
and UO_2171 (O_2171,N_29708,N_29829);
nand UO_2172 (O_2172,N_29955,N_29787);
xnor UO_2173 (O_2173,N_29707,N_29728);
nor UO_2174 (O_2174,N_29866,N_29738);
xor UO_2175 (O_2175,N_29770,N_29974);
nor UO_2176 (O_2176,N_29753,N_29901);
and UO_2177 (O_2177,N_29806,N_29740);
and UO_2178 (O_2178,N_29986,N_29989);
xnor UO_2179 (O_2179,N_29792,N_29880);
nand UO_2180 (O_2180,N_29862,N_29755);
nor UO_2181 (O_2181,N_29898,N_29827);
xor UO_2182 (O_2182,N_29753,N_29885);
and UO_2183 (O_2183,N_29719,N_29951);
xor UO_2184 (O_2184,N_29925,N_29880);
and UO_2185 (O_2185,N_29921,N_29898);
or UO_2186 (O_2186,N_29786,N_29782);
xnor UO_2187 (O_2187,N_29971,N_29942);
xnor UO_2188 (O_2188,N_29845,N_29851);
or UO_2189 (O_2189,N_29842,N_29957);
xnor UO_2190 (O_2190,N_29929,N_29907);
and UO_2191 (O_2191,N_29826,N_29848);
xnor UO_2192 (O_2192,N_29927,N_29920);
or UO_2193 (O_2193,N_29839,N_29704);
xnor UO_2194 (O_2194,N_29759,N_29951);
and UO_2195 (O_2195,N_29865,N_29829);
nand UO_2196 (O_2196,N_29869,N_29810);
xnor UO_2197 (O_2197,N_29772,N_29931);
or UO_2198 (O_2198,N_29721,N_29764);
and UO_2199 (O_2199,N_29939,N_29942);
or UO_2200 (O_2200,N_29703,N_29892);
xor UO_2201 (O_2201,N_29709,N_29913);
and UO_2202 (O_2202,N_29879,N_29850);
nand UO_2203 (O_2203,N_29807,N_29838);
or UO_2204 (O_2204,N_29983,N_29870);
nor UO_2205 (O_2205,N_29809,N_29991);
or UO_2206 (O_2206,N_29747,N_29765);
and UO_2207 (O_2207,N_29789,N_29818);
nor UO_2208 (O_2208,N_29869,N_29796);
nor UO_2209 (O_2209,N_29933,N_29814);
nor UO_2210 (O_2210,N_29891,N_29851);
nor UO_2211 (O_2211,N_29854,N_29738);
nor UO_2212 (O_2212,N_29930,N_29906);
xor UO_2213 (O_2213,N_29885,N_29704);
nand UO_2214 (O_2214,N_29920,N_29780);
or UO_2215 (O_2215,N_29868,N_29720);
or UO_2216 (O_2216,N_29967,N_29759);
and UO_2217 (O_2217,N_29922,N_29834);
or UO_2218 (O_2218,N_29853,N_29900);
nor UO_2219 (O_2219,N_29963,N_29858);
or UO_2220 (O_2220,N_29869,N_29742);
and UO_2221 (O_2221,N_29966,N_29810);
xnor UO_2222 (O_2222,N_29753,N_29747);
xor UO_2223 (O_2223,N_29757,N_29815);
xnor UO_2224 (O_2224,N_29805,N_29901);
and UO_2225 (O_2225,N_29865,N_29904);
xor UO_2226 (O_2226,N_29795,N_29708);
and UO_2227 (O_2227,N_29702,N_29987);
nor UO_2228 (O_2228,N_29817,N_29808);
and UO_2229 (O_2229,N_29826,N_29862);
nand UO_2230 (O_2230,N_29851,N_29812);
nor UO_2231 (O_2231,N_29772,N_29824);
or UO_2232 (O_2232,N_29886,N_29935);
nor UO_2233 (O_2233,N_29974,N_29702);
and UO_2234 (O_2234,N_29984,N_29887);
nand UO_2235 (O_2235,N_29759,N_29771);
or UO_2236 (O_2236,N_29839,N_29884);
xor UO_2237 (O_2237,N_29999,N_29861);
nor UO_2238 (O_2238,N_29741,N_29895);
and UO_2239 (O_2239,N_29906,N_29812);
and UO_2240 (O_2240,N_29992,N_29943);
nand UO_2241 (O_2241,N_29714,N_29961);
and UO_2242 (O_2242,N_29826,N_29824);
nor UO_2243 (O_2243,N_29730,N_29989);
xor UO_2244 (O_2244,N_29833,N_29901);
or UO_2245 (O_2245,N_29982,N_29911);
nor UO_2246 (O_2246,N_29871,N_29870);
or UO_2247 (O_2247,N_29756,N_29951);
and UO_2248 (O_2248,N_29955,N_29941);
nor UO_2249 (O_2249,N_29994,N_29744);
or UO_2250 (O_2250,N_29771,N_29762);
xnor UO_2251 (O_2251,N_29825,N_29722);
nand UO_2252 (O_2252,N_29737,N_29807);
or UO_2253 (O_2253,N_29945,N_29709);
or UO_2254 (O_2254,N_29791,N_29735);
and UO_2255 (O_2255,N_29961,N_29709);
or UO_2256 (O_2256,N_29841,N_29753);
xnor UO_2257 (O_2257,N_29915,N_29722);
and UO_2258 (O_2258,N_29768,N_29986);
nor UO_2259 (O_2259,N_29835,N_29865);
nand UO_2260 (O_2260,N_29928,N_29711);
nor UO_2261 (O_2261,N_29939,N_29855);
nor UO_2262 (O_2262,N_29752,N_29991);
and UO_2263 (O_2263,N_29855,N_29868);
nand UO_2264 (O_2264,N_29835,N_29961);
xnor UO_2265 (O_2265,N_29782,N_29918);
and UO_2266 (O_2266,N_29887,N_29926);
nand UO_2267 (O_2267,N_29723,N_29872);
nand UO_2268 (O_2268,N_29857,N_29799);
nor UO_2269 (O_2269,N_29722,N_29783);
nor UO_2270 (O_2270,N_29777,N_29770);
and UO_2271 (O_2271,N_29947,N_29886);
or UO_2272 (O_2272,N_29798,N_29893);
nand UO_2273 (O_2273,N_29793,N_29932);
xnor UO_2274 (O_2274,N_29834,N_29819);
xor UO_2275 (O_2275,N_29937,N_29961);
nand UO_2276 (O_2276,N_29976,N_29965);
nand UO_2277 (O_2277,N_29885,N_29945);
and UO_2278 (O_2278,N_29780,N_29965);
and UO_2279 (O_2279,N_29776,N_29772);
nand UO_2280 (O_2280,N_29751,N_29836);
nor UO_2281 (O_2281,N_29977,N_29910);
nor UO_2282 (O_2282,N_29978,N_29815);
nor UO_2283 (O_2283,N_29840,N_29924);
and UO_2284 (O_2284,N_29883,N_29807);
or UO_2285 (O_2285,N_29768,N_29938);
and UO_2286 (O_2286,N_29790,N_29723);
nand UO_2287 (O_2287,N_29708,N_29892);
and UO_2288 (O_2288,N_29880,N_29965);
xor UO_2289 (O_2289,N_29712,N_29791);
nor UO_2290 (O_2290,N_29894,N_29808);
and UO_2291 (O_2291,N_29825,N_29931);
xnor UO_2292 (O_2292,N_29813,N_29839);
or UO_2293 (O_2293,N_29958,N_29797);
nand UO_2294 (O_2294,N_29912,N_29863);
xnor UO_2295 (O_2295,N_29968,N_29822);
nand UO_2296 (O_2296,N_29778,N_29805);
and UO_2297 (O_2297,N_29873,N_29908);
xor UO_2298 (O_2298,N_29768,N_29952);
nor UO_2299 (O_2299,N_29843,N_29733);
or UO_2300 (O_2300,N_29761,N_29830);
nor UO_2301 (O_2301,N_29806,N_29827);
nor UO_2302 (O_2302,N_29955,N_29866);
nand UO_2303 (O_2303,N_29904,N_29908);
and UO_2304 (O_2304,N_29792,N_29778);
and UO_2305 (O_2305,N_29903,N_29819);
xor UO_2306 (O_2306,N_29944,N_29868);
or UO_2307 (O_2307,N_29864,N_29716);
nor UO_2308 (O_2308,N_29960,N_29867);
xnor UO_2309 (O_2309,N_29951,N_29829);
or UO_2310 (O_2310,N_29705,N_29751);
or UO_2311 (O_2311,N_29746,N_29718);
nand UO_2312 (O_2312,N_29967,N_29861);
nand UO_2313 (O_2313,N_29759,N_29703);
or UO_2314 (O_2314,N_29820,N_29834);
and UO_2315 (O_2315,N_29980,N_29927);
and UO_2316 (O_2316,N_29992,N_29925);
and UO_2317 (O_2317,N_29854,N_29808);
xor UO_2318 (O_2318,N_29776,N_29925);
and UO_2319 (O_2319,N_29934,N_29965);
nand UO_2320 (O_2320,N_29994,N_29738);
nand UO_2321 (O_2321,N_29956,N_29886);
xnor UO_2322 (O_2322,N_29884,N_29969);
nand UO_2323 (O_2323,N_29788,N_29710);
xor UO_2324 (O_2324,N_29713,N_29812);
nor UO_2325 (O_2325,N_29713,N_29924);
xnor UO_2326 (O_2326,N_29936,N_29902);
or UO_2327 (O_2327,N_29987,N_29933);
and UO_2328 (O_2328,N_29884,N_29797);
and UO_2329 (O_2329,N_29836,N_29736);
and UO_2330 (O_2330,N_29952,N_29893);
or UO_2331 (O_2331,N_29783,N_29990);
and UO_2332 (O_2332,N_29734,N_29876);
nand UO_2333 (O_2333,N_29976,N_29769);
nor UO_2334 (O_2334,N_29714,N_29849);
nor UO_2335 (O_2335,N_29918,N_29704);
nand UO_2336 (O_2336,N_29838,N_29798);
nand UO_2337 (O_2337,N_29796,N_29822);
nand UO_2338 (O_2338,N_29871,N_29826);
nand UO_2339 (O_2339,N_29711,N_29725);
or UO_2340 (O_2340,N_29940,N_29812);
or UO_2341 (O_2341,N_29819,N_29853);
nor UO_2342 (O_2342,N_29715,N_29778);
or UO_2343 (O_2343,N_29975,N_29715);
or UO_2344 (O_2344,N_29867,N_29756);
and UO_2345 (O_2345,N_29860,N_29844);
nor UO_2346 (O_2346,N_29752,N_29946);
or UO_2347 (O_2347,N_29752,N_29734);
and UO_2348 (O_2348,N_29703,N_29876);
or UO_2349 (O_2349,N_29863,N_29736);
nand UO_2350 (O_2350,N_29708,N_29750);
and UO_2351 (O_2351,N_29988,N_29937);
nand UO_2352 (O_2352,N_29997,N_29707);
and UO_2353 (O_2353,N_29752,N_29898);
and UO_2354 (O_2354,N_29866,N_29932);
and UO_2355 (O_2355,N_29773,N_29710);
and UO_2356 (O_2356,N_29987,N_29897);
and UO_2357 (O_2357,N_29741,N_29834);
and UO_2358 (O_2358,N_29991,N_29767);
xor UO_2359 (O_2359,N_29938,N_29839);
nor UO_2360 (O_2360,N_29830,N_29866);
and UO_2361 (O_2361,N_29921,N_29929);
and UO_2362 (O_2362,N_29906,N_29706);
xnor UO_2363 (O_2363,N_29943,N_29832);
xnor UO_2364 (O_2364,N_29962,N_29921);
and UO_2365 (O_2365,N_29989,N_29865);
xnor UO_2366 (O_2366,N_29808,N_29726);
xor UO_2367 (O_2367,N_29934,N_29823);
nor UO_2368 (O_2368,N_29896,N_29748);
and UO_2369 (O_2369,N_29752,N_29917);
and UO_2370 (O_2370,N_29825,N_29886);
nand UO_2371 (O_2371,N_29870,N_29755);
nor UO_2372 (O_2372,N_29870,N_29964);
xnor UO_2373 (O_2373,N_29748,N_29965);
and UO_2374 (O_2374,N_29782,N_29778);
and UO_2375 (O_2375,N_29933,N_29878);
xor UO_2376 (O_2376,N_29864,N_29881);
xor UO_2377 (O_2377,N_29930,N_29847);
xor UO_2378 (O_2378,N_29802,N_29810);
nand UO_2379 (O_2379,N_29917,N_29718);
nand UO_2380 (O_2380,N_29797,N_29804);
nor UO_2381 (O_2381,N_29822,N_29775);
nand UO_2382 (O_2382,N_29965,N_29758);
or UO_2383 (O_2383,N_29715,N_29783);
nor UO_2384 (O_2384,N_29960,N_29711);
or UO_2385 (O_2385,N_29817,N_29787);
xor UO_2386 (O_2386,N_29790,N_29952);
and UO_2387 (O_2387,N_29970,N_29905);
and UO_2388 (O_2388,N_29829,N_29894);
xnor UO_2389 (O_2389,N_29785,N_29803);
nand UO_2390 (O_2390,N_29902,N_29910);
xor UO_2391 (O_2391,N_29854,N_29865);
nor UO_2392 (O_2392,N_29900,N_29979);
and UO_2393 (O_2393,N_29987,N_29939);
or UO_2394 (O_2394,N_29811,N_29750);
nand UO_2395 (O_2395,N_29758,N_29734);
and UO_2396 (O_2396,N_29974,N_29898);
and UO_2397 (O_2397,N_29757,N_29983);
nor UO_2398 (O_2398,N_29804,N_29974);
nor UO_2399 (O_2399,N_29891,N_29709);
xnor UO_2400 (O_2400,N_29842,N_29849);
nor UO_2401 (O_2401,N_29867,N_29852);
or UO_2402 (O_2402,N_29911,N_29747);
or UO_2403 (O_2403,N_29997,N_29743);
nor UO_2404 (O_2404,N_29803,N_29814);
and UO_2405 (O_2405,N_29782,N_29821);
and UO_2406 (O_2406,N_29802,N_29894);
nand UO_2407 (O_2407,N_29722,N_29869);
xor UO_2408 (O_2408,N_29932,N_29865);
nand UO_2409 (O_2409,N_29815,N_29864);
nor UO_2410 (O_2410,N_29809,N_29832);
nor UO_2411 (O_2411,N_29971,N_29980);
or UO_2412 (O_2412,N_29965,N_29751);
or UO_2413 (O_2413,N_29922,N_29730);
xnor UO_2414 (O_2414,N_29743,N_29991);
nand UO_2415 (O_2415,N_29789,N_29872);
xnor UO_2416 (O_2416,N_29919,N_29934);
and UO_2417 (O_2417,N_29892,N_29815);
nand UO_2418 (O_2418,N_29977,N_29779);
nor UO_2419 (O_2419,N_29713,N_29964);
xor UO_2420 (O_2420,N_29717,N_29729);
nor UO_2421 (O_2421,N_29933,N_29813);
xor UO_2422 (O_2422,N_29824,N_29872);
and UO_2423 (O_2423,N_29897,N_29779);
nand UO_2424 (O_2424,N_29851,N_29770);
or UO_2425 (O_2425,N_29971,N_29865);
nor UO_2426 (O_2426,N_29801,N_29979);
and UO_2427 (O_2427,N_29965,N_29863);
nand UO_2428 (O_2428,N_29710,N_29714);
nand UO_2429 (O_2429,N_29764,N_29871);
or UO_2430 (O_2430,N_29929,N_29910);
nand UO_2431 (O_2431,N_29763,N_29983);
xor UO_2432 (O_2432,N_29993,N_29887);
xor UO_2433 (O_2433,N_29761,N_29942);
and UO_2434 (O_2434,N_29984,N_29893);
or UO_2435 (O_2435,N_29707,N_29999);
and UO_2436 (O_2436,N_29831,N_29707);
nor UO_2437 (O_2437,N_29796,N_29946);
or UO_2438 (O_2438,N_29877,N_29758);
or UO_2439 (O_2439,N_29861,N_29911);
or UO_2440 (O_2440,N_29702,N_29975);
nor UO_2441 (O_2441,N_29930,N_29796);
nor UO_2442 (O_2442,N_29763,N_29848);
nor UO_2443 (O_2443,N_29831,N_29712);
or UO_2444 (O_2444,N_29837,N_29815);
nor UO_2445 (O_2445,N_29771,N_29947);
nand UO_2446 (O_2446,N_29818,N_29920);
and UO_2447 (O_2447,N_29788,N_29703);
or UO_2448 (O_2448,N_29850,N_29859);
and UO_2449 (O_2449,N_29722,N_29908);
nor UO_2450 (O_2450,N_29876,N_29743);
or UO_2451 (O_2451,N_29855,N_29703);
or UO_2452 (O_2452,N_29739,N_29735);
nand UO_2453 (O_2453,N_29700,N_29983);
xor UO_2454 (O_2454,N_29971,N_29721);
nand UO_2455 (O_2455,N_29941,N_29983);
xor UO_2456 (O_2456,N_29750,N_29884);
xnor UO_2457 (O_2457,N_29809,N_29921);
or UO_2458 (O_2458,N_29815,N_29932);
nand UO_2459 (O_2459,N_29932,N_29708);
and UO_2460 (O_2460,N_29829,N_29838);
or UO_2461 (O_2461,N_29832,N_29726);
and UO_2462 (O_2462,N_29756,N_29786);
and UO_2463 (O_2463,N_29777,N_29920);
nand UO_2464 (O_2464,N_29898,N_29783);
xor UO_2465 (O_2465,N_29808,N_29906);
xor UO_2466 (O_2466,N_29904,N_29752);
xnor UO_2467 (O_2467,N_29834,N_29730);
and UO_2468 (O_2468,N_29702,N_29712);
nand UO_2469 (O_2469,N_29957,N_29776);
nand UO_2470 (O_2470,N_29977,N_29856);
nand UO_2471 (O_2471,N_29920,N_29723);
nand UO_2472 (O_2472,N_29709,N_29898);
or UO_2473 (O_2473,N_29967,N_29872);
and UO_2474 (O_2474,N_29836,N_29935);
or UO_2475 (O_2475,N_29885,N_29980);
or UO_2476 (O_2476,N_29896,N_29916);
and UO_2477 (O_2477,N_29773,N_29821);
xnor UO_2478 (O_2478,N_29955,N_29793);
and UO_2479 (O_2479,N_29908,N_29701);
and UO_2480 (O_2480,N_29911,N_29856);
and UO_2481 (O_2481,N_29751,N_29954);
nor UO_2482 (O_2482,N_29830,N_29997);
and UO_2483 (O_2483,N_29843,N_29988);
nand UO_2484 (O_2484,N_29993,N_29863);
nand UO_2485 (O_2485,N_29811,N_29935);
xnor UO_2486 (O_2486,N_29722,N_29791);
nand UO_2487 (O_2487,N_29963,N_29945);
xor UO_2488 (O_2488,N_29716,N_29775);
xnor UO_2489 (O_2489,N_29853,N_29946);
nand UO_2490 (O_2490,N_29882,N_29770);
xnor UO_2491 (O_2491,N_29750,N_29765);
nand UO_2492 (O_2492,N_29929,N_29876);
nand UO_2493 (O_2493,N_29857,N_29967);
xor UO_2494 (O_2494,N_29839,N_29984);
nand UO_2495 (O_2495,N_29985,N_29777);
and UO_2496 (O_2496,N_29790,N_29880);
or UO_2497 (O_2497,N_29772,N_29979);
or UO_2498 (O_2498,N_29910,N_29725);
nand UO_2499 (O_2499,N_29837,N_29956);
or UO_2500 (O_2500,N_29712,N_29984);
nor UO_2501 (O_2501,N_29973,N_29791);
nand UO_2502 (O_2502,N_29994,N_29966);
and UO_2503 (O_2503,N_29862,N_29970);
nor UO_2504 (O_2504,N_29893,N_29720);
nand UO_2505 (O_2505,N_29874,N_29981);
and UO_2506 (O_2506,N_29804,N_29749);
and UO_2507 (O_2507,N_29821,N_29930);
nand UO_2508 (O_2508,N_29899,N_29903);
nand UO_2509 (O_2509,N_29753,N_29748);
xor UO_2510 (O_2510,N_29713,N_29984);
or UO_2511 (O_2511,N_29853,N_29962);
and UO_2512 (O_2512,N_29706,N_29981);
or UO_2513 (O_2513,N_29954,N_29922);
xor UO_2514 (O_2514,N_29928,N_29872);
and UO_2515 (O_2515,N_29952,N_29914);
or UO_2516 (O_2516,N_29741,N_29904);
nor UO_2517 (O_2517,N_29996,N_29872);
nand UO_2518 (O_2518,N_29852,N_29873);
and UO_2519 (O_2519,N_29837,N_29809);
or UO_2520 (O_2520,N_29948,N_29922);
or UO_2521 (O_2521,N_29721,N_29783);
and UO_2522 (O_2522,N_29747,N_29706);
or UO_2523 (O_2523,N_29922,N_29886);
or UO_2524 (O_2524,N_29774,N_29768);
nor UO_2525 (O_2525,N_29812,N_29955);
nor UO_2526 (O_2526,N_29849,N_29823);
xnor UO_2527 (O_2527,N_29830,N_29961);
and UO_2528 (O_2528,N_29863,N_29821);
xor UO_2529 (O_2529,N_29753,N_29888);
or UO_2530 (O_2530,N_29719,N_29825);
nand UO_2531 (O_2531,N_29767,N_29796);
xor UO_2532 (O_2532,N_29870,N_29976);
and UO_2533 (O_2533,N_29866,N_29754);
or UO_2534 (O_2534,N_29992,N_29963);
nor UO_2535 (O_2535,N_29742,N_29984);
or UO_2536 (O_2536,N_29734,N_29908);
and UO_2537 (O_2537,N_29858,N_29750);
xnor UO_2538 (O_2538,N_29983,N_29854);
nand UO_2539 (O_2539,N_29996,N_29945);
nor UO_2540 (O_2540,N_29978,N_29784);
or UO_2541 (O_2541,N_29800,N_29736);
xnor UO_2542 (O_2542,N_29895,N_29962);
nand UO_2543 (O_2543,N_29789,N_29792);
or UO_2544 (O_2544,N_29832,N_29860);
or UO_2545 (O_2545,N_29866,N_29914);
xnor UO_2546 (O_2546,N_29771,N_29981);
and UO_2547 (O_2547,N_29802,N_29869);
xnor UO_2548 (O_2548,N_29806,N_29746);
and UO_2549 (O_2549,N_29885,N_29896);
xor UO_2550 (O_2550,N_29726,N_29977);
nand UO_2551 (O_2551,N_29795,N_29838);
xor UO_2552 (O_2552,N_29730,N_29831);
or UO_2553 (O_2553,N_29761,N_29940);
nor UO_2554 (O_2554,N_29731,N_29828);
and UO_2555 (O_2555,N_29734,N_29863);
and UO_2556 (O_2556,N_29740,N_29825);
and UO_2557 (O_2557,N_29755,N_29722);
nand UO_2558 (O_2558,N_29782,N_29755);
nor UO_2559 (O_2559,N_29839,N_29883);
nor UO_2560 (O_2560,N_29828,N_29861);
nand UO_2561 (O_2561,N_29801,N_29986);
xnor UO_2562 (O_2562,N_29897,N_29959);
or UO_2563 (O_2563,N_29884,N_29881);
and UO_2564 (O_2564,N_29938,N_29985);
or UO_2565 (O_2565,N_29723,N_29874);
nor UO_2566 (O_2566,N_29705,N_29753);
nand UO_2567 (O_2567,N_29976,N_29853);
nand UO_2568 (O_2568,N_29920,N_29897);
nor UO_2569 (O_2569,N_29880,N_29865);
and UO_2570 (O_2570,N_29789,N_29798);
and UO_2571 (O_2571,N_29906,N_29797);
xor UO_2572 (O_2572,N_29978,N_29896);
or UO_2573 (O_2573,N_29820,N_29940);
and UO_2574 (O_2574,N_29846,N_29751);
and UO_2575 (O_2575,N_29832,N_29864);
and UO_2576 (O_2576,N_29709,N_29739);
nand UO_2577 (O_2577,N_29956,N_29802);
nor UO_2578 (O_2578,N_29940,N_29999);
nor UO_2579 (O_2579,N_29984,N_29985);
and UO_2580 (O_2580,N_29978,N_29930);
nand UO_2581 (O_2581,N_29860,N_29762);
nor UO_2582 (O_2582,N_29872,N_29764);
nand UO_2583 (O_2583,N_29813,N_29765);
nor UO_2584 (O_2584,N_29796,N_29923);
or UO_2585 (O_2585,N_29909,N_29924);
and UO_2586 (O_2586,N_29784,N_29948);
nand UO_2587 (O_2587,N_29714,N_29770);
or UO_2588 (O_2588,N_29986,N_29718);
nor UO_2589 (O_2589,N_29847,N_29938);
xor UO_2590 (O_2590,N_29956,N_29734);
xor UO_2591 (O_2591,N_29973,N_29727);
or UO_2592 (O_2592,N_29833,N_29712);
and UO_2593 (O_2593,N_29998,N_29821);
xnor UO_2594 (O_2594,N_29909,N_29739);
nand UO_2595 (O_2595,N_29709,N_29971);
and UO_2596 (O_2596,N_29752,N_29701);
nor UO_2597 (O_2597,N_29763,N_29796);
xnor UO_2598 (O_2598,N_29753,N_29759);
and UO_2599 (O_2599,N_29821,N_29847);
nor UO_2600 (O_2600,N_29818,N_29866);
nand UO_2601 (O_2601,N_29726,N_29773);
nand UO_2602 (O_2602,N_29844,N_29726);
xor UO_2603 (O_2603,N_29802,N_29759);
nor UO_2604 (O_2604,N_29801,N_29914);
xnor UO_2605 (O_2605,N_29980,N_29860);
nor UO_2606 (O_2606,N_29749,N_29870);
and UO_2607 (O_2607,N_29995,N_29969);
and UO_2608 (O_2608,N_29854,N_29851);
xnor UO_2609 (O_2609,N_29705,N_29754);
or UO_2610 (O_2610,N_29942,N_29969);
or UO_2611 (O_2611,N_29927,N_29855);
and UO_2612 (O_2612,N_29934,N_29809);
nand UO_2613 (O_2613,N_29739,N_29856);
and UO_2614 (O_2614,N_29839,N_29736);
and UO_2615 (O_2615,N_29745,N_29804);
or UO_2616 (O_2616,N_29882,N_29782);
nand UO_2617 (O_2617,N_29716,N_29987);
or UO_2618 (O_2618,N_29999,N_29822);
nor UO_2619 (O_2619,N_29742,N_29714);
and UO_2620 (O_2620,N_29793,N_29887);
and UO_2621 (O_2621,N_29999,N_29892);
or UO_2622 (O_2622,N_29886,N_29834);
and UO_2623 (O_2623,N_29890,N_29911);
nor UO_2624 (O_2624,N_29761,N_29831);
nor UO_2625 (O_2625,N_29732,N_29727);
or UO_2626 (O_2626,N_29866,N_29996);
or UO_2627 (O_2627,N_29828,N_29733);
nand UO_2628 (O_2628,N_29837,N_29898);
nand UO_2629 (O_2629,N_29745,N_29877);
xor UO_2630 (O_2630,N_29946,N_29797);
and UO_2631 (O_2631,N_29932,N_29929);
xor UO_2632 (O_2632,N_29785,N_29789);
nor UO_2633 (O_2633,N_29769,N_29804);
nand UO_2634 (O_2634,N_29922,N_29956);
nand UO_2635 (O_2635,N_29716,N_29950);
nand UO_2636 (O_2636,N_29772,N_29923);
nor UO_2637 (O_2637,N_29762,N_29953);
nand UO_2638 (O_2638,N_29905,N_29867);
xnor UO_2639 (O_2639,N_29990,N_29879);
nor UO_2640 (O_2640,N_29842,N_29929);
nand UO_2641 (O_2641,N_29959,N_29945);
or UO_2642 (O_2642,N_29885,N_29772);
or UO_2643 (O_2643,N_29828,N_29926);
nor UO_2644 (O_2644,N_29879,N_29906);
nor UO_2645 (O_2645,N_29899,N_29825);
nor UO_2646 (O_2646,N_29879,N_29809);
nor UO_2647 (O_2647,N_29927,N_29901);
or UO_2648 (O_2648,N_29860,N_29878);
and UO_2649 (O_2649,N_29845,N_29813);
or UO_2650 (O_2650,N_29892,N_29903);
xnor UO_2651 (O_2651,N_29831,N_29980);
or UO_2652 (O_2652,N_29884,N_29940);
nor UO_2653 (O_2653,N_29821,N_29967);
xnor UO_2654 (O_2654,N_29780,N_29716);
nand UO_2655 (O_2655,N_29804,N_29993);
or UO_2656 (O_2656,N_29850,N_29952);
xor UO_2657 (O_2657,N_29704,N_29930);
nor UO_2658 (O_2658,N_29822,N_29987);
nand UO_2659 (O_2659,N_29839,N_29851);
nor UO_2660 (O_2660,N_29835,N_29887);
nand UO_2661 (O_2661,N_29922,N_29971);
and UO_2662 (O_2662,N_29847,N_29996);
and UO_2663 (O_2663,N_29768,N_29936);
or UO_2664 (O_2664,N_29935,N_29963);
or UO_2665 (O_2665,N_29869,N_29798);
or UO_2666 (O_2666,N_29917,N_29946);
or UO_2667 (O_2667,N_29782,N_29756);
nor UO_2668 (O_2668,N_29802,N_29965);
or UO_2669 (O_2669,N_29788,N_29705);
xor UO_2670 (O_2670,N_29700,N_29988);
and UO_2671 (O_2671,N_29705,N_29912);
or UO_2672 (O_2672,N_29889,N_29859);
and UO_2673 (O_2673,N_29994,N_29901);
nand UO_2674 (O_2674,N_29704,N_29773);
or UO_2675 (O_2675,N_29836,N_29992);
or UO_2676 (O_2676,N_29819,N_29720);
xor UO_2677 (O_2677,N_29991,N_29971);
and UO_2678 (O_2678,N_29997,N_29900);
xnor UO_2679 (O_2679,N_29796,N_29874);
nand UO_2680 (O_2680,N_29993,N_29971);
nor UO_2681 (O_2681,N_29974,N_29950);
nand UO_2682 (O_2682,N_29714,N_29828);
or UO_2683 (O_2683,N_29819,N_29805);
and UO_2684 (O_2684,N_29771,N_29761);
and UO_2685 (O_2685,N_29811,N_29707);
or UO_2686 (O_2686,N_29901,N_29855);
and UO_2687 (O_2687,N_29749,N_29849);
xor UO_2688 (O_2688,N_29876,N_29795);
xnor UO_2689 (O_2689,N_29891,N_29720);
xnor UO_2690 (O_2690,N_29912,N_29866);
or UO_2691 (O_2691,N_29860,N_29943);
nand UO_2692 (O_2692,N_29910,N_29847);
nand UO_2693 (O_2693,N_29929,N_29903);
or UO_2694 (O_2694,N_29941,N_29818);
nand UO_2695 (O_2695,N_29930,N_29922);
and UO_2696 (O_2696,N_29894,N_29797);
nor UO_2697 (O_2697,N_29972,N_29999);
or UO_2698 (O_2698,N_29884,N_29944);
nor UO_2699 (O_2699,N_29859,N_29813);
xnor UO_2700 (O_2700,N_29715,N_29816);
and UO_2701 (O_2701,N_29876,N_29874);
xor UO_2702 (O_2702,N_29913,N_29706);
xor UO_2703 (O_2703,N_29961,N_29859);
and UO_2704 (O_2704,N_29860,N_29942);
xor UO_2705 (O_2705,N_29833,N_29715);
or UO_2706 (O_2706,N_29751,N_29733);
xor UO_2707 (O_2707,N_29831,N_29770);
and UO_2708 (O_2708,N_29940,N_29890);
nor UO_2709 (O_2709,N_29896,N_29735);
or UO_2710 (O_2710,N_29838,N_29982);
and UO_2711 (O_2711,N_29854,N_29859);
nor UO_2712 (O_2712,N_29874,N_29868);
nand UO_2713 (O_2713,N_29927,N_29874);
and UO_2714 (O_2714,N_29919,N_29935);
nor UO_2715 (O_2715,N_29906,N_29782);
and UO_2716 (O_2716,N_29762,N_29852);
xnor UO_2717 (O_2717,N_29895,N_29886);
xor UO_2718 (O_2718,N_29701,N_29884);
nand UO_2719 (O_2719,N_29834,N_29892);
xor UO_2720 (O_2720,N_29781,N_29716);
nor UO_2721 (O_2721,N_29905,N_29753);
nand UO_2722 (O_2722,N_29955,N_29851);
and UO_2723 (O_2723,N_29864,N_29722);
and UO_2724 (O_2724,N_29992,N_29850);
and UO_2725 (O_2725,N_29975,N_29948);
nor UO_2726 (O_2726,N_29818,N_29853);
xor UO_2727 (O_2727,N_29802,N_29872);
or UO_2728 (O_2728,N_29891,N_29970);
or UO_2729 (O_2729,N_29959,N_29910);
nand UO_2730 (O_2730,N_29759,N_29882);
xnor UO_2731 (O_2731,N_29936,N_29762);
nand UO_2732 (O_2732,N_29870,N_29958);
nand UO_2733 (O_2733,N_29700,N_29996);
nand UO_2734 (O_2734,N_29827,N_29705);
and UO_2735 (O_2735,N_29928,N_29754);
nor UO_2736 (O_2736,N_29900,N_29720);
and UO_2737 (O_2737,N_29996,N_29839);
nand UO_2738 (O_2738,N_29716,N_29928);
or UO_2739 (O_2739,N_29949,N_29765);
nand UO_2740 (O_2740,N_29859,N_29956);
or UO_2741 (O_2741,N_29788,N_29877);
or UO_2742 (O_2742,N_29934,N_29834);
xnor UO_2743 (O_2743,N_29769,N_29737);
or UO_2744 (O_2744,N_29701,N_29802);
nand UO_2745 (O_2745,N_29725,N_29806);
nand UO_2746 (O_2746,N_29866,N_29952);
or UO_2747 (O_2747,N_29809,N_29721);
xnor UO_2748 (O_2748,N_29729,N_29823);
nand UO_2749 (O_2749,N_29944,N_29760);
and UO_2750 (O_2750,N_29913,N_29885);
xor UO_2751 (O_2751,N_29866,N_29959);
and UO_2752 (O_2752,N_29968,N_29838);
nand UO_2753 (O_2753,N_29759,N_29988);
and UO_2754 (O_2754,N_29891,N_29922);
xor UO_2755 (O_2755,N_29704,N_29909);
or UO_2756 (O_2756,N_29915,N_29732);
nand UO_2757 (O_2757,N_29961,N_29996);
or UO_2758 (O_2758,N_29710,N_29846);
xor UO_2759 (O_2759,N_29980,N_29820);
nand UO_2760 (O_2760,N_29912,N_29913);
xor UO_2761 (O_2761,N_29866,N_29721);
or UO_2762 (O_2762,N_29978,N_29750);
xnor UO_2763 (O_2763,N_29938,N_29904);
and UO_2764 (O_2764,N_29726,N_29949);
nand UO_2765 (O_2765,N_29967,N_29750);
and UO_2766 (O_2766,N_29759,N_29811);
or UO_2767 (O_2767,N_29703,N_29953);
nand UO_2768 (O_2768,N_29957,N_29756);
nand UO_2769 (O_2769,N_29733,N_29861);
nand UO_2770 (O_2770,N_29828,N_29739);
or UO_2771 (O_2771,N_29833,N_29867);
and UO_2772 (O_2772,N_29827,N_29733);
nand UO_2773 (O_2773,N_29733,N_29988);
nor UO_2774 (O_2774,N_29704,N_29735);
or UO_2775 (O_2775,N_29957,N_29884);
nor UO_2776 (O_2776,N_29993,N_29942);
nand UO_2777 (O_2777,N_29966,N_29751);
nor UO_2778 (O_2778,N_29921,N_29927);
and UO_2779 (O_2779,N_29836,N_29886);
xnor UO_2780 (O_2780,N_29852,N_29713);
xor UO_2781 (O_2781,N_29936,N_29892);
nor UO_2782 (O_2782,N_29838,N_29754);
nor UO_2783 (O_2783,N_29932,N_29967);
xor UO_2784 (O_2784,N_29796,N_29831);
nand UO_2785 (O_2785,N_29842,N_29748);
nor UO_2786 (O_2786,N_29812,N_29834);
and UO_2787 (O_2787,N_29703,N_29846);
xor UO_2788 (O_2788,N_29863,N_29927);
nor UO_2789 (O_2789,N_29845,N_29761);
xnor UO_2790 (O_2790,N_29776,N_29909);
xor UO_2791 (O_2791,N_29717,N_29869);
nand UO_2792 (O_2792,N_29719,N_29753);
or UO_2793 (O_2793,N_29886,N_29713);
xor UO_2794 (O_2794,N_29976,N_29999);
nand UO_2795 (O_2795,N_29847,N_29881);
and UO_2796 (O_2796,N_29747,N_29835);
and UO_2797 (O_2797,N_29787,N_29745);
nor UO_2798 (O_2798,N_29875,N_29975);
and UO_2799 (O_2799,N_29942,N_29789);
nor UO_2800 (O_2800,N_29883,N_29841);
nand UO_2801 (O_2801,N_29747,N_29743);
nand UO_2802 (O_2802,N_29928,N_29827);
and UO_2803 (O_2803,N_29858,N_29847);
nand UO_2804 (O_2804,N_29880,N_29817);
and UO_2805 (O_2805,N_29801,N_29787);
or UO_2806 (O_2806,N_29835,N_29962);
nand UO_2807 (O_2807,N_29849,N_29753);
and UO_2808 (O_2808,N_29995,N_29836);
nand UO_2809 (O_2809,N_29892,N_29792);
nor UO_2810 (O_2810,N_29714,N_29775);
nor UO_2811 (O_2811,N_29774,N_29750);
nand UO_2812 (O_2812,N_29986,N_29956);
and UO_2813 (O_2813,N_29818,N_29781);
xnor UO_2814 (O_2814,N_29803,N_29906);
nand UO_2815 (O_2815,N_29910,N_29743);
and UO_2816 (O_2816,N_29877,N_29836);
nor UO_2817 (O_2817,N_29765,N_29819);
or UO_2818 (O_2818,N_29860,N_29901);
xnor UO_2819 (O_2819,N_29847,N_29988);
and UO_2820 (O_2820,N_29974,N_29947);
nor UO_2821 (O_2821,N_29922,N_29783);
or UO_2822 (O_2822,N_29725,N_29787);
nor UO_2823 (O_2823,N_29977,N_29704);
nand UO_2824 (O_2824,N_29806,N_29764);
and UO_2825 (O_2825,N_29752,N_29964);
or UO_2826 (O_2826,N_29799,N_29802);
and UO_2827 (O_2827,N_29809,N_29957);
or UO_2828 (O_2828,N_29829,N_29959);
xor UO_2829 (O_2829,N_29993,N_29938);
or UO_2830 (O_2830,N_29994,N_29890);
and UO_2831 (O_2831,N_29993,N_29835);
nor UO_2832 (O_2832,N_29851,N_29960);
or UO_2833 (O_2833,N_29931,N_29734);
nand UO_2834 (O_2834,N_29848,N_29862);
nand UO_2835 (O_2835,N_29874,N_29730);
nor UO_2836 (O_2836,N_29912,N_29883);
or UO_2837 (O_2837,N_29904,N_29916);
or UO_2838 (O_2838,N_29897,N_29725);
xor UO_2839 (O_2839,N_29714,N_29871);
or UO_2840 (O_2840,N_29811,N_29712);
nand UO_2841 (O_2841,N_29855,N_29951);
nor UO_2842 (O_2842,N_29860,N_29786);
and UO_2843 (O_2843,N_29752,N_29710);
xor UO_2844 (O_2844,N_29749,N_29876);
or UO_2845 (O_2845,N_29841,N_29772);
or UO_2846 (O_2846,N_29956,N_29952);
and UO_2847 (O_2847,N_29756,N_29868);
or UO_2848 (O_2848,N_29912,N_29769);
and UO_2849 (O_2849,N_29870,N_29822);
nor UO_2850 (O_2850,N_29701,N_29841);
nor UO_2851 (O_2851,N_29767,N_29844);
nand UO_2852 (O_2852,N_29846,N_29810);
nand UO_2853 (O_2853,N_29767,N_29920);
or UO_2854 (O_2854,N_29968,N_29771);
nand UO_2855 (O_2855,N_29769,N_29729);
or UO_2856 (O_2856,N_29988,N_29824);
or UO_2857 (O_2857,N_29881,N_29825);
or UO_2858 (O_2858,N_29814,N_29865);
xnor UO_2859 (O_2859,N_29813,N_29996);
nand UO_2860 (O_2860,N_29830,N_29804);
nand UO_2861 (O_2861,N_29827,N_29938);
nor UO_2862 (O_2862,N_29791,N_29889);
nand UO_2863 (O_2863,N_29857,N_29995);
nand UO_2864 (O_2864,N_29824,N_29791);
and UO_2865 (O_2865,N_29937,N_29960);
nand UO_2866 (O_2866,N_29854,N_29850);
nor UO_2867 (O_2867,N_29969,N_29773);
and UO_2868 (O_2868,N_29750,N_29983);
or UO_2869 (O_2869,N_29960,N_29870);
nand UO_2870 (O_2870,N_29882,N_29983);
and UO_2871 (O_2871,N_29901,N_29929);
or UO_2872 (O_2872,N_29956,N_29950);
nor UO_2873 (O_2873,N_29935,N_29732);
xnor UO_2874 (O_2874,N_29771,N_29924);
or UO_2875 (O_2875,N_29949,N_29715);
nand UO_2876 (O_2876,N_29832,N_29706);
nor UO_2877 (O_2877,N_29912,N_29965);
and UO_2878 (O_2878,N_29823,N_29752);
and UO_2879 (O_2879,N_29768,N_29871);
xor UO_2880 (O_2880,N_29797,N_29994);
and UO_2881 (O_2881,N_29753,N_29792);
xor UO_2882 (O_2882,N_29992,N_29828);
nor UO_2883 (O_2883,N_29953,N_29893);
and UO_2884 (O_2884,N_29991,N_29834);
and UO_2885 (O_2885,N_29734,N_29756);
xor UO_2886 (O_2886,N_29915,N_29912);
xnor UO_2887 (O_2887,N_29813,N_29775);
nand UO_2888 (O_2888,N_29961,N_29781);
nor UO_2889 (O_2889,N_29794,N_29737);
and UO_2890 (O_2890,N_29881,N_29749);
or UO_2891 (O_2891,N_29806,N_29904);
xor UO_2892 (O_2892,N_29909,N_29729);
nor UO_2893 (O_2893,N_29915,N_29953);
nor UO_2894 (O_2894,N_29938,N_29924);
xor UO_2895 (O_2895,N_29757,N_29985);
nand UO_2896 (O_2896,N_29983,N_29893);
nor UO_2897 (O_2897,N_29937,N_29761);
or UO_2898 (O_2898,N_29993,N_29792);
nand UO_2899 (O_2899,N_29855,N_29937);
xnor UO_2900 (O_2900,N_29878,N_29844);
and UO_2901 (O_2901,N_29863,N_29909);
nor UO_2902 (O_2902,N_29976,N_29728);
and UO_2903 (O_2903,N_29908,N_29774);
nor UO_2904 (O_2904,N_29758,N_29746);
nand UO_2905 (O_2905,N_29827,N_29900);
nor UO_2906 (O_2906,N_29821,N_29834);
nor UO_2907 (O_2907,N_29896,N_29872);
xnor UO_2908 (O_2908,N_29766,N_29972);
or UO_2909 (O_2909,N_29998,N_29769);
xnor UO_2910 (O_2910,N_29961,N_29920);
xnor UO_2911 (O_2911,N_29857,N_29920);
nand UO_2912 (O_2912,N_29703,N_29795);
nor UO_2913 (O_2913,N_29847,N_29779);
and UO_2914 (O_2914,N_29782,N_29764);
or UO_2915 (O_2915,N_29967,N_29779);
nand UO_2916 (O_2916,N_29998,N_29913);
xor UO_2917 (O_2917,N_29926,N_29725);
nand UO_2918 (O_2918,N_29899,N_29841);
nor UO_2919 (O_2919,N_29933,N_29705);
nor UO_2920 (O_2920,N_29919,N_29869);
nand UO_2921 (O_2921,N_29822,N_29827);
nand UO_2922 (O_2922,N_29920,N_29948);
nor UO_2923 (O_2923,N_29909,N_29749);
nor UO_2924 (O_2924,N_29822,N_29860);
or UO_2925 (O_2925,N_29729,N_29815);
and UO_2926 (O_2926,N_29949,N_29731);
xnor UO_2927 (O_2927,N_29951,N_29760);
xor UO_2928 (O_2928,N_29777,N_29916);
or UO_2929 (O_2929,N_29738,N_29907);
and UO_2930 (O_2930,N_29894,N_29901);
and UO_2931 (O_2931,N_29767,N_29993);
or UO_2932 (O_2932,N_29794,N_29998);
and UO_2933 (O_2933,N_29839,N_29776);
nand UO_2934 (O_2934,N_29911,N_29979);
xor UO_2935 (O_2935,N_29776,N_29733);
nand UO_2936 (O_2936,N_29949,N_29819);
xnor UO_2937 (O_2937,N_29957,N_29910);
nor UO_2938 (O_2938,N_29942,N_29974);
nand UO_2939 (O_2939,N_29769,N_29985);
nand UO_2940 (O_2940,N_29969,N_29863);
or UO_2941 (O_2941,N_29926,N_29862);
and UO_2942 (O_2942,N_29982,N_29739);
nand UO_2943 (O_2943,N_29936,N_29795);
and UO_2944 (O_2944,N_29734,N_29986);
nor UO_2945 (O_2945,N_29722,N_29776);
nor UO_2946 (O_2946,N_29800,N_29866);
xor UO_2947 (O_2947,N_29977,N_29906);
xor UO_2948 (O_2948,N_29947,N_29838);
or UO_2949 (O_2949,N_29960,N_29907);
and UO_2950 (O_2950,N_29751,N_29936);
nand UO_2951 (O_2951,N_29817,N_29822);
or UO_2952 (O_2952,N_29830,N_29762);
xnor UO_2953 (O_2953,N_29783,N_29753);
and UO_2954 (O_2954,N_29994,N_29804);
nand UO_2955 (O_2955,N_29915,N_29832);
and UO_2956 (O_2956,N_29744,N_29945);
or UO_2957 (O_2957,N_29814,N_29951);
and UO_2958 (O_2958,N_29844,N_29990);
or UO_2959 (O_2959,N_29858,N_29816);
and UO_2960 (O_2960,N_29832,N_29932);
nor UO_2961 (O_2961,N_29918,N_29829);
nor UO_2962 (O_2962,N_29734,N_29865);
or UO_2963 (O_2963,N_29988,N_29726);
or UO_2964 (O_2964,N_29811,N_29912);
or UO_2965 (O_2965,N_29848,N_29881);
and UO_2966 (O_2966,N_29775,N_29998);
nor UO_2967 (O_2967,N_29810,N_29986);
and UO_2968 (O_2968,N_29795,N_29723);
xnor UO_2969 (O_2969,N_29723,N_29744);
nor UO_2970 (O_2970,N_29961,N_29851);
and UO_2971 (O_2971,N_29818,N_29700);
and UO_2972 (O_2972,N_29996,N_29734);
nor UO_2973 (O_2973,N_29765,N_29893);
or UO_2974 (O_2974,N_29732,N_29942);
nor UO_2975 (O_2975,N_29708,N_29759);
or UO_2976 (O_2976,N_29878,N_29753);
nor UO_2977 (O_2977,N_29994,N_29817);
or UO_2978 (O_2978,N_29702,N_29740);
or UO_2979 (O_2979,N_29802,N_29924);
nand UO_2980 (O_2980,N_29989,N_29953);
nor UO_2981 (O_2981,N_29766,N_29965);
or UO_2982 (O_2982,N_29998,N_29847);
nor UO_2983 (O_2983,N_29992,N_29951);
xnor UO_2984 (O_2984,N_29726,N_29954);
and UO_2985 (O_2985,N_29731,N_29880);
or UO_2986 (O_2986,N_29770,N_29725);
and UO_2987 (O_2987,N_29787,N_29850);
nor UO_2988 (O_2988,N_29961,N_29821);
xor UO_2989 (O_2989,N_29835,N_29728);
and UO_2990 (O_2990,N_29843,N_29923);
nand UO_2991 (O_2991,N_29976,N_29969);
and UO_2992 (O_2992,N_29951,N_29733);
or UO_2993 (O_2993,N_29817,N_29995);
nor UO_2994 (O_2994,N_29923,N_29842);
nand UO_2995 (O_2995,N_29826,N_29738);
or UO_2996 (O_2996,N_29758,N_29745);
and UO_2997 (O_2997,N_29931,N_29810);
and UO_2998 (O_2998,N_29705,N_29722);
nor UO_2999 (O_2999,N_29843,N_29904);
nand UO_3000 (O_3000,N_29827,N_29885);
nor UO_3001 (O_3001,N_29907,N_29916);
or UO_3002 (O_3002,N_29973,N_29839);
nor UO_3003 (O_3003,N_29871,N_29787);
and UO_3004 (O_3004,N_29832,N_29907);
or UO_3005 (O_3005,N_29865,N_29849);
or UO_3006 (O_3006,N_29814,N_29927);
nand UO_3007 (O_3007,N_29932,N_29764);
xor UO_3008 (O_3008,N_29919,N_29700);
and UO_3009 (O_3009,N_29864,N_29719);
nand UO_3010 (O_3010,N_29993,N_29981);
nor UO_3011 (O_3011,N_29706,N_29781);
and UO_3012 (O_3012,N_29877,N_29725);
and UO_3013 (O_3013,N_29755,N_29737);
xor UO_3014 (O_3014,N_29869,N_29764);
nor UO_3015 (O_3015,N_29905,N_29949);
nor UO_3016 (O_3016,N_29877,N_29817);
nand UO_3017 (O_3017,N_29728,N_29803);
nor UO_3018 (O_3018,N_29865,N_29737);
xor UO_3019 (O_3019,N_29771,N_29819);
nor UO_3020 (O_3020,N_29959,N_29801);
and UO_3021 (O_3021,N_29744,N_29884);
and UO_3022 (O_3022,N_29801,N_29910);
nand UO_3023 (O_3023,N_29994,N_29870);
or UO_3024 (O_3024,N_29917,N_29846);
and UO_3025 (O_3025,N_29950,N_29988);
nand UO_3026 (O_3026,N_29745,N_29887);
or UO_3027 (O_3027,N_29848,N_29755);
xor UO_3028 (O_3028,N_29910,N_29998);
and UO_3029 (O_3029,N_29702,N_29993);
and UO_3030 (O_3030,N_29971,N_29858);
nor UO_3031 (O_3031,N_29759,N_29887);
and UO_3032 (O_3032,N_29806,N_29870);
and UO_3033 (O_3033,N_29966,N_29762);
and UO_3034 (O_3034,N_29942,N_29944);
nand UO_3035 (O_3035,N_29838,N_29707);
or UO_3036 (O_3036,N_29856,N_29921);
or UO_3037 (O_3037,N_29955,N_29705);
nor UO_3038 (O_3038,N_29751,N_29925);
nand UO_3039 (O_3039,N_29711,N_29910);
xnor UO_3040 (O_3040,N_29885,N_29910);
nor UO_3041 (O_3041,N_29948,N_29716);
and UO_3042 (O_3042,N_29754,N_29977);
or UO_3043 (O_3043,N_29875,N_29850);
and UO_3044 (O_3044,N_29966,N_29724);
or UO_3045 (O_3045,N_29901,N_29706);
and UO_3046 (O_3046,N_29953,N_29991);
xor UO_3047 (O_3047,N_29865,N_29972);
nor UO_3048 (O_3048,N_29799,N_29937);
xnor UO_3049 (O_3049,N_29986,N_29905);
nor UO_3050 (O_3050,N_29863,N_29743);
nor UO_3051 (O_3051,N_29881,N_29762);
xnor UO_3052 (O_3052,N_29892,N_29935);
nand UO_3053 (O_3053,N_29792,N_29712);
or UO_3054 (O_3054,N_29734,N_29700);
nand UO_3055 (O_3055,N_29719,N_29995);
xor UO_3056 (O_3056,N_29918,N_29992);
xnor UO_3057 (O_3057,N_29823,N_29892);
and UO_3058 (O_3058,N_29796,N_29907);
nor UO_3059 (O_3059,N_29914,N_29970);
nand UO_3060 (O_3060,N_29749,N_29987);
nand UO_3061 (O_3061,N_29848,N_29962);
nor UO_3062 (O_3062,N_29843,N_29920);
xor UO_3063 (O_3063,N_29758,N_29780);
or UO_3064 (O_3064,N_29726,N_29734);
xnor UO_3065 (O_3065,N_29919,N_29983);
xnor UO_3066 (O_3066,N_29887,N_29813);
nor UO_3067 (O_3067,N_29910,N_29840);
nor UO_3068 (O_3068,N_29973,N_29873);
and UO_3069 (O_3069,N_29774,N_29983);
nand UO_3070 (O_3070,N_29945,N_29777);
nor UO_3071 (O_3071,N_29731,N_29761);
nand UO_3072 (O_3072,N_29916,N_29801);
or UO_3073 (O_3073,N_29770,N_29836);
xnor UO_3074 (O_3074,N_29824,N_29930);
or UO_3075 (O_3075,N_29901,N_29953);
and UO_3076 (O_3076,N_29864,N_29946);
nor UO_3077 (O_3077,N_29887,N_29820);
xor UO_3078 (O_3078,N_29866,N_29973);
xnor UO_3079 (O_3079,N_29840,N_29817);
nand UO_3080 (O_3080,N_29735,N_29943);
nand UO_3081 (O_3081,N_29937,N_29981);
or UO_3082 (O_3082,N_29863,N_29865);
and UO_3083 (O_3083,N_29993,N_29805);
nor UO_3084 (O_3084,N_29726,N_29935);
nand UO_3085 (O_3085,N_29930,N_29935);
nor UO_3086 (O_3086,N_29870,N_29798);
or UO_3087 (O_3087,N_29879,N_29823);
nand UO_3088 (O_3088,N_29725,N_29983);
and UO_3089 (O_3089,N_29945,N_29868);
or UO_3090 (O_3090,N_29959,N_29838);
or UO_3091 (O_3091,N_29818,N_29807);
nand UO_3092 (O_3092,N_29969,N_29772);
or UO_3093 (O_3093,N_29722,N_29981);
or UO_3094 (O_3094,N_29896,N_29732);
nor UO_3095 (O_3095,N_29784,N_29878);
nor UO_3096 (O_3096,N_29719,N_29950);
and UO_3097 (O_3097,N_29973,N_29943);
nor UO_3098 (O_3098,N_29807,N_29787);
or UO_3099 (O_3099,N_29732,N_29825);
xor UO_3100 (O_3100,N_29712,N_29925);
nor UO_3101 (O_3101,N_29987,N_29904);
xnor UO_3102 (O_3102,N_29879,N_29857);
or UO_3103 (O_3103,N_29906,N_29911);
or UO_3104 (O_3104,N_29928,N_29993);
and UO_3105 (O_3105,N_29828,N_29793);
and UO_3106 (O_3106,N_29909,N_29792);
or UO_3107 (O_3107,N_29810,N_29809);
nand UO_3108 (O_3108,N_29771,N_29766);
or UO_3109 (O_3109,N_29945,N_29892);
or UO_3110 (O_3110,N_29751,N_29782);
and UO_3111 (O_3111,N_29742,N_29827);
nand UO_3112 (O_3112,N_29707,N_29765);
xnor UO_3113 (O_3113,N_29969,N_29854);
and UO_3114 (O_3114,N_29869,N_29885);
nand UO_3115 (O_3115,N_29821,N_29966);
and UO_3116 (O_3116,N_29858,N_29982);
xor UO_3117 (O_3117,N_29950,N_29731);
nor UO_3118 (O_3118,N_29955,N_29828);
nor UO_3119 (O_3119,N_29884,N_29767);
and UO_3120 (O_3120,N_29759,N_29888);
nor UO_3121 (O_3121,N_29768,N_29955);
xor UO_3122 (O_3122,N_29891,N_29941);
nand UO_3123 (O_3123,N_29925,N_29936);
and UO_3124 (O_3124,N_29740,N_29774);
xnor UO_3125 (O_3125,N_29976,N_29716);
or UO_3126 (O_3126,N_29825,N_29943);
nand UO_3127 (O_3127,N_29974,N_29889);
nor UO_3128 (O_3128,N_29719,N_29954);
and UO_3129 (O_3129,N_29903,N_29727);
and UO_3130 (O_3130,N_29807,N_29724);
xor UO_3131 (O_3131,N_29823,N_29799);
xor UO_3132 (O_3132,N_29984,N_29843);
nor UO_3133 (O_3133,N_29759,N_29749);
and UO_3134 (O_3134,N_29851,N_29964);
nor UO_3135 (O_3135,N_29777,N_29780);
nor UO_3136 (O_3136,N_29770,N_29793);
nand UO_3137 (O_3137,N_29958,N_29861);
and UO_3138 (O_3138,N_29708,N_29706);
and UO_3139 (O_3139,N_29733,N_29702);
xor UO_3140 (O_3140,N_29824,N_29813);
nor UO_3141 (O_3141,N_29929,N_29859);
xor UO_3142 (O_3142,N_29909,N_29962);
xor UO_3143 (O_3143,N_29912,N_29784);
nand UO_3144 (O_3144,N_29811,N_29869);
or UO_3145 (O_3145,N_29802,N_29868);
or UO_3146 (O_3146,N_29840,N_29868);
or UO_3147 (O_3147,N_29866,N_29794);
xor UO_3148 (O_3148,N_29953,N_29994);
nand UO_3149 (O_3149,N_29723,N_29801);
nand UO_3150 (O_3150,N_29785,N_29954);
nor UO_3151 (O_3151,N_29790,N_29912);
nand UO_3152 (O_3152,N_29787,N_29987);
nand UO_3153 (O_3153,N_29767,N_29703);
nand UO_3154 (O_3154,N_29892,N_29793);
nor UO_3155 (O_3155,N_29810,N_29805);
nor UO_3156 (O_3156,N_29946,N_29953);
xor UO_3157 (O_3157,N_29865,N_29778);
and UO_3158 (O_3158,N_29954,N_29788);
or UO_3159 (O_3159,N_29976,N_29879);
and UO_3160 (O_3160,N_29921,N_29847);
or UO_3161 (O_3161,N_29944,N_29812);
xnor UO_3162 (O_3162,N_29862,N_29713);
nand UO_3163 (O_3163,N_29806,N_29910);
nor UO_3164 (O_3164,N_29702,N_29919);
nand UO_3165 (O_3165,N_29797,N_29800);
xor UO_3166 (O_3166,N_29913,N_29710);
xnor UO_3167 (O_3167,N_29932,N_29889);
nor UO_3168 (O_3168,N_29813,N_29740);
nor UO_3169 (O_3169,N_29933,N_29782);
and UO_3170 (O_3170,N_29855,N_29936);
nor UO_3171 (O_3171,N_29928,N_29934);
or UO_3172 (O_3172,N_29986,N_29703);
nor UO_3173 (O_3173,N_29943,N_29897);
or UO_3174 (O_3174,N_29780,N_29796);
nand UO_3175 (O_3175,N_29857,N_29911);
nand UO_3176 (O_3176,N_29758,N_29852);
nand UO_3177 (O_3177,N_29967,N_29928);
xnor UO_3178 (O_3178,N_29799,N_29888);
or UO_3179 (O_3179,N_29948,N_29878);
nor UO_3180 (O_3180,N_29717,N_29973);
xor UO_3181 (O_3181,N_29718,N_29954);
nor UO_3182 (O_3182,N_29876,N_29780);
nand UO_3183 (O_3183,N_29784,N_29777);
or UO_3184 (O_3184,N_29974,N_29979);
and UO_3185 (O_3185,N_29896,N_29984);
nand UO_3186 (O_3186,N_29763,N_29806);
or UO_3187 (O_3187,N_29825,N_29723);
and UO_3188 (O_3188,N_29742,N_29872);
nand UO_3189 (O_3189,N_29711,N_29868);
and UO_3190 (O_3190,N_29773,N_29818);
and UO_3191 (O_3191,N_29780,N_29955);
xor UO_3192 (O_3192,N_29801,N_29927);
xnor UO_3193 (O_3193,N_29944,N_29956);
and UO_3194 (O_3194,N_29835,N_29855);
and UO_3195 (O_3195,N_29863,N_29751);
nor UO_3196 (O_3196,N_29707,N_29814);
xor UO_3197 (O_3197,N_29872,N_29720);
nor UO_3198 (O_3198,N_29971,N_29724);
or UO_3199 (O_3199,N_29705,N_29890);
and UO_3200 (O_3200,N_29809,N_29949);
xnor UO_3201 (O_3201,N_29994,N_29928);
or UO_3202 (O_3202,N_29749,N_29836);
and UO_3203 (O_3203,N_29995,N_29838);
nor UO_3204 (O_3204,N_29949,N_29842);
xor UO_3205 (O_3205,N_29708,N_29967);
nor UO_3206 (O_3206,N_29726,N_29729);
xnor UO_3207 (O_3207,N_29865,N_29777);
nor UO_3208 (O_3208,N_29925,N_29781);
nand UO_3209 (O_3209,N_29861,N_29883);
and UO_3210 (O_3210,N_29937,N_29940);
and UO_3211 (O_3211,N_29703,N_29975);
nor UO_3212 (O_3212,N_29711,N_29818);
nor UO_3213 (O_3213,N_29782,N_29898);
or UO_3214 (O_3214,N_29807,N_29795);
and UO_3215 (O_3215,N_29765,N_29808);
nand UO_3216 (O_3216,N_29926,N_29822);
or UO_3217 (O_3217,N_29955,N_29701);
and UO_3218 (O_3218,N_29812,N_29890);
nand UO_3219 (O_3219,N_29910,N_29772);
and UO_3220 (O_3220,N_29961,N_29756);
xnor UO_3221 (O_3221,N_29824,N_29727);
nor UO_3222 (O_3222,N_29884,N_29890);
nor UO_3223 (O_3223,N_29714,N_29955);
or UO_3224 (O_3224,N_29764,N_29797);
and UO_3225 (O_3225,N_29916,N_29855);
nand UO_3226 (O_3226,N_29945,N_29841);
and UO_3227 (O_3227,N_29799,N_29739);
or UO_3228 (O_3228,N_29958,N_29827);
or UO_3229 (O_3229,N_29837,N_29912);
or UO_3230 (O_3230,N_29780,N_29865);
and UO_3231 (O_3231,N_29958,N_29833);
nor UO_3232 (O_3232,N_29870,N_29797);
nand UO_3233 (O_3233,N_29938,N_29931);
xnor UO_3234 (O_3234,N_29733,N_29950);
and UO_3235 (O_3235,N_29977,N_29897);
nor UO_3236 (O_3236,N_29920,N_29877);
and UO_3237 (O_3237,N_29847,N_29872);
or UO_3238 (O_3238,N_29993,N_29736);
xor UO_3239 (O_3239,N_29855,N_29772);
nor UO_3240 (O_3240,N_29881,N_29764);
nand UO_3241 (O_3241,N_29880,N_29754);
and UO_3242 (O_3242,N_29962,N_29982);
nor UO_3243 (O_3243,N_29801,N_29903);
or UO_3244 (O_3244,N_29936,N_29707);
nand UO_3245 (O_3245,N_29919,N_29958);
nor UO_3246 (O_3246,N_29759,N_29963);
or UO_3247 (O_3247,N_29959,N_29794);
or UO_3248 (O_3248,N_29905,N_29799);
and UO_3249 (O_3249,N_29841,N_29869);
or UO_3250 (O_3250,N_29780,N_29930);
or UO_3251 (O_3251,N_29984,N_29900);
and UO_3252 (O_3252,N_29730,N_29959);
xnor UO_3253 (O_3253,N_29816,N_29711);
and UO_3254 (O_3254,N_29845,N_29938);
nor UO_3255 (O_3255,N_29815,N_29869);
nand UO_3256 (O_3256,N_29828,N_29957);
nor UO_3257 (O_3257,N_29828,N_29905);
or UO_3258 (O_3258,N_29942,N_29881);
nand UO_3259 (O_3259,N_29738,N_29903);
nor UO_3260 (O_3260,N_29805,N_29771);
and UO_3261 (O_3261,N_29949,N_29804);
and UO_3262 (O_3262,N_29805,N_29712);
nor UO_3263 (O_3263,N_29883,N_29927);
xor UO_3264 (O_3264,N_29979,N_29896);
xnor UO_3265 (O_3265,N_29776,N_29998);
xor UO_3266 (O_3266,N_29972,N_29946);
nor UO_3267 (O_3267,N_29883,N_29711);
and UO_3268 (O_3268,N_29753,N_29934);
nor UO_3269 (O_3269,N_29781,N_29797);
nand UO_3270 (O_3270,N_29710,N_29774);
or UO_3271 (O_3271,N_29803,N_29913);
or UO_3272 (O_3272,N_29864,N_29970);
or UO_3273 (O_3273,N_29910,N_29735);
and UO_3274 (O_3274,N_29942,N_29995);
and UO_3275 (O_3275,N_29904,N_29968);
and UO_3276 (O_3276,N_29964,N_29952);
nand UO_3277 (O_3277,N_29867,N_29750);
and UO_3278 (O_3278,N_29849,N_29885);
xnor UO_3279 (O_3279,N_29857,N_29818);
or UO_3280 (O_3280,N_29987,N_29901);
and UO_3281 (O_3281,N_29776,N_29812);
or UO_3282 (O_3282,N_29789,N_29833);
or UO_3283 (O_3283,N_29728,N_29816);
nor UO_3284 (O_3284,N_29844,N_29953);
nand UO_3285 (O_3285,N_29733,N_29807);
xor UO_3286 (O_3286,N_29721,N_29733);
xnor UO_3287 (O_3287,N_29783,N_29865);
and UO_3288 (O_3288,N_29855,N_29919);
and UO_3289 (O_3289,N_29957,N_29838);
and UO_3290 (O_3290,N_29848,N_29807);
nor UO_3291 (O_3291,N_29841,N_29727);
xor UO_3292 (O_3292,N_29802,N_29961);
nor UO_3293 (O_3293,N_29737,N_29986);
nand UO_3294 (O_3294,N_29859,N_29796);
and UO_3295 (O_3295,N_29873,N_29722);
nand UO_3296 (O_3296,N_29925,N_29974);
nand UO_3297 (O_3297,N_29717,N_29963);
and UO_3298 (O_3298,N_29971,N_29947);
nor UO_3299 (O_3299,N_29905,N_29857);
or UO_3300 (O_3300,N_29914,N_29959);
or UO_3301 (O_3301,N_29869,N_29894);
nand UO_3302 (O_3302,N_29804,N_29985);
or UO_3303 (O_3303,N_29966,N_29778);
xor UO_3304 (O_3304,N_29907,N_29876);
or UO_3305 (O_3305,N_29995,N_29851);
xnor UO_3306 (O_3306,N_29851,N_29727);
nand UO_3307 (O_3307,N_29952,N_29913);
nor UO_3308 (O_3308,N_29907,N_29748);
xnor UO_3309 (O_3309,N_29995,N_29845);
and UO_3310 (O_3310,N_29804,N_29854);
nor UO_3311 (O_3311,N_29839,N_29788);
nor UO_3312 (O_3312,N_29794,N_29785);
nor UO_3313 (O_3313,N_29759,N_29741);
xor UO_3314 (O_3314,N_29797,N_29730);
nor UO_3315 (O_3315,N_29861,N_29921);
or UO_3316 (O_3316,N_29822,N_29764);
nand UO_3317 (O_3317,N_29950,N_29917);
xnor UO_3318 (O_3318,N_29936,N_29975);
or UO_3319 (O_3319,N_29952,N_29969);
and UO_3320 (O_3320,N_29763,N_29804);
or UO_3321 (O_3321,N_29789,N_29999);
and UO_3322 (O_3322,N_29954,N_29844);
nor UO_3323 (O_3323,N_29888,N_29990);
nor UO_3324 (O_3324,N_29770,N_29964);
xor UO_3325 (O_3325,N_29888,N_29948);
xnor UO_3326 (O_3326,N_29871,N_29745);
xor UO_3327 (O_3327,N_29758,N_29755);
and UO_3328 (O_3328,N_29904,N_29963);
or UO_3329 (O_3329,N_29930,N_29757);
and UO_3330 (O_3330,N_29722,N_29761);
nor UO_3331 (O_3331,N_29857,N_29888);
nor UO_3332 (O_3332,N_29986,N_29711);
xor UO_3333 (O_3333,N_29720,N_29853);
nand UO_3334 (O_3334,N_29843,N_29929);
nor UO_3335 (O_3335,N_29925,N_29850);
xor UO_3336 (O_3336,N_29900,N_29820);
or UO_3337 (O_3337,N_29965,N_29983);
and UO_3338 (O_3338,N_29853,N_29716);
or UO_3339 (O_3339,N_29962,N_29907);
and UO_3340 (O_3340,N_29744,N_29919);
or UO_3341 (O_3341,N_29800,N_29944);
nor UO_3342 (O_3342,N_29795,N_29940);
nor UO_3343 (O_3343,N_29700,N_29907);
nor UO_3344 (O_3344,N_29915,N_29977);
nor UO_3345 (O_3345,N_29935,N_29964);
and UO_3346 (O_3346,N_29890,N_29956);
or UO_3347 (O_3347,N_29908,N_29863);
and UO_3348 (O_3348,N_29778,N_29704);
or UO_3349 (O_3349,N_29896,N_29703);
xor UO_3350 (O_3350,N_29808,N_29969);
nor UO_3351 (O_3351,N_29888,N_29991);
xor UO_3352 (O_3352,N_29925,N_29834);
nor UO_3353 (O_3353,N_29726,N_29833);
and UO_3354 (O_3354,N_29958,N_29830);
nor UO_3355 (O_3355,N_29755,N_29965);
nor UO_3356 (O_3356,N_29784,N_29743);
nor UO_3357 (O_3357,N_29932,N_29814);
or UO_3358 (O_3358,N_29775,N_29717);
xnor UO_3359 (O_3359,N_29789,N_29844);
and UO_3360 (O_3360,N_29997,N_29881);
or UO_3361 (O_3361,N_29759,N_29822);
or UO_3362 (O_3362,N_29816,N_29824);
nand UO_3363 (O_3363,N_29735,N_29995);
nand UO_3364 (O_3364,N_29946,N_29982);
xnor UO_3365 (O_3365,N_29947,N_29848);
nor UO_3366 (O_3366,N_29820,N_29921);
nand UO_3367 (O_3367,N_29802,N_29874);
and UO_3368 (O_3368,N_29863,N_29763);
nor UO_3369 (O_3369,N_29801,N_29997);
nand UO_3370 (O_3370,N_29967,N_29915);
and UO_3371 (O_3371,N_29937,N_29998);
or UO_3372 (O_3372,N_29925,N_29898);
or UO_3373 (O_3373,N_29971,N_29852);
nand UO_3374 (O_3374,N_29866,N_29753);
or UO_3375 (O_3375,N_29942,N_29760);
nor UO_3376 (O_3376,N_29887,N_29937);
xnor UO_3377 (O_3377,N_29978,N_29845);
nor UO_3378 (O_3378,N_29738,N_29792);
or UO_3379 (O_3379,N_29721,N_29934);
or UO_3380 (O_3380,N_29854,N_29882);
or UO_3381 (O_3381,N_29849,N_29894);
and UO_3382 (O_3382,N_29964,N_29968);
and UO_3383 (O_3383,N_29795,N_29746);
and UO_3384 (O_3384,N_29708,N_29863);
nor UO_3385 (O_3385,N_29892,N_29866);
or UO_3386 (O_3386,N_29975,N_29957);
xnor UO_3387 (O_3387,N_29872,N_29718);
and UO_3388 (O_3388,N_29899,N_29759);
or UO_3389 (O_3389,N_29741,N_29769);
nor UO_3390 (O_3390,N_29894,N_29918);
nand UO_3391 (O_3391,N_29753,N_29999);
or UO_3392 (O_3392,N_29783,N_29841);
nor UO_3393 (O_3393,N_29798,N_29852);
nand UO_3394 (O_3394,N_29957,N_29939);
and UO_3395 (O_3395,N_29950,N_29805);
and UO_3396 (O_3396,N_29765,N_29725);
or UO_3397 (O_3397,N_29989,N_29748);
nor UO_3398 (O_3398,N_29845,N_29991);
nand UO_3399 (O_3399,N_29730,N_29844);
nand UO_3400 (O_3400,N_29921,N_29828);
nor UO_3401 (O_3401,N_29757,N_29890);
nor UO_3402 (O_3402,N_29926,N_29798);
nor UO_3403 (O_3403,N_29857,N_29982);
nor UO_3404 (O_3404,N_29777,N_29726);
nand UO_3405 (O_3405,N_29729,N_29941);
nor UO_3406 (O_3406,N_29739,N_29994);
and UO_3407 (O_3407,N_29748,N_29914);
xnor UO_3408 (O_3408,N_29953,N_29885);
and UO_3409 (O_3409,N_29741,N_29928);
and UO_3410 (O_3410,N_29959,N_29754);
nor UO_3411 (O_3411,N_29859,N_29846);
or UO_3412 (O_3412,N_29968,N_29839);
and UO_3413 (O_3413,N_29739,N_29911);
or UO_3414 (O_3414,N_29710,N_29938);
and UO_3415 (O_3415,N_29987,N_29929);
xor UO_3416 (O_3416,N_29855,N_29991);
xnor UO_3417 (O_3417,N_29813,N_29924);
xnor UO_3418 (O_3418,N_29772,N_29897);
and UO_3419 (O_3419,N_29719,N_29875);
xor UO_3420 (O_3420,N_29943,N_29971);
xnor UO_3421 (O_3421,N_29799,N_29701);
and UO_3422 (O_3422,N_29806,N_29829);
nor UO_3423 (O_3423,N_29792,N_29914);
and UO_3424 (O_3424,N_29912,N_29846);
nor UO_3425 (O_3425,N_29904,N_29710);
nor UO_3426 (O_3426,N_29707,N_29945);
and UO_3427 (O_3427,N_29860,N_29708);
and UO_3428 (O_3428,N_29960,N_29747);
and UO_3429 (O_3429,N_29840,N_29892);
or UO_3430 (O_3430,N_29943,N_29844);
and UO_3431 (O_3431,N_29987,N_29820);
nor UO_3432 (O_3432,N_29971,N_29820);
nand UO_3433 (O_3433,N_29829,N_29956);
nor UO_3434 (O_3434,N_29822,N_29936);
xnor UO_3435 (O_3435,N_29815,N_29853);
nand UO_3436 (O_3436,N_29844,N_29978);
or UO_3437 (O_3437,N_29932,N_29864);
and UO_3438 (O_3438,N_29948,N_29808);
nor UO_3439 (O_3439,N_29812,N_29804);
nand UO_3440 (O_3440,N_29747,N_29751);
xnor UO_3441 (O_3441,N_29820,N_29984);
xor UO_3442 (O_3442,N_29983,N_29980);
nand UO_3443 (O_3443,N_29994,N_29821);
and UO_3444 (O_3444,N_29879,N_29989);
or UO_3445 (O_3445,N_29934,N_29800);
xor UO_3446 (O_3446,N_29954,N_29962);
or UO_3447 (O_3447,N_29956,N_29849);
xnor UO_3448 (O_3448,N_29787,N_29882);
and UO_3449 (O_3449,N_29722,N_29843);
nor UO_3450 (O_3450,N_29755,N_29887);
nor UO_3451 (O_3451,N_29706,N_29862);
nor UO_3452 (O_3452,N_29729,N_29973);
or UO_3453 (O_3453,N_29821,N_29824);
nand UO_3454 (O_3454,N_29773,N_29778);
and UO_3455 (O_3455,N_29706,N_29970);
and UO_3456 (O_3456,N_29802,N_29812);
or UO_3457 (O_3457,N_29845,N_29841);
and UO_3458 (O_3458,N_29889,N_29869);
xor UO_3459 (O_3459,N_29948,N_29723);
nand UO_3460 (O_3460,N_29769,N_29913);
nor UO_3461 (O_3461,N_29978,N_29821);
and UO_3462 (O_3462,N_29918,N_29800);
and UO_3463 (O_3463,N_29828,N_29945);
nor UO_3464 (O_3464,N_29784,N_29844);
or UO_3465 (O_3465,N_29816,N_29718);
and UO_3466 (O_3466,N_29979,N_29841);
xor UO_3467 (O_3467,N_29711,N_29905);
and UO_3468 (O_3468,N_29993,N_29710);
nand UO_3469 (O_3469,N_29884,N_29921);
and UO_3470 (O_3470,N_29767,N_29922);
nor UO_3471 (O_3471,N_29771,N_29918);
xor UO_3472 (O_3472,N_29815,N_29739);
nor UO_3473 (O_3473,N_29999,N_29899);
nand UO_3474 (O_3474,N_29793,N_29992);
nor UO_3475 (O_3475,N_29768,N_29834);
or UO_3476 (O_3476,N_29866,N_29828);
and UO_3477 (O_3477,N_29944,N_29795);
nand UO_3478 (O_3478,N_29992,N_29950);
xor UO_3479 (O_3479,N_29805,N_29879);
nor UO_3480 (O_3480,N_29849,N_29855);
nand UO_3481 (O_3481,N_29841,N_29705);
nor UO_3482 (O_3482,N_29922,N_29980);
and UO_3483 (O_3483,N_29804,N_29867);
and UO_3484 (O_3484,N_29913,N_29787);
nor UO_3485 (O_3485,N_29872,N_29760);
nor UO_3486 (O_3486,N_29725,N_29744);
and UO_3487 (O_3487,N_29737,N_29710);
nand UO_3488 (O_3488,N_29902,N_29719);
or UO_3489 (O_3489,N_29850,N_29976);
or UO_3490 (O_3490,N_29825,N_29936);
nor UO_3491 (O_3491,N_29713,N_29701);
and UO_3492 (O_3492,N_29810,N_29948);
and UO_3493 (O_3493,N_29797,N_29947);
nand UO_3494 (O_3494,N_29803,N_29790);
nor UO_3495 (O_3495,N_29845,N_29749);
nand UO_3496 (O_3496,N_29939,N_29851);
and UO_3497 (O_3497,N_29886,N_29987);
nor UO_3498 (O_3498,N_29769,N_29792);
nand UO_3499 (O_3499,N_29947,N_29798);
endmodule