module basic_1000_10000_1500_10_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_91,In_441);
or U1 (N_1,In_452,In_532);
nor U2 (N_2,In_692,In_501);
nor U3 (N_3,In_348,In_940);
nand U4 (N_4,In_423,In_828);
and U5 (N_5,In_285,In_449);
xnor U6 (N_6,In_725,In_35);
xnor U7 (N_7,In_572,In_787);
or U8 (N_8,In_276,In_155);
xnor U9 (N_9,In_139,In_946);
nor U10 (N_10,In_502,In_862);
nor U11 (N_11,In_970,In_41);
nor U12 (N_12,In_972,In_173);
and U13 (N_13,In_614,In_621);
nor U14 (N_14,In_841,In_987);
or U15 (N_15,In_577,In_749);
nor U16 (N_16,In_683,In_172);
and U17 (N_17,In_873,In_542);
and U18 (N_18,In_758,In_989);
nand U19 (N_19,In_837,In_136);
nand U20 (N_20,In_631,In_229);
nor U21 (N_21,In_677,In_370);
xnor U22 (N_22,In_999,In_273);
nor U23 (N_23,In_9,In_905);
xor U24 (N_24,In_323,In_354);
nand U25 (N_25,In_521,In_96);
or U26 (N_26,In_295,In_208);
xor U27 (N_27,In_933,In_930);
and U28 (N_28,In_805,In_412);
nor U29 (N_29,In_639,In_986);
or U30 (N_30,In_942,In_798);
and U31 (N_31,In_55,In_153);
or U32 (N_32,In_187,In_777);
xor U33 (N_33,In_495,In_437);
xor U34 (N_34,In_813,In_255);
or U35 (N_35,In_498,In_536);
nor U36 (N_36,In_269,In_786);
nand U37 (N_37,In_839,In_253);
or U38 (N_38,In_890,In_235);
or U39 (N_39,In_699,In_410);
xor U40 (N_40,In_145,In_181);
xnor U41 (N_41,In_723,In_678);
nand U42 (N_42,In_360,In_247);
or U43 (N_43,In_53,In_591);
nor U44 (N_44,In_59,In_859);
and U45 (N_45,In_259,In_518);
nand U46 (N_46,In_779,In_979);
xor U47 (N_47,In_705,In_734);
nand U48 (N_48,In_543,In_847);
nand U49 (N_49,In_445,In_934);
xnor U50 (N_50,In_277,In_346);
and U51 (N_51,In_632,In_781);
or U52 (N_52,In_286,In_178);
or U53 (N_53,In_368,In_887);
or U54 (N_54,In_846,In_687);
nand U55 (N_55,In_119,In_160);
and U56 (N_56,In_559,In_328);
or U57 (N_57,In_785,In_684);
or U58 (N_58,In_802,In_857);
and U59 (N_59,In_922,In_806);
xnor U60 (N_60,In_949,In_988);
or U61 (N_61,In_243,In_199);
xor U62 (N_62,In_612,In_405);
and U63 (N_63,In_5,In_827);
or U64 (N_64,In_739,In_895);
nand U65 (N_65,In_533,In_820);
nor U66 (N_66,In_465,In_82);
nand U67 (N_67,In_822,In_225);
nor U68 (N_68,In_460,In_546);
nand U69 (N_69,In_38,In_48);
or U70 (N_70,In_404,In_448);
xnor U71 (N_71,In_417,In_27);
xor U72 (N_72,In_755,In_896);
xor U73 (N_73,In_603,In_158);
and U74 (N_74,In_192,In_224);
nand U75 (N_75,In_975,In_899);
nand U76 (N_76,In_171,In_945);
or U77 (N_77,In_668,In_525);
nand U78 (N_78,In_752,In_743);
and U79 (N_79,In_461,In_454);
nand U80 (N_80,In_369,In_455);
xor U81 (N_81,In_244,In_105);
and U82 (N_82,In_925,In_843);
and U83 (N_83,In_64,In_37);
and U84 (N_84,In_558,In_177);
or U85 (N_85,In_713,In_450);
nor U86 (N_86,In_117,In_914);
xnor U87 (N_87,In_304,In_485);
xnor U88 (N_88,In_353,In_505);
xnor U89 (N_89,In_983,In_362);
nand U90 (N_90,In_590,In_361);
and U91 (N_91,In_974,In_425);
nand U92 (N_92,In_241,In_409);
or U93 (N_93,In_651,In_990);
nand U94 (N_94,In_504,In_218);
xor U95 (N_95,In_729,In_977);
nor U96 (N_96,In_963,In_152);
nor U97 (N_97,In_951,In_645);
nand U98 (N_98,In_363,In_263);
and U99 (N_99,In_894,In_245);
xnor U100 (N_100,In_565,In_867);
nor U101 (N_101,In_341,In_732);
nand U102 (N_102,In_882,In_954);
nor U103 (N_103,In_99,In_955);
and U104 (N_104,In_54,In_724);
nand U105 (N_105,In_625,In_3);
xnor U106 (N_106,In_234,In_649);
and U107 (N_107,In_636,In_403);
and U108 (N_108,In_782,In_86);
or U109 (N_109,In_686,In_594);
xnor U110 (N_110,In_20,In_834);
or U111 (N_111,In_694,In_134);
and U112 (N_112,In_549,In_115);
nand U113 (N_113,In_670,In_297);
and U114 (N_114,In_903,In_650);
and U115 (N_115,In_811,In_588);
and U116 (N_116,In_201,In_855);
and U117 (N_117,In_500,In_489);
nor U118 (N_118,In_406,In_534);
and U119 (N_119,In_578,In_90);
nor U120 (N_120,In_167,In_142);
nor U121 (N_121,In_206,In_791);
or U122 (N_122,In_750,In_960);
or U123 (N_123,In_151,In_359);
and U124 (N_124,In_231,In_697);
nor U125 (N_125,In_561,In_540);
or U126 (N_126,In_667,In_967);
nand U127 (N_127,In_597,In_832);
xor U128 (N_128,In_763,In_716);
and U129 (N_129,In_608,In_672);
nand U130 (N_130,In_585,In_767);
and U131 (N_131,In_164,In_611);
nand U132 (N_132,In_110,In_522);
nand U133 (N_133,In_331,In_10);
and U134 (N_134,In_596,In_309);
and U135 (N_135,In_459,In_36);
or U136 (N_136,In_122,In_355);
nor U137 (N_137,In_49,In_2);
nand U138 (N_138,In_23,In_394);
and U139 (N_139,In_923,In_202);
xnor U140 (N_140,In_364,In_601);
or U141 (N_141,In_21,In_278);
or U142 (N_142,In_194,In_443);
nor U143 (N_143,In_97,In_108);
or U144 (N_144,In_529,In_275);
or U145 (N_145,In_961,In_642);
nor U146 (N_146,In_929,In_228);
nor U147 (N_147,In_124,In_127);
nor U148 (N_148,In_270,In_560);
or U149 (N_149,In_702,In_301);
or U150 (N_150,In_726,In_908);
xor U151 (N_151,In_6,In_200);
xor U152 (N_152,In_72,In_784);
nor U153 (N_153,In_290,In_736);
nand U154 (N_154,In_901,In_79);
nor U155 (N_155,In_809,In_400);
xnor U156 (N_156,In_288,In_366);
and U157 (N_157,In_95,In_681);
or U158 (N_158,In_907,In_324);
nor U159 (N_159,In_149,In_720);
xor U160 (N_160,In_126,In_89);
nor U161 (N_161,In_314,In_570);
xnor U162 (N_162,In_866,In_801);
xor U163 (N_163,In_858,In_321);
or U164 (N_164,In_250,In_204);
or U165 (N_165,In_146,In_11);
nand U166 (N_166,In_913,In_641);
nand U167 (N_167,In_804,In_302);
nor U168 (N_168,In_159,In_595);
nand U169 (N_169,In_60,In_564);
nor U170 (N_170,In_428,In_969);
or U171 (N_171,In_156,In_333);
and U172 (N_172,In_580,In_633);
nor U173 (N_173,In_438,In_757);
xor U174 (N_174,In_615,In_610);
or U175 (N_175,In_93,In_469);
nor U176 (N_176,In_640,In_952);
and U177 (N_177,In_329,In_327);
or U178 (N_178,In_481,In_212);
and U179 (N_179,In_180,In_818);
xor U180 (N_180,In_563,In_402);
and U181 (N_181,In_143,In_413);
xnor U182 (N_182,In_282,In_665);
nand U183 (N_183,In_8,In_797);
and U184 (N_184,In_807,In_795);
nor U185 (N_185,In_593,In_358);
and U186 (N_186,In_98,In_15);
nand U187 (N_187,In_22,In_680);
nor U188 (N_188,In_898,In_345);
and U189 (N_189,In_831,In_34);
nand U190 (N_190,In_819,In_81);
or U191 (N_191,In_685,In_148);
xor U192 (N_192,In_374,In_322);
xnor U193 (N_193,In_861,In_393);
nand U194 (N_194,In_131,In_966);
xnor U195 (N_195,In_874,In_917);
nor U196 (N_196,In_496,In_381);
or U197 (N_197,In_436,In_150);
xor U198 (N_198,In_503,In_185);
nand U199 (N_199,In_691,In_424);
xor U200 (N_200,In_814,In_372);
nand U201 (N_201,In_617,In_390);
or U202 (N_202,In_753,In_733);
or U203 (N_203,In_58,In_238);
nand U204 (N_204,In_926,In_770);
nor U205 (N_205,In_512,In_102);
nand U206 (N_206,In_56,In_63);
or U207 (N_207,In_499,In_161);
nand U208 (N_208,In_833,In_220);
and U209 (N_209,In_216,In_984);
or U210 (N_210,In_658,In_766);
nor U211 (N_211,In_884,In_384);
and U212 (N_212,In_464,In_936);
nand U213 (N_213,In_415,In_492);
nor U214 (N_214,In_69,In_24);
nand U215 (N_215,In_912,In_266);
xor U216 (N_216,In_386,In_271);
nor U217 (N_217,In_947,In_219);
and U218 (N_218,In_183,In_352);
xor U219 (N_219,In_62,In_104);
nand U220 (N_220,In_883,In_715);
nor U221 (N_221,In_399,In_12);
or U222 (N_222,In_256,In_65);
xor U223 (N_223,In_511,In_623);
and U224 (N_224,In_943,In_881);
nand U225 (N_225,In_125,In_919);
or U226 (N_226,In_682,In_526);
nand U227 (N_227,In_921,In_554);
nor U228 (N_228,In_87,In_457);
nand U229 (N_229,In_135,In_573);
nor U230 (N_230,In_109,In_854);
or U231 (N_231,In_924,In_848);
and U232 (N_232,In_427,In_78);
or U233 (N_233,In_196,In_287);
nand U234 (N_234,In_523,In_664);
or U235 (N_235,In_868,In_551);
nand U236 (N_236,In_154,In_392);
xnor U237 (N_237,In_293,In_85);
nand U238 (N_238,In_824,In_28);
or U239 (N_239,In_888,In_530);
xor U240 (N_240,In_137,In_637);
and U241 (N_241,In_175,In_812);
and U242 (N_242,In_43,In_872);
xnor U243 (N_243,In_429,In_274);
or U244 (N_244,In_738,In_773);
nor U245 (N_245,In_418,In_111);
or U246 (N_246,In_491,In_870);
nand U247 (N_247,In_928,In_607);
xnor U248 (N_248,In_19,In_982);
or U249 (N_249,In_176,In_434);
and U250 (N_250,In_391,In_476);
nor U251 (N_251,In_380,In_1);
nand U252 (N_252,In_996,In_182);
and U253 (N_253,In_864,In_584);
or U254 (N_254,In_67,In_299);
nor U255 (N_255,In_211,In_326);
or U256 (N_256,In_45,In_604);
and U257 (N_257,In_860,In_179);
or U258 (N_258,In_435,In_261);
and U259 (N_259,In_292,In_956);
nor U260 (N_260,In_655,In_83);
or U261 (N_261,In_193,In_889);
and U262 (N_262,In_973,In_215);
xnor U263 (N_263,In_432,In_774);
and U264 (N_264,In_576,In_877);
nand U265 (N_265,In_408,In_567);
nand U266 (N_266,In_959,In_316);
xor U267 (N_267,In_365,In_991);
nand U268 (N_268,In_772,In_927);
nand U269 (N_269,In_446,In_16);
or U270 (N_270,In_935,In_319);
nor U271 (N_271,In_138,In_467);
nand U272 (N_272,In_948,In_679);
and U273 (N_273,In_660,In_852);
or U274 (N_274,In_473,In_357);
and U275 (N_275,In_32,In_7);
nor U276 (N_276,In_902,In_994);
nor U277 (N_277,In_998,In_470);
or U278 (N_278,In_906,In_188);
xnor U279 (N_279,In_482,In_147);
nor U280 (N_280,In_606,In_307);
and U281 (N_281,In_688,In_373);
nand U282 (N_282,In_630,In_764);
and U283 (N_283,In_325,In_711);
and U284 (N_284,In_821,In_133);
and U285 (N_285,In_490,In_722);
or U286 (N_286,In_387,In_51);
nand U287 (N_287,In_94,In_33);
or U288 (N_288,In_447,In_652);
xnor U289 (N_289,In_26,In_466);
nand U290 (N_290,In_618,In_856);
nand U291 (N_291,In_426,In_265);
nand U292 (N_292,In_296,In_0);
xor U293 (N_293,In_57,In_792);
nand U294 (N_294,In_289,In_165);
nor U295 (N_295,In_789,In_221);
and U296 (N_296,In_579,In_592);
or U297 (N_297,In_574,In_396);
nand U298 (N_298,In_708,In_790);
xnor U299 (N_299,In_704,In_920);
xor U300 (N_300,In_283,In_748);
or U301 (N_301,In_507,In_941);
or U302 (N_302,In_456,In_968);
nand U303 (N_303,In_616,In_474);
nand U304 (N_304,In_629,In_422);
or U305 (N_305,In_581,In_262);
and U306 (N_306,In_31,In_510);
xor U307 (N_307,In_932,In_762);
or U308 (N_308,In_342,In_520);
nand U309 (N_309,In_128,In_897);
nand U310 (N_310,In_144,In_421);
nand U311 (N_311,In_214,In_953);
or U312 (N_312,In_203,In_728);
xnor U313 (N_313,In_132,In_350);
or U314 (N_314,In_398,In_783);
nand U315 (N_315,In_184,In_39);
or U316 (N_316,In_537,In_740);
xor U317 (N_317,In_291,In_971);
xnor U318 (N_318,In_318,In_416);
nand U319 (N_319,In_880,In_258);
and U320 (N_320,In_68,In_550);
nand U321 (N_321,In_674,In_524);
nand U322 (N_322,In_675,In_553);
nand U323 (N_323,In_628,In_844);
nor U324 (N_324,In_337,In_430);
and U325 (N_325,In_130,In_721);
or U326 (N_326,In_300,In_311);
nand U327 (N_327,In_508,In_205);
xor U328 (N_328,In_186,In_569);
xor U329 (N_329,In_483,In_622);
xnor U330 (N_330,In_92,In_746);
xnor U331 (N_331,In_817,In_778);
nor U332 (N_332,In_190,In_75);
xnor U333 (N_333,In_74,In_317);
xor U334 (N_334,In_433,In_237);
and U335 (N_335,In_810,In_871);
and U336 (N_336,In_442,In_700);
nor U337 (N_337,In_305,In_878);
and U338 (N_338,In_727,In_714);
or U339 (N_339,In_472,In_768);
nand U340 (N_340,In_599,In_440);
nor U341 (N_341,In_892,In_497);
nor U342 (N_342,In_118,In_842);
or U343 (N_343,In_635,In_479);
and U344 (N_344,In_571,In_937);
or U345 (N_345,In_251,In_545);
nand U346 (N_346,In_50,In_556);
or U347 (N_347,In_760,In_566);
nor U348 (N_348,In_965,In_775);
and U349 (N_349,In_869,In_835);
and U350 (N_350,In_539,In_227);
nor U351 (N_351,In_462,In_162);
nor U352 (N_352,In_661,In_771);
nor U353 (N_353,In_815,In_332);
or U354 (N_354,In_931,In_279);
xor U355 (N_355,In_382,In_958);
and U356 (N_356,In_379,In_646);
and U357 (N_357,In_562,In_647);
or U358 (N_358,In_347,In_166);
nand U359 (N_359,In_602,In_981);
nor U360 (N_360,In_825,In_303);
and U361 (N_361,In_793,In_915);
xor U362 (N_362,In_992,In_826);
xor U363 (N_363,In_336,In_663);
nor U364 (N_364,In_737,In_338);
nor U365 (N_365,In_385,In_875);
or U366 (N_366,In_803,In_910);
and U367 (N_367,In_306,In_264);
nand U368 (N_368,In_310,In_605);
xor U369 (N_369,In_76,In_918);
and U370 (N_370,In_140,In_718);
xnor U371 (N_371,In_197,In_344);
nand U372 (N_372,In_70,In_61);
and U373 (N_373,In_669,In_800);
and U374 (N_374,In_751,In_653);
or U375 (N_375,In_547,In_541);
xnor U376 (N_376,In_378,In_334);
nor U377 (N_377,In_463,In_643);
nor U378 (N_378,In_589,In_340);
nor U379 (N_379,In_414,In_313);
nand U380 (N_380,In_535,In_493);
xor U381 (N_381,In_349,In_985);
or U382 (N_382,In_850,In_356);
xnor U383 (N_383,In_52,In_478);
xor U384 (N_384,In_488,In_320);
nand U385 (N_385,In_281,In_233);
or U386 (N_386,In_308,In_213);
xnor U387 (N_387,In_169,In_788);
nor U388 (N_388,In_552,In_376);
xor U389 (N_389,In_916,In_477);
and U390 (N_390,In_648,In_769);
nor U391 (N_391,In_236,In_997);
xor U392 (N_392,In_246,In_30);
and U393 (N_393,In_717,In_745);
and U394 (N_394,In_829,In_619);
and U395 (N_395,In_239,In_252);
and U396 (N_396,In_315,In_557);
nand U397 (N_397,In_397,In_312);
nor U398 (N_398,In_853,In_885);
xnor U399 (N_399,In_84,In_849);
nor U400 (N_400,In_609,In_29);
xnor U401 (N_401,In_257,In_845);
or U402 (N_402,In_624,In_248);
and U403 (N_403,In_506,In_475);
and U404 (N_404,In_101,In_42);
nand U405 (N_405,In_575,In_389);
or U406 (N_406,In_367,In_710);
nor U407 (N_407,In_112,In_993);
nand U408 (N_408,In_480,In_747);
nand U409 (N_409,In_893,In_174);
nand U410 (N_410,In_453,In_189);
and U411 (N_411,In_695,In_88);
or U412 (N_412,In_383,In_904);
and U413 (N_413,In_226,In_731);
nor U414 (N_414,In_71,In_451);
or U415 (N_415,In_555,In_712);
nand U416 (N_416,In_582,In_528);
nand U417 (N_417,In_388,In_330);
xor U418 (N_418,In_47,In_494);
nand U419 (N_419,In_44,In_343);
xnor U420 (N_420,In_484,In_876);
and U421 (N_421,In_909,In_116);
and U422 (N_422,In_964,In_851);
nand U423 (N_423,In_657,In_780);
xor U424 (N_424,In_891,In_444);
nand U425 (N_425,In_170,In_911);
nand U426 (N_426,In_335,In_613);
nand U427 (N_427,In_207,In_163);
nand U428 (N_428,In_280,In_620);
nand U429 (N_429,In_701,In_249);
nand U430 (N_430,In_995,In_223);
nand U431 (N_431,In_458,In_268);
nor U432 (N_432,In_730,In_886);
or U433 (N_433,In_25,In_230);
or U434 (N_434,In_676,In_260);
nor U435 (N_435,In_962,In_209);
xnor U436 (N_436,In_698,In_598);
xor U437 (N_437,In_950,In_531);
nor U438 (N_438,In_836,In_298);
nor U439 (N_439,In_754,In_939);
and U440 (N_440,In_107,In_375);
nor U441 (N_441,In_420,In_18);
or U442 (N_442,In_100,In_794);
nand U443 (N_443,In_538,In_816);
or U444 (N_444,In_519,In_863);
or U445 (N_445,In_690,In_759);
nor U446 (N_446,In_395,In_267);
nor U447 (N_447,In_123,In_671);
nor U448 (N_448,In_401,In_627);
and U449 (N_449,In_13,In_106);
and U450 (N_450,In_976,In_865);
and U451 (N_451,In_516,In_113);
nor U452 (N_452,In_294,In_656);
nor U453 (N_453,In_900,In_129);
xnor U454 (N_454,In_696,In_742);
xnor U455 (N_455,In_634,In_411);
or U456 (N_456,In_14,In_487);
xor U457 (N_457,In_761,In_808);
xor U458 (N_458,In_548,In_586);
or U459 (N_459,In_513,In_222);
nor U460 (N_460,In_254,In_644);
or U461 (N_461,In_776,In_689);
nand U462 (N_462,In_103,In_735);
xnor U463 (N_463,In_600,In_756);
and U464 (N_464,In_114,In_938);
nand U465 (N_465,In_707,In_486);
nor U466 (N_466,In_40,In_240);
and U467 (N_467,In_823,In_799);
and U468 (N_468,In_944,In_583);
nor U469 (N_469,In_471,In_765);
xnor U470 (N_470,In_796,In_527);
xnor U471 (N_471,In_17,In_741);
nor U472 (N_472,In_73,In_232);
or U473 (N_473,In_377,In_351);
and U474 (N_474,In_709,In_439);
or U475 (N_475,In_879,In_957);
nand U476 (N_476,In_66,In_168);
nand U477 (N_477,In_121,In_514);
nor U478 (N_478,In_744,In_719);
nand U479 (N_479,In_830,In_659);
and U480 (N_480,In_654,In_568);
nor U481 (N_481,In_4,In_80);
and U482 (N_482,In_77,In_666);
nor U483 (N_483,In_120,In_339);
or U484 (N_484,In_673,In_468);
and U485 (N_485,In_210,In_217);
nand U486 (N_486,In_980,In_517);
and U487 (N_487,In_431,In_703);
nor U488 (N_488,In_419,In_157);
nand U489 (N_489,In_198,In_626);
nor U490 (N_490,In_407,In_587);
and U491 (N_491,In_706,In_46);
xnor U492 (N_492,In_693,In_371);
nand U493 (N_493,In_191,In_662);
and U494 (N_494,In_840,In_141);
or U495 (N_495,In_284,In_515);
xor U496 (N_496,In_509,In_838);
or U497 (N_497,In_638,In_195);
nand U498 (N_498,In_242,In_978);
xor U499 (N_499,In_272,In_544);
or U500 (N_500,In_57,In_943);
nor U501 (N_501,In_921,In_21);
nand U502 (N_502,In_492,In_145);
or U503 (N_503,In_548,In_161);
xnor U504 (N_504,In_878,In_672);
and U505 (N_505,In_170,In_359);
and U506 (N_506,In_151,In_760);
xnor U507 (N_507,In_64,In_282);
nand U508 (N_508,In_705,In_524);
and U509 (N_509,In_831,In_835);
and U510 (N_510,In_780,In_106);
nor U511 (N_511,In_267,In_211);
or U512 (N_512,In_591,In_90);
nor U513 (N_513,In_919,In_716);
nand U514 (N_514,In_537,In_385);
xnor U515 (N_515,In_96,In_816);
or U516 (N_516,In_664,In_351);
nor U517 (N_517,In_756,In_408);
nand U518 (N_518,In_213,In_894);
nand U519 (N_519,In_327,In_157);
or U520 (N_520,In_401,In_62);
nand U521 (N_521,In_13,In_916);
xor U522 (N_522,In_48,In_173);
nor U523 (N_523,In_904,In_941);
or U524 (N_524,In_938,In_885);
and U525 (N_525,In_199,In_798);
nand U526 (N_526,In_658,In_516);
or U527 (N_527,In_673,In_59);
nand U528 (N_528,In_369,In_61);
nor U529 (N_529,In_691,In_310);
and U530 (N_530,In_967,In_741);
nand U531 (N_531,In_552,In_541);
or U532 (N_532,In_653,In_478);
nor U533 (N_533,In_509,In_161);
xnor U534 (N_534,In_875,In_892);
xor U535 (N_535,In_142,In_330);
nor U536 (N_536,In_609,In_352);
or U537 (N_537,In_375,In_867);
nand U538 (N_538,In_591,In_717);
xor U539 (N_539,In_385,In_764);
or U540 (N_540,In_541,In_563);
xor U541 (N_541,In_719,In_804);
and U542 (N_542,In_817,In_753);
nand U543 (N_543,In_298,In_468);
xor U544 (N_544,In_65,In_637);
nor U545 (N_545,In_967,In_691);
and U546 (N_546,In_975,In_87);
nor U547 (N_547,In_610,In_15);
xnor U548 (N_548,In_833,In_551);
xnor U549 (N_549,In_548,In_627);
and U550 (N_550,In_335,In_584);
or U551 (N_551,In_890,In_332);
or U552 (N_552,In_661,In_869);
and U553 (N_553,In_475,In_499);
or U554 (N_554,In_881,In_977);
or U555 (N_555,In_2,In_527);
nand U556 (N_556,In_790,In_368);
nor U557 (N_557,In_516,In_288);
or U558 (N_558,In_849,In_95);
xnor U559 (N_559,In_5,In_221);
nand U560 (N_560,In_802,In_397);
nor U561 (N_561,In_422,In_572);
xor U562 (N_562,In_332,In_874);
nand U563 (N_563,In_41,In_575);
nand U564 (N_564,In_642,In_119);
or U565 (N_565,In_662,In_913);
or U566 (N_566,In_803,In_143);
nand U567 (N_567,In_315,In_777);
and U568 (N_568,In_553,In_996);
nand U569 (N_569,In_43,In_61);
or U570 (N_570,In_654,In_367);
nor U571 (N_571,In_110,In_367);
or U572 (N_572,In_145,In_629);
nor U573 (N_573,In_532,In_548);
and U574 (N_574,In_540,In_78);
or U575 (N_575,In_498,In_560);
xnor U576 (N_576,In_728,In_505);
nand U577 (N_577,In_137,In_459);
or U578 (N_578,In_523,In_257);
nor U579 (N_579,In_380,In_245);
nor U580 (N_580,In_240,In_963);
nor U581 (N_581,In_163,In_274);
xor U582 (N_582,In_532,In_483);
and U583 (N_583,In_74,In_924);
or U584 (N_584,In_605,In_193);
and U585 (N_585,In_643,In_248);
or U586 (N_586,In_64,In_182);
nand U587 (N_587,In_869,In_935);
and U588 (N_588,In_82,In_703);
or U589 (N_589,In_34,In_842);
and U590 (N_590,In_119,In_998);
and U591 (N_591,In_17,In_469);
or U592 (N_592,In_547,In_774);
xor U593 (N_593,In_514,In_970);
nand U594 (N_594,In_822,In_842);
or U595 (N_595,In_630,In_539);
nor U596 (N_596,In_485,In_49);
nor U597 (N_597,In_610,In_441);
xor U598 (N_598,In_929,In_120);
and U599 (N_599,In_506,In_818);
nand U600 (N_600,In_574,In_444);
or U601 (N_601,In_280,In_941);
nand U602 (N_602,In_154,In_564);
xnor U603 (N_603,In_253,In_433);
and U604 (N_604,In_757,In_119);
or U605 (N_605,In_968,In_43);
and U606 (N_606,In_85,In_818);
and U607 (N_607,In_553,In_864);
nor U608 (N_608,In_137,In_485);
or U609 (N_609,In_269,In_730);
or U610 (N_610,In_825,In_62);
nand U611 (N_611,In_387,In_633);
xnor U612 (N_612,In_982,In_210);
xnor U613 (N_613,In_381,In_847);
nand U614 (N_614,In_630,In_877);
or U615 (N_615,In_88,In_621);
and U616 (N_616,In_21,In_138);
and U617 (N_617,In_812,In_744);
xor U618 (N_618,In_400,In_96);
or U619 (N_619,In_335,In_579);
or U620 (N_620,In_541,In_471);
nand U621 (N_621,In_538,In_341);
xor U622 (N_622,In_233,In_621);
xnor U623 (N_623,In_385,In_204);
nand U624 (N_624,In_10,In_791);
or U625 (N_625,In_991,In_395);
and U626 (N_626,In_14,In_646);
xor U627 (N_627,In_574,In_598);
and U628 (N_628,In_215,In_234);
and U629 (N_629,In_137,In_979);
xor U630 (N_630,In_136,In_821);
or U631 (N_631,In_438,In_769);
and U632 (N_632,In_345,In_219);
nor U633 (N_633,In_18,In_857);
nand U634 (N_634,In_929,In_332);
nor U635 (N_635,In_702,In_265);
nor U636 (N_636,In_382,In_230);
nor U637 (N_637,In_503,In_597);
nor U638 (N_638,In_892,In_607);
and U639 (N_639,In_883,In_684);
and U640 (N_640,In_405,In_530);
nand U641 (N_641,In_989,In_934);
xnor U642 (N_642,In_161,In_388);
xor U643 (N_643,In_134,In_275);
and U644 (N_644,In_58,In_935);
or U645 (N_645,In_25,In_748);
nand U646 (N_646,In_439,In_467);
nor U647 (N_647,In_888,In_100);
and U648 (N_648,In_374,In_121);
and U649 (N_649,In_7,In_90);
nor U650 (N_650,In_593,In_368);
xnor U651 (N_651,In_817,In_453);
nor U652 (N_652,In_653,In_287);
nor U653 (N_653,In_737,In_923);
nand U654 (N_654,In_387,In_824);
or U655 (N_655,In_356,In_825);
and U656 (N_656,In_605,In_839);
or U657 (N_657,In_216,In_250);
nor U658 (N_658,In_764,In_341);
or U659 (N_659,In_298,In_457);
nor U660 (N_660,In_632,In_951);
nor U661 (N_661,In_860,In_834);
or U662 (N_662,In_303,In_466);
or U663 (N_663,In_81,In_865);
or U664 (N_664,In_169,In_167);
nand U665 (N_665,In_666,In_456);
or U666 (N_666,In_965,In_628);
nand U667 (N_667,In_240,In_251);
xor U668 (N_668,In_673,In_264);
xor U669 (N_669,In_476,In_372);
and U670 (N_670,In_672,In_609);
nor U671 (N_671,In_377,In_673);
nand U672 (N_672,In_842,In_361);
nor U673 (N_673,In_789,In_706);
nand U674 (N_674,In_455,In_865);
nand U675 (N_675,In_793,In_110);
or U676 (N_676,In_791,In_355);
nor U677 (N_677,In_503,In_736);
or U678 (N_678,In_143,In_972);
or U679 (N_679,In_502,In_567);
nor U680 (N_680,In_29,In_980);
xor U681 (N_681,In_523,In_660);
nor U682 (N_682,In_644,In_56);
and U683 (N_683,In_765,In_806);
and U684 (N_684,In_849,In_396);
nor U685 (N_685,In_787,In_647);
and U686 (N_686,In_285,In_855);
or U687 (N_687,In_174,In_411);
and U688 (N_688,In_955,In_339);
xor U689 (N_689,In_121,In_635);
and U690 (N_690,In_491,In_403);
nand U691 (N_691,In_360,In_609);
xnor U692 (N_692,In_476,In_754);
and U693 (N_693,In_954,In_495);
or U694 (N_694,In_724,In_14);
xor U695 (N_695,In_801,In_586);
or U696 (N_696,In_804,In_64);
and U697 (N_697,In_626,In_58);
nand U698 (N_698,In_880,In_950);
or U699 (N_699,In_28,In_126);
nand U700 (N_700,In_25,In_913);
nor U701 (N_701,In_267,In_596);
and U702 (N_702,In_875,In_664);
nor U703 (N_703,In_377,In_196);
nor U704 (N_704,In_155,In_346);
xor U705 (N_705,In_22,In_502);
or U706 (N_706,In_264,In_561);
or U707 (N_707,In_337,In_419);
or U708 (N_708,In_131,In_495);
and U709 (N_709,In_368,In_852);
and U710 (N_710,In_654,In_239);
or U711 (N_711,In_100,In_443);
xor U712 (N_712,In_461,In_913);
and U713 (N_713,In_612,In_288);
nand U714 (N_714,In_754,In_700);
and U715 (N_715,In_429,In_661);
and U716 (N_716,In_777,In_734);
nand U717 (N_717,In_150,In_998);
xor U718 (N_718,In_61,In_523);
nand U719 (N_719,In_101,In_867);
xor U720 (N_720,In_815,In_563);
xor U721 (N_721,In_117,In_601);
nand U722 (N_722,In_886,In_354);
or U723 (N_723,In_451,In_607);
or U724 (N_724,In_536,In_500);
and U725 (N_725,In_942,In_205);
xor U726 (N_726,In_684,In_235);
xnor U727 (N_727,In_126,In_903);
xor U728 (N_728,In_573,In_271);
nand U729 (N_729,In_177,In_172);
nor U730 (N_730,In_337,In_278);
nand U731 (N_731,In_19,In_95);
nor U732 (N_732,In_245,In_592);
and U733 (N_733,In_548,In_758);
xor U734 (N_734,In_992,In_828);
or U735 (N_735,In_647,In_387);
nor U736 (N_736,In_902,In_890);
nand U737 (N_737,In_37,In_678);
or U738 (N_738,In_293,In_764);
and U739 (N_739,In_492,In_141);
xnor U740 (N_740,In_712,In_612);
nand U741 (N_741,In_808,In_478);
nand U742 (N_742,In_674,In_969);
and U743 (N_743,In_686,In_176);
nand U744 (N_744,In_464,In_886);
or U745 (N_745,In_877,In_81);
nand U746 (N_746,In_956,In_487);
xor U747 (N_747,In_792,In_640);
or U748 (N_748,In_539,In_431);
and U749 (N_749,In_451,In_438);
xor U750 (N_750,In_132,In_643);
xnor U751 (N_751,In_926,In_228);
nand U752 (N_752,In_157,In_998);
xnor U753 (N_753,In_803,In_161);
and U754 (N_754,In_173,In_444);
and U755 (N_755,In_230,In_943);
or U756 (N_756,In_628,In_25);
nand U757 (N_757,In_432,In_365);
and U758 (N_758,In_374,In_10);
or U759 (N_759,In_404,In_966);
xnor U760 (N_760,In_300,In_516);
and U761 (N_761,In_73,In_346);
nand U762 (N_762,In_873,In_19);
or U763 (N_763,In_598,In_194);
or U764 (N_764,In_489,In_422);
nand U765 (N_765,In_396,In_905);
or U766 (N_766,In_545,In_661);
nor U767 (N_767,In_744,In_556);
and U768 (N_768,In_158,In_619);
and U769 (N_769,In_204,In_722);
nand U770 (N_770,In_384,In_532);
nand U771 (N_771,In_964,In_110);
or U772 (N_772,In_53,In_950);
nand U773 (N_773,In_538,In_972);
nand U774 (N_774,In_723,In_68);
nand U775 (N_775,In_217,In_980);
or U776 (N_776,In_162,In_110);
and U777 (N_777,In_433,In_88);
nor U778 (N_778,In_682,In_160);
and U779 (N_779,In_794,In_387);
xnor U780 (N_780,In_225,In_16);
nand U781 (N_781,In_634,In_673);
or U782 (N_782,In_987,In_233);
nor U783 (N_783,In_979,In_788);
xor U784 (N_784,In_123,In_565);
xor U785 (N_785,In_543,In_540);
and U786 (N_786,In_377,In_69);
nor U787 (N_787,In_364,In_703);
nand U788 (N_788,In_949,In_74);
and U789 (N_789,In_344,In_725);
nor U790 (N_790,In_937,In_863);
xor U791 (N_791,In_917,In_837);
nor U792 (N_792,In_875,In_585);
and U793 (N_793,In_622,In_337);
or U794 (N_794,In_506,In_454);
nand U795 (N_795,In_409,In_780);
or U796 (N_796,In_529,In_133);
xor U797 (N_797,In_286,In_804);
xnor U798 (N_798,In_808,In_633);
nor U799 (N_799,In_164,In_188);
and U800 (N_800,In_587,In_418);
and U801 (N_801,In_101,In_506);
nor U802 (N_802,In_805,In_103);
xor U803 (N_803,In_287,In_895);
or U804 (N_804,In_597,In_63);
and U805 (N_805,In_70,In_368);
nand U806 (N_806,In_926,In_120);
nand U807 (N_807,In_142,In_434);
nor U808 (N_808,In_667,In_438);
nand U809 (N_809,In_413,In_550);
or U810 (N_810,In_863,In_924);
nand U811 (N_811,In_428,In_220);
or U812 (N_812,In_594,In_40);
xor U813 (N_813,In_304,In_96);
and U814 (N_814,In_389,In_878);
nand U815 (N_815,In_303,In_137);
nor U816 (N_816,In_388,In_488);
or U817 (N_817,In_806,In_60);
xor U818 (N_818,In_553,In_969);
nor U819 (N_819,In_649,In_537);
or U820 (N_820,In_699,In_957);
nand U821 (N_821,In_354,In_609);
xor U822 (N_822,In_709,In_155);
xnor U823 (N_823,In_880,In_588);
or U824 (N_824,In_265,In_346);
or U825 (N_825,In_332,In_147);
and U826 (N_826,In_748,In_331);
xnor U827 (N_827,In_562,In_818);
nor U828 (N_828,In_572,In_350);
or U829 (N_829,In_138,In_178);
nor U830 (N_830,In_111,In_87);
nor U831 (N_831,In_658,In_70);
nand U832 (N_832,In_961,In_189);
nand U833 (N_833,In_341,In_37);
and U834 (N_834,In_934,In_654);
xor U835 (N_835,In_410,In_675);
and U836 (N_836,In_254,In_33);
xnor U837 (N_837,In_998,In_252);
and U838 (N_838,In_905,In_914);
or U839 (N_839,In_787,In_553);
nand U840 (N_840,In_367,In_821);
or U841 (N_841,In_523,In_98);
nor U842 (N_842,In_288,In_971);
nand U843 (N_843,In_672,In_353);
and U844 (N_844,In_771,In_743);
or U845 (N_845,In_242,In_432);
nand U846 (N_846,In_85,In_9);
or U847 (N_847,In_120,In_875);
nor U848 (N_848,In_586,In_50);
nand U849 (N_849,In_202,In_698);
or U850 (N_850,In_710,In_11);
or U851 (N_851,In_405,In_908);
and U852 (N_852,In_490,In_499);
and U853 (N_853,In_344,In_921);
nand U854 (N_854,In_375,In_128);
nand U855 (N_855,In_316,In_963);
xnor U856 (N_856,In_417,In_428);
and U857 (N_857,In_396,In_202);
or U858 (N_858,In_958,In_520);
nor U859 (N_859,In_994,In_159);
and U860 (N_860,In_500,In_440);
nand U861 (N_861,In_651,In_674);
nand U862 (N_862,In_362,In_466);
xor U863 (N_863,In_393,In_941);
xor U864 (N_864,In_369,In_909);
nand U865 (N_865,In_176,In_99);
nor U866 (N_866,In_464,In_880);
and U867 (N_867,In_848,In_454);
nand U868 (N_868,In_439,In_680);
or U869 (N_869,In_309,In_541);
or U870 (N_870,In_452,In_90);
or U871 (N_871,In_23,In_788);
or U872 (N_872,In_940,In_775);
nand U873 (N_873,In_359,In_53);
and U874 (N_874,In_489,In_945);
nor U875 (N_875,In_824,In_991);
or U876 (N_876,In_410,In_356);
or U877 (N_877,In_325,In_278);
nand U878 (N_878,In_81,In_125);
nor U879 (N_879,In_481,In_397);
nor U880 (N_880,In_13,In_107);
and U881 (N_881,In_824,In_275);
and U882 (N_882,In_643,In_364);
xnor U883 (N_883,In_538,In_362);
and U884 (N_884,In_292,In_206);
nand U885 (N_885,In_648,In_266);
xor U886 (N_886,In_621,In_247);
nand U887 (N_887,In_226,In_899);
nand U888 (N_888,In_996,In_912);
and U889 (N_889,In_93,In_433);
and U890 (N_890,In_686,In_410);
nor U891 (N_891,In_618,In_357);
xnor U892 (N_892,In_380,In_644);
or U893 (N_893,In_711,In_759);
and U894 (N_894,In_999,In_326);
xor U895 (N_895,In_27,In_703);
nand U896 (N_896,In_516,In_605);
nor U897 (N_897,In_296,In_882);
nor U898 (N_898,In_459,In_37);
nor U899 (N_899,In_369,In_239);
nor U900 (N_900,In_268,In_663);
nor U901 (N_901,In_525,In_758);
nor U902 (N_902,In_916,In_937);
nor U903 (N_903,In_185,In_528);
or U904 (N_904,In_444,In_912);
or U905 (N_905,In_956,In_210);
nand U906 (N_906,In_780,In_104);
and U907 (N_907,In_904,In_647);
and U908 (N_908,In_615,In_422);
nand U909 (N_909,In_507,In_454);
and U910 (N_910,In_470,In_93);
nand U911 (N_911,In_69,In_292);
or U912 (N_912,In_700,In_679);
or U913 (N_913,In_449,In_5);
nor U914 (N_914,In_468,In_655);
xor U915 (N_915,In_748,In_691);
nor U916 (N_916,In_563,In_99);
xnor U917 (N_917,In_888,In_734);
xnor U918 (N_918,In_301,In_541);
nand U919 (N_919,In_21,In_996);
or U920 (N_920,In_898,In_389);
and U921 (N_921,In_739,In_977);
or U922 (N_922,In_857,In_440);
xnor U923 (N_923,In_944,In_105);
nor U924 (N_924,In_967,In_727);
and U925 (N_925,In_259,In_995);
and U926 (N_926,In_138,In_134);
nand U927 (N_927,In_10,In_169);
nor U928 (N_928,In_797,In_869);
xnor U929 (N_929,In_922,In_297);
and U930 (N_930,In_996,In_196);
and U931 (N_931,In_44,In_301);
and U932 (N_932,In_336,In_309);
xor U933 (N_933,In_398,In_124);
or U934 (N_934,In_959,In_803);
nand U935 (N_935,In_479,In_208);
and U936 (N_936,In_66,In_471);
or U937 (N_937,In_462,In_911);
xor U938 (N_938,In_232,In_365);
nor U939 (N_939,In_242,In_357);
nor U940 (N_940,In_273,In_596);
or U941 (N_941,In_882,In_327);
and U942 (N_942,In_599,In_797);
nor U943 (N_943,In_691,In_959);
nand U944 (N_944,In_446,In_630);
xnor U945 (N_945,In_13,In_905);
and U946 (N_946,In_445,In_93);
xnor U947 (N_947,In_666,In_881);
nand U948 (N_948,In_490,In_242);
nand U949 (N_949,In_489,In_828);
or U950 (N_950,In_507,In_94);
or U951 (N_951,In_183,In_676);
xor U952 (N_952,In_609,In_449);
nor U953 (N_953,In_283,In_974);
xor U954 (N_954,In_911,In_114);
nand U955 (N_955,In_443,In_264);
and U956 (N_956,In_301,In_323);
nand U957 (N_957,In_49,In_796);
nand U958 (N_958,In_175,In_385);
nand U959 (N_959,In_356,In_988);
nor U960 (N_960,In_599,In_246);
nand U961 (N_961,In_41,In_642);
or U962 (N_962,In_555,In_618);
nor U963 (N_963,In_795,In_540);
or U964 (N_964,In_227,In_725);
nand U965 (N_965,In_93,In_802);
nor U966 (N_966,In_403,In_561);
nor U967 (N_967,In_351,In_864);
nand U968 (N_968,In_254,In_73);
and U969 (N_969,In_737,In_537);
or U970 (N_970,In_93,In_88);
or U971 (N_971,In_768,In_216);
xor U972 (N_972,In_410,In_183);
nand U973 (N_973,In_499,In_221);
nor U974 (N_974,In_687,In_117);
xor U975 (N_975,In_715,In_829);
nor U976 (N_976,In_121,In_127);
or U977 (N_977,In_572,In_261);
nor U978 (N_978,In_663,In_259);
nor U979 (N_979,In_27,In_887);
nand U980 (N_980,In_270,In_646);
and U981 (N_981,In_44,In_659);
or U982 (N_982,In_506,In_180);
nor U983 (N_983,In_304,In_545);
and U984 (N_984,In_245,In_285);
xor U985 (N_985,In_889,In_110);
or U986 (N_986,In_364,In_811);
and U987 (N_987,In_368,In_34);
xnor U988 (N_988,In_76,In_516);
and U989 (N_989,In_104,In_867);
or U990 (N_990,In_125,In_513);
xor U991 (N_991,In_641,In_153);
nand U992 (N_992,In_673,In_75);
nor U993 (N_993,In_733,In_364);
and U994 (N_994,In_977,In_710);
nor U995 (N_995,In_732,In_831);
nor U996 (N_996,In_962,In_777);
nand U997 (N_997,In_322,In_700);
nor U998 (N_998,In_776,In_307);
nor U999 (N_999,In_870,In_268);
xor U1000 (N_1000,N_426,N_923);
xnor U1001 (N_1001,N_585,N_641);
or U1002 (N_1002,N_770,N_237);
and U1003 (N_1003,N_971,N_69);
xnor U1004 (N_1004,N_310,N_706);
nand U1005 (N_1005,N_647,N_338);
or U1006 (N_1006,N_775,N_672);
nand U1007 (N_1007,N_262,N_528);
or U1008 (N_1008,N_210,N_83);
nand U1009 (N_1009,N_625,N_119);
and U1010 (N_1010,N_140,N_70);
xor U1011 (N_1011,N_193,N_747);
or U1012 (N_1012,N_78,N_959);
nand U1013 (N_1013,N_243,N_912);
xnor U1014 (N_1014,N_392,N_0);
xor U1015 (N_1015,N_280,N_578);
nand U1016 (N_1016,N_963,N_900);
xnor U1017 (N_1017,N_327,N_571);
and U1018 (N_1018,N_487,N_254);
nand U1019 (N_1019,N_395,N_544);
xnor U1020 (N_1020,N_215,N_635);
nand U1021 (N_1021,N_9,N_835);
xor U1022 (N_1022,N_199,N_377);
or U1023 (N_1023,N_779,N_349);
and U1024 (N_1024,N_823,N_861);
nand U1025 (N_1025,N_208,N_686);
nand U1026 (N_1026,N_153,N_333);
or U1027 (N_1027,N_159,N_227);
or U1028 (N_1028,N_760,N_551);
and U1029 (N_1029,N_359,N_548);
and U1030 (N_1030,N_86,N_356);
or U1031 (N_1031,N_555,N_54);
xnor U1032 (N_1032,N_462,N_320);
nor U1033 (N_1033,N_977,N_894);
nor U1034 (N_1034,N_344,N_231);
nand U1035 (N_1035,N_51,N_309);
or U1036 (N_1036,N_476,N_577);
and U1037 (N_1037,N_403,N_61);
or U1038 (N_1038,N_794,N_157);
nand U1039 (N_1039,N_351,N_347);
xor U1040 (N_1040,N_37,N_474);
xor U1041 (N_1041,N_965,N_873);
and U1042 (N_1042,N_658,N_903);
xor U1043 (N_1043,N_381,N_465);
nand U1044 (N_1044,N_650,N_855);
and U1045 (N_1045,N_205,N_366);
or U1046 (N_1046,N_717,N_987);
xor U1047 (N_1047,N_453,N_557);
nor U1048 (N_1048,N_224,N_492);
nor U1049 (N_1049,N_608,N_530);
nand U1050 (N_1050,N_270,N_1);
and U1051 (N_1051,N_568,N_122);
xnor U1052 (N_1052,N_805,N_979);
nor U1053 (N_1053,N_33,N_831);
and U1054 (N_1054,N_564,N_216);
and U1055 (N_1055,N_287,N_284);
and U1056 (N_1056,N_456,N_917);
xnor U1057 (N_1057,N_891,N_135);
and U1058 (N_1058,N_107,N_168);
nand U1059 (N_1059,N_605,N_631);
and U1060 (N_1060,N_670,N_689);
and U1061 (N_1061,N_793,N_459);
nand U1062 (N_1062,N_654,N_211);
nand U1063 (N_1063,N_16,N_429);
and U1064 (N_1064,N_316,N_245);
or U1065 (N_1065,N_758,N_265);
or U1066 (N_1066,N_713,N_525);
xor U1067 (N_1067,N_276,N_685);
or U1068 (N_1068,N_537,N_506);
xnor U1069 (N_1069,N_481,N_936);
nor U1070 (N_1070,N_125,N_897);
xnor U1071 (N_1071,N_712,N_859);
or U1072 (N_1072,N_606,N_680);
or U1073 (N_1073,N_961,N_597);
and U1074 (N_1074,N_81,N_782);
nand U1075 (N_1075,N_445,N_498);
or U1076 (N_1076,N_688,N_721);
and U1077 (N_1077,N_534,N_306);
and U1078 (N_1078,N_454,N_348);
and U1079 (N_1079,N_129,N_192);
and U1080 (N_1080,N_136,N_709);
or U1081 (N_1081,N_165,N_698);
and U1082 (N_1082,N_504,N_870);
xor U1083 (N_1083,N_879,N_217);
nor U1084 (N_1084,N_575,N_632);
xnor U1085 (N_1085,N_483,N_353);
and U1086 (N_1086,N_74,N_708);
nor U1087 (N_1087,N_864,N_666);
and U1088 (N_1088,N_375,N_693);
nand U1089 (N_1089,N_82,N_194);
nor U1090 (N_1090,N_535,N_253);
nand U1091 (N_1091,N_704,N_98);
and U1092 (N_1092,N_120,N_479);
or U1093 (N_1093,N_662,N_300);
and U1094 (N_1094,N_840,N_540);
nor U1095 (N_1095,N_803,N_931);
or U1096 (N_1096,N_892,N_679);
nor U1097 (N_1097,N_77,N_640);
nand U1098 (N_1098,N_991,N_878);
or U1099 (N_1099,N_602,N_437);
nand U1100 (N_1100,N_185,N_556);
nor U1101 (N_1101,N_108,N_390);
nor U1102 (N_1102,N_281,N_282);
or U1103 (N_1103,N_186,N_283);
nor U1104 (N_1104,N_611,N_370);
xor U1105 (N_1105,N_110,N_567);
and U1106 (N_1106,N_66,N_893);
nand U1107 (N_1107,N_741,N_142);
nand U1108 (N_1108,N_363,N_905);
nor U1109 (N_1109,N_545,N_410);
nand U1110 (N_1110,N_887,N_671);
and U1111 (N_1111,N_79,N_695);
or U1112 (N_1112,N_862,N_21);
nand U1113 (N_1113,N_612,N_924);
or U1114 (N_1114,N_178,N_497);
nand U1115 (N_1115,N_304,N_19);
and U1116 (N_1116,N_49,N_984);
and U1117 (N_1117,N_649,N_702);
nor U1118 (N_1118,N_983,N_179);
or U1119 (N_1119,N_720,N_251);
xor U1120 (N_1120,N_357,N_990);
xor U1121 (N_1121,N_238,N_885);
or U1122 (N_1122,N_904,N_967);
nor U1123 (N_1123,N_371,N_918);
or U1124 (N_1124,N_11,N_810);
nand U1125 (N_1125,N_6,N_895);
nor U1126 (N_1126,N_188,N_549);
xor U1127 (N_1127,N_707,N_538);
or U1128 (N_1128,N_778,N_152);
xnor U1129 (N_1129,N_952,N_146);
xor U1130 (N_1130,N_814,N_527);
nor U1131 (N_1131,N_560,N_850);
xnor U1132 (N_1132,N_723,N_774);
nand U1133 (N_1133,N_547,N_313);
or U1134 (N_1134,N_875,N_500);
nor U1135 (N_1135,N_854,N_884);
and U1136 (N_1136,N_232,N_415);
nand U1137 (N_1137,N_665,N_992);
nand U1138 (N_1138,N_522,N_235);
nand U1139 (N_1139,N_920,N_834);
nand U1140 (N_1140,N_75,N_446);
nand U1141 (N_1141,N_113,N_801);
and U1142 (N_1142,N_826,N_480);
or U1143 (N_1143,N_439,N_112);
or U1144 (N_1144,N_323,N_105);
and U1145 (N_1145,N_123,N_914);
nor U1146 (N_1146,N_8,N_674);
or U1147 (N_1147,N_218,N_877);
xor U1148 (N_1148,N_43,N_729);
nor U1149 (N_1149,N_566,N_2);
nand U1150 (N_1150,N_792,N_493);
nor U1151 (N_1151,N_812,N_268);
nand U1152 (N_1152,N_223,N_418);
nor U1153 (N_1153,N_876,N_848);
nor U1154 (N_1154,N_334,N_956);
nand U1155 (N_1155,N_394,N_24);
nor U1156 (N_1156,N_501,N_815);
nor U1157 (N_1157,N_329,N_833);
xor U1158 (N_1158,N_841,N_962);
nand U1159 (N_1159,N_511,N_637);
xor U1160 (N_1160,N_749,N_807);
nand U1161 (N_1161,N_628,N_63);
and U1162 (N_1162,N_190,N_145);
xnor U1163 (N_1163,N_633,N_378);
nor U1164 (N_1164,N_646,N_790);
and U1165 (N_1165,N_246,N_572);
and U1166 (N_1166,N_412,N_350);
xnor U1167 (N_1167,N_407,N_839);
or U1168 (N_1168,N_594,N_935);
nand U1169 (N_1169,N_402,N_328);
nor U1170 (N_1170,N_554,N_871);
xnor U1171 (N_1171,N_851,N_288);
xnor U1172 (N_1172,N_322,N_89);
or U1173 (N_1173,N_582,N_523);
and U1174 (N_1174,N_467,N_408);
nand U1175 (N_1175,N_198,N_664);
xor U1176 (N_1176,N_14,N_922);
xnor U1177 (N_1177,N_71,N_659);
xnor U1178 (N_1178,N_515,N_62);
and U1179 (N_1179,N_667,N_700);
nand U1180 (N_1180,N_425,N_907);
nand U1181 (N_1181,N_899,N_845);
nand U1182 (N_1182,N_274,N_824);
nand U1183 (N_1183,N_913,N_393);
and U1184 (N_1184,N_960,N_431);
nor U1185 (N_1185,N_951,N_844);
xor U1186 (N_1186,N_85,N_417);
nand U1187 (N_1187,N_180,N_590);
nand U1188 (N_1188,N_367,N_289);
and U1189 (N_1189,N_463,N_99);
nor U1190 (N_1190,N_336,N_266);
xor U1191 (N_1191,N_273,N_451);
or U1192 (N_1192,N_829,N_822);
and U1193 (N_1193,N_365,N_745);
and U1194 (N_1194,N_669,N_277);
xnor U1195 (N_1195,N_94,N_644);
nand U1196 (N_1196,N_10,N_312);
nand U1197 (N_1197,N_615,N_499);
xor U1198 (N_1198,N_624,N_653);
nor U1199 (N_1199,N_28,N_795);
xnor U1200 (N_1200,N_255,N_295);
nand U1201 (N_1201,N_678,N_989);
nor U1202 (N_1202,N_259,N_866);
and U1203 (N_1203,N_648,N_477);
and U1204 (N_1204,N_837,N_380);
or U1205 (N_1205,N_318,N_342);
and U1206 (N_1206,N_733,N_627);
and U1207 (N_1207,N_128,N_233);
nor U1208 (N_1208,N_716,N_55);
nor U1209 (N_1209,N_17,N_638);
nor U1210 (N_1210,N_311,N_789);
nand U1211 (N_1211,N_915,N_888);
or U1212 (N_1212,N_710,N_532);
nand U1213 (N_1213,N_604,N_67);
xnor U1214 (N_1214,N_818,N_516);
xor U1215 (N_1215,N_106,N_821);
and U1216 (N_1216,N_470,N_746);
nor U1217 (N_1217,N_673,N_943);
nor U1218 (N_1218,N_734,N_744);
or U1219 (N_1219,N_510,N_561);
and U1220 (N_1220,N_214,N_59);
xnor U1221 (N_1221,N_502,N_396);
nand U1222 (N_1222,N_26,N_175);
xor U1223 (N_1223,N_763,N_229);
xor U1224 (N_1224,N_932,N_315);
nor U1225 (N_1225,N_278,N_44);
nor U1226 (N_1226,N_852,N_642);
xor U1227 (N_1227,N_629,N_292);
nor U1228 (N_1228,N_491,N_221);
nor U1229 (N_1229,N_41,N_297);
nand U1230 (N_1230,N_47,N_101);
or U1231 (N_1231,N_427,N_768);
and U1232 (N_1232,N_222,N_738);
nor U1233 (N_1233,N_847,N_23);
nor U1234 (N_1234,N_676,N_442);
xor U1235 (N_1235,N_766,N_996);
nor U1236 (N_1236,N_452,N_409);
or U1237 (N_1237,N_7,N_589);
or U1238 (N_1238,N_569,N_387);
or U1239 (N_1239,N_335,N_869);
xor U1240 (N_1240,N_27,N_405);
and U1241 (N_1241,N_668,N_937);
nor U1242 (N_1242,N_986,N_478);
nand U1243 (N_1243,N_115,N_727);
or U1244 (N_1244,N_326,N_767);
nand U1245 (N_1245,N_660,N_574);
and U1246 (N_1246,N_958,N_406);
or U1247 (N_1247,N_724,N_111);
and U1248 (N_1248,N_754,N_154);
or U1249 (N_1249,N_969,N_539);
xnor U1250 (N_1250,N_621,N_882);
xnor U1251 (N_1251,N_401,N_583);
and U1252 (N_1252,N_505,N_250);
nand U1253 (N_1253,N_374,N_189);
nand U1254 (N_1254,N_469,N_360);
xnor U1255 (N_1255,N_677,N_715);
nand U1256 (N_1256,N_422,N_182);
or U1257 (N_1257,N_966,N_331);
xor U1258 (N_1258,N_441,N_519);
xor U1259 (N_1259,N_118,N_22);
and U1260 (N_1260,N_60,N_430);
and U1261 (N_1261,N_619,N_683);
xor U1262 (N_1262,N_620,N_457);
xnor U1263 (N_1263,N_939,N_448);
nor U1264 (N_1264,N_865,N_204);
and U1265 (N_1265,N_234,N_562);
and U1266 (N_1266,N_80,N_352);
and U1267 (N_1267,N_581,N_843);
and U1268 (N_1268,N_933,N_132);
nor U1269 (N_1269,N_161,N_616);
nor U1270 (N_1270,N_225,N_368);
nor U1271 (N_1271,N_719,N_35);
and U1272 (N_1272,N_432,N_414);
nand U1273 (N_1273,N_298,N_813);
and U1274 (N_1274,N_275,N_764);
xnor U1275 (N_1275,N_114,N_65);
xnor U1276 (N_1276,N_319,N_880);
nand U1277 (N_1277,N_771,N_769);
or U1278 (N_1278,N_472,N_379);
xnor U1279 (N_1279,N_898,N_603);
xnor U1280 (N_1280,N_345,N_308);
and U1281 (N_1281,N_696,N_264);
and U1282 (N_1282,N_346,N_927);
xor U1283 (N_1283,N_141,N_599);
xnor U1284 (N_1284,N_321,N_906);
nor U1285 (N_1285,N_985,N_711);
or U1286 (N_1286,N_860,N_692);
or U1287 (N_1287,N_699,N_748);
xnor U1288 (N_1288,N_701,N_202);
nand U1289 (N_1289,N_925,N_187);
or U1290 (N_1290,N_765,N_400);
xnor U1291 (N_1291,N_520,N_388);
and U1292 (N_1292,N_751,N_543);
nor U1293 (N_1293,N_240,N_798);
nor U1294 (N_1294,N_656,N_513);
xor U1295 (N_1295,N_4,N_750);
xor U1296 (N_1296,N_171,N_314);
xnor U1297 (N_1297,N_421,N_389);
nor U1298 (N_1298,N_718,N_916);
nand U1299 (N_1299,N_20,N_832);
nor U1300 (N_1300,N_87,N_76);
nor U1301 (N_1301,N_858,N_148);
xnor U1302 (N_1302,N_438,N_58);
and U1303 (N_1303,N_868,N_116);
nor U1304 (N_1304,N_15,N_303);
xnor U1305 (N_1305,N_397,N_435);
and U1306 (N_1306,N_271,N_138);
and U1307 (N_1307,N_294,N_518);
nor U1308 (N_1308,N_596,N_39);
nor U1309 (N_1309,N_941,N_974);
or U1310 (N_1310,N_325,N_428);
xor U1311 (N_1311,N_970,N_299);
nor U1312 (N_1312,N_220,N_53);
nand U1313 (N_1313,N_496,N_489);
nand U1314 (N_1314,N_610,N_420);
xor U1315 (N_1315,N_507,N_836);
nand U1316 (N_1316,N_601,N_780);
nand U1317 (N_1317,N_291,N_819);
nor U1318 (N_1318,N_12,N_607);
or U1319 (N_1319,N_732,N_736);
nor U1320 (N_1320,N_170,N_143);
nor U1321 (N_1321,N_372,N_296);
nor U1322 (N_1322,N_846,N_752);
xor U1323 (N_1323,N_928,N_946);
nor U1324 (N_1324,N_443,N_48);
or U1325 (N_1325,N_761,N_68);
or U1326 (N_1326,N_816,N_163);
xor U1327 (N_1327,N_285,N_100);
nand U1328 (N_1328,N_286,N_293);
nor U1329 (N_1329,N_173,N_784);
xnor U1330 (N_1330,N_881,N_570);
and U1331 (N_1331,N_383,N_827);
nor U1332 (N_1332,N_639,N_503);
and U1333 (N_1333,N_623,N_473);
or U1334 (N_1334,N_384,N_485);
xnor U1335 (N_1335,N_584,N_301);
nor U1336 (N_1336,N_484,N_30);
nand U1337 (N_1337,N_825,N_757);
or U1338 (N_1338,N_651,N_64);
or U1339 (N_1339,N_137,N_791);
nor U1340 (N_1340,N_867,N_18);
nor U1341 (N_1341,N_96,N_740);
nor U1342 (N_1342,N_684,N_786);
xor U1343 (N_1343,N_756,N_863);
or U1344 (N_1344,N_995,N_226);
or U1345 (N_1345,N_697,N_104);
or U1346 (N_1346,N_842,N_948);
xnor U1347 (N_1347,N_725,N_109);
nand U1348 (N_1348,N_200,N_743);
nor U1349 (N_1349,N_25,N_514);
nor U1350 (N_1350,N_52,N_447);
nor U1351 (N_1351,N_942,N_130);
nor U1352 (N_1352,N_126,N_978);
nor U1353 (N_1353,N_636,N_46);
or U1354 (N_1354,N_509,N_358);
or U1355 (N_1355,N_341,N_926);
or U1356 (N_1356,N_444,N_460);
and U1357 (N_1357,N_468,N_434);
xnor U1358 (N_1358,N_391,N_626);
or U1359 (N_1359,N_901,N_339);
xnor U1360 (N_1360,N_808,N_531);
nand U1361 (N_1361,N_177,N_207);
and U1362 (N_1362,N_994,N_828);
nor U1363 (N_1363,N_703,N_797);
xnor U1364 (N_1364,N_964,N_455);
nor U1365 (N_1365,N_645,N_183);
nand U1366 (N_1366,N_973,N_279);
and U1367 (N_1367,N_102,N_436);
and U1368 (N_1368,N_919,N_737);
nor U1369 (N_1369,N_124,N_369);
or U1370 (N_1370,N_800,N_934);
or U1371 (N_1371,N_890,N_643);
xnor U1372 (N_1372,N_248,N_482);
nor U1373 (N_1373,N_988,N_340);
or U1374 (N_1374,N_3,N_411);
xor U1375 (N_1375,N_857,N_413);
or U1376 (N_1376,N_600,N_849);
and U1377 (N_1377,N_36,N_305);
nor U1378 (N_1378,N_464,N_630);
nand U1379 (N_1379,N_362,N_526);
or U1380 (N_1380,N_853,N_586);
or U1381 (N_1381,N_576,N_546);
and U1382 (N_1382,N_458,N_373);
or U1383 (N_1383,N_197,N_993);
nand U1384 (N_1384,N_486,N_386);
and U1385 (N_1385,N_239,N_999);
nand U1386 (N_1386,N_663,N_617);
nor U1387 (N_1387,N_728,N_419);
nor U1388 (N_1388,N_799,N_38);
nand U1389 (N_1389,N_802,N_31);
or U1390 (N_1390,N_595,N_587);
or U1391 (N_1391,N_954,N_598);
xnor U1392 (N_1392,N_921,N_34);
and U1393 (N_1393,N_755,N_263);
nand U1394 (N_1394,N_440,N_290);
and U1395 (N_1395,N_127,N_950);
or U1396 (N_1396,N_559,N_886);
and U1397 (N_1397,N_343,N_252);
nand U1398 (N_1398,N_156,N_45);
nor U1399 (N_1399,N_260,N_133);
nand U1400 (N_1400,N_158,N_622);
and U1401 (N_1401,N_675,N_788);
xor U1402 (N_1402,N_772,N_57);
nand U1403 (N_1403,N_247,N_940);
nor U1404 (N_1404,N_687,N_195);
or U1405 (N_1405,N_817,N_258);
xor U1406 (N_1406,N_50,N_657);
or U1407 (N_1407,N_206,N_166);
and U1408 (N_1408,N_257,N_307);
nand U1409 (N_1409,N_196,N_242);
xnor U1410 (N_1410,N_521,N_730);
nand U1411 (N_1411,N_785,N_953);
xnor U1412 (N_1412,N_781,N_416);
nand U1413 (N_1413,N_618,N_139);
and U1414 (N_1414,N_42,N_488);
or U1415 (N_1415,N_580,N_889);
nand U1416 (N_1416,N_512,N_261);
nand U1417 (N_1417,N_471,N_806);
xor U1418 (N_1418,N_976,N_466);
or U1419 (N_1419,N_524,N_144);
and U1420 (N_1420,N_324,N_376);
and U1421 (N_1421,N_883,N_552);
or U1422 (N_1422,N_694,N_796);
and U1423 (N_1423,N_404,N_475);
nor U1424 (N_1424,N_90,N_655);
nand U1425 (N_1425,N_783,N_553);
nand U1426 (N_1426,N_731,N_423);
or U1427 (N_1427,N_944,N_614);
and U1428 (N_1428,N_588,N_579);
xor U1429 (N_1429,N_981,N_980);
nand U1430 (N_1430,N_73,N_735);
or U1431 (N_1431,N_330,N_820);
or U1432 (N_1432,N_955,N_661);
and U1433 (N_1433,N_201,N_896);
nor U1434 (N_1434,N_149,N_908);
and U1435 (N_1435,N_541,N_508);
nor U1436 (N_1436,N_529,N_609);
or U1437 (N_1437,N_563,N_212);
or U1438 (N_1438,N_911,N_929);
nor U1439 (N_1439,N_164,N_29);
or U1440 (N_1440,N_147,N_691);
xor U1441 (N_1441,N_150,N_722);
nand U1442 (N_1442,N_830,N_84);
and U1443 (N_1443,N_753,N_241);
nand U1444 (N_1444,N_236,N_681);
and U1445 (N_1445,N_998,N_317);
nand U1446 (N_1446,N_181,N_13);
xor U1447 (N_1447,N_167,N_162);
xnor U1448 (N_1448,N_997,N_909);
or U1449 (N_1449,N_424,N_949);
nand U1450 (N_1450,N_490,N_945);
or U1451 (N_1451,N_968,N_573);
xnor U1452 (N_1452,N_874,N_856);
or U1453 (N_1453,N_495,N_726);
nand U1454 (N_1454,N_209,N_219);
or U1455 (N_1455,N_902,N_652);
nand U1456 (N_1456,N_256,N_382);
and U1457 (N_1457,N_714,N_385);
nor U1458 (N_1458,N_244,N_355);
or U1459 (N_1459,N_361,N_947);
and U1460 (N_1460,N_450,N_494);
nand U1461 (N_1461,N_776,N_174);
or U1462 (N_1462,N_131,N_364);
or U1463 (N_1463,N_982,N_809);
or U1464 (N_1464,N_176,N_739);
nor U1465 (N_1465,N_91,N_267);
xor U1466 (N_1466,N_705,N_591);
or U1467 (N_1467,N_593,N_32);
or U1468 (N_1468,N_461,N_172);
xor U1469 (N_1469,N_203,N_930);
nand U1470 (N_1470,N_742,N_533);
nand U1471 (N_1471,N_56,N_88);
nand U1472 (N_1472,N_759,N_938);
nand U1473 (N_1473,N_399,N_184);
and U1474 (N_1474,N_558,N_269);
and U1475 (N_1475,N_337,N_40);
nand U1476 (N_1476,N_213,N_634);
and U1477 (N_1477,N_592,N_160);
nand U1478 (N_1478,N_302,N_169);
nand U1479 (N_1479,N_804,N_230);
xor U1480 (N_1480,N_134,N_517);
nand U1481 (N_1481,N_272,N_5);
nor U1482 (N_1482,N_762,N_690);
and U1483 (N_1483,N_191,N_151);
and U1484 (N_1484,N_332,N_682);
xor U1485 (N_1485,N_975,N_536);
and U1486 (N_1486,N_542,N_228);
nand U1487 (N_1487,N_354,N_249);
xor U1488 (N_1488,N_550,N_773);
or U1489 (N_1489,N_910,N_838);
nand U1490 (N_1490,N_872,N_92);
or U1491 (N_1491,N_777,N_72);
xnor U1492 (N_1492,N_972,N_117);
nand U1493 (N_1493,N_398,N_93);
xor U1494 (N_1494,N_121,N_103);
nand U1495 (N_1495,N_433,N_613);
or U1496 (N_1496,N_787,N_449);
and U1497 (N_1497,N_811,N_95);
nor U1498 (N_1498,N_957,N_565);
xnor U1499 (N_1499,N_97,N_155);
nor U1500 (N_1500,N_637,N_103);
or U1501 (N_1501,N_39,N_718);
nor U1502 (N_1502,N_944,N_843);
and U1503 (N_1503,N_537,N_158);
or U1504 (N_1504,N_442,N_170);
nor U1505 (N_1505,N_38,N_371);
and U1506 (N_1506,N_219,N_437);
nor U1507 (N_1507,N_8,N_454);
xnor U1508 (N_1508,N_358,N_366);
xnor U1509 (N_1509,N_729,N_550);
nand U1510 (N_1510,N_272,N_416);
nand U1511 (N_1511,N_464,N_914);
nor U1512 (N_1512,N_98,N_556);
or U1513 (N_1513,N_3,N_800);
xnor U1514 (N_1514,N_384,N_109);
or U1515 (N_1515,N_418,N_47);
nand U1516 (N_1516,N_459,N_934);
nor U1517 (N_1517,N_281,N_602);
nand U1518 (N_1518,N_702,N_176);
xnor U1519 (N_1519,N_679,N_105);
xnor U1520 (N_1520,N_216,N_85);
or U1521 (N_1521,N_214,N_800);
nand U1522 (N_1522,N_815,N_556);
or U1523 (N_1523,N_736,N_299);
nand U1524 (N_1524,N_9,N_867);
xor U1525 (N_1525,N_407,N_63);
nor U1526 (N_1526,N_41,N_305);
xor U1527 (N_1527,N_528,N_239);
nand U1528 (N_1528,N_424,N_37);
and U1529 (N_1529,N_24,N_337);
nand U1530 (N_1530,N_733,N_822);
nor U1531 (N_1531,N_793,N_156);
or U1532 (N_1532,N_27,N_371);
nor U1533 (N_1533,N_110,N_537);
xor U1534 (N_1534,N_591,N_878);
xnor U1535 (N_1535,N_136,N_44);
nor U1536 (N_1536,N_548,N_303);
or U1537 (N_1537,N_851,N_168);
nand U1538 (N_1538,N_583,N_100);
xor U1539 (N_1539,N_31,N_928);
nor U1540 (N_1540,N_721,N_459);
xor U1541 (N_1541,N_514,N_659);
nor U1542 (N_1542,N_765,N_673);
nand U1543 (N_1543,N_561,N_926);
xor U1544 (N_1544,N_35,N_258);
nand U1545 (N_1545,N_266,N_338);
or U1546 (N_1546,N_669,N_748);
nor U1547 (N_1547,N_391,N_107);
and U1548 (N_1548,N_553,N_462);
nand U1549 (N_1549,N_149,N_860);
or U1550 (N_1550,N_918,N_461);
xnor U1551 (N_1551,N_678,N_42);
or U1552 (N_1552,N_771,N_882);
or U1553 (N_1553,N_194,N_928);
nor U1554 (N_1554,N_621,N_551);
and U1555 (N_1555,N_967,N_469);
or U1556 (N_1556,N_74,N_388);
or U1557 (N_1557,N_5,N_576);
nand U1558 (N_1558,N_943,N_355);
nand U1559 (N_1559,N_208,N_294);
nor U1560 (N_1560,N_151,N_177);
xor U1561 (N_1561,N_485,N_231);
and U1562 (N_1562,N_694,N_109);
nor U1563 (N_1563,N_617,N_493);
and U1564 (N_1564,N_546,N_977);
nor U1565 (N_1565,N_775,N_648);
xnor U1566 (N_1566,N_157,N_445);
and U1567 (N_1567,N_490,N_652);
or U1568 (N_1568,N_374,N_489);
nor U1569 (N_1569,N_221,N_601);
xnor U1570 (N_1570,N_366,N_226);
and U1571 (N_1571,N_262,N_610);
or U1572 (N_1572,N_58,N_913);
or U1573 (N_1573,N_204,N_425);
nor U1574 (N_1574,N_820,N_767);
nand U1575 (N_1575,N_729,N_436);
nor U1576 (N_1576,N_808,N_335);
and U1577 (N_1577,N_539,N_581);
nand U1578 (N_1578,N_894,N_616);
and U1579 (N_1579,N_832,N_135);
nor U1580 (N_1580,N_954,N_12);
xnor U1581 (N_1581,N_544,N_870);
xor U1582 (N_1582,N_684,N_96);
and U1583 (N_1583,N_451,N_620);
nor U1584 (N_1584,N_542,N_117);
nor U1585 (N_1585,N_363,N_92);
and U1586 (N_1586,N_966,N_530);
or U1587 (N_1587,N_830,N_905);
or U1588 (N_1588,N_206,N_534);
nor U1589 (N_1589,N_568,N_418);
nand U1590 (N_1590,N_921,N_366);
and U1591 (N_1591,N_510,N_652);
xor U1592 (N_1592,N_14,N_618);
and U1593 (N_1593,N_136,N_886);
xor U1594 (N_1594,N_753,N_546);
and U1595 (N_1595,N_725,N_359);
and U1596 (N_1596,N_120,N_957);
nand U1597 (N_1597,N_641,N_805);
xnor U1598 (N_1598,N_722,N_315);
and U1599 (N_1599,N_335,N_978);
and U1600 (N_1600,N_178,N_626);
nand U1601 (N_1601,N_554,N_827);
nand U1602 (N_1602,N_913,N_307);
nor U1603 (N_1603,N_141,N_912);
nand U1604 (N_1604,N_356,N_608);
xor U1605 (N_1605,N_879,N_776);
nand U1606 (N_1606,N_115,N_219);
xnor U1607 (N_1607,N_61,N_68);
and U1608 (N_1608,N_90,N_654);
and U1609 (N_1609,N_207,N_112);
nor U1610 (N_1610,N_859,N_898);
and U1611 (N_1611,N_600,N_853);
or U1612 (N_1612,N_480,N_6);
xor U1613 (N_1613,N_835,N_613);
nor U1614 (N_1614,N_684,N_731);
xor U1615 (N_1615,N_552,N_39);
and U1616 (N_1616,N_677,N_307);
and U1617 (N_1617,N_771,N_395);
nor U1618 (N_1618,N_64,N_21);
xnor U1619 (N_1619,N_36,N_293);
and U1620 (N_1620,N_618,N_388);
nor U1621 (N_1621,N_125,N_880);
nand U1622 (N_1622,N_655,N_158);
nand U1623 (N_1623,N_579,N_769);
xor U1624 (N_1624,N_254,N_498);
xor U1625 (N_1625,N_899,N_593);
xor U1626 (N_1626,N_331,N_377);
or U1627 (N_1627,N_937,N_174);
or U1628 (N_1628,N_180,N_900);
nand U1629 (N_1629,N_641,N_509);
and U1630 (N_1630,N_911,N_947);
nand U1631 (N_1631,N_450,N_158);
xnor U1632 (N_1632,N_932,N_288);
or U1633 (N_1633,N_687,N_823);
xnor U1634 (N_1634,N_460,N_289);
or U1635 (N_1635,N_51,N_514);
xor U1636 (N_1636,N_212,N_740);
or U1637 (N_1637,N_330,N_546);
nand U1638 (N_1638,N_557,N_941);
and U1639 (N_1639,N_946,N_776);
nand U1640 (N_1640,N_528,N_755);
and U1641 (N_1641,N_506,N_636);
xor U1642 (N_1642,N_451,N_59);
nor U1643 (N_1643,N_651,N_599);
xnor U1644 (N_1644,N_904,N_770);
nand U1645 (N_1645,N_553,N_49);
or U1646 (N_1646,N_322,N_58);
or U1647 (N_1647,N_583,N_708);
and U1648 (N_1648,N_451,N_461);
and U1649 (N_1649,N_694,N_385);
nand U1650 (N_1650,N_828,N_468);
nor U1651 (N_1651,N_844,N_679);
or U1652 (N_1652,N_795,N_909);
nand U1653 (N_1653,N_861,N_29);
nor U1654 (N_1654,N_687,N_801);
or U1655 (N_1655,N_897,N_884);
xor U1656 (N_1656,N_677,N_661);
and U1657 (N_1657,N_559,N_943);
nor U1658 (N_1658,N_901,N_826);
nand U1659 (N_1659,N_733,N_27);
nor U1660 (N_1660,N_269,N_623);
nor U1661 (N_1661,N_998,N_258);
nand U1662 (N_1662,N_189,N_477);
or U1663 (N_1663,N_220,N_417);
or U1664 (N_1664,N_43,N_308);
nor U1665 (N_1665,N_429,N_247);
nand U1666 (N_1666,N_358,N_841);
xnor U1667 (N_1667,N_13,N_660);
and U1668 (N_1668,N_576,N_242);
nand U1669 (N_1669,N_969,N_603);
or U1670 (N_1670,N_915,N_419);
nor U1671 (N_1671,N_176,N_238);
nand U1672 (N_1672,N_139,N_36);
xor U1673 (N_1673,N_643,N_112);
and U1674 (N_1674,N_965,N_138);
or U1675 (N_1675,N_229,N_745);
or U1676 (N_1676,N_701,N_325);
and U1677 (N_1677,N_608,N_807);
nor U1678 (N_1678,N_318,N_993);
nor U1679 (N_1679,N_397,N_269);
nand U1680 (N_1680,N_453,N_925);
and U1681 (N_1681,N_671,N_220);
xor U1682 (N_1682,N_650,N_610);
xnor U1683 (N_1683,N_999,N_742);
xnor U1684 (N_1684,N_869,N_271);
or U1685 (N_1685,N_728,N_61);
xnor U1686 (N_1686,N_443,N_474);
or U1687 (N_1687,N_800,N_636);
xnor U1688 (N_1688,N_878,N_509);
or U1689 (N_1689,N_69,N_685);
nor U1690 (N_1690,N_221,N_809);
nor U1691 (N_1691,N_122,N_742);
and U1692 (N_1692,N_305,N_621);
xnor U1693 (N_1693,N_978,N_423);
or U1694 (N_1694,N_45,N_844);
xor U1695 (N_1695,N_477,N_652);
or U1696 (N_1696,N_546,N_15);
xnor U1697 (N_1697,N_143,N_96);
xnor U1698 (N_1698,N_244,N_919);
xor U1699 (N_1699,N_389,N_565);
and U1700 (N_1700,N_992,N_264);
xor U1701 (N_1701,N_523,N_436);
xor U1702 (N_1702,N_435,N_526);
or U1703 (N_1703,N_612,N_581);
nand U1704 (N_1704,N_171,N_960);
xnor U1705 (N_1705,N_724,N_548);
and U1706 (N_1706,N_215,N_432);
nor U1707 (N_1707,N_977,N_3);
nor U1708 (N_1708,N_588,N_885);
nand U1709 (N_1709,N_585,N_249);
or U1710 (N_1710,N_51,N_18);
or U1711 (N_1711,N_23,N_133);
nand U1712 (N_1712,N_668,N_615);
or U1713 (N_1713,N_861,N_962);
nor U1714 (N_1714,N_294,N_297);
xor U1715 (N_1715,N_781,N_742);
nand U1716 (N_1716,N_10,N_642);
nand U1717 (N_1717,N_343,N_14);
and U1718 (N_1718,N_470,N_591);
or U1719 (N_1719,N_720,N_569);
xnor U1720 (N_1720,N_684,N_404);
xnor U1721 (N_1721,N_879,N_450);
and U1722 (N_1722,N_343,N_658);
nand U1723 (N_1723,N_646,N_556);
nand U1724 (N_1724,N_900,N_68);
or U1725 (N_1725,N_436,N_642);
nand U1726 (N_1726,N_422,N_107);
and U1727 (N_1727,N_740,N_564);
nor U1728 (N_1728,N_819,N_345);
and U1729 (N_1729,N_813,N_179);
or U1730 (N_1730,N_65,N_388);
or U1731 (N_1731,N_238,N_923);
or U1732 (N_1732,N_18,N_888);
nand U1733 (N_1733,N_89,N_565);
or U1734 (N_1734,N_381,N_489);
or U1735 (N_1735,N_801,N_372);
xnor U1736 (N_1736,N_482,N_397);
and U1737 (N_1737,N_252,N_620);
xor U1738 (N_1738,N_425,N_12);
or U1739 (N_1739,N_433,N_372);
xor U1740 (N_1740,N_253,N_617);
nand U1741 (N_1741,N_772,N_379);
or U1742 (N_1742,N_93,N_450);
nand U1743 (N_1743,N_831,N_293);
or U1744 (N_1744,N_354,N_446);
and U1745 (N_1745,N_296,N_744);
xnor U1746 (N_1746,N_954,N_976);
and U1747 (N_1747,N_730,N_687);
xnor U1748 (N_1748,N_236,N_824);
nor U1749 (N_1749,N_565,N_227);
xor U1750 (N_1750,N_483,N_230);
and U1751 (N_1751,N_894,N_175);
and U1752 (N_1752,N_102,N_887);
or U1753 (N_1753,N_69,N_530);
nor U1754 (N_1754,N_300,N_806);
and U1755 (N_1755,N_90,N_412);
or U1756 (N_1756,N_318,N_798);
xnor U1757 (N_1757,N_55,N_171);
or U1758 (N_1758,N_117,N_36);
nand U1759 (N_1759,N_794,N_891);
or U1760 (N_1760,N_700,N_7);
and U1761 (N_1761,N_880,N_886);
nor U1762 (N_1762,N_255,N_706);
xnor U1763 (N_1763,N_814,N_167);
and U1764 (N_1764,N_579,N_154);
nand U1765 (N_1765,N_414,N_124);
or U1766 (N_1766,N_594,N_451);
or U1767 (N_1767,N_839,N_915);
nand U1768 (N_1768,N_106,N_693);
or U1769 (N_1769,N_250,N_65);
nand U1770 (N_1770,N_892,N_480);
or U1771 (N_1771,N_996,N_307);
nor U1772 (N_1772,N_589,N_775);
or U1773 (N_1773,N_839,N_335);
or U1774 (N_1774,N_957,N_653);
nand U1775 (N_1775,N_974,N_407);
and U1776 (N_1776,N_53,N_854);
and U1777 (N_1777,N_140,N_725);
nor U1778 (N_1778,N_665,N_955);
xnor U1779 (N_1779,N_639,N_166);
nand U1780 (N_1780,N_70,N_984);
xor U1781 (N_1781,N_651,N_589);
and U1782 (N_1782,N_775,N_781);
xnor U1783 (N_1783,N_919,N_323);
xor U1784 (N_1784,N_193,N_712);
and U1785 (N_1785,N_919,N_768);
xnor U1786 (N_1786,N_29,N_357);
or U1787 (N_1787,N_894,N_110);
and U1788 (N_1788,N_499,N_483);
and U1789 (N_1789,N_251,N_666);
xnor U1790 (N_1790,N_118,N_989);
or U1791 (N_1791,N_330,N_790);
and U1792 (N_1792,N_165,N_76);
or U1793 (N_1793,N_536,N_266);
xnor U1794 (N_1794,N_49,N_702);
and U1795 (N_1795,N_783,N_20);
nor U1796 (N_1796,N_341,N_382);
nand U1797 (N_1797,N_550,N_166);
xor U1798 (N_1798,N_601,N_274);
nand U1799 (N_1799,N_628,N_489);
nor U1800 (N_1800,N_955,N_932);
and U1801 (N_1801,N_619,N_453);
nand U1802 (N_1802,N_583,N_774);
nand U1803 (N_1803,N_740,N_813);
nand U1804 (N_1804,N_329,N_215);
nand U1805 (N_1805,N_250,N_667);
and U1806 (N_1806,N_260,N_592);
nor U1807 (N_1807,N_676,N_994);
xor U1808 (N_1808,N_856,N_301);
xor U1809 (N_1809,N_655,N_525);
nor U1810 (N_1810,N_704,N_964);
or U1811 (N_1811,N_666,N_77);
nor U1812 (N_1812,N_972,N_162);
or U1813 (N_1813,N_493,N_671);
xnor U1814 (N_1814,N_824,N_410);
and U1815 (N_1815,N_400,N_968);
nor U1816 (N_1816,N_597,N_519);
xnor U1817 (N_1817,N_764,N_199);
nand U1818 (N_1818,N_165,N_187);
or U1819 (N_1819,N_394,N_314);
and U1820 (N_1820,N_649,N_188);
nor U1821 (N_1821,N_231,N_390);
nand U1822 (N_1822,N_11,N_791);
or U1823 (N_1823,N_705,N_886);
or U1824 (N_1824,N_581,N_121);
and U1825 (N_1825,N_466,N_374);
xnor U1826 (N_1826,N_177,N_283);
nor U1827 (N_1827,N_474,N_19);
nand U1828 (N_1828,N_703,N_872);
and U1829 (N_1829,N_243,N_771);
or U1830 (N_1830,N_374,N_791);
and U1831 (N_1831,N_84,N_292);
xor U1832 (N_1832,N_271,N_127);
or U1833 (N_1833,N_545,N_784);
or U1834 (N_1834,N_940,N_798);
and U1835 (N_1835,N_469,N_572);
xnor U1836 (N_1836,N_956,N_327);
nand U1837 (N_1837,N_963,N_403);
xnor U1838 (N_1838,N_717,N_154);
nor U1839 (N_1839,N_382,N_653);
xor U1840 (N_1840,N_151,N_697);
xor U1841 (N_1841,N_458,N_84);
xor U1842 (N_1842,N_83,N_581);
nand U1843 (N_1843,N_965,N_733);
nor U1844 (N_1844,N_221,N_693);
nand U1845 (N_1845,N_152,N_68);
or U1846 (N_1846,N_126,N_487);
xor U1847 (N_1847,N_214,N_564);
xor U1848 (N_1848,N_204,N_473);
nand U1849 (N_1849,N_859,N_644);
and U1850 (N_1850,N_824,N_775);
nor U1851 (N_1851,N_76,N_589);
or U1852 (N_1852,N_66,N_989);
xor U1853 (N_1853,N_5,N_483);
nand U1854 (N_1854,N_578,N_311);
nand U1855 (N_1855,N_281,N_787);
nor U1856 (N_1856,N_353,N_486);
nor U1857 (N_1857,N_529,N_650);
nand U1858 (N_1858,N_97,N_711);
nor U1859 (N_1859,N_755,N_845);
xnor U1860 (N_1860,N_339,N_359);
and U1861 (N_1861,N_630,N_123);
nand U1862 (N_1862,N_145,N_728);
and U1863 (N_1863,N_156,N_733);
nand U1864 (N_1864,N_226,N_505);
and U1865 (N_1865,N_677,N_477);
nand U1866 (N_1866,N_70,N_418);
nand U1867 (N_1867,N_835,N_596);
or U1868 (N_1868,N_448,N_823);
nand U1869 (N_1869,N_943,N_981);
or U1870 (N_1870,N_969,N_720);
nor U1871 (N_1871,N_996,N_400);
xor U1872 (N_1872,N_669,N_560);
nor U1873 (N_1873,N_818,N_978);
nor U1874 (N_1874,N_78,N_686);
nand U1875 (N_1875,N_790,N_406);
xnor U1876 (N_1876,N_519,N_681);
nand U1877 (N_1877,N_651,N_883);
or U1878 (N_1878,N_326,N_452);
nand U1879 (N_1879,N_389,N_96);
nand U1880 (N_1880,N_540,N_606);
nor U1881 (N_1881,N_459,N_314);
nand U1882 (N_1882,N_302,N_747);
xor U1883 (N_1883,N_590,N_153);
or U1884 (N_1884,N_379,N_151);
and U1885 (N_1885,N_356,N_3);
xor U1886 (N_1886,N_610,N_340);
or U1887 (N_1887,N_841,N_746);
and U1888 (N_1888,N_66,N_543);
or U1889 (N_1889,N_583,N_684);
xnor U1890 (N_1890,N_342,N_906);
xnor U1891 (N_1891,N_326,N_413);
nor U1892 (N_1892,N_47,N_525);
nor U1893 (N_1893,N_562,N_156);
nand U1894 (N_1894,N_236,N_477);
and U1895 (N_1895,N_133,N_624);
nand U1896 (N_1896,N_887,N_829);
nor U1897 (N_1897,N_408,N_804);
nor U1898 (N_1898,N_418,N_305);
xor U1899 (N_1899,N_196,N_832);
nand U1900 (N_1900,N_215,N_556);
and U1901 (N_1901,N_363,N_664);
nor U1902 (N_1902,N_211,N_246);
nor U1903 (N_1903,N_875,N_328);
or U1904 (N_1904,N_111,N_678);
or U1905 (N_1905,N_140,N_197);
nand U1906 (N_1906,N_628,N_263);
nand U1907 (N_1907,N_445,N_610);
or U1908 (N_1908,N_193,N_217);
or U1909 (N_1909,N_705,N_17);
and U1910 (N_1910,N_220,N_426);
or U1911 (N_1911,N_750,N_645);
xnor U1912 (N_1912,N_738,N_196);
and U1913 (N_1913,N_259,N_557);
or U1914 (N_1914,N_877,N_862);
xnor U1915 (N_1915,N_709,N_559);
nor U1916 (N_1916,N_671,N_371);
and U1917 (N_1917,N_343,N_55);
xor U1918 (N_1918,N_975,N_484);
nand U1919 (N_1919,N_12,N_926);
and U1920 (N_1920,N_182,N_626);
xnor U1921 (N_1921,N_750,N_377);
and U1922 (N_1922,N_835,N_689);
or U1923 (N_1923,N_209,N_506);
nand U1924 (N_1924,N_855,N_45);
nand U1925 (N_1925,N_415,N_85);
nor U1926 (N_1926,N_958,N_76);
nor U1927 (N_1927,N_534,N_423);
nor U1928 (N_1928,N_614,N_752);
and U1929 (N_1929,N_521,N_545);
nor U1930 (N_1930,N_807,N_412);
xor U1931 (N_1931,N_785,N_277);
or U1932 (N_1932,N_927,N_971);
or U1933 (N_1933,N_736,N_634);
and U1934 (N_1934,N_795,N_858);
or U1935 (N_1935,N_863,N_227);
nand U1936 (N_1936,N_830,N_728);
or U1937 (N_1937,N_392,N_776);
nand U1938 (N_1938,N_645,N_145);
nor U1939 (N_1939,N_702,N_312);
and U1940 (N_1940,N_875,N_219);
nand U1941 (N_1941,N_93,N_748);
nor U1942 (N_1942,N_375,N_916);
and U1943 (N_1943,N_391,N_868);
or U1944 (N_1944,N_359,N_633);
xnor U1945 (N_1945,N_48,N_263);
nor U1946 (N_1946,N_473,N_756);
and U1947 (N_1947,N_187,N_792);
or U1948 (N_1948,N_528,N_154);
or U1949 (N_1949,N_348,N_767);
nor U1950 (N_1950,N_58,N_300);
xnor U1951 (N_1951,N_206,N_501);
or U1952 (N_1952,N_222,N_138);
nor U1953 (N_1953,N_466,N_15);
or U1954 (N_1954,N_641,N_955);
and U1955 (N_1955,N_718,N_544);
nor U1956 (N_1956,N_610,N_782);
nor U1957 (N_1957,N_261,N_3);
and U1958 (N_1958,N_51,N_721);
xor U1959 (N_1959,N_581,N_240);
and U1960 (N_1960,N_284,N_409);
or U1961 (N_1961,N_51,N_814);
or U1962 (N_1962,N_516,N_162);
or U1963 (N_1963,N_278,N_892);
xor U1964 (N_1964,N_555,N_662);
xor U1965 (N_1965,N_139,N_445);
or U1966 (N_1966,N_74,N_457);
nor U1967 (N_1967,N_673,N_888);
xor U1968 (N_1968,N_345,N_6);
xnor U1969 (N_1969,N_629,N_67);
nand U1970 (N_1970,N_950,N_56);
nor U1971 (N_1971,N_359,N_644);
and U1972 (N_1972,N_925,N_354);
xnor U1973 (N_1973,N_380,N_833);
nand U1974 (N_1974,N_739,N_293);
and U1975 (N_1975,N_868,N_854);
xor U1976 (N_1976,N_651,N_913);
or U1977 (N_1977,N_48,N_922);
nor U1978 (N_1978,N_766,N_867);
nor U1979 (N_1979,N_792,N_889);
and U1980 (N_1980,N_727,N_621);
and U1981 (N_1981,N_846,N_734);
nor U1982 (N_1982,N_928,N_839);
or U1983 (N_1983,N_841,N_588);
or U1984 (N_1984,N_855,N_939);
nor U1985 (N_1985,N_303,N_546);
or U1986 (N_1986,N_707,N_31);
nand U1987 (N_1987,N_816,N_783);
xnor U1988 (N_1988,N_668,N_649);
nand U1989 (N_1989,N_517,N_798);
or U1990 (N_1990,N_577,N_33);
nand U1991 (N_1991,N_532,N_815);
nand U1992 (N_1992,N_200,N_677);
nor U1993 (N_1993,N_735,N_411);
xor U1994 (N_1994,N_202,N_20);
or U1995 (N_1995,N_213,N_364);
or U1996 (N_1996,N_557,N_339);
nand U1997 (N_1997,N_395,N_402);
nand U1998 (N_1998,N_945,N_159);
nor U1999 (N_1999,N_808,N_127);
nor U2000 (N_2000,N_1364,N_1376);
nor U2001 (N_2001,N_1015,N_1433);
nand U2002 (N_2002,N_1793,N_1182);
nand U2003 (N_2003,N_1621,N_1692);
or U2004 (N_2004,N_1505,N_1372);
or U2005 (N_2005,N_1881,N_1730);
xor U2006 (N_2006,N_1788,N_1844);
and U2007 (N_2007,N_1579,N_1446);
nor U2008 (N_2008,N_1922,N_1590);
and U2009 (N_2009,N_1003,N_1865);
xor U2010 (N_2010,N_1029,N_1897);
nor U2011 (N_2011,N_1195,N_1175);
nor U2012 (N_2012,N_1550,N_1190);
nor U2013 (N_2013,N_1752,N_1496);
or U2014 (N_2014,N_1271,N_1463);
xor U2015 (N_2015,N_1298,N_1597);
nand U2016 (N_2016,N_1246,N_1239);
nand U2017 (N_2017,N_1030,N_1201);
nor U2018 (N_2018,N_1088,N_1458);
nand U2019 (N_2019,N_1371,N_1420);
and U2020 (N_2020,N_1279,N_1722);
or U2021 (N_2021,N_1207,N_1936);
nand U2022 (N_2022,N_1316,N_1028);
and U2023 (N_2023,N_1381,N_1598);
nor U2024 (N_2024,N_1322,N_1642);
xnor U2025 (N_2025,N_1146,N_1720);
and U2026 (N_2026,N_1506,N_1724);
nor U2027 (N_2027,N_1554,N_1929);
and U2028 (N_2028,N_1901,N_1985);
or U2029 (N_2029,N_1685,N_1112);
nor U2030 (N_2030,N_1711,N_1065);
or U2031 (N_2031,N_1221,N_1935);
and U2032 (N_2032,N_1084,N_1682);
or U2033 (N_2033,N_1532,N_1052);
nand U2034 (N_2034,N_1803,N_1244);
nor U2035 (N_2035,N_1307,N_1157);
nand U2036 (N_2036,N_1672,N_1773);
xor U2037 (N_2037,N_1904,N_1600);
nand U2038 (N_2038,N_1938,N_1261);
or U2039 (N_2039,N_1409,N_1868);
nand U2040 (N_2040,N_1323,N_1305);
xnor U2041 (N_2041,N_1884,N_1419);
nor U2042 (N_2042,N_1217,N_1510);
and U2043 (N_2043,N_1796,N_1679);
xor U2044 (N_2044,N_1194,N_1330);
xor U2045 (N_2045,N_1304,N_1238);
xor U2046 (N_2046,N_1442,N_1066);
xnor U2047 (N_2047,N_1222,N_1866);
or U2048 (N_2048,N_1961,N_1278);
nor U2049 (N_2049,N_1768,N_1824);
nor U2050 (N_2050,N_1129,N_1503);
nand U2051 (N_2051,N_1426,N_1893);
nor U2052 (N_2052,N_1523,N_1368);
or U2053 (N_2053,N_1185,N_1334);
or U2054 (N_2054,N_1257,N_1125);
nor U2055 (N_2055,N_1815,N_1921);
and U2056 (N_2056,N_1563,N_1749);
xor U2057 (N_2057,N_1662,N_1604);
and U2058 (N_2058,N_1348,N_1913);
and U2059 (N_2059,N_1220,N_1297);
or U2060 (N_2060,N_1111,N_1591);
and U2061 (N_2061,N_1704,N_1601);
nand U2062 (N_2062,N_1219,N_1694);
nand U2063 (N_2063,N_1500,N_1115);
nor U2064 (N_2064,N_1101,N_1479);
or U2065 (N_2065,N_1417,N_1610);
or U2066 (N_2066,N_1161,N_1451);
nand U2067 (N_2067,N_1860,N_1189);
and U2068 (N_2068,N_1080,N_1646);
and U2069 (N_2069,N_1756,N_1117);
nand U2070 (N_2070,N_1141,N_1949);
xnor U2071 (N_2071,N_1365,N_1840);
xnor U2072 (N_2072,N_1018,N_1128);
nor U2073 (N_2073,N_1567,N_1605);
xor U2074 (N_2074,N_1122,N_1719);
nand U2075 (N_2075,N_1648,N_1394);
xor U2076 (N_2076,N_1032,N_1039);
and U2077 (N_2077,N_1887,N_1953);
nand U2078 (N_2078,N_1202,N_1483);
xnor U2079 (N_2079,N_1143,N_1634);
and U2080 (N_2080,N_1068,N_1245);
and U2081 (N_2081,N_1250,N_1658);
and U2082 (N_2082,N_1502,N_1940);
xnor U2083 (N_2083,N_1732,N_1671);
xnor U2084 (N_2084,N_1772,N_1176);
nand U2085 (N_2085,N_1465,N_1745);
nand U2086 (N_2086,N_1274,N_1275);
xnor U2087 (N_2087,N_1665,N_1613);
and U2088 (N_2088,N_1331,N_1473);
nand U2089 (N_2089,N_1937,N_1355);
xnor U2090 (N_2090,N_1551,N_1235);
and U2091 (N_2091,N_1888,N_1301);
nand U2092 (N_2092,N_1814,N_1431);
and U2093 (N_2093,N_1262,N_1294);
nand U2094 (N_2094,N_1624,N_1452);
nor U2095 (N_2095,N_1973,N_1863);
or U2096 (N_2096,N_1078,N_1050);
and U2097 (N_2097,N_1499,N_1413);
xnor U2098 (N_2098,N_1676,N_1954);
xnor U2099 (N_2099,N_1459,N_1988);
and U2100 (N_2100,N_1821,N_1236);
nand U2101 (N_2101,N_1638,N_1025);
or U2102 (N_2102,N_1046,N_1683);
or U2103 (N_2103,N_1491,N_1461);
nor U2104 (N_2104,N_1325,N_1769);
and U2105 (N_2105,N_1209,N_1789);
nand U2106 (N_2106,N_1708,N_1492);
xnor U2107 (N_2107,N_1012,N_1467);
nor U2108 (N_2108,N_1177,N_1609);
nand U2109 (N_2109,N_1964,N_1771);
xnor U2110 (N_2110,N_1472,N_1873);
and U2111 (N_2111,N_1540,N_1140);
nor U2112 (N_2112,N_1932,N_1854);
xor U2113 (N_2113,N_1688,N_1059);
nand U2114 (N_2114,N_1623,N_1317);
and U2115 (N_2115,N_1537,N_1418);
nor U2116 (N_2116,N_1268,N_1170);
xor U2117 (N_2117,N_1852,N_1497);
nand U2118 (N_2118,N_1121,N_1941);
nand U2119 (N_2119,N_1074,N_1763);
nand U2120 (N_2120,N_1741,N_1819);
or U2121 (N_2121,N_1572,N_1526);
and U2122 (N_2122,N_1747,N_1515);
nor U2123 (N_2123,N_1790,N_1971);
and U2124 (N_2124,N_1280,N_1197);
and U2125 (N_2125,N_1020,N_1920);
and U2126 (N_2126,N_1583,N_1155);
xor U2127 (N_2127,N_1192,N_1234);
and U2128 (N_2128,N_1669,N_1160);
xor U2129 (N_2129,N_1549,N_1438);
nand U2130 (N_2130,N_1454,N_1653);
or U2131 (N_2131,N_1931,N_1726);
xnor U2132 (N_2132,N_1594,N_1535);
nand U2133 (N_2133,N_1064,N_1849);
xor U2134 (N_2134,N_1809,N_1460);
xor U2135 (N_2135,N_1343,N_1149);
xor U2136 (N_2136,N_1797,N_1320);
and U2137 (N_2137,N_1909,N_1488);
nor U2138 (N_2138,N_1341,N_1043);
nand U2139 (N_2139,N_1620,N_1309);
or U2140 (N_2140,N_1543,N_1282);
nand U2141 (N_2141,N_1373,N_1783);
or U2142 (N_2142,N_1260,N_1955);
xor U2143 (N_2143,N_1359,N_1782);
nand U2144 (N_2144,N_1384,N_1163);
xor U2145 (N_2145,N_1017,N_1392);
nor U2146 (N_2146,N_1389,N_1753);
and U2147 (N_2147,N_1332,N_1478);
nand U2148 (N_2148,N_1013,N_1135);
and U2149 (N_2149,N_1344,N_1486);
nand U2150 (N_2150,N_1009,N_1794);
nor U2151 (N_2151,N_1541,N_1210);
nand U2152 (N_2152,N_1205,N_1952);
nor U2153 (N_2153,N_1437,N_1237);
nand U2154 (N_2154,N_1660,N_1379);
xnor U2155 (N_2155,N_1656,N_1837);
nand U2156 (N_2156,N_1686,N_1524);
xor U2157 (N_2157,N_1213,N_1361);
or U2158 (N_2158,N_1233,N_1657);
and U2159 (N_2159,N_1630,N_1617);
nor U2160 (N_2160,N_1681,N_1761);
or U2161 (N_2161,N_1200,N_1870);
xor U2162 (N_2162,N_1619,N_1536);
nand U2163 (N_2163,N_1928,N_1443);
and U2164 (N_2164,N_1996,N_1659);
xnor U2165 (N_2165,N_1021,N_1575);
xnor U2166 (N_2166,N_1900,N_1310);
xnor U2167 (N_2167,N_1602,N_1340);
nand U2168 (N_2168,N_1303,N_1053);
xor U2169 (N_2169,N_1559,N_1725);
xnor U2170 (N_2170,N_1777,N_1586);
or U2171 (N_2171,N_1640,N_1440);
or U2172 (N_2172,N_1022,N_1926);
nand U2173 (N_2173,N_1302,N_1089);
nand U2174 (N_2174,N_1919,N_1315);
and U2175 (N_2175,N_1166,N_1739);
or U2176 (N_2176,N_1407,N_1010);
nor U2177 (N_2177,N_1891,N_1716);
nor U2178 (N_2178,N_1116,N_1487);
nand U2179 (N_2179,N_1999,N_1430);
or U2180 (N_2180,N_1918,N_1987);
nor U2181 (N_2181,N_1830,N_1435);
xnor U2182 (N_2182,N_1896,N_1707);
and U2183 (N_2183,N_1829,N_1277);
and U2184 (N_2184,N_1061,N_1810);
nor U2185 (N_2185,N_1637,N_1589);
xor U2186 (N_2186,N_1108,N_1758);
or U2187 (N_2187,N_1951,N_1718);
nor U2188 (N_2188,N_1740,N_1156);
and U2189 (N_2189,N_1049,N_1023);
and U2190 (N_2190,N_1085,N_1026);
xor U2191 (N_2191,N_1997,N_1991);
and U2192 (N_2192,N_1073,N_1511);
nor U2193 (N_2193,N_1054,N_1568);
or U2194 (N_2194,N_1075,N_1818);
and U2195 (N_2195,N_1946,N_1784);
nand U2196 (N_2196,N_1110,N_1983);
nor U2197 (N_2197,N_1979,N_1570);
xor U2198 (N_2198,N_1415,N_1915);
or U2199 (N_2199,N_1705,N_1391);
xnor U2200 (N_2200,N_1071,N_1173);
or U2201 (N_2201,N_1070,N_1436);
xor U2202 (N_2202,N_1000,N_1644);
nand U2203 (N_2203,N_1147,N_1456);
xnor U2204 (N_2204,N_1930,N_1346);
nor U2205 (N_2205,N_1060,N_1569);
nor U2206 (N_2206,N_1853,N_1048);
and U2207 (N_2207,N_1848,N_1347);
nor U2208 (N_2208,N_1103,N_1948);
xor U2209 (N_2209,N_1943,N_1318);
nand U2210 (N_2210,N_1399,N_1336);
xnor U2211 (N_2211,N_1910,N_1240);
xor U2212 (N_2212,N_1269,N_1735);
nand U2213 (N_2213,N_1998,N_1780);
nor U2214 (N_2214,N_1545,N_1882);
and U2215 (N_2215,N_1556,N_1828);
and U2216 (N_2216,N_1158,N_1475);
and U2217 (N_2217,N_1847,N_1776);
nor U2218 (N_2218,N_1151,N_1357);
or U2219 (N_2219,N_1203,N_1811);
nand U2220 (N_2220,N_1327,N_1193);
nor U2221 (N_2221,N_1611,N_1041);
nand U2222 (N_2222,N_1291,N_1011);
nand U2223 (N_2223,N_1034,N_1582);
and U2224 (N_2224,N_1516,N_1077);
and U2225 (N_2225,N_1970,N_1558);
xnor U2226 (N_2226,N_1104,N_1944);
xor U2227 (N_2227,N_1875,N_1764);
xnor U2228 (N_2228,N_1124,N_1801);
and U2229 (N_2229,N_1286,N_1527);
xnor U2230 (N_2230,N_1138,N_1664);
nor U2231 (N_2231,N_1639,N_1733);
nor U2232 (N_2232,N_1967,N_1565);
nand U2233 (N_2233,N_1227,N_1439);
xor U2234 (N_2234,N_1521,N_1595);
xnor U2235 (N_2235,N_1636,N_1787);
or U2236 (N_2236,N_1014,N_1514);
or U2237 (N_2237,N_1395,N_1670);
nor U2238 (N_2238,N_1468,N_1889);
xor U2239 (N_2239,N_1522,N_1218);
and U2240 (N_2240,N_1062,N_1287);
and U2241 (N_2241,N_1493,N_1040);
and U2242 (N_2242,N_1518,N_1765);
nor U2243 (N_2243,N_1480,N_1106);
nor U2244 (N_2244,N_1421,N_1629);
nor U2245 (N_2245,N_1786,N_1383);
nand U2246 (N_2246,N_1120,N_1877);
nor U2247 (N_2247,N_1416,N_1299);
xor U2248 (N_2248,N_1546,N_1878);
xnor U2249 (N_2249,N_1845,N_1817);
xor U2250 (N_2250,N_1584,N_1661);
and U2251 (N_2251,N_1172,N_1666);
nand U2252 (N_2252,N_1641,N_1804);
nor U2253 (N_2253,N_1547,N_1827);
nand U2254 (N_2254,N_1615,N_1180);
and U2255 (N_2255,N_1469,N_1693);
xor U2256 (N_2256,N_1016,N_1097);
xor U2257 (N_2257,N_1126,N_1035);
nor U2258 (N_2258,N_1295,N_1553);
nor U2259 (N_2259,N_1574,N_1649);
xor U2260 (N_2260,N_1750,N_1127);
or U2261 (N_2261,N_1628,N_1880);
or U2262 (N_2262,N_1945,N_1476);
nand U2263 (N_2263,N_1531,N_1335);
or U2264 (N_2264,N_1485,N_1678);
or U2265 (N_2265,N_1706,N_1037);
nor U2266 (N_2266,N_1489,N_1164);
xor U2267 (N_2267,N_1313,N_1230);
xnor U2268 (N_2268,N_1215,N_1775);
xor U2269 (N_2269,N_1975,N_1051);
or U2270 (N_2270,N_1822,N_1337);
nor U2271 (N_2271,N_1593,N_1248);
xnor U2272 (N_2272,N_1603,N_1162);
and U2273 (N_2273,N_1872,N_1288);
nor U2274 (N_2274,N_1224,N_1731);
or U2275 (N_2275,N_1957,N_1885);
or U2276 (N_2276,N_1131,N_1984);
xnor U2277 (N_2277,N_1153,N_1963);
nand U2278 (N_2278,N_1429,N_1767);
nand U2279 (N_2279,N_1960,N_1802);
nor U2280 (N_2280,N_1701,N_1422);
xor U2281 (N_2281,N_1779,N_1191);
or U2282 (N_2282,N_1861,N_1695);
nor U2283 (N_2283,N_1807,N_1328);
and U2284 (N_2284,N_1912,N_1862);
nand U2285 (N_2285,N_1241,N_1256);
nand U2286 (N_2286,N_1843,N_1186);
and U2287 (N_2287,N_1424,N_1007);
xnor U2288 (N_2288,N_1857,N_1895);
xnor U2289 (N_2289,N_1044,N_1375);
nor U2290 (N_2290,N_1805,N_1006);
xor U2291 (N_2291,N_1552,N_1380);
and U2292 (N_2292,N_1905,N_1178);
and U2293 (N_2293,N_1923,N_1374);
nor U2294 (N_2294,N_1482,N_1585);
or U2295 (N_2295,N_1367,N_1942);
nor U2296 (N_2296,N_1181,N_1076);
xor U2297 (N_2297,N_1211,N_1806);
xnor U2298 (N_2298,N_1036,N_1414);
or U2299 (N_2299,N_1114,N_1632);
xor U2300 (N_2300,N_1995,N_1455);
xnor U2301 (N_2301,N_1512,N_1292);
nand U2302 (N_2302,N_1377,N_1539);
or U2303 (N_2303,N_1816,N_1981);
nand U2304 (N_2304,N_1136,N_1994);
nor U2305 (N_2305,N_1069,N_1762);
nand U2306 (N_2306,N_1850,N_1154);
nand U2307 (N_2307,N_1742,N_1027);
nor U2308 (N_2308,N_1466,N_1226);
xnor U2309 (N_2309,N_1091,N_1618);
nor U2310 (N_2310,N_1864,N_1319);
and U2311 (N_2311,N_1107,N_1736);
or U2312 (N_2312,N_1339,N_1096);
nor U2313 (N_2313,N_1974,N_1557);
xnor U2314 (N_2314,N_1703,N_1883);
nand U2315 (N_2315,N_1564,N_1766);
nor U2316 (N_2316,N_1823,N_1754);
and U2317 (N_2317,N_1792,N_1675);
and U2318 (N_2318,N_1699,N_1024);
nand U2319 (N_2319,N_1696,N_1321);
nand U2320 (N_2320,N_1168,N_1498);
nand U2321 (N_2321,N_1836,N_1687);
xnor U2322 (N_2322,N_1428,N_1859);
or U2323 (N_2323,N_1738,N_1312);
and U2324 (N_2324,N_1100,N_1353);
or U2325 (N_2325,N_1174,N_1925);
or U2326 (N_2326,N_1133,N_1102);
nor U2327 (N_2327,N_1571,N_1179);
nor U2328 (N_2328,N_1019,N_1993);
nand U2329 (N_2329,N_1145,N_1093);
xnor U2330 (N_2330,N_1588,N_1229);
and U2331 (N_2331,N_1423,N_1966);
or U2332 (N_2332,N_1517,N_1989);
xnor U2333 (N_2333,N_1907,N_1072);
nor U2334 (N_2334,N_1232,N_1614);
or U2335 (N_2335,N_1728,N_1587);
nand U2336 (N_2336,N_1652,N_1338);
xnor U2337 (N_2337,N_1791,N_1978);
nand U2338 (N_2338,N_1729,N_1757);
nor U2339 (N_2339,N_1002,N_1902);
and U2340 (N_2340,N_1645,N_1962);
nand U2341 (N_2341,N_1228,N_1898);
nor U2342 (N_2342,N_1311,N_1643);
nand U2343 (N_2343,N_1055,N_1401);
nand U2344 (N_2344,N_1734,N_1408);
xor U2345 (N_2345,N_1231,N_1406);
and U2346 (N_2346,N_1410,N_1281);
xnor U2347 (N_2347,N_1434,N_1087);
and U2348 (N_2348,N_1171,N_1698);
xnor U2349 (N_2349,N_1358,N_1047);
nor U2350 (N_2350,N_1977,N_1223);
xor U2351 (N_2351,N_1284,N_1684);
xor U2352 (N_2352,N_1714,N_1090);
nand U2353 (N_2353,N_1300,N_1225);
and U2354 (N_2354,N_1362,N_1566);
nand U2355 (N_2355,N_1042,N_1654);
or U2356 (N_2356,N_1033,N_1109);
nand U2357 (N_2357,N_1599,N_1397);
nor U2358 (N_2358,N_1204,N_1134);
or U2359 (N_2359,N_1691,N_1132);
nand U2360 (N_2360,N_1118,N_1917);
nor U2361 (N_2361,N_1249,N_1958);
and U2362 (N_2362,N_1095,N_1382);
or U2363 (N_2363,N_1031,N_1378);
and U2364 (N_2364,N_1519,N_1462);
and U2365 (N_2365,N_1445,N_1533);
and U2366 (N_2366,N_1390,N_1148);
nand U2367 (N_2367,N_1785,N_1137);
and U2368 (N_2368,N_1504,N_1908);
and U2369 (N_2369,N_1717,N_1534);
nand U2370 (N_2370,N_1258,N_1270);
and U2371 (N_2371,N_1755,N_1259);
xor U2372 (N_2372,N_1965,N_1581);
and U2373 (N_2373,N_1525,N_1214);
nand U2374 (N_2374,N_1251,N_1825);
or U2375 (N_2375,N_1079,N_1247);
nor U2376 (N_2376,N_1289,N_1555);
nor U2377 (N_2377,N_1871,N_1663);
and U2378 (N_2378,N_1266,N_1188);
and U2379 (N_2379,N_1737,N_1254);
nand U2380 (N_2380,N_1577,N_1832);
xnor U2381 (N_2381,N_1142,N_1838);
nand U2382 (N_2382,N_1253,N_1184);
xnor U2383 (N_2383,N_1899,N_1008);
and U2384 (N_2384,N_1094,N_1911);
xor U2385 (N_2385,N_1464,N_1529);
nor U2386 (N_2386,N_1723,N_1252);
xor U2387 (N_2387,N_1976,N_1744);
or U2388 (N_2388,N_1083,N_1573);
nor U2389 (N_2389,N_1130,N_1612);
nor U2390 (N_2390,N_1842,N_1086);
or U2391 (N_2391,N_1934,N_1352);
nand U2392 (N_2392,N_1308,N_1360);
nand U2393 (N_2393,N_1990,N_1808);
nor U2394 (N_2394,N_1199,N_1982);
nand U2395 (N_2395,N_1856,N_1324);
and U2396 (N_2396,N_1712,N_1082);
xnor U2397 (N_2397,N_1329,N_1306);
nor U2398 (N_2398,N_1349,N_1947);
xnor U2399 (N_2399,N_1702,N_1187);
nor U2400 (N_2400,N_1448,N_1333);
and U2401 (N_2401,N_1677,N_1385);
nor U2402 (N_2402,N_1820,N_1798);
or U2403 (N_2403,N_1484,N_1916);
and U2404 (N_2404,N_1625,N_1152);
xor U2405 (N_2405,N_1879,N_1432);
or U2406 (N_2406,N_1063,N_1759);
nand U2407 (N_2407,N_1580,N_1933);
nand U2408 (N_2408,N_1606,N_1139);
and U2409 (N_2409,N_1099,N_1903);
nor U2410 (N_2410,N_1405,N_1273);
xnor U2411 (N_2411,N_1813,N_1631);
nand U2412 (N_2412,N_1490,N_1457);
nand U2413 (N_2413,N_1835,N_1781);
or U2414 (N_2414,N_1393,N_1208);
xor U2415 (N_2415,N_1098,N_1616);
and U2416 (N_2416,N_1400,N_1800);
nand U2417 (N_2417,N_1528,N_1370);
nor U2418 (N_2418,N_1548,N_1746);
xor U2419 (N_2419,N_1561,N_1650);
or U2420 (N_2420,N_1959,N_1892);
or U2421 (N_2421,N_1402,N_1004);
xnor U2422 (N_2422,N_1647,N_1544);
or U2423 (N_2423,N_1412,N_1255);
xor U2424 (N_2424,N_1542,N_1427);
or U2425 (N_2425,N_1351,N_1474);
or U2426 (N_2426,N_1283,N_1560);
nand U2427 (N_2427,N_1263,N_1388);
and U2428 (N_2428,N_1495,N_1450);
nand U2429 (N_2429,N_1715,N_1092);
nand U2430 (N_2430,N_1354,N_1369);
xor U2431 (N_2431,N_1627,N_1869);
nor U2432 (N_2432,N_1285,N_1150);
xnor U2433 (N_2433,N_1453,N_1607);
or U2434 (N_2434,N_1196,N_1774);
xor U2435 (N_2435,N_1481,N_1894);
nand U2436 (N_2436,N_1342,N_1626);
nor U2437 (N_2437,N_1356,N_1169);
or U2438 (N_2438,N_1363,N_1045);
and U2439 (N_2439,N_1513,N_1538);
or U2440 (N_2440,N_1350,N_1673);
nand U2441 (N_2441,N_1743,N_1846);
nand U2442 (N_2442,N_1326,N_1710);
or U2443 (N_2443,N_1890,N_1058);
or U2444 (N_2444,N_1855,N_1345);
xor U2445 (N_2445,N_1276,N_1449);
or U2446 (N_2446,N_1144,N_1296);
nor U2447 (N_2447,N_1206,N_1709);
nor U2448 (N_2448,N_1471,N_1576);
xnor U2449 (N_2449,N_1697,N_1387);
and U2450 (N_2450,N_1167,N_1212);
nor U2451 (N_2451,N_1633,N_1690);
and U2452 (N_2452,N_1608,N_1198);
nand U2453 (N_2453,N_1596,N_1470);
xnor U2454 (N_2454,N_1293,N_1839);
nor U2455 (N_2455,N_1727,N_1924);
and U2456 (N_2456,N_1939,N_1113);
or U2457 (N_2457,N_1980,N_1562);
and U2458 (N_2458,N_1986,N_1056);
or U2459 (N_2459,N_1906,N_1314);
and U2460 (N_2460,N_1770,N_1183);
xnor U2461 (N_2461,N_1441,N_1038);
or U2462 (N_2462,N_1760,N_1700);
nand U2463 (N_2463,N_1081,N_1680);
or U2464 (N_2464,N_1950,N_1005);
or U2465 (N_2465,N_1655,N_1216);
nand U2466 (N_2466,N_1105,N_1477);
xnor U2467 (N_2467,N_1841,N_1123);
nand U2468 (N_2468,N_1290,N_1403);
nor U2469 (N_2469,N_1667,N_1411);
and U2470 (N_2470,N_1159,N_1858);
and U2471 (N_2471,N_1165,N_1243);
and U2472 (N_2472,N_1578,N_1398);
and U2473 (N_2473,N_1886,N_1404);
or U2474 (N_2474,N_1799,N_1520);
nand U2475 (N_2475,N_1651,N_1444);
or U2476 (N_2476,N_1968,N_1851);
nand U2477 (N_2477,N_1867,N_1119);
xnor U2478 (N_2478,N_1956,N_1509);
or U2479 (N_2479,N_1067,N_1833);
nand U2480 (N_2480,N_1927,N_1622);
nand U2481 (N_2481,N_1874,N_1507);
and U2482 (N_2482,N_1876,N_1501);
nor U2483 (N_2483,N_1494,N_1425);
nor U2484 (N_2484,N_1713,N_1831);
and U2485 (N_2485,N_1826,N_1992);
or U2486 (N_2486,N_1969,N_1386);
nand U2487 (N_2487,N_1674,N_1001);
or U2488 (N_2488,N_1751,N_1972);
nand U2489 (N_2489,N_1267,N_1530);
and U2490 (N_2490,N_1812,N_1592);
and U2491 (N_2491,N_1057,N_1272);
and U2492 (N_2492,N_1508,N_1914);
or U2493 (N_2493,N_1778,N_1447);
and U2494 (N_2494,N_1689,N_1721);
xor U2495 (N_2495,N_1795,N_1635);
and U2496 (N_2496,N_1242,N_1748);
nand U2497 (N_2497,N_1396,N_1668);
and U2498 (N_2498,N_1265,N_1366);
and U2499 (N_2499,N_1834,N_1264);
and U2500 (N_2500,N_1032,N_1129);
nor U2501 (N_2501,N_1623,N_1994);
nand U2502 (N_2502,N_1905,N_1975);
xor U2503 (N_2503,N_1739,N_1888);
and U2504 (N_2504,N_1332,N_1347);
nor U2505 (N_2505,N_1303,N_1491);
xor U2506 (N_2506,N_1067,N_1419);
and U2507 (N_2507,N_1847,N_1737);
or U2508 (N_2508,N_1388,N_1652);
nand U2509 (N_2509,N_1884,N_1494);
and U2510 (N_2510,N_1626,N_1728);
or U2511 (N_2511,N_1849,N_1199);
nor U2512 (N_2512,N_1838,N_1739);
nand U2513 (N_2513,N_1477,N_1870);
or U2514 (N_2514,N_1044,N_1058);
nand U2515 (N_2515,N_1135,N_1902);
nand U2516 (N_2516,N_1067,N_1217);
and U2517 (N_2517,N_1288,N_1168);
nand U2518 (N_2518,N_1628,N_1800);
nor U2519 (N_2519,N_1913,N_1668);
or U2520 (N_2520,N_1089,N_1504);
and U2521 (N_2521,N_1862,N_1715);
or U2522 (N_2522,N_1825,N_1835);
nand U2523 (N_2523,N_1925,N_1374);
nor U2524 (N_2524,N_1530,N_1507);
nor U2525 (N_2525,N_1130,N_1973);
xor U2526 (N_2526,N_1944,N_1542);
nand U2527 (N_2527,N_1247,N_1603);
nand U2528 (N_2528,N_1727,N_1319);
or U2529 (N_2529,N_1146,N_1941);
and U2530 (N_2530,N_1350,N_1380);
nor U2531 (N_2531,N_1290,N_1114);
nand U2532 (N_2532,N_1648,N_1319);
xor U2533 (N_2533,N_1184,N_1431);
and U2534 (N_2534,N_1692,N_1364);
nor U2535 (N_2535,N_1363,N_1034);
nor U2536 (N_2536,N_1798,N_1887);
or U2537 (N_2537,N_1151,N_1130);
and U2538 (N_2538,N_1643,N_1981);
or U2539 (N_2539,N_1931,N_1517);
or U2540 (N_2540,N_1414,N_1686);
nand U2541 (N_2541,N_1531,N_1646);
and U2542 (N_2542,N_1108,N_1948);
nor U2543 (N_2543,N_1185,N_1754);
nand U2544 (N_2544,N_1977,N_1933);
xnor U2545 (N_2545,N_1275,N_1643);
or U2546 (N_2546,N_1368,N_1132);
nor U2547 (N_2547,N_1376,N_1895);
nor U2548 (N_2548,N_1702,N_1188);
and U2549 (N_2549,N_1131,N_1320);
or U2550 (N_2550,N_1715,N_1789);
nand U2551 (N_2551,N_1440,N_1566);
or U2552 (N_2552,N_1284,N_1519);
nor U2553 (N_2553,N_1786,N_1888);
or U2554 (N_2554,N_1619,N_1475);
nor U2555 (N_2555,N_1318,N_1094);
nor U2556 (N_2556,N_1736,N_1806);
and U2557 (N_2557,N_1339,N_1857);
and U2558 (N_2558,N_1443,N_1152);
nand U2559 (N_2559,N_1794,N_1912);
or U2560 (N_2560,N_1177,N_1627);
nor U2561 (N_2561,N_1150,N_1560);
and U2562 (N_2562,N_1186,N_1414);
or U2563 (N_2563,N_1198,N_1097);
xor U2564 (N_2564,N_1780,N_1416);
and U2565 (N_2565,N_1891,N_1386);
or U2566 (N_2566,N_1689,N_1936);
nand U2567 (N_2567,N_1758,N_1966);
nor U2568 (N_2568,N_1845,N_1220);
nand U2569 (N_2569,N_1338,N_1759);
nand U2570 (N_2570,N_1928,N_1551);
or U2571 (N_2571,N_1180,N_1621);
or U2572 (N_2572,N_1657,N_1371);
nand U2573 (N_2573,N_1359,N_1301);
nand U2574 (N_2574,N_1644,N_1423);
nor U2575 (N_2575,N_1208,N_1703);
nand U2576 (N_2576,N_1323,N_1030);
xor U2577 (N_2577,N_1122,N_1002);
and U2578 (N_2578,N_1659,N_1339);
xor U2579 (N_2579,N_1115,N_1499);
nor U2580 (N_2580,N_1014,N_1405);
nor U2581 (N_2581,N_1445,N_1429);
and U2582 (N_2582,N_1823,N_1613);
xnor U2583 (N_2583,N_1303,N_1572);
or U2584 (N_2584,N_1255,N_1903);
nand U2585 (N_2585,N_1329,N_1068);
nor U2586 (N_2586,N_1395,N_1282);
or U2587 (N_2587,N_1660,N_1120);
xor U2588 (N_2588,N_1081,N_1983);
or U2589 (N_2589,N_1068,N_1303);
or U2590 (N_2590,N_1869,N_1452);
nor U2591 (N_2591,N_1508,N_1075);
nor U2592 (N_2592,N_1633,N_1964);
xnor U2593 (N_2593,N_1007,N_1601);
xor U2594 (N_2594,N_1390,N_1765);
or U2595 (N_2595,N_1758,N_1045);
or U2596 (N_2596,N_1647,N_1478);
nor U2597 (N_2597,N_1177,N_1855);
and U2598 (N_2598,N_1296,N_1669);
nor U2599 (N_2599,N_1546,N_1492);
nor U2600 (N_2600,N_1063,N_1262);
nor U2601 (N_2601,N_1815,N_1262);
xor U2602 (N_2602,N_1950,N_1021);
or U2603 (N_2603,N_1959,N_1935);
xnor U2604 (N_2604,N_1233,N_1938);
and U2605 (N_2605,N_1043,N_1120);
xor U2606 (N_2606,N_1878,N_1989);
nand U2607 (N_2607,N_1495,N_1830);
nand U2608 (N_2608,N_1598,N_1604);
and U2609 (N_2609,N_1897,N_1810);
xnor U2610 (N_2610,N_1848,N_1733);
nand U2611 (N_2611,N_1780,N_1157);
xnor U2612 (N_2612,N_1779,N_1106);
or U2613 (N_2613,N_1996,N_1919);
nor U2614 (N_2614,N_1447,N_1192);
nand U2615 (N_2615,N_1098,N_1556);
or U2616 (N_2616,N_1371,N_1530);
and U2617 (N_2617,N_1624,N_1629);
xor U2618 (N_2618,N_1345,N_1932);
and U2619 (N_2619,N_1608,N_1658);
xnor U2620 (N_2620,N_1846,N_1852);
and U2621 (N_2621,N_1145,N_1802);
xnor U2622 (N_2622,N_1673,N_1971);
nand U2623 (N_2623,N_1118,N_1394);
xnor U2624 (N_2624,N_1843,N_1755);
nor U2625 (N_2625,N_1849,N_1880);
and U2626 (N_2626,N_1470,N_1571);
nor U2627 (N_2627,N_1143,N_1109);
nand U2628 (N_2628,N_1310,N_1132);
or U2629 (N_2629,N_1054,N_1255);
nor U2630 (N_2630,N_1816,N_1079);
and U2631 (N_2631,N_1451,N_1756);
nand U2632 (N_2632,N_1698,N_1649);
xor U2633 (N_2633,N_1723,N_1426);
and U2634 (N_2634,N_1790,N_1026);
nor U2635 (N_2635,N_1009,N_1991);
nand U2636 (N_2636,N_1236,N_1841);
and U2637 (N_2637,N_1477,N_1388);
nand U2638 (N_2638,N_1783,N_1750);
xor U2639 (N_2639,N_1806,N_1300);
nand U2640 (N_2640,N_1095,N_1532);
or U2641 (N_2641,N_1604,N_1435);
xnor U2642 (N_2642,N_1707,N_1617);
or U2643 (N_2643,N_1858,N_1442);
nand U2644 (N_2644,N_1757,N_1495);
and U2645 (N_2645,N_1406,N_1049);
nor U2646 (N_2646,N_1659,N_1631);
xnor U2647 (N_2647,N_1603,N_1360);
nor U2648 (N_2648,N_1841,N_1886);
and U2649 (N_2649,N_1770,N_1393);
or U2650 (N_2650,N_1082,N_1446);
nand U2651 (N_2651,N_1024,N_1873);
xor U2652 (N_2652,N_1048,N_1952);
xnor U2653 (N_2653,N_1428,N_1631);
nand U2654 (N_2654,N_1954,N_1608);
nand U2655 (N_2655,N_1012,N_1702);
and U2656 (N_2656,N_1922,N_1086);
and U2657 (N_2657,N_1519,N_1199);
xnor U2658 (N_2658,N_1651,N_1099);
nand U2659 (N_2659,N_1307,N_1515);
nor U2660 (N_2660,N_1889,N_1511);
or U2661 (N_2661,N_1791,N_1007);
and U2662 (N_2662,N_1799,N_1397);
or U2663 (N_2663,N_1893,N_1467);
or U2664 (N_2664,N_1205,N_1944);
nor U2665 (N_2665,N_1383,N_1005);
nor U2666 (N_2666,N_1910,N_1082);
nand U2667 (N_2667,N_1588,N_1110);
or U2668 (N_2668,N_1440,N_1400);
and U2669 (N_2669,N_1441,N_1751);
or U2670 (N_2670,N_1379,N_1135);
xor U2671 (N_2671,N_1551,N_1636);
nand U2672 (N_2672,N_1483,N_1441);
or U2673 (N_2673,N_1248,N_1892);
or U2674 (N_2674,N_1597,N_1347);
or U2675 (N_2675,N_1094,N_1005);
nand U2676 (N_2676,N_1933,N_1698);
or U2677 (N_2677,N_1227,N_1960);
and U2678 (N_2678,N_1650,N_1771);
and U2679 (N_2679,N_1982,N_1560);
nor U2680 (N_2680,N_1186,N_1021);
nand U2681 (N_2681,N_1560,N_1007);
xor U2682 (N_2682,N_1216,N_1426);
nor U2683 (N_2683,N_1874,N_1856);
xor U2684 (N_2684,N_1529,N_1340);
nand U2685 (N_2685,N_1735,N_1763);
xor U2686 (N_2686,N_1250,N_1949);
xor U2687 (N_2687,N_1511,N_1589);
nand U2688 (N_2688,N_1854,N_1137);
nor U2689 (N_2689,N_1971,N_1087);
xnor U2690 (N_2690,N_1727,N_1126);
nand U2691 (N_2691,N_1853,N_1139);
nor U2692 (N_2692,N_1557,N_1166);
nand U2693 (N_2693,N_1639,N_1020);
nand U2694 (N_2694,N_1828,N_1810);
and U2695 (N_2695,N_1591,N_1449);
and U2696 (N_2696,N_1017,N_1390);
nand U2697 (N_2697,N_1445,N_1819);
nand U2698 (N_2698,N_1569,N_1851);
nand U2699 (N_2699,N_1677,N_1042);
and U2700 (N_2700,N_1763,N_1186);
nand U2701 (N_2701,N_1546,N_1836);
nor U2702 (N_2702,N_1864,N_1913);
and U2703 (N_2703,N_1162,N_1290);
and U2704 (N_2704,N_1498,N_1776);
nand U2705 (N_2705,N_1221,N_1445);
or U2706 (N_2706,N_1214,N_1796);
xnor U2707 (N_2707,N_1234,N_1124);
nand U2708 (N_2708,N_1599,N_1870);
and U2709 (N_2709,N_1508,N_1657);
nor U2710 (N_2710,N_1697,N_1242);
xnor U2711 (N_2711,N_1255,N_1035);
or U2712 (N_2712,N_1633,N_1903);
nor U2713 (N_2713,N_1702,N_1367);
nor U2714 (N_2714,N_1046,N_1107);
and U2715 (N_2715,N_1375,N_1453);
and U2716 (N_2716,N_1904,N_1606);
and U2717 (N_2717,N_1888,N_1948);
or U2718 (N_2718,N_1480,N_1909);
nor U2719 (N_2719,N_1592,N_1420);
or U2720 (N_2720,N_1425,N_1844);
nor U2721 (N_2721,N_1894,N_1116);
xor U2722 (N_2722,N_1209,N_1518);
nand U2723 (N_2723,N_1064,N_1210);
nand U2724 (N_2724,N_1716,N_1044);
or U2725 (N_2725,N_1600,N_1530);
nand U2726 (N_2726,N_1680,N_1718);
xor U2727 (N_2727,N_1201,N_1489);
and U2728 (N_2728,N_1252,N_1952);
or U2729 (N_2729,N_1947,N_1545);
xor U2730 (N_2730,N_1452,N_1684);
and U2731 (N_2731,N_1827,N_1079);
nor U2732 (N_2732,N_1212,N_1541);
and U2733 (N_2733,N_1664,N_1183);
and U2734 (N_2734,N_1115,N_1333);
nand U2735 (N_2735,N_1937,N_1820);
nand U2736 (N_2736,N_1892,N_1390);
nor U2737 (N_2737,N_1383,N_1001);
and U2738 (N_2738,N_1663,N_1324);
nand U2739 (N_2739,N_1226,N_1333);
nand U2740 (N_2740,N_1521,N_1658);
xor U2741 (N_2741,N_1981,N_1726);
and U2742 (N_2742,N_1589,N_1685);
nor U2743 (N_2743,N_1025,N_1789);
and U2744 (N_2744,N_1596,N_1260);
and U2745 (N_2745,N_1103,N_1301);
and U2746 (N_2746,N_1340,N_1933);
and U2747 (N_2747,N_1313,N_1889);
or U2748 (N_2748,N_1885,N_1491);
and U2749 (N_2749,N_1048,N_1959);
and U2750 (N_2750,N_1744,N_1465);
and U2751 (N_2751,N_1899,N_1512);
and U2752 (N_2752,N_1951,N_1175);
or U2753 (N_2753,N_1791,N_1071);
and U2754 (N_2754,N_1437,N_1590);
nor U2755 (N_2755,N_1190,N_1595);
xor U2756 (N_2756,N_1343,N_1847);
nor U2757 (N_2757,N_1954,N_1547);
nor U2758 (N_2758,N_1893,N_1353);
and U2759 (N_2759,N_1345,N_1899);
or U2760 (N_2760,N_1567,N_1466);
nor U2761 (N_2761,N_1471,N_1361);
or U2762 (N_2762,N_1965,N_1763);
nor U2763 (N_2763,N_1245,N_1236);
nor U2764 (N_2764,N_1530,N_1585);
nor U2765 (N_2765,N_1592,N_1424);
nor U2766 (N_2766,N_1029,N_1448);
nand U2767 (N_2767,N_1199,N_1977);
nor U2768 (N_2768,N_1502,N_1929);
or U2769 (N_2769,N_1431,N_1787);
or U2770 (N_2770,N_1905,N_1493);
nand U2771 (N_2771,N_1527,N_1939);
and U2772 (N_2772,N_1140,N_1904);
nand U2773 (N_2773,N_1669,N_1899);
or U2774 (N_2774,N_1683,N_1984);
and U2775 (N_2775,N_1323,N_1893);
and U2776 (N_2776,N_1515,N_1563);
nor U2777 (N_2777,N_1940,N_1275);
xnor U2778 (N_2778,N_1495,N_1401);
nand U2779 (N_2779,N_1917,N_1924);
nor U2780 (N_2780,N_1008,N_1644);
and U2781 (N_2781,N_1698,N_1174);
xnor U2782 (N_2782,N_1602,N_1499);
xor U2783 (N_2783,N_1499,N_1752);
xor U2784 (N_2784,N_1000,N_1737);
or U2785 (N_2785,N_1301,N_1370);
or U2786 (N_2786,N_1828,N_1233);
xor U2787 (N_2787,N_1608,N_1839);
and U2788 (N_2788,N_1292,N_1372);
or U2789 (N_2789,N_1232,N_1687);
xor U2790 (N_2790,N_1716,N_1306);
nand U2791 (N_2791,N_1109,N_1168);
nor U2792 (N_2792,N_1556,N_1495);
xor U2793 (N_2793,N_1917,N_1871);
and U2794 (N_2794,N_1428,N_1127);
and U2795 (N_2795,N_1195,N_1511);
nand U2796 (N_2796,N_1969,N_1174);
or U2797 (N_2797,N_1753,N_1978);
nor U2798 (N_2798,N_1712,N_1553);
nor U2799 (N_2799,N_1241,N_1599);
nor U2800 (N_2800,N_1823,N_1713);
nor U2801 (N_2801,N_1312,N_1748);
and U2802 (N_2802,N_1191,N_1432);
xnor U2803 (N_2803,N_1098,N_1912);
nand U2804 (N_2804,N_1824,N_1847);
and U2805 (N_2805,N_1058,N_1343);
nand U2806 (N_2806,N_1244,N_1240);
nor U2807 (N_2807,N_1759,N_1384);
xnor U2808 (N_2808,N_1924,N_1159);
or U2809 (N_2809,N_1375,N_1522);
and U2810 (N_2810,N_1424,N_1231);
xor U2811 (N_2811,N_1707,N_1928);
xnor U2812 (N_2812,N_1503,N_1137);
xor U2813 (N_2813,N_1958,N_1944);
or U2814 (N_2814,N_1833,N_1626);
nor U2815 (N_2815,N_1560,N_1371);
nand U2816 (N_2816,N_1252,N_1404);
nand U2817 (N_2817,N_1659,N_1870);
xor U2818 (N_2818,N_1817,N_1627);
or U2819 (N_2819,N_1805,N_1800);
and U2820 (N_2820,N_1037,N_1238);
xnor U2821 (N_2821,N_1104,N_1986);
xor U2822 (N_2822,N_1733,N_1113);
nor U2823 (N_2823,N_1626,N_1163);
nor U2824 (N_2824,N_1021,N_1196);
xor U2825 (N_2825,N_1181,N_1180);
and U2826 (N_2826,N_1113,N_1622);
nor U2827 (N_2827,N_1095,N_1450);
nor U2828 (N_2828,N_1187,N_1301);
and U2829 (N_2829,N_1662,N_1916);
nand U2830 (N_2830,N_1488,N_1993);
nor U2831 (N_2831,N_1900,N_1468);
nand U2832 (N_2832,N_1038,N_1934);
nor U2833 (N_2833,N_1128,N_1721);
xnor U2834 (N_2834,N_1231,N_1775);
nand U2835 (N_2835,N_1902,N_1604);
xnor U2836 (N_2836,N_1363,N_1806);
or U2837 (N_2837,N_1624,N_1660);
and U2838 (N_2838,N_1298,N_1412);
or U2839 (N_2839,N_1882,N_1575);
nand U2840 (N_2840,N_1678,N_1239);
or U2841 (N_2841,N_1066,N_1039);
or U2842 (N_2842,N_1925,N_1245);
or U2843 (N_2843,N_1553,N_1225);
or U2844 (N_2844,N_1919,N_1520);
or U2845 (N_2845,N_1641,N_1348);
xnor U2846 (N_2846,N_1437,N_1430);
or U2847 (N_2847,N_1117,N_1634);
xnor U2848 (N_2848,N_1838,N_1275);
or U2849 (N_2849,N_1668,N_1494);
and U2850 (N_2850,N_1081,N_1561);
and U2851 (N_2851,N_1501,N_1589);
nand U2852 (N_2852,N_1780,N_1700);
and U2853 (N_2853,N_1008,N_1909);
and U2854 (N_2854,N_1625,N_1364);
xor U2855 (N_2855,N_1210,N_1926);
nor U2856 (N_2856,N_1997,N_1690);
and U2857 (N_2857,N_1792,N_1094);
and U2858 (N_2858,N_1699,N_1865);
xor U2859 (N_2859,N_1723,N_1647);
or U2860 (N_2860,N_1484,N_1240);
nand U2861 (N_2861,N_1716,N_1859);
nand U2862 (N_2862,N_1508,N_1809);
nor U2863 (N_2863,N_1486,N_1801);
nor U2864 (N_2864,N_1672,N_1737);
xnor U2865 (N_2865,N_1467,N_1093);
nor U2866 (N_2866,N_1437,N_1478);
and U2867 (N_2867,N_1072,N_1727);
nand U2868 (N_2868,N_1413,N_1672);
or U2869 (N_2869,N_1494,N_1303);
nand U2870 (N_2870,N_1428,N_1887);
nor U2871 (N_2871,N_1040,N_1229);
or U2872 (N_2872,N_1907,N_1542);
nand U2873 (N_2873,N_1703,N_1413);
xnor U2874 (N_2874,N_1627,N_1415);
xor U2875 (N_2875,N_1063,N_1633);
and U2876 (N_2876,N_1917,N_1665);
nand U2877 (N_2877,N_1490,N_1657);
xnor U2878 (N_2878,N_1790,N_1583);
nand U2879 (N_2879,N_1969,N_1238);
or U2880 (N_2880,N_1095,N_1077);
xnor U2881 (N_2881,N_1833,N_1887);
nor U2882 (N_2882,N_1215,N_1880);
or U2883 (N_2883,N_1016,N_1621);
nor U2884 (N_2884,N_1021,N_1051);
nand U2885 (N_2885,N_1833,N_1999);
nor U2886 (N_2886,N_1242,N_1563);
nor U2887 (N_2887,N_1409,N_1961);
or U2888 (N_2888,N_1501,N_1388);
and U2889 (N_2889,N_1014,N_1866);
xor U2890 (N_2890,N_1817,N_1012);
or U2891 (N_2891,N_1905,N_1982);
and U2892 (N_2892,N_1934,N_1734);
and U2893 (N_2893,N_1966,N_1480);
nand U2894 (N_2894,N_1240,N_1755);
and U2895 (N_2895,N_1279,N_1264);
nor U2896 (N_2896,N_1426,N_1572);
and U2897 (N_2897,N_1389,N_1359);
nand U2898 (N_2898,N_1125,N_1141);
and U2899 (N_2899,N_1525,N_1092);
nand U2900 (N_2900,N_1024,N_1077);
and U2901 (N_2901,N_1303,N_1791);
and U2902 (N_2902,N_1915,N_1771);
nand U2903 (N_2903,N_1931,N_1606);
nand U2904 (N_2904,N_1912,N_1230);
nand U2905 (N_2905,N_1227,N_1539);
nand U2906 (N_2906,N_1003,N_1140);
nor U2907 (N_2907,N_1913,N_1978);
xor U2908 (N_2908,N_1466,N_1390);
and U2909 (N_2909,N_1947,N_1708);
nand U2910 (N_2910,N_1048,N_1579);
and U2911 (N_2911,N_1991,N_1728);
nor U2912 (N_2912,N_1022,N_1780);
and U2913 (N_2913,N_1086,N_1161);
nand U2914 (N_2914,N_1213,N_1898);
or U2915 (N_2915,N_1907,N_1215);
nand U2916 (N_2916,N_1327,N_1691);
xnor U2917 (N_2917,N_1509,N_1399);
nor U2918 (N_2918,N_1117,N_1755);
nor U2919 (N_2919,N_1961,N_1248);
nor U2920 (N_2920,N_1322,N_1780);
or U2921 (N_2921,N_1192,N_1940);
or U2922 (N_2922,N_1536,N_1741);
and U2923 (N_2923,N_1149,N_1993);
and U2924 (N_2924,N_1373,N_1832);
or U2925 (N_2925,N_1935,N_1761);
nor U2926 (N_2926,N_1184,N_1884);
xor U2927 (N_2927,N_1576,N_1033);
or U2928 (N_2928,N_1791,N_1045);
xor U2929 (N_2929,N_1355,N_1249);
nor U2930 (N_2930,N_1373,N_1671);
nand U2931 (N_2931,N_1587,N_1244);
and U2932 (N_2932,N_1374,N_1833);
xor U2933 (N_2933,N_1113,N_1097);
and U2934 (N_2934,N_1693,N_1370);
xnor U2935 (N_2935,N_1332,N_1890);
xnor U2936 (N_2936,N_1772,N_1768);
nor U2937 (N_2937,N_1049,N_1630);
nor U2938 (N_2938,N_1832,N_1199);
nand U2939 (N_2939,N_1091,N_1748);
nor U2940 (N_2940,N_1796,N_1464);
nor U2941 (N_2941,N_1759,N_1325);
nor U2942 (N_2942,N_1719,N_1974);
nor U2943 (N_2943,N_1233,N_1442);
nor U2944 (N_2944,N_1902,N_1537);
xnor U2945 (N_2945,N_1738,N_1962);
nand U2946 (N_2946,N_1698,N_1226);
or U2947 (N_2947,N_1897,N_1340);
xnor U2948 (N_2948,N_1343,N_1732);
nor U2949 (N_2949,N_1381,N_1034);
or U2950 (N_2950,N_1087,N_1361);
and U2951 (N_2951,N_1916,N_1789);
nand U2952 (N_2952,N_1118,N_1983);
xor U2953 (N_2953,N_1970,N_1309);
xnor U2954 (N_2954,N_1866,N_1055);
and U2955 (N_2955,N_1884,N_1707);
xnor U2956 (N_2956,N_1158,N_1869);
nor U2957 (N_2957,N_1058,N_1365);
or U2958 (N_2958,N_1731,N_1674);
nor U2959 (N_2959,N_1274,N_1834);
or U2960 (N_2960,N_1406,N_1700);
xnor U2961 (N_2961,N_1308,N_1775);
nand U2962 (N_2962,N_1890,N_1077);
nand U2963 (N_2963,N_1805,N_1156);
and U2964 (N_2964,N_1993,N_1343);
or U2965 (N_2965,N_1589,N_1298);
or U2966 (N_2966,N_1855,N_1208);
and U2967 (N_2967,N_1819,N_1683);
or U2968 (N_2968,N_1392,N_1325);
xnor U2969 (N_2969,N_1674,N_1144);
xor U2970 (N_2970,N_1590,N_1774);
nor U2971 (N_2971,N_1121,N_1660);
nand U2972 (N_2972,N_1836,N_1164);
nand U2973 (N_2973,N_1938,N_1369);
xor U2974 (N_2974,N_1485,N_1101);
or U2975 (N_2975,N_1711,N_1414);
or U2976 (N_2976,N_1075,N_1102);
xnor U2977 (N_2977,N_1120,N_1383);
xor U2978 (N_2978,N_1958,N_1150);
and U2979 (N_2979,N_1633,N_1448);
and U2980 (N_2980,N_1426,N_1045);
xor U2981 (N_2981,N_1202,N_1885);
nand U2982 (N_2982,N_1168,N_1213);
and U2983 (N_2983,N_1276,N_1989);
and U2984 (N_2984,N_1318,N_1777);
xor U2985 (N_2985,N_1277,N_1612);
nand U2986 (N_2986,N_1638,N_1190);
and U2987 (N_2987,N_1035,N_1107);
xnor U2988 (N_2988,N_1690,N_1166);
xnor U2989 (N_2989,N_1100,N_1201);
nand U2990 (N_2990,N_1965,N_1977);
or U2991 (N_2991,N_1478,N_1227);
nand U2992 (N_2992,N_1577,N_1070);
xor U2993 (N_2993,N_1189,N_1715);
xor U2994 (N_2994,N_1512,N_1677);
or U2995 (N_2995,N_1920,N_1598);
and U2996 (N_2996,N_1899,N_1895);
and U2997 (N_2997,N_1235,N_1587);
nand U2998 (N_2998,N_1987,N_1860);
or U2999 (N_2999,N_1346,N_1601);
nor U3000 (N_3000,N_2857,N_2910);
nand U3001 (N_3001,N_2337,N_2202);
and U3002 (N_3002,N_2347,N_2112);
and U3003 (N_3003,N_2691,N_2843);
or U3004 (N_3004,N_2904,N_2236);
or U3005 (N_3005,N_2056,N_2139);
or U3006 (N_3006,N_2512,N_2585);
nor U3007 (N_3007,N_2958,N_2976);
xor U3008 (N_3008,N_2987,N_2468);
xnor U3009 (N_3009,N_2162,N_2802);
and U3010 (N_3010,N_2306,N_2426);
xor U3011 (N_3011,N_2445,N_2128);
and U3012 (N_3012,N_2997,N_2535);
nand U3013 (N_3013,N_2772,N_2725);
nor U3014 (N_3014,N_2416,N_2927);
xor U3015 (N_3015,N_2825,N_2200);
nor U3016 (N_3016,N_2109,N_2875);
and U3017 (N_3017,N_2149,N_2562);
nor U3018 (N_3018,N_2052,N_2407);
or U3019 (N_3019,N_2751,N_2208);
nand U3020 (N_3020,N_2756,N_2786);
and U3021 (N_3021,N_2061,N_2113);
or U3022 (N_3022,N_2408,N_2321);
nand U3023 (N_3023,N_2338,N_2980);
nand U3024 (N_3024,N_2260,N_2367);
nand U3025 (N_3025,N_2131,N_2308);
or U3026 (N_3026,N_2066,N_2862);
nand U3027 (N_3027,N_2286,N_2495);
or U3028 (N_3028,N_2433,N_2929);
nor U3029 (N_3029,N_2784,N_2329);
nand U3030 (N_3030,N_2753,N_2489);
nand U3031 (N_3031,N_2313,N_2093);
nor U3032 (N_3032,N_2838,N_2783);
nand U3033 (N_3033,N_2741,N_2292);
and U3034 (N_3034,N_2203,N_2287);
xnor U3035 (N_3035,N_2371,N_2404);
nor U3036 (N_3036,N_2546,N_2595);
xnor U3037 (N_3037,N_2581,N_2606);
or U3038 (N_3038,N_2799,N_2171);
or U3039 (N_3039,N_2041,N_2881);
nor U3040 (N_3040,N_2948,N_2818);
xnor U3041 (N_3041,N_2637,N_2084);
xor U3042 (N_3042,N_2919,N_2339);
nor U3043 (N_3043,N_2536,N_2365);
or U3044 (N_3044,N_2004,N_2739);
nand U3045 (N_3045,N_2370,N_2067);
and U3046 (N_3046,N_2985,N_2696);
and U3047 (N_3047,N_2280,N_2971);
nand U3048 (N_3048,N_2269,N_2608);
nor U3049 (N_3049,N_2417,N_2749);
nor U3050 (N_3050,N_2704,N_2024);
nand U3051 (N_3051,N_2928,N_2110);
and U3052 (N_3052,N_2556,N_2373);
or U3053 (N_3053,N_2392,N_2653);
or U3054 (N_3054,N_2632,N_2310);
xnor U3055 (N_3055,N_2973,N_2516);
or U3056 (N_3056,N_2558,N_2156);
and U3057 (N_3057,N_2678,N_2685);
nor U3058 (N_3058,N_2413,N_2053);
and U3059 (N_3059,N_2335,N_2713);
xor U3060 (N_3060,N_2554,N_2430);
and U3061 (N_3061,N_2796,N_2146);
or U3062 (N_3062,N_2577,N_2550);
nand U3063 (N_3063,N_2646,N_2226);
nor U3064 (N_3064,N_2745,N_2301);
nand U3065 (N_3065,N_2791,N_2450);
xnor U3066 (N_3066,N_2331,N_2220);
and U3067 (N_3067,N_2769,N_2458);
nand U3068 (N_3068,N_2587,N_2641);
xor U3069 (N_3069,N_2699,N_2240);
xnor U3070 (N_3070,N_2356,N_2094);
nor U3071 (N_3071,N_2455,N_2659);
nand U3072 (N_3072,N_2000,N_2435);
and U3073 (N_3073,N_2235,N_2628);
xnor U3074 (N_3074,N_2410,N_2199);
and U3075 (N_3075,N_2573,N_2603);
xor U3076 (N_3076,N_2654,N_2572);
xnor U3077 (N_3077,N_2798,N_2499);
nand U3078 (N_3078,N_2531,N_2873);
or U3079 (N_3079,N_2528,N_2377);
or U3080 (N_3080,N_2174,N_2995);
or U3081 (N_3081,N_2831,N_2944);
or U3082 (N_3082,N_2490,N_2500);
or U3083 (N_3083,N_2661,N_2736);
nor U3084 (N_3084,N_2157,N_2049);
xnor U3085 (N_3085,N_2775,N_2609);
and U3086 (N_3086,N_2778,N_2497);
xor U3087 (N_3087,N_2938,N_2349);
xnor U3088 (N_3088,N_2780,N_2728);
xor U3089 (N_3089,N_2115,N_2075);
nand U3090 (N_3090,N_2185,N_2925);
nand U3091 (N_3091,N_2465,N_2544);
nor U3092 (N_3092,N_2690,N_2363);
nor U3093 (N_3093,N_2529,N_2820);
nor U3094 (N_3094,N_2727,N_2770);
xor U3095 (N_3095,N_2511,N_2350);
and U3096 (N_3096,N_2627,N_2255);
nor U3097 (N_3097,N_2635,N_2638);
nor U3098 (N_3098,N_2817,N_2334);
nor U3099 (N_3099,N_2640,N_2238);
nor U3100 (N_3100,N_2452,N_2340);
and U3101 (N_3101,N_2719,N_2265);
xor U3102 (N_3102,N_2785,N_2126);
or U3103 (N_3103,N_2908,N_2001);
and U3104 (N_3104,N_2057,N_2506);
nor U3105 (N_3105,N_2853,N_2823);
and U3106 (N_3106,N_2933,N_2808);
nor U3107 (N_3107,N_2989,N_2117);
or U3108 (N_3108,N_2935,N_2723);
xor U3109 (N_3109,N_2805,N_2724);
xor U3110 (N_3110,N_2328,N_2680);
nor U3111 (N_3111,N_2731,N_2836);
nand U3112 (N_3112,N_2038,N_2217);
or U3113 (N_3113,N_2423,N_2742);
and U3114 (N_3114,N_2624,N_2754);
or U3115 (N_3115,N_2906,N_2574);
or U3116 (N_3116,N_2681,N_2854);
xor U3117 (N_3117,N_2463,N_2721);
nor U3118 (N_3118,N_2237,N_2806);
nor U3119 (N_3119,N_2257,N_2522);
and U3120 (N_3120,N_2387,N_2332);
and U3121 (N_3121,N_2002,N_2341);
nand U3122 (N_3122,N_2912,N_2104);
and U3123 (N_3123,N_2323,N_2224);
xor U3124 (N_3124,N_2982,N_2665);
and U3125 (N_3125,N_2402,N_2955);
nor U3126 (N_3126,N_2856,N_2144);
nor U3127 (N_3127,N_2429,N_2623);
xor U3128 (N_3128,N_2662,N_2504);
or U3129 (N_3129,N_2846,N_2384);
or U3130 (N_3130,N_2524,N_2896);
nand U3131 (N_3131,N_2189,N_2582);
or U3132 (N_3132,N_2801,N_2663);
xor U3133 (N_3133,N_2390,N_2018);
xor U3134 (N_3134,N_2172,N_2821);
xor U3135 (N_3135,N_2372,N_2954);
and U3136 (N_3136,N_2295,N_2999);
xor U3137 (N_3137,N_2277,N_2447);
nand U3138 (N_3138,N_2108,N_2601);
and U3139 (N_3139,N_2893,N_2949);
nor U3140 (N_3140,N_2619,N_2448);
or U3141 (N_3141,N_2466,N_2814);
xnor U3142 (N_3142,N_2686,N_2182);
and U3143 (N_3143,N_2412,N_2965);
nand U3144 (N_3144,N_2563,N_2752);
nor U3145 (N_3145,N_2552,N_2884);
and U3146 (N_3146,N_2205,N_2923);
and U3147 (N_3147,N_2121,N_2660);
and U3148 (N_3148,N_2300,N_2311);
or U3149 (N_3149,N_2254,N_2122);
or U3150 (N_3150,N_2688,N_2030);
and U3151 (N_3151,N_2243,N_2193);
nor U3152 (N_3152,N_2682,N_2278);
or U3153 (N_3153,N_2209,N_2726);
or U3154 (N_3154,N_2969,N_2705);
nand U3155 (N_3155,N_2656,N_2083);
nor U3156 (N_3156,N_2730,N_2293);
nor U3157 (N_3157,N_2936,N_2568);
and U3158 (N_3158,N_2848,N_2178);
and U3159 (N_3159,N_2720,N_2086);
xor U3160 (N_3160,N_2503,N_2451);
and U3161 (N_3161,N_2129,N_2716);
and U3162 (N_3162,N_2596,N_2434);
and U3163 (N_3163,N_2667,N_2441);
xor U3164 (N_3164,N_2670,N_2180);
nand U3165 (N_3165,N_2732,N_2618);
nand U3166 (N_3166,N_2953,N_2625);
and U3167 (N_3167,N_2080,N_2557);
or U3168 (N_3168,N_2804,N_2258);
xor U3169 (N_3169,N_2227,N_2461);
nand U3170 (N_3170,N_2526,N_2011);
nand U3171 (N_3171,N_2211,N_2252);
xnor U3172 (N_3172,N_2829,N_2366);
nand U3173 (N_3173,N_2124,N_2270);
or U3174 (N_3174,N_2415,N_2324);
xnor U3175 (N_3175,N_2879,N_2797);
xor U3176 (N_3176,N_2963,N_2476);
nand U3177 (N_3177,N_2070,N_2263);
and U3178 (N_3178,N_2352,N_2613);
or U3179 (N_3179,N_2414,N_2368);
nor U3180 (N_3180,N_2871,N_2034);
xor U3181 (N_3181,N_2859,N_2855);
nand U3182 (N_3182,N_2941,N_2822);
or U3183 (N_3183,N_2702,N_2042);
and U3184 (N_3184,N_2133,N_2216);
or U3185 (N_3185,N_2147,N_2130);
nor U3186 (N_3186,N_2249,N_2863);
nand U3187 (N_3187,N_2920,N_2065);
nor U3188 (N_3188,N_2584,N_2251);
and U3189 (N_3189,N_2138,N_2865);
nor U3190 (N_3190,N_2677,N_2136);
xor U3191 (N_3191,N_2790,N_2816);
and U3192 (N_3192,N_2343,N_2118);
nand U3193 (N_3193,N_2082,N_2733);
nand U3194 (N_3194,N_2353,N_2488);
and U3195 (N_3195,N_2326,N_2210);
xor U3196 (N_3196,N_2959,N_2593);
xnor U3197 (N_3197,N_2446,N_2457);
or U3198 (N_3198,N_2247,N_2355);
nor U3199 (N_3199,N_2917,N_2740);
or U3200 (N_3200,N_2703,N_2974);
xnor U3201 (N_3201,N_2545,N_2116);
nor U3202 (N_3202,N_2089,N_2899);
and U3203 (N_3203,N_2932,N_2234);
xnor U3204 (N_3204,N_2222,N_2979);
and U3205 (N_3205,N_2383,N_2943);
xnor U3206 (N_3206,N_2394,N_2764);
and U3207 (N_3207,N_2327,N_2271);
and U3208 (N_3208,N_2244,N_2901);
xnor U3209 (N_3209,N_2267,N_2945);
and U3210 (N_3210,N_2962,N_2657);
xor U3211 (N_3211,N_2225,N_2239);
nand U3212 (N_3212,N_2847,N_2968);
or U3213 (N_3213,N_2097,N_2296);
nand U3214 (N_3214,N_2760,N_2456);
nor U3215 (N_3215,N_2059,N_2464);
nand U3216 (N_3216,N_2190,N_2651);
and U3217 (N_3217,N_2718,N_2420);
xnor U3218 (N_3218,N_2253,N_2330);
nor U3219 (N_3219,N_2406,N_2792);
or U3220 (N_3220,N_2709,N_2614);
or U3221 (N_3221,N_2622,N_2275);
or U3222 (N_3222,N_2044,N_2081);
and U3223 (N_3223,N_2553,N_2409);
nand U3224 (N_3224,N_2167,N_2787);
and U3225 (N_3225,N_2400,N_2824);
nor U3226 (N_3226,N_2914,N_2187);
nor U3227 (N_3227,N_2303,N_2348);
xnor U3228 (N_3228,N_2826,N_2501);
xor U3229 (N_3229,N_2592,N_2950);
nand U3230 (N_3230,N_2639,N_2570);
or U3231 (N_3231,N_2530,N_2523);
nor U3232 (N_3232,N_2679,N_2119);
nor U3233 (N_3233,N_2284,N_2454);
nor U3234 (N_3234,N_2360,N_2107);
nor U3235 (N_3235,N_2135,N_2812);
nand U3236 (N_3236,N_2045,N_2207);
nor U3237 (N_3237,N_2514,N_2842);
nor U3238 (N_3238,N_2449,N_2715);
xor U3239 (N_3239,N_2915,N_2421);
nor U3240 (N_3240,N_2378,N_2706);
nand U3241 (N_3241,N_2977,N_2469);
xnor U3242 (N_3242,N_2453,N_2695);
nand U3243 (N_3243,N_2114,N_2777);
nand U3244 (N_3244,N_2970,N_2440);
and U3245 (N_3245,N_2380,N_2892);
and U3246 (N_3246,N_2229,N_2898);
nor U3247 (N_3247,N_2642,N_2100);
nor U3248 (N_3248,N_2242,N_2694);
xor U3249 (N_3249,N_2984,N_2233);
nor U3250 (N_3250,N_2291,N_2096);
and U3251 (N_3251,N_2911,N_2050);
or U3252 (N_3252,N_2960,N_2576);
nor U3253 (N_3253,N_2425,N_2273);
nand U3254 (N_3254,N_2611,N_2776);
xnor U3255 (N_3255,N_2975,N_2201);
and U3256 (N_3256,N_2714,N_2054);
nand U3257 (N_3257,N_2027,N_2952);
nand U3258 (N_3258,N_2035,N_2781);
xor U3259 (N_3259,N_2532,N_2895);
xor U3260 (N_3260,N_2290,N_2850);
or U3261 (N_3261,N_2946,N_2498);
nand U3262 (N_3262,N_2598,N_2722);
nor U3263 (N_3263,N_2548,N_2106);
and U3264 (N_3264,N_2525,N_2362);
or U3265 (N_3265,N_2262,N_2833);
nor U3266 (N_3266,N_2259,N_2837);
nand U3267 (N_3267,N_2612,N_2849);
or U3268 (N_3268,N_2840,N_2886);
nor U3269 (N_3269,N_2245,N_2605);
or U3270 (N_3270,N_2029,N_2077);
nor U3271 (N_3271,N_2020,N_2674);
and U3272 (N_3272,N_2230,N_2708);
and U3273 (N_3273,N_2496,N_2759);
and U3274 (N_3274,N_2386,N_2513);
xnor U3275 (N_3275,N_2757,N_2521);
nand U3276 (N_3276,N_2482,N_2068);
xnor U3277 (N_3277,N_2540,N_2916);
or U3278 (N_3278,N_2747,N_2160);
and U3279 (N_3279,N_2502,N_2152);
or U3280 (N_3280,N_2811,N_2462);
and U3281 (N_3281,N_2852,N_2918);
or U3282 (N_3282,N_2697,N_2650);
nor U3283 (N_3283,N_2023,N_2994);
nand U3284 (N_3284,N_2436,N_2610);
xnor U3285 (N_3285,N_2891,N_2957);
and U3286 (N_3286,N_2173,N_2604);
nand U3287 (N_3287,N_2634,N_2319);
xor U3288 (N_3288,N_2900,N_2008);
and U3289 (N_3289,N_2062,N_2316);
xnor U3290 (N_3290,N_2483,N_2256);
nor U3291 (N_3291,N_2515,N_2346);
nor U3292 (N_3292,N_2459,N_2830);
or U3293 (N_3293,N_2844,N_2834);
xor U3294 (N_3294,N_2687,N_2388);
nor U3295 (N_3295,N_2396,N_2698);
or U3296 (N_3296,N_2672,N_2212);
xnor U3297 (N_3297,N_2154,N_2494);
xnor U3298 (N_3298,N_2005,N_2307);
nand U3299 (N_3299,N_2551,N_2771);
or U3300 (N_3300,N_2880,N_2539);
xnor U3301 (N_3301,N_2439,N_2748);
nor U3302 (N_3302,N_2376,N_2064);
or U3303 (N_3303,N_2336,N_2033);
or U3304 (N_3304,N_2851,N_2250);
and U3305 (N_3305,N_2766,N_2897);
nand U3306 (N_3306,N_2047,N_2542);
and U3307 (N_3307,N_2549,N_2333);
and U3308 (N_3308,N_2092,N_2145);
nand U3309 (N_3309,N_2750,N_2951);
and U3310 (N_3310,N_2069,N_2990);
or U3311 (N_3311,N_2175,N_2538);
nand U3312 (N_3312,N_2214,N_2248);
nor U3313 (N_3313,N_2014,N_2602);
and U3314 (N_3314,N_2076,N_2013);
or U3315 (N_3315,N_2972,N_2304);
and U3316 (N_3316,N_2475,N_2046);
and U3317 (N_3317,N_2734,N_2031);
nor U3318 (N_3318,N_2314,N_2399);
nor U3319 (N_3319,N_2141,N_2675);
nor U3320 (N_3320,N_2357,N_2071);
xor U3321 (N_3321,N_2078,N_2302);
nand U3322 (N_3322,N_2398,N_2591);
and U3323 (N_3323,N_2342,N_2206);
xnor U3324 (N_3324,N_2810,N_2102);
nor U3325 (N_3325,N_2658,N_2120);
nor U3326 (N_3326,N_2246,N_2105);
nor U3327 (N_3327,N_2003,N_2391);
nor U3328 (N_3328,N_2197,N_2931);
xnor U3329 (N_3329,N_2939,N_2767);
xnor U3330 (N_3330,N_2937,N_2085);
nand U3331 (N_3331,N_2712,N_2298);
nand U3332 (N_3332,N_2707,N_2907);
and U3333 (N_3333,N_2924,N_2424);
nand U3334 (N_3334,N_2992,N_2317);
and U3335 (N_3335,N_2845,N_2779);
nor U3336 (N_3336,N_2794,N_2288);
and U3337 (N_3337,N_2858,N_2009);
and U3338 (N_3338,N_2079,N_2882);
and U3339 (N_3339,N_2789,N_2991);
and U3340 (N_3340,N_2527,N_2294);
nor U3341 (N_3341,N_2866,N_2921);
and U3342 (N_3342,N_2519,N_2534);
nand U3343 (N_3343,N_2431,N_2579);
nor U3344 (N_3344,N_2183,N_2888);
xnor U3345 (N_3345,N_2633,N_2729);
nand U3346 (N_3346,N_2043,N_2998);
nor U3347 (N_3347,N_2617,N_2223);
or U3348 (N_3348,N_2701,N_2583);
xnor U3349 (N_3349,N_2192,N_2996);
nor U3350 (N_3350,N_2671,N_2813);
nor U3351 (N_3351,N_2509,N_2876);
and U3352 (N_3352,N_2015,N_2600);
xnor U3353 (N_3353,N_2491,N_2913);
or U3354 (N_3354,N_2241,N_2282);
nor U3355 (N_3355,N_2091,N_2644);
xor U3356 (N_3356,N_2518,N_2397);
xor U3357 (N_3357,N_2176,N_2165);
or U3358 (N_3358,N_2123,N_2285);
xnor U3359 (N_3359,N_2442,N_2166);
nor U3360 (N_3360,N_2379,N_2902);
or U3361 (N_3361,N_2221,N_2835);
nand U3362 (N_3362,N_2484,N_2215);
and U3363 (N_3363,N_2039,N_2652);
nand U3364 (N_3364,N_2219,N_2422);
or U3365 (N_3365,N_2782,N_2669);
nand U3366 (N_3366,N_2381,N_2385);
xor U3367 (N_3367,N_2564,N_2983);
nand U3368 (N_3368,N_2443,N_2763);
nor U3369 (N_3369,N_2058,N_2063);
xnor U3370 (N_3370,N_2839,N_2607);
nor U3371 (N_3371,N_2673,N_2153);
xnor U3372 (N_3372,N_2692,N_2143);
xor U3373 (N_3373,N_2827,N_2101);
or U3374 (N_3374,N_2649,N_2345);
xor U3375 (N_3375,N_2737,N_2666);
and U3376 (N_3376,N_2274,N_2427);
and U3377 (N_3377,N_2322,N_2344);
and U3378 (N_3378,N_2590,N_2492);
nand U3379 (N_3379,N_2127,N_2472);
nand U3380 (N_3380,N_2832,N_2710);
and U3381 (N_3381,N_2025,N_2305);
and U3382 (N_3382,N_2676,N_2664);
or U3383 (N_3383,N_2098,N_2389);
nand U3384 (N_3384,N_2807,N_2037);
nand U3385 (N_3385,N_2382,N_2485);
xor U3386 (N_3386,N_2578,N_2717);
nand U3387 (N_3387,N_2877,N_2986);
nand U3388 (N_3388,N_2964,N_2318);
nand U3389 (N_3389,N_2700,N_2683);
or U3390 (N_3390,N_2191,N_2022);
xnor U3391 (N_3391,N_2374,N_2177);
xor U3392 (N_3392,N_2418,N_2668);
xnor U3393 (N_3393,N_2021,N_2621);
or U3394 (N_3394,N_2571,N_2874);
and U3395 (N_3395,N_2647,N_2620);
or U3396 (N_3396,N_2048,N_2051);
or U3397 (N_3397,N_2885,N_2547);
or U3398 (N_3398,N_2636,N_2090);
nor U3399 (N_3399,N_2510,N_2134);
nand U3400 (N_3400,N_2213,N_2281);
and U3401 (N_3401,N_2905,N_2087);
xor U3402 (N_3402,N_2159,N_2218);
and U3403 (N_3403,N_2615,N_2878);
nor U3404 (N_3404,N_2169,N_2507);
nand U3405 (N_3405,N_2819,N_2204);
nor U3406 (N_3406,N_2470,N_2872);
xnor U3407 (N_3407,N_2477,N_2616);
xor U3408 (N_3408,N_2711,N_2868);
and U3409 (N_3409,N_2403,N_2815);
nand U3410 (N_3410,N_2148,N_2566);
nor U3411 (N_3411,N_2693,N_2629);
nand U3412 (N_3412,N_2351,N_2055);
nand U3413 (N_3413,N_2283,N_2993);
and U3414 (N_3414,N_2630,N_2060);
or U3415 (N_3415,N_2861,N_2555);
nand U3416 (N_3416,N_2575,N_2432);
xor U3417 (N_3417,N_2560,N_2181);
and U3418 (N_3418,N_2164,N_2474);
or U3419 (N_3419,N_2419,N_2184);
and U3420 (N_3420,N_2561,N_2765);
nand U3421 (N_3421,N_2631,N_2361);
nand U3422 (N_3422,N_2354,N_2569);
nand U3423 (N_3423,N_2393,N_2762);
nand U3424 (N_3424,N_2887,N_2161);
nor U3425 (N_3425,N_2867,N_2428);
nand U3426 (N_3426,N_2588,N_2198);
and U3427 (N_3427,N_2168,N_2228);
nor U3428 (N_3428,N_2320,N_2883);
nand U3429 (N_3429,N_2276,N_2774);
nand U3430 (N_3430,N_2309,N_2299);
and U3431 (N_3431,N_2947,N_2032);
or U3432 (N_3432,N_2232,N_2132);
and U3433 (N_3433,N_2163,N_2864);
xnor U3434 (N_3434,N_2395,N_2297);
nand U3435 (N_3435,N_2599,N_2961);
xor U3436 (N_3436,N_2981,N_2312);
and U3437 (N_3437,N_2155,N_2272);
or U3438 (N_3438,N_2364,N_2158);
and U3439 (N_3439,N_2940,N_2520);
xnor U3440 (N_3440,N_2279,N_2026);
xor U3441 (N_3441,N_2375,N_2179);
xnor U3442 (N_3442,N_2643,N_2479);
nand U3443 (N_3443,N_2942,N_2074);
nor U3444 (N_3444,N_2738,N_2761);
and U3445 (N_3445,N_2266,N_2437);
nor U3446 (N_3446,N_2072,N_2978);
nor U3447 (N_3447,N_2125,N_2010);
nor U3448 (N_3448,N_2988,N_2231);
or U3449 (N_3449,N_2142,N_2019);
xor U3450 (N_3450,N_2016,N_2481);
xnor U3451 (N_3451,N_2800,N_2405);
and U3452 (N_3452,N_2788,N_2150);
nand U3453 (N_3453,N_2028,N_2006);
or U3454 (N_3454,N_2589,N_2111);
and U3455 (N_3455,N_2543,N_2170);
and U3456 (N_3456,N_2140,N_2088);
and U3457 (N_3457,N_2746,N_2487);
and U3458 (N_3458,N_2007,N_2744);
xnor U3459 (N_3459,N_2099,N_2684);
and U3460 (N_3460,N_2758,N_2768);
xor U3461 (N_3461,N_2315,N_2095);
and U3462 (N_3462,N_2358,N_2467);
or U3463 (N_3463,N_2478,N_2196);
and U3464 (N_3464,N_2359,N_2967);
nand U3465 (N_3465,N_2580,N_2325);
nor U3466 (N_3466,N_2533,N_2012);
xor U3467 (N_3467,N_2655,N_2743);
and U3468 (N_3468,N_2017,N_2803);
nand U3469 (N_3469,N_2438,N_2471);
nand U3470 (N_3470,N_2594,N_2073);
or U3471 (N_3471,N_2809,N_2793);
nor U3472 (N_3472,N_2541,N_2922);
xnor U3473 (N_3473,N_2411,N_2505);
nand U3474 (N_3474,N_2934,N_2537);
and U3475 (N_3475,N_2186,N_2188);
nand U3476 (N_3476,N_2689,N_2597);
nand U3477 (N_3477,N_2890,N_2473);
and U3478 (N_3478,N_2903,N_2648);
or U3479 (N_3479,N_2956,N_2909);
nor U3480 (N_3480,N_2869,N_2586);
xnor U3481 (N_3481,N_2828,N_2795);
or U3482 (N_3482,N_2264,N_2040);
or U3483 (N_3483,N_2369,N_2444);
or U3484 (N_3484,N_2755,N_2261);
xnor U3485 (N_3485,N_2966,N_2870);
nand U3486 (N_3486,N_2894,N_2480);
xor U3487 (N_3487,N_2841,N_2930);
or U3488 (N_3488,N_2151,N_2565);
or U3489 (N_3489,N_2103,N_2567);
nor U3490 (N_3490,N_2626,N_2773);
xor U3491 (N_3491,N_2645,N_2926);
nand U3492 (N_3492,N_2194,N_2860);
nand U3493 (N_3493,N_2195,N_2559);
nor U3494 (N_3494,N_2508,N_2486);
or U3495 (N_3495,N_2401,N_2889);
or U3496 (N_3496,N_2493,N_2460);
xor U3497 (N_3497,N_2289,N_2517);
nand U3498 (N_3498,N_2036,N_2268);
xor U3499 (N_3499,N_2735,N_2137);
and U3500 (N_3500,N_2042,N_2777);
and U3501 (N_3501,N_2983,N_2457);
and U3502 (N_3502,N_2971,N_2286);
or U3503 (N_3503,N_2070,N_2660);
xor U3504 (N_3504,N_2793,N_2796);
xor U3505 (N_3505,N_2672,N_2137);
xor U3506 (N_3506,N_2438,N_2130);
and U3507 (N_3507,N_2439,N_2410);
and U3508 (N_3508,N_2949,N_2137);
nand U3509 (N_3509,N_2546,N_2039);
xnor U3510 (N_3510,N_2295,N_2523);
nand U3511 (N_3511,N_2106,N_2365);
or U3512 (N_3512,N_2676,N_2802);
xor U3513 (N_3513,N_2928,N_2651);
xnor U3514 (N_3514,N_2082,N_2244);
xnor U3515 (N_3515,N_2542,N_2501);
xnor U3516 (N_3516,N_2593,N_2398);
or U3517 (N_3517,N_2065,N_2887);
or U3518 (N_3518,N_2367,N_2342);
and U3519 (N_3519,N_2955,N_2398);
xor U3520 (N_3520,N_2434,N_2303);
xnor U3521 (N_3521,N_2882,N_2332);
xor U3522 (N_3522,N_2574,N_2455);
xnor U3523 (N_3523,N_2906,N_2307);
nand U3524 (N_3524,N_2218,N_2375);
or U3525 (N_3525,N_2019,N_2366);
xnor U3526 (N_3526,N_2874,N_2679);
or U3527 (N_3527,N_2995,N_2385);
nand U3528 (N_3528,N_2391,N_2515);
nand U3529 (N_3529,N_2731,N_2182);
xor U3530 (N_3530,N_2662,N_2559);
nor U3531 (N_3531,N_2324,N_2855);
xnor U3532 (N_3532,N_2675,N_2435);
xor U3533 (N_3533,N_2322,N_2069);
nand U3534 (N_3534,N_2623,N_2581);
or U3535 (N_3535,N_2016,N_2318);
and U3536 (N_3536,N_2116,N_2916);
and U3537 (N_3537,N_2421,N_2005);
or U3538 (N_3538,N_2999,N_2729);
and U3539 (N_3539,N_2555,N_2784);
nand U3540 (N_3540,N_2697,N_2917);
nor U3541 (N_3541,N_2189,N_2132);
or U3542 (N_3542,N_2623,N_2150);
and U3543 (N_3543,N_2475,N_2705);
or U3544 (N_3544,N_2569,N_2583);
or U3545 (N_3545,N_2541,N_2182);
or U3546 (N_3546,N_2688,N_2522);
or U3547 (N_3547,N_2675,N_2626);
or U3548 (N_3548,N_2057,N_2312);
or U3549 (N_3549,N_2347,N_2157);
nor U3550 (N_3550,N_2394,N_2959);
or U3551 (N_3551,N_2332,N_2948);
nor U3552 (N_3552,N_2333,N_2778);
and U3553 (N_3553,N_2259,N_2372);
or U3554 (N_3554,N_2813,N_2936);
and U3555 (N_3555,N_2252,N_2698);
nor U3556 (N_3556,N_2608,N_2423);
xor U3557 (N_3557,N_2863,N_2048);
or U3558 (N_3558,N_2071,N_2351);
xnor U3559 (N_3559,N_2468,N_2173);
nand U3560 (N_3560,N_2999,N_2593);
and U3561 (N_3561,N_2812,N_2209);
and U3562 (N_3562,N_2178,N_2431);
nor U3563 (N_3563,N_2570,N_2552);
nor U3564 (N_3564,N_2074,N_2311);
nand U3565 (N_3565,N_2500,N_2549);
or U3566 (N_3566,N_2630,N_2681);
or U3567 (N_3567,N_2204,N_2056);
nor U3568 (N_3568,N_2195,N_2132);
nor U3569 (N_3569,N_2530,N_2098);
xor U3570 (N_3570,N_2887,N_2690);
xor U3571 (N_3571,N_2784,N_2988);
xnor U3572 (N_3572,N_2133,N_2932);
or U3573 (N_3573,N_2676,N_2377);
and U3574 (N_3574,N_2855,N_2883);
nor U3575 (N_3575,N_2736,N_2665);
nor U3576 (N_3576,N_2916,N_2064);
nor U3577 (N_3577,N_2097,N_2881);
xor U3578 (N_3578,N_2658,N_2699);
nor U3579 (N_3579,N_2643,N_2587);
nor U3580 (N_3580,N_2811,N_2793);
and U3581 (N_3581,N_2168,N_2802);
and U3582 (N_3582,N_2104,N_2597);
nand U3583 (N_3583,N_2747,N_2887);
and U3584 (N_3584,N_2053,N_2421);
nor U3585 (N_3585,N_2787,N_2781);
and U3586 (N_3586,N_2958,N_2188);
nand U3587 (N_3587,N_2568,N_2561);
nor U3588 (N_3588,N_2879,N_2379);
or U3589 (N_3589,N_2697,N_2469);
and U3590 (N_3590,N_2851,N_2971);
and U3591 (N_3591,N_2708,N_2711);
and U3592 (N_3592,N_2520,N_2244);
nand U3593 (N_3593,N_2438,N_2150);
or U3594 (N_3594,N_2583,N_2540);
or U3595 (N_3595,N_2389,N_2210);
and U3596 (N_3596,N_2099,N_2288);
nor U3597 (N_3597,N_2246,N_2264);
nand U3598 (N_3598,N_2270,N_2457);
or U3599 (N_3599,N_2572,N_2219);
nor U3600 (N_3600,N_2663,N_2157);
nand U3601 (N_3601,N_2912,N_2149);
nor U3602 (N_3602,N_2343,N_2506);
nor U3603 (N_3603,N_2690,N_2649);
xnor U3604 (N_3604,N_2247,N_2953);
or U3605 (N_3605,N_2403,N_2792);
or U3606 (N_3606,N_2875,N_2247);
nand U3607 (N_3607,N_2779,N_2264);
and U3608 (N_3608,N_2647,N_2670);
nor U3609 (N_3609,N_2060,N_2225);
and U3610 (N_3610,N_2985,N_2262);
xor U3611 (N_3611,N_2761,N_2805);
nand U3612 (N_3612,N_2878,N_2584);
nor U3613 (N_3613,N_2758,N_2425);
nor U3614 (N_3614,N_2469,N_2000);
nor U3615 (N_3615,N_2248,N_2511);
nand U3616 (N_3616,N_2038,N_2148);
and U3617 (N_3617,N_2233,N_2120);
xnor U3618 (N_3618,N_2844,N_2997);
or U3619 (N_3619,N_2613,N_2171);
and U3620 (N_3620,N_2194,N_2043);
and U3621 (N_3621,N_2994,N_2603);
nor U3622 (N_3622,N_2500,N_2801);
nand U3623 (N_3623,N_2167,N_2721);
and U3624 (N_3624,N_2464,N_2825);
xor U3625 (N_3625,N_2320,N_2459);
xnor U3626 (N_3626,N_2452,N_2295);
nor U3627 (N_3627,N_2205,N_2504);
or U3628 (N_3628,N_2113,N_2510);
and U3629 (N_3629,N_2511,N_2863);
or U3630 (N_3630,N_2432,N_2999);
or U3631 (N_3631,N_2326,N_2523);
and U3632 (N_3632,N_2659,N_2167);
and U3633 (N_3633,N_2785,N_2681);
or U3634 (N_3634,N_2696,N_2205);
xnor U3635 (N_3635,N_2988,N_2442);
xnor U3636 (N_3636,N_2940,N_2727);
or U3637 (N_3637,N_2925,N_2102);
xor U3638 (N_3638,N_2372,N_2633);
or U3639 (N_3639,N_2044,N_2955);
nand U3640 (N_3640,N_2884,N_2808);
xnor U3641 (N_3641,N_2600,N_2895);
nor U3642 (N_3642,N_2984,N_2121);
nand U3643 (N_3643,N_2140,N_2523);
nor U3644 (N_3644,N_2937,N_2422);
xor U3645 (N_3645,N_2880,N_2532);
or U3646 (N_3646,N_2450,N_2726);
nor U3647 (N_3647,N_2005,N_2196);
nor U3648 (N_3648,N_2698,N_2637);
nand U3649 (N_3649,N_2672,N_2742);
nor U3650 (N_3650,N_2422,N_2453);
xor U3651 (N_3651,N_2131,N_2867);
nand U3652 (N_3652,N_2389,N_2596);
nor U3653 (N_3653,N_2151,N_2601);
or U3654 (N_3654,N_2504,N_2137);
and U3655 (N_3655,N_2210,N_2373);
xnor U3656 (N_3656,N_2405,N_2890);
nand U3657 (N_3657,N_2073,N_2775);
or U3658 (N_3658,N_2368,N_2384);
xor U3659 (N_3659,N_2469,N_2889);
nand U3660 (N_3660,N_2391,N_2920);
or U3661 (N_3661,N_2688,N_2146);
nor U3662 (N_3662,N_2856,N_2521);
nand U3663 (N_3663,N_2063,N_2325);
nor U3664 (N_3664,N_2286,N_2362);
nand U3665 (N_3665,N_2981,N_2660);
and U3666 (N_3666,N_2599,N_2889);
nor U3667 (N_3667,N_2226,N_2153);
and U3668 (N_3668,N_2383,N_2537);
and U3669 (N_3669,N_2173,N_2747);
nor U3670 (N_3670,N_2237,N_2502);
or U3671 (N_3671,N_2644,N_2869);
and U3672 (N_3672,N_2825,N_2292);
and U3673 (N_3673,N_2177,N_2826);
nand U3674 (N_3674,N_2919,N_2626);
nand U3675 (N_3675,N_2552,N_2294);
and U3676 (N_3676,N_2879,N_2961);
xnor U3677 (N_3677,N_2908,N_2022);
or U3678 (N_3678,N_2389,N_2577);
nor U3679 (N_3679,N_2312,N_2433);
and U3680 (N_3680,N_2419,N_2919);
nor U3681 (N_3681,N_2453,N_2980);
and U3682 (N_3682,N_2832,N_2558);
nor U3683 (N_3683,N_2420,N_2689);
and U3684 (N_3684,N_2985,N_2990);
or U3685 (N_3685,N_2401,N_2706);
xnor U3686 (N_3686,N_2939,N_2236);
xnor U3687 (N_3687,N_2799,N_2327);
nand U3688 (N_3688,N_2617,N_2095);
nor U3689 (N_3689,N_2401,N_2280);
or U3690 (N_3690,N_2861,N_2674);
nand U3691 (N_3691,N_2297,N_2532);
and U3692 (N_3692,N_2309,N_2945);
xnor U3693 (N_3693,N_2063,N_2520);
and U3694 (N_3694,N_2436,N_2829);
nor U3695 (N_3695,N_2173,N_2461);
xor U3696 (N_3696,N_2117,N_2248);
nor U3697 (N_3697,N_2822,N_2189);
or U3698 (N_3698,N_2015,N_2247);
xor U3699 (N_3699,N_2505,N_2510);
or U3700 (N_3700,N_2801,N_2813);
nand U3701 (N_3701,N_2636,N_2264);
or U3702 (N_3702,N_2867,N_2096);
or U3703 (N_3703,N_2758,N_2193);
xor U3704 (N_3704,N_2846,N_2462);
and U3705 (N_3705,N_2195,N_2330);
nand U3706 (N_3706,N_2189,N_2473);
xor U3707 (N_3707,N_2927,N_2712);
nor U3708 (N_3708,N_2340,N_2974);
and U3709 (N_3709,N_2982,N_2384);
and U3710 (N_3710,N_2669,N_2699);
and U3711 (N_3711,N_2969,N_2788);
xor U3712 (N_3712,N_2798,N_2144);
xor U3713 (N_3713,N_2350,N_2427);
and U3714 (N_3714,N_2810,N_2403);
nor U3715 (N_3715,N_2010,N_2765);
and U3716 (N_3716,N_2993,N_2773);
nor U3717 (N_3717,N_2826,N_2870);
and U3718 (N_3718,N_2926,N_2495);
nor U3719 (N_3719,N_2212,N_2662);
nor U3720 (N_3720,N_2836,N_2905);
or U3721 (N_3721,N_2570,N_2109);
or U3722 (N_3722,N_2256,N_2187);
nand U3723 (N_3723,N_2862,N_2644);
or U3724 (N_3724,N_2215,N_2252);
and U3725 (N_3725,N_2567,N_2444);
nor U3726 (N_3726,N_2036,N_2163);
nor U3727 (N_3727,N_2893,N_2774);
nand U3728 (N_3728,N_2722,N_2487);
or U3729 (N_3729,N_2668,N_2657);
xor U3730 (N_3730,N_2148,N_2754);
and U3731 (N_3731,N_2416,N_2302);
xor U3732 (N_3732,N_2714,N_2416);
xnor U3733 (N_3733,N_2276,N_2813);
or U3734 (N_3734,N_2768,N_2245);
nor U3735 (N_3735,N_2549,N_2898);
and U3736 (N_3736,N_2680,N_2891);
nand U3737 (N_3737,N_2161,N_2281);
xor U3738 (N_3738,N_2130,N_2131);
or U3739 (N_3739,N_2492,N_2131);
xnor U3740 (N_3740,N_2695,N_2346);
xor U3741 (N_3741,N_2998,N_2036);
nand U3742 (N_3742,N_2795,N_2935);
or U3743 (N_3743,N_2275,N_2166);
and U3744 (N_3744,N_2588,N_2743);
nor U3745 (N_3745,N_2391,N_2326);
or U3746 (N_3746,N_2851,N_2833);
or U3747 (N_3747,N_2517,N_2988);
and U3748 (N_3748,N_2363,N_2408);
nor U3749 (N_3749,N_2481,N_2709);
and U3750 (N_3750,N_2181,N_2328);
and U3751 (N_3751,N_2138,N_2596);
nor U3752 (N_3752,N_2604,N_2187);
or U3753 (N_3753,N_2934,N_2441);
nor U3754 (N_3754,N_2122,N_2860);
and U3755 (N_3755,N_2361,N_2758);
nor U3756 (N_3756,N_2786,N_2265);
xor U3757 (N_3757,N_2834,N_2867);
nand U3758 (N_3758,N_2492,N_2672);
or U3759 (N_3759,N_2303,N_2398);
or U3760 (N_3760,N_2887,N_2431);
nor U3761 (N_3761,N_2868,N_2549);
nor U3762 (N_3762,N_2356,N_2809);
nor U3763 (N_3763,N_2283,N_2219);
xnor U3764 (N_3764,N_2598,N_2575);
xnor U3765 (N_3765,N_2430,N_2928);
and U3766 (N_3766,N_2425,N_2561);
and U3767 (N_3767,N_2908,N_2220);
xnor U3768 (N_3768,N_2264,N_2194);
nand U3769 (N_3769,N_2056,N_2633);
and U3770 (N_3770,N_2764,N_2014);
or U3771 (N_3771,N_2459,N_2979);
nor U3772 (N_3772,N_2606,N_2516);
nand U3773 (N_3773,N_2754,N_2854);
or U3774 (N_3774,N_2343,N_2256);
or U3775 (N_3775,N_2545,N_2737);
or U3776 (N_3776,N_2704,N_2779);
or U3777 (N_3777,N_2723,N_2991);
or U3778 (N_3778,N_2781,N_2280);
or U3779 (N_3779,N_2012,N_2460);
xor U3780 (N_3780,N_2720,N_2283);
nor U3781 (N_3781,N_2464,N_2405);
xor U3782 (N_3782,N_2385,N_2044);
nand U3783 (N_3783,N_2549,N_2982);
and U3784 (N_3784,N_2374,N_2459);
nor U3785 (N_3785,N_2228,N_2922);
nor U3786 (N_3786,N_2901,N_2953);
and U3787 (N_3787,N_2669,N_2140);
or U3788 (N_3788,N_2396,N_2428);
and U3789 (N_3789,N_2006,N_2470);
nand U3790 (N_3790,N_2685,N_2698);
xnor U3791 (N_3791,N_2593,N_2881);
xor U3792 (N_3792,N_2803,N_2503);
or U3793 (N_3793,N_2746,N_2730);
xor U3794 (N_3794,N_2541,N_2328);
and U3795 (N_3795,N_2147,N_2596);
nand U3796 (N_3796,N_2675,N_2027);
or U3797 (N_3797,N_2168,N_2090);
nor U3798 (N_3798,N_2230,N_2887);
xor U3799 (N_3799,N_2593,N_2714);
and U3800 (N_3800,N_2374,N_2531);
nand U3801 (N_3801,N_2459,N_2146);
nor U3802 (N_3802,N_2633,N_2765);
xnor U3803 (N_3803,N_2775,N_2729);
or U3804 (N_3804,N_2429,N_2452);
and U3805 (N_3805,N_2316,N_2386);
xor U3806 (N_3806,N_2241,N_2030);
nand U3807 (N_3807,N_2408,N_2465);
nor U3808 (N_3808,N_2882,N_2235);
xor U3809 (N_3809,N_2689,N_2184);
or U3810 (N_3810,N_2899,N_2357);
and U3811 (N_3811,N_2334,N_2369);
and U3812 (N_3812,N_2814,N_2524);
xor U3813 (N_3813,N_2480,N_2374);
or U3814 (N_3814,N_2048,N_2907);
or U3815 (N_3815,N_2254,N_2618);
nand U3816 (N_3816,N_2460,N_2530);
and U3817 (N_3817,N_2169,N_2035);
nor U3818 (N_3818,N_2564,N_2451);
nor U3819 (N_3819,N_2394,N_2724);
xnor U3820 (N_3820,N_2050,N_2480);
xor U3821 (N_3821,N_2659,N_2430);
nand U3822 (N_3822,N_2910,N_2267);
and U3823 (N_3823,N_2973,N_2068);
nand U3824 (N_3824,N_2136,N_2400);
xor U3825 (N_3825,N_2574,N_2418);
and U3826 (N_3826,N_2746,N_2669);
xor U3827 (N_3827,N_2320,N_2058);
xnor U3828 (N_3828,N_2666,N_2637);
or U3829 (N_3829,N_2740,N_2638);
nand U3830 (N_3830,N_2976,N_2085);
xnor U3831 (N_3831,N_2513,N_2146);
and U3832 (N_3832,N_2195,N_2648);
and U3833 (N_3833,N_2703,N_2881);
nand U3834 (N_3834,N_2272,N_2727);
xor U3835 (N_3835,N_2192,N_2390);
nand U3836 (N_3836,N_2416,N_2293);
or U3837 (N_3837,N_2822,N_2306);
and U3838 (N_3838,N_2483,N_2781);
and U3839 (N_3839,N_2597,N_2857);
nand U3840 (N_3840,N_2360,N_2874);
nor U3841 (N_3841,N_2171,N_2576);
or U3842 (N_3842,N_2725,N_2845);
and U3843 (N_3843,N_2262,N_2033);
xor U3844 (N_3844,N_2877,N_2856);
and U3845 (N_3845,N_2467,N_2959);
and U3846 (N_3846,N_2866,N_2984);
nor U3847 (N_3847,N_2226,N_2107);
nand U3848 (N_3848,N_2448,N_2466);
or U3849 (N_3849,N_2689,N_2679);
or U3850 (N_3850,N_2624,N_2469);
nand U3851 (N_3851,N_2882,N_2087);
xor U3852 (N_3852,N_2261,N_2057);
nand U3853 (N_3853,N_2017,N_2383);
nand U3854 (N_3854,N_2418,N_2834);
or U3855 (N_3855,N_2566,N_2012);
or U3856 (N_3856,N_2154,N_2937);
nand U3857 (N_3857,N_2306,N_2680);
and U3858 (N_3858,N_2640,N_2788);
xnor U3859 (N_3859,N_2122,N_2770);
nor U3860 (N_3860,N_2165,N_2952);
and U3861 (N_3861,N_2030,N_2777);
nor U3862 (N_3862,N_2136,N_2309);
and U3863 (N_3863,N_2186,N_2630);
and U3864 (N_3864,N_2183,N_2964);
xnor U3865 (N_3865,N_2732,N_2545);
nor U3866 (N_3866,N_2881,N_2740);
xnor U3867 (N_3867,N_2335,N_2553);
nand U3868 (N_3868,N_2008,N_2769);
and U3869 (N_3869,N_2515,N_2171);
nand U3870 (N_3870,N_2555,N_2810);
xnor U3871 (N_3871,N_2847,N_2437);
or U3872 (N_3872,N_2548,N_2992);
and U3873 (N_3873,N_2071,N_2750);
and U3874 (N_3874,N_2678,N_2739);
xnor U3875 (N_3875,N_2821,N_2814);
or U3876 (N_3876,N_2809,N_2170);
nand U3877 (N_3877,N_2414,N_2074);
xor U3878 (N_3878,N_2160,N_2520);
xnor U3879 (N_3879,N_2028,N_2564);
and U3880 (N_3880,N_2396,N_2132);
nand U3881 (N_3881,N_2139,N_2337);
or U3882 (N_3882,N_2488,N_2921);
and U3883 (N_3883,N_2666,N_2840);
xnor U3884 (N_3884,N_2621,N_2904);
or U3885 (N_3885,N_2006,N_2022);
xor U3886 (N_3886,N_2959,N_2430);
or U3887 (N_3887,N_2947,N_2864);
xor U3888 (N_3888,N_2956,N_2722);
nand U3889 (N_3889,N_2305,N_2060);
or U3890 (N_3890,N_2840,N_2102);
or U3891 (N_3891,N_2100,N_2721);
xnor U3892 (N_3892,N_2912,N_2202);
nor U3893 (N_3893,N_2848,N_2051);
xnor U3894 (N_3894,N_2730,N_2064);
or U3895 (N_3895,N_2631,N_2492);
xor U3896 (N_3896,N_2352,N_2254);
xnor U3897 (N_3897,N_2058,N_2274);
xor U3898 (N_3898,N_2846,N_2176);
nor U3899 (N_3899,N_2906,N_2702);
nand U3900 (N_3900,N_2835,N_2070);
xor U3901 (N_3901,N_2676,N_2090);
nand U3902 (N_3902,N_2404,N_2755);
and U3903 (N_3903,N_2921,N_2990);
nand U3904 (N_3904,N_2341,N_2103);
nand U3905 (N_3905,N_2928,N_2862);
or U3906 (N_3906,N_2205,N_2220);
xor U3907 (N_3907,N_2163,N_2266);
nand U3908 (N_3908,N_2214,N_2488);
and U3909 (N_3909,N_2101,N_2176);
nand U3910 (N_3910,N_2324,N_2420);
or U3911 (N_3911,N_2314,N_2915);
and U3912 (N_3912,N_2020,N_2515);
and U3913 (N_3913,N_2044,N_2655);
or U3914 (N_3914,N_2894,N_2672);
nand U3915 (N_3915,N_2779,N_2618);
or U3916 (N_3916,N_2341,N_2142);
nor U3917 (N_3917,N_2407,N_2050);
nand U3918 (N_3918,N_2322,N_2973);
or U3919 (N_3919,N_2542,N_2942);
nor U3920 (N_3920,N_2880,N_2110);
nor U3921 (N_3921,N_2362,N_2560);
and U3922 (N_3922,N_2442,N_2375);
or U3923 (N_3923,N_2932,N_2105);
xor U3924 (N_3924,N_2002,N_2512);
xnor U3925 (N_3925,N_2797,N_2165);
or U3926 (N_3926,N_2302,N_2289);
nand U3927 (N_3927,N_2388,N_2435);
nor U3928 (N_3928,N_2332,N_2264);
or U3929 (N_3929,N_2824,N_2894);
xnor U3930 (N_3930,N_2454,N_2676);
nand U3931 (N_3931,N_2291,N_2790);
and U3932 (N_3932,N_2037,N_2689);
and U3933 (N_3933,N_2228,N_2589);
or U3934 (N_3934,N_2827,N_2456);
and U3935 (N_3935,N_2151,N_2654);
xor U3936 (N_3936,N_2899,N_2891);
nand U3937 (N_3937,N_2819,N_2136);
nand U3938 (N_3938,N_2660,N_2302);
and U3939 (N_3939,N_2519,N_2856);
nand U3940 (N_3940,N_2735,N_2783);
nor U3941 (N_3941,N_2933,N_2109);
nand U3942 (N_3942,N_2130,N_2268);
xor U3943 (N_3943,N_2496,N_2490);
nand U3944 (N_3944,N_2674,N_2392);
nor U3945 (N_3945,N_2791,N_2456);
xor U3946 (N_3946,N_2491,N_2568);
nand U3947 (N_3947,N_2684,N_2521);
nand U3948 (N_3948,N_2549,N_2255);
nand U3949 (N_3949,N_2519,N_2506);
or U3950 (N_3950,N_2902,N_2782);
and U3951 (N_3951,N_2916,N_2532);
and U3952 (N_3952,N_2229,N_2764);
and U3953 (N_3953,N_2937,N_2320);
nand U3954 (N_3954,N_2043,N_2567);
or U3955 (N_3955,N_2971,N_2811);
nand U3956 (N_3956,N_2868,N_2031);
or U3957 (N_3957,N_2404,N_2563);
nand U3958 (N_3958,N_2194,N_2190);
and U3959 (N_3959,N_2768,N_2161);
or U3960 (N_3960,N_2204,N_2467);
nand U3961 (N_3961,N_2365,N_2526);
nor U3962 (N_3962,N_2554,N_2933);
or U3963 (N_3963,N_2816,N_2539);
nor U3964 (N_3964,N_2652,N_2617);
nor U3965 (N_3965,N_2426,N_2566);
nor U3966 (N_3966,N_2868,N_2059);
xnor U3967 (N_3967,N_2638,N_2245);
xnor U3968 (N_3968,N_2829,N_2876);
or U3969 (N_3969,N_2519,N_2331);
nor U3970 (N_3970,N_2594,N_2534);
xor U3971 (N_3971,N_2612,N_2239);
or U3972 (N_3972,N_2360,N_2548);
nor U3973 (N_3973,N_2229,N_2712);
and U3974 (N_3974,N_2291,N_2073);
nor U3975 (N_3975,N_2659,N_2173);
nand U3976 (N_3976,N_2698,N_2559);
or U3977 (N_3977,N_2450,N_2176);
nand U3978 (N_3978,N_2396,N_2266);
nand U3979 (N_3979,N_2734,N_2199);
nor U3980 (N_3980,N_2394,N_2630);
xor U3981 (N_3981,N_2881,N_2468);
or U3982 (N_3982,N_2710,N_2507);
or U3983 (N_3983,N_2620,N_2966);
or U3984 (N_3984,N_2033,N_2635);
nand U3985 (N_3985,N_2130,N_2627);
xor U3986 (N_3986,N_2460,N_2775);
nor U3987 (N_3987,N_2652,N_2386);
xnor U3988 (N_3988,N_2056,N_2787);
xnor U3989 (N_3989,N_2356,N_2641);
nand U3990 (N_3990,N_2999,N_2294);
nand U3991 (N_3991,N_2869,N_2086);
xor U3992 (N_3992,N_2191,N_2441);
nand U3993 (N_3993,N_2696,N_2481);
nor U3994 (N_3994,N_2667,N_2597);
and U3995 (N_3995,N_2243,N_2063);
nand U3996 (N_3996,N_2586,N_2086);
xor U3997 (N_3997,N_2031,N_2233);
nand U3998 (N_3998,N_2735,N_2662);
xnor U3999 (N_3999,N_2143,N_2207);
and U4000 (N_4000,N_3527,N_3808);
or U4001 (N_4001,N_3170,N_3693);
xor U4002 (N_4002,N_3692,N_3861);
nand U4003 (N_4003,N_3632,N_3002);
and U4004 (N_4004,N_3863,N_3975);
nor U4005 (N_4005,N_3958,N_3371);
nand U4006 (N_4006,N_3666,N_3589);
or U4007 (N_4007,N_3049,N_3866);
nor U4008 (N_4008,N_3557,N_3925);
xor U4009 (N_4009,N_3685,N_3740);
and U4010 (N_4010,N_3443,N_3508);
xnor U4011 (N_4011,N_3826,N_3630);
xnor U4012 (N_4012,N_3191,N_3536);
nor U4013 (N_4013,N_3389,N_3003);
nand U4014 (N_4014,N_3552,N_3806);
xor U4015 (N_4015,N_3071,N_3533);
and U4016 (N_4016,N_3553,N_3103);
xor U4017 (N_4017,N_3864,N_3821);
nor U4018 (N_4018,N_3922,N_3151);
or U4019 (N_4019,N_3481,N_3137);
or U4020 (N_4020,N_3383,N_3700);
nand U4021 (N_4021,N_3026,N_3878);
or U4022 (N_4022,N_3231,N_3426);
xnor U4023 (N_4023,N_3627,N_3949);
and U4024 (N_4024,N_3273,N_3939);
or U4025 (N_4025,N_3992,N_3354);
or U4026 (N_4026,N_3794,N_3235);
or U4027 (N_4027,N_3368,N_3653);
nor U4028 (N_4028,N_3737,N_3787);
nor U4029 (N_4029,N_3683,N_3633);
and U4030 (N_4030,N_3118,N_3884);
xor U4031 (N_4031,N_3624,N_3255);
xor U4032 (N_4032,N_3807,N_3597);
and U4033 (N_4033,N_3476,N_3460);
or U4034 (N_4034,N_3429,N_3046);
nand U4035 (N_4035,N_3620,N_3375);
nand U4036 (N_4036,N_3233,N_3778);
or U4037 (N_4037,N_3576,N_3648);
xnor U4038 (N_4038,N_3813,N_3898);
and U4039 (N_4039,N_3133,N_3337);
xnor U4040 (N_4040,N_3546,N_3293);
nor U4041 (N_4041,N_3247,N_3523);
or U4042 (N_4042,N_3823,N_3355);
xor U4043 (N_4043,N_3680,N_3607);
and U4044 (N_4044,N_3328,N_3849);
or U4045 (N_4045,N_3098,N_3467);
or U4046 (N_4046,N_3268,N_3917);
and U4047 (N_4047,N_3444,N_3580);
nand U4048 (N_4048,N_3838,N_3466);
nand U4049 (N_4049,N_3815,N_3634);
nor U4050 (N_4050,N_3927,N_3441);
or U4051 (N_4051,N_3437,N_3631);
nand U4052 (N_4052,N_3540,N_3637);
and U4053 (N_4053,N_3261,N_3168);
nand U4054 (N_4054,N_3198,N_3165);
nand U4055 (N_4055,N_3645,N_3831);
or U4056 (N_4056,N_3901,N_3773);
or U4057 (N_4057,N_3131,N_3083);
xor U4058 (N_4058,N_3801,N_3294);
and U4059 (N_4059,N_3459,N_3208);
xnor U4060 (N_4060,N_3760,N_3820);
nor U4061 (N_4061,N_3169,N_3753);
nor U4062 (N_4062,N_3875,N_3491);
or U4063 (N_4063,N_3391,N_3257);
xnor U4064 (N_4064,N_3800,N_3453);
nor U4065 (N_4065,N_3916,N_3431);
nor U4066 (N_4066,N_3499,N_3783);
xor U4067 (N_4067,N_3140,N_3872);
xor U4068 (N_4068,N_3993,N_3771);
and U4069 (N_4069,N_3784,N_3111);
nand U4070 (N_4070,N_3068,N_3542);
xor U4071 (N_4071,N_3281,N_3341);
or U4072 (N_4072,N_3613,N_3554);
xnor U4073 (N_4073,N_3979,N_3021);
or U4074 (N_4074,N_3192,N_3636);
nand U4075 (N_4075,N_3754,N_3360);
or U4076 (N_4076,N_3125,N_3709);
or U4077 (N_4077,N_3547,N_3988);
xnor U4078 (N_4078,N_3428,N_3042);
and U4079 (N_4079,N_3007,N_3644);
xor U4080 (N_4080,N_3918,N_3020);
xor U4081 (N_4081,N_3910,N_3019);
or U4082 (N_4082,N_3749,N_3144);
or U4083 (N_4083,N_3171,N_3315);
or U4084 (N_4084,N_3908,N_3104);
nor U4085 (N_4085,N_3238,N_3870);
and U4086 (N_4086,N_3660,N_3674);
or U4087 (N_4087,N_3819,N_3578);
nor U4088 (N_4088,N_3503,N_3586);
and U4089 (N_4089,N_3618,N_3909);
and U4090 (N_4090,N_3659,N_3848);
xor U4091 (N_4091,N_3505,N_3498);
or U4092 (N_4092,N_3719,N_3507);
xnor U4093 (N_4093,N_3654,N_3851);
and U4094 (N_4094,N_3403,N_3983);
nand U4095 (N_4095,N_3926,N_3359);
nand U4096 (N_4096,N_3405,N_3350);
xnor U4097 (N_4097,N_3130,N_3640);
xnor U4098 (N_4098,N_3526,N_3480);
nor U4099 (N_4099,N_3642,N_3722);
or U4100 (N_4100,N_3410,N_3432);
xnor U4101 (N_4101,N_3162,N_3905);
nor U4102 (N_4102,N_3677,N_3469);
or U4103 (N_4103,N_3101,N_3073);
or U4104 (N_4104,N_3197,N_3698);
xnor U4105 (N_4105,N_3253,N_3306);
nand U4106 (N_4106,N_3729,N_3406);
nor U4107 (N_4107,N_3195,N_3183);
nand U4108 (N_4108,N_3221,N_3770);
xnor U4109 (N_4109,N_3063,N_3574);
nor U4110 (N_4110,N_3928,N_3564);
nor U4111 (N_4111,N_3996,N_3040);
xnor U4112 (N_4112,N_3216,N_3070);
and U4113 (N_4113,N_3414,N_3489);
xor U4114 (N_4114,N_3969,N_3639);
or U4115 (N_4115,N_3768,N_3731);
and U4116 (N_4116,N_3114,N_3756);
xor U4117 (N_4117,N_3055,N_3282);
and U4118 (N_4118,N_3423,N_3710);
nand U4119 (N_4119,N_3088,N_3513);
and U4120 (N_4120,N_3832,N_3834);
and U4121 (N_4121,N_3803,N_3960);
nor U4122 (N_4122,N_3248,N_3575);
and U4123 (N_4123,N_3978,N_3177);
and U4124 (N_4124,N_3260,N_3193);
and U4125 (N_4125,N_3920,N_3448);
nand U4126 (N_4126,N_3242,N_3043);
nor U4127 (N_4127,N_3963,N_3959);
xor U4128 (N_4128,N_3881,N_3132);
xor U4129 (N_4129,N_3774,N_3655);
and U4130 (N_4130,N_3516,N_3903);
or U4131 (N_4131,N_3682,N_3712);
nand U4132 (N_4132,N_3464,N_3651);
nor U4133 (N_4133,N_3135,N_3529);
nand U4134 (N_4134,N_3329,N_3146);
nand U4135 (N_4135,N_3027,N_3269);
and U4136 (N_4136,N_3500,N_3089);
nor U4137 (N_4137,N_3924,N_3822);
and U4138 (N_4138,N_3810,N_3343);
nand U4139 (N_4139,N_3038,N_3695);
xor U4140 (N_4140,N_3211,N_3080);
or U4141 (N_4141,N_3887,N_3549);
xor U4142 (N_4142,N_3723,N_3560);
or U4143 (N_4143,N_3950,N_3204);
xnor U4144 (N_4144,N_3150,N_3537);
or U4145 (N_4145,N_3156,N_3424);
or U4146 (N_4146,N_3841,N_3859);
xnor U4147 (N_4147,N_3025,N_3891);
or U4148 (N_4148,N_3658,N_3715);
and U4149 (N_4149,N_3782,N_3041);
nand U4150 (N_4150,N_3474,N_3409);
and U4151 (N_4151,N_3694,N_3187);
xnor U4152 (N_4152,N_3099,N_3128);
nor U4153 (N_4153,N_3495,N_3907);
and U4154 (N_4154,N_3713,N_3596);
and U4155 (N_4155,N_3097,N_3577);
and U4156 (N_4156,N_3867,N_3280);
and U4157 (N_4157,N_3054,N_3289);
or U4158 (N_4158,N_3264,N_3696);
nand U4159 (N_4159,N_3327,N_3532);
nand U4160 (N_4160,N_3301,N_3129);
nand U4161 (N_4161,N_3045,N_3422);
or U4162 (N_4162,N_3805,N_3034);
or U4163 (N_4163,N_3450,N_3015);
and U4164 (N_4164,N_3229,N_3452);
xor U4165 (N_4165,N_3830,N_3739);
nor U4166 (N_4166,N_3716,N_3387);
and U4167 (N_4167,N_3646,N_3797);
nand U4168 (N_4168,N_3276,N_3342);
and U4169 (N_4169,N_3374,N_3930);
xnor U4170 (N_4170,N_3445,N_3203);
nor U4171 (N_4171,N_3766,N_3100);
xor U4172 (N_4172,N_3243,N_3854);
nand U4173 (N_4173,N_3862,N_3181);
nor U4174 (N_4174,N_3944,N_3581);
or U4175 (N_4175,N_3973,N_3417);
or U4176 (N_4176,N_3430,N_3093);
or U4177 (N_4177,N_3724,N_3163);
xor U4178 (N_4178,N_3940,N_3900);
nand U4179 (N_4179,N_3483,N_3955);
nand U4180 (N_4180,N_3291,N_3284);
xnor U4181 (N_4181,N_3600,N_3688);
xor U4182 (N_4182,N_3590,N_3148);
nand U4183 (N_4183,N_3829,N_3323);
nor U4184 (N_4184,N_3643,N_3656);
or U4185 (N_4185,N_3159,N_3117);
xnor U4186 (N_4186,N_3468,N_3962);
or U4187 (N_4187,N_3364,N_3297);
and U4188 (N_4188,N_3401,N_3811);
or U4189 (N_4189,N_3515,N_3224);
nand U4190 (N_4190,N_3012,N_3657);
xnor U4191 (N_4191,N_3732,N_3601);
and U4192 (N_4192,N_3220,N_3947);
and U4193 (N_4193,N_3490,N_3175);
xnor U4194 (N_4194,N_3933,N_3828);
or U4195 (N_4195,N_3090,N_3971);
xor U4196 (N_4196,N_3018,N_3890);
xnor U4197 (N_4197,N_3667,N_3697);
nor U4198 (N_4198,N_3721,N_3869);
nand U4199 (N_4199,N_3091,N_3079);
nor U4200 (N_4200,N_3519,N_3296);
and U4201 (N_4201,N_3957,N_3661);
xor U4202 (N_4202,N_3395,N_3488);
or U4203 (N_4203,N_3571,N_3687);
or U4204 (N_4204,N_3568,N_3384);
nand U4205 (N_4205,N_3970,N_3461);
nor U4206 (N_4206,N_3048,N_3230);
nor U4207 (N_4207,N_3392,N_3030);
or U4208 (N_4208,N_3110,N_3663);
nand U4209 (N_4209,N_3369,N_3702);
and U4210 (N_4210,N_3608,N_3772);
nand U4211 (N_4211,N_3029,N_3011);
nor U4212 (N_4212,N_3116,N_3635);
nand U4213 (N_4213,N_3853,N_3598);
and U4214 (N_4214,N_3477,N_3736);
and U4215 (N_4215,N_3013,N_3792);
and U4216 (N_4216,N_3485,N_3275);
nor U4217 (N_4217,N_3134,N_3565);
nor U4218 (N_4218,N_3455,N_3954);
nor U4219 (N_4219,N_3393,N_3381);
nand U4220 (N_4220,N_3790,N_3934);
xnor U4221 (N_4221,N_3769,N_3705);
xnor U4222 (N_4222,N_3956,N_3338);
or U4223 (N_4223,N_3899,N_3943);
or U4224 (N_4224,N_3398,N_3283);
nor U4225 (N_4225,N_3244,N_3186);
or U4226 (N_4226,N_3595,N_3475);
nand U4227 (N_4227,N_3584,N_3166);
nand U4228 (N_4228,N_3113,N_3427);
or U4229 (N_4229,N_3082,N_3107);
nor U4230 (N_4230,N_3764,N_3497);
or U4231 (N_4231,N_3254,N_3977);
xor U4232 (N_4232,N_3404,N_3741);
nand U4233 (N_4233,N_3031,N_3016);
nor U4234 (N_4234,N_3077,N_3250);
or U4235 (N_4235,N_3326,N_3835);
xor U4236 (N_4236,N_3416,N_3743);
nand U4237 (N_4237,N_3122,N_3921);
and U4238 (N_4238,N_3000,N_3791);
and U4239 (N_4239,N_3272,N_3484);
nand U4240 (N_4240,N_3748,N_3390);
nand U4241 (N_4241,N_3999,N_3747);
xor U4242 (N_4242,N_3793,N_3885);
and U4243 (N_4243,N_3086,N_3278);
xor U4244 (N_4244,N_3435,N_3896);
and U4245 (N_4245,N_3858,N_3312);
xnor U4246 (N_4246,N_3961,N_3524);
nor U4247 (N_4247,N_3436,N_3592);
xor U4248 (N_4248,N_3377,N_3067);
and U4249 (N_4249,N_3616,N_3874);
nor U4250 (N_4250,N_3981,N_3256);
or U4251 (N_4251,N_3447,N_3017);
nor U4252 (N_4252,N_3232,N_3897);
nand U4253 (N_4253,N_3096,N_3370);
nor U4254 (N_4254,N_3691,N_3583);
or U4255 (N_4255,N_3434,N_3157);
nand U4256 (N_4256,N_3202,N_3923);
nand U4257 (N_4257,N_3102,N_3902);
and U4258 (N_4258,N_3671,N_3520);
nor U4259 (N_4259,N_3775,N_3010);
nand U4260 (N_4260,N_3378,N_3109);
nand U4261 (N_4261,N_3836,N_3263);
nand U4262 (N_4262,N_3201,N_3078);
nand U4263 (N_4263,N_3147,N_3185);
nor U4264 (N_4264,N_3946,N_3214);
and U4265 (N_4265,N_3628,N_3473);
or U4266 (N_4266,N_3703,N_3174);
xor U4267 (N_4267,N_3543,N_3788);
nor U4268 (N_4268,N_3415,N_3809);
nand U4269 (N_4269,N_3711,N_3362);
nor U4270 (N_4270,N_3388,N_3911);
and U4271 (N_4271,N_3738,N_3511);
nand U4272 (N_4272,N_3952,N_3143);
xnor U4273 (N_4273,N_3941,N_3176);
or U4274 (N_4274,N_3298,N_3153);
nor U4275 (N_4275,N_3039,N_3539);
nand U4276 (N_4276,N_3249,N_3462);
nand U4277 (N_4277,N_3120,N_3676);
or U4278 (N_4278,N_3295,N_3210);
or U4279 (N_4279,N_3964,N_3471);
and U4280 (N_4280,N_3065,N_3912);
or U4281 (N_4281,N_3223,N_3799);
nand U4282 (N_4282,N_3457,N_3798);
and U4283 (N_4283,N_3309,N_3084);
and U4284 (N_4284,N_3412,N_3846);
and U4285 (N_4285,N_3320,N_3126);
xnor U4286 (N_4286,N_3479,N_3440);
and U4287 (N_4287,N_3419,N_3847);
and U4288 (N_4288,N_3115,N_3382);
and U4289 (N_4289,N_3287,N_3142);
nor U4290 (N_4290,N_3421,N_3812);
xor U4291 (N_4291,N_3744,N_3161);
and U4292 (N_4292,N_3307,N_3056);
and U4293 (N_4293,N_3517,N_3604);
and U4294 (N_4294,N_3108,N_3189);
xor U4295 (N_4295,N_3196,N_3014);
or U4296 (N_4296,N_3347,N_3689);
nor U4297 (N_4297,N_3865,N_3967);
and U4298 (N_4298,N_3718,N_3779);
or U4299 (N_4299,N_3611,N_3514);
or U4300 (N_4300,N_3325,N_3334);
or U4301 (N_4301,N_3913,N_3209);
nand U4302 (N_4302,N_3180,N_3622);
nand U4303 (N_4303,N_3945,N_3681);
nand U4304 (N_4304,N_3619,N_3271);
or U4305 (N_4305,N_3534,N_3585);
nand U4306 (N_4306,N_3501,N_3259);
xnor U4307 (N_4307,N_3037,N_3496);
or U4308 (N_4308,N_3121,N_3302);
or U4309 (N_4309,N_3033,N_3892);
xor U4310 (N_4310,N_3837,N_3332);
nor U4311 (N_4311,N_3840,N_3313);
nor U4312 (N_4312,N_3124,N_3614);
or U4313 (N_4313,N_3331,N_3545);
nor U4314 (N_4314,N_3236,N_3786);
nor U4315 (N_4315,N_3300,N_3504);
xor U4316 (N_4316,N_3879,N_3478);
or U4317 (N_4317,N_3182,N_3953);
xor U4318 (N_4318,N_3408,N_3759);
or U4319 (N_4319,N_3615,N_3767);
or U4320 (N_4320,N_3670,N_3673);
and U4321 (N_4321,N_3868,N_3699);
nor U4322 (N_4322,N_3968,N_3623);
or U4323 (N_4323,N_3538,N_3518);
nand U4324 (N_4324,N_3512,N_3252);
xor U4325 (N_4325,N_3980,N_3050);
and U4326 (N_4326,N_3985,N_3245);
nor U4327 (N_4327,N_3366,N_3028);
nor U4328 (N_4328,N_3087,N_3976);
or U4329 (N_4329,N_3136,N_3758);
nand U4330 (N_4330,N_3871,N_3548);
and U4331 (N_4331,N_3966,N_3817);
and U4332 (N_4332,N_3385,N_3638);
or U4333 (N_4333,N_3222,N_3207);
and U4334 (N_4334,N_3446,N_3839);
nor U4335 (N_4335,N_3987,N_3734);
nand U4336 (N_4336,N_3857,N_3824);
xnor U4337 (N_4337,N_3785,N_3882);
xnor U4338 (N_4338,N_3986,N_3752);
xor U4339 (N_4339,N_3234,N_3762);
nor U4340 (N_4340,N_3376,N_3047);
xor U4341 (N_4341,N_3893,N_3356);
nand U4342 (N_4342,N_3679,N_3407);
and U4343 (N_4343,N_3746,N_3206);
and U4344 (N_4344,N_3394,N_3528);
nand U4345 (N_4345,N_3727,N_3367);
nor U4346 (N_4346,N_3397,N_3361);
and U4347 (N_4347,N_3842,N_3579);
xor U4348 (N_4348,N_3314,N_3594);
and U4349 (N_4349,N_3262,N_3668);
or U4350 (N_4350,N_3106,N_3818);
and U4351 (N_4351,N_3707,N_3246);
nand U4352 (N_4352,N_3451,N_3119);
nor U4353 (N_4353,N_3825,N_3123);
nand U4354 (N_4354,N_3069,N_3777);
and U4355 (N_4355,N_3396,N_3051);
or U4356 (N_4356,N_3551,N_3781);
and U4357 (N_4357,N_3708,N_3267);
and U4358 (N_4358,N_3802,N_3009);
xnor U4359 (N_4359,N_3138,N_3915);
and U4360 (N_4360,N_3974,N_3288);
nand U4361 (N_4361,N_3399,N_3023);
xnor U4362 (N_4362,N_3733,N_3032);
and U4363 (N_4363,N_3860,N_3544);
or U4364 (N_4364,N_3587,N_3761);
and U4365 (N_4365,N_3965,N_3277);
nor U4366 (N_4366,N_3463,N_3605);
and U4367 (N_4367,N_3531,N_3843);
or U4368 (N_4368,N_3530,N_3562);
or U4369 (N_4369,N_3158,N_3062);
nor U4370 (N_4370,N_3035,N_3714);
nand U4371 (N_4371,N_3588,N_3873);
and U4372 (N_4372,N_3606,N_3270);
or U4373 (N_4373,N_3386,N_3285);
and U4374 (N_4374,N_3188,N_3239);
xnor U4375 (N_4375,N_3349,N_3219);
nor U4376 (N_4376,N_3199,N_3363);
and U4377 (N_4377,N_3804,N_3152);
and U4378 (N_4378,N_3621,N_3717);
xnor U4379 (N_4379,N_3650,N_3227);
xnor U4380 (N_4380,N_3827,N_3292);
nor U4381 (N_4381,N_3336,N_3936);
or U4382 (N_4382,N_3241,N_3998);
or U4383 (N_4383,N_3351,N_3745);
or U4384 (N_4384,N_3626,N_3052);
xor U4385 (N_4385,N_3190,N_3995);
or U4386 (N_4386,N_3470,N_3855);
nor U4387 (N_4387,N_3305,N_3888);
and U4388 (N_4388,N_3454,N_3442);
nand U4389 (N_4389,N_3665,N_3664);
xor U4390 (N_4390,N_3572,N_3603);
nand U4391 (N_4391,N_3330,N_3373);
and U4392 (N_4392,N_3690,N_3525);
nor U4393 (N_4393,N_3509,N_3317);
or U4394 (N_4394,N_3561,N_3726);
nor U4395 (N_4395,N_3982,N_3776);
xnor U4396 (N_4396,N_3889,N_3647);
nand U4397 (N_4397,N_3880,N_3678);
nand U4398 (N_4398,N_3036,N_3059);
nand U4399 (N_4399,N_3567,N_3906);
xnor U4400 (N_4400,N_3570,N_3629);
nand U4401 (N_4401,N_3563,N_3876);
xor U4402 (N_4402,N_3856,N_3228);
nor U4403 (N_4403,N_3456,N_3725);
nor U4404 (N_4404,N_3990,N_3433);
xor U4405 (N_4405,N_3217,N_3994);
or U4406 (N_4406,N_3686,N_3487);
or U4407 (N_4407,N_3931,N_3265);
or U4408 (N_4408,N_3612,N_3742);
xor U4409 (N_4409,N_3886,N_3439);
or U4410 (N_4410,N_3550,N_3173);
nand U4411 (N_4411,N_3044,N_3662);
xnor U4412 (N_4412,N_3652,N_3322);
nand U4413 (N_4413,N_3060,N_3184);
nor U4414 (N_4414,N_3730,N_3092);
xor U4415 (N_4415,N_3318,N_3053);
and U4416 (N_4416,N_3154,N_3582);
or U4417 (N_4417,N_3502,N_3672);
or U4418 (N_4418,N_3178,N_3085);
and U4419 (N_4419,N_3279,N_3304);
nand U4420 (N_4420,N_3796,N_3081);
or U4421 (N_4421,N_3522,N_3352);
and U4422 (N_4422,N_3991,N_3929);
nor U4423 (N_4423,N_3155,N_3061);
xor U4424 (N_4424,N_3308,N_3266);
or U4425 (N_4425,N_3095,N_3625);
or U4426 (N_4426,N_3573,N_3482);
xor U4427 (N_4427,N_3558,N_3609);
xnor U4428 (N_4428,N_3472,N_3348);
or U4429 (N_4429,N_3833,N_3064);
nor U4430 (N_4430,N_3215,N_3164);
nand U4431 (N_4431,N_3149,N_3075);
xnor U4432 (N_4432,N_3877,N_3486);
or U4433 (N_4433,N_3641,N_3139);
nand U4434 (N_4434,N_3310,N_3521);
or U4435 (N_4435,N_3795,N_3942);
xor U4436 (N_4436,N_3494,N_3321);
nand U4437 (N_4437,N_3346,N_3345);
and U4438 (N_4438,N_3172,N_3458);
or U4439 (N_4439,N_3602,N_3105);
and U4440 (N_4440,N_3559,N_3465);
nor U4441 (N_4441,N_3311,N_3225);
xnor U4442 (N_4442,N_3057,N_3425);
and U4443 (N_4443,N_3006,N_3932);
nor U4444 (N_4444,N_3757,N_3948);
or U4445 (N_4445,N_3218,N_3720);
xor U4446 (N_4446,N_3290,N_3365);
nor U4447 (N_4447,N_3413,N_3704);
and U4448 (N_4448,N_3194,N_3763);
xnor U4449 (N_4449,N_3258,N_3212);
and U4450 (N_4450,N_3205,N_3005);
nor U4451 (N_4451,N_3400,N_3420);
xor U4452 (N_4452,N_3200,N_3141);
and U4453 (N_4453,N_3535,N_3160);
or U4454 (N_4454,N_3735,N_3755);
or U4455 (N_4455,N_3591,N_3076);
nor U4456 (N_4456,N_3684,N_3286);
or U4457 (N_4457,N_3324,N_3989);
or U4458 (N_4458,N_3213,N_3179);
nand U4459 (N_4459,N_3816,N_3316);
nor U4460 (N_4460,N_3226,N_3914);
nor U4461 (N_4461,N_3555,N_3984);
nand U4462 (N_4462,N_3506,N_3617);
and U4463 (N_4463,N_3845,N_3649);
and U4464 (N_4464,N_3701,N_3344);
and U4465 (N_4465,N_3339,N_3299);
and U4466 (N_4466,N_3814,N_3599);
nor U4467 (N_4467,N_3951,N_3353);
or U4468 (N_4468,N_3340,N_3358);
and U4469 (N_4469,N_3127,N_3541);
xnor U4470 (N_4470,N_3335,N_3492);
nor U4471 (N_4471,N_3895,N_3493);
xor U4472 (N_4472,N_3894,N_3972);
nor U4473 (N_4473,N_3852,N_3850);
nor U4474 (N_4474,N_3883,N_3937);
nor U4475 (N_4475,N_3780,N_3438);
nand U4476 (N_4476,N_3379,N_3058);
nand U4477 (N_4477,N_3402,N_3240);
nand U4478 (N_4478,N_3094,N_3610);
and U4479 (N_4479,N_3001,N_3997);
xor U4480 (N_4480,N_3074,N_3145);
or U4481 (N_4481,N_3411,N_3938);
nor U4482 (N_4482,N_3418,N_3380);
xnor U4483 (N_4483,N_3904,N_3319);
nor U4484 (N_4484,N_3251,N_3274);
and U4485 (N_4485,N_3675,N_3510);
and U4486 (N_4486,N_3765,N_3022);
xnor U4487 (N_4487,N_3569,N_3669);
and U4488 (N_4488,N_3844,N_3789);
and U4489 (N_4489,N_3066,N_3004);
or U4490 (N_4490,N_3237,N_3372);
xor U4491 (N_4491,N_3024,N_3728);
nand U4492 (N_4492,N_3593,N_3167);
xnor U4493 (N_4493,N_3706,N_3303);
xnor U4494 (N_4494,N_3449,N_3919);
xnor U4495 (N_4495,N_3112,N_3072);
and U4496 (N_4496,N_3935,N_3556);
and U4497 (N_4497,N_3333,N_3008);
nand U4498 (N_4498,N_3566,N_3751);
and U4499 (N_4499,N_3357,N_3750);
or U4500 (N_4500,N_3050,N_3600);
nand U4501 (N_4501,N_3648,N_3930);
nor U4502 (N_4502,N_3461,N_3739);
nor U4503 (N_4503,N_3720,N_3127);
nand U4504 (N_4504,N_3252,N_3066);
or U4505 (N_4505,N_3790,N_3675);
and U4506 (N_4506,N_3172,N_3570);
and U4507 (N_4507,N_3795,N_3471);
and U4508 (N_4508,N_3596,N_3490);
xor U4509 (N_4509,N_3129,N_3168);
xor U4510 (N_4510,N_3903,N_3458);
xnor U4511 (N_4511,N_3849,N_3901);
and U4512 (N_4512,N_3423,N_3803);
nor U4513 (N_4513,N_3566,N_3189);
and U4514 (N_4514,N_3063,N_3318);
nand U4515 (N_4515,N_3861,N_3462);
nor U4516 (N_4516,N_3869,N_3550);
or U4517 (N_4517,N_3934,N_3704);
xor U4518 (N_4518,N_3333,N_3056);
or U4519 (N_4519,N_3308,N_3669);
nand U4520 (N_4520,N_3504,N_3325);
and U4521 (N_4521,N_3657,N_3513);
nor U4522 (N_4522,N_3185,N_3529);
or U4523 (N_4523,N_3201,N_3253);
or U4524 (N_4524,N_3981,N_3213);
xor U4525 (N_4525,N_3698,N_3771);
or U4526 (N_4526,N_3628,N_3437);
nand U4527 (N_4527,N_3430,N_3562);
or U4528 (N_4528,N_3662,N_3104);
or U4529 (N_4529,N_3440,N_3179);
and U4530 (N_4530,N_3413,N_3046);
nor U4531 (N_4531,N_3948,N_3488);
nor U4532 (N_4532,N_3777,N_3976);
xnor U4533 (N_4533,N_3462,N_3020);
nand U4534 (N_4534,N_3457,N_3539);
and U4535 (N_4535,N_3513,N_3185);
and U4536 (N_4536,N_3851,N_3070);
xnor U4537 (N_4537,N_3690,N_3817);
or U4538 (N_4538,N_3131,N_3890);
or U4539 (N_4539,N_3285,N_3750);
or U4540 (N_4540,N_3322,N_3075);
xor U4541 (N_4541,N_3248,N_3355);
nand U4542 (N_4542,N_3184,N_3437);
or U4543 (N_4543,N_3362,N_3964);
or U4544 (N_4544,N_3285,N_3563);
or U4545 (N_4545,N_3582,N_3609);
and U4546 (N_4546,N_3684,N_3307);
nand U4547 (N_4547,N_3893,N_3978);
xnor U4548 (N_4548,N_3505,N_3101);
and U4549 (N_4549,N_3057,N_3675);
nand U4550 (N_4550,N_3143,N_3418);
xnor U4551 (N_4551,N_3875,N_3786);
nor U4552 (N_4552,N_3452,N_3825);
or U4553 (N_4553,N_3402,N_3494);
xnor U4554 (N_4554,N_3252,N_3476);
nand U4555 (N_4555,N_3838,N_3344);
nor U4556 (N_4556,N_3374,N_3041);
or U4557 (N_4557,N_3128,N_3861);
and U4558 (N_4558,N_3638,N_3460);
or U4559 (N_4559,N_3019,N_3707);
or U4560 (N_4560,N_3860,N_3162);
xnor U4561 (N_4561,N_3951,N_3728);
and U4562 (N_4562,N_3537,N_3761);
xor U4563 (N_4563,N_3440,N_3205);
or U4564 (N_4564,N_3877,N_3301);
nand U4565 (N_4565,N_3675,N_3371);
nor U4566 (N_4566,N_3523,N_3639);
or U4567 (N_4567,N_3451,N_3730);
and U4568 (N_4568,N_3663,N_3212);
and U4569 (N_4569,N_3975,N_3770);
and U4570 (N_4570,N_3302,N_3297);
xor U4571 (N_4571,N_3700,N_3484);
xnor U4572 (N_4572,N_3209,N_3983);
nand U4573 (N_4573,N_3977,N_3637);
xor U4574 (N_4574,N_3939,N_3539);
and U4575 (N_4575,N_3069,N_3897);
xor U4576 (N_4576,N_3116,N_3626);
and U4577 (N_4577,N_3447,N_3072);
nor U4578 (N_4578,N_3806,N_3439);
xor U4579 (N_4579,N_3028,N_3434);
nand U4580 (N_4580,N_3633,N_3960);
or U4581 (N_4581,N_3937,N_3873);
nand U4582 (N_4582,N_3112,N_3473);
nand U4583 (N_4583,N_3284,N_3871);
nor U4584 (N_4584,N_3109,N_3616);
nor U4585 (N_4585,N_3686,N_3564);
nor U4586 (N_4586,N_3609,N_3125);
nand U4587 (N_4587,N_3932,N_3463);
nor U4588 (N_4588,N_3066,N_3171);
and U4589 (N_4589,N_3561,N_3252);
nor U4590 (N_4590,N_3208,N_3449);
xnor U4591 (N_4591,N_3826,N_3112);
nand U4592 (N_4592,N_3901,N_3054);
nor U4593 (N_4593,N_3698,N_3295);
xnor U4594 (N_4594,N_3528,N_3335);
xor U4595 (N_4595,N_3169,N_3276);
nand U4596 (N_4596,N_3937,N_3468);
and U4597 (N_4597,N_3269,N_3418);
xor U4598 (N_4598,N_3882,N_3538);
xnor U4599 (N_4599,N_3058,N_3019);
nand U4600 (N_4600,N_3140,N_3591);
and U4601 (N_4601,N_3701,N_3247);
xor U4602 (N_4602,N_3273,N_3020);
xor U4603 (N_4603,N_3222,N_3811);
and U4604 (N_4604,N_3912,N_3272);
and U4605 (N_4605,N_3985,N_3369);
nor U4606 (N_4606,N_3311,N_3702);
or U4607 (N_4607,N_3857,N_3993);
nand U4608 (N_4608,N_3995,N_3503);
and U4609 (N_4609,N_3761,N_3526);
and U4610 (N_4610,N_3506,N_3507);
or U4611 (N_4611,N_3200,N_3895);
xor U4612 (N_4612,N_3749,N_3970);
nor U4613 (N_4613,N_3817,N_3327);
and U4614 (N_4614,N_3676,N_3173);
nand U4615 (N_4615,N_3510,N_3103);
nand U4616 (N_4616,N_3503,N_3067);
or U4617 (N_4617,N_3388,N_3700);
nor U4618 (N_4618,N_3200,N_3656);
nor U4619 (N_4619,N_3112,N_3280);
xor U4620 (N_4620,N_3304,N_3394);
and U4621 (N_4621,N_3070,N_3532);
xor U4622 (N_4622,N_3997,N_3654);
and U4623 (N_4623,N_3230,N_3988);
or U4624 (N_4624,N_3466,N_3619);
xnor U4625 (N_4625,N_3558,N_3570);
nor U4626 (N_4626,N_3801,N_3593);
xnor U4627 (N_4627,N_3304,N_3496);
nor U4628 (N_4628,N_3155,N_3722);
xor U4629 (N_4629,N_3943,N_3418);
nand U4630 (N_4630,N_3465,N_3595);
nor U4631 (N_4631,N_3368,N_3560);
xor U4632 (N_4632,N_3486,N_3215);
and U4633 (N_4633,N_3744,N_3331);
and U4634 (N_4634,N_3670,N_3480);
or U4635 (N_4635,N_3514,N_3121);
xor U4636 (N_4636,N_3087,N_3441);
nand U4637 (N_4637,N_3244,N_3651);
nor U4638 (N_4638,N_3238,N_3497);
nand U4639 (N_4639,N_3908,N_3533);
nor U4640 (N_4640,N_3074,N_3260);
nand U4641 (N_4641,N_3859,N_3170);
and U4642 (N_4642,N_3985,N_3851);
nor U4643 (N_4643,N_3330,N_3438);
xnor U4644 (N_4644,N_3087,N_3523);
or U4645 (N_4645,N_3715,N_3110);
or U4646 (N_4646,N_3290,N_3468);
nor U4647 (N_4647,N_3333,N_3113);
nor U4648 (N_4648,N_3619,N_3193);
xnor U4649 (N_4649,N_3707,N_3219);
xnor U4650 (N_4650,N_3586,N_3275);
and U4651 (N_4651,N_3783,N_3756);
and U4652 (N_4652,N_3520,N_3916);
or U4653 (N_4653,N_3975,N_3177);
xor U4654 (N_4654,N_3389,N_3409);
or U4655 (N_4655,N_3461,N_3149);
nand U4656 (N_4656,N_3688,N_3139);
nor U4657 (N_4657,N_3796,N_3836);
and U4658 (N_4658,N_3890,N_3884);
xor U4659 (N_4659,N_3294,N_3449);
and U4660 (N_4660,N_3033,N_3713);
and U4661 (N_4661,N_3018,N_3249);
xor U4662 (N_4662,N_3531,N_3314);
nor U4663 (N_4663,N_3667,N_3580);
or U4664 (N_4664,N_3335,N_3741);
nor U4665 (N_4665,N_3542,N_3388);
and U4666 (N_4666,N_3599,N_3777);
nand U4667 (N_4667,N_3076,N_3706);
nor U4668 (N_4668,N_3253,N_3777);
xor U4669 (N_4669,N_3414,N_3539);
or U4670 (N_4670,N_3485,N_3476);
or U4671 (N_4671,N_3772,N_3167);
or U4672 (N_4672,N_3948,N_3674);
nor U4673 (N_4673,N_3987,N_3858);
or U4674 (N_4674,N_3213,N_3413);
nand U4675 (N_4675,N_3535,N_3780);
xor U4676 (N_4676,N_3260,N_3653);
nor U4677 (N_4677,N_3075,N_3131);
or U4678 (N_4678,N_3283,N_3353);
nor U4679 (N_4679,N_3760,N_3006);
or U4680 (N_4680,N_3494,N_3682);
nor U4681 (N_4681,N_3039,N_3371);
nand U4682 (N_4682,N_3326,N_3425);
and U4683 (N_4683,N_3695,N_3500);
or U4684 (N_4684,N_3897,N_3598);
nand U4685 (N_4685,N_3490,N_3122);
xnor U4686 (N_4686,N_3690,N_3889);
xnor U4687 (N_4687,N_3294,N_3115);
and U4688 (N_4688,N_3841,N_3232);
or U4689 (N_4689,N_3507,N_3022);
xor U4690 (N_4690,N_3431,N_3840);
and U4691 (N_4691,N_3942,N_3392);
xnor U4692 (N_4692,N_3552,N_3128);
nor U4693 (N_4693,N_3517,N_3311);
and U4694 (N_4694,N_3183,N_3927);
nand U4695 (N_4695,N_3420,N_3164);
nand U4696 (N_4696,N_3067,N_3944);
xnor U4697 (N_4697,N_3367,N_3822);
nand U4698 (N_4698,N_3329,N_3817);
or U4699 (N_4699,N_3415,N_3073);
nor U4700 (N_4700,N_3898,N_3035);
and U4701 (N_4701,N_3624,N_3714);
xnor U4702 (N_4702,N_3747,N_3179);
nor U4703 (N_4703,N_3592,N_3067);
or U4704 (N_4704,N_3948,N_3735);
nor U4705 (N_4705,N_3238,N_3163);
and U4706 (N_4706,N_3211,N_3246);
nor U4707 (N_4707,N_3007,N_3776);
or U4708 (N_4708,N_3295,N_3713);
nor U4709 (N_4709,N_3128,N_3179);
xnor U4710 (N_4710,N_3320,N_3778);
or U4711 (N_4711,N_3749,N_3772);
nor U4712 (N_4712,N_3545,N_3620);
or U4713 (N_4713,N_3592,N_3130);
nor U4714 (N_4714,N_3125,N_3606);
nand U4715 (N_4715,N_3057,N_3131);
xor U4716 (N_4716,N_3979,N_3239);
nor U4717 (N_4717,N_3089,N_3092);
nand U4718 (N_4718,N_3191,N_3059);
or U4719 (N_4719,N_3119,N_3181);
nand U4720 (N_4720,N_3249,N_3314);
nor U4721 (N_4721,N_3512,N_3095);
nor U4722 (N_4722,N_3833,N_3075);
xor U4723 (N_4723,N_3462,N_3961);
nand U4724 (N_4724,N_3255,N_3251);
xor U4725 (N_4725,N_3036,N_3142);
nand U4726 (N_4726,N_3053,N_3093);
and U4727 (N_4727,N_3577,N_3492);
or U4728 (N_4728,N_3169,N_3148);
xnor U4729 (N_4729,N_3969,N_3745);
nand U4730 (N_4730,N_3293,N_3750);
nor U4731 (N_4731,N_3750,N_3650);
xnor U4732 (N_4732,N_3712,N_3272);
or U4733 (N_4733,N_3173,N_3964);
and U4734 (N_4734,N_3694,N_3659);
or U4735 (N_4735,N_3210,N_3600);
or U4736 (N_4736,N_3485,N_3078);
and U4737 (N_4737,N_3570,N_3235);
nor U4738 (N_4738,N_3616,N_3716);
nand U4739 (N_4739,N_3812,N_3395);
and U4740 (N_4740,N_3198,N_3076);
and U4741 (N_4741,N_3503,N_3841);
and U4742 (N_4742,N_3477,N_3794);
and U4743 (N_4743,N_3167,N_3013);
or U4744 (N_4744,N_3822,N_3752);
nor U4745 (N_4745,N_3323,N_3516);
nor U4746 (N_4746,N_3056,N_3920);
and U4747 (N_4747,N_3296,N_3258);
nor U4748 (N_4748,N_3273,N_3393);
nor U4749 (N_4749,N_3288,N_3024);
nor U4750 (N_4750,N_3222,N_3394);
nand U4751 (N_4751,N_3552,N_3455);
xnor U4752 (N_4752,N_3671,N_3977);
and U4753 (N_4753,N_3575,N_3705);
and U4754 (N_4754,N_3491,N_3200);
nand U4755 (N_4755,N_3105,N_3398);
nor U4756 (N_4756,N_3072,N_3867);
nor U4757 (N_4757,N_3072,N_3693);
xor U4758 (N_4758,N_3655,N_3296);
and U4759 (N_4759,N_3486,N_3012);
or U4760 (N_4760,N_3751,N_3464);
and U4761 (N_4761,N_3854,N_3850);
nand U4762 (N_4762,N_3841,N_3681);
xnor U4763 (N_4763,N_3506,N_3366);
xor U4764 (N_4764,N_3069,N_3482);
nand U4765 (N_4765,N_3425,N_3451);
or U4766 (N_4766,N_3775,N_3567);
and U4767 (N_4767,N_3156,N_3783);
and U4768 (N_4768,N_3597,N_3404);
nand U4769 (N_4769,N_3293,N_3121);
nand U4770 (N_4770,N_3198,N_3776);
nor U4771 (N_4771,N_3744,N_3935);
nor U4772 (N_4772,N_3755,N_3733);
or U4773 (N_4773,N_3568,N_3862);
and U4774 (N_4774,N_3103,N_3005);
nand U4775 (N_4775,N_3178,N_3271);
xor U4776 (N_4776,N_3265,N_3028);
or U4777 (N_4777,N_3536,N_3255);
or U4778 (N_4778,N_3727,N_3172);
nor U4779 (N_4779,N_3687,N_3359);
xor U4780 (N_4780,N_3117,N_3125);
and U4781 (N_4781,N_3359,N_3271);
xnor U4782 (N_4782,N_3952,N_3275);
or U4783 (N_4783,N_3492,N_3432);
or U4784 (N_4784,N_3038,N_3313);
nand U4785 (N_4785,N_3709,N_3494);
xnor U4786 (N_4786,N_3126,N_3795);
and U4787 (N_4787,N_3744,N_3795);
xor U4788 (N_4788,N_3151,N_3884);
nand U4789 (N_4789,N_3506,N_3482);
nand U4790 (N_4790,N_3834,N_3382);
or U4791 (N_4791,N_3644,N_3396);
nand U4792 (N_4792,N_3057,N_3523);
and U4793 (N_4793,N_3602,N_3771);
and U4794 (N_4794,N_3482,N_3590);
xor U4795 (N_4795,N_3316,N_3031);
and U4796 (N_4796,N_3246,N_3853);
or U4797 (N_4797,N_3390,N_3804);
nand U4798 (N_4798,N_3567,N_3223);
xnor U4799 (N_4799,N_3332,N_3844);
nand U4800 (N_4800,N_3543,N_3309);
xnor U4801 (N_4801,N_3991,N_3968);
nand U4802 (N_4802,N_3785,N_3054);
and U4803 (N_4803,N_3900,N_3867);
xnor U4804 (N_4804,N_3482,N_3708);
or U4805 (N_4805,N_3239,N_3904);
xnor U4806 (N_4806,N_3125,N_3619);
and U4807 (N_4807,N_3162,N_3241);
nor U4808 (N_4808,N_3499,N_3814);
xnor U4809 (N_4809,N_3739,N_3639);
nand U4810 (N_4810,N_3372,N_3975);
nand U4811 (N_4811,N_3906,N_3293);
nand U4812 (N_4812,N_3632,N_3478);
or U4813 (N_4813,N_3374,N_3785);
and U4814 (N_4814,N_3568,N_3415);
or U4815 (N_4815,N_3683,N_3216);
nand U4816 (N_4816,N_3670,N_3380);
or U4817 (N_4817,N_3946,N_3658);
nand U4818 (N_4818,N_3282,N_3841);
nor U4819 (N_4819,N_3306,N_3539);
or U4820 (N_4820,N_3903,N_3522);
and U4821 (N_4821,N_3534,N_3002);
nor U4822 (N_4822,N_3240,N_3413);
or U4823 (N_4823,N_3359,N_3933);
and U4824 (N_4824,N_3946,N_3323);
xnor U4825 (N_4825,N_3241,N_3589);
and U4826 (N_4826,N_3222,N_3803);
or U4827 (N_4827,N_3756,N_3321);
or U4828 (N_4828,N_3149,N_3697);
xnor U4829 (N_4829,N_3940,N_3730);
nor U4830 (N_4830,N_3941,N_3373);
xnor U4831 (N_4831,N_3001,N_3072);
and U4832 (N_4832,N_3579,N_3808);
nor U4833 (N_4833,N_3565,N_3603);
nand U4834 (N_4834,N_3979,N_3632);
nor U4835 (N_4835,N_3212,N_3325);
or U4836 (N_4836,N_3293,N_3067);
xor U4837 (N_4837,N_3859,N_3882);
xor U4838 (N_4838,N_3201,N_3371);
nand U4839 (N_4839,N_3541,N_3097);
or U4840 (N_4840,N_3061,N_3738);
and U4841 (N_4841,N_3982,N_3203);
nand U4842 (N_4842,N_3333,N_3456);
nor U4843 (N_4843,N_3952,N_3405);
xnor U4844 (N_4844,N_3044,N_3354);
or U4845 (N_4845,N_3766,N_3285);
and U4846 (N_4846,N_3935,N_3453);
or U4847 (N_4847,N_3003,N_3510);
nand U4848 (N_4848,N_3591,N_3137);
and U4849 (N_4849,N_3175,N_3815);
nor U4850 (N_4850,N_3261,N_3369);
and U4851 (N_4851,N_3627,N_3440);
or U4852 (N_4852,N_3052,N_3972);
nor U4853 (N_4853,N_3694,N_3264);
xor U4854 (N_4854,N_3144,N_3586);
nand U4855 (N_4855,N_3761,N_3447);
nor U4856 (N_4856,N_3757,N_3136);
and U4857 (N_4857,N_3551,N_3369);
nor U4858 (N_4858,N_3158,N_3518);
nor U4859 (N_4859,N_3955,N_3241);
or U4860 (N_4860,N_3889,N_3225);
nor U4861 (N_4861,N_3428,N_3199);
nor U4862 (N_4862,N_3756,N_3497);
or U4863 (N_4863,N_3352,N_3619);
nand U4864 (N_4864,N_3928,N_3420);
and U4865 (N_4865,N_3794,N_3271);
or U4866 (N_4866,N_3846,N_3952);
nand U4867 (N_4867,N_3197,N_3602);
nand U4868 (N_4868,N_3933,N_3668);
nor U4869 (N_4869,N_3831,N_3428);
nand U4870 (N_4870,N_3991,N_3741);
xor U4871 (N_4871,N_3376,N_3117);
nor U4872 (N_4872,N_3237,N_3207);
nand U4873 (N_4873,N_3631,N_3504);
nor U4874 (N_4874,N_3510,N_3376);
and U4875 (N_4875,N_3448,N_3205);
and U4876 (N_4876,N_3287,N_3669);
nand U4877 (N_4877,N_3754,N_3788);
xnor U4878 (N_4878,N_3640,N_3351);
nor U4879 (N_4879,N_3571,N_3997);
nor U4880 (N_4880,N_3680,N_3877);
nand U4881 (N_4881,N_3956,N_3069);
nand U4882 (N_4882,N_3646,N_3633);
or U4883 (N_4883,N_3903,N_3927);
nor U4884 (N_4884,N_3758,N_3034);
and U4885 (N_4885,N_3655,N_3035);
nand U4886 (N_4886,N_3219,N_3997);
and U4887 (N_4887,N_3092,N_3040);
nor U4888 (N_4888,N_3130,N_3505);
xor U4889 (N_4889,N_3139,N_3212);
or U4890 (N_4890,N_3035,N_3542);
and U4891 (N_4891,N_3221,N_3533);
or U4892 (N_4892,N_3445,N_3831);
xnor U4893 (N_4893,N_3395,N_3298);
xor U4894 (N_4894,N_3934,N_3262);
nor U4895 (N_4895,N_3393,N_3767);
nor U4896 (N_4896,N_3158,N_3246);
xor U4897 (N_4897,N_3857,N_3331);
xnor U4898 (N_4898,N_3964,N_3482);
or U4899 (N_4899,N_3466,N_3386);
or U4900 (N_4900,N_3872,N_3985);
xnor U4901 (N_4901,N_3982,N_3232);
xnor U4902 (N_4902,N_3215,N_3872);
and U4903 (N_4903,N_3623,N_3242);
xor U4904 (N_4904,N_3634,N_3691);
xor U4905 (N_4905,N_3243,N_3571);
xnor U4906 (N_4906,N_3035,N_3827);
or U4907 (N_4907,N_3436,N_3315);
xor U4908 (N_4908,N_3521,N_3082);
and U4909 (N_4909,N_3128,N_3558);
or U4910 (N_4910,N_3354,N_3876);
nor U4911 (N_4911,N_3601,N_3086);
nand U4912 (N_4912,N_3065,N_3074);
or U4913 (N_4913,N_3491,N_3150);
and U4914 (N_4914,N_3371,N_3427);
nor U4915 (N_4915,N_3122,N_3989);
xor U4916 (N_4916,N_3722,N_3279);
xnor U4917 (N_4917,N_3276,N_3699);
xnor U4918 (N_4918,N_3998,N_3302);
nor U4919 (N_4919,N_3975,N_3301);
and U4920 (N_4920,N_3912,N_3557);
nor U4921 (N_4921,N_3364,N_3969);
or U4922 (N_4922,N_3013,N_3274);
xnor U4923 (N_4923,N_3434,N_3598);
and U4924 (N_4924,N_3605,N_3253);
and U4925 (N_4925,N_3276,N_3779);
nand U4926 (N_4926,N_3415,N_3916);
and U4927 (N_4927,N_3301,N_3557);
and U4928 (N_4928,N_3858,N_3814);
or U4929 (N_4929,N_3275,N_3563);
nor U4930 (N_4930,N_3061,N_3076);
and U4931 (N_4931,N_3176,N_3836);
or U4932 (N_4932,N_3204,N_3040);
xor U4933 (N_4933,N_3562,N_3837);
xnor U4934 (N_4934,N_3887,N_3376);
nand U4935 (N_4935,N_3216,N_3386);
nor U4936 (N_4936,N_3949,N_3619);
nand U4937 (N_4937,N_3438,N_3638);
nor U4938 (N_4938,N_3130,N_3482);
or U4939 (N_4939,N_3605,N_3241);
or U4940 (N_4940,N_3815,N_3229);
and U4941 (N_4941,N_3220,N_3771);
nand U4942 (N_4942,N_3888,N_3233);
xnor U4943 (N_4943,N_3956,N_3774);
nor U4944 (N_4944,N_3846,N_3969);
or U4945 (N_4945,N_3513,N_3116);
nor U4946 (N_4946,N_3257,N_3617);
or U4947 (N_4947,N_3687,N_3084);
xnor U4948 (N_4948,N_3414,N_3595);
or U4949 (N_4949,N_3948,N_3142);
and U4950 (N_4950,N_3104,N_3503);
nor U4951 (N_4951,N_3549,N_3139);
or U4952 (N_4952,N_3856,N_3301);
nor U4953 (N_4953,N_3222,N_3560);
or U4954 (N_4954,N_3331,N_3672);
xnor U4955 (N_4955,N_3227,N_3823);
nand U4956 (N_4956,N_3233,N_3524);
nand U4957 (N_4957,N_3296,N_3805);
xor U4958 (N_4958,N_3823,N_3522);
nand U4959 (N_4959,N_3809,N_3103);
nand U4960 (N_4960,N_3032,N_3761);
xor U4961 (N_4961,N_3097,N_3902);
xnor U4962 (N_4962,N_3151,N_3378);
xnor U4963 (N_4963,N_3752,N_3064);
nand U4964 (N_4964,N_3812,N_3509);
or U4965 (N_4965,N_3184,N_3511);
nor U4966 (N_4966,N_3915,N_3215);
or U4967 (N_4967,N_3316,N_3354);
or U4968 (N_4968,N_3104,N_3549);
nand U4969 (N_4969,N_3001,N_3092);
or U4970 (N_4970,N_3744,N_3049);
nand U4971 (N_4971,N_3814,N_3208);
nand U4972 (N_4972,N_3359,N_3026);
xnor U4973 (N_4973,N_3418,N_3621);
xor U4974 (N_4974,N_3682,N_3731);
nor U4975 (N_4975,N_3446,N_3761);
nand U4976 (N_4976,N_3950,N_3277);
nand U4977 (N_4977,N_3612,N_3888);
or U4978 (N_4978,N_3587,N_3785);
or U4979 (N_4979,N_3195,N_3137);
nor U4980 (N_4980,N_3871,N_3017);
nor U4981 (N_4981,N_3386,N_3177);
and U4982 (N_4982,N_3639,N_3755);
and U4983 (N_4983,N_3533,N_3842);
or U4984 (N_4984,N_3564,N_3892);
or U4985 (N_4985,N_3104,N_3922);
xnor U4986 (N_4986,N_3806,N_3793);
nand U4987 (N_4987,N_3617,N_3580);
or U4988 (N_4988,N_3488,N_3596);
or U4989 (N_4989,N_3921,N_3027);
and U4990 (N_4990,N_3943,N_3749);
and U4991 (N_4991,N_3233,N_3217);
and U4992 (N_4992,N_3644,N_3047);
nor U4993 (N_4993,N_3952,N_3003);
nor U4994 (N_4994,N_3923,N_3110);
xor U4995 (N_4995,N_3707,N_3140);
nor U4996 (N_4996,N_3684,N_3198);
or U4997 (N_4997,N_3059,N_3237);
and U4998 (N_4998,N_3395,N_3245);
xnor U4999 (N_4999,N_3792,N_3511);
xor U5000 (N_5000,N_4754,N_4136);
or U5001 (N_5001,N_4057,N_4684);
xnor U5002 (N_5002,N_4573,N_4047);
nor U5003 (N_5003,N_4264,N_4553);
nand U5004 (N_5004,N_4256,N_4990);
nand U5005 (N_5005,N_4963,N_4392);
nand U5006 (N_5006,N_4725,N_4055);
and U5007 (N_5007,N_4132,N_4336);
or U5008 (N_5008,N_4560,N_4289);
or U5009 (N_5009,N_4751,N_4495);
and U5010 (N_5010,N_4121,N_4109);
or U5011 (N_5011,N_4740,N_4664);
or U5012 (N_5012,N_4155,N_4983);
or U5013 (N_5013,N_4561,N_4004);
nand U5014 (N_5014,N_4158,N_4802);
or U5015 (N_5015,N_4532,N_4451);
and U5016 (N_5016,N_4596,N_4605);
nand U5017 (N_5017,N_4301,N_4753);
nor U5018 (N_5018,N_4575,N_4512);
and U5019 (N_5019,N_4654,N_4290);
nand U5020 (N_5020,N_4675,N_4000);
nor U5021 (N_5021,N_4460,N_4316);
nand U5022 (N_5022,N_4978,N_4120);
nor U5023 (N_5023,N_4080,N_4430);
xor U5024 (N_5024,N_4717,N_4019);
and U5025 (N_5025,N_4199,N_4036);
nand U5026 (N_5026,N_4448,N_4953);
xor U5027 (N_5027,N_4169,N_4240);
nor U5028 (N_5028,N_4563,N_4422);
nand U5029 (N_5029,N_4239,N_4462);
nand U5030 (N_5030,N_4585,N_4966);
or U5031 (N_5031,N_4639,N_4022);
xnor U5032 (N_5032,N_4069,N_4837);
xor U5033 (N_5033,N_4649,N_4646);
xor U5034 (N_5034,N_4304,N_4117);
nand U5035 (N_5035,N_4008,N_4708);
nor U5036 (N_5036,N_4307,N_4214);
nand U5037 (N_5037,N_4326,N_4042);
or U5038 (N_5038,N_4072,N_4190);
and U5039 (N_5039,N_4597,N_4703);
nor U5040 (N_5040,N_4672,N_4181);
and U5041 (N_5041,N_4710,N_4828);
and U5042 (N_5042,N_4403,N_4295);
nor U5043 (N_5043,N_4712,N_4020);
or U5044 (N_5044,N_4807,N_4817);
and U5045 (N_5045,N_4051,N_4883);
nor U5046 (N_5046,N_4350,N_4258);
and U5047 (N_5047,N_4997,N_4780);
and U5048 (N_5048,N_4067,N_4732);
nand U5049 (N_5049,N_4523,N_4651);
nand U5050 (N_5050,N_4085,N_4416);
or U5051 (N_5051,N_4232,N_4777);
nor U5052 (N_5052,N_4506,N_4074);
and U5053 (N_5053,N_4477,N_4794);
or U5054 (N_5054,N_4832,N_4433);
nand U5055 (N_5055,N_4478,N_4619);
or U5056 (N_5056,N_4901,N_4251);
nand U5057 (N_5057,N_4156,N_4040);
or U5058 (N_5058,N_4670,N_4682);
and U5059 (N_5059,N_4125,N_4935);
nor U5060 (N_5060,N_4611,N_4988);
xor U5061 (N_5061,N_4458,N_4891);
nand U5062 (N_5062,N_4886,N_4441);
or U5063 (N_5063,N_4442,N_4187);
nand U5064 (N_5064,N_4185,N_4804);
nor U5065 (N_5065,N_4348,N_4652);
and U5066 (N_5066,N_4113,N_4438);
or U5067 (N_5067,N_4772,N_4513);
nand U5068 (N_5068,N_4775,N_4756);
and U5069 (N_5069,N_4905,N_4849);
nand U5070 (N_5070,N_4582,N_4724);
nor U5071 (N_5071,N_4218,N_4009);
nor U5072 (N_5072,N_4618,N_4558);
or U5073 (N_5073,N_4546,N_4273);
xnor U5074 (N_5074,N_4183,N_4936);
nand U5075 (N_5075,N_4059,N_4137);
nor U5076 (N_5076,N_4706,N_4736);
nand U5077 (N_5077,N_4249,N_4328);
nor U5078 (N_5078,N_4267,N_4269);
xnor U5079 (N_5079,N_4409,N_4954);
and U5080 (N_5080,N_4789,N_4228);
or U5081 (N_5081,N_4956,N_4788);
and U5082 (N_5082,N_4571,N_4225);
nor U5083 (N_5083,N_4075,N_4310);
or U5084 (N_5084,N_4327,N_4680);
and U5085 (N_5085,N_4588,N_4134);
xor U5086 (N_5086,N_4406,N_4146);
xor U5087 (N_5087,N_4078,N_4948);
nand U5088 (N_5088,N_4421,N_4385);
or U5089 (N_5089,N_4656,N_4705);
nor U5090 (N_5090,N_4130,N_4970);
nand U5091 (N_5091,N_4445,N_4917);
or U5092 (N_5092,N_4131,N_4084);
nand U5093 (N_5093,N_4070,N_4800);
or U5094 (N_5094,N_4398,N_4859);
or U5095 (N_5095,N_4115,N_4220);
xor U5096 (N_5096,N_4095,N_4524);
xor U5097 (N_5097,N_4037,N_4168);
nor U5098 (N_5098,N_4728,N_4570);
and U5099 (N_5099,N_4830,N_4241);
or U5100 (N_5100,N_4629,N_4707);
or U5101 (N_5101,N_4872,N_4016);
and U5102 (N_5102,N_4104,N_4870);
and U5103 (N_5103,N_4673,N_4934);
or U5104 (N_5104,N_4030,N_4925);
nor U5105 (N_5105,N_4400,N_4812);
nand U5106 (N_5106,N_4294,N_4052);
or U5107 (N_5107,N_4720,N_4973);
and U5108 (N_5108,N_4363,N_4873);
nor U5109 (N_5109,N_4292,N_4068);
and U5110 (N_5110,N_4391,N_4843);
xor U5111 (N_5111,N_4189,N_4617);
nor U5112 (N_5112,N_4029,N_4986);
nor U5113 (N_5113,N_4580,N_4345);
xor U5114 (N_5114,N_4894,N_4816);
or U5115 (N_5115,N_4315,N_4094);
and U5116 (N_5116,N_4924,N_4467);
nor U5117 (N_5117,N_4951,N_4144);
xnor U5118 (N_5118,N_4535,N_4834);
and U5119 (N_5119,N_4309,N_4425);
nand U5120 (N_5120,N_4965,N_4915);
or U5121 (N_5121,N_4152,N_4662);
xor U5122 (N_5122,N_4599,N_4469);
nand U5123 (N_5123,N_4685,N_4114);
nand U5124 (N_5124,N_4248,N_4261);
nor U5125 (N_5125,N_4919,N_4209);
xnor U5126 (N_5126,N_4317,N_4364);
xor U5127 (N_5127,N_4929,N_4669);
nor U5128 (N_5128,N_4922,N_4731);
or U5129 (N_5129,N_4291,N_4519);
nand U5130 (N_5130,N_4176,N_4063);
nor U5131 (N_5131,N_4449,N_4744);
and U5132 (N_5132,N_4244,N_4205);
nor U5133 (N_5133,N_4274,N_4033);
and U5134 (N_5134,N_4767,N_4394);
nor U5135 (N_5135,N_4116,N_4697);
or U5136 (N_5136,N_4481,N_4658);
xnor U5137 (N_5137,N_4921,N_4034);
nand U5138 (N_5138,N_4981,N_4982);
and U5139 (N_5139,N_4536,N_4678);
nor U5140 (N_5140,N_4738,N_4005);
nor U5141 (N_5141,N_4098,N_4322);
nand U5142 (N_5142,N_4522,N_4359);
xnor U5143 (N_5143,N_4444,N_4382);
and U5144 (N_5144,N_4024,N_4108);
and U5145 (N_5145,N_4056,N_4021);
nand U5146 (N_5146,N_4941,N_4340);
nand U5147 (N_5147,N_4845,N_4083);
nand U5148 (N_5148,N_4206,N_4112);
nand U5149 (N_5149,N_4607,N_4939);
nor U5150 (N_5150,N_4993,N_4610);
xnor U5151 (N_5151,N_4139,N_4353);
nand U5152 (N_5152,N_4344,N_4041);
nand U5153 (N_5153,N_4967,N_4552);
nand U5154 (N_5154,N_4930,N_4174);
nand U5155 (N_5155,N_4012,N_4170);
or U5156 (N_5156,N_4674,N_4735);
nand U5157 (N_5157,N_4857,N_4861);
and U5158 (N_5158,N_4491,N_4791);
xnor U5159 (N_5159,N_4479,N_4647);
xnor U5160 (N_5160,N_4908,N_4747);
nand U5161 (N_5161,N_4539,N_4025);
nand U5162 (N_5162,N_4381,N_4324);
or U5163 (N_5163,N_4903,N_4866);
nor U5164 (N_5164,N_4138,N_4395);
nor U5165 (N_5165,N_4200,N_4633);
and U5166 (N_5166,N_4475,N_4959);
or U5167 (N_5167,N_4334,N_4230);
or U5168 (N_5168,N_4171,N_4949);
or U5169 (N_5169,N_4792,N_4480);
nand U5170 (N_5170,N_4683,N_4627);
nand U5171 (N_5171,N_4361,N_4231);
and U5172 (N_5172,N_4823,N_4813);
nor U5173 (N_5173,N_4411,N_4691);
and U5174 (N_5174,N_4160,N_4594);
or U5175 (N_5175,N_4165,N_4003);
nand U5176 (N_5176,N_4124,N_4297);
xor U5177 (N_5177,N_4848,N_4592);
xor U5178 (N_5178,N_4579,N_4931);
nand U5179 (N_5179,N_4254,N_4383);
xor U5180 (N_5180,N_4219,N_4637);
xnor U5181 (N_5181,N_4825,N_4329);
and U5182 (N_5182,N_4100,N_4771);
nand U5183 (N_5183,N_4871,N_4576);
xor U5184 (N_5184,N_4975,N_4150);
nand U5185 (N_5185,N_4810,N_4584);
or U5186 (N_5186,N_4360,N_4096);
xnor U5187 (N_5187,N_4829,N_4679);
xor U5188 (N_5188,N_4201,N_4537);
and U5189 (N_5189,N_4408,N_4889);
nand U5190 (N_5190,N_4374,N_4060);
and U5191 (N_5191,N_4275,N_4314);
and U5192 (N_5192,N_4102,N_4636);
and U5193 (N_5193,N_4574,N_4803);
xor U5194 (N_5194,N_4958,N_4293);
xor U5195 (N_5195,N_4023,N_4841);
nor U5196 (N_5196,N_4875,N_4140);
and U5197 (N_5197,N_4373,N_4760);
nand U5198 (N_5198,N_4472,N_4991);
xor U5199 (N_5199,N_4362,N_4123);
xor U5200 (N_5200,N_4073,N_4884);
or U5201 (N_5201,N_4192,N_4031);
nand U5202 (N_5202,N_4427,N_4907);
and U5203 (N_5203,N_4699,N_4106);
nor U5204 (N_5204,N_4839,N_4370);
or U5205 (N_5205,N_4892,N_4835);
xor U5206 (N_5206,N_4867,N_4860);
or U5207 (N_5207,N_4711,N_4824);
or U5208 (N_5208,N_4577,N_4126);
nor U5209 (N_5209,N_4399,N_4818);
nand U5210 (N_5210,N_4940,N_4049);
xnor U5211 (N_5211,N_4904,N_4259);
or U5212 (N_5212,N_4628,N_4286);
nand U5213 (N_5213,N_4620,N_4253);
and U5214 (N_5214,N_4914,N_4271);
nor U5215 (N_5215,N_4238,N_4701);
and U5216 (N_5216,N_4644,N_4492);
nor U5217 (N_5217,N_4893,N_4497);
and U5218 (N_5218,N_4500,N_4581);
xnor U5219 (N_5219,N_4153,N_4962);
xor U5220 (N_5220,N_4346,N_4050);
and U5221 (N_5221,N_4105,N_4616);
nor U5222 (N_5222,N_4902,N_4053);
nor U5223 (N_5223,N_4635,N_4676);
or U5224 (N_5224,N_4811,N_4700);
and U5225 (N_5225,N_4778,N_4419);
xor U5226 (N_5226,N_4842,N_4226);
or U5227 (N_5227,N_4779,N_4081);
or U5228 (N_5228,N_4511,N_4013);
or U5229 (N_5229,N_4704,N_4531);
nand U5230 (N_5230,N_4739,N_4145);
nand U5231 (N_5231,N_4815,N_4749);
nor U5232 (N_5232,N_4526,N_4805);
xor U5233 (N_5233,N_4039,N_4379);
and U5234 (N_5234,N_4401,N_4452);
nand U5235 (N_5235,N_4543,N_4007);
xor U5236 (N_5236,N_4847,N_4242);
or U5237 (N_5237,N_4687,N_4957);
xor U5238 (N_5238,N_4337,N_4011);
or U5239 (N_5239,N_4177,N_4538);
and U5240 (N_5240,N_4509,N_4722);
nor U5241 (N_5241,N_4572,N_4061);
or U5242 (N_5242,N_4482,N_4439);
and U5243 (N_5243,N_4280,N_4974);
nor U5244 (N_5244,N_4786,N_4655);
or U5245 (N_5245,N_4721,N_4319);
nor U5246 (N_5246,N_4623,N_4766);
xnor U5247 (N_5247,N_4118,N_4376);
and U5248 (N_5248,N_4366,N_4955);
nor U5249 (N_5249,N_4626,N_4785);
and U5250 (N_5250,N_4456,N_4709);
xor U5251 (N_5251,N_4440,N_4593);
nor U5252 (N_5252,N_4354,N_4723);
and U5253 (N_5253,N_4947,N_4862);
nor U5254 (N_5254,N_4564,N_4799);
or U5255 (N_5255,N_4943,N_4534);
and U5256 (N_5256,N_4881,N_4255);
nand U5257 (N_5257,N_4279,N_4148);
xor U5258 (N_5258,N_4591,N_4417);
nor U5259 (N_5259,N_4303,N_4435);
nor U5260 (N_5260,N_4737,N_4562);
and U5261 (N_5261,N_4470,N_4542);
or U5262 (N_5262,N_4494,N_4496);
nand U5263 (N_5263,N_4236,N_4349);
and U5264 (N_5264,N_4393,N_4208);
and U5265 (N_5265,N_4686,N_4390);
or U5266 (N_5266,N_4634,N_4998);
nor U5267 (N_5267,N_4755,N_4846);
nand U5268 (N_5268,N_4550,N_4938);
xnor U5269 (N_5269,N_4787,N_4920);
and U5270 (N_5270,N_4325,N_4695);
nor U5271 (N_5271,N_4621,N_4426);
and U5272 (N_5272,N_4645,N_4223);
or U5273 (N_5273,N_4781,N_4485);
and U5274 (N_5274,N_4089,N_4266);
and U5275 (N_5275,N_4302,N_4412);
and U5276 (N_5276,N_4714,N_4850);
or U5277 (N_5277,N_4487,N_4194);
and U5278 (N_5278,N_4827,N_4882);
and U5279 (N_5279,N_4216,N_4224);
xnor U5280 (N_5280,N_4961,N_4263);
xor U5281 (N_5281,N_4899,N_4282);
or U5282 (N_5282,N_4630,N_4916);
nor U5283 (N_5283,N_4071,N_4260);
nor U5284 (N_5284,N_4567,N_4122);
or U5285 (N_5285,N_4151,N_4801);
nand U5286 (N_5286,N_4356,N_4471);
nor U5287 (N_5287,N_4212,N_4167);
nand U5288 (N_5288,N_4147,N_4418);
xnor U5289 (N_5289,N_4358,N_4368);
nand U5290 (N_5290,N_4213,N_4741);
or U5291 (N_5291,N_4520,N_4510);
nand U5292 (N_5292,N_4796,N_4692);
nand U5293 (N_5293,N_4643,N_4926);
xnor U5294 (N_5294,N_4141,N_4600);
xor U5295 (N_5295,N_4992,N_4461);
xnor U5296 (N_5296,N_4898,N_4525);
xor U5297 (N_5297,N_4343,N_4002);
and U5298 (N_5298,N_4864,N_4135);
nor U5299 (N_5299,N_4097,N_4854);
nand U5300 (N_5300,N_4589,N_4942);
or U5301 (N_5301,N_4464,N_4387);
or U5302 (N_5302,N_4198,N_4410);
nand U5303 (N_5303,N_4603,N_4615);
or U5304 (N_5304,N_4545,N_4027);
nand U5305 (N_5305,N_4822,N_4932);
xor U5306 (N_5306,N_4702,N_4038);
nand U5307 (N_5307,N_4838,N_4128);
nand U5308 (N_5308,N_4661,N_4046);
or U5309 (N_5309,N_4338,N_4006);
nand U5310 (N_5310,N_4308,N_4437);
or U5311 (N_5311,N_4878,N_4980);
or U5312 (N_5312,N_4272,N_4179);
or U5313 (N_5313,N_4415,N_4608);
or U5314 (N_5314,N_4809,N_4203);
or U5315 (N_5315,N_4484,N_4428);
or U5316 (N_5316,N_4378,N_4443);
nor U5317 (N_5317,N_4045,N_4770);
nor U5318 (N_5318,N_4602,N_4332);
or U5319 (N_5319,N_4587,N_4614);
and U5320 (N_5320,N_4211,N_4154);
nand U5321 (N_5321,N_4320,N_4210);
nand U5322 (N_5322,N_4950,N_4498);
nor U5323 (N_5323,N_4648,N_4227);
or U5324 (N_5324,N_4900,N_4222);
or U5325 (N_5325,N_4321,N_4129);
and U5326 (N_5326,N_4665,N_4668);
or U5327 (N_5327,N_4985,N_4814);
or U5328 (N_5328,N_4197,N_4969);
and U5329 (N_5329,N_4650,N_4434);
xnor U5330 (N_5330,N_4960,N_4971);
nor U5331 (N_5331,N_4119,N_4653);
xnor U5332 (N_5332,N_4195,N_4305);
and U5333 (N_5333,N_4166,N_4014);
nor U5334 (N_5334,N_4182,N_4952);
nor U5335 (N_5335,N_4968,N_4270);
xor U5336 (N_5336,N_4836,N_4143);
xor U5337 (N_5337,N_4331,N_4681);
xnor U5338 (N_5338,N_4516,N_4065);
nand U5339 (N_5339,N_4713,N_4459);
and U5340 (N_5340,N_4161,N_4554);
or U5341 (N_5341,N_4657,N_4099);
or U5342 (N_5342,N_4043,N_4734);
nand U5343 (N_5343,N_4312,N_4514);
nor U5344 (N_5344,N_4865,N_4501);
xor U5345 (N_5345,N_4246,N_4436);
or U5346 (N_5346,N_4624,N_4423);
nor U5347 (N_5347,N_4808,N_4396);
xor U5348 (N_5348,N_4503,N_4493);
and U5349 (N_5349,N_4162,N_4079);
nand U5350 (N_5350,N_4397,N_4429);
nor U5351 (N_5351,N_4609,N_4913);
nand U5352 (N_5352,N_4318,N_4508);
xnor U5353 (N_5353,N_4404,N_4698);
nor U5354 (N_5354,N_4660,N_4693);
and U5355 (N_5355,N_4107,N_4583);
and U5356 (N_5356,N_4278,N_4551);
or U5357 (N_5357,N_4446,N_4371);
and U5358 (N_5358,N_4111,N_4377);
and U5359 (N_5359,N_4869,N_4093);
nor U5360 (N_5360,N_4765,N_4530);
or U5361 (N_5361,N_4157,N_4001);
nand U5362 (N_5362,N_4405,N_4369);
and U5363 (N_5363,N_4262,N_4895);
and U5364 (N_5364,N_4752,N_4101);
xor U5365 (N_5365,N_4489,N_4245);
nand U5366 (N_5366,N_4910,N_4507);
nor U5367 (N_5367,N_4844,N_4795);
or U5368 (N_5368,N_4159,N_4454);
or U5369 (N_5369,N_4976,N_4880);
nor U5370 (N_5370,N_4759,N_4757);
and U5371 (N_5371,N_4298,N_4641);
xnor U5372 (N_5372,N_4287,N_4028);
or U5373 (N_5373,N_4252,N_4663);
and U5374 (N_5374,N_4389,N_4018);
and U5375 (N_5375,N_4745,N_4716);
nor U5376 (N_5376,N_4402,N_4521);
nand U5377 (N_5377,N_4424,N_4833);
and U5378 (N_5378,N_4384,N_4798);
and U5379 (N_5379,N_4453,N_4288);
and U5380 (N_5380,N_4149,N_4090);
nor U5381 (N_5381,N_4586,N_4659);
nand U5382 (N_5382,N_4887,N_4386);
and U5383 (N_5383,N_4927,N_4351);
xor U5384 (N_5384,N_4928,N_4933);
or U5385 (N_5385,N_4557,N_4502);
nand U5386 (N_5386,N_4622,N_4196);
nand U5387 (N_5387,N_4082,N_4533);
or U5388 (N_5388,N_4339,N_4549);
xnor U5389 (N_5389,N_4909,N_4284);
and U5390 (N_5390,N_4746,N_4473);
or U5391 (N_5391,N_4556,N_4776);
xnor U5392 (N_5392,N_4774,N_4868);
xnor U5393 (N_5393,N_4715,N_4568);
or U5394 (N_5394,N_4234,N_4946);
nor U5395 (N_5395,N_4504,N_4569);
nor U5396 (N_5396,N_4696,N_4235);
nand U5397 (N_5397,N_4186,N_4726);
nor U5398 (N_5398,N_4127,N_4979);
and U5399 (N_5399,N_4667,N_4207);
nor U5400 (N_5400,N_4215,N_4283);
xnor U5401 (N_5401,N_4202,N_4483);
nor U5402 (N_5402,N_4265,N_4595);
nand U5403 (N_5403,N_4229,N_4897);
and U5404 (N_5404,N_4335,N_4355);
nor U5405 (N_5405,N_4277,N_4996);
xnor U5406 (N_5406,N_4555,N_4853);
xnor U5407 (N_5407,N_4888,N_4413);
nor U5408 (N_5408,N_4247,N_4450);
nand U5409 (N_5409,N_4233,N_4937);
nor U5410 (N_5410,N_4341,N_4468);
xnor U5411 (N_5411,N_4515,N_4086);
and U5412 (N_5412,N_4333,N_4856);
xnor U5413 (N_5413,N_4528,N_4819);
or U5414 (N_5414,N_4300,N_4237);
nand U5415 (N_5415,N_4764,N_4945);
xor U5416 (N_5416,N_4598,N_4110);
and U5417 (N_5417,N_4163,N_4742);
nor U5418 (N_5418,N_4457,N_4133);
xnor U5419 (N_5419,N_4944,N_4642);
xnor U5420 (N_5420,N_4748,N_4727);
nand U5421 (N_5421,N_4268,N_4204);
xnor U5422 (N_5422,N_4173,N_4342);
xnor U5423 (N_5423,N_4694,N_4250);
xor U5424 (N_5424,N_4999,N_4761);
nor U5425 (N_5425,N_4407,N_4763);
and U5426 (N_5426,N_4311,N_4414);
and U5427 (N_5427,N_4994,N_4666);
nor U5428 (N_5428,N_4372,N_4688);
xnor U5429 (N_5429,N_4730,N_4590);
nand U5430 (N_5430,N_4540,N_4172);
or U5431 (N_5431,N_4578,N_4911);
or U5432 (N_5432,N_4306,N_4296);
xor U5433 (N_5433,N_4631,N_4347);
nand U5434 (N_5434,N_4719,N_4505);
nor U5435 (N_5435,N_4517,N_4476);
nor U5436 (N_5436,N_4601,N_4367);
xor U5437 (N_5437,N_4010,N_4299);
nand U5438 (N_5438,N_4465,N_4048);
and U5439 (N_5439,N_4750,N_4768);
nor U5440 (N_5440,N_4490,N_4918);
or U5441 (N_5441,N_4032,N_4323);
nor U5442 (N_5442,N_4486,N_4964);
and U5443 (N_5443,N_4625,N_4455);
nor U5444 (N_5444,N_4026,N_4840);
or U5445 (N_5445,N_4221,N_4180);
xor U5446 (N_5446,N_4826,N_4066);
nor U5447 (N_5447,N_4175,N_4874);
or U5448 (N_5448,N_4877,N_4863);
nand U5449 (N_5449,N_4743,N_4671);
nor U5450 (N_5450,N_4977,N_4357);
nor U5451 (N_5451,N_4054,N_4548);
xnor U5452 (N_5452,N_4906,N_4447);
nor U5453 (N_5453,N_4474,N_4017);
or U5454 (N_5454,N_4432,N_4015);
and U5455 (N_5455,N_4488,N_4077);
nand U5456 (N_5456,N_4064,N_4879);
and U5457 (N_5457,N_4890,N_4689);
and U5458 (N_5458,N_4784,N_4518);
nor U5459 (N_5459,N_4876,N_4923);
or U5460 (N_5460,N_4544,N_4035);
or U5461 (N_5461,N_4547,N_4420);
or U5462 (N_5462,N_4885,N_4793);
or U5463 (N_5463,N_4790,N_4606);
and U5464 (N_5464,N_4638,N_4612);
nor U5465 (N_5465,N_4690,N_4380);
nor U5466 (N_5466,N_4821,N_4820);
and U5467 (N_5467,N_4529,N_4103);
xor U5468 (N_5468,N_4995,N_4188);
and U5469 (N_5469,N_4613,N_4718);
or U5470 (N_5470,N_4640,N_4257);
and U5471 (N_5471,N_4896,N_4388);
nor U5472 (N_5472,N_4044,N_4062);
nand U5473 (N_5473,N_4758,N_4851);
xor U5474 (N_5474,N_4769,N_4806);
xnor U5475 (N_5475,N_4058,N_4217);
xnor U5476 (N_5476,N_4729,N_4142);
or U5477 (N_5477,N_4912,N_4184);
or U5478 (N_5478,N_4285,N_4632);
nand U5479 (N_5479,N_4855,N_4375);
xor U5480 (N_5480,N_4565,N_4559);
nand U5481 (N_5481,N_4783,N_4677);
and U5482 (N_5482,N_4178,N_4831);
or U5483 (N_5483,N_4858,N_4852);
and U5484 (N_5484,N_4733,N_4527);
or U5485 (N_5485,N_4087,N_4276);
nor U5486 (N_5486,N_4541,N_4365);
nand U5487 (N_5487,N_4782,N_4313);
and U5488 (N_5488,N_4092,N_4193);
or U5489 (N_5489,N_4164,N_4243);
or U5490 (N_5490,N_4604,N_4281);
or U5491 (N_5491,N_4431,N_4797);
nand U5492 (N_5492,N_4352,N_4984);
or U5493 (N_5493,N_4773,N_4972);
xnor U5494 (N_5494,N_4330,N_4091);
or U5495 (N_5495,N_4566,N_4762);
or U5496 (N_5496,N_4499,N_4466);
or U5497 (N_5497,N_4987,N_4076);
nand U5498 (N_5498,N_4463,N_4191);
nor U5499 (N_5499,N_4989,N_4088);
nand U5500 (N_5500,N_4577,N_4704);
or U5501 (N_5501,N_4959,N_4786);
xnor U5502 (N_5502,N_4183,N_4997);
nor U5503 (N_5503,N_4132,N_4918);
xor U5504 (N_5504,N_4972,N_4901);
xor U5505 (N_5505,N_4167,N_4511);
or U5506 (N_5506,N_4983,N_4385);
xnor U5507 (N_5507,N_4745,N_4084);
nor U5508 (N_5508,N_4143,N_4429);
nand U5509 (N_5509,N_4286,N_4193);
and U5510 (N_5510,N_4296,N_4670);
nor U5511 (N_5511,N_4985,N_4291);
or U5512 (N_5512,N_4456,N_4648);
nor U5513 (N_5513,N_4055,N_4372);
nor U5514 (N_5514,N_4223,N_4921);
nand U5515 (N_5515,N_4230,N_4339);
nand U5516 (N_5516,N_4891,N_4551);
or U5517 (N_5517,N_4635,N_4208);
nand U5518 (N_5518,N_4616,N_4463);
xnor U5519 (N_5519,N_4178,N_4758);
nor U5520 (N_5520,N_4304,N_4725);
nand U5521 (N_5521,N_4056,N_4245);
nand U5522 (N_5522,N_4518,N_4046);
nand U5523 (N_5523,N_4614,N_4912);
xnor U5524 (N_5524,N_4590,N_4655);
nor U5525 (N_5525,N_4466,N_4032);
nand U5526 (N_5526,N_4151,N_4963);
and U5527 (N_5527,N_4186,N_4994);
or U5528 (N_5528,N_4261,N_4768);
nor U5529 (N_5529,N_4818,N_4476);
xor U5530 (N_5530,N_4811,N_4530);
nor U5531 (N_5531,N_4655,N_4025);
or U5532 (N_5532,N_4701,N_4398);
nor U5533 (N_5533,N_4594,N_4425);
or U5534 (N_5534,N_4666,N_4480);
and U5535 (N_5535,N_4067,N_4959);
and U5536 (N_5536,N_4380,N_4742);
or U5537 (N_5537,N_4979,N_4052);
nor U5538 (N_5538,N_4666,N_4675);
nor U5539 (N_5539,N_4684,N_4340);
and U5540 (N_5540,N_4227,N_4910);
nor U5541 (N_5541,N_4653,N_4782);
nand U5542 (N_5542,N_4659,N_4815);
and U5543 (N_5543,N_4362,N_4916);
nand U5544 (N_5544,N_4210,N_4136);
or U5545 (N_5545,N_4722,N_4583);
xnor U5546 (N_5546,N_4035,N_4239);
or U5547 (N_5547,N_4684,N_4098);
or U5548 (N_5548,N_4160,N_4778);
xor U5549 (N_5549,N_4637,N_4544);
and U5550 (N_5550,N_4292,N_4853);
and U5551 (N_5551,N_4427,N_4769);
or U5552 (N_5552,N_4069,N_4194);
and U5553 (N_5553,N_4044,N_4717);
and U5554 (N_5554,N_4039,N_4578);
xnor U5555 (N_5555,N_4344,N_4939);
nor U5556 (N_5556,N_4428,N_4371);
or U5557 (N_5557,N_4415,N_4328);
or U5558 (N_5558,N_4021,N_4389);
xor U5559 (N_5559,N_4677,N_4482);
and U5560 (N_5560,N_4952,N_4668);
nor U5561 (N_5561,N_4269,N_4037);
nand U5562 (N_5562,N_4664,N_4480);
and U5563 (N_5563,N_4660,N_4406);
or U5564 (N_5564,N_4835,N_4929);
xor U5565 (N_5565,N_4858,N_4011);
nand U5566 (N_5566,N_4859,N_4248);
or U5567 (N_5567,N_4366,N_4871);
and U5568 (N_5568,N_4796,N_4140);
or U5569 (N_5569,N_4854,N_4247);
and U5570 (N_5570,N_4847,N_4568);
or U5571 (N_5571,N_4743,N_4683);
xnor U5572 (N_5572,N_4143,N_4912);
or U5573 (N_5573,N_4656,N_4250);
and U5574 (N_5574,N_4874,N_4065);
and U5575 (N_5575,N_4269,N_4060);
nand U5576 (N_5576,N_4535,N_4821);
nor U5577 (N_5577,N_4812,N_4880);
and U5578 (N_5578,N_4628,N_4706);
nand U5579 (N_5579,N_4185,N_4229);
xor U5580 (N_5580,N_4679,N_4194);
or U5581 (N_5581,N_4350,N_4528);
or U5582 (N_5582,N_4996,N_4557);
nor U5583 (N_5583,N_4445,N_4771);
nand U5584 (N_5584,N_4908,N_4387);
or U5585 (N_5585,N_4021,N_4014);
xnor U5586 (N_5586,N_4621,N_4249);
and U5587 (N_5587,N_4802,N_4529);
and U5588 (N_5588,N_4632,N_4967);
nor U5589 (N_5589,N_4314,N_4242);
nor U5590 (N_5590,N_4477,N_4472);
nor U5591 (N_5591,N_4745,N_4010);
or U5592 (N_5592,N_4115,N_4628);
and U5593 (N_5593,N_4292,N_4759);
or U5594 (N_5594,N_4159,N_4449);
and U5595 (N_5595,N_4062,N_4704);
xnor U5596 (N_5596,N_4568,N_4073);
nand U5597 (N_5597,N_4800,N_4750);
or U5598 (N_5598,N_4378,N_4025);
nor U5599 (N_5599,N_4821,N_4983);
xor U5600 (N_5600,N_4875,N_4651);
nor U5601 (N_5601,N_4187,N_4788);
nand U5602 (N_5602,N_4714,N_4096);
xnor U5603 (N_5603,N_4154,N_4865);
and U5604 (N_5604,N_4488,N_4675);
xnor U5605 (N_5605,N_4739,N_4661);
xor U5606 (N_5606,N_4084,N_4413);
and U5607 (N_5607,N_4640,N_4368);
xor U5608 (N_5608,N_4779,N_4906);
and U5609 (N_5609,N_4232,N_4337);
or U5610 (N_5610,N_4784,N_4998);
nand U5611 (N_5611,N_4556,N_4613);
nor U5612 (N_5612,N_4007,N_4907);
xor U5613 (N_5613,N_4196,N_4634);
nor U5614 (N_5614,N_4350,N_4436);
xnor U5615 (N_5615,N_4579,N_4243);
nand U5616 (N_5616,N_4504,N_4044);
xor U5617 (N_5617,N_4688,N_4562);
xnor U5618 (N_5618,N_4610,N_4150);
nor U5619 (N_5619,N_4833,N_4601);
nor U5620 (N_5620,N_4801,N_4177);
nand U5621 (N_5621,N_4263,N_4118);
xnor U5622 (N_5622,N_4522,N_4653);
nor U5623 (N_5623,N_4009,N_4788);
nor U5624 (N_5624,N_4627,N_4054);
xnor U5625 (N_5625,N_4671,N_4643);
nand U5626 (N_5626,N_4589,N_4440);
xor U5627 (N_5627,N_4395,N_4878);
xnor U5628 (N_5628,N_4245,N_4433);
nand U5629 (N_5629,N_4945,N_4983);
nand U5630 (N_5630,N_4084,N_4682);
or U5631 (N_5631,N_4390,N_4098);
nand U5632 (N_5632,N_4116,N_4837);
and U5633 (N_5633,N_4983,N_4869);
nor U5634 (N_5634,N_4239,N_4583);
or U5635 (N_5635,N_4560,N_4861);
and U5636 (N_5636,N_4319,N_4260);
nand U5637 (N_5637,N_4084,N_4287);
or U5638 (N_5638,N_4962,N_4252);
nor U5639 (N_5639,N_4601,N_4841);
and U5640 (N_5640,N_4433,N_4788);
and U5641 (N_5641,N_4091,N_4241);
and U5642 (N_5642,N_4323,N_4246);
or U5643 (N_5643,N_4829,N_4338);
or U5644 (N_5644,N_4868,N_4822);
or U5645 (N_5645,N_4157,N_4511);
nand U5646 (N_5646,N_4871,N_4304);
nor U5647 (N_5647,N_4770,N_4713);
nand U5648 (N_5648,N_4769,N_4754);
or U5649 (N_5649,N_4469,N_4742);
and U5650 (N_5650,N_4127,N_4977);
nand U5651 (N_5651,N_4839,N_4022);
and U5652 (N_5652,N_4098,N_4937);
nor U5653 (N_5653,N_4216,N_4842);
nor U5654 (N_5654,N_4006,N_4269);
or U5655 (N_5655,N_4323,N_4268);
nor U5656 (N_5656,N_4753,N_4715);
nand U5657 (N_5657,N_4930,N_4387);
nand U5658 (N_5658,N_4501,N_4613);
nor U5659 (N_5659,N_4357,N_4573);
nor U5660 (N_5660,N_4979,N_4745);
nor U5661 (N_5661,N_4913,N_4968);
nand U5662 (N_5662,N_4289,N_4245);
xnor U5663 (N_5663,N_4018,N_4433);
and U5664 (N_5664,N_4897,N_4587);
and U5665 (N_5665,N_4613,N_4802);
nor U5666 (N_5666,N_4726,N_4747);
or U5667 (N_5667,N_4365,N_4305);
xnor U5668 (N_5668,N_4456,N_4368);
xor U5669 (N_5669,N_4239,N_4635);
nor U5670 (N_5670,N_4752,N_4660);
nor U5671 (N_5671,N_4694,N_4746);
nand U5672 (N_5672,N_4189,N_4049);
and U5673 (N_5673,N_4923,N_4310);
and U5674 (N_5674,N_4462,N_4045);
xor U5675 (N_5675,N_4624,N_4242);
xnor U5676 (N_5676,N_4589,N_4318);
nand U5677 (N_5677,N_4289,N_4559);
nor U5678 (N_5678,N_4855,N_4962);
and U5679 (N_5679,N_4903,N_4801);
and U5680 (N_5680,N_4190,N_4697);
and U5681 (N_5681,N_4702,N_4890);
and U5682 (N_5682,N_4210,N_4623);
nand U5683 (N_5683,N_4628,N_4076);
nor U5684 (N_5684,N_4690,N_4773);
and U5685 (N_5685,N_4935,N_4444);
or U5686 (N_5686,N_4649,N_4284);
and U5687 (N_5687,N_4550,N_4071);
and U5688 (N_5688,N_4522,N_4666);
or U5689 (N_5689,N_4015,N_4376);
nand U5690 (N_5690,N_4122,N_4452);
nand U5691 (N_5691,N_4252,N_4318);
nor U5692 (N_5692,N_4331,N_4793);
or U5693 (N_5693,N_4973,N_4997);
and U5694 (N_5694,N_4223,N_4692);
or U5695 (N_5695,N_4823,N_4192);
xor U5696 (N_5696,N_4448,N_4410);
nand U5697 (N_5697,N_4508,N_4452);
xor U5698 (N_5698,N_4376,N_4559);
nand U5699 (N_5699,N_4802,N_4496);
and U5700 (N_5700,N_4314,N_4468);
or U5701 (N_5701,N_4949,N_4052);
and U5702 (N_5702,N_4512,N_4141);
or U5703 (N_5703,N_4102,N_4722);
xnor U5704 (N_5704,N_4566,N_4123);
xnor U5705 (N_5705,N_4130,N_4882);
and U5706 (N_5706,N_4353,N_4757);
nor U5707 (N_5707,N_4408,N_4110);
or U5708 (N_5708,N_4391,N_4733);
nand U5709 (N_5709,N_4023,N_4335);
or U5710 (N_5710,N_4901,N_4296);
or U5711 (N_5711,N_4582,N_4217);
or U5712 (N_5712,N_4523,N_4657);
and U5713 (N_5713,N_4622,N_4814);
nor U5714 (N_5714,N_4234,N_4455);
or U5715 (N_5715,N_4144,N_4439);
and U5716 (N_5716,N_4015,N_4193);
nand U5717 (N_5717,N_4669,N_4645);
nor U5718 (N_5718,N_4012,N_4786);
and U5719 (N_5719,N_4802,N_4524);
and U5720 (N_5720,N_4457,N_4675);
xnor U5721 (N_5721,N_4358,N_4311);
nand U5722 (N_5722,N_4056,N_4214);
and U5723 (N_5723,N_4550,N_4524);
xor U5724 (N_5724,N_4214,N_4910);
and U5725 (N_5725,N_4304,N_4621);
nand U5726 (N_5726,N_4178,N_4316);
nand U5727 (N_5727,N_4082,N_4229);
nand U5728 (N_5728,N_4445,N_4498);
xor U5729 (N_5729,N_4328,N_4716);
nand U5730 (N_5730,N_4521,N_4954);
xor U5731 (N_5731,N_4968,N_4130);
nand U5732 (N_5732,N_4776,N_4145);
and U5733 (N_5733,N_4862,N_4840);
or U5734 (N_5734,N_4177,N_4254);
xnor U5735 (N_5735,N_4944,N_4665);
nand U5736 (N_5736,N_4622,N_4123);
and U5737 (N_5737,N_4715,N_4559);
and U5738 (N_5738,N_4150,N_4736);
and U5739 (N_5739,N_4126,N_4211);
or U5740 (N_5740,N_4740,N_4784);
nor U5741 (N_5741,N_4069,N_4517);
or U5742 (N_5742,N_4656,N_4467);
or U5743 (N_5743,N_4479,N_4396);
xnor U5744 (N_5744,N_4593,N_4330);
and U5745 (N_5745,N_4762,N_4037);
or U5746 (N_5746,N_4554,N_4516);
nand U5747 (N_5747,N_4345,N_4189);
xor U5748 (N_5748,N_4571,N_4123);
nor U5749 (N_5749,N_4246,N_4660);
xnor U5750 (N_5750,N_4795,N_4810);
xnor U5751 (N_5751,N_4138,N_4385);
xor U5752 (N_5752,N_4035,N_4231);
nand U5753 (N_5753,N_4240,N_4929);
nand U5754 (N_5754,N_4818,N_4563);
and U5755 (N_5755,N_4547,N_4419);
nand U5756 (N_5756,N_4163,N_4030);
nor U5757 (N_5757,N_4176,N_4276);
or U5758 (N_5758,N_4486,N_4321);
and U5759 (N_5759,N_4356,N_4747);
nand U5760 (N_5760,N_4280,N_4886);
or U5761 (N_5761,N_4628,N_4567);
xnor U5762 (N_5762,N_4315,N_4264);
nor U5763 (N_5763,N_4051,N_4153);
nor U5764 (N_5764,N_4567,N_4736);
xnor U5765 (N_5765,N_4371,N_4157);
and U5766 (N_5766,N_4824,N_4849);
or U5767 (N_5767,N_4668,N_4907);
nand U5768 (N_5768,N_4716,N_4055);
and U5769 (N_5769,N_4667,N_4823);
nand U5770 (N_5770,N_4907,N_4544);
nand U5771 (N_5771,N_4497,N_4037);
nand U5772 (N_5772,N_4825,N_4192);
xor U5773 (N_5773,N_4309,N_4928);
xnor U5774 (N_5774,N_4639,N_4398);
nor U5775 (N_5775,N_4514,N_4016);
and U5776 (N_5776,N_4720,N_4630);
nor U5777 (N_5777,N_4248,N_4047);
and U5778 (N_5778,N_4825,N_4332);
nor U5779 (N_5779,N_4011,N_4127);
nand U5780 (N_5780,N_4477,N_4609);
nand U5781 (N_5781,N_4892,N_4285);
or U5782 (N_5782,N_4873,N_4565);
and U5783 (N_5783,N_4013,N_4657);
xor U5784 (N_5784,N_4751,N_4955);
and U5785 (N_5785,N_4696,N_4029);
nand U5786 (N_5786,N_4061,N_4660);
or U5787 (N_5787,N_4079,N_4207);
or U5788 (N_5788,N_4705,N_4945);
xnor U5789 (N_5789,N_4662,N_4527);
nand U5790 (N_5790,N_4001,N_4978);
and U5791 (N_5791,N_4949,N_4068);
or U5792 (N_5792,N_4197,N_4131);
xor U5793 (N_5793,N_4770,N_4894);
xnor U5794 (N_5794,N_4478,N_4558);
nor U5795 (N_5795,N_4485,N_4129);
or U5796 (N_5796,N_4446,N_4294);
nor U5797 (N_5797,N_4308,N_4090);
or U5798 (N_5798,N_4525,N_4472);
nand U5799 (N_5799,N_4551,N_4897);
and U5800 (N_5800,N_4864,N_4764);
xor U5801 (N_5801,N_4089,N_4006);
xnor U5802 (N_5802,N_4607,N_4192);
nor U5803 (N_5803,N_4732,N_4277);
xnor U5804 (N_5804,N_4420,N_4184);
and U5805 (N_5805,N_4017,N_4271);
xor U5806 (N_5806,N_4540,N_4733);
or U5807 (N_5807,N_4267,N_4826);
nor U5808 (N_5808,N_4081,N_4559);
xor U5809 (N_5809,N_4042,N_4360);
nor U5810 (N_5810,N_4393,N_4960);
xor U5811 (N_5811,N_4910,N_4278);
or U5812 (N_5812,N_4832,N_4307);
nand U5813 (N_5813,N_4151,N_4479);
xor U5814 (N_5814,N_4213,N_4112);
nor U5815 (N_5815,N_4257,N_4802);
or U5816 (N_5816,N_4522,N_4401);
nor U5817 (N_5817,N_4904,N_4244);
xnor U5818 (N_5818,N_4633,N_4959);
nor U5819 (N_5819,N_4694,N_4725);
or U5820 (N_5820,N_4448,N_4873);
or U5821 (N_5821,N_4564,N_4381);
nand U5822 (N_5822,N_4792,N_4328);
or U5823 (N_5823,N_4849,N_4066);
or U5824 (N_5824,N_4065,N_4403);
nor U5825 (N_5825,N_4687,N_4316);
and U5826 (N_5826,N_4495,N_4191);
and U5827 (N_5827,N_4739,N_4268);
and U5828 (N_5828,N_4014,N_4897);
and U5829 (N_5829,N_4285,N_4604);
or U5830 (N_5830,N_4628,N_4899);
xor U5831 (N_5831,N_4255,N_4063);
nand U5832 (N_5832,N_4657,N_4297);
xnor U5833 (N_5833,N_4194,N_4490);
nand U5834 (N_5834,N_4182,N_4513);
and U5835 (N_5835,N_4488,N_4047);
nor U5836 (N_5836,N_4697,N_4556);
nor U5837 (N_5837,N_4959,N_4882);
nor U5838 (N_5838,N_4861,N_4425);
xor U5839 (N_5839,N_4970,N_4612);
nor U5840 (N_5840,N_4988,N_4524);
nor U5841 (N_5841,N_4950,N_4601);
nand U5842 (N_5842,N_4590,N_4794);
xor U5843 (N_5843,N_4391,N_4904);
nor U5844 (N_5844,N_4365,N_4731);
xnor U5845 (N_5845,N_4084,N_4665);
nor U5846 (N_5846,N_4902,N_4651);
nor U5847 (N_5847,N_4024,N_4799);
nand U5848 (N_5848,N_4984,N_4716);
and U5849 (N_5849,N_4502,N_4454);
and U5850 (N_5850,N_4983,N_4580);
xnor U5851 (N_5851,N_4609,N_4041);
and U5852 (N_5852,N_4297,N_4444);
and U5853 (N_5853,N_4569,N_4853);
xnor U5854 (N_5854,N_4421,N_4128);
and U5855 (N_5855,N_4675,N_4441);
nand U5856 (N_5856,N_4392,N_4716);
xnor U5857 (N_5857,N_4391,N_4729);
nand U5858 (N_5858,N_4047,N_4515);
or U5859 (N_5859,N_4034,N_4020);
nor U5860 (N_5860,N_4621,N_4899);
or U5861 (N_5861,N_4521,N_4766);
nor U5862 (N_5862,N_4092,N_4185);
and U5863 (N_5863,N_4533,N_4869);
nand U5864 (N_5864,N_4474,N_4215);
nor U5865 (N_5865,N_4093,N_4347);
nand U5866 (N_5866,N_4424,N_4571);
nor U5867 (N_5867,N_4236,N_4534);
or U5868 (N_5868,N_4445,N_4824);
xor U5869 (N_5869,N_4759,N_4708);
nand U5870 (N_5870,N_4402,N_4602);
or U5871 (N_5871,N_4434,N_4299);
xor U5872 (N_5872,N_4640,N_4326);
xor U5873 (N_5873,N_4959,N_4316);
nand U5874 (N_5874,N_4999,N_4612);
nor U5875 (N_5875,N_4706,N_4976);
or U5876 (N_5876,N_4391,N_4870);
or U5877 (N_5877,N_4788,N_4266);
and U5878 (N_5878,N_4706,N_4376);
nor U5879 (N_5879,N_4233,N_4840);
nor U5880 (N_5880,N_4959,N_4570);
or U5881 (N_5881,N_4066,N_4728);
and U5882 (N_5882,N_4265,N_4234);
nand U5883 (N_5883,N_4102,N_4094);
nor U5884 (N_5884,N_4608,N_4439);
nor U5885 (N_5885,N_4752,N_4836);
xnor U5886 (N_5886,N_4612,N_4071);
or U5887 (N_5887,N_4968,N_4336);
nand U5888 (N_5888,N_4056,N_4402);
nor U5889 (N_5889,N_4077,N_4292);
nand U5890 (N_5890,N_4262,N_4844);
xnor U5891 (N_5891,N_4282,N_4345);
or U5892 (N_5892,N_4068,N_4093);
xor U5893 (N_5893,N_4858,N_4630);
or U5894 (N_5894,N_4922,N_4170);
or U5895 (N_5895,N_4117,N_4131);
nand U5896 (N_5896,N_4790,N_4198);
or U5897 (N_5897,N_4899,N_4187);
or U5898 (N_5898,N_4655,N_4465);
nor U5899 (N_5899,N_4036,N_4743);
nor U5900 (N_5900,N_4195,N_4312);
and U5901 (N_5901,N_4695,N_4826);
nor U5902 (N_5902,N_4622,N_4687);
nand U5903 (N_5903,N_4571,N_4101);
and U5904 (N_5904,N_4182,N_4722);
and U5905 (N_5905,N_4394,N_4075);
nand U5906 (N_5906,N_4939,N_4605);
nand U5907 (N_5907,N_4736,N_4917);
and U5908 (N_5908,N_4421,N_4261);
xnor U5909 (N_5909,N_4761,N_4379);
and U5910 (N_5910,N_4952,N_4056);
nor U5911 (N_5911,N_4315,N_4406);
xor U5912 (N_5912,N_4927,N_4694);
nor U5913 (N_5913,N_4478,N_4686);
nand U5914 (N_5914,N_4411,N_4165);
and U5915 (N_5915,N_4212,N_4955);
and U5916 (N_5916,N_4071,N_4204);
nor U5917 (N_5917,N_4816,N_4699);
nor U5918 (N_5918,N_4992,N_4423);
xnor U5919 (N_5919,N_4655,N_4292);
nor U5920 (N_5920,N_4070,N_4701);
or U5921 (N_5921,N_4638,N_4036);
nand U5922 (N_5922,N_4582,N_4604);
xnor U5923 (N_5923,N_4226,N_4785);
nor U5924 (N_5924,N_4066,N_4918);
and U5925 (N_5925,N_4355,N_4628);
or U5926 (N_5926,N_4643,N_4795);
nor U5927 (N_5927,N_4601,N_4592);
and U5928 (N_5928,N_4992,N_4152);
or U5929 (N_5929,N_4337,N_4760);
nor U5930 (N_5930,N_4693,N_4102);
and U5931 (N_5931,N_4014,N_4657);
nand U5932 (N_5932,N_4464,N_4632);
nand U5933 (N_5933,N_4695,N_4257);
xor U5934 (N_5934,N_4692,N_4345);
nand U5935 (N_5935,N_4622,N_4118);
and U5936 (N_5936,N_4117,N_4210);
or U5937 (N_5937,N_4426,N_4267);
and U5938 (N_5938,N_4164,N_4838);
and U5939 (N_5939,N_4661,N_4073);
and U5940 (N_5940,N_4563,N_4743);
nand U5941 (N_5941,N_4031,N_4767);
nor U5942 (N_5942,N_4323,N_4203);
nor U5943 (N_5943,N_4752,N_4830);
xnor U5944 (N_5944,N_4326,N_4597);
and U5945 (N_5945,N_4583,N_4778);
and U5946 (N_5946,N_4529,N_4064);
and U5947 (N_5947,N_4607,N_4763);
or U5948 (N_5948,N_4789,N_4749);
nor U5949 (N_5949,N_4768,N_4100);
and U5950 (N_5950,N_4143,N_4656);
and U5951 (N_5951,N_4471,N_4391);
or U5952 (N_5952,N_4274,N_4539);
xnor U5953 (N_5953,N_4452,N_4086);
or U5954 (N_5954,N_4595,N_4273);
nor U5955 (N_5955,N_4266,N_4237);
xnor U5956 (N_5956,N_4568,N_4469);
and U5957 (N_5957,N_4917,N_4150);
nand U5958 (N_5958,N_4313,N_4000);
or U5959 (N_5959,N_4105,N_4137);
nand U5960 (N_5960,N_4724,N_4898);
and U5961 (N_5961,N_4130,N_4994);
xor U5962 (N_5962,N_4084,N_4961);
nor U5963 (N_5963,N_4443,N_4621);
or U5964 (N_5964,N_4259,N_4372);
nor U5965 (N_5965,N_4825,N_4068);
and U5966 (N_5966,N_4890,N_4749);
nor U5967 (N_5967,N_4152,N_4920);
or U5968 (N_5968,N_4427,N_4066);
nand U5969 (N_5969,N_4395,N_4004);
or U5970 (N_5970,N_4212,N_4819);
and U5971 (N_5971,N_4412,N_4423);
or U5972 (N_5972,N_4210,N_4959);
and U5973 (N_5973,N_4825,N_4208);
and U5974 (N_5974,N_4779,N_4799);
or U5975 (N_5975,N_4868,N_4344);
nand U5976 (N_5976,N_4655,N_4163);
or U5977 (N_5977,N_4276,N_4263);
and U5978 (N_5978,N_4948,N_4630);
and U5979 (N_5979,N_4072,N_4549);
nand U5980 (N_5980,N_4012,N_4767);
and U5981 (N_5981,N_4396,N_4874);
and U5982 (N_5982,N_4086,N_4509);
or U5983 (N_5983,N_4770,N_4353);
and U5984 (N_5984,N_4751,N_4740);
and U5985 (N_5985,N_4637,N_4676);
xor U5986 (N_5986,N_4523,N_4456);
or U5987 (N_5987,N_4270,N_4516);
nor U5988 (N_5988,N_4679,N_4364);
or U5989 (N_5989,N_4541,N_4265);
and U5990 (N_5990,N_4984,N_4497);
nor U5991 (N_5991,N_4616,N_4185);
nand U5992 (N_5992,N_4071,N_4266);
xnor U5993 (N_5993,N_4555,N_4549);
and U5994 (N_5994,N_4561,N_4419);
xnor U5995 (N_5995,N_4894,N_4010);
nand U5996 (N_5996,N_4634,N_4241);
or U5997 (N_5997,N_4617,N_4084);
or U5998 (N_5998,N_4820,N_4403);
xnor U5999 (N_5999,N_4278,N_4617);
nor U6000 (N_6000,N_5802,N_5608);
or U6001 (N_6001,N_5236,N_5685);
and U6002 (N_6002,N_5010,N_5956);
nor U6003 (N_6003,N_5492,N_5564);
or U6004 (N_6004,N_5738,N_5360);
nand U6005 (N_6005,N_5675,N_5044);
nor U6006 (N_6006,N_5633,N_5673);
xor U6007 (N_6007,N_5262,N_5448);
nand U6008 (N_6008,N_5334,N_5298);
nor U6009 (N_6009,N_5772,N_5770);
nand U6010 (N_6010,N_5018,N_5844);
or U6011 (N_6011,N_5367,N_5748);
or U6012 (N_6012,N_5677,N_5246);
xor U6013 (N_6013,N_5648,N_5720);
or U6014 (N_6014,N_5257,N_5346);
nor U6015 (N_6015,N_5701,N_5900);
nor U6016 (N_6016,N_5927,N_5891);
and U6017 (N_6017,N_5531,N_5939);
nand U6018 (N_6018,N_5807,N_5830);
nor U6019 (N_6019,N_5887,N_5949);
or U6020 (N_6020,N_5189,N_5994);
nor U6021 (N_6021,N_5102,N_5694);
nor U6022 (N_6022,N_5328,N_5489);
xor U6023 (N_6023,N_5136,N_5274);
and U6024 (N_6024,N_5307,N_5993);
or U6025 (N_6025,N_5013,N_5631);
or U6026 (N_6026,N_5460,N_5740);
nor U6027 (N_6027,N_5594,N_5568);
nand U6028 (N_6028,N_5170,N_5174);
and U6029 (N_6029,N_5599,N_5221);
nand U6030 (N_6030,N_5666,N_5235);
xnor U6031 (N_6031,N_5829,N_5182);
xnor U6032 (N_6032,N_5764,N_5981);
or U6033 (N_6033,N_5555,N_5906);
xnor U6034 (N_6034,N_5124,N_5946);
xnor U6035 (N_6035,N_5324,N_5687);
nand U6036 (N_6036,N_5790,N_5926);
or U6037 (N_6037,N_5545,N_5569);
or U6038 (N_6038,N_5417,N_5398);
or U6039 (N_6039,N_5483,N_5913);
or U6040 (N_6040,N_5425,N_5924);
or U6041 (N_6041,N_5261,N_5114);
or U6042 (N_6042,N_5281,N_5625);
and U6043 (N_6043,N_5813,N_5305);
xnor U6044 (N_6044,N_5996,N_5245);
or U6045 (N_6045,N_5252,N_5026);
xnor U6046 (N_6046,N_5186,N_5881);
xnor U6047 (N_6047,N_5263,N_5839);
or U6048 (N_6048,N_5300,N_5809);
nand U6049 (N_6049,N_5350,N_5032);
nand U6050 (N_6050,N_5297,N_5513);
nor U6051 (N_6051,N_5356,N_5962);
nand U6052 (N_6052,N_5200,N_5856);
nor U6053 (N_6053,N_5787,N_5724);
nor U6054 (N_6054,N_5179,N_5447);
or U6055 (N_6055,N_5624,N_5269);
or U6056 (N_6056,N_5522,N_5501);
or U6057 (N_6057,N_5659,N_5444);
xor U6058 (N_6058,N_5070,N_5317);
nand U6059 (N_6059,N_5875,N_5636);
nor U6060 (N_6060,N_5537,N_5651);
nand U6061 (N_6061,N_5079,N_5143);
and U6062 (N_6062,N_5185,N_5794);
nor U6063 (N_6063,N_5394,N_5241);
or U6064 (N_6064,N_5231,N_5977);
nand U6065 (N_6065,N_5431,N_5093);
or U6066 (N_6066,N_5818,N_5497);
and U6067 (N_6067,N_5105,N_5155);
nor U6068 (N_6068,N_5979,N_5291);
or U6069 (N_6069,N_5468,N_5602);
and U6070 (N_6070,N_5965,N_5584);
nor U6071 (N_6071,N_5661,N_5744);
and U6072 (N_6072,N_5530,N_5150);
nor U6073 (N_6073,N_5556,N_5288);
and U6074 (N_6074,N_5978,N_5571);
xnor U6075 (N_6075,N_5126,N_5353);
xnor U6076 (N_6076,N_5475,N_5258);
nand U6077 (N_6077,N_5495,N_5583);
nand U6078 (N_6078,N_5162,N_5730);
nor U6079 (N_6079,N_5760,N_5311);
xnor U6080 (N_6080,N_5240,N_5922);
and U6081 (N_6081,N_5299,N_5751);
xor U6082 (N_6082,N_5512,N_5154);
nor U6083 (N_6083,N_5715,N_5959);
xnor U6084 (N_6084,N_5643,N_5723);
xor U6085 (N_6085,N_5777,N_5708);
nand U6086 (N_6086,N_5786,N_5304);
and U6087 (N_6087,N_5826,N_5035);
or U6088 (N_6088,N_5253,N_5341);
and U6089 (N_6089,N_5396,N_5039);
and U6090 (N_6090,N_5464,N_5273);
and U6091 (N_6091,N_5414,N_5438);
xor U6092 (N_6092,N_5050,N_5002);
xor U6093 (N_6093,N_5190,N_5637);
nand U6094 (N_6094,N_5816,N_5115);
or U6095 (N_6095,N_5045,N_5542);
xor U6096 (N_6096,N_5947,N_5628);
or U6097 (N_6097,N_5316,N_5808);
or U6098 (N_6098,N_5422,N_5478);
nor U6099 (N_6099,N_5128,N_5208);
nor U6100 (N_6100,N_5644,N_5423);
or U6101 (N_6101,N_5742,N_5575);
xnor U6102 (N_6102,N_5156,N_5033);
nor U6103 (N_6103,N_5111,N_5178);
and U6104 (N_6104,N_5523,N_5498);
nand U6105 (N_6105,N_5535,N_5340);
nand U6106 (N_6106,N_5401,N_5151);
nand U6107 (N_6107,N_5707,N_5428);
xnor U6108 (N_6108,N_5792,N_5243);
nand U6109 (N_6109,N_5543,N_5137);
xnor U6110 (N_6110,N_5023,N_5799);
xnor U6111 (N_6111,N_5435,N_5558);
xor U6112 (N_6112,N_5488,N_5203);
nor U6113 (N_6113,N_5911,N_5160);
nand U6114 (N_6114,N_5385,N_5862);
xor U6115 (N_6115,N_5477,N_5695);
and U6116 (N_6116,N_5217,N_5219);
nor U6117 (N_6117,N_5713,N_5604);
xnor U6118 (N_6118,N_5060,N_5548);
or U6119 (N_6119,N_5158,N_5017);
and U6120 (N_6120,N_5974,N_5655);
and U6121 (N_6121,N_5019,N_5528);
nand U6122 (N_6122,N_5879,N_5817);
xor U6123 (N_6123,N_5941,N_5597);
nand U6124 (N_6124,N_5653,N_5780);
or U6125 (N_6125,N_5506,N_5667);
nor U6126 (N_6126,N_5074,N_5953);
and U6127 (N_6127,N_5954,N_5987);
and U6128 (N_6128,N_5763,N_5616);
xnor U6129 (N_6129,N_5302,N_5419);
or U6130 (N_6130,N_5333,N_5177);
and U6131 (N_6131,N_5827,N_5952);
xnor U6132 (N_6132,N_5061,N_5592);
nor U6133 (N_6133,N_5199,N_5016);
xnor U6134 (N_6134,N_5502,N_5146);
or U6135 (N_6135,N_5581,N_5226);
nor U6136 (N_6136,N_5679,N_5649);
nand U6137 (N_6137,N_5216,N_5822);
or U6138 (N_6138,N_5593,N_5280);
nand U6139 (N_6139,N_5140,N_5538);
nand U6140 (N_6140,N_5944,N_5097);
nor U6141 (N_6141,N_5073,N_5663);
nand U6142 (N_6142,N_5553,N_5629);
or U6143 (N_6143,N_5138,N_5833);
and U6144 (N_6144,N_5391,N_5860);
xnor U6145 (N_6145,N_5481,N_5938);
nor U6146 (N_6146,N_5450,N_5020);
and U6147 (N_6147,N_5206,N_5493);
nor U6148 (N_6148,N_5968,N_5868);
or U6149 (N_6149,N_5758,N_5218);
nand U6150 (N_6150,N_5194,N_5966);
and U6151 (N_6151,N_5089,N_5410);
nand U6152 (N_6152,N_5165,N_5390);
or U6153 (N_6153,N_5008,N_5539);
nor U6154 (N_6154,N_5198,N_5640);
nand U6155 (N_6155,N_5113,N_5885);
or U6156 (N_6156,N_5296,N_5865);
nand U6157 (N_6157,N_5957,N_5267);
nand U6158 (N_6158,N_5322,N_5042);
xor U6159 (N_6159,N_5612,N_5570);
nor U6160 (N_6160,N_5632,N_5265);
or U6161 (N_6161,N_5840,N_5169);
or U6162 (N_6162,N_5188,N_5015);
nor U6163 (N_6163,N_5842,N_5846);
xnor U6164 (N_6164,N_5825,N_5117);
xor U6165 (N_6165,N_5365,N_5439);
and U6166 (N_6166,N_5755,N_5287);
and U6167 (N_6167,N_5192,N_5167);
xnor U6168 (N_6168,N_5040,N_5903);
nand U6169 (N_6169,N_5164,N_5133);
xnor U6170 (N_6170,N_5387,N_5482);
nand U6171 (N_6171,N_5735,N_5331);
nor U6172 (N_6172,N_5517,N_5187);
and U6173 (N_6173,N_5348,N_5940);
nor U6174 (N_6174,N_5511,N_5769);
nor U6175 (N_6175,N_5585,N_5622);
nand U6176 (N_6176,N_5639,N_5092);
or U6177 (N_6177,N_5344,N_5992);
nand U6178 (N_6178,N_5270,N_5472);
or U6179 (N_6179,N_5849,N_5430);
nor U6180 (N_6180,N_5916,N_5456);
nor U6181 (N_6181,N_5275,N_5980);
or U6182 (N_6182,N_5699,N_5732);
or U6183 (N_6183,N_5765,N_5323);
and U6184 (N_6184,N_5931,N_5239);
nor U6185 (N_6185,N_5209,N_5054);
nand U6186 (N_6186,N_5999,N_5918);
nor U6187 (N_6187,N_5036,N_5393);
nor U6188 (N_6188,N_5437,N_5686);
xnor U6189 (N_6189,N_5181,N_5180);
or U6190 (N_6190,N_5249,N_5610);
nor U6191 (N_6191,N_5355,N_5507);
or U6192 (N_6192,N_5869,N_5434);
or U6193 (N_6193,N_5034,N_5386);
nor U6194 (N_6194,N_5682,N_5122);
or U6195 (N_6195,N_5768,N_5873);
and U6196 (N_6196,N_5746,N_5726);
nor U6197 (N_6197,N_5620,N_5131);
nand U6198 (N_6198,N_5232,N_5909);
xor U6199 (N_6199,N_5351,N_5657);
xnor U6200 (N_6200,N_5948,N_5576);
nand U6201 (N_6201,N_5471,N_5496);
xnor U6202 (N_6202,N_5046,N_5697);
nand U6203 (N_6203,N_5429,N_5526);
and U6204 (N_6204,N_5835,N_5377);
and U6205 (N_6205,N_5374,N_5251);
nor U6206 (N_6206,N_5009,N_5831);
and U6207 (N_6207,N_5282,N_5867);
nor U6208 (N_6208,N_5793,N_5025);
xor U6209 (N_6209,N_5491,N_5562);
or U6210 (N_6210,N_5857,N_5458);
or U6211 (N_6211,N_5065,N_5470);
nand U6212 (N_6212,N_5985,N_5255);
and U6213 (N_6213,N_5806,N_5621);
and U6214 (N_6214,N_5301,N_5877);
nand U6215 (N_6215,N_5838,N_5905);
nor U6216 (N_6216,N_5370,N_5658);
xor U6217 (N_6217,N_5843,N_5915);
nand U6218 (N_6218,N_5883,N_5424);
xnor U6219 (N_6219,N_5889,N_5567);
nand U6220 (N_6220,N_5784,N_5656);
nand U6221 (N_6221,N_5103,N_5795);
or U6222 (N_6222,N_5991,N_5823);
and U6223 (N_6223,N_5084,N_5413);
or U6224 (N_6224,N_5782,N_5973);
or U6225 (N_6225,N_5005,N_5284);
nand U6226 (N_6226,N_5728,N_5392);
nor U6227 (N_6227,N_5847,N_5509);
xor U6228 (N_6228,N_5369,N_5309);
or U6229 (N_6229,N_5554,N_5573);
and U6230 (N_6230,N_5157,N_5363);
nand U6231 (N_6231,N_5774,N_5762);
and U6232 (N_6232,N_5778,N_5233);
nor U6233 (N_6233,N_5731,N_5250);
and U6234 (N_6234,N_5088,N_5880);
xor U6235 (N_6235,N_5967,N_5714);
nor U6236 (N_6236,N_5866,N_5318);
xnor U6237 (N_6237,N_5963,N_5988);
nor U6238 (N_6238,N_5698,N_5173);
nor U6239 (N_6239,N_5547,N_5395);
nand U6240 (N_6240,N_5004,N_5135);
nor U6241 (N_6241,N_5615,N_5626);
or U6242 (N_6242,N_5971,N_5098);
xor U6243 (N_6243,N_5163,N_5238);
nor U6244 (N_6244,N_5404,N_5814);
nand U6245 (N_6245,N_5120,N_5453);
or U6246 (N_6246,N_5619,N_5082);
and U6247 (N_6247,N_5466,N_5202);
or U6248 (N_6248,N_5759,N_5159);
and U6249 (N_6249,N_5645,N_5166);
and U6250 (N_6250,N_5750,N_5696);
nor U6251 (N_6251,N_5407,N_5196);
nand U6252 (N_6252,N_5406,N_5935);
xor U6253 (N_6253,N_5021,N_5094);
or U6254 (N_6254,N_5609,N_5692);
or U6255 (N_6255,N_5729,N_5705);
nor U6256 (N_6256,N_5733,N_5719);
xnor U6257 (N_6257,N_5925,N_5244);
nor U6258 (N_6258,N_5349,N_5864);
or U6259 (N_6259,N_5718,N_5402);
and U6260 (N_6260,N_5161,N_5669);
xnor U6261 (N_6261,N_5912,N_5734);
nand U6262 (N_6262,N_5123,N_5230);
xor U6263 (N_6263,N_5215,N_5725);
xnor U6264 (N_6264,N_5749,N_5929);
nor U6265 (N_6265,N_5071,N_5798);
nor U6266 (N_6266,N_5047,N_5711);
and U6267 (N_6267,N_5572,N_5358);
and U6268 (N_6268,N_5898,N_5557);
or U6269 (N_6269,N_5508,N_5076);
nand U6270 (N_6270,N_5660,N_5641);
nor U6271 (N_6271,N_5003,N_5066);
xor U6272 (N_6272,N_5736,N_5934);
xnor U6273 (N_6273,N_5559,N_5998);
and U6274 (N_6274,N_5381,N_5872);
nor U6275 (N_6275,N_5320,N_5853);
or U6276 (N_6276,N_5290,N_5797);
xnor U6277 (N_6277,N_5459,N_5433);
or U6278 (N_6278,N_5201,N_5152);
nor U6279 (N_6279,N_5613,N_5279);
and U6280 (N_6280,N_5081,N_5229);
or U6281 (N_6281,N_5688,N_5519);
and U6282 (N_6282,N_5022,N_5693);
or U6283 (N_6283,N_5310,N_5306);
or U6284 (N_6284,N_5969,N_5684);
nor U6285 (N_6285,N_5532,N_5587);
nand U6286 (N_6286,N_5607,N_5756);
xnor U6287 (N_6287,N_5197,N_5056);
nor U6288 (N_6288,N_5006,N_5789);
and U6289 (N_6289,N_5476,N_5247);
nor U6290 (N_6290,N_5551,N_5212);
nor U6291 (N_6291,N_5141,N_5691);
and U6292 (N_6292,N_5266,N_5104);
or U6293 (N_6293,N_5264,N_5504);
nor U6294 (N_6294,N_5525,N_5646);
and U6295 (N_6295,N_5462,N_5888);
and U6296 (N_6296,N_5960,N_5380);
and U6297 (N_6297,N_5937,N_5024);
xnor U6298 (N_6298,N_5500,N_5767);
or U6299 (N_6299,N_5709,N_5982);
nor U6300 (N_6300,N_5172,N_5440);
or U6301 (N_6301,N_5063,N_5541);
and U6302 (N_6302,N_5662,N_5222);
nor U6303 (N_6303,N_5330,N_5144);
or U6304 (N_6304,N_5086,N_5283);
or U6305 (N_6305,N_5514,N_5776);
nor U6306 (N_6306,N_5052,N_5921);
xnor U6307 (N_6307,N_5781,N_5049);
and U6308 (N_6308,N_5832,N_5038);
or U6309 (N_6309,N_5409,N_5565);
or U6310 (N_6310,N_5108,N_5127);
nand U6311 (N_6311,N_5067,N_5361);
xnor U6312 (N_6312,N_5227,N_5213);
or U6313 (N_6313,N_5053,N_5970);
nor U6314 (N_6314,N_5800,N_5454);
and U6315 (N_6315,N_5618,N_5801);
or U6316 (N_6316,N_5077,N_5383);
nor U6317 (N_6317,N_5455,N_5722);
nand U6318 (N_6318,N_5225,N_5145);
and U6319 (N_6319,N_5582,N_5321);
nor U6320 (N_6320,N_5384,N_5418);
nand U6321 (N_6321,N_5861,N_5256);
nand U6322 (N_6322,N_5596,N_5958);
nor U6323 (N_6323,N_5577,N_5175);
nor U6324 (N_6324,N_5234,N_5884);
nor U6325 (N_6325,N_5205,N_5057);
xnor U6326 (N_6326,N_5183,N_5739);
nand U6327 (N_6327,N_5214,N_5886);
xnor U6328 (N_6328,N_5055,N_5623);
and U6329 (N_6329,N_5757,N_5589);
nor U6330 (N_6330,N_5805,N_5578);
nand U6331 (N_6331,N_5271,N_5095);
and U6332 (N_6332,N_5943,N_5518);
xor U6333 (N_6333,N_5503,N_5119);
and U6334 (N_6334,N_5819,N_5012);
xnor U6335 (N_6335,N_5896,N_5107);
nand U6336 (N_6336,N_5529,N_5579);
or U6337 (N_6337,N_5964,N_5989);
nor U6338 (N_6338,N_5520,N_5210);
xor U6339 (N_6339,N_5870,N_5836);
and U6340 (N_6340,N_5563,N_5371);
or U6341 (N_6341,N_5876,N_5654);
and U6342 (N_6342,N_5951,N_5457);
or U6343 (N_6343,N_5902,N_5540);
nor U6344 (N_6344,N_5706,N_5485);
xor U6345 (N_6345,N_5907,N_5863);
or U6346 (N_6346,N_5552,N_5950);
nor U6347 (N_6347,N_5325,N_5373);
nor U6348 (N_6348,N_5783,N_5441);
and U6349 (N_6349,N_5388,N_5779);
xnor U6350 (N_6350,N_5101,N_5260);
xor U6351 (N_6351,N_5990,N_5408);
xor U6352 (N_6352,N_5588,N_5364);
nor U6353 (N_6353,N_5338,N_5352);
nand U6354 (N_6354,N_5224,N_5617);
nor U6355 (N_6355,N_5339,N_5294);
and U6356 (N_6356,N_5195,N_5112);
nand U6357 (N_6357,N_5499,N_5897);
or U6358 (N_6358,N_5841,N_5812);
or U6359 (N_6359,N_5908,N_5892);
nand U6360 (N_6360,N_5796,N_5465);
nand U6361 (N_6361,N_5930,N_5854);
nor U6362 (N_6362,N_5375,N_5041);
and U6363 (N_6363,N_5191,N_5343);
and U6364 (N_6364,N_5727,N_5319);
nor U6365 (N_6365,N_5521,N_5118);
or U6366 (N_6366,N_5277,N_5399);
and U6367 (N_6367,N_5936,N_5064);
nand U6368 (N_6368,N_5248,N_5403);
nor U6369 (N_6369,N_5449,N_5139);
or U6370 (N_6370,N_5810,N_5920);
nor U6371 (N_6371,N_5027,N_5125);
xnor U6372 (N_6372,N_5761,N_5741);
and U6373 (N_6373,N_5536,N_5359);
and U6374 (N_6374,N_5893,N_5834);
xor U6375 (N_6375,N_5972,N_5129);
or U6376 (N_6376,N_5516,N_5773);
nand U6377 (N_6377,N_5515,N_5904);
nor U6378 (N_6378,N_5031,N_5347);
nor U6379 (N_6379,N_5204,N_5171);
nor U6380 (N_6380,N_5544,N_5919);
or U6381 (N_6381,N_5580,N_5775);
xnor U6382 (N_6382,N_5614,N_5932);
and U6383 (N_6383,N_5745,N_5852);
xor U6384 (N_6384,N_5335,N_5001);
xnor U6385 (N_6385,N_5804,N_5362);
nor U6386 (N_6386,N_5574,N_5443);
nor U6387 (N_6387,N_5803,N_5600);
or U6388 (N_6388,N_5671,N_5176);
nor U6389 (N_6389,N_5630,N_5882);
and U6390 (N_6390,N_5480,N_5820);
nand U6391 (N_6391,N_5986,N_5037);
nand U6392 (N_6392,N_5590,N_5858);
nand U6393 (N_6393,N_5085,N_5678);
or U6394 (N_6394,N_5132,N_5389);
nand U6395 (N_6395,N_5116,N_5068);
nand U6396 (N_6396,N_5223,N_5894);
and U6397 (N_6397,N_5442,N_5411);
and U6398 (N_6398,N_5228,N_5487);
xor U6399 (N_6399,N_5717,N_5368);
nand U6400 (N_6400,N_5753,N_5043);
nand U6401 (N_6401,N_5665,N_5961);
and U6402 (N_6402,N_5148,N_5672);
or U6403 (N_6403,N_5376,N_5561);
xor U6404 (N_6404,N_5083,N_5933);
nand U6405 (N_6405,N_5327,N_5062);
nor U6406 (N_6406,N_5011,N_5534);
nand U6407 (N_6407,N_5664,N_5848);
nand U6408 (N_6408,N_5785,N_5704);
nor U6409 (N_6409,N_5550,N_5895);
xor U6410 (N_6410,N_5689,N_5072);
and U6411 (N_6411,N_5451,N_5976);
or U6412 (N_6412,N_5674,N_5329);
or U6413 (N_6413,N_5436,N_5153);
and U6414 (N_6414,N_5586,N_5087);
nor U6415 (N_6415,N_5000,N_5983);
and U6416 (N_6416,N_5942,N_5293);
and U6417 (N_6417,N_5560,N_5754);
nand U6418 (N_6418,N_5121,N_5670);
nor U6419 (N_6419,N_5242,N_5168);
xor U6420 (N_6420,N_5193,N_5527);
and U6421 (N_6421,N_5130,N_5710);
or U6422 (N_6422,N_5995,N_5851);
xor U6423 (N_6423,N_5308,N_5075);
xnor U6424 (N_6424,N_5743,N_5254);
or U6425 (N_6425,N_5627,N_5286);
xnor U6426 (N_6426,N_5533,N_5652);
nor U6427 (N_6427,N_5871,N_5285);
and U6428 (N_6428,N_5314,N_5791);
nor U6429 (N_6429,N_5859,N_5313);
and U6430 (N_6430,N_5357,N_5345);
nand U6431 (N_6431,N_5716,N_5681);
xnor U6432 (N_6432,N_5473,N_5815);
xnor U6433 (N_6433,N_5220,N_5703);
xnor U6434 (N_6434,N_5766,N_5700);
or U6435 (N_6435,N_5690,N_5326);
or U6436 (N_6436,N_5494,N_5788);
nand U6437 (N_6437,N_5917,N_5342);
nor U6438 (N_6438,N_5091,N_5014);
xnor U6439 (N_6439,N_5474,N_5315);
and U6440 (N_6440,N_5821,N_5426);
xor U6441 (N_6441,N_5379,N_5292);
nor U6442 (N_6442,N_5997,N_5650);
xor U6443 (N_6443,N_5611,N_5874);
or U6444 (N_6444,N_5452,N_5490);
xnor U6445 (N_6445,N_5099,N_5303);
nand U6446 (N_6446,N_5461,N_5747);
or U6447 (N_6447,N_5901,N_5680);
nand U6448 (N_6448,N_5336,N_5445);
nand U6449 (N_6449,N_5484,N_5211);
or U6450 (N_6450,N_5090,N_5184);
or U6451 (N_6451,N_5855,N_5914);
xor U6452 (N_6452,N_5059,N_5400);
and U6453 (N_6453,N_5824,N_5147);
and U6454 (N_6454,N_5149,N_5421);
nand U6455 (N_6455,N_5603,N_5598);
or U6456 (N_6456,N_5635,N_5427);
nand U6457 (N_6457,N_5134,N_5647);
and U6458 (N_6458,N_5524,N_5259);
and U6459 (N_6459,N_5432,N_5007);
or U6460 (N_6460,N_5605,N_5486);
nand U6461 (N_6461,N_5899,N_5467);
or U6462 (N_6462,N_5676,N_5928);
or U6463 (N_6463,N_5668,N_5366);
and U6464 (N_6464,N_5058,N_5712);
nand U6465 (N_6465,N_5721,N_5268);
nand U6466 (N_6466,N_5811,N_5463);
or U6467 (N_6467,N_5096,N_5415);
and U6468 (N_6468,N_5837,N_5510);
and U6469 (N_6469,N_5354,N_5028);
nand U6470 (N_6470,N_5412,N_5566);
or U6471 (N_6471,N_5595,N_5276);
and U6472 (N_6472,N_5080,N_5078);
or U6473 (N_6473,N_5278,N_5048);
nand U6474 (N_6474,N_5142,N_5029);
nor U6475 (N_6475,N_5638,N_5642);
nor U6476 (N_6476,N_5601,N_5207);
nand U6477 (N_6477,N_5984,N_5069);
nor U6478 (N_6478,N_5030,N_5945);
or U6479 (N_6479,N_5109,N_5752);
xor U6480 (N_6480,N_5416,N_5591);
xor U6481 (N_6481,N_5850,N_5332);
nand U6482 (N_6482,N_5737,N_5420);
or U6483 (N_6483,N_5469,N_5100);
or U6484 (N_6484,N_5312,N_5771);
and U6485 (N_6485,N_5378,N_5923);
and U6486 (N_6486,N_5337,N_5106);
xnor U6487 (N_6487,N_5505,N_5683);
and U6488 (N_6488,N_5397,N_5479);
nand U6489 (N_6489,N_5237,N_5890);
and U6490 (N_6490,N_5702,N_5295);
nand U6491 (N_6491,N_5634,N_5289);
xor U6492 (N_6492,N_5382,N_5546);
and U6493 (N_6493,N_5372,N_5549);
xor U6494 (N_6494,N_5110,N_5606);
nor U6495 (N_6495,N_5975,N_5955);
and U6496 (N_6496,N_5446,N_5910);
xnor U6497 (N_6497,N_5845,N_5405);
xor U6498 (N_6498,N_5828,N_5878);
nor U6499 (N_6499,N_5051,N_5272);
nand U6500 (N_6500,N_5653,N_5758);
nor U6501 (N_6501,N_5490,N_5256);
and U6502 (N_6502,N_5576,N_5956);
or U6503 (N_6503,N_5073,N_5940);
xor U6504 (N_6504,N_5085,N_5138);
nor U6505 (N_6505,N_5864,N_5381);
or U6506 (N_6506,N_5143,N_5057);
nor U6507 (N_6507,N_5895,N_5670);
nand U6508 (N_6508,N_5746,N_5477);
xor U6509 (N_6509,N_5782,N_5859);
or U6510 (N_6510,N_5550,N_5734);
or U6511 (N_6511,N_5641,N_5913);
nor U6512 (N_6512,N_5151,N_5266);
and U6513 (N_6513,N_5229,N_5730);
nor U6514 (N_6514,N_5799,N_5295);
nand U6515 (N_6515,N_5768,N_5761);
nand U6516 (N_6516,N_5477,N_5537);
nand U6517 (N_6517,N_5776,N_5979);
or U6518 (N_6518,N_5455,N_5440);
or U6519 (N_6519,N_5686,N_5824);
and U6520 (N_6520,N_5545,N_5941);
and U6521 (N_6521,N_5375,N_5297);
xnor U6522 (N_6522,N_5132,N_5071);
nand U6523 (N_6523,N_5375,N_5464);
xor U6524 (N_6524,N_5922,N_5182);
nand U6525 (N_6525,N_5481,N_5451);
or U6526 (N_6526,N_5278,N_5243);
nand U6527 (N_6527,N_5775,N_5360);
nor U6528 (N_6528,N_5186,N_5488);
or U6529 (N_6529,N_5160,N_5353);
nand U6530 (N_6530,N_5322,N_5898);
nor U6531 (N_6531,N_5547,N_5079);
xor U6532 (N_6532,N_5909,N_5679);
nand U6533 (N_6533,N_5413,N_5735);
xor U6534 (N_6534,N_5581,N_5336);
nand U6535 (N_6535,N_5108,N_5174);
and U6536 (N_6536,N_5298,N_5588);
or U6537 (N_6537,N_5404,N_5872);
xor U6538 (N_6538,N_5836,N_5213);
nor U6539 (N_6539,N_5344,N_5811);
and U6540 (N_6540,N_5332,N_5219);
nor U6541 (N_6541,N_5510,N_5244);
nor U6542 (N_6542,N_5093,N_5619);
nor U6543 (N_6543,N_5136,N_5898);
nor U6544 (N_6544,N_5096,N_5948);
nand U6545 (N_6545,N_5085,N_5258);
or U6546 (N_6546,N_5107,N_5387);
or U6547 (N_6547,N_5095,N_5398);
xnor U6548 (N_6548,N_5017,N_5678);
nor U6549 (N_6549,N_5948,N_5309);
nor U6550 (N_6550,N_5563,N_5876);
nand U6551 (N_6551,N_5064,N_5033);
and U6552 (N_6552,N_5309,N_5653);
nand U6553 (N_6553,N_5201,N_5951);
xnor U6554 (N_6554,N_5211,N_5942);
and U6555 (N_6555,N_5469,N_5754);
xnor U6556 (N_6556,N_5452,N_5025);
nand U6557 (N_6557,N_5793,N_5420);
nor U6558 (N_6558,N_5802,N_5992);
nand U6559 (N_6559,N_5224,N_5893);
and U6560 (N_6560,N_5586,N_5657);
nand U6561 (N_6561,N_5903,N_5541);
xnor U6562 (N_6562,N_5221,N_5956);
nor U6563 (N_6563,N_5878,N_5677);
or U6564 (N_6564,N_5162,N_5608);
nor U6565 (N_6565,N_5637,N_5062);
xor U6566 (N_6566,N_5052,N_5912);
nand U6567 (N_6567,N_5341,N_5140);
xor U6568 (N_6568,N_5689,N_5473);
and U6569 (N_6569,N_5478,N_5282);
nand U6570 (N_6570,N_5259,N_5690);
nor U6571 (N_6571,N_5493,N_5845);
or U6572 (N_6572,N_5006,N_5507);
or U6573 (N_6573,N_5315,N_5662);
xnor U6574 (N_6574,N_5551,N_5919);
or U6575 (N_6575,N_5908,N_5443);
xnor U6576 (N_6576,N_5623,N_5019);
xnor U6577 (N_6577,N_5008,N_5468);
or U6578 (N_6578,N_5808,N_5353);
or U6579 (N_6579,N_5462,N_5793);
and U6580 (N_6580,N_5633,N_5909);
nor U6581 (N_6581,N_5078,N_5236);
xor U6582 (N_6582,N_5604,N_5623);
xor U6583 (N_6583,N_5252,N_5269);
nand U6584 (N_6584,N_5881,N_5374);
and U6585 (N_6585,N_5734,N_5501);
nand U6586 (N_6586,N_5637,N_5371);
nor U6587 (N_6587,N_5179,N_5893);
or U6588 (N_6588,N_5098,N_5297);
and U6589 (N_6589,N_5093,N_5045);
nand U6590 (N_6590,N_5191,N_5742);
nand U6591 (N_6591,N_5087,N_5751);
xnor U6592 (N_6592,N_5362,N_5063);
or U6593 (N_6593,N_5018,N_5498);
and U6594 (N_6594,N_5214,N_5582);
and U6595 (N_6595,N_5850,N_5112);
nand U6596 (N_6596,N_5217,N_5573);
nand U6597 (N_6597,N_5191,N_5474);
xor U6598 (N_6598,N_5903,N_5127);
and U6599 (N_6599,N_5189,N_5438);
and U6600 (N_6600,N_5967,N_5812);
or U6601 (N_6601,N_5095,N_5039);
or U6602 (N_6602,N_5162,N_5260);
or U6603 (N_6603,N_5562,N_5383);
and U6604 (N_6604,N_5481,N_5631);
nor U6605 (N_6605,N_5211,N_5625);
or U6606 (N_6606,N_5207,N_5830);
nor U6607 (N_6607,N_5225,N_5223);
nor U6608 (N_6608,N_5890,N_5509);
xnor U6609 (N_6609,N_5318,N_5854);
nor U6610 (N_6610,N_5393,N_5585);
and U6611 (N_6611,N_5435,N_5453);
or U6612 (N_6612,N_5567,N_5205);
nand U6613 (N_6613,N_5478,N_5035);
and U6614 (N_6614,N_5917,N_5767);
nor U6615 (N_6615,N_5566,N_5266);
nor U6616 (N_6616,N_5086,N_5706);
xnor U6617 (N_6617,N_5298,N_5628);
nand U6618 (N_6618,N_5847,N_5159);
xnor U6619 (N_6619,N_5050,N_5821);
and U6620 (N_6620,N_5564,N_5225);
nor U6621 (N_6621,N_5296,N_5533);
or U6622 (N_6622,N_5172,N_5002);
nor U6623 (N_6623,N_5694,N_5386);
nand U6624 (N_6624,N_5281,N_5029);
or U6625 (N_6625,N_5929,N_5412);
nand U6626 (N_6626,N_5121,N_5047);
nor U6627 (N_6627,N_5174,N_5332);
nor U6628 (N_6628,N_5860,N_5096);
nor U6629 (N_6629,N_5966,N_5543);
xnor U6630 (N_6630,N_5054,N_5775);
xnor U6631 (N_6631,N_5638,N_5853);
and U6632 (N_6632,N_5335,N_5667);
nand U6633 (N_6633,N_5239,N_5326);
nand U6634 (N_6634,N_5089,N_5325);
nand U6635 (N_6635,N_5086,N_5237);
nor U6636 (N_6636,N_5368,N_5469);
xor U6637 (N_6637,N_5046,N_5431);
or U6638 (N_6638,N_5413,N_5770);
xnor U6639 (N_6639,N_5888,N_5306);
nand U6640 (N_6640,N_5707,N_5161);
or U6641 (N_6641,N_5153,N_5043);
or U6642 (N_6642,N_5206,N_5846);
or U6643 (N_6643,N_5377,N_5759);
and U6644 (N_6644,N_5450,N_5976);
nand U6645 (N_6645,N_5844,N_5520);
or U6646 (N_6646,N_5426,N_5454);
and U6647 (N_6647,N_5999,N_5160);
nand U6648 (N_6648,N_5771,N_5310);
or U6649 (N_6649,N_5164,N_5093);
nand U6650 (N_6650,N_5793,N_5845);
and U6651 (N_6651,N_5788,N_5221);
or U6652 (N_6652,N_5857,N_5355);
nor U6653 (N_6653,N_5005,N_5133);
and U6654 (N_6654,N_5004,N_5095);
and U6655 (N_6655,N_5036,N_5070);
xnor U6656 (N_6656,N_5213,N_5396);
xnor U6657 (N_6657,N_5115,N_5612);
or U6658 (N_6658,N_5114,N_5441);
or U6659 (N_6659,N_5033,N_5190);
and U6660 (N_6660,N_5868,N_5515);
nand U6661 (N_6661,N_5139,N_5181);
xnor U6662 (N_6662,N_5823,N_5090);
or U6663 (N_6663,N_5386,N_5303);
and U6664 (N_6664,N_5363,N_5687);
nor U6665 (N_6665,N_5903,N_5734);
nand U6666 (N_6666,N_5091,N_5984);
and U6667 (N_6667,N_5190,N_5697);
xnor U6668 (N_6668,N_5563,N_5465);
or U6669 (N_6669,N_5584,N_5885);
nor U6670 (N_6670,N_5104,N_5911);
and U6671 (N_6671,N_5144,N_5480);
nand U6672 (N_6672,N_5425,N_5829);
nor U6673 (N_6673,N_5982,N_5768);
nor U6674 (N_6674,N_5462,N_5703);
and U6675 (N_6675,N_5344,N_5710);
or U6676 (N_6676,N_5415,N_5007);
xor U6677 (N_6677,N_5530,N_5549);
nand U6678 (N_6678,N_5065,N_5289);
nand U6679 (N_6679,N_5148,N_5311);
or U6680 (N_6680,N_5097,N_5892);
or U6681 (N_6681,N_5606,N_5225);
nand U6682 (N_6682,N_5903,N_5431);
nand U6683 (N_6683,N_5690,N_5951);
xnor U6684 (N_6684,N_5416,N_5044);
or U6685 (N_6685,N_5224,N_5868);
and U6686 (N_6686,N_5347,N_5646);
xor U6687 (N_6687,N_5211,N_5190);
or U6688 (N_6688,N_5183,N_5175);
xnor U6689 (N_6689,N_5398,N_5855);
xor U6690 (N_6690,N_5188,N_5676);
and U6691 (N_6691,N_5225,N_5464);
nor U6692 (N_6692,N_5141,N_5766);
xor U6693 (N_6693,N_5713,N_5821);
nor U6694 (N_6694,N_5067,N_5376);
or U6695 (N_6695,N_5067,N_5801);
and U6696 (N_6696,N_5348,N_5038);
xor U6697 (N_6697,N_5188,N_5791);
xnor U6698 (N_6698,N_5680,N_5278);
xor U6699 (N_6699,N_5805,N_5610);
nor U6700 (N_6700,N_5792,N_5452);
nor U6701 (N_6701,N_5047,N_5332);
or U6702 (N_6702,N_5483,N_5648);
nand U6703 (N_6703,N_5502,N_5560);
nor U6704 (N_6704,N_5426,N_5608);
nor U6705 (N_6705,N_5215,N_5974);
nor U6706 (N_6706,N_5484,N_5848);
nand U6707 (N_6707,N_5823,N_5038);
nand U6708 (N_6708,N_5525,N_5124);
and U6709 (N_6709,N_5490,N_5787);
or U6710 (N_6710,N_5335,N_5505);
and U6711 (N_6711,N_5070,N_5267);
nand U6712 (N_6712,N_5281,N_5810);
nand U6713 (N_6713,N_5400,N_5056);
nand U6714 (N_6714,N_5847,N_5421);
nand U6715 (N_6715,N_5058,N_5323);
nand U6716 (N_6716,N_5952,N_5791);
nor U6717 (N_6717,N_5341,N_5502);
and U6718 (N_6718,N_5440,N_5299);
nor U6719 (N_6719,N_5070,N_5804);
xnor U6720 (N_6720,N_5730,N_5893);
nor U6721 (N_6721,N_5635,N_5303);
xnor U6722 (N_6722,N_5402,N_5801);
nand U6723 (N_6723,N_5778,N_5128);
nor U6724 (N_6724,N_5329,N_5280);
and U6725 (N_6725,N_5253,N_5923);
or U6726 (N_6726,N_5738,N_5112);
and U6727 (N_6727,N_5657,N_5557);
nor U6728 (N_6728,N_5598,N_5145);
nor U6729 (N_6729,N_5584,N_5629);
xor U6730 (N_6730,N_5880,N_5099);
nor U6731 (N_6731,N_5265,N_5975);
or U6732 (N_6732,N_5465,N_5618);
or U6733 (N_6733,N_5674,N_5829);
and U6734 (N_6734,N_5698,N_5449);
or U6735 (N_6735,N_5005,N_5811);
and U6736 (N_6736,N_5944,N_5270);
and U6737 (N_6737,N_5231,N_5352);
nand U6738 (N_6738,N_5438,N_5505);
nor U6739 (N_6739,N_5100,N_5444);
nor U6740 (N_6740,N_5949,N_5793);
xnor U6741 (N_6741,N_5171,N_5435);
xnor U6742 (N_6742,N_5026,N_5343);
or U6743 (N_6743,N_5550,N_5620);
or U6744 (N_6744,N_5850,N_5225);
or U6745 (N_6745,N_5201,N_5271);
and U6746 (N_6746,N_5779,N_5412);
and U6747 (N_6747,N_5614,N_5044);
and U6748 (N_6748,N_5441,N_5913);
or U6749 (N_6749,N_5102,N_5504);
nand U6750 (N_6750,N_5111,N_5353);
or U6751 (N_6751,N_5859,N_5429);
or U6752 (N_6752,N_5849,N_5326);
or U6753 (N_6753,N_5019,N_5702);
or U6754 (N_6754,N_5141,N_5493);
nor U6755 (N_6755,N_5189,N_5579);
nand U6756 (N_6756,N_5855,N_5471);
or U6757 (N_6757,N_5064,N_5945);
and U6758 (N_6758,N_5880,N_5933);
nand U6759 (N_6759,N_5188,N_5567);
xor U6760 (N_6760,N_5154,N_5290);
nor U6761 (N_6761,N_5301,N_5065);
and U6762 (N_6762,N_5410,N_5604);
xor U6763 (N_6763,N_5625,N_5869);
xnor U6764 (N_6764,N_5910,N_5409);
nand U6765 (N_6765,N_5797,N_5615);
nand U6766 (N_6766,N_5280,N_5263);
and U6767 (N_6767,N_5813,N_5115);
and U6768 (N_6768,N_5221,N_5266);
xnor U6769 (N_6769,N_5254,N_5461);
xor U6770 (N_6770,N_5100,N_5774);
and U6771 (N_6771,N_5682,N_5277);
xnor U6772 (N_6772,N_5049,N_5454);
xor U6773 (N_6773,N_5683,N_5093);
xor U6774 (N_6774,N_5182,N_5760);
nand U6775 (N_6775,N_5771,N_5516);
or U6776 (N_6776,N_5963,N_5088);
nand U6777 (N_6777,N_5008,N_5018);
nor U6778 (N_6778,N_5577,N_5273);
and U6779 (N_6779,N_5664,N_5528);
xor U6780 (N_6780,N_5701,N_5048);
or U6781 (N_6781,N_5769,N_5098);
nand U6782 (N_6782,N_5544,N_5752);
nand U6783 (N_6783,N_5301,N_5659);
or U6784 (N_6784,N_5775,N_5762);
or U6785 (N_6785,N_5496,N_5266);
or U6786 (N_6786,N_5581,N_5015);
and U6787 (N_6787,N_5503,N_5282);
or U6788 (N_6788,N_5380,N_5663);
nor U6789 (N_6789,N_5894,N_5488);
nor U6790 (N_6790,N_5714,N_5888);
nor U6791 (N_6791,N_5245,N_5698);
xnor U6792 (N_6792,N_5833,N_5618);
and U6793 (N_6793,N_5822,N_5946);
and U6794 (N_6794,N_5076,N_5935);
nand U6795 (N_6795,N_5672,N_5323);
and U6796 (N_6796,N_5457,N_5601);
nor U6797 (N_6797,N_5820,N_5963);
xnor U6798 (N_6798,N_5882,N_5362);
xnor U6799 (N_6799,N_5391,N_5977);
nand U6800 (N_6800,N_5726,N_5650);
xor U6801 (N_6801,N_5667,N_5440);
nand U6802 (N_6802,N_5428,N_5790);
and U6803 (N_6803,N_5300,N_5247);
nor U6804 (N_6804,N_5388,N_5800);
or U6805 (N_6805,N_5114,N_5757);
and U6806 (N_6806,N_5773,N_5811);
and U6807 (N_6807,N_5701,N_5901);
nor U6808 (N_6808,N_5925,N_5561);
xor U6809 (N_6809,N_5987,N_5115);
and U6810 (N_6810,N_5381,N_5389);
or U6811 (N_6811,N_5413,N_5570);
xnor U6812 (N_6812,N_5849,N_5954);
xnor U6813 (N_6813,N_5346,N_5350);
and U6814 (N_6814,N_5662,N_5524);
or U6815 (N_6815,N_5389,N_5393);
nand U6816 (N_6816,N_5718,N_5394);
xnor U6817 (N_6817,N_5156,N_5106);
nand U6818 (N_6818,N_5999,N_5577);
nor U6819 (N_6819,N_5072,N_5961);
or U6820 (N_6820,N_5143,N_5190);
xor U6821 (N_6821,N_5256,N_5244);
nand U6822 (N_6822,N_5938,N_5066);
and U6823 (N_6823,N_5776,N_5886);
or U6824 (N_6824,N_5371,N_5308);
nor U6825 (N_6825,N_5667,N_5007);
nor U6826 (N_6826,N_5433,N_5280);
and U6827 (N_6827,N_5277,N_5893);
nor U6828 (N_6828,N_5142,N_5801);
nor U6829 (N_6829,N_5165,N_5180);
nor U6830 (N_6830,N_5636,N_5038);
and U6831 (N_6831,N_5588,N_5552);
or U6832 (N_6832,N_5787,N_5531);
nor U6833 (N_6833,N_5009,N_5930);
or U6834 (N_6834,N_5140,N_5167);
nand U6835 (N_6835,N_5122,N_5613);
xnor U6836 (N_6836,N_5360,N_5322);
xor U6837 (N_6837,N_5578,N_5140);
xnor U6838 (N_6838,N_5229,N_5166);
nand U6839 (N_6839,N_5385,N_5111);
and U6840 (N_6840,N_5485,N_5156);
or U6841 (N_6841,N_5282,N_5584);
nand U6842 (N_6842,N_5907,N_5114);
xor U6843 (N_6843,N_5872,N_5064);
xor U6844 (N_6844,N_5803,N_5083);
or U6845 (N_6845,N_5680,N_5084);
nor U6846 (N_6846,N_5696,N_5350);
and U6847 (N_6847,N_5696,N_5192);
nand U6848 (N_6848,N_5960,N_5470);
nand U6849 (N_6849,N_5883,N_5447);
nor U6850 (N_6850,N_5315,N_5924);
nand U6851 (N_6851,N_5521,N_5247);
xor U6852 (N_6852,N_5911,N_5147);
xnor U6853 (N_6853,N_5118,N_5381);
nor U6854 (N_6854,N_5519,N_5704);
or U6855 (N_6855,N_5571,N_5914);
or U6856 (N_6856,N_5985,N_5855);
xnor U6857 (N_6857,N_5774,N_5293);
nor U6858 (N_6858,N_5424,N_5467);
nor U6859 (N_6859,N_5752,N_5209);
nand U6860 (N_6860,N_5147,N_5126);
and U6861 (N_6861,N_5008,N_5742);
xnor U6862 (N_6862,N_5021,N_5123);
xor U6863 (N_6863,N_5200,N_5831);
xnor U6864 (N_6864,N_5810,N_5217);
or U6865 (N_6865,N_5124,N_5826);
nor U6866 (N_6866,N_5536,N_5363);
nand U6867 (N_6867,N_5051,N_5788);
and U6868 (N_6868,N_5680,N_5299);
nor U6869 (N_6869,N_5172,N_5745);
xnor U6870 (N_6870,N_5883,N_5435);
nand U6871 (N_6871,N_5519,N_5418);
and U6872 (N_6872,N_5359,N_5451);
xor U6873 (N_6873,N_5788,N_5189);
or U6874 (N_6874,N_5936,N_5684);
and U6875 (N_6875,N_5655,N_5461);
and U6876 (N_6876,N_5587,N_5373);
xnor U6877 (N_6877,N_5578,N_5854);
xor U6878 (N_6878,N_5516,N_5398);
xor U6879 (N_6879,N_5231,N_5540);
nor U6880 (N_6880,N_5809,N_5524);
and U6881 (N_6881,N_5993,N_5666);
nand U6882 (N_6882,N_5360,N_5220);
nand U6883 (N_6883,N_5758,N_5729);
and U6884 (N_6884,N_5286,N_5144);
nor U6885 (N_6885,N_5789,N_5757);
nor U6886 (N_6886,N_5703,N_5968);
xnor U6887 (N_6887,N_5960,N_5383);
nand U6888 (N_6888,N_5726,N_5906);
nand U6889 (N_6889,N_5146,N_5557);
xor U6890 (N_6890,N_5200,N_5622);
nand U6891 (N_6891,N_5157,N_5695);
or U6892 (N_6892,N_5942,N_5014);
or U6893 (N_6893,N_5577,N_5029);
xnor U6894 (N_6894,N_5133,N_5447);
xnor U6895 (N_6895,N_5205,N_5485);
or U6896 (N_6896,N_5932,N_5337);
and U6897 (N_6897,N_5888,N_5072);
xor U6898 (N_6898,N_5934,N_5833);
and U6899 (N_6899,N_5211,N_5748);
and U6900 (N_6900,N_5136,N_5645);
nor U6901 (N_6901,N_5036,N_5143);
and U6902 (N_6902,N_5725,N_5637);
nand U6903 (N_6903,N_5621,N_5228);
nand U6904 (N_6904,N_5938,N_5366);
and U6905 (N_6905,N_5322,N_5698);
and U6906 (N_6906,N_5650,N_5326);
nand U6907 (N_6907,N_5891,N_5430);
nor U6908 (N_6908,N_5844,N_5855);
nand U6909 (N_6909,N_5938,N_5982);
or U6910 (N_6910,N_5341,N_5966);
nand U6911 (N_6911,N_5247,N_5546);
nand U6912 (N_6912,N_5001,N_5339);
xor U6913 (N_6913,N_5851,N_5303);
xnor U6914 (N_6914,N_5273,N_5123);
nor U6915 (N_6915,N_5795,N_5919);
or U6916 (N_6916,N_5221,N_5149);
nor U6917 (N_6917,N_5295,N_5237);
nor U6918 (N_6918,N_5594,N_5872);
xor U6919 (N_6919,N_5795,N_5334);
or U6920 (N_6920,N_5550,N_5772);
or U6921 (N_6921,N_5869,N_5384);
xor U6922 (N_6922,N_5842,N_5296);
nand U6923 (N_6923,N_5406,N_5946);
xnor U6924 (N_6924,N_5905,N_5130);
nor U6925 (N_6925,N_5017,N_5738);
nand U6926 (N_6926,N_5229,N_5164);
nand U6927 (N_6927,N_5734,N_5097);
or U6928 (N_6928,N_5604,N_5655);
nand U6929 (N_6929,N_5613,N_5492);
nand U6930 (N_6930,N_5477,N_5293);
and U6931 (N_6931,N_5181,N_5522);
nand U6932 (N_6932,N_5368,N_5530);
and U6933 (N_6933,N_5601,N_5316);
xnor U6934 (N_6934,N_5654,N_5446);
and U6935 (N_6935,N_5953,N_5743);
nor U6936 (N_6936,N_5636,N_5098);
or U6937 (N_6937,N_5173,N_5294);
or U6938 (N_6938,N_5695,N_5244);
nor U6939 (N_6939,N_5532,N_5165);
or U6940 (N_6940,N_5958,N_5289);
or U6941 (N_6941,N_5081,N_5689);
or U6942 (N_6942,N_5752,N_5427);
and U6943 (N_6943,N_5314,N_5761);
or U6944 (N_6944,N_5993,N_5071);
nor U6945 (N_6945,N_5073,N_5556);
and U6946 (N_6946,N_5691,N_5614);
or U6947 (N_6947,N_5290,N_5004);
xnor U6948 (N_6948,N_5185,N_5179);
nand U6949 (N_6949,N_5999,N_5231);
and U6950 (N_6950,N_5718,N_5689);
nand U6951 (N_6951,N_5572,N_5316);
xor U6952 (N_6952,N_5592,N_5809);
and U6953 (N_6953,N_5740,N_5979);
nand U6954 (N_6954,N_5443,N_5539);
and U6955 (N_6955,N_5828,N_5309);
nor U6956 (N_6956,N_5851,N_5778);
or U6957 (N_6957,N_5576,N_5674);
xor U6958 (N_6958,N_5212,N_5936);
and U6959 (N_6959,N_5246,N_5755);
and U6960 (N_6960,N_5089,N_5320);
xor U6961 (N_6961,N_5458,N_5680);
or U6962 (N_6962,N_5791,N_5790);
nor U6963 (N_6963,N_5868,N_5958);
xnor U6964 (N_6964,N_5665,N_5873);
or U6965 (N_6965,N_5420,N_5694);
nor U6966 (N_6966,N_5837,N_5747);
or U6967 (N_6967,N_5522,N_5955);
xnor U6968 (N_6968,N_5107,N_5625);
or U6969 (N_6969,N_5388,N_5253);
or U6970 (N_6970,N_5170,N_5405);
or U6971 (N_6971,N_5434,N_5288);
nand U6972 (N_6972,N_5189,N_5551);
and U6973 (N_6973,N_5402,N_5704);
nor U6974 (N_6974,N_5251,N_5267);
xor U6975 (N_6975,N_5788,N_5425);
xor U6976 (N_6976,N_5013,N_5054);
nor U6977 (N_6977,N_5563,N_5351);
nand U6978 (N_6978,N_5528,N_5113);
or U6979 (N_6979,N_5506,N_5660);
nor U6980 (N_6980,N_5982,N_5528);
xor U6981 (N_6981,N_5296,N_5766);
and U6982 (N_6982,N_5188,N_5453);
xnor U6983 (N_6983,N_5513,N_5112);
nor U6984 (N_6984,N_5227,N_5929);
nand U6985 (N_6985,N_5418,N_5707);
or U6986 (N_6986,N_5597,N_5305);
or U6987 (N_6987,N_5291,N_5741);
and U6988 (N_6988,N_5338,N_5378);
nand U6989 (N_6989,N_5853,N_5167);
nor U6990 (N_6990,N_5673,N_5988);
nand U6991 (N_6991,N_5548,N_5239);
xor U6992 (N_6992,N_5598,N_5157);
and U6993 (N_6993,N_5257,N_5799);
or U6994 (N_6994,N_5448,N_5059);
nand U6995 (N_6995,N_5189,N_5302);
or U6996 (N_6996,N_5655,N_5986);
nor U6997 (N_6997,N_5670,N_5735);
nand U6998 (N_6998,N_5393,N_5497);
nand U6999 (N_6999,N_5769,N_5800);
xor U7000 (N_7000,N_6585,N_6117);
xnor U7001 (N_7001,N_6554,N_6630);
or U7002 (N_7002,N_6744,N_6518);
or U7003 (N_7003,N_6959,N_6365);
nor U7004 (N_7004,N_6688,N_6353);
nand U7005 (N_7005,N_6780,N_6083);
nand U7006 (N_7006,N_6437,N_6927);
or U7007 (N_7007,N_6604,N_6726);
and U7008 (N_7008,N_6636,N_6860);
and U7009 (N_7009,N_6292,N_6398);
and U7010 (N_7010,N_6031,N_6799);
nor U7011 (N_7011,N_6017,N_6970);
nor U7012 (N_7012,N_6277,N_6490);
nand U7013 (N_7013,N_6038,N_6296);
or U7014 (N_7014,N_6946,N_6281);
nand U7015 (N_7015,N_6596,N_6136);
nand U7016 (N_7016,N_6323,N_6521);
nand U7017 (N_7017,N_6449,N_6631);
nor U7018 (N_7018,N_6489,N_6987);
nor U7019 (N_7019,N_6240,N_6219);
xnor U7020 (N_7020,N_6293,N_6516);
or U7021 (N_7021,N_6078,N_6924);
and U7022 (N_7022,N_6629,N_6070);
xnor U7023 (N_7023,N_6790,N_6994);
and U7024 (N_7024,N_6395,N_6053);
and U7025 (N_7025,N_6522,N_6228);
xnor U7026 (N_7026,N_6304,N_6874);
nor U7027 (N_7027,N_6366,N_6607);
and U7028 (N_7028,N_6798,N_6039);
nand U7029 (N_7029,N_6127,N_6124);
nor U7030 (N_7030,N_6947,N_6656);
xnor U7031 (N_7031,N_6652,N_6092);
and U7032 (N_7032,N_6741,N_6737);
or U7033 (N_7033,N_6718,N_6575);
and U7034 (N_7034,N_6103,N_6900);
and U7035 (N_7035,N_6878,N_6133);
and U7036 (N_7036,N_6479,N_6176);
or U7037 (N_7037,N_6020,N_6517);
nand U7038 (N_7038,N_6760,N_6699);
or U7039 (N_7039,N_6894,N_6451);
xnor U7040 (N_7040,N_6976,N_6907);
xor U7041 (N_7041,N_6553,N_6601);
nand U7042 (N_7042,N_6658,N_6137);
or U7043 (N_7043,N_6319,N_6423);
or U7044 (N_7044,N_6359,N_6742);
or U7045 (N_7045,N_6581,N_6386);
nand U7046 (N_7046,N_6996,N_6298);
and U7047 (N_7047,N_6331,N_6580);
nand U7048 (N_7048,N_6873,N_6975);
nand U7049 (N_7049,N_6301,N_6480);
and U7050 (N_7050,N_6108,N_6569);
xnor U7051 (N_7051,N_6081,N_6122);
nand U7052 (N_7052,N_6379,N_6226);
nor U7053 (N_7053,N_6843,N_6307);
nand U7054 (N_7054,N_6134,N_6837);
xor U7055 (N_7055,N_6797,N_6417);
xor U7056 (N_7056,N_6795,N_6671);
xor U7057 (N_7057,N_6220,N_6368);
xnor U7058 (N_7058,N_6154,N_6239);
or U7059 (N_7059,N_6833,N_6495);
or U7060 (N_7060,N_6146,N_6863);
xnor U7061 (N_7061,N_6785,N_6236);
nand U7062 (N_7062,N_6338,N_6888);
nor U7063 (N_7063,N_6700,N_6121);
or U7064 (N_7064,N_6761,N_6381);
nor U7065 (N_7065,N_6993,N_6642);
nor U7066 (N_7066,N_6838,N_6257);
xnor U7067 (N_7067,N_6937,N_6327);
nand U7068 (N_7068,N_6118,N_6782);
nand U7069 (N_7069,N_6261,N_6675);
nand U7070 (N_7070,N_6592,N_6267);
nand U7071 (N_7071,N_6141,N_6617);
and U7072 (N_7072,N_6673,N_6767);
xor U7073 (N_7073,N_6965,N_6275);
nor U7074 (N_7074,N_6135,N_6171);
and U7075 (N_7075,N_6724,N_6579);
and U7076 (N_7076,N_6251,N_6558);
nand U7077 (N_7077,N_6457,N_6500);
nor U7078 (N_7078,N_6345,N_6311);
nand U7079 (N_7079,N_6882,N_6619);
xnor U7080 (N_7080,N_6082,N_6434);
xor U7081 (N_7081,N_6541,N_6828);
nor U7082 (N_7082,N_6035,N_6650);
nand U7083 (N_7083,N_6736,N_6126);
nand U7084 (N_7084,N_6628,N_6986);
xor U7085 (N_7085,N_6485,N_6729);
nand U7086 (N_7086,N_6163,N_6106);
and U7087 (N_7087,N_6546,N_6041);
nand U7088 (N_7088,N_6145,N_6022);
or U7089 (N_7089,N_6661,N_6404);
nor U7090 (N_7090,N_6291,N_6599);
nor U7091 (N_7091,N_6356,N_6060);
nand U7092 (N_7092,N_6635,N_6468);
or U7093 (N_7093,N_6094,N_6271);
nor U7094 (N_7094,N_6476,N_6250);
or U7095 (N_7095,N_6730,N_6189);
xnor U7096 (N_7096,N_6354,N_6416);
xor U7097 (N_7097,N_6602,N_6861);
or U7098 (N_7098,N_6979,N_6960);
xnor U7099 (N_7099,N_6977,N_6971);
nor U7100 (N_7100,N_6701,N_6911);
and U7101 (N_7101,N_6152,N_6034);
or U7102 (N_7102,N_6571,N_6586);
nand U7103 (N_7103,N_6225,N_6180);
nand U7104 (N_7104,N_6009,N_6156);
and U7105 (N_7105,N_6640,N_6711);
xnor U7106 (N_7106,N_6666,N_6218);
xnor U7107 (N_7107,N_6390,N_6567);
nor U7108 (N_7108,N_6932,N_6100);
nor U7109 (N_7109,N_6668,N_6549);
xor U7110 (N_7110,N_6821,N_6274);
nor U7111 (N_7111,N_6066,N_6295);
and U7112 (N_7112,N_6852,N_6004);
xor U7113 (N_7113,N_6392,N_6372);
nor U7114 (N_7114,N_6660,N_6164);
nor U7115 (N_7115,N_6680,N_6046);
xor U7116 (N_7116,N_6371,N_6346);
nand U7117 (N_7117,N_6936,N_6459);
or U7118 (N_7118,N_6535,N_6028);
or U7119 (N_7119,N_6374,N_6101);
xnor U7120 (N_7120,N_6119,N_6923);
xnor U7121 (N_7121,N_6641,N_6887);
or U7122 (N_7122,N_6759,N_6877);
xor U7123 (N_7123,N_6938,N_6032);
and U7124 (N_7124,N_6400,N_6095);
nand U7125 (N_7125,N_6132,N_6322);
and U7126 (N_7126,N_6804,N_6445);
nor U7127 (N_7127,N_6144,N_6123);
nand U7128 (N_7128,N_6065,N_6564);
nor U7129 (N_7129,N_6462,N_6672);
nand U7130 (N_7130,N_6857,N_6363);
nand U7131 (N_7131,N_6069,N_6183);
nor U7132 (N_7132,N_6308,N_6576);
nand U7133 (N_7133,N_6502,N_6870);
nor U7134 (N_7134,N_6318,N_6254);
or U7135 (N_7135,N_6234,N_6647);
xnor U7136 (N_7136,N_6302,N_6347);
or U7137 (N_7137,N_6011,N_6273);
and U7138 (N_7138,N_6283,N_6375);
xor U7139 (N_7139,N_6568,N_6844);
nor U7140 (N_7140,N_6683,N_6201);
nand U7141 (N_7141,N_6173,N_6488);
or U7142 (N_7142,N_6279,N_6620);
and U7143 (N_7143,N_6350,N_6955);
nand U7144 (N_7144,N_6403,N_6950);
xor U7145 (N_7145,N_6868,N_6645);
or U7146 (N_7146,N_6875,N_6869);
or U7147 (N_7147,N_6942,N_6505);
or U7148 (N_7148,N_6918,N_6786);
nand U7149 (N_7149,N_6191,N_6633);
xor U7150 (N_7150,N_6775,N_6627);
nand U7151 (N_7151,N_6836,N_6985);
and U7152 (N_7152,N_6847,N_6961);
nand U7153 (N_7153,N_6320,N_6430);
nand U7154 (N_7154,N_6952,N_6036);
or U7155 (N_7155,N_6482,N_6845);
nor U7156 (N_7156,N_6334,N_6886);
nor U7157 (N_7157,N_6461,N_6526);
or U7158 (N_7158,N_6026,N_6948);
xor U7159 (N_7159,N_6249,N_6397);
nand U7160 (N_7160,N_6899,N_6625);
nor U7161 (N_7161,N_6754,N_6727);
or U7162 (N_7162,N_6380,N_6357);
xor U7163 (N_7163,N_6056,N_6590);
xnor U7164 (N_7164,N_6084,N_6957);
xnor U7165 (N_7165,N_6194,N_6367);
and U7166 (N_7166,N_6897,N_6045);
or U7167 (N_7167,N_6405,N_6895);
nor U7168 (N_7168,N_6475,N_6207);
nor U7169 (N_7169,N_6755,N_6494);
or U7170 (N_7170,N_6704,N_6533);
xnor U7171 (N_7171,N_6665,N_6051);
nor U7172 (N_7172,N_6452,N_6120);
xnor U7173 (N_7173,N_6536,N_6075);
nor U7174 (N_7174,N_6543,N_6231);
nor U7175 (N_7175,N_6678,N_6829);
and U7176 (N_7176,N_6953,N_6128);
or U7177 (N_7177,N_6259,N_6916);
and U7178 (N_7178,N_6284,N_6248);
or U7179 (N_7179,N_6618,N_6548);
or U7180 (N_7180,N_6968,N_6687);
nor U7181 (N_7181,N_6890,N_6748);
nand U7182 (N_7182,N_6740,N_6995);
nand U7183 (N_7183,N_6615,N_6393);
or U7184 (N_7184,N_6603,N_6040);
and U7185 (N_7185,N_6424,N_6030);
nand U7186 (N_7186,N_6098,N_6179);
nor U7187 (N_7187,N_6426,N_6150);
xor U7188 (N_7188,N_6988,N_6088);
nor U7189 (N_7189,N_6112,N_6401);
or U7190 (N_7190,N_6238,N_6871);
xor U7191 (N_7191,N_6733,N_6697);
nor U7192 (N_7192,N_6728,N_6012);
nand U7193 (N_7193,N_6486,N_6364);
or U7194 (N_7194,N_6824,N_6657);
nor U7195 (N_7195,N_6605,N_6949);
or U7196 (N_7196,N_6966,N_6609);
nand U7197 (N_7197,N_6632,N_6382);
xnor U7198 (N_7198,N_6165,N_6243);
and U7199 (N_7199,N_6503,N_6547);
or U7200 (N_7200,N_6309,N_6738);
and U7201 (N_7201,N_6922,N_6802);
xnor U7202 (N_7202,N_6974,N_6578);
or U7203 (N_7203,N_6204,N_6872);
nor U7204 (N_7204,N_6743,N_6206);
nor U7205 (N_7205,N_6749,N_6278);
or U7206 (N_7206,N_6623,N_6529);
xor U7207 (N_7207,N_6450,N_6634);
or U7208 (N_7208,N_6787,N_6762);
nor U7209 (N_7209,N_6174,N_6102);
xor U7210 (N_7210,N_6637,N_6825);
nor U7211 (N_7211,N_6235,N_6294);
or U7212 (N_7212,N_6385,N_6941);
and U7213 (N_7213,N_6280,N_6429);
nand U7214 (N_7214,N_6286,N_6812);
and U7215 (N_7215,N_6209,N_6160);
and U7216 (N_7216,N_6244,N_6667);
nor U7217 (N_7217,N_6138,N_6674);
or U7218 (N_7218,N_6407,N_6989);
nor U7219 (N_7219,N_6999,N_6085);
nand U7220 (N_7220,N_6693,N_6444);
and U7221 (N_7221,N_6747,N_6972);
xnor U7222 (N_7222,N_6614,N_6469);
nand U7223 (N_7223,N_6440,N_6708);
nor U7224 (N_7224,N_6792,N_6458);
nand U7225 (N_7225,N_6007,N_6698);
nor U7226 (N_7226,N_6545,N_6597);
and U7227 (N_7227,N_6717,N_6481);
nand U7228 (N_7228,N_6893,N_6958);
nand U7229 (N_7229,N_6187,N_6441);
and U7230 (N_7230,N_6770,N_6841);
and U7231 (N_7231,N_6981,N_6202);
nor U7232 (N_7232,N_6252,N_6501);
or U7233 (N_7233,N_6467,N_6655);
nand U7234 (N_7234,N_6373,N_6559);
or U7235 (N_7235,N_6216,N_6776);
xor U7236 (N_7236,N_6969,N_6344);
or U7237 (N_7237,N_6313,N_6791);
or U7238 (N_7238,N_6237,N_6919);
nor U7239 (N_7239,N_6879,N_6714);
nor U7240 (N_7240,N_6910,N_6933);
xnor U7241 (N_7241,N_6456,N_6734);
or U7242 (N_7242,N_6624,N_6422);
nand U7243 (N_7243,N_6925,N_6842);
nand U7244 (N_7244,N_6091,N_6431);
or U7245 (N_7245,N_6352,N_6362);
xor U7246 (N_7246,N_6396,N_6266);
nor U7247 (N_7247,N_6210,N_6412);
or U7248 (N_7248,N_6814,N_6677);
xnor U7249 (N_7249,N_6856,N_6834);
and U7250 (N_7250,N_6303,N_6794);
xnor U7251 (N_7251,N_6466,N_6622);
or U7252 (N_7252,N_6169,N_6783);
and U7253 (N_7253,N_6528,N_6214);
and U7254 (N_7254,N_6534,N_6884);
or U7255 (N_7255,N_6768,N_6185);
or U7256 (N_7256,N_6341,N_6720);
xor U7257 (N_7257,N_6757,N_6316);
nand U7258 (N_7258,N_6142,N_6491);
and U7259 (N_7259,N_6565,N_6453);
and U7260 (N_7260,N_6213,N_6696);
or U7261 (N_7261,N_6913,N_6351);
and U7262 (N_7262,N_6676,N_6846);
and U7263 (N_7263,N_6167,N_6333);
and U7264 (N_7264,N_6161,N_6756);
nor U7265 (N_7265,N_6713,N_6954);
nand U7266 (N_7266,N_6241,N_6027);
nor U7267 (N_7267,N_6073,N_6312);
xnor U7268 (N_7268,N_6653,N_6514);
nand U7269 (N_7269,N_6175,N_6264);
nand U7270 (N_7270,N_6096,N_6473);
xor U7271 (N_7271,N_6663,N_6914);
nor U7272 (N_7272,N_6725,N_6552);
and U7273 (N_7273,N_6811,N_6892);
or U7274 (N_7274,N_6116,N_6731);
xor U7275 (N_7275,N_6413,N_6439);
and U7276 (N_7276,N_6832,N_6143);
and U7277 (N_7277,N_6212,N_6158);
xnor U7278 (N_7278,N_6391,N_6686);
and U7279 (N_7279,N_6796,N_6903);
and U7280 (N_7280,N_6735,N_6325);
nor U7281 (N_7281,N_6172,N_6186);
nor U7282 (N_7282,N_6583,N_6931);
or U7283 (N_7283,N_6550,N_6463);
nor U7284 (N_7284,N_6348,N_6166);
nand U7285 (N_7285,N_6662,N_6613);
and U7286 (N_7286,N_6399,N_6355);
nor U7287 (N_7287,N_6561,N_6648);
xnor U7288 (N_7288,N_6818,N_6710);
or U7289 (N_7289,N_6556,N_6052);
nor U7290 (N_7290,N_6600,N_6854);
nand U7291 (N_7291,N_6067,N_6509);
nand U7292 (N_7292,N_6448,N_6498);
and U7293 (N_7293,N_6059,N_6200);
xor U7294 (N_7294,N_6008,N_6507);
nand U7295 (N_7295,N_6643,N_6370);
and U7296 (N_7296,N_6419,N_6188);
nor U7297 (N_7297,N_6420,N_6940);
xor U7298 (N_7298,N_6800,N_6433);
nor U7299 (N_7299,N_6902,N_6428);
xor U7300 (N_7300,N_6898,N_6998);
xnor U7301 (N_7301,N_6807,N_6840);
or U7302 (N_7302,N_6808,N_6848);
and U7303 (N_7303,N_6061,N_6584);
xor U7304 (N_7304,N_6654,N_6793);
nor U7305 (N_7305,N_6010,N_6182);
or U7306 (N_7306,N_6992,N_6157);
and U7307 (N_7307,N_6197,N_6835);
nand U7308 (N_7308,N_6669,N_6025);
xor U7309 (N_7309,N_6520,N_6511);
xor U7310 (N_7310,N_6506,N_6722);
nor U7311 (N_7311,N_6865,N_6178);
or U7312 (N_7312,N_6224,N_6616);
xor U7313 (N_7313,N_6497,N_6709);
nand U7314 (N_7314,N_6018,N_6287);
nand U7315 (N_7315,N_6229,N_6855);
nor U7316 (N_7316,N_6033,N_6258);
and U7317 (N_7317,N_6064,N_6199);
or U7318 (N_7318,N_6523,N_6299);
nand U7319 (N_7319,N_6504,N_6317);
nor U7320 (N_7320,N_6268,N_6908);
nor U7321 (N_7321,N_6750,N_6255);
xnor U7322 (N_7322,N_6525,N_6074);
or U7323 (N_7323,N_6029,N_6148);
and U7324 (N_7324,N_6217,N_6436);
or U7325 (N_7325,N_6080,N_6823);
nand U7326 (N_7326,N_6377,N_6086);
nor U7327 (N_7327,N_6880,N_6378);
or U7328 (N_7328,N_6072,N_6774);
nor U7329 (N_7329,N_6245,N_6198);
nor U7330 (N_7330,N_6184,N_6766);
xor U7331 (N_7331,N_6827,N_6021);
xnor U7332 (N_7332,N_6926,N_6589);
nand U7333 (N_7333,N_6315,N_6336);
nor U7334 (N_7334,N_6001,N_6510);
and U7335 (N_7335,N_6772,N_6256);
nand U7336 (N_7336,N_6048,N_6705);
or U7337 (N_7337,N_6360,N_6421);
nand U7338 (N_7338,N_6232,N_6773);
or U7339 (N_7339,N_6649,N_6889);
and U7340 (N_7340,N_6015,N_6626);
nor U7341 (N_7341,N_6651,N_6883);
and U7342 (N_7342,N_6104,N_6867);
or U7343 (N_7343,N_6002,N_6097);
xor U7344 (N_7344,N_6659,N_6111);
xnor U7345 (N_7345,N_6830,N_6990);
nand U7346 (N_7346,N_6109,N_6443);
nand U7347 (N_7347,N_6915,N_6765);
or U7348 (N_7348,N_6859,N_6904);
or U7349 (N_7349,N_6695,N_6858);
nor U7350 (N_7350,N_6447,N_6415);
xnor U7351 (N_7351,N_6263,N_6964);
nor U7352 (N_7352,N_6876,N_6909);
nand U7353 (N_7353,N_6920,N_6557);
nand U7354 (N_7354,N_6771,N_6023);
xnor U7355 (N_7355,N_6921,N_6905);
nor U7356 (N_7356,N_6788,N_6777);
nor U7357 (N_7357,N_6276,N_6442);
nor U7358 (N_7358,N_6591,N_6570);
nand U7359 (N_7359,N_6153,N_6820);
nand U7360 (N_7360,N_6973,N_6131);
and U7361 (N_7361,N_6538,N_6155);
nor U7362 (N_7362,N_6418,N_6044);
and U7363 (N_7363,N_6929,N_6991);
and U7364 (N_7364,N_6000,N_6297);
or U7365 (N_7365,N_6712,N_6435);
xor U7366 (N_7366,N_6384,N_6037);
nor U7367 (N_7367,N_6896,N_6732);
xor U7368 (N_7368,N_6751,N_6049);
xnor U7369 (N_7369,N_6068,N_6269);
xnor U7370 (N_7370,N_6335,N_6980);
and U7371 (N_7371,N_6935,N_6555);
and U7372 (N_7372,N_6478,N_6409);
nand U7373 (N_7373,N_6881,N_6057);
or U7374 (N_7374,N_6956,N_6162);
xor U7375 (N_7375,N_6809,N_6260);
or U7376 (N_7376,N_6944,N_6050);
nand U7377 (N_7377,N_6912,N_6129);
and U7378 (N_7378,N_6196,N_6388);
nor U7379 (N_7379,N_6310,N_6901);
or U7380 (N_7380,N_6472,N_6389);
nor U7381 (N_7381,N_6850,N_6272);
nor U7382 (N_7382,N_6906,N_6764);
or U7383 (N_7383,N_6321,N_6242);
nand U7384 (N_7384,N_6723,N_6519);
xor U7385 (N_7385,N_6438,N_6527);
nor U7386 (N_7386,N_6611,N_6329);
or U7387 (N_7387,N_6513,N_6125);
or U7388 (N_7388,N_6679,N_6151);
and U7389 (N_7389,N_6512,N_6917);
or U7390 (N_7390,N_6691,N_6531);
or U7391 (N_7391,N_6071,N_6464);
nand U7392 (N_7392,N_6997,N_6427);
or U7393 (N_7393,N_6460,N_6684);
and U7394 (N_7394,N_6962,N_6951);
and U7395 (N_7395,N_6746,N_6265);
nor U7396 (N_7396,N_6606,N_6769);
or U7397 (N_7397,N_6005,N_6815);
and U7398 (N_7398,N_6978,N_6573);
or U7399 (N_7399,N_6465,N_6483);
xnor U7400 (N_7400,N_6562,N_6337);
nand U7401 (N_7401,N_6499,N_6168);
xnor U7402 (N_7402,N_6721,N_6147);
xnor U7403 (N_7403,N_6484,N_6703);
nor U7404 (N_7404,N_6690,N_6339);
nand U7405 (N_7405,N_6934,N_6864);
and U7406 (N_7406,N_6411,N_6612);
or U7407 (N_7407,N_6816,N_6230);
nor U7408 (N_7408,N_6587,N_6719);
nand U7409 (N_7409,N_6387,N_6945);
nor U7410 (N_7410,N_6247,N_6582);
or U7411 (N_7411,N_6406,N_6332);
nand U7412 (N_7412,N_6190,N_6984);
or U7413 (N_7413,N_6446,N_6099);
or U7414 (N_7414,N_6801,N_6328);
or U7415 (N_7415,N_6493,N_6539);
or U7416 (N_7416,N_6314,N_6193);
and U7417 (N_7417,N_6928,N_6054);
xor U7418 (N_7418,N_6402,N_6849);
and U7419 (N_7419,N_6208,N_6544);
or U7420 (N_7420,N_6885,N_6745);
or U7421 (N_7421,N_6983,N_6306);
nor U7422 (N_7422,N_6043,N_6227);
nand U7423 (N_7423,N_6326,N_6817);
and U7424 (N_7424,N_6716,N_6159);
nand U7425 (N_7425,N_6560,N_6595);
nor U7426 (N_7426,N_6805,N_6810);
nor U7427 (N_7427,N_6967,N_6608);
nand U7428 (N_7428,N_6866,N_6508);
or U7429 (N_7429,N_6530,N_6089);
nand U7430 (N_7430,N_6223,N_6891);
and U7431 (N_7431,N_6140,N_6246);
and U7432 (N_7432,N_6682,N_6290);
xnor U7433 (N_7433,N_6047,N_6340);
nor U7434 (N_7434,N_6361,N_6685);
and U7435 (N_7435,N_6639,N_6003);
nand U7436 (N_7436,N_6542,N_6621);
xor U7437 (N_7437,N_6113,N_6288);
nor U7438 (N_7438,N_6215,N_6107);
nor U7439 (N_7439,N_6537,N_6789);
nor U7440 (N_7440,N_6692,N_6644);
nand U7441 (N_7441,N_6851,N_6487);
nor U7442 (N_7442,N_6532,N_6016);
nor U7443 (N_7443,N_6262,N_6598);
and U7444 (N_7444,N_6285,N_6753);
xor U7445 (N_7445,N_6130,N_6055);
xor U7446 (N_7446,N_6058,N_6110);
xnor U7447 (N_7447,N_6282,N_6170);
nand U7448 (N_7448,N_6819,N_6139);
nand U7449 (N_7449,N_6087,N_6982);
or U7450 (N_7450,N_6253,N_6638);
nand U7451 (N_7451,N_6149,N_6563);
and U7452 (N_7452,N_6572,N_6455);
xnor U7453 (N_7453,N_6474,N_6177);
xnor U7454 (N_7454,N_6862,N_6681);
or U7455 (N_7455,N_6477,N_6063);
nand U7456 (N_7456,N_6524,N_6019);
nand U7457 (N_7457,N_6289,N_6577);
nand U7458 (N_7458,N_6454,N_6414);
and U7459 (N_7459,N_6707,N_6079);
nand U7460 (N_7460,N_6963,N_6305);
nand U7461 (N_7461,N_6062,N_6014);
nand U7462 (N_7462,N_6930,N_6376);
nand U7463 (N_7463,N_6211,N_6181);
and U7464 (N_7464,N_6042,N_6076);
and U7465 (N_7465,N_6105,N_6383);
or U7466 (N_7466,N_6831,N_6222);
or U7467 (N_7467,N_6784,N_6471);
nor U7468 (N_7468,N_6822,N_6192);
or U7469 (N_7469,N_6646,N_6943);
nor U7470 (N_7470,N_6574,N_6551);
nor U7471 (N_7471,N_6470,N_6939);
nand U7472 (N_7472,N_6593,N_6758);
or U7473 (N_7473,N_6839,N_6739);
and U7474 (N_7474,N_6115,N_6689);
and U7475 (N_7475,N_6205,N_6706);
nor U7476 (N_7476,N_6515,N_6013);
and U7477 (N_7477,N_6610,N_6492);
xor U7478 (N_7478,N_6566,N_6233);
nor U7479 (N_7479,N_6752,N_6853);
xnor U7480 (N_7480,N_6432,N_6813);
nand U7481 (N_7481,N_6342,N_6203);
nand U7482 (N_7482,N_6195,N_6806);
nand U7483 (N_7483,N_6781,N_6093);
nor U7484 (N_7484,N_6330,N_6410);
or U7485 (N_7485,N_6221,N_6702);
nand U7486 (N_7486,N_6803,N_6540);
nand U7487 (N_7487,N_6694,N_6826);
xor U7488 (N_7488,N_6090,N_6594);
nor U7489 (N_7489,N_6006,N_6077);
and U7490 (N_7490,N_6349,N_6343);
nor U7491 (N_7491,N_6270,N_6408);
and U7492 (N_7492,N_6778,N_6300);
or U7493 (N_7493,N_6715,N_6670);
and U7494 (N_7494,N_6496,N_6358);
nor U7495 (N_7495,N_6324,N_6369);
or U7496 (N_7496,N_6394,N_6779);
xnor U7497 (N_7497,N_6664,N_6425);
nand U7498 (N_7498,N_6763,N_6588);
nor U7499 (N_7499,N_6114,N_6024);
and U7500 (N_7500,N_6050,N_6817);
nand U7501 (N_7501,N_6276,N_6056);
xor U7502 (N_7502,N_6293,N_6563);
nor U7503 (N_7503,N_6721,N_6837);
xor U7504 (N_7504,N_6986,N_6790);
or U7505 (N_7505,N_6857,N_6521);
xnor U7506 (N_7506,N_6523,N_6207);
nand U7507 (N_7507,N_6105,N_6004);
xnor U7508 (N_7508,N_6630,N_6774);
nor U7509 (N_7509,N_6832,N_6241);
nand U7510 (N_7510,N_6667,N_6450);
or U7511 (N_7511,N_6086,N_6671);
or U7512 (N_7512,N_6230,N_6479);
nor U7513 (N_7513,N_6240,N_6814);
nand U7514 (N_7514,N_6877,N_6115);
and U7515 (N_7515,N_6431,N_6594);
or U7516 (N_7516,N_6726,N_6302);
nor U7517 (N_7517,N_6559,N_6750);
nor U7518 (N_7518,N_6774,N_6802);
or U7519 (N_7519,N_6128,N_6037);
and U7520 (N_7520,N_6603,N_6508);
nor U7521 (N_7521,N_6428,N_6345);
or U7522 (N_7522,N_6201,N_6878);
and U7523 (N_7523,N_6496,N_6877);
xnor U7524 (N_7524,N_6257,N_6723);
nor U7525 (N_7525,N_6397,N_6105);
and U7526 (N_7526,N_6742,N_6116);
and U7527 (N_7527,N_6302,N_6111);
nor U7528 (N_7528,N_6435,N_6739);
or U7529 (N_7529,N_6349,N_6791);
nor U7530 (N_7530,N_6026,N_6798);
or U7531 (N_7531,N_6078,N_6038);
xnor U7532 (N_7532,N_6106,N_6800);
nand U7533 (N_7533,N_6098,N_6541);
nor U7534 (N_7534,N_6266,N_6693);
xor U7535 (N_7535,N_6524,N_6692);
nor U7536 (N_7536,N_6727,N_6810);
or U7537 (N_7537,N_6635,N_6582);
or U7538 (N_7538,N_6707,N_6500);
or U7539 (N_7539,N_6032,N_6513);
xor U7540 (N_7540,N_6555,N_6872);
and U7541 (N_7541,N_6207,N_6608);
nor U7542 (N_7542,N_6590,N_6357);
xnor U7543 (N_7543,N_6708,N_6349);
nor U7544 (N_7544,N_6211,N_6323);
and U7545 (N_7545,N_6204,N_6358);
nor U7546 (N_7546,N_6722,N_6765);
xor U7547 (N_7547,N_6834,N_6231);
and U7548 (N_7548,N_6821,N_6697);
nor U7549 (N_7549,N_6380,N_6600);
or U7550 (N_7550,N_6969,N_6957);
or U7551 (N_7551,N_6373,N_6052);
nor U7552 (N_7552,N_6098,N_6064);
nand U7553 (N_7553,N_6017,N_6125);
or U7554 (N_7554,N_6327,N_6270);
xnor U7555 (N_7555,N_6279,N_6449);
and U7556 (N_7556,N_6822,N_6041);
or U7557 (N_7557,N_6923,N_6773);
xnor U7558 (N_7558,N_6922,N_6112);
nand U7559 (N_7559,N_6845,N_6494);
nor U7560 (N_7560,N_6792,N_6252);
nand U7561 (N_7561,N_6992,N_6460);
nor U7562 (N_7562,N_6429,N_6879);
nand U7563 (N_7563,N_6870,N_6266);
or U7564 (N_7564,N_6461,N_6960);
nor U7565 (N_7565,N_6193,N_6191);
xnor U7566 (N_7566,N_6642,N_6766);
and U7567 (N_7567,N_6065,N_6821);
nor U7568 (N_7568,N_6052,N_6357);
nor U7569 (N_7569,N_6623,N_6207);
and U7570 (N_7570,N_6997,N_6460);
and U7571 (N_7571,N_6332,N_6927);
xnor U7572 (N_7572,N_6201,N_6519);
xor U7573 (N_7573,N_6253,N_6560);
nor U7574 (N_7574,N_6033,N_6945);
and U7575 (N_7575,N_6721,N_6450);
and U7576 (N_7576,N_6211,N_6604);
nand U7577 (N_7577,N_6261,N_6454);
nor U7578 (N_7578,N_6974,N_6991);
and U7579 (N_7579,N_6989,N_6178);
and U7580 (N_7580,N_6139,N_6360);
xor U7581 (N_7581,N_6052,N_6620);
nand U7582 (N_7582,N_6395,N_6538);
nor U7583 (N_7583,N_6967,N_6674);
nor U7584 (N_7584,N_6720,N_6849);
nand U7585 (N_7585,N_6547,N_6480);
nor U7586 (N_7586,N_6866,N_6522);
and U7587 (N_7587,N_6424,N_6860);
nand U7588 (N_7588,N_6890,N_6583);
or U7589 (N_7589,N_6821,N_6747);
xor U7590 (N_7590,N_6971,N_6233);
and U7591 (N_7591,N_6042,N_6538);
nor U7592 (N_7592,N_6402,N_6541);
or U7593 (N_7593,N_6494,N_6833);
and U7594 (N_7594,N_6926,N_6384);
xor U7595 (N_7595,N_6299,N_6132);
nand U7596 (N_7596,N_6085,N_6585);
nand U7597 (N_7597,N_6980,N_6518);
and U7598 (N_7598,N_6083,N_6436);
nand U7599 (N_7599,N_6693,N_6996);
or U7600 (N_7600,N_6663,N_6441);
xor U7601 (N_7601,N_6915,N_6044);
and U7602 (N_7602,N_6505,N_6225);
nand U7603 (N_7603,N_6324,N_6674);
nand U7604 (N_7604,N_6167,N_6911);
or U7605 (N_7605,N_6568,N_6472);
and U7606 (N_7606,N_6799,N_6830);
and U7607 (N_7607,N_6675,N_6938);
xor U7608 (N_7608,N_6146,N_6286);
nor U7609 (N_7609,N_6304,N_6677);
xnor U7610 (N_7610,N_6870,N_6366);
nand U7611 (N_7611,N_6152,N_6648);
nor U7612 (N_7612,N_6541,N_6829);
and U7613 (N_7613,N_6504,N_6006);
or U7614 (N_7614,N_6816,N_6958);
nand U7615 (N_7615,N_6276,N_6988);
or U7616 (N_7616,N_6841,N_6943);
xnor U7617 (N_7617,N_6638,N_6203);
nand U7618 (N_7618,N_6999,N_6624);
nand U7619 (N_7619,N_6873,N_6963);
or U7620 (N_7620,N_6497,N_6739);
xor U7621 (N_7621,N_6978,N_6577);
xnor U7622 (N_7622,N_6145,N_6819);
xor U7623 (N_7623,N_6427,N_6105);
and U7624 (N_7624,N_6162,N_6742);
and U7625 (N_7625,N_6857,N_6296);
and U7626 (N_7626,N_6335,N_6221);
and U7627 (N_7627,N_6438,N_6096);
or U7628 (N_7628,N_6545,N_6049);
and U7629 (N_7629,N_6503,N_6551);
xor U7630 (N_7630,N_6944,N_6013);
nand U7631 (N_7631,N_6796,N_6951);
xor U7632 (N_7632,N_6184,N_6594);
and U7633 (N_7633,N_6065,N_6898);
nand U7634 (N_7634,N_6993,N_6402);
nor U7635 (N_7635,N_6782,N_6887);
nand U7636 (N_7636,N_6578,N_6080);
nand U7637 (N_7637,N_6638,N_6955);
nand U7638 (N_7638,N_6875,N_6157);
nand U7639 (N_7639,N_6048,N_6269);
and U7640 (N_7640,N_6641,N_6207);
nand U7641 (N_7641,N_6473,N_6938);
nand U7642 (N_7642,N_6259,N_6187);
and U7643 (N_7643,N_6271,N_6701);
nor U7644 (N_7644,N_6823,N_6856);
xnor U7645 (N_7645,N_6671,N_6488);
xnor U7646 (N_7646,N_6248,N_6701);
and U7647 (N_7647,N_6135,N_6410);
or U7648 (N_7648,N_6488,N_6209);
nor U7649 (N_7649,N_6929,N_6885);
or U7650 (N_7650,N_6727,N_6131);
nor U7651 (N_7651,N_6732,N_6506);
nor U7652 (N_7652,N_6465,N_6265);
or U7653 (N_7653,N_6237,N_6434);
nor U7654 (N_7654,N_6036,N_6233);
or U7655 (N_7655,N_6073,N_6636);
or U7656 (N_7656,N_6122,N_6067);
xnor U7657 (N_7657,N_6907,N_6404);
xor U7658 (N_7658,N_6344,N_6950);
and U7659 (N_7659,N_6541,N_6404);
nand U7660 (N_7660,N_6646,N_6412);
or U7661 (N_7661,N_6722,N_6092);
nand U7662 (N_7662,N_6227,N_6756);
nor U7663 (N_7663,N_6096,N_6372);
xor U7664 (N_7664,N_6795,N_6390);
or U7665 (N_7665,N_6680,N_6020);
nand U7666 (N_7666,N_6299,N_6492);
nand U7667 (N_7667,N_6426,N_6897);
nand U7668 (N_7668,N_6292,N_6317);
or U7669 (N_7669,N_6314,N_6338);
and U7670 (N_7670,N_6862,N_6528);
or U7671 (N_7671,N_6386,N_6121);
and U7672 (N_7672,N_6562,N_6090);
and U7673 (N_7673,N_6052,N_6685);
or U7674 (N_7674,N_6058,N_6323);
xnor U7675 (N_7675,N_6641,N_6769);
nand U7676 (N_7676,N_6812,N_6485);
xnor U7677 (N_7677,N_6601,N_6888);
or U7678 (N_7678,N_6102,N_6347);
or U7679 (N_7679,N_6937,N_6649);
and U7680 (N_7680,N_6571,N_6649);
nand U7681 (N_7681,N_6433,N_6553);
xor U7682 (N_7682,N_6849,N_6055);
nand U7683 (N_7683,N_6679,N_6884);
and U7684 (N_7684,N_6289,N_6036);
and U7685 (N_7685,N_6574,N_6839);
and U7686 (N_7686,N_6341,N_6262);
and U7687 (N_7687,N_6667,N_6981);
and U7688 (N_7688,N_6968,N_6964);
nand U7689 (N_7689,N_6581,N_6665);
xnor U7690 (N_7690,N_6105,N_6378);
xnor U7691 (N_7691,N_6721,N_6500);
xor U7692 (N_7692,N_6045,N_6486);
xor U7693 (N_7693,N_6228,N_6179);
nand U7694 (N_7694,N_6669,N_6516);
or U7695 (N_7695,N_6516,N_6417);
nand U7696 (N_7696,N_6590,N_6042);
xor U7697 (N_7697,N_6034,N_6510);
nand U7698 (N_7698,N_6414,N_6563);
and U7699 (N_7699,N_6924,N_6809);
nor U7700 (N_7700,N_6063,N_6984);
xnor U7701 (N_7701,N_6616,N_6834);
nand U7702 (N_7702,N_6226,N_6776);
nor U7703 (N_7703,N_6537,N_6057);
or U7704 (N_7704,N_6921,N_6752);
and U7705 (N_7705,N_6253,N_6601);
or U7706 (N_7706,N_6299,N_6662);
xor U7707 (N_7707,N_6083,N_6018);
nor U7708 (N_7708,N_6207,N_6431);
and U7709 (N_7709,N_6619,N_6238);
xnor U7710 (N_7710,N_6169,N_6830);
or U7711 (N_7711,N_6406,N_6859);
nand U7712 (N_7712,N_6325,N_6474);
xor U7713 (N_7713,N_6948,N_6164);
or U7714 (N_7714,N_6495,N_6628);
xnor U7715 (N_7715,N_6608,N_6543);
and U7716 (N_7716,N_6925,N_6593);
xor U7717 (N_7717,N_6918,N_6326);
nor U7718 (N_7718,N_6137,N_6426);
and U7719 (N_7719,N_6315,N_6509);
nor U7720 (N_7720,N_6942,N_6972);
nor U7721 (N_7721,N_6524,N_6690);
and U7722 (N_7722,N_6586,N_6555);
xor U7723 (N_7723,N_6190,N_6508);
xor U7724 (N_7724,N_6887,N_6262);
and U7725 (N_7725,N_6144,N_6479);
nor U7726 (N_7726,N_6204,N_6827);
nor U7727 (N_7727,N_6567,N_6523);
or U7728 (N_7728,N_6610,N_6547);
and U7729 (N_7729,N_6977,N_6363);
or U7730 (N_7730,N_6641,N_6406);
and U7731 (N_7731,N_6501,N_6612);
and U7732 (N_7732,N_6037,N_6051);
nor U7733 (N_7733,N_6309,N_6306);
xnor U7734 (N_7734,N_6738,N_6660);
xor U7735 (N_7735,N_6400,N_6420);
nand U7736 (N_7736,N_6886,N_6636);
nand U7737 (N_7737,N_6936,N_6499);
xor U7738 (N_7738,N_6477,N_6719);
nand U7739 (N_7739,N_6551,N_6967);
nor U7740 (N_7740,N_6474,N_6654);
xnor U7741 (N_7741,N_6094,N_6783);
and U7742 (N_7742,N_6391,N_6330);
or U7743 (N_7743,N_6717,N_6101);
and U7744 (N_7744,N_6769,N_6818);
nand U7745 (N_7745,N_6966,N_6518);
or U7746 (N_7746,N_6422,N_6366);
and U7747 (N_7747,N_6667,N_6644);
nand U7748 (N_7748,N_6107,N_6940);
nor U7749 (N_7749,N_6085,N_6811);
nand U7750 (N_7750,N_6969,N_6338);
nor U7751 (N_7751,N_6749,N_6030);
nand U7752 (N_7752,N_6614,N_6094);
or U7753 (N_7753,N_6663,N_6540);
nor U7754 (N_7754,N_6363,N_6947);
nor U7755 (N_7755,N_6853,N_6758);
nand U7756 (N_7756,N_6962,N_6172);
or U7757 (N_7757,N_6012,N_6477);
xor U7758 (N_7758,N_6906,N_6960);
nor U7759 (N_7759,N_6381,N_6409);
nor U7760 (N_7760,N_6865,N_6898);
nand U7761 (N_7761,N_6881,N_6493);
or U7762 (N_7762,N_6822,N_6318);
and U7763 (N_7763,N_6566,N_6900);
or U7764 (N_7764,N_6007,N_6489);
nor U7765 (N_7765,N_6999,N_6016);
nor U7766 (N_7766,N_6824,N_6342);
nand U7767 (N_7767,N_6724,N_6858);
and U7768 (N_7768,N_6185,N_6872);
xnor U7769 (N_7769,N_6316,N_6106);
nor U7770 (N_7770,N_6602,N_6681);
nand U7771 (N_7771,N_6000,N_6348);
and U7772 (N_7772,N_6216,N_6618);
nor U7773 (N_7773,N_6379,N_6115);
and U7774 (N_7774,N_6568,N_6695);
xor U7775 (N_7775,N_6757,N_6539);
and U7776 (N_7776,N_6673,N_6386);
xor U7777 (N_7777,N_6254,N_6290);
and U7778 (N_7778,N_6819,N_6956);
xnor U7779 (N_7779,N_6207,N_6339);
xor U7780 (N_7780,N_6734,N_6203);
or U7781 (N_7781,N_6334,N_6754);
and U7782 (N_7782,N_6508,N_6744);
nor U7783 (N_7783,N_6706,N_6015);
or U7784 (N_7784,N_6484,N_6535);
xnor U7785 (N_7785,N_6128,N_6855);
nor U7786 (N_7786,N_6118,N_6078);
nor U7787 (N_7787,N_6813,N_6020);
or U7788 (N_7788,N_6951,N_6273);
nand U7789 (N_7789,N_6602,N_6813);
and U7790 (N_7790,N_6744,N_6780);
nand U7791 (N_7791,N_6789,N_6745);
nand U7792 (N_7792,N_6071,N_6584);
xnor U7793 (N_7793,N_6950,N_6958);
nor U7794 (N_7794,N_6711,N_6981);
nor U7795 (N_7795,N_6387,N_6220);
and U7796 (N_7796,N_6768,N_6155);
nand U7797 (N_7797,N_6502,N_6115);
nor U7798 (N_7798,N_6113,N_6082);
or U7799 (N_7799,N_6194,N_6492);
and U7800 (N_7800,N_6606,N_6657);
and U7801 (N_7801,N_6615,N_6574);
xnor U7802 (N_7802,N_6586,N_6017);
xnor U7803 (N_7803,N_6012,N_6279);
or U7804 (N_7804,N_6153,N_6230);
xor U7805 (N_7805,N_6410,N_6329);
nor U7806 (N_7806,N_6214,N_6539);
nand U7807 (N_7807,N_6250,N_6896);
or U7808 (N_7808,N_6880,N_6386);
and U7809 (N_7809,N_6648,N_6284);
and U7810 (N_7810,N_6683,N_6067);
or U7811 (N_7811,N_6664,N_6932);
and U7812 (N_7812,N_6634,N_6563);
nor U7813 (N_7813,N_6153,N_6567);
and U7814 (N_7814,N_6926,N_6037);
nor U7815 (N_7815,N_6736,N_6289);
or U7816 (N_7816,N_6537,N_6494);
or U7817 (N_7817,N_6803,N_6238);
xnor U7818 (N_7818,N_6143,N_6996);
or U7819 (N_7819,N_6229,N_6492);
and U7820 (N_7820,N_6455,N_6497);
or U7821 (N_7821,N_6498,N_6004);
nor U7822 (N_7822,N_6626,N_6285);
xnor U7823 (N_7823,N_6790,N_6716);
or U7824 (N_7824,N_6641,N_6606);
or U7825 (N_7825,N_6369,N_6965);
nor U7826 (N_7826,N_6720,N_6695);
nand U7827 (N_7827,N_6768,N_6760);
nor U7828 (N_7828,N_6469,N_6372);
or U7829 (N_7829,N_6845,N_6674);
nor U7830 (N_7830,N_6920,N_6241);
xor U7831 (N_7831,N_6686,N_6379);
nand U7832 (N_7832,N_6916,N_6430);
or U7833 (N_7833,N_6400,N_6855);
or U7834 (N_7834,N_6496,N_6250);
and U7835 (N_7835,N_6756,N_6532);
nand U7836 (N_7836,N_6835,N_6127);
nand U7837 (N_7837,N_6876,N_6545);
xor U7838 (N_7838,N_6644,N_6884);
xnor U7839 (N_7839,N_6891,N_6291);
or U7840 (N_7840,N_6569,N_6483);
or U7841 (N_7841,N_6037,N_6960);
nand U7842 (N_7842,N_6515,N_6657);
nand U7843 (N_7843,N_6727,N_6006);
nand U7844 (N_7844,N_6659,N_6764);
and U7845 (N_7845,N_6812,N_6456);
nand U7846 (N_7846,N_6577,N_6830);
or U7847 (N_7847,N_6532,N_6021);
or U7848 (N_7848,N_6954,N_6703);
and U7849 (N_7849,N_6170,N_6753);
nor U7850 (N_7850,N_6243,N_6276);
nand U7851 (N_7851,N_6549,N_6501);
xor U7852 (N_7852,N_6097,N_6578);
xnor U7853 (N_7853,N_6369,N_6969);
xor U7854 (N_7854,N_6418,N_6534);
or U7855 (N_7855,N_6511,N_6863);
or U7856 (N_7856,N_6604,N_6571);
nand U7857 (N_7857,N_6986,N_6730);
and U7858 (N_7858,N_6510,N_6891);
xor U7859 (N_7859,N_6772,N_6709);
xor U7860 (N_7860,N_6330,N_6121);
nand U7861 (N_7861,N_6846,N_6809);
xor U7862 (N_7862,N_6317,N_6489);
and U7863 (N_7863,N_6737,N_6384);
nand U7864 (N_7864,N_6265,N_6184);
and U7865 (N_7865,N_6704,N_6271);
nor U7866 (N_7866,N_6231,N_6981);
and U7867 (N_7867,N_6584,N_6197);
and U7868 (N_7868,N_6829,N_6267);
xor U7869 (N_7869,N_6755,N_6486);
nor U7870 (N_7870,N_6918,N_6973);
nand U7871 (N_7871,N_6655,N_6619);
or U7872 (N_7872,N_6807,N_6018);
and U7873 (N_7873,N_6095,N_6132);
xor U7874 (N_7874,N_6916,N_6787);
nand U7875 (N_7875,N_6367,N_6557);
and U7876 (N_7876,N_6694,N_6836);
nor U7877 (N_7877,N_6273,N_6172);
xnor U7878 (N_7878,N_6277,N_6727);
nand U7879 (N_7879,N_6334,N_6981);
nand U7880 (N_7880,N_6644,N_6948);
nand U7881 (N_7881,N_6720,N_6229);
xor U7882 (N_7882,N_6662,N_6282);
nor U7883 (N_7883,N_6127,N_6535);
and U7884 (N_7884,N_6933,N_6198);
and U7885 (N_7885,N_6660,N_6585);
nor U7886 (N_7886,N_6800,N_6884);
xor U7887 (N_7887,N_6884,N_6345);
nand U7888 (N_7888,N_6434,N_6526);
or U7889 (N_7889,N_6771,N_6069);
nand U7890 (N_7890,N_6648,N_6757);
and U7891 (N_7891,N_6738,N_6363);
or U7892 (N_7892,N_6953,N_6959);
nand U7893 (N_7893,N_6413,N_6324);
and U7894 (N_7894,N_6767,N_6794);
xor U7895 (N_7895,N_6091,N_6477);
xnor U7896 (N_7896,N_6122,N_6409);
nor U7897 (N_7897,N_6932,N_6308);
or U7898 (N_7898,N_6261,N_6509);
nor U7899 (N_7899,N_6798,N_6906);
or U7900 (N_7900,N_6510,N_6292);
or U7901 (N_7901,N_6273,N_6228);
and U7902 (N_7902,N_6358,N_6511);
nor U7903 (N_7903,N_6765,N_6621);
and U7904 (N_7904,N_6082,N_6854);
and U7905 (N_7905,N_6916,N_6762);
nand U7906 (N_7906,N_6805,N_6677);
or U7907 (N_7907,N_6133,N_6998);
nand U7908 (N_7908,N_6935,N_6968);
nor U7909 (N_7909,N_6522,N_6180);
nand U7910 (N_7910,N_6157,N_6814);
or U7911 (N_7911,N_6172,N_6182);
nand U7912 (N_7912,N_6411,N_6705);
or U7913 (N_7913,N_6078,N_6099);
nand U7914 (N_7914,N_6238,N_6774);
and U7915 (N_7915,N_6392,N_6202);
or U7916 (N_7916,N_6631,N_6923);
and U7917 (N_7917,N_6367,N_6461);
nand U7918 (N_7918,N_6146,N_6629);
and U7919 (N_7919,N_6758,N_6929);
or U7920 (N_7920,N_6417,N_6821);
and U7921 (N_7921,N_6866,N_6752);
xnor U7922 (N_7922,N_6426,N_6707);
or U7923 (N_7923,N_6662,N_6701);
xnor U7924 (N_7924,N_6175,N_6974);
nor U7925 (N_7925,N_6439,N_6416);
xnor U7926 (N_7926,N_6784,N_6300);
nand U7927 (N_7927,N_6392,N_6153);
nor U7928 (N_7928,N_6066,N_6279);
or U7929 (N_7929,N_6798,N_6004);
and U7930 (N_7930,N_6362,N_6744);
and U7931 (N_7931,N_6993,N_6168);
or U7932 (N_7932,N_6171,N_6414);
nand U7933 (N_7933,N_6035,N_6439);
or U7934 (N_7934,N_6261,N_6057);
xnor U7935 (N_7935,N_6464,N_6260);
or U7936 (N_7936,N_6423,N_6781);
or U7937 (N_7937,N_6274,N_6401);
nand U7938 (N_7938,N_6329,N_6934);
or U7939 (N_7939,N_6908,N_6534);
or U7940 (N_7940,N_6381,N_6339);
or U7941 (N_7941,N_6294,N_6030);
nor U7942 (N_7942,N_6839,N_6134);
nand U7943 (N_7943,N_6930,N_6175);
and U7944 (N_7944,N_6896,N_6799);
or U7945 (N_7945,N_6156,N_6146);
or U7946 (N_7946,N_6021,N_6424);
nor U7947 (N_7947,N_6632,N_6639);
or U7948 (N_7948,N_6064,N_6033);
or U7949 (N_7949,N_6594,N_6434);
nor U7950 (N_7950,N_6135,N_6874);
and U7951 (N_7951,N_6792,N_6514);
and U7952 (N_7952,N_6086,N_6816);
xor U7953 (N_7953,N_6580,N_6364);
xnor U7954 (N_7954,N_6007,N_6495);
and U7955 (N_7955,N_6029,N_6964);
and U7956 (N_7956,N_6296,N_6974);
or U7957 (N_7957,N_6668,N_6289);
and U7958 (N_7958,N_6127,N_6545);
and U7959 (N_7959,N_6690,N_6410);
or U7960 (N_7960,N_6905,N_6120);
nor U7961 (N_7961,N_6222,N_6429);
nand U7962 (N_7962,N_6258,N_6809);
and U7963 (N_7963,N_6322,N_6824);
nand U7964 (N_7964,N_6389,N_6280);
nand U7965 (N_7965,N_6948,N_6928);
nor U7966 (N_7966,N_6561,N_6470);
and U7967 (N_7967,N_6850,N_6508);
nand U7968 (N_7968,N_6065,N_6972);
nor U7969 (N_7969,N_6585,N_6444);
nand U7970 (N_7970,N_6294,N_6364);
xor U7971 (N_7971,N_6215,N_6531);
nor U7972 (N_7972,N_6472,N_6130);
xor U7973 (N_7973,N_6344,N_6726);
nand U7974 (N_7974,N_6010,N_6150);
nor U7975 (N_7975,N_6897,N_6915);
nand U7976 (N_7976,N_6344,N_6265);
and U7977 (N_7977,N_6322,N_6246);
nor U7978 (N_7978,N_6066,N_6774);
and U7979 (N_7979,N_6264,N_6864);
nor U7980 (N_7980,N_6268,N_6993);
nor U7981 (N_7981,N_6588,N_6756);
nand U7982 (N_7982,N_6179,N_6895);
nand U7983 (N_7983,N_6977,N_6415);
nand U7984 (N_7984,N_6390,N_6310);
nor U7985 (N_7985,N_6048,N_6813);
nor U7986 (N_7986,N_6447,N_6990);
nand U7987 (N_7987,N_6548,N_6963);
and U7988 (N_7988,N_6325,N_6756);
xnor U7989 (N_7989,N_6574,N_6816);
nand U7990 (N_7990,N_6981,N_6173);
nor U7991 (N_7991,N_6629,N_6041);
nand U7992 (N_7992,N_6231,N_6749);
or U7993 (N_7993,N_6506,N_6874);
nand U7994 (N_7994,N_6185,N_6084);
nand U7995 (N_7995,N_6586,N_6681);
nand U7996 (N_7996,N_6048,N_6984);
nand U7997 (N_7997,N_6077,N_6850);
nand U7998 (N_7998,N_6165,N_6805);
and U7999 (N_7999,N_6469,N_6027);
or U8000 (N_8000,N_7122,N_7626);
or U8001 (N_8001,N_7853,N_7939);
xnor U8002 (N_8002,N_7146,N_7461);
or U8003 (N_8003,N_7749,N_7035);
xnor U8004 (N_8004,N_7164,N_7265);
nand U8005 (N_8005,N_7020,N_7321);
xor U8006 (N_8006,N_7854,N_7133);
or U8007 (N_8007,N_7151,N_7501);
xnor U8008 (N_8008,N_7315,N_7834);
nand U8009 (N_8009,N_7410,N_7706);
or U8010 (N_8010,N_7629,N_7062);
and U8011 (N_8011,N_7992,N_7733);
nor U8012 (N_8012,N_7666,N_7227);
nand U8013 (N_8013,N_7096,N_7003);
and U8014 (N_8014,N_7181,N_7421);
nor U8015 (N_8015,N_7283,N_7211);
nand U8016 (N_8016,N_7068,N_7998);
xor U8017 (N_8017,N_7687,N_7288);
and U8018 (N_8018,N_7500,N_7643);
xor U8019 (N_8019,N_7638,N_7140);
nand U8020 (N_8020,N_7174,N_7021);
and U8021 (N_8021,N_7158,N_7284);
or U8022 (N_8022,N_7117,N_7595);
nor U8023 (N_8023,N_7273,N_7754);
nor U8024 (N_8024,N_7736,N_7898);
or U8025 (N_8025,N_7816,N_7921);
xor U8026 (N_8026,N_7098,N_7540);
or U8027 (N_8027,N_7730,N_7072);
and U8028 (N_8028,N_7884,N_7607);
nand U8029 (N_8029,N_7427,N_7585);
nor U8030 (N_8030,N_7069,N_7752);
or U8031 (N_8031,N_7539,N_7946);
xnor U8032 (N_8032,N_7195,N_7506);
xor U8033 (N_8033,N_7510,N_7938);
or U8034 (N_8034,N_7641,N_7570);
xnor U8035 (N_8035,N_7739,N_7502);
or U8036 (N_8036,N_7080,N_7823);
xnor U8037 (N_8037,N_7051,N_7490);
and U8038 (N_8038,N_7023,N_7779);
nand U8039 (N_8039,N_7449,N_7059);
and U8040 (N_8040,N_7339,N_7791);
xor U8041 (N_8041,N_7204,N_7916);
or U8042 (N_8042,N_7477,N_7362);
or U8043 (N_8043,N_7678,N_7968);
nor U8044 (N_8044,N_7577,N_7868);
or U8045 (N_8045,N_7030,N_7147);
and U8046 (N_8046,N_7392,N_7246);
nand U8047 (N_8047,N_7012,N_7932);
nor U8048 (N_8048,N_7919,N_7085);
nand U8049 (N_8049,N_7793,N_7381);
or U8050 (N_8050,N_7341,N_7159);
nand U8051 (N_8051,N_7416,N_7826);
nand U8052 (N_8052,N_7574,N_7034);
nor U8053 (N_8053,N_7877,N_7950);
xor U8054 (N_8054,N_7922,N_7179);
nand U8055 (N_8055,N_7657,N_7469);
and U8056 (N_8056,N_7157,N_7546);
or U8057 (N_8057,N_7267,N_7378);
nor U8058 (N_8058,N_7380,N_7497);
and U8059 (N_8059,N_7252,N_7617);
nand U8060 (N_8060,N_7930,N_7361);
or U8061 (N_8061,N_7698,N_7822);
or U8062 (N_8062,N_7905,N_7937);
nand U8063 (N_8063,N_7832,N_7766);
xor U8064 (N_8064,N_7060,N_7317);
or U8065 (N_8065,N_7013,N_7408);
xor U8066 (N_8066,N_7785,N_7987);
nand U8067 (N_8067,N_7705,N_7525);
or U8068 (N_8068,N_7512,N_7223);
and U8069 (N_8069,N_7763,N_7266);
or U8070 (N_8070,N_7241,N_7686);
nand U8071 (N_8071,N_7166,N_7444);
nand U8072 (N_8072,N_7095,N_7256);
nand U8073 (N_8073,N_7640,N_7611);
nor U8074 (N_8074,N_7802,N_7615);
nand U8075 (N_8075,N_7374,N_7821);
or U8076 (N_8076,N_7774,N_7828);
xnor U8077 (N_8077,N_7960,N_7353);
nor U8078 (N_8078,N_7304,N_7936);
xor U8079 (N_8079,N_7772,N_7695);
nand U8080 (N_8080,N_7762,N_7735);
nor U8081 (N_8081,N_7890,N_7104);
and U8082 (N_8082,N_7446,N_7907);
or U8083 (N_8083,N_7747,N_7505);
or U8084 (N_8084,N_7230,N_7818);
or U8085 (N_8085,N_7769,N_7126);
or U8086 (N_8086,N_7160,N_7584);
xor U8087 (N_8087,N_7533,N_7306);
nor U8088 (N_8088,N_7142,N_7670);
nand U8089 (N_8089,N_7679,N_7795);
nand U8090 (N_8090,N_7819,N_7291);
xnor U8091 (N_8091,N_7553,N_7172);
nand U8092 (N_8092,N_7168,N_7872);
xor U8093 (N_8093,N_7492,N_7295);
nand U8094 (N_8094,N_7005,N_7900);
nor U8095 (N_8095,N_7066,N_7229);
xor U8096 (N_8096,N_7709,N_7326);
nand U8097 (N_8097,N_7977,N_7677);
nor U8098 (N_8098,N_7419,N_7015);
nand U8099 (N_8099,N_7789,N_7524);
nand U8100 (N_8100,N_7849,N_7278);
nand U8101 (N_8101,N_7487,N_7485);
xor U8102 (N_8102,N_7097,N_7714);
xor U8103 (N_8103,N_7275,N_7084);
xor U8104 (N_8104,N_7484,N_7162);
or U8105 (N_8105,N_7409,N_7475);
xor U8106 (N_8106,N_7741,N_7055);
or U8107 (N_8107,N_7951,N_7047);
or U8108 (N_8108,N_7141,N_7548);
or U8109 (N_8109,N_7587,N_7206);
nand U8110 (N_8110,N_7778,N_7010);
xnor U8111 (N_8111,N_7384,N_7797);
or U8112 (N_8112,N_7594,N_7568);
and U8113 (N_8113,N_7811,N_7559);
and U8114 (N_8114,N_7131,N_7282);
nand U8115 (N_8115,N_7031,N_7787);
and U8116 (N_8116,N_7780,N_7812);
nor U8117 (N_8117,N_7330,N_7001);
nor U8118 (N_8118,N_7534,N_7642);
nand U8119 (N_8119,N_7809,N_7620);
xnor U8120 (N_8120,N_7507,N_7776);
xnor U8121 (N_8121,N_7351,N_7447);
and U8122 (N_8122,N_7183,N_7239);
or U8123 (N_8123,N_7116,N_7700);
nor U8124 (N_8124,N_7026,N_7254);
and U8125 (N_8125,N_7891,N_7786);
and U8126 (N_8126,N_7926,N_7481);
or U8127 (N_8127,N_7025,N_7293);
nand U8128 (N_8128,N_7850,N_7324);
nand U8129 (N_8129,N_7990,N_7984);
nor U8130 (N_8130,N_7966,N_7532);
and U8131 (N_8131,N_7280,N_7250);
nand U8132 (N_8132,N_7573,N_7222);
and U8133 (N_8133,N_7794,N_7719);
xnor U8134 (N_8134,N_7903,N_7494);
nand U8135 (N_8135,N_7541,N_7048);
nor U8136 (N_8136,N_7301,N_7463);
or U8137 (N_8137,N_7344,N_7258);
or U8138 (N_8138,N_7989,N_7673);
nor U8139 (N_8139,N_7653,N_7137);
nor U8140 (N_8140,N_7155,N_7445);
nand U8141 (N_8141,N_7527,N_7486);
and U8142 (N_8142,N_7139,N_7336);
xnor U8143 (N_8143,N_7895,N_7543);
nand U8144 (N_8144,N_7008,N_7654);
nor U8145 (N_8145,N_7110,N_7127);
and U8146 (N_8146,N_7043,N_7090);
nor U8147 (N_8147,N_7333,N_7002);
nand U8148 (N_8148,N_7560,N_7129);
or U8149 (N_8149,N_7773,N_7053);
xor U8150 (N_8150,N_7439,N_7808);
nand U8151 (N_8151,N_7978,N_7400);
xor U8152 (N_8152,N_7651,N_7077);
xor U8153 (N_8153,N_7598,N_7526);
nor U8154 (N_8154,N_7454,N_7969);
or U8155 (N_8155,N_7833,N_7228);
and U8156 (N_8156,N_7894,N_7871);
or U8157 (N_8157,N_7307,N_7269);
or U8158 (N_8158,N_7661,N_7538);
nor U8159 (N_8159,N_7892,N_7609);
or U8160 (N_8160,N_7176,N_7369);
nand U8161 (N_8161,N_7221,N_7063);
nand U8162 (N_8162,N_7993,N_7799);
xor U8163 (N_8163,N_7563,N_7264);
or U8164 (N_8164,N_7655,N_7180);
and U8165 (N_8165,N_7323,N_7352);
nand U8166 (N_8166,N_7556,N_7508);
and U8167 (N_8167,N_7057,N_7581);
nand U8168 (N_8168,N_7014,N_7671);
xnor U8169 (N_8169,N_7564,N_7478);
nor U8170 (N_8170,N_7999,N_7857);
and U8171 (N_8171,N_7414,N_7418);
xor U8172 (N_8172,N_7422,N_7200);
nand U8173 (N_8173,N_7467,N_7839);
nand U8174 (N_8174,N_7521,N_7310);
nand U8175 (N_8175,N_7088,N_7184);
or U8176 (N_8176,N_7495,N_7796);
nor U8177 (N_8177,N_7913,N_7764);
or U8178 (N_8178,N_7782,N_7253);
nand U8179 (N_8179,N_7688,N_7106);
nor U8180 (N_8180,N_7198,N_7980);
or U8181 (N_8181,N_7986,N_7610);
nand U8182 (N_8182,N_7017,N_7509);
and U8183 (N_8183,N_7457,N_7619);
nor U8184 (N_8184,N_7842,N_7759);
or U8185 (N_8185,N_7875,N_7314);
nand U8186 (N_8186,N_7914,N_7976);
xnor U8187 (N_8187,N_7044,N_7437);
and U8188 (N_8188,N_7451,N_7149);
nand U8189 (N_8189,N_7386,N_7196);
and U8190 (N_8190,N_7215,N_7727);
or U8191 (N_8191,N_7983,N_7726);
or U8192 (N_8192,N_7544,N_7649);
nor U8193 (N_8193,N_7711,N_7287);
or U8194 (N_8194,N_7628,N_7255);
and U8195 (N_8195,N_7466,N_7420);
xor U8196 (N_8196,N_7878,N_7128);
xnor U8197 (N_8197,N_7309,N_7399);
or U8198 (N_8198,N_7562,N_7864);
xnor U8199 (N_8199,N_7579,N_7516);
or U8200 (N_8200,N_7262,N_7218);
nand U8201 (N_8201,N_7197,N_7332);
or U8202 (N_8202,N_7476,N_7858);
nand U8203 (N_8203,N_7429,N_7800);
xnor U8204 (N_8204,N_7558,N_7886);
xor U8205 (N_8205,N_7675,N_7103);
nor U8206 (N_8206,N_7364,N_7245);
nor U8207 (N_8207,N_7366,N_7390);
nand U8208 (N_8208,N_7716,N_7949);
or U8209 (N_8209,N_7458,N_7817);
and U8210 (N_8210,N_7929,N_7441);
xnor U8211 (N_8211,N_7313,N_7389);
nor U8212 (N_8212,N_7135,N_7667);
xor U8213 (N_8213,N_7674,N_7058);
xor U8214 (N_8214,N_7820,N_7303);
nor U8215 (N_8215,N_7708,N_7479);
nor U8216 (N_8216,N_7233,N_7879);
or U8217 (N_8217,N_7647,N_7571);
or U8218 (N_8218,N_7528,N_7566);
nand U8219 (N_8219,N_7347,N_7046);
xnor U8220 (N_8220,N_7616,N_7728);
nand U8221 (N_8221,N_7472,N_7555);
nand U8222 (N_8222,N_7075,N_7433);
or U8223 (N_8223,N_7311,N_7710);
and U8224 (N_8224,N_7806,N_7580);
nor U8225 (N_8225,N_7367,N_7713);
or U8226 (N_8226,N_7279,N_7056);
or U8227 (N_8227,N_7078,N_7318);
or U8228 (N_8228,N_7226,N_7639);
nand U8229 (N_8229,N_7635,N_7007);
nand U8230 (N_8230,N_7109,N_7193);
xor U8231 (N_8231,N_7632,N_7165);
or U8232 (N_8232,N_7153,N_7788);
nor U8233 (N_8233,N_7599,N_7426);
and U8234 (N_8234,N_7320,N_7112);
or U8235 (N_8235,N_7372,N_7851);
nor U8236 (N_8236,N_7702,N_7957);
xnor U8237 (N_8237,N_7552,N_7285);
nor U8238 (N_8238,N_7964,N_7974);
or U8239 (N_8239,N_7319,N_7623);
and U8240 (N_8240,N_7920,N_7867);
and U8241 (N_8241,N_7417,N_7236);
or U8242 (N_8242,N_7908,N_7561);
or U8243 (N_8243,N_7248,N_7652);
xor U8244 (N_8244,N_7356,N_7880);
nor U8245 (N_8245,N_7425,N_7603);
nand U8246 (N_8246,N_7994,N_7814);
and U8247 (N_8247,N_7606,N_7470);
xnor U8248 (N_8248,N_7442,N_7979);
nand U8249 (N_8249,N_7387,N_7807);
or U8250 (N_8250,N_7308,N_7092);
or U8251 (N_8251,N_7115,N_7973);
or U8252 (N_8252,N_7268,N_7411);
xnor U8253 (N_8253,N_7480,N_7186);
nand U8254 (N_8254,N_7455,N_7397);
or U8255 (N_8255,N_7912,N_7037);
or U8256 (N_8256,N_7083,N_7520);
or U8257 (N_8257,N_7413,N_7996);
and U8258 (N_8258,N_7931,N_7125);
and U8259 (N_8259,N_7750,N_7294);
and U8260 (N_8260,N_7790,N_7038);
nor U8261 (N_8261,N_7270,N_7093);
nand U8262 (N_8262,N_7523,N_7721);
and U8263 (N_8263,N_7346,N_7859);
nor U8264 (N_8264,N_7150,N_7770);
nand U8265 (N_8265,N_7605,N_7107);
and U8266 (N_8266,N_7554,N_7328);
or U8267 (N_8267,N_7910,N_7316);
xnor U8268 (N_8268,N_7371,N_7187);
and U8269 (N_8269,N_7202,N_7132);
xnor U8270 (N_8270,N_7199,N_7402);
nand U8271 (N_8271,N_7586,N_7395);
nand U8272 (N_8272,N_7612,N_7435);
and U8273 (N_8273,N_7840,N_7971);
nand U8274 (N_8274,N_7843,N_7359);
or U8275 (N_8275,N_7407,N_7342);
nand U8276 (N_8276,N_7684,N_7448);
or U8277 (N_8277,N_7909,N_7173);
nor U8278 (N_8278,N_7627,N_7876);
nand U8279 (N_8279,N_7054,N_7237);
xnor U8280 (N_8280,N_7614,N_7847);
nand U8281 (N_8281,N_7163,N_7967);
and U8282 (N_8282,N_7915,N_7290);
nor U8283 (N_8283,N_7076,N_7746);
nor U8284 (N_8284,N_7838,N_7720);
nand U8285 (N_8285,N_7499,N_7234);
nand U8286 (N_8286,N_7701,N_7844);
nor U8287 (N_8287,N_7464,N_7636);
nand U8288 (N_8288,N_7870,N_7074);
xor U8289 (N_8289,N_7777,N_7136);
nor U8290 (N_8290,N_7217,N_7535);
and U8291 (N_8291,N_7201,N_7690);
xnor U8292 (N_8292,N_7855,N_7775);
nor U8293 (N_8293,N_7622,N_7831);
xnor U8294 (N_8294,N_7680,N_7216);
xor U8295 (N_8295,N_7496,N_7032);
and U8296 (N_8296,N_7804,N_7664);
and U8297 (N_8297,N_7219,N_7436);
nand U8298 (N_8298,N_7744,N_7385);
nor U8299 (N_8299,N_7988,N_7911);
nand U8300 (N_8300,N_7207,N_7856);
or U8301 (N_8301,N_7064,N_7517);
nor U8302 (N_8302,N_7203,N_7019);
xnor U8303 (N_8303,N_7224,N_7712);
or U8304 (N_8304,N_7731,N_7656);
xor U8305 (N_8305,N_7934,N_7423);
xnor U8306 (N_8306,N_7404,N_7918);
xnor U8307 (N_8307,N_7578,N_7511);
xor U8308 (N_8308,N_7190,N_7662);
and U8309 (N_8309,N_7665,N_7829);
nor U8310 (N_8310,N_7343,N_7345);
or U8311 (N_8311,N_7515,N_7134);
xnor U8312 (N_8312,N_7928,N_7760);
nor U8313 (N_8313,N_7257,N_7593);
nor U8314 (N_8314,N_7145,N_7178);
nand U8315 (N_8315,N_7491,N_7208);
and U8316 (N_8316,N_7531,N_7751);
nor U8317 (N_8317,N_7592,N_7975);
nor U8318 (N_8318,N_7784,N_7659);
or U8319 (N_8319,N_7242,N_7123);
nor U8320 (N_8320,N_7363,N_7933);
or U8321 (N_8321,N_7557,N_7238);
nor U8322 (N_8322,N_7953,N_7355);
nor U8323 (N_8323,N_7755,N_7302);
nand U8324 (N_8324,N_7171,N_7298);
nor U8325 (N_8325,N_7565,N_7765);
xnor U8326 (N_8326,N_7272,N_7590);
nand U8327 (N_8327,N_7130,N_7009);
nor U8328 (N_8328,N_7111,N_7862);
and U8329 (N_8329,N_7925,N_7668);
xor U8330 (N_8330,N_7379,N_7985);
or U8331 (N_8331,N_7089,N_7572);
nor U8332 (N_8332,N_7672,N_7917);
and U8333 (N_8333,N_7835,N_7944);
and U8334 (N_8334,N_7452,N_7474);
and U8335 (N_8335,N_7781,N_7697);
nor U8336 (N_8336,N_7740,N_7837);
nand U8337 (N_8337,N_7039,N_7600);
nand U8338 (N_8338,N_7191,N_7065);
or U8339 (N_8339,N_7645,N_7432);
or U8340 (N_8340,N_7182,N_7335);
xnor U8341 (N_8341,N_7569,N_7893);
nor U8342 (N_8342,N_7175,N_7589);
nand U8343 (N_8343,N_7803,N_7036);
or U8344 (N_8344,N_7613,N_7887);
nor U8345 (N_8345,N_7660,N_7300);
and U8346 (N_8346,N_7071,N_7923);
nand U8347 (N_8347,N_7401,N_7018);
and U8348 (N_8348,N_7995,N_7338);
nand U8349 (N_8349,N_7483,N_7597);
nor U8350 (N_8350,N_7368,N_7049);
nor U8351 (N_8351,N_7329,N_7276);
nor U8352 (N_8352,N_7991,N_7551);
and U8353 (N_8353,N_7882,N_7514);
xnor U8354 (N_8354,N_7798,N_7885);
nor U8355 (N_8355,N_7841,N_7576);
nand U8356 (N_8356,N_7846,N_7596);
or U8357 (N_8357,N_7438,N_7383);
nand U8358 (N_8358,N_7482,N_7365);
nor U8359 (N_8359,N_7830,N_7468);
nor U8360 (N_8360,N_7340,N_7753);
xor U8361 (N_8361,N_7696,N_7067);
or U8362 (N_8362,N_7948,N_7286);
and U8363 (N_8363,N_7881,N_7724);
and U8364 (N_8364,N_7440,N_7225);
nor U8365 (N_8365,N_7567,N_7997);
xor U8366 (N_8366,N_7631,N_7896);
or U8367 (N_8367,N_7119,N_7102);
nor U8368 (N_8368,N_7575,N_7958);
and U8369 (N_8369,N_7658,N_7382);
nor U8370 (N_8370,N_7742,N_7027);
nor U8371 (N_8371,N_7942,N_7070);
or U8372 (N_8372,N_7982,N_7801);
or U8373 (N_8373,N_7260,N_7274);
and U8374 (N_8374,N_7488,N_7170);
nor U8375 (N_8375,N_7000,N_7042);
nor U8376 (N_8376,N_7296,N_7683);
xor U8377 (N_8377,N_7052,N_7456);
nand U8378 (N_8378,N_7443,N_7783);
or U8379 (N_8379,N_7079,N_7016);
or U8380 (N_8380,N_7194,N_7434);
xor U8381 (N_8381,N_7406,N_7963);
or U8382 (N_8382,N_7732,N_7970);
and U8383 (N_8383,N_7836,N_7348);
xnor U8384 (N_8384,N_7428,N_7232);
or U8385 (N_8385,N_7729,N_7815);
or U8386 (N_8386,N_7462,N_7860);
and U8387 (N_8387,N_7504,N_7715);
nand U8388 (N_8388,N_7334,N_7943);
xor U8389 (N_8389,N_7415,N_7022);
and U8390 (N_8390,N_7120,N_7412);
nand U8391 (N_8391,N_7725,N_7604);
or U8392 (N_8392,N_7518,N_7358);
nor U8393 (N_8393,N_7213,N_7646);
or U8394 (N_8394,N_7403,N_7869);
and U8395 (N_8395,N_7874,N_7312);
and U8396 (N_8396,N_7935,N_7493);
or U8397 (N_8397,N_7322,N_7952);
nor U8398 (N_8398,N_7460,N_7825);
or U8399 (N_8399,N_7289,N_7924);
nand U8400 (N_8400,N_7393,N_7082);
or U8401 (N_8401,N_7618,N_7734);
nor U8402 (N_8402,N_7277,N_7707);
and U8403 (N_8403,N_7703,N_7827);
and U8404 (N_8404,N_7325,N_7588);
nor U8405 (N_8405,N_7167,N_7169);
nand U8406 (N_8406,N_7972,N_7738);
xor U8407 (N_8407,N_7350,N_7861);
nand U8408 (N_8408,N_7757,N_7143);
xnor U8409 (N_8409,N_7029,N_7522);
or U8410 (N_8410,N_7327,N_7945);
nor U8411 (N_8411,N_7865,N_7954);
and U8412 (N_8412,N_7549,N_7743);
nand U8413 (N_8413,N_7431,N_7086);
and U8414 (N_8414,N_7489,N_7899);
nor U8415 (N_8415,N_7685,N_7471);
xnor U8416 (N_8416,N_7693,N_7981);
nand U8417 (N_8417,N_7124,N_7863);
nand U8418 (N_8418,N_7608,N_7375);
nor U8419 (N_8419,N_7723,N_7377);
or U8420 (N_8420,N_7583,N_7941);
and U8421 (N_8421,N_7370,N_7848);
nor U8422 (N_8422,N_7040,N_7240);
nor U8423 (N_8423,N_7717,N_7061);
and U8424 (N_8424,N_7177,N_7398);
xor U8425 (N_8425,N_7758,N_7542);
nand U8426 (N_8426,N_7845,N_7529);
or U8427 (N_8427,N_7214,N_7152);
and U8428 (N_8428,N_7154,N_7637);
and U8429 (N_8429,N_7810,N_7259);
or U8430 (N_8430,N_7901,N_7231);
nor U8431 (N_8431,N_7331,N_7114);
and U8432 (N_8432,N_7357,N_7081);
nor U8433 (N_8433,N_7852,N_7465);
and U8434 (N_8434,N_7621,N_7210);
nand U8435 (N_8435,N_7767,N_7354);
nand U8436 (N_8436,N_7873,N_7940);
xnor U8437 (N_8437,N_7249,N_7205);
nor U8438 (N_8438,N_7756,N_7883);
or U8439 (N_8439,N_7699,N_7121);
xor U8440 (N_8440,N_7722,N_7011);
nand U8441 (N_8441,N_7768,N_7633);
nand U8442 (N_8442,N_7373,N_7545);
xor U8443 (N_8443,N_7189,N_7192);
nand U8444 (N_8444,N_7247,N_7530);
nor U8445 (N_8445,N_7947,N_7681);
or U8446 (N_8446,N_7737,N_7138);
xor U8447 (N_8447,N_7956,N_7694);
nand U8448 (N_8448,N_7396,N_7004);
and U8449 (N_8449,N_7888,N_7292);
nand U8450 (N_8450,N_7897,N_7349);
nor U8451 (N_8451,N_7261,N_7718);
xor U8452 (N_8452,N_7536,N_7748);
and U8453 (N_8453,N_7161,N_7959);
xor U8454 (N_8454,N_7624,N_7251);
or U8455 (N_8455,N_7669,N_7243);
or U8456 (N_8456,N_7244,N_7962);
and U8457 (N_8457,N_7792,N_7113);
xnor U8458 (N_8458,N_7118,N_7281);
nor U8459 (N_8459,N_7689,N_7188);
or U8460 (N_8460,N_7156,N_7209);
xnor U8461 (N_8461,N_7271,N_7394);
xnor U8462 (N_8462,N_7498,N_7144);
and U8463 (N_8463,N_7473,N_7360);
nand U8464 (N_8464,N_7235,N_7100);
or U8465 (N_8465,N_7024,N_7813);
nor U8466 (N_8466,N_7537,N_7503);
nand U8467 (N_8467,N_7692,N_7644);
or U8468 (N_8468,N_7927,N_7087);
xor U8469 (N_8469,N_7676,N_7634);
xnor U8470 (N_8470,N_7045,N_7745);
nor U8471 (N_8471,N_7704,N_7591);
nand U8472 (N_8472,N_7391,N_7108);
nor U8473 (N_8473,N_7961,N_7602);
xor U8474 (N_8474,N_7299,N_7889);
or U8475 (N_8475,N_7033,N_7771);
xor U8476 (N_8476,N_7388,N_7650);
or U8477 (N_8477,N_7866,N_7091);
or U8478 (N_8478,N_7094,N_7185);
xor U8479 (N_8479,N_7050,N_7453);
nor U8480 (N_8480,N_7028,N_7006);
or U8481 (N_8481,N_7263,N_7305);
xor U8482 (N_8482,N_7824,N_7101);
and U8483 (N_8483,N_7582,N_7906);
or U8484 (N_8484,N_7682,N_7099);
xnor U8485 (N_8485,N_7601,N_7459);
and U8486 (N_8486,N_7513,N_7041);
and U8487 (N_8487,N_7105,N_7212);
and U8488 (N_8488,N_7663,N_7691);
nor U8489 (N_8489,N_7805,N_7337);
and U8490 (N_8490,N_7902,N_7904);
and U8491 (N_8491,N_7625,N_7648);
or U8492 (N_8492,N_7073,N_7630);
xnor U8493 (N_8493,N_7220,N_7430);
nand U8494 (N_8494,N_7550,N_7297);
or U8495 (N_8495,N_7376,N_7761);
xnor U8496 (N_8496,N_7547,N_7450);
nor U8497 (N_8497,N_7955,N_7519);
nand U8498 (N_8498,N_7965,N_7405);
xnor U8499 (N_8499,N_7424,N_7148);
nor U8500 (N_8500,N_7276,N_7664);
and U8501 (N_8501,N_7519,N_7444);
xor U8502 (N_8502,N_7574,N_7449);
nand U8503 (N_8503,N_7112,N_7372);
xor U8504 (N_8504,N_7181,N_7906);
and U8505 (N_8505,N_7425,N_7459);
or U8506 (N_8506,N_7243,N_7867);
nor U8507 (N_8507,N_7172,N_7797);
or U8508 (N_8508,N_7454,N_7460);
and U8509 (N_8509,N_7640,N_7118);
xor U8510 (N_8510,N_7579,N_7561);
nor U8511 (N_8511,N_7967,N_7335);
nand U8512 (N_8512,N_7642,N_7363);
nor U8513 (N_8513,N_7908,N_7881);
nand U8514 (N_8514,N_7616,N_7684);
nand U8515 (N_8515,N_7234,N_7646);
or U8516 (N_8516,N_7588,N_7799);
and U8517 (N_8517,N_7102,N_7802);
nor U8518 (N_8518,N_7174,N_7270);
and U8519 (N_8519,N_7606,N_7471);
xnor U8520 (N_8520,N_7171,N_7516);
or U8521 (N_8521,N_7959,N_7776);
xnor U8522 (N_8522,N_7419,N_7516);
xnor U8523 (N_8523,N_7180,N_7979);
and U8524 (N_8524,N_7406,N_7068);
or U8525 (N_8525,N_7373,N_7333);
nor U8526 (N_8526,N_7757,N_7298);
or U8527 (N_8527,N_7008,N_7315);
nor U8528 (N_8528,N_7160,N_7910);
or U8529 (N_8529,N_7618,N_7557);
or U8530 (N_8530,N_7978,N_7446);
and U8531 (N_8531,N_7618,N_7154);
xor U8532 (N_8532,N_7538,N_7541);
nor U8533 (N_8533,N_7158,N_7175);
nand U8534 (N_8534,N_7579,N_7270);
and U8535 (N_8535,N_7918,N_7871);
nand U8536 (N_8536,N_7514,N_7184);
or U8537 (N_8537,N_7017,N_7137);
or U8538 (N_8538,N_7723,N_7976);
nor U8539 (N_8539,N_7835,N_7533);
or U8540 (N_8540,N_7271,N_7436);
nand U8541 (N_8541,N_7884,N_7327);
nand U8542 (N_8542,N_7033,N_7133);
and U8543 (N_8543,N_7230,N_7309);
and U8544 (N_8544,N_7663,N_7464);
and U8545 (N_8545,N_7659,N_7954);
xnor U8546 (N_8546,N_7901,N_7408);
xnor U8547 (N_8547,N_7449,N_7211);
xnor U8548 (N_8548,N_7374,N_7732);
nor U8549 (N_8549,N_7943,N_7059);
or U8550 (N_8550,N_7980,N_7928);
nand U8551 (N_8551,N_7677,N_7307);
or U8552 (N_8552,N_7395,N_7172);
nor U8553 (N_8553,N_7662,N_7122);
nor U8554 (N_8554,N_7529,N_7418);
and U8555 (N_8555,N_7810,N_7657);
nand U8556 (N_8556,N_7901,N_7735);
nor U8557 (N_8557,N_7570,N_7441);
or U8558 (N_8558,N_7506,N_7283);
and U8559 (N_8559,N_7496,N_7220);
and U8560 (N_8560,N_7218,N_7704);
xnor U8561 (N_8561,N_7880,N_7425);
nor U8562 (N_8562,N_7622,N_7959);
nand U8563 (N_8563,N_7352,N_7119);
or U8564 (N_8564,N_7355,N_7352);
nor U8565 (N_8565,N_7709,N_7773);
nor U8566 (N_8566,N_7975,N_7268);
and U8567 (N_8567,N_7014,N_7186);
and U8568 (N_8568,N_7113,N_7753);
xor U8569 (N_8569,N_7383,N_7878);
or U8570 (N_8570,N_7195,N_7101);
and U8571 (N_8571,N_7551,N_7568);
nor U8572 (N_8572,N_7227,N_7708);
or U8573 (N_8573,N_7326,N_7301);
nand U8574 (N_8574,N_7911,N_7530);
or U8575 (N_8575,N_7015,N_7461);
and U8576 (N_8576,N_7120,N_7747);
or U8577 (N_8577,N_7588,N_7219);
xnor U8578 (N_8578,N_7403,N_7633);
nand U8579 (N_8579,N_7985,N_7544);
nand U8580 (N_8580,N_7094,N_7402);
nand U8581 (N_8581,N_7925,N_7073);
nor U8582 (N_8582,N_7045,N_7495);
xnor U8583 (N_8583,N_7781,N_7549);
and U8584 (N_8584,N_7532,N_7499);
or U8585 (N_8585,N_7120,N_7165);
nor U8586 (N_8586,N_7320,N_7820);
nand U8587 (N_8587,N_7674,N_7323);
and U8588 (N_8588,N_7988,N_7826);
and U8589 (N_8589,N_7953,N_7185);
nand U8590 (N_8590,N_7098,N_7259);
nor U8591 (N_8591,N_7051,N_7421);
and U8592 (N_8592,N_7768,N_7990);
nor U8593 (N_8593,N_7405,N_7095);
or U8594 (N_8594,N_7057,N_7476);
xnor U8595 (N_8595,N_7517,N_7521);
xnor U8596 (N_8596,N_7592,N_7769);
nor U8597 (N_8597,N_7828,N_7843);
nor U8598 (N_8598,N_7763,N_7751);
xnor U8599 (N_8599,N_7621,N_7895);
nand U8600 (N_8600,N_7674,N_7409);
nor U8601 (N_8601,N_7050,N_7068);
nor U8602 (N_8602,N_7313,N_7209);
xor U8603 (N_8603,N_7781,N_7134);
nand U8604 (N_8604,N_7975,N_7871);
nand U8605 (N_8605,N_7349,N_7771);
nand U8606 (N_8606,N_7557,N_7434);
nor U8607 (N_8607,N_7456,N_7028);
xnor U8608 (N_8608,N_7437,N_7345);
and U8609 (N_8609,N_7709,N_7256);
xnor U8610 (N_8610,N_7180,N_7752);
xor U8611 (N_8611,N_7389,N_7898);
nand U8612 (N_8612,N_7553,N_7929);
nor U8613 (N_8613,N_7267,N_7661);
and U8614 (N_8614,N_7712,N_7801);
or U8615 (N_8615,N_7046,N_7391);
nor U8616 (N_8616,N_7982,N_7358);
xnor U8617 (N_8617,N_7488,N_7760);
xnor U8618 (N_8618,N_7171,N_7816);
or U8619 (N_8619,N_7681,N_7282);
nand U8620 (N_8620,N_7262,N_7886);
or U8621 (N_8621,N_7437,N_7499);
and U8622 (N_8622,N_7201,N_7212);
nor U8623 (N_8623,N_7577,N_7536);
and U8624 (N_8624,N_7608,N_7514);
nand U8625 (N_8625,N_7726,N_7624);
nor U8626 (N_8626,N_7031,N_7371);
and U8627 (N_8627,N_7109,N_7818);
nand U8628 (N_8628,N_7942,N_7517);
nand U8629 (N_8629,N_7393,N_7028);
and U8630 (N_8630,N_7744,N_7008);
xor U8631 (N_8631,N_7969,N_7147);
and U8632 (N_8632,N_7576,N_7971);
or U8633 (N_8633,N_7753,N_7763);
xor U8634 (N_8634,N_7450,N_7776);
xnor U8635 (N_8635,N_7099,N_7275);
nor U8636 (N_8636,N_7625,N_7417);
or U8637 (N_8637,N_7489,N_7786);
xor U8638 (N_8638,N_7967,N_7525);
nand U8639 (N_8639,N_7973,N_7165);
nor U8640 (N_8640,N_7818,N_7126);
and U8641 (N_8641,N_7533,N_7075);
or U8642 (N_8642,N_7314,N_7059);
nor U8643 (N_8643,N_7785,N_7568);
or U8644 (N_8644,N_7690,N_7746);
nand U8645 (N_8645,N_7154,N_7920);
nor U8646 (N_8646,N_7191,N_7657);
xnor U8647 (N_8647,N_7508,N_7384);
nor U8648 (N_8648,N_7481,N_7484);
and U8649 (N_8649,N_7430,N_7980);
xnor U8650 (N_8650,N_7355,N_7425);
and U8651 (N_8651,N_7529,N_7803);
or U8652 (N_8652,N_7559,N_7767);
or U8653 (N_8653,N_7463,N_7697);
nand U8654 (N_8654,N_7204,N_7458);
or U8655 (N_8655,N_7372,N_7266);
or U8656 (N_8656,N_7572,N_7381);
and U8657 (N_8657,N_7790,N_7069);
xnor U8658 (N_8658,N_7825,N_7651);
or U8659 (N_8659,N_7661,N_7515);
and U8660 (N_8660,N_7307,N_7054);
nand U8661 (N_8661,N_7289,N_7685);
or U8662 (N_8662,N_7185,N_7044);
nand U8663 (N_8663,N_7852,N_7265);
or U8664 (N_8664,N_7062,N_7532);
and U8665 (N_8665,N_7883,N_7754);
xor U8666 (N_8666,N_7676,N_7049);
nand U8667 (N_8667,N_7777,N_7235);
and U8668 (N_8668,N_7225,N_7095);
nand U8669 (N_8669,N_7776,N_7111);
xor U8670 (N_8670,N_7614,N_7795);
xnor U8671 (N_8671,N_7905,N_7998);
nand U8672 (N_8672,N_7275,N_7589);
xnor U8673 (N_8673,N_7135,N_7515);
nand U8674 (N_8674,N_7082,N_7067);
nor U8675 (N_8675,N_7697,N_7851);
or U8676 (N_8676,N_7145,N_7665);
nand U8677 (N_8677,N_7377,N_7179);
or U8678 (N_8678,N_7388,N_7364);
and U8679 (N_8679,N_7755,N_7293);
and U8680 (N_8680,N_7403,N_7400);
xnor U8681 (N_8681,N_7015,N_7984);
nor U8682 (N_8682,N_7300,N_7450);
xor U8683 (N_8683,N_7849,N_7988);
xor U8684 (N_8684,N_7990,N_7550);
xnor U8685 (N_8685,N_7421,N_7745);
or U8686 (N_8686,N_7533,N_7128);
or U8687 (N_8687,N_7349,N_7373);
and U8688 (N_8688,N_7589,N_7818);
nand U8689 (N_8689,N_7143,N_7479);
and U8690 (N_8690,N_7911,N_7870);
and U8691 (N_8691,N_7975,N_7556);
xnor U8692 (N_8692,N_7972,N_7959);
nand U8693 (N_8693,N_7982,N_7612);
nand U8694 (N_8694,N_7156,N_7816);
nor U8695 (N_8695,N_7258,N_7101);
xor U8696 (N_8696,N_7875,N_7113);
nor U8697 (N_8697,N_7236,N_7665);
nand U8698 (N_8698,N_7804,N_7513);
and U8699 (N_8699,N_7878,N_7570);
xnor U8700 (N_8700,N_7922,N_7108);
or U8701 (N_8701,N_7783,N_7298);
nand U8702 (N_8702,N_7142,N_7961);
nor U8703 (N_8703,N_7519,N_7246);
and U8704 (N_8704,N_7581,N_7505);
xnor U8705 (N_8705,N_7658,N_7109);
nor U8706 (N_8706,N_7104,N_7644);
xnor U8707 (N_8707,N_7519,N_7862);
and U8708 (N_8708,N_7927,N_7641);
nand U8709 (N_8709,N_7733,N_7438);
xor U8710 (N_8710,N_7436,N_7429);
and U8711 (N_8711,N_7066,N_7833);
nor U8712 (N_8712,N_7931,N_7650);
nand U8713 (N_8713,N_7304,N_7760);
nor U8714 (N_8714,N_7416,N_7785);
and U8715 (N_8715,N_7586,N_7869);
and U8716 (N_8716,N_7559,N_7462);
and U8717 (N_8717,N_7793,N_7399);
nor U8718 (N_8718,N_7445,N_7990);
xor U8719 (N_8719,N_7860,N_7638);
nor U8720 (N_8720,N_7589,N_7932);
and U8721 (N_8721,N_7906,N_7162);
nand U8722 (N_8722,N_7479,N_7491);
and U8723 (N_8723,N_7102,N_7871);
nand U8724 (N_8724,N_7564,N_7947);
xor U8725 (N_8725,N_7518,N_7499);
or U8726 (N_8726,N_7145,N_7766);
nor U8727 (N_8727,N_7226,N_7352);
and U8728 (N_8728,N_7670,N_7027);
and U8729 (N_8729,N_7721,N_7580);
or U8730 (N_8730,N_7715,N_7912);
xor U8731 (N_8731,N_7384,N_7981);
or U8732 (N_8732,N_7769,N_7604);
xor U8733 (N_8733,N_7034,N_7179);
and U8734 (N_8734,N_7940,N_7100);
or U8735 (N_8735,N_7894,N_7875);
or U8736 (N_8736,N_7911,N_7859);
xor U8737 (N_8737,N_7324,N_7500);
and U8738 (N_8738,N_7489,N_7164);
or U8739 (N_8739,N_7623,N_7585);
or U8740 (N_8740,N_7105,N_7113);
xor U8741 (N_8741,N_7309,N_7043);
or U8742 (N_8742,N_7090,N_7011);
and U8743 (N_8743,N_7154,N_7823);
nand U8744 (N_8744,N_7869,N_7881);
nand U8745 (N_8745,N_7605,N_7330);
nor U8746 (N_8746,N_7218,N_7580);
or U8747 (N_8747,N_7110,N_7202);
xor U8748 (N_8748,N_7282,N_7213);
xor U8749 (N_8749,N_7455,N_7609);
nor U8750 (N_8750,N_7825,N_7174);
or U8751 (N_8751,N_7024,N_7925);
nand U8752 (N_8752,N_7531,N_7183);
nand U8753 (N_8753,N_7944,N_7811);
nand U8754 (N_8754,N_7873,N_7881);
nand U8755 (N_8755,N_7976,N_7043);
nor U8756 (N_8756,N_7715,N_7964);
nor U8757 (N_8757,N_7647,N_7234);
xor U8758 (N_8758,N_7902,N_7973);
and U8759 (N_8759,N_7507,N_7184);
or U8760 (N_8760,N_7592,N_7299);
or U8761 (N_8761,N_7310,N_7935);
xor U8762 (N_8762,N_7521,N_7718);
and U8763 (N_8763,N_7502,N_7920);
nor U8764 (N_8764,N_7760,N_7179);
nor U8765 (N_8765,N_7646,N_7522);
or U8766 (N_8766,N_7071,N_7520);
nand U8767 (N_8767,N_7027,N_7017);
xor U8768 (N_8768,N_7530,N_7696);
or U8769 (N_8769,N_7440,N_7053);
or U8770 (N_8770,N_7029,N_7333);
or U8771 (N_8771,N_7155,N_7245);
nand U8772 (N_8772,N_7339,N_7448);
and U8773 (N_8773,N_7931,N_7875);
nor U8774 (N_8774,N_7131,N_7768);
xor U8775 (N_8775,N_7655,N_7899);
nor U8776 (N_8776,N_7013,N_7133);
nor U8777 (N_8777,N_7530,N_7451);
nand U8778 (N_8778,N_7978,N_7661);
and U8779 (N_8779,N_7262,N_7540);
nor U8780 (N_8780,N_7105,N_7758);
xor U8781 (N_8781,N_7266,N_7073);
nand U8782 (N_8782,N_7051,N_7510);
and U8783 (N_8783,N_7662,N_7069);
and U8784 (N_8784,N_7083,N_7512);
nor U8785 (N_8785,N_7144,N_7045);
nand U8786 (N_8786,N_7323,N_7555);
xor U8787 (N_8787,N_7580,N_7197);
xor U8788 (N_8788,N_7657,N_7626);
or U8789 (N_8789,N_7514,N_7991);
and U8790 (N_8790,N_7788,N_7290);
or U8791 (N_8791,N_7725,N_7698);
xnor U8792 (N_8792,N_7518,N_7040);
and U8793 (N_8793,N_7423,N_7300);
xor U8794 (N_8794,N_7185,N_7354);
and U8795 (N_8795,N_7478,N_7833);
or U8796 (N_8796,N_7357,N_7167);
nand U8797 (N_8797,N_7840,N_7071);
and U8798 (N_8798,N_7330,N_7407);
nor U8799 (N_8799,N_7412,N_7707);
or U8800 (N_8800,N_7637,N_7476);
and U8801 (N_8801,N_7711,N_7821);
nor U8802 (N_8802,N_7064,N_7172);
nor U8803 (N_8803,N_7646,N_7335);
xor U8804 (N_8804,N_7675,N_7071);
or U8805 (N_8805,N_7664,N_7481);
nand U8806 (N_8806,N_7728,N_7096);
or U8807 (N_8807,N_7629,N_7836);
nor U8808 (N_8808,N_7273,N_7991);
nand U8809 (N_8809,N_7379,N_7879);
nor U8810 (N_8810,N_7914,N_7784);
and U8811 (N_8811,N_7306,N_7024);
or U8812 (N_8812,N_7504,N_7052);
xnor U8813 (N_8813,N_7289,N_7630);
and U8814 (N_8814,N_7264,N_7868);
or U8815 (N_8815,N_7461,N_7634);
xnor U8816 (N_8816,N_7881,N_7947);
or U8817 (N_8817,N_7623,N_7897);
and U8818 (N_8818,N_7901,N_7906);
or U8819 (N_8819,N_7375,N_7396);
xor U8820 (N_8820,N_7302,N_7724);
nor U8821 (N_8821,N_7925,N_7086);
nand U8822 (N_8822,N_7624,N_7559);
and U8823 (N_8823,N_7224,N_7973);
and U8824 (N_8824,N_7916,N_7696);
nand U8825 (N_8825,N_7399,N_7083);
nand U8826 (N_8826,N_7157,N_7669);
nor U8827 (N_8827,N_7802,N_7996);
nor U8828 (N_8828,N_7788,N_7754);
and U8829 (N_8829,N_7926,N_7928);
and U8830 (N_8830,N_7769,N_7764);
nand U8831 (N_8831,N_7947,N_7318);
nand U8832 (N_8832,N_7552,N_7043);
nor U8833 (N_8833,N_7239,N_7569);
or U8834 (N_8834,N_7640,N_7322);
or U8835 (N_8835,N_7929,N_7889);
nand U8836 (N_8836,N_7544,N_7764);
nand U8837 (N_8837,N_7603,N_7205);
xor U8838 (N_8838,N_7372,N_7748);
or U8839 (N_8839,N_7696,N_7279);
nand U8840 (N_8840,N_7057,N_7020);
nand U8841 (N_8841,N_7856,N_7047);
xor U8842 (N_8842,N_7251,N_7034);
and U8843 (N_8843,N_7895,N_7491);
nor U8844 (N_8844,N_7674,N_7729);
nand U8845 (N_8845,N_7650,N_7850);
and U8846 (N_8846,N_7888,N_7965);
nand U8847 (N_8847,N_7167,N_7729);
nand U8848 (N_8848,N_7802,N_7709);
and U8849 (N_8849,N_7434,N_7828);
nor U8850 (N_8850,N_7281,N_7484);
nor U8851 (N_8851,N_7717,N_7914);
xor U8852 (N_8852,N_7519,N_7311);
and U8853 (N_8853,N_7981,N_7235);
nor U8854 (N_8854,N_7321,N_7695);
or U8855 (N_8855,N_7663,N_7888);
or U8856 (N_8856,N_7946,N_7008);
nand U8857 (N_8857,N_7442,N_7891);
and U8858 (N_8858,N_7214,N_7278);
xnor U8859 (N_8859,N_7534,N_7160);
xnor U8860 (N_8860,N_7657,N_7298);
or U8861 (N_8861,N_7230,N_7356);
and U8862 (N_8862,N_7499,N_7597);
nor U8863 (N_8863,N_7518,N_7384);
nand U8864 (N_8864,N_7022,N_7641);
or U8865 (N_8865,N_7858,N_7067);
and U8866 (N_8866,N_7182,N_7038);
and U8867 (N_8867,N_7672,N_7549);
nand U8868 (N_8868,N_7873,N_7161);
nand U8869 (N_8869,N_7682,N_7514);
or U8870 (N_8870,N_7496,N_7186);
nand U8871 (N_8871,N_7941,N_7968);
xor U8872 (N_8872,N_7304,N_7614);
or U8873 (N_8873,N_7950,N_7032);
and U8874 (N_8874,N_7198,N_7748);
and U8875 (N_8875,N_7608,N_7239);
xor U8876 (N_8876,N_7102,N_7844);
nor U8877 (N_8877,N_7208,N_7630);
or U8878 (N_8878,N_7751,N_7212);
or U8879 (N_8879,N_7628,N_7035);
nand U8880 (N_8880,N_7324,N_7149);
nor U8881 (N_8881,N_7592,N_7153);
nand U8882 (N_8882,N_7160,N_7911);
nor U8883 (N_8883,N_7827,N_7514);
or U8884 (N_8884,N_7742,N_7561);
nor U8885 (N_8885,N_7224,N_7418);
xor U8886 (N_8886,N_7436,N_7614);
nor U8887 (N_8887,N_7376,N_7129);
xor U8888 (N_8888,N_7612,N_7551);
nor U8889 (N_8889,N_7352,N_7302);
and U8890 (N_8890,N_7434,N_7573);
or U8891 (N_8891,N_7465,N_7587);
nand U8892 (N_8892,N_7155,N_7293);
nor U8893 (N_8893,N_7018,N_7319);
xor U8894 (N_8894,N_7536,N_7795);
nor U8895 (N_8895,N_7371,N_7618);
xnor U8896 (N_8896,N_7098,N_7494);
nand U8897 (N_8897,N_7758,N_7541);
nand U8898 (N_8898,N_7125,N_7382);
nand U8899 (N_8899,N_7089,N_7055);
nand U8900 (N_8900,N_7781,N_7077);
or U8901 (N_8901,N_7972,N_7486);
xor U8902 (N_8902,N_7362,N_7456);
or U8903 (N_8903,N_7304,N_7286);
xor U8904 (N_8904,N_7836,N_7522);
nor U8905 (N_8905,N_7655,N_7916);
nand U8906 (N_8906,N_7498,N_7199);
and U8907 (N_8907,N_7326,N_7840);
xnor U8908 (N_8908,N_7407,N_7552);
nand U8909 (N_8909,N_7798,N_7199);
nand U8910 (N_8910,N_7652,N_7556);
and U8911 (N_8911,N_7936,N_7347);
or U8912 (N_8912,N_7141,N_7019);
nand U8913 (N_8913,N_7272,N_7393);
nand U8914 (N_8914,N_7943,N_7081);
nand U8915 (N_8915,N_7757,N_7495);
nand U8916 (N_8916,N_7655,N_7501);
nor U8917 (N_8917,N_7272,N_7142);
nand U8918 (N_8918,N_7357,N_7201);
or U8919 (N_8919,N_7843,N_7291);
nand U8920 (N_8920,N_7161,N_7173);
nor U8921 (N_8921,N_7773,N_7441);
nand U8922 (N_8922,N_7754,N_7640);
nand U8923 (N_8923,N_7907,N_7416);
nor U8924 (N_8924,N_7259,N_7741);
xnor U8925 (N_8925,N_7290,N_7299);
xnor U8926 (N_8926,N_7023,N_7903);
or U8927 (N_8927,N_7224,N_7184);
or U8928 (N_8928,N_7421,N_7785);
or U8929 (N_8929,N_7360,N_7855);
nor U8930 (N_8930,N_7112,N_7886);
nor U8931 (N_8931,N_7624,N_7131);
or U8932 (N_8932,N_7991,N_7518);
xor U8933 (N_8933,N_7467,N_7309);
xor U8934 (N_8934,N_7610,N_7316);
xor U8935 (N_8935,N_7397,N_7407);
xnor U8936 (N_8936,N_7481,N_7029);
or U8937 (N_8937,N_7603,N_7559);
and U8938 (N_8938,N_7022,N_7001);
nor U8939 (N_8939,N_7735,N_7825);
and U8940 (N_8940,N_7015,N_7965);
and U8941 (N_8941,N_7229,N_7728);
nand U8942 (N_8942,N_7588,N_7270);
nand U8943 (N_8943,N_7719,N_7354);
or U8944 (N_8944,N_7742,N_7941);
nor U8945 (N_8945,N_7138,N_7238);
xor U8946 (N_8946,N_7659,N_7206);
nand U8947 (N_8947,N_7277,N_7615);
and U8948 (N_8948,N_7517,N_7658);
nand U8949 (N_8949,N_7976,N_7546);
nand U8950 (N_8950,N_7515,N_7489);
and U8951 (N_8951,N_7359,N_7284);
nand U8952 (N_8952,N_7794,N_7712);
or U8953 (N_8953,N_7926,N_7764);
and U8954 (N_8954,N_7789,N_7839);
nand U8955 (N_8955,N_7933,N_7975);
xor U8956 (N_8956,N_7507,N_7818);
nand U8957 (N_8957,N_7995,N_7247);
or U8958 (N_8958,N_7774,N_7181);
and U8959 (N_8959,N_7742,N_7335);
or U8960 (N_8960,N_7937,N_7218);
nor U8961 (N_8961,N_7861,N_7541);
nand U8962 (N_8962,N_7914,N_7175);
and U8963 (N_8963,N_7339,N_7887);
nor U8964 (N_8964,N_7932,N_7619);
or U8965 (N_8965,N_7250,N_7572);
xor U8966 (N_8966,N_7847,N_7290);
xnor U8967 (N_8967,N_7595,N_7212);
nand U8968 (N_8968,N_7938,N_7126);
nor U8969 (N_8969,N_7697,N_7181);
or U8970 (N_8970,N_7115,N_7084);
nand U8971 (N_8971,N_7614,N_7287);
nand U8972 (N_8972,N_7669,N_7495);
nor U8973 (N_8973,N_7951,N_7442);
nand U8974 (N_8974,N_7301,N_7620);
nand U8975 (N_8975,N_7134,N_7500);
and U8976 (N_8976,N_7089,N_7544);
nor U8977 (N_8977,N_7873,N_7770);
nand U8978 (N_8978,N_7210,N_7441);
nand U8979 (N_8979,N_7832,N_7532);
nor U8980 (N_8980,N_7417,N_7970);
and U8981 (N_8981,N_7576,N_7544);
nand U8982 (N_8982,N_7701,N_7419);
nor U8983 (N_8983,N_7440,N_7286);
nor U8984 (N_8984,N_7355,N_7846);
and U8985 (N_8985,N_7832,N_7123);
nand U8986 (N_8986,N_7260,N_7001);
and U8987 (N_8987,N_7591,N_7547);
or U8988 (N_8988,N_7219,N_7650);
and U8989 (N_8989,N_7461,N_7395);
or U8990 (N_8990,N_7897,N_7974);
nor U8991 (N_8991,N_7789,N_7503);
nor U8992 (N_8992,N_7019,N_7356);
xor U8993 (N_8993,N_7021,N_7813);
or U8994 (N_8994,N_7988,N_7767);
or U8995 (N_8995,N_7829,N_7876);
or U8996 (N_8996,N_7780,N_7359);
nor U8997 (N_8997,N_7042,N_7156);
or U8998 (N_8998,N_7983,N_7949);
and U8999 (N_8999,N_7251,N_7235);
xor U9000 (N_9000,N_8896,N_8783);
or U9001 (N_9001,N_8170,N_8611);
nor U9002 (N_9002,N_8181,N_8395);
or U9003 (N_9003,N_8668,N_8087);
nand U9004 (N_9004,N_8810,N_8563);
and U9005 (N_9005,N_8126,N_8808);
and U9006 (N_9006,N_8275,N_8415);
or U9007 (N_9007,N_8665,N_8912);
xor U9008 (N_9008,N_8632,N_8554);
nor U9009 (N_9009,N_8673,N_8357);
xor U9010 (N_9010,N_8319,N_8637);
or U9011 (N_9011,N_8648,N_8515);
or U9012 (N_9012,N_8557,N_8830);
and U9013 (N_9013,N_8393,N_8477);
nand U9014 (N_9014,N_8725,N_8151);
and U9015 (N_9015,N_8465,N_8754);
nor U9016 (N_9016,N_8659,N_8696);
nand U9017 (N_9017,N_8268,N_8813);
and U9018 (N_9018,N_8821,N_8675);
and U9019 (N_9019,N_8689,N_8840);
nor U9020 (N_9020,N_8957,N_8748);
xnor U9021 (N_9021,N_8186,N_8054);
nor U9022 (N_9022,N_8401,N_8392);
nor U9023 (N_9023,N_8372,N_8095);
xor U9024 (N_9024,N_8751,N_8092);
nand U9025 (N_9025,N_8997,N_8968);
xor U9026 (N_9026,N_8291,N_8025);
nand U9027 (N_9027,N_8592,N_8738);
nor U9028 (N_9028,N_8265,N_8380);
and U9029 (N_9029,N_8405,N_8327);
and U9030 (N_9030,N_8773,N_8888);
nor U9031 (N_9031,N_8114,N_8222);
nand U9032 (N_9032,N_8692,N_8003);
or U9033 (N_9033,N_8883,N_8556);
xnor U9034 (N_9034,N_8449,N_8103);
and U9035 (N_9035,N_8086,N_8803);
nand U9036 (N_9036,N_8278,N_8424);
xnor U9037 (N_9037,N_8919,N_8490);
nand U9038 (N_9038,N_8132,N_8743);
nor U9039 (N_9039,N_8476,N_8062);
nor U9040 (N_9040,N_8300,N_8261);
nand U9041 (N_9041,N_8289,N_8038);
and U9042 (N_9042,N_8165,N_8464);
nand U9043 (N_9043,N_8493,N_8811);
xnor U9044 (N_9044,N_8963,N_8468);
xnor U9045 (N_9045,N_8544,N_8273);
xor U9046 (N_9046,N_8138,N_8863);
nor U9047 (N_9047,N_8658,N_8566);
nand U9048 (N_9048,N_8943,N_8995);
nor U9049 (N_9049,N_8982,N_8535);
nor U9050 (N_9050,N_8894,N_8647);
nand U9051 (N_9051,N_8175,N_8364);
nand U9052 (N_9052,N_8721,N_8428);
xnor U9053 (N_9053,N_8009,N_8026);
or U9054 (N_9054,N_8891,N_8441);
or U9055 (N_9055,N_8605,N_8260);
xor U9056 (N_9056,N_8055,N_8010);
or U9057 (N_9057,N_8510,N_8924);
nand U9058 (N_9058,N_8407,N_8248);
nor U9059 (N_9059,N_8644,N_8501);
nand U9060 (N_9060,N_8686,N_8683);
and U9061 (N_9061,N_8005,N_8693);
nand U9062 (N_9062,N_8500,N_8100);
nor U9063 (N_9063,N_8842,N_8817);
or U9064 (N_9064,N_8416,N_8741);
xnor U9065 (N_9065,N_8506,N_8908);
nor U9066 (N_9066,N_8189,N_8917);
xnor U9067 (N_9067,N_8885,N_8220);
nor U9068 (N_9068,N_8340,N_8074);
nand U9069 (N_9069,N_8561,N_8097);
nand U9070 (N_9070,N_8367,N_8844);
nor U9071 (N_9071,N_8984,N_8002);
and U9072 (N_9072,N_8128,N_8240);
xor U9073 (N_9073,N_8085,N_8656);
or U9074 (N_9074,N_8358,N_8767);
nand U9075 (N_9075,N_8244,N_8871);
or U9076 (N_9076,N_8410,N_8606);
nor U9077 (N_9077,N_8852,N_8022);
or U9078 (N_9078,N_8524,N_8188);
nor U9079 (N_9079,N_8270,N_8429);
or U9080 (N_9080,N_8909,N_8564);
xnor U9081 (N_9081,N_8112,N_8223);
xnor U9082 (N_9082,N_8547,N_8569);
xnor U9083 (N_9083,N_8672,N_8822);
xnor U9084 (N_9084,N_8595,N_8843);
nor U9085 (N_9085,N_8150,N_8450);
nor U9086 (N_9086,N_8483,N_8518);
nor U9087 (N_9087,N_8215,N_8430);
or U9088 (N_9088,N_8120,N_8122);
or U9089 (N_9089,N_8812,N_8080);
or U9090 (N_9090,N_8172,N_8516);
and U9091 (N_9091,N_8245,N_8800);
nor U9092 (N_9092,N_8777,N_8230);
and U9093 (N_9093,N_8940,N_8243);
nand U9094 (N_9094,N_8333,N_8434);
nand U9095 (N_9095,N_8373,N_8107);
xor U9096 (N_9096,N_8104,N_8938);
xnor U9097 (N_9097,N_8178,N_8084);
xnor U9098 (N_9098,N_8484,N_8666);
and U9099 (N_9099,N_8109,N_8035);
nand U9100 (N_9100,N_8682,N_8847);
nor U9101 (N_9101,N_8155,N_8412);
and U9102 (N_9102,N_8130,N_8988);
nor U9103 (N_9103,N_8839,N_8201);
or U9104 (N_9104,N_8024,N_8798);
nand U9105 (N_9105,N_8902,N_8949);
and U9106 (N_9106,N_8855,N_8713);
nand U9107 (N_9107,N_8528,N_8915);
xor U9108 (N_9108,N_8323,N_8717);
nand U9109 (N_9109,N_8094,N_8420);
nor U9110 (N_9110,N_8562,N_8599);
nor U9111 (N_9111,N_8200,N_8694);
or U9112 (N_9112,N_8508,N_8971);
xor U9113 (N_9113,N_8772,N_8481);
nor U9114 (N_9114,N_8046,N_8900);
or U9115 (N_9115,N_8073,N_8755);
xor U9116 (N_9116,N_8318,N_8571);
xor U9117 (N_9117,N_8377,N_8942);
nand U9118 (N_9118,N_8704,N_8118);
nand U9119 (N_9119,N_8457,N_8498);
xnor U9120 (N_9120,N_8050,N_8448);
nor U9121 (N_9121,N_8669,N_8173);
nand U9122 (N_9122,N_8676,N_8347);
nor U9123 (N_9123,N_8198,N_8731);
xor U9124 (N_9124,N_8332,N_8487);
xnor U9125 (N_9125,N_8509,N_8570);
and U9126 (N_9126,N_8017,N_8491);
xnor U9127 (N_9127,N_8296,N_8343);
xor U9128 (N_9128,N_8989,N_8496);
nor U9129 (N_9129,N_8784,N_8145);
nor U9130 (N_9130,N_8388,N_8264);
and U9131 (N_9131,N_8633,N_8030);
nor U9132 (N_9132,N_8306,N_8207);
nand U9133 (N_9133,N_8786,N_8670);
nand U9134 (N_9134,N_8687,N_8579);
xnor U9135 (N_9135,N_8023,N_8251);
nor U9136 (N_9136,N_8652,N_8685);
xnor U9137 (N_9137,N_8252,N_8060);
or U9138 (N_9138,N_8397,N_8106);
and U9139 (N_9139,N_8931,N_8801);
nand U9140 (N_9140,N_8019,N_8699);
or U9141 (N_9141,N_8444,N_8432);
nand U9142 (N_9142,N_8714,N_8044);
xor U9143 (N_9143,N_8753,N_8301);
nor U9144 (N_9144,N_8948,N_8070);
or U9145 (N_9145,N_8763,N_8622);
and U9146 (N_9146,N_8654,N_8905);
nand U9147 (N_9147,N_8258,N_8646);
nor U9148 (N_9148,N_8629,N_8199);
nor U9149 (N_9149,N_8361,N_8475);
nand U9150 (N_9150,N_8869,N_8585);
nor U9151 (N_9151,N_8166,N_8108);
nand U9152 (N_9152,N_8892,N_8697);
nand U9153 (N_9153,N_8951,N_8287);
and U9154 (N_9154,N_8954,N_8310);
or U9155 (N_9155,N_8495,N_8987);
nand U9156 (N_9156,N_8004,N_8276);
or U9157 (N_9157,N_8077,N_8964);
nand U9158 (N_9158,N_8488,N_8907);
nor U9159 (N_9159,N_8182,N_8423);
xor U9160 (N_9160,N_8775,N_8376);
and U9161 (N_9161,N_8848,N_8338);
nand U9162 (N_9162,N_8001,N_8521);
and U9163 (N_9163,N_8887,N_8121);
nor U9164 (N_9164,N_8959,N_8180);
nand U9165 (N_9165,N_8460,N_8572);
or U9166 (N_9166,N_8400,N_8131);
nor U9167 (N_9167,N_8433,N_8414);
nand U9168 (N_9168,N_8833,N_8255);
or U9169 (N_9169,N_8643,N_8136);
and U9170 (N_9170,N_8174,N_8816);
or U9171 (N_9171,N_8041,N_8337);
nor U9172 (N_9172,N_8870,N_8806);
and U9173 (N_9173,N_8443,N_8016);
nand U9174 (N_9174,N_8614,N_8679);
xor U9175 (N_9175,N_8079,N_8425);
xnor U9176 (N_9176,N_8911,N_8799);
or U9177 (N_9177,N_8246,N_8466);
xor U9178 (N_9178,N_8071,N_8582);
xor U9179 (N_9179,N_8978,N_8903);
or U9180 (N_9180,N_8913,N_8378);
nand U9181 (N_9181,N_8758,N_8729);
nand U9182 (N_9182,N_8101,N_8470);
nor U9183 (N_9183,N_8546,N_8661);
nor U9184 (N_9184,N_8083,N_8880);
or U9185 (N_9185,N_8053,N_8899);
and U9186 (N_9186,N_8774,N_8418);
xnor U9187 (N_9187,N_8156,N_8567);
and U9188 (N_9188,N_8574,N_8792);
or U9189 (N_9189,N_8761,N_8322);
and U9190 (N_9190,N_8630,N_8550);
or U9191 (N_9191,N_8163,N_8113);
and U9192 (N_9192,N_8921,N_8922);
xnor U9193 (N_9193,N_8727,N_8194);
xor U9194 (N_9194,N_8916,N_8720);
and U9195 (N_9195,N_8503,N_8304);
and U9196 (N_9196,N_8618,N_8785);
nand U9197 (N_9197,N_8527,N_8147);
and U9198 (N_9198,N_8820,N_8872);
nand U9199 (N_9199,N_8063,N_8797);
and U9200 (N_9200,N_8043,N_8625);
nand U9201 (N_9201,N_8012,N_8075);
and U9202 (N_9202,N_8970,N_8382);
nand U9203 (N_9203,N_8828,N_8355);
xnor U9204 (N_9204,N_8752,N_8297);
xnor U9205 (N_9205,N_8762,N_8048);
nor U9206 (N_9206,N_8531,N_8655);
xor U9207 (N_9207,N_8237,N_8231);
nor U9208 (N_9208,N_8235,N_8667);
nor U9209 (N_9209,N_8144,N_8294);
and U9210 (N_9210,N_8218,N_8967);
xnor U9211 (N_9211,N_8617,N_8953);
xnor U9212 (N_9212,N_8241,N_8233);
nand U9213 (N_9213,N_8375,N_8489);
or U9214 (N_9214,N_8525,N_8756);
and U9215 (N_9215,N_8209,N_8886);
xor U9216 (N_9216,N_8950,N_8853);
and U9217 (N_9217,N_8941,N_8417);
xor U9218 (N_9218,N_8650,N_8932);
xnor U9219 (N_9219,N_8387,N_8526);
nand U9220 (N_9220,N_8795,N_8134);
and U9221 (N_9221,N_8782,N_8250);
nor U9222 (N_9222,N_8153,N_8893);
and U9223 (N_9223,N_8735,N_8920);
and U9224 (N_9224,N_8143,N_8581);
xor U9225 (N_9225,N_8119,N_8836);
nor U9226 (N_9226,N_8623,N_8624);
and U9227 (N_9227,N_8316,N_8545);
nand U9228 (N_9228,N_8739,N_8286);
nand U9229 (N_9229,N_8018,N_8224);
nand U9230 (N_9230,N_8285,N_8141);
xor U9231 (N_9231,N_8292,N_8344);
and U9232 (N_9232,N_8615,N_8918);
and U9233 (N_9233,N_8446,N_8593);
xnor U9234 (N_9234,N_8972,N_8081);
xnor U9235 (N_9235,N_8356,N_8635);
and U9236 (N_9236,N_8733,N_8639);
and U9237 (N_9237,N_8945,N_8242);
and U9238 (N_9238,N_8602,N_8641);
nand U9239 (N_9239,N_8184,N_8402);
and U9240 (N_9240,N_8815,N_8052);
xor U9241 (N_9241,N_8159,N_8015);
and U9242 (N_9242,N_8396,N_8642);
and U9243 (N_9243,N_8703,N_8875);
nand U9244 (N_9244,N_8671,N_8616);
nand U9245 (N_9245,N_8860,N_8542);
and U9246 (N_9246,N_8927,N_8440);
xor U9247 (N_9247,N_8365,N_8031);
nand U9248 (N_9248,N_8190,N_8162);
or U9249 (N_9249,N_8790,N_8723);
xor U9250 (N_9250,N_8154,N_8776);
nor U9251 (N_9251,N_8631,N_8677);
xor U9252 (N_9252,N_8197,N_8975);
xnor U9253 (N_9253,N_8161,N_8539);
and U9254 (N_9254,N_8897,N_8834);
or U9255 (N_9255,N_8436,N_8827);
nor U9256 (N_9256,N_8099,N_8933);
xnor U9257 (N_9257,N_8791,N_8719);
nand U9258 (N_9258,N_8326,N_8311);
or U9259 (N_9259,N_8091,N_8486);
nor U9260 (N_9260,N_8926,N_8837);
nand U9261 (N_9261,N_8691,N_8479);
or U9262 (N_9262,N_8369,N_8601);
xnor U9263 (N_9263,N_8507,N_8923);
and U9264 (N_9264,N_8598,N_8711);
nand U9265 (N_9265,N_8504,N_8040);
or U9266 (N_9266,N_8341,N_8226);
or U9267 (N_9267,N_8505,N_8314);
or U9268 (N_9268,N_8657,N_8980);
nor U9269 (N_9269,N_8502,N_8051);
and U9270 (N_9270,N_8353,N_8459);
nand U9271 (N_9271,N_8330,N_8514);
xor U9272 (N_9272,N_8409,N_8014);
nand U9273 (N_9273,N_8740,N_8334);
nor U9274 (N_9274,N_8690,N_8193);
and U9275 (N_9275,N_8568,N_8110);
xnor U9276 (N_9276,N_8728,N_8320);
nor U9277 (N_9277,N_8914,N_8435);
xor U9278 (N_9278,N_8033,N_8447);
or U9279 (N_9279,N_8191,N_8594);
nand U9280 (N_9280,N_8851,N_8976);
nand U9281 (N_9281,N_8841,N_8823);
xnor U9282 (N_9282,N_8471,N_8536);
nand U9283 (N_9283,N_8331,N_8354);
and U9284 (N_9284,N_8455,N_8472);
and U9285 (N_9285,N_8196,N_8403);
and U9286 (N_9286,N_8497,N_8293);
nand U9287 (N_9287,N_8249,N_8346);
or U9288 (N_9288,N_8160,N_8478);
nor U9289 (N_9289,N_8882,N_8591);
and U9290 (N_9290,N_8212,N_8036);
nand U9291 (N_9291,N_8149,N_8283);
and U9292 (N_9292,N_8148,N_8700);
xnor U9293 (N_9293,N_8764,N_8499);
xor U9294 (N_9294,N_8047,N_8965);
xnor U9295 (N_9295,N_8530,N_8519);
xnor U9296 (N_9296,N_8638,N_8956);
nand U9297 (N_9297,N_8379,N_8575);
and U9298 (N_9298,N_8558,N_8398);
and U9299 (N_9299,N_8538,N_8442);
nand U9300 (N_9300,N_8688,N_8814);
or U9301 (N_9301,N_8759,N_8111);
and U9302 (N_9302,N_8467,N_8979);
xnor U9303 (N_9303,N_8211,N_8849);
nor U9304 (N_9304,N_8007,N_8494);
nor U9305 (N_9305,N_8187,N_8370);
nor U9306 (N_9306,N_8302,N_8826);
xor U9307 (N_9307,N_8277,N_8221);
or U9308 (N_9308,N_8889,N_8553);
nand U9309 (N_9309,N_8049,N_8303);
or U9310 (N_9310,N_8256,N_8000);
nand U9311 (N_9311,N_8308,N_8213);
nor U9312 (N_9312,N_8269,N_8645);
nand U9313 (N_9313,N_8279,N_8861);
xor U9314 (N_9314,N_8955,N_8802);
or U9315 (N_9315,N_8068,N_8431);
or U9316 (N_9316,N_8208,N_8267);
and U9317 (N_9317,N_8008,N_8192);
or U9318 (N_9318,N_8272,N_8088);
or U9319 (N_9319,N_8555,N_8288);
nor U9320 (N_9320,N_8227,N_8253);
nor U9321 (N_9321,N_8020,N_8426);
and U9322 (N_9322,N_8736,N_8098);
xor U9323 (N_9323,N_8996,N_8456);
and U9324 (N_9324,N_8280,N_8824);
nor U9325 (N_9325,N_8146,N_8168);
and U9326 (N_9326,N_8124,N_8925);
nor U9327 (N_9327,N_8082,N_8680);
and U9328 (N_9328,N_8698,N_8158);
xnor U9329 (N_9329,N_8974,N_8634);
nor U9330 (N_9330,N_8946,N_8307);
or U9331 (N_9331,N_8452,N_8363);
nand U9332 (N_9332,N_8877,N_8990);
and U9333 (N_9333,N_8281,N_8981);
nand U9334 (N_9334,N_8093,N_8474);
xor U9335 (N_9335,N_8734,N_8133);
and U9336 (N_9336,N_8749,N_8463);
xnor U9337 (N_9337,N_8072,N_8305);
and U9338 (N_9338,N_8710,N_8219);
and U9339 (N_9339,N_8983,N_8177);
or U9340 (N_9340,N_8708,N_8865);
nand U9341 (N_9341,N_8006,N_8766);
xnor U9342 (N_9342,N_8309,N_8993);
nor U9343 (N_9343,N_8804,N_8422);
or U9344 (N_9344,N_8588,N_8778);
xnor U9345 (N_9345,N_8236,N_8576);
nor U9346 (N_9346,N_8257,N_8262);
xnor U9347 (N_9347,N_8284,N_8862);
or U9348 (N_9348,N_8878,N_8712);
nand U9349 (N_9349,N_8716,N_8835);
or U9350 (N_9350,N_8511,N_8078);
nand U9351 (N_9351,N_8707,N_8684);
nor U9352 (N_9352,N_8724,N_8769);
xor U9353 (N_9353,N_8626,N_8930);
nor U9354 (N_9354,N_8850,N_8383);
or U9355 (N_9355,N_8747,N_8247);
nor U9356 (N_9356,N_8274,N_8421);
and U9357 (N_9357,N_8858,N_8389);
or U9358 (N_9358,N_8169,N_8117);
nand U9359 (N_9359,N_8868,N_8620);
nand U9360 (N_9360,N_8517,N_8540);
and U9361 (N_9361,N_8013,N_8884);
or U9362 (N_9362,N_8259,N_8064);
xor U9363 (N_9363,N_8619,N_8328);
and U9364 (N_9364,N_8454,N_8873);
and U9365 (N_9365,N_8335,N_8135);
nand U9366 (N_9366,N_8583,N_8578);
nand U9367 (N_9367,N_8042,N_8312);
and U9368 (N_9368,N_8368,N_8947);
xor U9369 (N_9369,N_8779,N_8404);
and U9370 (N_9370,N_8730,N_8898);
xnor U9371 (N_9371,N_8999,N_8139);
and U9372 (N_9372,N_8371,N_8204);
and U9373 (N_9373,N_8856,N_8966);
nor U9374 (N_9374,N_8028,N_8105);
or U9375 (N_9375,N_8298,N_8045);
xnor U9376 (N_9376,N_8552,N_8164);
nand U9377 (N_9377,N_8482,N_8998);
xnor U9378 (N_9378,N_8973,N_8351);
or U9379 (N_9379,N_8385,N_8548);
nand U9380 (N_9380,N_8329,N_8640);
xor U9381 (N_9381,N_8039,N_8610);
nor U9382 (N_9382,N_8458,N_8462);
and U9383 (N_9383,N_8750,N_8607);
nor U9384 (N_9384,N_8952,N_8934);
nand U9385 (N_9385,N_8928,N_8681);
or U9386 (N_9386,N_8621,N_8350);
nor U9387 (N_9387,N_8961,N_8202);
nand U9388 (N_9388,N_8857,N_8781);
nand U9389 (N_9389,N_8362,N_8746);
nand U9390 (N_9390,N_8890,N_8461);
or U9391 (N_9391,N_8573,N_8229);
xor U9392 (N_9392,N_8203,N_8076);
xor U9393 (N_9393,N_8701,N_8613);
and U9394 (N_9394,N_8176,N_8225);
nor U9395 (N_9395,N_8744,N_8879);
or U9396 (N_9396,N_8770,N_8771);
or U9397 (N_9397,N_8381,N_8768);
nand U9398 (N_9398,N_8867,N_8529);
nor U9399 (N_9399,N_8492,N_8485);
nand U9400 (N_9400,N_8254,N_8290);
xnor U9401 (N_9401,N_8663,N_8427);
and U9402 (N_9402,N_8451,N_8437);
and U9403 (N_9403,N_8239,N_8859);
and U9404 (N_9404,N_8939,N_8413);
or U9405 (N_9405,N_8394,N_8406);
nor U9406 (N_9406,N_8991,N_8805);
and U9407 (N_9407,N_8061,N_8419);
and U9408 (N_9408,N_8167,N_8994);
nand U9409 (N_9409,N_8709,N_8021);
xor U9410 (N_9410,N_8628,N_8185);
or U9411 (N_9411,N_8532,N_8807);
or U9412 (N_9412,N_8263,N_8513);
and U9413 (N_9413,N_8678,N_8090);
xnor U9414 (N_9414,N_8787,N_8793);
or U9415 (N_9415,N_8587,N_8216);
nand U9416 (N_9416,N_8818,N_8765);
nor U9417 (N_9417,N_8520,N_8011);
and U9418 (N_9418,N_8317,N_8969);
and U9419 (N_9419,N_8027,N_8349);
nand U9420 (N_9420,N_8608,N_8232);
nor U9421 (N_9421,N_8217,N_8565);
and U9422 (N_9422,N_8102,N_8559);
xor U9423 (N_9423,N_8958,N_8664);
nor U9424 (N_9424,N_8874,N_8066);
xor U9425 (N_9425,N_8390,N_8597);
xor U9426 (N_9426,N_8142,N_8876);
xnor U9427 (N_9427,N_8829,N_8152);
or U9428 (N_9428,N_8985,N_8904);
xnor U9429 (N_9429,N_8183,N_8195);
or U9430 (N_9430,N_8604,N_8819);
nor U9431 (N_9431,N_8705,N_8612);
or U9432 (N_9432,N_8069,N_8522);
nor U9433 (N_9433,N_8295,N_8937);
nor U9434 (N_9434,N_8864,N_8726);
nor U9435 (N_9435,N_8534,N_8742);
and U9436 (N_9436,N_8391,N_8551);
nand U9437 (N_9437,N_8649,N_8589);
and U9438 (N_9438,N_8137,N_8473);
nor U9439 (N_9439,N_8234,N_8116);
and U9440 (N_9440,N_8523,N_8936);
nor U9441 (N_9441,N_8127,N_8636);
and U9442 (N_9442,N_8386,N_8339);
and U9443 (N_9443,N_8760,N_8706);
nand U9444 (N_9444,N_8745,N_8342);
xnor U9445 (N_9445,N_8089,N_8321);
or U9446 (N_9446,N_8067,N_8935);
nand U9447 (N_9447,N_8282,N_8651);
nor U9448 (N_9448,N_8206,N_8171);
nand U9449 (N_9449,N_8838,N_8057);
or U9450 (N_9450,N_8123,N_8299);
or U9451 (N_9451,N_8205,N_8845);
xnor U9452 (N_9452,N_8129,N_8315);
xnor U9453 (N_9453,N_8214,N_8718);
xnor U9454 (N_9454,N_8832,N_8140);
nor U9455 (N_9455,N_8715,N_8702);
or U9456 (N_9456,N_8662,N_8266);
xnor U9457 (N_9457,N_8737,N_8157);
and U9458 (N_9458,N_8794,N_8453);
nand U9459 (N_9459,N_8596,N_8058);
nor U9460 (N_9460,N_8345,N_8895);
and U9461 (N_9461,N_8034,N_8929);
nand U9462 (N_9462,N_8992,N_8480);
and U9463 (N_9463,N_8584,N_8788);
or U9464 (N_9464,N_8059,N_8032);
and U9465 (N_9465,N_8469,N_8537);
nor U9466 (N_9466,N_8960,N_8037);
nand U9467 (N_9467,N_8512,N_8910);
nand U9468 (N_9468,N_8586,N_8445);
or U9469 (N_9469,N_8438,N_8881);
nand U9470 (N_9470,N_8348,N_8809);
xnor U9471 (N_9471,N_8541,N_8660);
and U9472 (N_9472,N_8825,N_8901);
or U9473 (N_9473,N_8796,N_8399);
or U9474 (N_9474,N_8352,N_8653);
nand U9475 (N_9475,N_8695,N_8580);
xnor U9476 (N_9476,N_8411,N_8210);
and U9477 (N_9477,N_8439,N_8271);
nand U9478 (N_9478,N_8366,N_8757);
nor U9479 (N_9479,N_8590,N_8609);
nor U9480 (N_9480,N_8179,N_8977);
or U9481 (N_9481,N_8780,N_8115);
xor U9482 (N_9482,N_8029,N_8238);
or U9483 (N_9483,N_8374,N_8384);
nor U9484 (N_9484,N_8962,N_8986);
nand U9485 (N_9485,N_8560,N_8722);
xor U9486 (N_9486,N_8854,N_8360);
and U9487 (N_9487,N_8627,N_8056);
and U9488 (N_9488,N_8228,N_8846);
or U9489 (N_9489,N_8577,N_8533);
and U9490 (N_9490,N_8789,N_8674);
xor U9491 (N_9491,N_8313,N_8096);
xnor U9492 (N_9492,N_8944,N_8359);
nor U9493 (N_9493,N_8065,N_8906);
xor U9494 (N_9494,N_8600,N_8125);
or U9495 (N_9495,N_8336,N_8549);
and U9496 (N_9496,N_8325,N_8831);
xor U9497 (N_9497,N_8866,N_8543);
nand U9498 (N_9498,N_8603,N_8324);
nand U9499 (N_9499,N_8408,N_8732);
nor U9500 (N_9500,N_8781,N_8375);
nor U9501 (N_9501,N_8846,N_8014);
nand U9502 (N_9502,N_8243,N_8258);
xor U9503 (N_9503,N_8538,N_8060);
xnor U9504 (N_9504,N_8299,N_8081);
xnor U9505 (N_9505,N_8248,N_8262);
and U9506 (N_9506,N_8419,N_8653);
and U9507 (N_9507,N_8854,N_8548);
nor U9508 (N_9508,N_8530,N_8382);
nand U9509 (N_9509,N_8236,N_8811);
nand U9510 (N_9510,N_8826,N_8655);
xor U9511 (N_9511,N_8558,N_8529);
nand U9512 (N_9512,N_8358,N_8046);
and U9513 (N_9513,N_8084,N_8324);
nor U9514 (N_9514,N_8026,N_8804);
or U9515 (N_9515,N_8312,N_8765);
xor U9516 (N_9516,N_8028,N_8557);
nand U9517 (N_9517,N_8252,N_8061);
nor U9518 (N_9518,N_8547,N_8261);
nand U9519 (N_9519,N_8197,N_8248);
xor U9520 (N_9520,N_8806,N_8872);
nor U9521 (N_9521,N_8633,N_8435);
or U9522 (N_9522,N_8813,N_8894);
nand U9523 (N_9523,N_8233,N_8680);
and U9524 (N_9524,N_8887,N_8024);
or U9525 (N_9525,N_8209,N_8166);
nor U9526 (N_9526,N_8155,N_8368);
nand U9527 (N_9527,N_8670,N_8391);
nor U9528 (N_9528,N_8729,N_8749);
and U9529 (N_9529,N_8634,N_8674);
or U9530 (N_9530,N_8592,N_8115);
nor U9531 (N_9531,N_8596,N_8152);
xor U9532 (N_9532,N_8174,N_8165);
or U9533 (N_9533,N_8463,N_8319);
and U9534 (N_9534,N_8449,N_8425);
or U9535 (N_9535,N_8758,N_8398);
nor U9536 (N_9536,N_8445,N_8425);
or U9537 (N_9537,N_8363,N_8880);
nand U9538 (N_9538,N_8316,N_8824);
nor U9539 (N_9539,N_8146,N_8936);
nor U9540 (N_9540,N_8003,N_8875);
xor U9541 (N_9541,N_8211,N_8367);
and U9542 (N_9542,N_8112,N_8887);
xor U9543 (N_9543,N_8515,N_8276);
and U9544 (N_9544,N_8842,N_8190);
or U9545 (N_9545,N_8538,N_8409);
and U9546 (N_9546,N_8825,N_8865);
and U9547 (N_9547,N_8566,N_8753);
nor U9548 (N_9548,N_8454,N_8785);
nor U9549 (N_9549,N_8058,N_8662);
and U9550 (N_9550,N_8946,N_8715);
nor U9551 (N_9551,N_8437,N_8998);
nor U9552 (N_9552,N_8864,N_8272);
xor U9553 (N_9553,N_8213,N_8686);
or U9554 (N_9554,N_8278,N_8617);
xnor U9555 (N_9555,N_8432,N_8237);
nand U9556 (N_9556,N_8710,N_8283);
and U9557 (N_9557,N_8277,N_8199);
nor U9558 (N_9558,N_8606,N_8739);
xnor U9559 (N_9559,N_8978,N_8151);
nor U9560 (N_9560,N_8173,N_8458);
xor U9561 (N_9561,N_8179,N_8289);
and U9562 (N_9562,N_8411,N_8955);
nand U9563 (N_9563,N_8614,N_8590);
or U9564 (N_9564,N_8949,N_8304);
nand U9565 (N_9565,N_8894,N_8261);
nor U9566 (N_9566,N_8374,N_8624);
and U9567 (N_9567,N_8036,N_8649);
and U9568 (N_9568,N_8663,N_8083);
and U9569 (N_9569,N_8626,N_8133);
nor U9570 (N_9570,N_8747,N_8050);
or U9571 (N_9571,N_8280,N_8230);
xnor U9572 (N_9572,N_8420,N_8005);
nand U9573 (N_9573,N_8925,N_8555);
and U9574 (N_9574,N_8963,N_8976);
and U9575 (N_9575,N_8637,N_8648);
nor U9576 (N_9576,N_8398,N_8348);
and U9577 (N_9577,N_8702,N_8881);
nor U9578 (N_9578,N_8914,N_8705);
nor U9579 (N_9579,N_8581,N_8738);
xnor U9580 (N_9580,N_8831,N_8797);
and U9581 (N_9581,N_8849,N_8087);
nor U9582 (N_9582,N_8237,N_8534);
or U9583 (N_9583,N_8546,N_8147);
nand U9584 (N_9584,N_8475,N_8880);
or U9585 (N_9585,N_8549,N_8808);
nand U9586 (N_9586,N_8416,N_8966);
nor U9587 (N_9587,N_8359,N_8089);
and U9588 (N_9588,N_8603,N_8645);
nand U9589 (N_9589,N_8599,N_8051);
or U9590 (N_9590,N_8455,N_8794);
and U9591 (N_9591,N_8664,N_8257);
nor U9592 (N_9592,N_8579,N_8868);
xor U9593 (N_9593,N_8556,N_8094);
and U9594 (N_9594,N_8579,N_8499);
nand U9595 (N_9595,N_8337,N_8823);
xor U9596 (N_9596,N_8808,N_8909);
and U9597 (N_9597,N_8381,N_8517);
and U9598 (N_9598,N_8159,N_8392);
nor U9599 (N_9599,N_8543,N_8912);
xor U9600 (N_9600,N_8691,N_8098);
nor U9601 (N_9601,N_8162,N_8158);
and U9602 (N_9602,N_8065,N_8291);
nor U9603 (N_9603,N_8737,N_8030);
or U9604 (N_9604,N_8165,N_8665);
or U9605 (N_9605,N_8249,N_8856);
and U9606 (N_9606,N_8623,N_8312);
or U9607 (N_9607,N_8056,N_8271);
xnor U9608 (N_9608,N_8525,N_8946);
and U9609 (N_9609,N_8725,N_8808);
and U9610 (N_9610,N_8483,N_8073);
xor U9611 (N_9611,N_8931,N_8720);
nor U9612 (N_9612,N_8122,N_8892);
nor U9613 (N_9613,N_8800,N_8199);
and U9614 (N_9614,N_8510,N_8391);
nor U9615 (N_9615,N_8966,N_8735);
nand U9616 (N_9616,N_8336,N_8571);
and U9617 (N_9617,N_8842,N_8346);
nor U9618 (N_9618,N_8381,N_8439);
or U9619 (N_9619,N_8840,N_8569);
nand U9620 (N_9620,N_8033,N_8905);
nor U9621 (N_9621,N_8967,N_8248);
xnor U9622 (N_9622,N_8186,N_8698);
and U9623 (N_9623,N_8493,N_8069);
or U9624 (N_9624,N_8294,N_8343);
xnor U9625 (N_9625,N_8728,N_8060);
and U9626 (N_9626,N_8241,N_8197);
nor U9627 (N_9627,N_8594,N_8643);
and U9628 (N_9628,N_8903,N_8317);
and U9629 (N_9629,N_8071,N_8276);
nor U9630 (N_9630,N_8765,N_8606);
or U9631 (N_9631,N_8534,N_8822);
or U9632 (N_9632,N_8887,N_8950);
and U9633 (N_9633,N_8450,N_8819);
or U9634 (N_9634,N_8173,N_8936);
and U9635 (N_9635,N_8023,N_8792);
nand U9636 (N_9636,N_8523,N_8632);
or U9637 (N_9637,N_8741,N_8774);
or U9638 (N_9638,N_8064,N_8888);
nand U9639 (N_9639,N_8945,N_8478);
and U9640 (N_9640,N_8405,N_8018);
xor U9641 (N_9641,N_8830,N_8136);
nand U9642 (N_9642,N_8098,N_8307);
or U9643 (N_9643,N_8398,N_8640);
xor U9644 (N_9644,N_8255,N_8611);
and U9645 (N_9645,N_8440,N_8960);
nor U9646 (N_9646,N_8415,N_8971);
nand U9647 (N_9647,N_8750,N_8473);
or U9648 (N_9648,N_8283,N_8440);
or U9649 (N_9649,N_8573,N_8585);
nor U9650 (N_9650,N_8839,N_8185);
xor U9651 (N_9651,N_8995,N_8883);
nand U9652 (N_9652,N_8102,N_8161);
nand U9653 (N_9653,N_8879,N_8968);
nand U9654 (N_9654,N_8284,N_8003);
nor U9655 (N_9655,N_8134,N_8325);
or U9656 (N_9656,N_8195,N_8602);
and U9657 (N_9657,N_8982,N_8147);
xnor U9658 (N_9658,N_8727,N_8333);
xor U9659 (N_9659,N_8691,N_8115);
and U9660 (N_9660,N_8818,N_8985);
nand U9661 (N_9661,N_8059,N_8004);
nand U9662 (N_9662,N_8880,N_8487);
and U9663 (N_9663,N_8640,N_8587);
or U9664 (N_9664,N_8303,N_8823);
nand U9665 (N_9665,N_8445,N_8616);
and U9666 (N_9666,N_8395,N_8940);
and U9667 (N_9667,N_8734,N_8880);
nor U9668 (N_9668,N_8784,N_8651);
and U9669 (N_9669,N_8669,N_8416);
xor U9670 (N_9670,N_8998,N_8371);
xnor U9671 (N_9671,N_8802,N_8611);
and U9672 (N_9672,N_8859,N_8823);
and U9673 (N_9673,N_8250,N_8603);
nor U9674 (N_9674,N_8421,N_8010);
and U9675 (N_9675,N_8759,N_8477);
nor U9676 (N_9676,N_8014,N_8090);
nand U9677 (N_9677,N_8335,N_8468);
or U9678 (N_9678,N_8706,N_8594);
or U9679 (N_9679,N_8171,N_8469);
nand U9680 (N_9680,N_8260,N_8689);
xor U9681 (N_9681,N_8509,N_8720);
or U9682 (N_9682,N_8663,N_8897);
xor U9683 (N_9683,N_8509,N_8013);
xor U9684 (N_9684,N_8506,N_8197);
and U9685 (N_9685,N_8992,N_8118);
or U9686 (N_9686,N_8750,N_8717);
and U9687 (N_9687,N_8964,N_8242);
nand U9688 (N_9688,N_8459,N_8633);
or U9689 (N_9689,N_8335,N_8294);
and U9690 (N_9690,N_8296,N_8247);
nand U9691 (N_9691,N_8097,N_8779);
and U9692 (N_9692,N_8465,N_8945);
and U9693 (N_9693,N_8821,N_8994);
or U9694 (N_9694,N_8774,N_8880);
nor U9695 (N_9695,N_8684,N_8887);
nor U9696 (N_9696,N_8025,N_8370);
nor U9697 (N_9697,N_8699,N_8897);
nand U9698 (N_9698,N_8991,N_8299);
xor U9699 (N_9699,N_8910,N_8566);
xor U9700 (N_9700,N_8122,N_8541);
nor U9701 (N_9701,N_8151,N_8192);
and U9702 (N_9702,N_8022,N_8887);
xor U9703 (N_9703,N_8934,N_8045);
and U9704 (N_9704,N_8562,N_8473);
and U9705 (N_9705,N_8018,N_8974);
nor U9706 (N_9706,N_8905,N_8093);
xnor U9707 (N_9707,N_8277,N_8603);
nor U9708 (N_9708,N_8107,N_8723);
nor U9709 (N_9709,N_8666,N_8878);
nand U9710 (N_9710,N_8176,N_8996);
nand U9711 (N_9711,N_8883,N_8492);
nor U9712 (N_9712,N_8062,N_8968);
nor U9713 (N_9713,N_8755,N_8391);
or U9714 (N_9714,N_8134,N_8801);
and U9715 (N_9715,N_8437,N_8504);
xor U9716 (N_9716,N_8337,N_8227);
or U9717 (N_9717,N_8477,N_8896);
nand U9718 (N_9718,N_8569,N_8990);
xor U9719 (N_9719,N_8584,N_8240);
xor U9720 (N_9720,N_8896,N_8530);
nand U9721 (N_9721,N_8196,N_8325);
or U9722 (N_9722,N_8761,N_8508);
xor U9723 (N_9723,N_8915,N_8499);
nor U9724 (N_9724,N_8248,N_8881);
and U9725 (N_9725,N_8716,N_8998);
xor U9726 (N_9726,N_8771,N_8667);
nor U9727 (N_9727,N_8304,N_8679);
or U9728 (N_9728,N_8106,N_8792);
xor U9729 (N_9729,N_8020,N_8058);
nor U9730 (N_9730,N_8231,N_8288);
nor U9731 (N_9731,N_8123,N_8196);
and U9732 (N_9732,N_8992,N_8918);
or U9733 (N_9733,N_8574,N_8130);
or U9734 (N_9734,N_8663,N_8593);
or U9735 (N_9735,N_8869,N_8848);
nor U9736 (N_9736,N_8425,N_8405);
nor U9737 (N_9737,N_8283,N_8988);
and U9738 (N_9738,N_8808,N_8239);
or U9739 (N_9739,N_8317,N_8746);
or U9740 (N_9740,N_8875,N_8991);
nand U9741 (N_9741,N_8936,N_8042);
and U9742 (N_9742,N_8051,N_8065);
nand U9743 (N_9743,N_8136,N_8277);
or U9744 (N_9744,N_8832,N_8934);
or U9745 (N_9745,N_8274,N_8304);
and U9746 (N_9746,N_8805,N_8664);
xor U9747 (N_9747,N_8373,N_8456);
xor U9748 (N_9748,N_8471,N_8191);
and U9749 (N_9749,N_8098,N_8442);
xnor U9750 (N_9750,N_8877,N_8288);
xnor U9751 (N_9751,N_8706,N_8973);
nand U9752 (N_9752,N_8460,N_8036);
or U9753 (N_9753,N_8565,N_8662);
and U9754 (N_9754,N_8112,N_8305);
nor U9755 (N_9755,N_8119,N_8674);
or U9756 (N_9756,N_8781,N_8250);
nand U9757 (N_9757,N_8743,N_8381);
or U9758 (N_9758,N_8122,N_8084);
xnor U9759 (N_9759,N_8523,N_8025);
nor U9760 (N_9760,N_8999,N_8395);
nor U9761 (N_9761,N_8952,N_8587);
nand U9762 (N_9762,N_8473,N_8604);
nand U9763 (N_9763,N_8514,N_8570);
nor U9764 (N_9764,N_8547,N_8439);
nor U9765 (N_9765,N_8043,N_8064);
and U9766 (N_9766,N_8457,N_8534);
nor U9767 (N_9767,N_8724,N_8039);
nor U9768 (N_9768,N_8106,N_8378);
and U9769 (N_9769,N_8255,N_8672);
xor U9770 (N_9770,N_8910,N_8155);
nand U9771 (N_9771,N_8193,N_8022);
or U9772 (N_9772,N_8787,N_8212);
nand U9773 (N_9773,N_8179,N_8600);
or U9774 (N_9774,N_8058,N_8642);
nand U9775 (N_9775,N_8187,N_8495);
and U9776 (N_9776,N_8077,N_8353);
or U9777 (N_9777,N_8889,N_8186);
and U9778 (N_9778,N_8416,N_8331);
nand U9779 (N_9779,N_8765,N_8644);
nor U9780 (N_9780,N_8821,N_8926);
nand U9781 (N_9781,N_8912,N_8608);
or U9782 (N_9782,N_8905,N_8424);
xnor U9783 (N_9783,N_8604,N_8270);
nand U9784 (N_9784,N_8975,N_8762);
and U9785 (N_9785,N_8582,N_8472);
xor U9786 (N_9786,N_8623,N_8055);
nor U9787 (N_9787,N_8545,N_8778);
xnor U9788 (N_9788,N_8501,N_8282);
and U9789 (N_9789,N_8962,N_8115);
nand U9790 (N_9790,N_8978,N_8952);
nand U9791 (N_9791,N_8580,N_8644);
nand U9792 (N_9792,N_8807,N_8571);
nor U9793 (N_9793,N_8522,N_8705);
nor U9794 (N_9794,N_8090,N_8704);
nand U9795 (N_9795,N_8216,N_8367);
nand U9796 (N_9796,N_8303,N_8196);
and U9797 (N_9797,N_8229,N_8079);
nand U9798 (N_9798,N_8823,N_8266);
nor U9799 (N_9799,N_8818,N_8740);
nor U9800 (N_9800,N_8650,N_8696);
and U9801 (N_9801,N_8705,N_8048);
nor U9802 (N_9802,N_8424,N_8889);
and U9803 (N_9803,N_8383,N_8984);
nand U9804 (N_9804,N_8005,N_8009);
and U9805 (N_9805,N_8655,N_8059);
xor U9806 (N_9806,N_8969,N_8356);
or U9807 (N_9807,N_8857,N_8293);
xor U9808 (N_9808,N_8133,N_8457);
nand U9809 (N_9809,N_8652,N_8348);
and U9810 (N_9810,N_8880,N_8020);
nor U9811 (N_9811,N_8123,N_8492);
or U9812 (N_9812,N_8316,N_8682);
xor U9813 (N_9813,N_8250,N_8692);
and U9814 (N_9814,N_8118,N_8230);
and U9815 (N_9815,N_8533,N_8300);
or U9816 (N_9816,N_8539,N_8477);
and U9817 (N_9817,N_8466,N_8268);
and U9818 (N_9818,N_8988,N_8275);
nor U9819 (N_9819,N_8508,N_8902);
and U9820 (N_9820,N_8342,N_8256);
nor U9821 (N_9821,N_8103,N_8044);
and U9822 (N_9822,N_8578,N_8600);
xor U9823 (N_9823,N_8919,N_8556);
and U9824 (N_9824,N_8405,N_8082);
nand U9825 (N_9825,N_8711,N_8133);
or U9826 (N_9826,N_8936,N_8577);
nor U9827 (N_9827,N_8657,N_8209);
or U9828 (N_9828,N_8003,N_8696);
and U9829 (N_9829,N_8199,N_8099);
and U9830 (N_9830,N_8522,N_8818);
nor U9831 (N_9831,N_8348,N_8619);
and U9832 (N_9832,N_8823,N_8348);
xor U9833 (N_9833,N_8800,N_8591);
nor U9834 (N_9834,N_8212,N_8325);
nand U9835 (N_9835,N_8289,N_8078);
xor U9836 (N_9836,N_8665,N_8055);
nand U9837 (N_9837,N_8627,N_8358);
nor U9838 (N_9838,N_8335,N_8964);
xnor U9839 (N_9839,N_8786,N_8158);
nand U9840 (N_9840,N_8547,N_8358);
or U9841 (N_9841,N_8492,N_8563);
nand U9842 (N_9842,N_8627,N_8212);
xor U9843 (N_9843,N_8565,N_8151);
and U9844 (N_9844,N_8273,N_8623);
nand U9845 (N_9845,N_8405,N_8756);
and U9846 (N_9846,N_8107,N_8272);
xnor U9847 (N_9847,N_8757,N_8247);
nand U9848 (N_9848,N_8669,N_8835);
and U9849 (N_9849,N_8407,N_8531);
nor U9850 (N_9850,N_8185,N_8369);
xor U9851 (N_9851,N_8603,N_8850);
xor U9852 (N_9852,N_8622,N_8047);
nand U9853 (N_9853,N_8784,N_8271);
xor U9854 (N_9854,N_8033,N_8242);
and U9855 (N_9855,N_8068,N_8644);
xnor U9856 (N_9856,N_8399,N_8617);
or U9857 (N_9857,N_8670,N_8971);
nand U9858 (N_9858,N_8312,N_8638);
and U9859 (N_9859,N_8970,N_8799);
and U9860 (N_9860,N_8142,N_8346);
nand U9861 (N_9861,N_8589,N_8725);
and U9862 (N_9862,N_8771,N_8181);
nand U9863 (N_9863,N_8670,N_8538);
nand U9864 (N_9864,N_8079,N_8226);
or U9865 (N_9865,N_8307,N_8897);
and U9866 (N_9866,N_8415,N_8577);
and U9867 (N_9867,N_8414,N_8920);
or U9868 (N_9868,N_8294,N_8575);
and U9869 (N_9869,N_8197,N_8480);
nor U9870 (N_9870,N_8859,N_8104);
xnor U9871 (N_9871,N_8104,N_8274);
nand U9872 (N_9872,N_8480,N_8472);
or U9873 (N_9873,N_8177,N_8999);
nand U9874 (N_9874,N_8048,N_8361);
nand U9875 (N_9875,N_8490,N_8405);
nand U9876 (N_9876,N_8160,N_8639);
xnor U9877 (N_9877,N_8238,N_8944);
nor U9878 (N_9878,N_8693,N_8841);
and U9879 (N_9879,N_8284,N_8447);
nand U9880 (N_9880,N_8579,N_8935);
and U9881 (N_9881,N_8791,N_8443);
xnor U9882 (N_9882,N_8719,N_8318);
or U9883 (N_9883,N_8622,N_8612);
or U9884 (N_9884,N_8738,N_8481);
nand U9885 (N_9885,N_8969,N_8917);
and U9886 (N_9886,N_8266,N_8599);
or U9887 (N_9887,N_8148,N_8697);
xnor U9888 (N_9888,N_8098,N_8785);
nand U9889 (N_9889,N_8582,N_8257);
or U9890 (N_9890,N_8534,N_8031);
nor U9891 (N_9891,N_8719,N_8245);
xnor U9892 (N_9892,N_8822,N_8973);
or U9893 (N_9893,N_8276,N_8030);
xnor U9894 (N_9894,N_8869,N_8922);
and U9895 (N_9895,N_8173,N_8175);
and U9896 (N_9896,N_8579,N_8083);
xor U9897 (N_9897,N_8327,N_8506);
nor U9898 (N_9898,N_8619,N_8699);
or U9899 (N_9899,N_8942,N_8738);
nor U9900 (N_9900,N_8565,N_8481);
xnor U9901 (N_9901,N_8507,N_8976);
nor U9902 (N_9902,N_8227,N_8268);
nor U9903 (N_9903,N_8024,N_8052);
nand U9904 (N_9904,N_8283,N_8704);
or U9905 (N_9905,N_8706,N_8641);
nand U9906 (N_9906,N_8512,N_8173);
and U9907 (N_9907,N_8706,N_8255);
nand U9908 (N_9908,N_8547,N_8290);
nor U9909 (N_9909,N_8950,N_8743);
or U9910 (N_9910,N_8792,N_8979);
and U9911 (N_9911,N_8522,N_8820);
and U9912 (N_9912,N_8996,N_8935);
or U9913 (N_9913,N_8631,N_8403);
nand U9914 (N_9914,N_8478,N_8352);
nor U9915 (N_9915,N_8501,N_8190);
nor U9916 (N_9916,N_8934,N_8847);
nor U9917 (N_9917,N_8214,N_8480);
or U9918 (N_9918,N_8065,N_8016);
nand U9919 (N_9919,N_8419,N_8027);
nand U9920 (N_9920,N_8362,N_8049);
and U9921 (N_9921,N_8351,N_8042);
nor U9922 (N_9922,N_8678,N_8826);
xor U9923 (N_9923,N_8378,N_8618);
and U9924 (N_9924,N_8473,N_8299);
nand U9925 (N_9925,N_8663,N_8122);
or U9926 (N_9926,N_8997,N_8653);
or U9927 (N_9927,N_8973,N_8281);
or U9928 (N_9928,N_8360,N_8897);
and U9929 (N_9929,N_8597,N_8078);
nand U9930 (N_9930,N_8018,N_8419);
nand U9931 (N_9931,N_8604,N_8632);
nand U9932 (N_9932,N_8022,N_8231);
xor U9933 (N_9933,N_8056,N_8939);
and U9934 (N_9934,N_8650,N_8706);
or U9935 (N_9935,N_8446,N_8826);
xnor U9936 (N_9936,N_8342,N_8617);
or U9937 (N_9937,N_8096,N_8029);
and U9938 (N_9938,N_8528,N_8106);
xnor U9939 (N_9939,N_8637,N_8933);
and U9940 (N_9940,N_8965,N_8467);
and U9941 (N_9941,N_8131,N_8743);
and U9942 (N_9942,N_8856,N_8333);
xnor U9943 (N_9943,N_8490,N_8246);
and U9944 (N_9944,N_8193,N_8276);
nor U9945 (N_9945,N_8261,N_8746);
nor U9946 (N_9946,N_8878,N_8174);
nand U9947 (N_9947,N_8549,N_8446);
nor U9948 (N_9948,N_8517,N_8356);
xnor U9949 (N_9949,N_8160,N_8116);
xnor U9950 (N_9950,N_8899,N_8534);
xor U9951 (N_9951,N_8162,N_8611);
or U9952 (N_9952,N_8870,N_8043);
or U9953 (N_9953,N_8523,N_8069);
xnor U9954 (N_9954,N_8405,N_8279);
nor U9955 (N_9955,N_8591,N_8732);
and U9956 (N_9956,N_8134,N_8649);
xor U9957 (N_9957,N_8112,N_8641);
or U9958 (N_9958,N_8235,N_8406);
and U9959 (N_9959,N_8606,N_8226);
xor U9960 (N_9960,N_8213,N_8867);
or U9961 (N_9961,N_8096,N_8624);
or U9962 (N_9962,N_8811,N_8448);
nand U9963 (N_9963,N_8769,N_8352);
nand U9964 (N_9964,N_8863,N_8734);
and U9965 (N_9965,N_8956,N_8658);
and U9966 (N_9966,N_8157,N_8353);
and U9967 (N_9967,N_8289,N_8761);
or U9968 (N_9968,N_8841,N_8521);
nor U9969 (N_9969,N_8385,N_8258);
and U9970 (N_9970,N_8375,N_8552);
xnor U9971 (N_9971,N_8711,N_8176);
and U9972 (N_9972,N_8600,N_8024);
and U9973 (N_9973,N_8272,N_8554);
or U9974 (N_9974,N_8106,N_8681);
nand U9975 (N_9975,N_8594,N_8532);
xnor U9976 (N_9976,N_8654,N_8746);
nor U9977 (N_9977,N_8205,N_8297);
nor U9978 (N_9978,N_8467,N_8953);
or U9979 (N_9979,N_8743,N_8402);
or U9980 (N_9980,N_8501,N_8240);
nor U9981 (N_9981,N_8469,N_8633);
and U9982 (N_9982,N_8643,N_8604);
or U9983 (N_9983,N_8460,N_8768);
nor U9984 (N_9984,N_8277,N_8536);
nand U9985 (N_9985,N_8116,N_8430);
nand U9986 (N_9986,N_8143,N_8813);
and U9987 (N_9987,N_8589,N_8419);
nor U9988 (N_9988,N_8077,N_8595);
nand U9989 (N_9989,N_8253,N_8286);
or U9990 (N_9990,N_8963,N_8995);
xor U9991 (N_9991,N_8680,N_8125);
nand U9992 (N_9992,N_8484,N_8383);
or U9993 (N_9993,N_8193,N_8318);
nand U9994 (N_9994,N_8774,N_8689);
or U9995 (N_9995,N_8227,N_8422);
and U9996 (N_9996,N_8844,N_8754);
nor U9997 (N_9997,N_8049,N_8889);
and U9998 (N_9998,N_8586,N_8829);
xor U9999 (N_9999,N_8278,N_8613);
and UO_0 (O_0,N_9784,N_9526);
xor UO_1 (O_1,N_9482,N_9453);
and UO_2 (O_2,N_9387,N_9576);
or UO_3 (O_3,N_9334,N_9016);
or UO_4 (O_4,N_9092,N_9851);
and UO_5 (O_5,N_9332,N_9008);
and UO_6 (O_6,N_9204,N_9376);
nor UO_7 (O_7,N_9281,N_9375);
or UO_8 (O_8,N_9998,N_9487);
or UO_9 (O_9,N_9400,N_9327);
nand UO_10 (O_10,N_9450,N_9781);
or UO_11 (O_11,N_9091,N_9255);
nand UO_12 (O_12,N_9074,N_9750);
and UO_13 (O_13,N_9904,N_9672);
xor UO_14 (O_14,N_9635,N_9017);
nor UO_15 (O_15,N_9059,N_9643);
nand UO_16 (O_16,N_9339,N_9166);
nand UO_17 (O_17,N_9201,N_9637);
xor UO_18 (O_18,N_9262,N_9593);
xor UO_19 (O_19,N_9795,N_9258);
xor UO_20 (O_20,N_9523,N_9289);
and UO_21 (O_21,N_9473,N_9377);
nand UO_22 (O_22,N_9514,N_9757);
and UO_23 (O_23,N_9737,N_9922);
and UO_24 (O_24,N_9032,N_9519);
nand UO_25 (O_25,N_9568,N_9597);
xnor UO_26 (O_26,N_9690,N_9290);
nor UO_27 (O_27,N_9251,N_9649);
or UO_28 (O_28,N_9942,N_9900);
and UO_29 (O_29,N_9037,N_9570);
nor UO_30 (O_30,N_9828,N_9476);
nor UO_31 (O_31,N_9411,N_9174);
nand UO_32 (O_32,N_9239,N_9625);
or UO_33 (O_33,N_9064,N_9391);
or UO_34 (O_34,N_9292,N_9536);
nor UO_35 (O_35,N_9312,N_9645);
nand UO_36 (O_36,N_9628,N_9596);
nand UO_37 (O_37,N_9126,N_9783);
and UO_38 (O_38,N_9704,N_9924);
or UO_39 (O_39,N_9427,N_9517);
xor UO_40 (O_40,N_9782,N_9002);
nor UO_41 (O_41,N_9322,N_9222);
or UO_42 (O_42,N_9124,N_9192);
xor UO_43 (O_43,N_9586,N_9865);
or UO_44 (O_44,N_9574,N_9972);
and UO_45 (O_45,N_9683,N_9238);
nor UO_46 (O_46,N_9849,N_9026);
nor UO_47 (O_47,N_9767,N_9793);
nand UO_48 (O_48,N_9565,N_9600);
and UO_49 (O_49,N_9745,N_9727);
nor UO_50 (O_50,N_9545,N_9345);
nand UO_51 (O_51,N_9320,N_9392);
nand UO_52 (O_52,N_9601,N_9956);
nand UO_53 (O_53,N_9451,N_9671);
and UO_54 (O_54,N_9491,N_9226);
and UO_55 (O_55,N_9522,N_9455);
and UO_56 (O_56,N_9532,N_9742);
nand UO_57 (O_57,N_9443,N_9558);
or UO_58 (O_58,N_9903,N_9407);
nor UO_59 (O_59,N_9996,N_9010);
nor UO_60 (O_60,N_9073,N_9662);
xor UO_61 (O_61,N_9354,N_9584);
nand UO_62 (O_62,N_9694,N_9121);
nor UO_63 (O_63,N_9449,N_9713);
or UO_64 (O_64,N_9705,N_9624);
nand UO_65 (O_65,N_9120,N_9142);
or UO_66 (O_66,N_9004,N_9196);
xor UO_67 (O_67,N_9083,N_9066);
nor UO_68 (O_68,N_9110,N_9677);
nor UO_69 (O_69,N_9069,N_9931);
nor UO_70 (O_70,N_9118,N_9716);
and UO_71 (O_71,N_9182,N_9504);
and UO_72 (O_72,N_9462,N_9819);
nand UO_73 (O_73,N_9787,N_9766);
or UO_74 (O_74,N_9642,N_9145);
or UO_75 (O_75,N_9952,N_9317);
xnor UO_76 (O_76,N_9484,N_9210);
xor UO_77 (O_77,N_9508,N_9477);
or UO_78 (O_78,N_9493,N_9501);
nand UO_79 (O_79,N_9208,N_9739);
or UO_80 (O_80,N_9548,N_9914);
nand UO_81 (O_81,N_9567,N_9552);
nand UO_82 (O_82,N_9815,N_9200);
and UO_83 (O_83,N_9919,N_9318);
nor UO_84 (O_84,N_9464,N_9304);
and UO_85 (O_85,N_9138,N_9214);
nand UO_86 (O_86,N_9641,N_9697);
nor UO_87 (O_87,N_9941,N_9755);
nor UO_88 (O_88,N_9897,N_9753);
and UO_89 (O_89,N_9060,N_9505);
nor UO_90 (O_90,N_9583,N_9890);
xor UO_91 (O_91,N_9235,N_9151);
xnor UO_92 (O_92,N_9144,N_9820);
xor UO_93 (O_93,N_9836,N_9316);
nor UO_94 (O_94,N_9539,N_9046);
nand UO_95 (O_95,N_9360,N_9306);
and UO_96 (O_96,N_9163,N_9445);
nand UO_97 (O_97,N_9562,N_9609);
nand UO_98 (O_98,N_9190,N_9472);
and UO_99 (O_99,N_9911,N_9043);
and UO_100 (O_100,N_9520,N_9018);
nand UO_101 (O_101,N_9847,N_9398);
or UO_102 (O_102,N_9324,N_9102);
nand UO_103 (O_103,N_9825,N_9627);
nand UO_104 (O_104,N_9419,N_9711);
and UO_105 (O_105,N_9668,N_9866);
or UO_106 (O_106,N_9412,N_9676);
nand UO_107 (O_107,N_9237,N_9219);
or UO_108 (O_108,N_9005,N_9986);
xnor UO_109 (O_109,N_9081,N_9287);
or UO_110 (O_110,N_9225,N_9198);
nand UO_111 (O_111,N_9093,N_9724);
or UO_112 (O_112,N_9114,N_9802);
nor UO_113 (O_113,N_9632,N_9420);
nand UO_114 (O_114,N_9152,N_9042);
xnor UO_115 (O_115,N_9158,N_9068);
nor UO_116 (O_116,N_9580,N_9966);
and UO_117 (O_117,N_9095,N_9809);
or UO_118 (O_118,N_9143,N_9748);
xor UO_119 (O_119,N_9803,N_9211);
and UO_120 (O_120,N_9045,N_9626);
xor UO_121 (O_121,N_9156,N_9698);
nand UO_122 (O_122,N_9232,N_9775);
nand UO_123 (O_123,N_9488,N_9348);
or UO_124 (O_124,N_9154,N_9774);
nor UO_125 (O_125,N_9185,N_9389);
or UO_126 (O_126,N_9760,N_9314);
or UO_127 (O_127,N_9796,N_9240);
nand UO_128 (O_128,N_9041,N_9157);
nand UO_129 (O_129,N_9329,N_9305);
xnor UO_130 (O_130,N_9763,N_9181);
and UO_131 (O_131,N_9710,N_9833);
or UO_132 (O_132,N_9194,N_9301);
and UO_133 (O_133,N_9893,N_9414);
nand UO_134 (O_134,N_9758,N_9957);
and UO_135 (O_135,N_9850,N_9249);
or UO_136 (O_136,N_9667,N_9685);
xnor UO_137 (O_137,N_9933,N_9492);
or UO_138 (O_138,N_9104,N_9653);
and UO_139 (O_139,N_9646,N_9738);
nor UO_140 (O_140,N_9468,N_9835);
and UO_141 (O_141,N_9561,N_9977);
nor UO_142 (O_142,N_9009,N_9117);
nor UO_143 (O_143,N_9457,N_9466);
or UO_144 (O_144,N_9257,N_9003);
or UO_145 (O_145,N_9437,N_9132);
xor UO_146 (O_146,N_9050,N_9669);
and UO_147 (O_147,N_9338,N_9298);
nor UO_148 (O_148,N_9469,N_9871);
and UO_149 (O_149,N_9213,N_9541);
xnor UO_150 (O_150,N_9598,N_9302);
and UO_151 (O_151,N_9939,N_9528);
and UO_152 (O_152,N_9342,N_9463);
nand UO_153 (O_153,N_9830,N_9907);
xnor UO_154 (O_154,N_9278,N_9652);
and UO_155 (O_155,N_9971,N_9859);
or UO_156 (O_156,N_9243,N_9707);
or UO_157 (O_157,N_9533,N_9250);
and UO_158 (O_158,N_9892,N_9319);
xor UO_159 (O_159,N_9681,N_9441);
and UO_160 (O_160,N_9682,N_9806);
or UO_161 (O_161,N_9875,N_9581);
nand UO_162 (O_162,N_9734,N_9428);
or UO_163 (O_163,N_9184,N_9277);
xor UO_164 (O_164,N_9894,N_9658);
and UO_165 (O_165,N_9885,N_9722);
xor UO_166 (O_166,N_9031,N_9726);
nand UO_167 (O_167,N_9822,N_9665);
xnor UO_168 (O_168,N_9368,N_9430);
xnor UO_169 (O_169,N_9364,N_9128);
nor UO_170 (O_170,N_9864,N_9034);
or UO_171 (O_171,N_9741,N_9309);
xnor UO_172 (O_172,N_9053,N_9221);
nand UO_173 (O_173,N_9877,N_9358);
nor UO_174 (O_174,N_9740,N_9097);
or UO_175 (O_175,N_9406,N_9267);
xor UO_176 (O_176,N_9995,N_9512);
xor UO_177 (O_177,N_9055,N_9197);
or UO_178 (O_178,N_9300,N_9982);
or UO_179 (O_179,N_9486,N_9880);
or UO_180 (O_180,N_9834,N_9715);
nand UO_181 (O_181,N_9779,N_9647);
or UO_182 (O_182,N_9888,N_9374);
xor UO_183 (O_183,N_9489,N_9498);
xor UO_184 (O_184,N_9103,N_9276);
and UO_185 (O_185,N_9279,N_9631);
xnor UO_186 (O_186,N_9186,N_9183);
or UO_187 (O_187,N_9659,N_9917);
or UO_188 (O_188,N_9096,N_9577);
xnor UO_189 (O_189,N_9199,N_9854);
and UO_190 (O_190,N_9044,N_9729);
nand UO_191 (O_191,N_9134,N_9180);
xnor UO_192 (O_192,N_9950,N_9867);
xor UO_193 (O_193,N_9856,N_9530);
xor UO_194 (O_194,N_9664,N_9930);
and UO_195 (O_195,N_9088,N_9790);
nand UO_196 (O_196,N_9882,N_9759);
nor UO_197 (O_197,N_9841,N_9953);
nand UO_198 (O_198,N_9233,N_9780);
nand UO_199 (O_199,N_9351,N_9418);
xor UO_200 (O_200,N_9554,N_9065);
nand UO_201 (O_201,N_9490,N_9357);
or UO_202 (O_202,N_9703,N_9299);
nor UO_203 (O_203,N_9997,N_9452);
or UO_204 (O_204,N_9136,N_9051);
nand UO_205 (O_205,N_9988,N_9507);
nor UO_206 (O_206,N_9310,N_9800);
nor UO_207 (O_207,N_9030,N_9303);
or UO_208 (O_208,N_9797,N_9785);
or UO_209 (O_209,N_9951,N_9960);
nor UO_210 (O_210,N_9858,N_9695);
nand UO_211 (O_211,N_9550,N_9435);
or UO_212 (O_212,N_9928,N_9161);
and UO_213 (O_213,N_9109,N_9896);
or UO_214 (O_214,N_9460,N_9344);
nand UO_215 (O_215,N_9876,N_9639);
or UO_216 (O_216,N_9191,N_9612);
and UO_217 (O_217,N_9693,N_9948);
nand UO_218 (O_218,N_9636,N_9993);
xor UO_219 (O_219,N_9560,N_9230);
and UO_220 (O_220,N_9105,N_9321);
nand UO_221 (O_221,N_9638,N_9475);
nor UO_222 (O_222,N_9661,N_9122);
and UO_223 (O_223,N_9777,N_9193);
and UO_224 (O_224,N_9404,N_9608);
nand UO_225 (O_225,N_9129,N_9973);
nor UO_226 (O_226,N_9421,N_9663);
and UO_227 (O_227,N_9401,N_9934);
or UO_228 (O_228,N_9119,N_9330);
or UO_229 (O_229,N_9910,N_9614);
or UO_230 (O_230,N_9206,N_9746);
xnor UO_231 (O_231,N_9818,N_9853);
and UO_232 (O_232,N_9023,N_9990);
nor UO_233 (O_233,N_9747,N_9112);
nor UO_234 (O_234,N_9355,N_9630);
nand UO_235 (O_235,N_9012,N_9970);
nor UO_236 (O_236,N_9666,N_9169);
or UO_237 (O_237,N_9162,N_9680);
and UO_238 (O_238,N_9699,N_9778);
xnor UO_239 (O_239,N_9730,N_9606);
nand UO_240 (O_240,N_9816,N_9688);
nor UO_241 (O_241,N_9657,N_9605);
nor UO_242 (O_242,N_9706,N_9599);
nand UO_243 (O_243,N_9634,N_9063);
nor UO_244 (O_244,N_9502,N_9307);
and UO_245 (O_245,N_9607,N_9969);
xor UO_246 (O_246,N_9650,N_9629);
nor UO_247 (O_247,N_9131,N_9263);
nor UO_248 (O_248,N_9901,N_9826);
and UO_249 (O_249,N_9280,N_9968);
nor UO_250 (O_250,N_9503,N_9378);
and UO_251 (O_251,N_9510,N_9337);
nor UO_252 (O_252,N_9524,N_9242);
or UO_253 (O_253,N_9436,N_9481);
or UO_254 (O_254,N_9167,N_9000);
nor UO_255 (O_255,N_9860,N_9821);
xnor UO_256 (O_256,N_9980,N_9992);
nor UO_257 (O_257,N_9228,N_9438);
nor UO_258 (O_258,N_9165,N_9518);
and UO_259 (O_259,N_9273,N_9149);
nor UO_260 (O_260,N_9424,N_9178);
nor UO_261 (O_261,N_9135,N_9732);
nor UO_262 (O_262,N_9383,N_9403);
and UO_263 (O_263,N_9842,N_9979);
and UO_264 (O_264,N_9013,N_9623);
nand UO_265 (O_265,N_9981,N_9616);
xor UO_266 (O_266,N_9071,N_9592);
nand UO_267 (O_267,N_9147,N_9656);
xor UO_268 (O_268,N_9223,N_9862);
nor UO_269 (O_269,N_9975,N_9878);
xor UO_270 (O_270,N_9347,N_9229);
nand UO_271 (O_271,N_9429,N_9870);
or UO_272 (O_272,N_9153,N_9067);
or UO_273 (O_273,N_9844,N_9772);
and UO_274 (O_274,N_9485,N_9513);
nand UO_275 (O_275,N_9813,N_9367);
and UO_276 (O_276,N_9720,N_9079);
or UO_277 (O_277,N_9923,N_9380);
nand UO_278 (O_278,N_9341,N_9805);
nand UO_279 (O_279,N_9852,N_9585);
nand UO_280 (O_280,N_9525,N_9189);
nor UO_281 (O_281,N_9220,N_9409);
nand UO_282 (O_282,N_9399,N_9113);
nor UO_283 (O_283,N_9308,N_9547);
or UO_284 (O_284,N_9215,N_9660);
nand UO_285 (O_285,N_9293,N_9056);
xor UO_286 (O_286,N_9028,N_9610);
nor UO_287 (O_287,N_9447,N_9076);
and UO_288 (O_288,N_9569,N_9094);
and UO_289 (O_289,N_9555,N_9648);
xnor UO_290 (O_290,N_9617,N_9670);
and UO_291 (O_291,N_9684,N_9495);
and UO_292 (O_292,N_9227,N_9687);
and UO_293 (O_293,N_9195,N_9288);
nor UO_294 (O_294,N_9515,N_9007);
nor UO_295 (O_295,N_9719,N_9212);
and UO_296 (O_296,N_9432,N_9072);
and UO_297 (O_297,N_9170,N_9395);
xor UO_298 (O_298,N_9423,N_9909);
or UO_299 (O_299,N_9171,N_9036);
nor UO_300 (O_300,N_9286,N_9543);
and UO_301 (O_301,N_9831,N_9804);
and UO_302 (O_302,N_9408,N_9070);
or UO_303 (O_303,N_9947,N_9540);
and UO_304 (O_304,N_9285,N_9001);
nor UO_305 (O_305,N_9356,N_9175);
and UO_306 (O_306,N_9461,N_9701);
nand UO_307 (O_307,N_9448,N_9439);
xor UO_308 (O_308,N_9579,N_9203);
and UO_309 (O_309,N_9937,N_9762);
or UO_310 (O_310,N_9619,N_9573);
nor UO_311 (O_311,N_9075,N_9396);
xor UO_312 (O_312,N_9899,N_9497);
or UO_313 (O_313,N_9062,N_9019);
xnor UO_314 (O_314,N_9218,N_9291);
or UO_315 (O_315,N_9839,N_9718);
nand UO_316 (O_316,N_9405,N_9352);
nor UO_317 (O_317,N_9478,N_9426);
and UO_318 (O_318,N_9792,N_9736);
or UO_319 (O_319,N_9544,N_9594);
xnor UO_320 (O_320,N_9021,N_9516);
and UO_321 (O_321,N_9700,N_9111);
nor UO_322 (O_322,N_9801,N_9604);
or UO_323 (O_323,N_9209,N_9381);
nand UO_324 (O_324,N_9905,N_9259);
and UO_325 (O_325,N_9234,N_9365);
nand UO_326 (O_326,N_9049,N_9538);
and UO_327 (O_327,N_9786,N_9768);
nand UO_328 (O_328,N_9906,N_9902);
nand UO_329 (O_329,N_9480,N_9578);
or UO_330 (O_330,N_9884,N_9271);
nor UO_331 (O_331,N_9689,N_9390);
or UO_332 (O_332,N_9921,N_9458);
nor UO_333 (O_333,N_9618,N_9294);
xor UO_334 (O_334,N_9678,N_9446);
and UO_335 (O_335,N_9529,N_9633);
xor UO_336 (O_336,N_9253,N_9959);
or UO_337 (O_337,N_9824,N_9838);
nor UO_338 (O_338,N_9984,N_9654);
or UO_339 (O_339,N_9177,N_9615);
nand UO_340 (O_340,N_9417,N_9089);
xor UO_341 (O_341,N_9350,N_9098);
or UO_342 (O_342,N_9874,N_9873);
or UO_343 (O_343,N_9949,N_9247);
or UO_344 (O_344,N_9014,N_9440);
nand UO_345 (O_345,N_9471,N_9467);
nand UO_346 (O_346,N_9602,N_9557);
xnor UO_347 (O_347,N_9099,N_9024);
xor UO_348 (O_348,N_9721,N_9817);
and UO_349 (O_349,N_9236,N_9749);
xor UO_350 (O_350,N_9108,N_9511);
or UO_351 (O_351,N_9895,N_9549);
nand UO_352 (O_352,N_9978,N_9848);
nand UO_353 (O_353,N_9613,N_9296);
and UO_354 (O_354,N_9246,N_9994);
nand UO_355 (O_355,N_9974,N_9187);
nor UO_356 (O_356,N_9384,N_9708);
or UO_357 (O_357,N_9837,N_9313);
and UO_358 (O_358,N_9137,N_9723);
nor UO_359 (O_359,N_9620,N_9509);
nor UO_360 (O_360,N_9537,N_9349);
or UO_361 (O_361,N_9125,N_9571);
and UO_362 (O_362,N_9465,N_9843);
and UO_363 (O_363,N_9496,N_9940);
xor UO_364 (O_364,N_9370,N_9361);
or UO_365 (O_365,N_9394,N_9216);
xor UO_366 (O_366,N_9926,N_9252);
xnor UO_367 (O_367,N_9869,N_9047);
nand UO_368 (O_368,N_9331,N_9855);
and UO_369 (O_369,N_9991,N_9916);
and UO_370 (O_370,N_9020,N_9958);
nand UO_371 (O_371,N_9770,N_9393);
xnor UO_372 (O_372,N_9590,N_9891);
nand UO_373 (O_373,N_9733,N_9265);
or UO_374 (O_374,N_9572,N_9611);
nand UO_375 (O_375,N_9202,N_9872);
nand UO_376 (O_376,N_9743,N_9454);
nand UO_377 (O_377,N_9139,N_9260);
xnor UO_378 (O_378,N_9556,N_9640);
and UO_379 (O_379,N_9133,N_9025);
or UO_380 (O_380,N_9415,N_9256);
xor UO_381 (O_381,N_9591,N_9422);
nor UO_382 (O_382,N_9266,N_9832);
nand UO_383 (O_383,N_9379,N_9735);
nor UO_384 (O_384,N_9692,N_9932);
and UO_385 (O_385,N_9771,N_9150);
nor UO_386 (O_386,N_9886,N_9311);
or UO_387 (O_387,N_9696,N_9945);
xor UO_388 (O_388,N_9807,N_9127);
nor UO_389 (O_389,N_9651,N_9366);
nor UO_390 (O_390,N_9107,N_9521);
nor UO_391 (O_391,N_9863,N_9140);
xnor UO_392 (O_392,N_9373,N_9328);
xor UO_393 (O_393,N_9146,N_9048);
or UO_394 (O_394,N_9675,N_9954);
xnor UO_395 (O_395,N_9535,N_9588);
and UO_396 (O_396,N_9861,N_9725);
and UO_397 (O_397,N_9343,N_9534);
or UO_398 (O_398,N_9898,N_9474);
or UO_399 (O_399,N_9333,N_9765);
nor UO_400 (O_400,N_9148,N_9754);
xor UO_401 (O_401,N_9101,N_9918);
nor UO_402 (O_402,N_9912,N_9929);
nand UO_403 (O_403,N_9717,N_9788);
nand UO_404 (O_404,N_9057,N_9444);
nand UO_405 (O_405,N_9589,N_9346);
and UO_406 (O_406,N_9168,N_9085);
xor UO_407 (O_407,N_9433,N_9116);
or UO_408 (O_408,N_9702,N_9621);
nand UO_409 (O_409,N_9386,N_9315);
nand UO_410 (O_410,N_9479,N_9983);
or UO_411 (O_411,N_9106,N_9622);
or UO_412 (O_412,N_9673,N_9231);
nor UO_413 (O_413,N_9679,N_9179);
nor UO_414 (O_414,N_9087,N_9714);
or UO_415 (O_415,N_9987,N_9058);
or UO_416 (O_416,N_9823,N_9967);
nor UO_417 (O_417,N_9938,N_9728);
nand UO_418 (O_418,N_9082,N_9494);
nor UO_419 (O_419,N_9090,N_9744);
nand UO_420 (O_420,N_9925,N_9382);
xnor UO_421 (O_421,N_9155,N_9814);
and UO_422 (O_422,N_9965,N_9188);
nand UO_423 (O_423,N_9546,N_9022);
nand UO_424 (O_424,N_9791,N_9470);
or UO_425 (O_425,N_9936,N_9410);
and UO_426 (O_426,N_9371,N_9274);
and UO_427 (O_427,N_9935,N_9595);
and UO_428 (O_428,N_9799,N_9015);
nand UO_429 (O_429,N_9086,N_9846);
nand UO_430 (O_430,N_9054,N_9264);
nand UO_431 (O_431,N_9811,N_9883);
or UO_432 (O_432,N_9176,N_9751);
nor UO_433 (O_433,N_9808,N_9284);
xor UO_434 (O_434,N_9459,N_9961);
nor UO_435 (O_435,N_9431,N_9413);
nand UO_436 (O_436,N_9542,N_9962);
and UO_437 (O_437,N_9955,N_9944);
or UO_438 (O_438,N_9434,N_9575);
xor UO_439 (O_439,N_9323,N_9130);
and UO_440 (O_440,N_9159,N_9674);
nor UO_441 (O_441,N_9325,N_9483);
nor UO_442 (O_442,N_9908,N_9442);
nor UO_443 (O_443,N_9141,N_9686);
nor UO_444 (O_444,N_9100,N_9964);
nor UO_445 (O_445,N_9340,N_9644);
nand UO_446 (O_446,N_9563,N_9603);
nand UO_447 (O_447,N_9709,N_9241);
nor UO_448 (O_448,N_9587,N_9353);
xor UO_449 (O_449,N_9416,N_9029);
or UO_450 (O_450,N_9500,N_9566);
or UO_451 (O_451,N_9551,N_9040);
nor UO_452 (O_452,N_9261,N_9985);
and UO_453 (O_453,N_9268,N_9397);
and UO_454 (O_454,N_9655,N_9039);
nor UO_455 (O_455,N_9691,N_9531);
nor UO_456 (O_456,N_9499,N_9244);
and UO_457 (O_457,N_9077,N_9033);
or UO_458 (O_458,N_9999,N_9812);
nor UO_459 (O_459,N_9335,N_9559);
xnor UO_460 (O_460,N_9297,N_9425);
or UO_461 (O_461,N_9756,N_9270);
nor UO_462 (O_462,N_9840,N_9731);
nand UO_463 (O_463,N_9868,N_9205);
xnor UO_464 (O_464,N_9035,N_9456);
nand UO_465 (O_465,N_9164,N_9172);
or UO_466 (O_466,N_9963,N_9402);
and UO_467 (O_467,N_9943,N_9506);
and UO_468 (O_468,N_9372,N_9789);
xnor UO_469 (O_469,N_9369,N_9810);
nor UO_470 (O_470,N_9224,N_9388);
nand UO_471 (O_471,N_9363,N_9553);
or UO_472 (O_472,N_9798,N_9752);
nand UO_473 (O_473,N_9946,N_9887);
nor UO_474 (O_474,N_9115,N_9027);
nor UO_475 (O_475,N_9881,N_9359);
nor UO_476 (O_476,N_9295,N_9326);
nand UO_477 (O_477,N_9794,N_9160);
xnor UO_478 (O_478,N_9245,N_9052);
nor UO_479 (O_479,N_9269,N_9913);
nor UO_480 (O_480,N_9845,N_9084);
nor UO_481 (O_481,N_9173,N_9078);
or UO_482 (O_482,N_9776,N_9712);
nand UO_483 (O_483,N_9254,N_9879);
and UO_484 (O_484,N_9275,N_9764);
nor UO_485 (O_485,N_9889,N_9976);
or UO_486 (O_486,N_9217,N_9385);
nor UO_487 (O_487,N_9207,N_9827);
nand UO_488 (O_488,N_9915,N_9829);
nand UO_489 (O_489,N_9564,N_9006);
xor UO_490 (O_490,N_9011,N_9527);
and UO_491 (O_491,N_9761,N_9283);
nand UO_492 (O_492,N_9920,N_9769);
nand UO_493 (O_493,N_9038,N_9272);
and UO_494 (O_494,N_9582,N_9773);
nor UO_495 (O_495,N_9282,N_9061);
nand UO_496 (O_496,N_9123,N_9248);
nor UO_497 (O_497,N_9336,N_9927);
nor UO_498 (O_498,N_9080,N_9989);
xor UO_499 (O_499,N_9362,N_9857);
and UO_500 (O_500,N_9340,N_9780);
or UO_501 (O_501,N_9128,N_9757);
and UO_502 (O_502,N_9029,N_9139);
or UO_503 (O_503,N_9210,N_9385);
or UO_504 (O_504,N_9195,N_9046);
nor UO_505 (O_505,N_9876,N_9046);
xor UO_506 (O_506,N_9601,N_9604);
and UO_507 (O_507,N_9600,N_9769);
or UO_508 (O_508,N_9651,N_9118);
and UO_509 (O_509,N_9028,N_9039);
nand UO_510 (O_510,N_9841,N_9827);
and UO_511 (O_511,N_9151,N_9566);
nor UO_512 (O_512,N_9448,N_9106);
or UO_513 (O_513,N_9432,N_9457);
and UO_514 (O_514,N_9761,N_9745);
nor UO_515 (O_515,N_9206,N_9601);
nor UO_516 (O_516,N_9774,N_9027);
xnor UO_517 (O_517,N_9438,N_9097);
nand UO_518 (O_518,N_9237,N_9591);
and UO_519 (O_519,N_9644,N_9145);
xnor UO_520 (O_520,N_9069,N_9990);
nor UO_521 (O_521,N_9381,N_9990);
xnor UO_522 (O_522,N_9679,N_9180);
or UO_523 (O_523,N_9747,N_9298);
or UO_524 (O_524,N_9711,N_9602);
nor UO_525 (O_525,N_9384,N_9875);
or UO_526 (O_526,N_9849,N_9436);
xor UO_527 (O_527,N_9486,N_9950);
or UO_528 (O_528,N_9318,N_9352);
nand UO_529 (O_529,N_9734,N_9589);
and UO_530 (O_530,N_9356,N_9703);
or UO_531 (O_531,N_9815,N_9121);
nand UO_532 (O_532,N_9476,N_9739);
nand UO_533 (O_533,N_9939,N_9112);
and UO_534 (O_534,N_9990,N_9665);
and UO_535 (O_535,N_9850,N_9118);
nor UO_536 (O_536,N_9284,N_9163);
and UO_537 (O_537,N_9638,N_9584);
nand UO_538 (O_538,N_9580,N_9013);
or UO_539 (O_539,N_9792,N_9209);
xor UO_540 (O_540,N_9523,N_9231);
xor UO_541 (O_541,N_9752,N_9593);
xor UO_542 (O_542,N_9548,N_9748);
nand UO_543 (O_543,N_9517,N_9704);
nand UO_544 (O_544,N_9868,N_9112);
and UO_545 (O_545,N_9080,N_9277);
or UO_546 (O_546,N_9544,N_9179);
or UO_547 (O_547,N_9464,N_9744);
xnor UO_548 (O_548,N_9915,N_9932);
or UO_549 (O_549,N_9422,N_9489);
and UO_550 (O_550,N_9426,N_9211);
nor UO_551 (O_551,N_9506,N_9322);
xnor UO_552 (O_552,N_9005,N_9805);
nor UO_553 (O_553,N_9989,N_9742);
nor UO_554 (O_554,N_9970,N_9596);
or UO_555 (O_555,N_9085,N_9121);
and UO_556 (O_556,N_9051,N_9249);
nand UO_557 (O_557,N_9927,N_9663);
xnor UO_558 (O_558,N_9653,N_9141);
xor UO_559 (O_559,N_9390,N_9801);
and UO_560 (O_560,N_9662,N_9864);
or UO_561 (O_561,N_9281,N_9566);
or UO_562 (O_562,N_9216,N_9260);
xor UO_563 (O_563,N_9742,N_9200);
nor UO_564 (O_564,N_9238,N_9331);
nand UO_565 (O_565,N_9980,N_9478);
nor UO_566 (O_566,N_9801,N_9444);
xnor UO_567 (O_567,N_9053,N_9532);
or UO_568 (O_568,N_9321,N_9600);
and UO_569 (O_569,N_9982,N_9588);
or UO_570 (O_570,N_9580,N_9829);
and UO_571 (O_571,N_9872,N_9582);
xnor UO_572 (O_572,N_9867,N_9235);
nor UO_573 (O_573,N_9172,N_9505);
nand UO_574 (O_574,N_9760,N_9089);
nand UO_575 (O_575,N_9625,N_9127);
or UO_576 (O_576,N_9617,N_9373);
nand UO_577 (O_577,N_9181,N_9977);
xor UO_578 (O_578,N_9588,N_9138);
nand UO_579 (O_579,N_9009,N_9832);
or UO_580 (O_580,N_9935,N_9496);
nor UO_581 (O_581,N_9803,N_9448);
nand UO_582 (O_582,N_9476,N_9630);
nor UO_583 (O_583,N_9099,N_9506);
xor UO_584 (O_584,N_9968,N_9527);
xnor UO_585 (O_585,N_9299,N_9141);
xnor UO_586 (O_586,N_9364,N_9922);
or UO_587 (O_587,N_9780,N_9180);
nand UO_588 (O_588,N_9138,N_9610);
and UO_589 (O_589,N_9283,N_9727);
xor UO_590 (O_590,N_9693,N_9408);
and UO_591 (O_591,N_9835,N_9990);
and UO_592 (O_592,N_9909,N_9897);
nand UO_593 (O_593,N_9012,N_9893);
nor UO_594 (O_594,N_9085,N_9374);
xor UO_595 (O_595,N_9460,N_9090);
nand UO_596 (O_596,N_9566,N_9129);
and UO_597 (O_597,N_9709,N_9217);
or UO_598 (O_598,N_9797,N_9060);
xnor UO_599 (O_599,N_9882,N_9240);
or UO_600 (O_600,N_9308,N_9514);
nor UO_601 (O_601,N_9717,N_9976);
nand UO_602 (O_602,N_9016,N_9791);
nor UO_603 (O_603,N_9436,N_9284);
and UO_604 (O_604,N_9944,N_9512);
xor UO_605 (O_605,N_9817,N_9751);
or UO_606 (O_606,N_9881,N_9961);
nor UO_607 (O_607,N_9959,N_9209);
or UO_608 (O_608,N_9936,N_9086);
xnor UO_609 (O_609,N_9057,N_9898);
nand UO_610 (O_610,N_9431,N_9034);
and UO_611 (O_611,N_9959,N_9133);
xor UO_612 (O_612,N_9580,N_9803);
nand UO_613 (O_613,N_9686,N_9852);
xnor UO_614 (O_614,N_9890,N_9922);
nor UO_615 (O_615,N_9610,N_9089);
nor UO_616 (O_616,N_9884,N_9660);
or UO_617 (O_617,N_9458,N_9706);
xor UO_618 (O_618,N_9927,N_9506);
nand UO_619 (O_619,N_9224,N_9302);
nand UO_620 (O_620,N_9876,N_9075);
xnor UO_621 (O_621,N_9151,N_9359);
xor UO_622 (O_622,N_9214,N_9096);
nand UO_623 (O_623,N_9122,N_9458);
nor UO_624 (O_624,N_9310,N_9366);
and UO_625 (O_625,N_9663,N_9039);
xnor UO_626 (O_626,N_9041,N_9301);
xnor UO_627 (O_627,N_9230,N_9227);
nand UO_628 (O_628,N_9130,N_9850);
or UO_629 (O_629,N_9324,N_9545);
and UO_630 (O_630,N_9852,N_9501);
and UO_631 (O_631,N_9276,N_9734);
nor UO_632 (O_632,N_9444,N_9615);
nor UO_633 (O_633,N_9541,N_9905);
xor UO_634 (O_634,N_9495,N_9992);
or UO_635 (O_635,N_9958,N_9933);
and UO_636 (O_636,N_9850,N_9729);
nor UO_637 (O_637,N_9418,N_9042);
and UO_638 (O_638,N_9441,N_9596);
nand UO_639 (O_639,N_9748,N_9154);
xnor UO_640 (O_640,N_9172,N_9175);
or UO_641 (O_641,N_9221,N_9540);
and UO_642 (O_642,N_9886,N_9098);
or UO_643 (O_643,N_9264,N_9376);
or UO_644 (O_644,N_9051,N_9033);
nand UO_645 (O_645,N_9049,N_9414);
nor UO_646 (O_646,N_9078,N_9534);
xor UO_647 (O_647,N_9402,N_9834);
or UO_648 (O_648,N_9991,N_9287);
nor UO_649 (O_649,N_9623,N_9565);
or UO_650 (O_650,N_9463,N_9914);
and UO_651 (O_651,N_9616,N_9457);
and UO_652 (O_652,N_9165,N_9700);
or UO_653 (O_653,N_9029,N_9190);
nand UO_654 (O_654,N_9134,N_9611);
nand UO_655 (O_655,N_9205,N_9371);
and UO_656 (O_656,N_9798,N_9853);
nand UO_657 (O_657,N_9553,N_9158);
and UO_658 (O_658,N_9764,N_9505);
nand UO_659 (O_659,N_9821,N_9153);
xnor UO_660 (O_660,N_9156,N_9254);
xnor UO_661 (O_661,N_9279,N_9424);
nand UO_662 (O_662,N_9128,N_9996);
nor UO_663 (O_663,N_9063,N_9018);
and UO_664 (O_664,N_9413,N_9569);
nand UO_665 (O_665,N_9486,N_9008);
nor UO_666 (O_666,N_9433,N_9184);
and UO_667 (O_667,N_9912,N_9868);
or UO_668 (O_668,N_9320,N_9592);
and UO_669 (O_669,N_9622,N_9020);
or UO_670 (O_670,N_9006,N_9513);
nand UO_671 (O_671,N_9666,N_9977);
and UO_672 (O_672,N_9633,N_9113);
nand UO_673 (O_673,N_9807,N_9998);
nand UO_674 (O_674,N_9593,N_9676);
nand UO_675 (O_675,N_9676,N_9792);
and UO_676 (O_676,N_9863,N_9954);
nand UO_677 (O_677,N_9727,N_9900);
nand UO_678 (O_678,N_9761,N_9757);
nand UO_679 (O_679,N_9157,N_9885);
or UO_680 (O_680,N_9774,N_9282);
nand UO_681 (O_681,N_9722,N_9076);
nor UO_682 (O_682,N_9436,N_9530);
nand UO_683 (O_683,N_9567,N_9720);
nand UO_684 (O_684,N_9412,N_9214);
nand UO_685 (O_685,N_9031,N_9960);
nand UO_686 (O_686,N_9317,N_9744);
nand UO_687 (O_687,N_9171,N_9448);
nor UO_688 (O_688,N_9843,N_9273);
and UO_689 (O_689,N_9087,N_9879);
xor UO_690 (O_690,N_9471,N_9728);
nor UO_691 (O_691,N_9978,N_9322);
and UO_692 (O_692,N_9043,N_9943);
nor UO_693 (O_693,N_9749,N_9476);
xor UO_694 (O_694,N_9210,N_9268);
nand UO_695 (O_695,N_9322,N_9156);
and UO_696 (O_696,N_9973,N_9603);
nor UO_697 (O_697,N_9881,N_9733);
nand UO_698 (O_698,N_9145,N_9598);
xnor UO_699 (O_699,N_9659,N_9213);
and UO_700 (O_700,N_9198,N_9539);
xor UO_701 (O_701,N_9647,N_9958);
or UO_702 (O_702,N_9524,N_9360);
and UO_703 (O_703,N_9805,N_9831);
and UO_704 (O_704,N_9766,N_9229);
xor UO_705 (O_705,N_9507,N_9697);
nand UO_706 (O_706,N_9189,N_9698);
nand UO_707 (O_707,N_9035,N_9866);
or UO_708 (O_708,N_9589,N_9819);
or UO_709 (O_709,N_9241,N_9811);
xor UO_710 (O_710,N_9277,N_9294);
nor UO_711 (O_711,N_9601,N_9098);
nand UO_712 (O_712,N_9615,N_9619);
nor UO_713 (O_713,N_9484,N_9352);
and UO_714 (O_714,N_9155,N_9648);
nor UO_715 (O_715,N_9055,N_9669);
and UO_716 (O_716,N_9249,N_9055);
or UO_717 (O_717,N_9462,N_9595);
or UO_718 (O_718,N_9222,N_9198);
nor UO_719 (O_719,N_9774,N_9974);
xor UO_720 (O_720,N_9431,N_9077);
or UO_721 (O_721,N_9336,N_9782);
xor UO_722 (O_722,N_9393,N_9752);
nor UO_723 (O_723,N_9375,N_9069);
xor UO_724 (O_724,N_9511,N_9936);
or UO_725 (O_725,N_9694,N_9523);
nand UO_726 (O_726,N_9368,N_9353);
nand UO_727 (O_727,N_9927,N_9051);
nor UO_728 (O_728,N_9136,N_9439);
or UO_729 (O_729,N_9156,N_9026);
nand UO_730 (O_730,N_9335,N_9076);
or UO_731 (O_731,N_9565,N_9555);
nand UO_732 (O_732,N_9192,N_9429);
nand UO_733 (O_733,N_9190,N_9903);
nand UO_734 (O_734,N_9067,N_9054);
nand UO_735 (O_735,N_9382,N_9468);
and UO_736 (O_736,N_9801,N_9065);
or UO_737 (O_737,N_9660,N_9926);
xor UO_738 (O_738,N_9041,N_9079);
nand UO_739 (O_739,N_9683,N_9244);
xnor UO_740 (O_740,N_9120,N_9792);
or UO_741 (O_741,N_9087,N_9338);
and UO_742 (O_742,N_9088,N_9076);
nor UO_743 (O_743,N_9197,N_9689);
xnor UO_744 (O_744,N_9391,N_9672);
or UO_745 (O_745,N_9114,N_9783);
xnor UO_746 (O_746,N_9598,N_9097);
nor UO_747 (O_747,N_9964,N_9661);
nor UO_748 (O_748,N_9444,N_9350);
or UO_749 (O_749,N_9675,N_9219);
nor UO_750 (O_750,N_9593,N_9479);
and UO_751 (O_751,N_9517,N_9469);
nand UO_752 (O_752,N_9629,N_9194);
nand UO_753 (O_753,N_9810,N_9793);
nand UO_754 (O_754,N_9689,N_9186);
and UO_755 (O_755,N_9556,N_9485);
xnor UO_756 (O_756,N_9441,N_9924);
nor UO_757 (O_757,N_9336,N_9966);
or UO_758 (O_758,N_9962,N_9350);
nor UO_759 (O_759,N_9899,N_9127);
and UO_760 (O_760,N_9785,N_9205);
xor UO_761 (O_761,N_9161,N_9373);
xnor UO_762 (O_762,N_9254,N_9073);
or UO_763 (O_763,N_9587,N_9947);
and UO_764 (O_764,N_9185,N_9842);
or UO_765 (O_765,N_9168,N_9208);
xnor UO_766 (O_766,N_9474,N_9829);
or UO_767 (O_767,N_9806,N_9095);
and UO_768 (O_768,N_9862,N_9034);
xnor UO_769 (O_769,N_9311,N_9468);
xor UO_770 (O_770,N_9505,N_9773);
nor UO_771 (O_771,N_9166,N_9713);
xnor UO_772 (O_772,N_9052,N_9552);
or UO_773 (O_773,N_9755,N_9695);
xor UO_774 (O_774,N_9773,N_9118);
or UO_775 (O_775,N_9088,N_9593);
xnor UO_776 (O_776,N_9492,N_9338);
nand UO_777 (O_777,N_9705,N_9714);
nand UO_778 (O_778,N_9861,N_9146);
nand UO_779 (O_779,N_9200,N_9563);
nand UO_780 (O_780,N_9890,N_9485);
nand UO_781 (O_781,N_9023,N_9858);
nand UO_782 (O_782,N_9887,N_9209);
or UO_783 (O_783,N_9630,N_9582);
or UO_784 (O_784,N_9212,N_9024);
nand UO_785 (O_785,N_9573,N_9673);
and UO_786 (O_786,N_9379,N_9648);
or UO_787 (O_787,N_9191,N_9412);
nor UO_788 (O_788,N_9671,N_9678);
nor UO_789 (O_789,N_9858,N_9426);
or UO_790 (O_790,N_9259,N_9135);
or UO_791 (O_791,N_9486,N_9673);
nor UO_792 (O_792,N_9853,N_9406);
nor UO_793 (O_793,N_9599,N_9236);
and UO_794 (O_794,N_9381,N_9776);
xor UO_795 (O_795,N_9518,N_9977);
xnor UO_796 (O_796,N_9213,N_9914);
nand UO_797 (O_797,N_9708,N_9363);
and UO_798 (O_798,N_9969,N_9079);
nor UO_799 (O_799,N_9411,N_9878);
and UO_800 (O_800,N_9807,N_9851);
or UO_801 (O_801,N_9160,N_9452);
nand UO_802 (O_802,N_9086,N_9177);
or UO_803 (O_803,N_9903,N_9944);
nor UO_804 (O_804,N_9170,N_9733);
and UO_805 (O_805,N_9163,N_9882);
and UO_806 (O_806,N_9679,N_9378);
xnor UO_807 (O_807,N_9031,N_9054);
nand UO_808 (O_808,N_9600,N_9443);
and UO_809 (O_809,N_9281,N_9379);
nor UO_810 (O_810,N_9845,N_9691);
and UO_811 (O_811,N_9718,N_9843);
and UO_812 (O_812,N_9492,N_9706);
or UO_813 (O_813,N_9777,N_9752);
or UO_814 (O_814,N_9030,N_9967);
or UO_815 (O_815,N_9552,N_9005);
xor UO_816 (O_816,N_9556,N_9346);
nand UO_817 (O_817,N_9683,N_9051);
xor UO_818 (O_818,N_9897,N_9047);
nor UO_819 (O_819,N_9694,N_9616);
or UO_820 (O_820,N_9926,N_9883);
xnor UO_821 (O_821,N_9347,N_9335);
or UO_822 (O_822,N_9785,N_9966);
or UO_823 (O_823,N_9252,N_9109);
nand UO_824 (O_824,N_9728,N_9137);
xor UO_825 (O_825,N_9691,N_9547);
and UO_826 (O_826,N_9470,N_9672);
nand UO_827 (O_827,N_9504,N_9198);
or UO_828 (O_828,N_9636,N_9807);
xnor UO_829 (O_829,N_9387,N_9282);
xor UO_830 (O_830,N_9899,N_9353);
xnor UO_831 (O_831,N_9057,N_9899);
or UO_832 (O_832,N_9767,N_9740);
or UO_833 (O_833,N_9708,N_9797);
nand UO_834 (O_834,N_9206,N_9834);
or UO_835 (O_835,N_9220,N_9982);
or UO_836 (O_836,N_9922,N_9277);
and UO_837 (O_837,N_9548,N_9701);
and UO_838 (O_838,N_9165,N_9423);
and UO_839 (O_839,N_9079,N_9855);
nor UO_840 (O_840,N_9041,N_9768);
nand UO_841 (O_841,N_9873,N_9640);
xnor UO_842 (O_842,N_9631,N_9219);
xor UO_843 (O_843,N_9945,N_9657);
and UO_844 (O_844,N_9337,N_9939);
or UO_845 (O_845,N_9646,N_9035);
or UO_846 (O_846,N_9930,N_9767);
nand UO_847 (O_847,N_9613,N_9065);
and UO_848 (O_848,N_9799,N_9819);
and UO_849 (O_849,N_9291,N_9464);
and UO_850 (O_850,N_9863,N_9476);
xnor UO_851 (O_851,N_9768,N_9181);
or UO_852 (O_852,N_9583,N_9280);
or UO_853 (O_853,N_9426,N_9156);
or UO_854 (O_854,N_9963,N_9338);
xnor UO_855 (O_855,N_9340,N_9833);
nor UO_856 (O_856,N_9854,N_9137);
xnor UO_857 (O_857,N_9543,N_9880);
or UO_858 (O_858,N_9411,N_9150);
nand UO_859 (O_859,N_9945,N_9403);
xnor UO_860 (O_860,N_9534,N_9034);
nor UO_861 (O_861,N_9076,N_9217);
nor UO_862 (O_862,N_9117,N_9392);
xor UO_863 (O_863,N_9959,N_9464);
nor UO_864 (O_864,N_9611,N_9281);
and UO_865 (O_865,N_9410,N_9122);
or UO_866 (O_866,N_9710,N_9367);
and UO_867 (O_867,N_9896,N_9336);
and UO_868 (O_868,N_9235,N_9806);
nand UO_869 (O_869,N_9203,N_9650);
nand UO_870 (O_870,N_9963,N_9955);
nor UO_871 (O_871,N_9311,N_9072);
or UO_872 (O_872,N_9035,N_9539);
xnor UO_873 (O_873,N_9474,N_9890);
xnor UO_874 (O_874,N_9402,N_9340);
and UO_875 (O_875,N_9740,N_9159);
xnor UO_876 (O_876,N_9845,N_9620);
or UO_877 (O_877,N_9264,N_9680);
nand UO_878 (O_878,N_9475,N_9957);
nor UO_879 (O_879,N_9044,N_9961);
xor UO_880 (O_880,N_9430,N_9646);
or UO_881 (O_881,N_9362,N_9359);
xor UO_882 (O_882,N_9574,N_9333);
nor UO_883 (O_883,N_9945,N_9396);
or UO_884 (O_884,N_9639,N_9427);
xor UO_885 (O_885,N_9006,N_9164);
or UO_886 (O_886,N_9491,N_9065);
nor UO_887 (O_887,N_9737,N_9067);
nor UO_888 (O_888,N_9327,N_9916);
xor UO_889 (O_889,N_9225,N_9226);
or UO_890 (O_890,N_9767,N_9617);
xnor UO_891 (O_891,N_9020,N_9013);
nor UO_892 (O_892,N_9617,N_9691);
and UO_893 (O_893,N_9398,N_9184);
or UO_894 (O_894,N_9018,N_9830);
nor UO_895 (O_895,N_9393,N_9997);
xnor UO_896 (O_896,N_9814,N_9713);
xnor UO_897 (O_897,N_9041,N_9987);
nor UO_898 (O_898,N_9479,N_9342);
nand UO_899 (O_899,N_9915,N_9836);
and UO_900 (O_900,N_9620,N_9722);
nor UO_901 (O_901,N_9419,N_9126);
or UO_902 (O_902,N_9137,N_9398);
or UO_903 (O_903,N_9888,N_9088);
nand UO_904 (O_904,N_9729,N_9912);
nor UO_905 (O_905,N_9294,N_9743);
nor UO_906 (O_906,N_9616,N_9439);
nor UO_907 (O_907,N_9734,N_9029);
nand UO_908 (O_908,N_9444,N_9782);
or UO_909 (O_909,N_9597,N_9440);
xnor UO_910 (O_910,N_9920,N_9729);
xor UO_911 (O_911,N_9880,N_9990);
nor UO_912 (O_912,N_9396,N_9514);
and UO_913 (O_913,N_9929,N_9256);
xor UO_914 (O_914,N_9025,N_9639);
nor UO_915 (O_915,N_9625,N_9865);
or UO_916 (O_916,N_9913,N_9633);
or UO_917 (O_917,N_9138,N_9115);
nand UO_918 (O_918,N_9636,N_9683);
and UO_919 (O_919,N_9286,N_9235);
xor UO_920 (O_920,N_9132,N_9888);
nor UO_921 (O_921,N_9048,N_9960);
nor UO_922 (O_922,N_9614,N_9093);
and UO_923 (O_923,N_9361,N_9475);
nand UO_924 (O_924,N_9031,N_9027);
or UO_925 (O_925,N_9195,N_9540);
or UO_926 (O_926,N_9885,N_9276);
nand UO_927 (O_927,N_9528,N_9255);
and UO_928 (O_928,N_9639,N_9183);
nand UO_929 (O_929,N_9211,N_9500);
nand UO_930 (O_930,N_9510,N_9452);
nor UO_931 (O_931,N_9921,N_9314);
xor UO_932 (O_932,N_9208,N_9145);
xnor UO_933 (O_933,N_9288,N_9950);
and UO_934 (O_934,N_9438,N_9616);
nand UO_935 (O_935,N_9865,N_9366);
or UO_936 (O_936,N_9504,N_9903);
and UO_937 (O_937,N_9035,N_9132);
or UO_938 (O_938,N_9347,N_9687);
and UO_939 (O_939,N_9382,N_9767);
or UO_940 (O_940,N_9186,N_9021);
or UO_941 (O_941,N_9358,N_9464);
nor UO_942 (O_942,N_9544,N_9777);
and UO_943 (O_943,N_9943,N_9497);
xnor UO_944 (O_944,N_9110,N_9163);
or UO_945 (O_945,N_9302,N_9475);
xor UO_946 (O_946,N_9140,N_9043);
nand UO_947 (O_947,N_9535,N_9780);
nand UO_948 (O_948,N_9908,N_9037);
nand UO_949 (O_949,N_9234,N_9547);
or UO_950 (O_950,N_9152,N_9982);
xnor UO_951 (O_951,N_9361,N_9044);
xor UO_952 (O_952,N_9888,N_9799);
xor UO_953 (O_953,N_9929,N_9735);
xnor UO_954 (O_954,N_9262,N_9707);
xnor UO_955 (O_955,N_9734,N_9969);
xnor UO_956 (O_956,N_9699,N_9653);
and UO_957 (O_957,N_9334,N_9610);
nor UO_958 (O_958,N_9837,N_9598);
or UO_959 (O_959,N_9353,N_9910);
xor UO_960 (O_960,N_9695,N_9111);
xor UO_961 (O_961,N_9212,N_9299);
and UO_962 (O_962,N_9047,N_9344);
xnor UO_963 (O_963,N_9066,N_9804);
and UO_964 (O_964,N_9350,N_9944);
or UO_965 (O_965,N_9086,N_9490);
or UO_966 (O_966,N_9441,N_9339);
nand UO_967 (O_967,N_9573,N_9889);
or UO_968 (O_968,N_9522,N_9959);
xnor UO_969 (O_969,N_9160,N_9559);
or UO_970 (O_970,N_9733,N_9293);
xor UO_971 (O_971,N_9129,N_9331);
nor UO_972 (O_972,N_9378,N_9759);
nand UO_973 (O_973,N_9138,N_9845);
nand UO_974 (O_974,N_9462,N_9418);
nor UO_975 (O_975,N_9980,N_9959);
and UO_976 (O_976,N_9833,N_9405);
nor UO_977 (O_977,N_9757,N_9453);
xor UO_978 (O_978,N_9444,N_9843);
xor UO_979 (O_979,N_9917,N_9315);
or UO_980 (O_980,N_9267,N_9338);
and UO_981 (O_981,N_9727,N_9992);
xnor UO_982 (O_982,N_9449,N_9424);
xor UO_983 (O_983,N_9764,N_9917);
nand UO_984 (O_984,N_9381,N_9485);
or UO_985 (O_985,N_9594,N_9549);
nand UO_986 (O_986,N_9667,N_9201);
or UO_987 (O_987,N_9286,N_9509);
nor UO_988 (O_988,N_9091,N_9928);
or UO_989 (O_989,N_9603,N_9184);
nor UO_990 (O_990,N_9059,N_9691);
nand UO_991 (O_991,N_9392,N_9695);
and UO_992 (O_992,N_9511,N_9410);
or UO_993 (O_993,N_9656,N_9954);
and UO_994 (O_994,N_9525,N_9533);
and UO_995 (O_995,N_9106,N_9262);
nand UO_996 (O_996,N_9348,N_9800);
nand UO_997 (O_997,N_9999,N_9324);
nand UO_998 (O_998,N_9184,N_9807);
xnor UO_999 (O_999,N_9520,N_9054);
nor UO_1000 (O_1000,N_9387,N_9272);
nor UO_1001 (O_1001,N_9557,N_9033);
or UO_1002 (O_1002,N_9382,N_9133);
nand UO_1003 (O_1003,N_9964,N_9182);
nand UO_1004 (O_1004,N_9233,N_9157);
xor UO_1005 (O_1005,N_9184,N_9880);
nor UO_1006 (O_1006,N_9287,N_9558);
and UO_1007 (O_1007,N_9020,N_9152);
or UO_1008 (O_1008,N_9771,N_9839);
nand UO_1009 (O_1009,N_9952,N_9239);
xnor UO_1010 (O_1010,N_9982,N_9254);
or UO_1011 (O_1011,N_9610,N_9056);
and UO_1012 (O_1012,N_9948,N_9691);
nand UO_1013 (O_1013,N_9924,N_9641);
xnor UO_1014 (O_1014,N_9753,N_9762);
and UO_1015 (O_1015,N_9628,N_9687);
nand UO_1016 (O_1016,N_9626,N_9814);
xnor UO_1017 (O_1017,N_9508,N_9007);
nand UO_1018 (O_1018,N_9870,N_9347);
nor UO_1019 (O_1019,N_9810,N_9483);
nand UO_1020 (O_1020,N_9179,N_9821);
xnor UO_1021 (O_1021,N_9198,N_9732);
and UO_1022 (O_1022,N_9172,N_9868);
nand UO_1023 (O_1023,N_9883,N_9577);
and UO_1024 (O_1024,N_9564,N_9135);
xor UO_1025 (O_1025,N_9801,N_9288);
nand UO_1026 (O_1026,N_9433,N_9134);
nand UO_1027 (O_1027,N_9100,N_9336);
xor UO_1028 (O_1028,N_9132,N_9095);
nand UO_1029 (O_1029,N_9884,N_9999);
or UO_1030 (O_1030,N_9616,N_9327);
and UO_1031 (O_1031,N_9340,N_9282);
nor UO_1032 (O_1032,N_9294,N_9628);
or UO_1033 (O_1033,N_9101,N_9281);
nor UO_1034 (O_1034,N_9850,N_9849);
nor UO_1035 (O_1035,N_9533,N_9962);
or UO_1036 (O_1036,N_9884,N_9402);
and UO_1037 (O_1037,N_9884,N_9728);
xor UO_1038 (O_1038,N_9488,N_9361);
or UO_1039 (O_1039,N_9025,N_9233);
and UO_1040 (O_1040,N_9948,N_9035);
nand UO_1041 (O_1041,N_9433,N_9423);
nor UO_1042 (O_1042,N_9234,N_9641);
or UO_1043 (O_1043,N_9487,N_9905);
nand UO_1044 (O_1044,N_9412,N_9052);
or UO_1045 (O_1045,N_9236,N_9288);
nand UO_1046 (O_1046,N_9450,N_9672);
nand UO_1047 (O_1047,N_9328,N_9174);
xor UO_1048 (O_1048,N_9473,N_9433);
and UO_1049 (O_1049,N_9083,N_9013);
nor UO_1050 (O_1050,N_9144,N_9239);
nand UO_1051 (O_1051,N_9860,N_9922);
nor UO_1052 (O_1052,N_9145,N_9592);
xor UO_1053 (O_1053,N_9726,N_9385);
nor UO_1054 (O_1054,N_9399,N_9603);
and UO_1055 (O_1055,N_9397,N_9478);
nor UO_1056 (O_1056,N_9278,N_9277);
nand UO_1057 (O_1057,N_9370,N_9456);
or UO_1058 (O_1058,N_9142,N_9717);
or UO_1059 (O_1059,N_9175,N_9942);
and UO_1060 (O_1060,N_9840,N_9068);
xor UO_1061 (O_1061,N_9122,N_9203);
nor UO_1062 (O_1062,N_9033,N_9797);
and UO_1063 (O_1063,N_9409,N_9775);
nand UO_1064 (O_1064,N_9689,N_9215);
xor UO_1065 (O_1065,N_9593,N_9651);
and UO_1066 (O_1066,N_9893,N_9483);
nor UO_1067 (O_1067,N_9092,N_9807);
nand UO_1068 (O_1068,N_9258,N_9643);
or UO_1069 (O_1069,N_9593,N_9392);
or UO_1070 (O_1070,N_9862,N_9267);
xor UO_1071 (O_1071,N_9868,N_9723);
and UO_1072 (O_1072,N_9013,N_9424);
xnor UO_1073 (O_1073,N_9086,N_9366);
nor UO_1074 (O_1074,N_9949,N_9548);
nand UO_1075 (O_1075,N_9056,N_9931);
or UO_1076 (O_1076,N_9487,N_9022);
nand UO_1077 (O_1077,N_9738,N_9049);
nand UO_1078 (O_1078,N_9583,N_9745);
nand UO_1079 (O_1079,N_9831,N_9862);
xnor UO_1080 (O_1080,N_9656,N_9425);
xnor UO_1081 (O_1081,N_9628,N_9511);
nor UO_1082 (O_1082,N_9774,N_9286);
nor UO_1083 (O_1083,N_9739,N_9807);
xnor UO_1084 (O_1084,N_9604,N_9236);
and UO_1085 (O_1085,N_9911,N_9655);
nand UO_1086 (O_1086,N_9460,N_9907);
or UO_1087 (O_1087,N_9000,N_9723);
and UO_1088 (O_1088,N_9016,N_9206);
nor UO_1089 (O_1089,N_9554,N_9172);
nor UO_1090 (O_1090,N_9796,N_9441);
or UO_1091 (O_1091,N_9517,N_9136);
and UO_1092 (O_1092,N_9115,N_9838);
nor UO_1093 (O_1093,N_9639,N_9883);
or UO_1094 (O_1094,N_9454,N_9213);
or UO_1095 (O_1095,N_9071,N_9480);
xnor UO_1096 (O_1096,N_9196,N_9611);
and UO_1097 (O_1097,N_9182,N_9164);
and UO_1098 (O_1098,N_9775,N_9324);
nor UO_1099 (O_1099,N_9397,N_9227);
xor UO_1100 (O_1100,N_9074,N_9659);
nor UO_1101 (O_1101,N_9045,N_9785);
xnor UO_1102 (O_1102,N_9020,N_9255);
xnor UO_1103 (O_1103,N_9304,N_9311);
nand UO_1104 (O_1104,N_9423,N_9520);
xor UO_1105 (O_1105,N_9962,N_9428);
or UO_1106 (O_1106,N_9929,N_9951);
or UO_1107 (O_1107,N_9461,N_9197);
nand UO_1108 (O_1108,N_9879,N_9048);
nand UO_1109 (O_1109,N_9786,N_9634);
xor UO_1110 (O_1110,N_9309,N_9180);
nand UO_1111 (O_1111,N_9135,N_9432);
nor UO_1112 (O_1112,N_9640,N_9379);
nor UO_1113 (O_1113,N_9138,N_9337);
nor UO_1114 (O_1114,N_9146,N_9608);
and UO_1115 (O_1115,N_9466,N_9684);
or UO_1116 (O_1116,N_9285,N_9598);
nor UO_1117 (O_1117,N_9123,N_9091);
xor UO_1118 (O_1118,N_9552,N_9454);
nand UO_1119 (O_1119,N_9896,N_9944);
or UO_1120 (O_1120,N_9806,N_9346);
nor UO_1121 (O_1121,N_9346,N_9931);
nor UO_1122 (O_1122,N_9029,N_9239);
or UO_1123 (O_1123,N_9075,N_9869);
nand UO_1124 (O_1124,N_9403,N_9216);
nand UO_1125 (O_1125,N_9370,N_9958);
or UO_1126 (O_1126,N_9385,N_9064);
or UO_1127 (O_1127,N_9524,N_9742);
and UO_1128 (O_1128,N_9632,N_9373);
nand UO_1129 (O_1129,N_9834,N_9773);
nor UO_1130 (O_1130,N_9103,N_9731);
xnor UO_1131 (O_1131,N_9828,N_9783);
nand UO_1132 (O_1132,N_9340,N_9627);
or UO_1133 (O_1133,N_9697,N_9178);
xnor UO_1134 (O_1134,N_9090,N_9526);
nor UO_1135 (O_1135,N_9963,N_9118);
or UO_1136 (O_1136,N_9691,N_9729);
and UO_1137 (O_1137,N_9856,N_9216);
xnor UO_1138 (O_1138,N_9152,N_9102);
nand UO_1139 (O_1139,N_9100,N_9713);
or UO_1140 (O_1140,N_9011,N_9225);
and UO_1141 (O_1141,N_9174,N_9313);
or UO_1142 (O_1142,N_9263,N_9708);
xor UO_1143 (O_1143,N_9725,N_9357);
or UO_1144 (O_1144,N_9072,N_9572);
nor UO_1145 (O_1145,N_9236,N_9110);
nand UO_1146 (O_1146,N_9327,N_9149);
nor UO_1147 (O_1147,N_9822,N_9731);
or UO_1148 (O_1148,N_9717,N_9247);
and UO_1149 (O_1149,N_9567,N_9717);
nor UO_1150 (O_1150,N_9875,N_9524);
and UO_1151 (O_1151,N_9253,N_9919);
or UO_1152 (O_1152,N_9286,N_9010);
nor UO_1153 (O_1153,N_9775,N_9594);
nand UO_1154 (O_1154,N_9871,N_9748);
or UO_1155 (O_1155,N_9365,N_9054);
and UO_1156 (O_1156,N_9137,N_9204);
and UO_1157 (O_1157,N_9606,N_9253);
and UO_1158 (O_1158,N_9979,N_9368);
or UO_1159 (O_1159,N_9486,N_9047);
nand UO_1160 (O_1160,N_9870,N_9436);
or UO_1161 (O_1161,N_9189,N_9045);
or UO_1162 (O_1162,N_9995,N_9705);
xor UO_1163 (O_1163,N_9331,N_9455);
xor UO_1164 (O_1164,N_9542,N_9490);
nor UO_1165 (O_1165,N_9095,N_9690);
or UO_1166 (O_1166,N_9058,N_9375);
and UO_1167 (O_1167,N_9712,N_9332);
xnor UO_1168 (O_1168,N_9925,N_9996);
xnor UO_1169 (O_1169,N_9076,N_9944);
and UO_1170 (O_1170,N_9208,N_9866);
or UO_1171 (O_1171,N_9491,N_9424);
xnor UO_1172 (O_1172,N_9955,N_9440);
xnor UO_1173 (O_1173,N_9703,N_9858);
or UO_1174 (O_1174,N_9691,N_9376);
xnor UO_1175 (O_1175,N_9036,N_9333);
xor UO_1176 (O_1176,N_9779,N_9272);
nor UO_1177 (O_1177,N_9776,N_9623);
or UO_1178 (O_1178,N_9175,N_9742);
nor UO_1179 (O_1179,N_9325,N_9456);
nand UO_1180 (O_1180,N_9581,N_9611);
or UO_1181 (O_1181,N_9794,N_9614);
nand UO_1182 (O_1182,N_9720,N_9404);
or UO_1183 (O_1183,N_9038,N_9843);
nor UO_1184 (O_1184,N_9495,N_9419);
and UO_1185 (O_1185,N_9830,N_9392);
nor UO_1186 (O_1186,N_9825,N_9390);
and UO_1187 (O_1187,N_9900,N_9559);
nor UO_1188 (O_1188,N_9715,N_9413);
nor UO_1189 (O_1189,N_9566,N_9735);
nand UO_1190 (O_1190,N_9950,N_9054);
nor UO_1191 (O_1191,N_9577,N_9013);
nor UO_1192 (O_1192,N_9014,N_9825);
or UO_1193 (O_1193,N_9794,N_9475);
nand UO_1194 (O_1194,N_9734,N_9130);
nand UO_1195 (O_1195,N_9888,N_9267);
or UO_1196 (O_1196,N_9595,N_9852);
nand UO_1197 (O_1197,N_9857,N_9128);
or UO_1198 (O_1198,N_9868,N_9340);
and UO_1199 (O_1199,N_9511,N_9187);
and UO_1200 (O_1200,N_9972,N_9901);
or UO_1201 (O_1201,N_9419,N_9696);
and UO_1202 (O_1202,N_9980,N_9098);
or UO_1203 (O_1203,N_9554,N_9804);
or UO_1204 (O_1204,N_9866,N_9623);
nand UO_1205 (O_1205,N_9773,N_9333);
nor UO_1206 (O_1206,N_9614,N_9383);
or UO_1207 (O_1207,N_9958,N_9392);
nand UO_1208 (O_1208,N_9205,N_9625);
or UO_1209 (O_1209,N_9828,N_9548);
or UO_1210 (O_1210,N_9783,N_9684);
and UO_1211 (O_1211,N_9412,N_9644);
or UO_1212 (O_1212,N_9271,N_9763);
xnor UO_1213 (O_1213,N_9728,N_9731);
nor UO_1214 (O_1214,N_9176,N_9834);
nor UO_1215 (O_1215,N_9891,N_9594);
nor UO_1216 (O_1216,N_9325,N_9956);
or UO_1217 (O_1217,N_9101,N_9074);
and UO_1218 (O_1218,N_9341,N_9952);
xnor UO_1219 (O_1219,N_9082,N_9370);
nor UO_1220 (O_1220,N_9106,N_9996);
nand UO_1221 (O_1221,N_9107,N_9970);
or UO_1222 (O_1222,N_9949,N_9950);
or UO_1223 (O_1223,N_9973,N_9304);
and UO_1224 (O_1224,N_9224,N_9203);
nor UO_1225 (O_1225,N_9936,N_9130);
and UO_1226 (O_1226,N_9292,N_9624);
nand UO_1227 (O_1227,N_9757,N_9942);
or UO_1228 (O_1228,N_9964,N_9392);
and UO_1229 (O_1229,N_9813,N_9975);
and UO_1230 (O_1230,N_9150,N_9230);
nor UO_1231 (O_1231,N_9266,N_9215);
or UO_1232 (O_1232,N_9390,N_9261);
nand UO_1233 (O_1233,N_9076,N_9440);
xnor UO_1234 (O_1234,N_9931,N_9596);
and UO_1235 (O_1235,N_9792,N_9587);
and UO_1236 (O_1236,N_9772,N_9364);
or UO_1237 (O_1237,N_9936,N_9685);
or UO_1238 (O_1238,N_9173,N_9982);
and UO_1239 (O_1239,N_9781,N_9913);
nor UO_1240 (O_1240,N_9491,N_9317);
nor UO_1241 (O_1241,N_9356,N_9103);
and UO_1242 (O_1242,N_9796,N_9079);
nand UO_1243 (O_1243,N_9557,N_9893);
and UO_1244 (O_1244,N_9746,N_9425);
nand UO_1245 (O_1245,N_9112,N_9571);
or UO_1246 (O_1246,N_9528,N_9911);
nor UO_1247 (O_1247,N_9580,N_9930);
xnor UO_1248 (O_1248,N_9780,N_9131);
or UO_1249 (O_1249,N_9479,N_9669);
nand UO_1250 (O_1250,N_9846,N_9991);
or UO_1251 (O_1251,N_9052,N_9440);
and UO_1252 (O_1252,N_9543,N_9829);
nand UO_1253 (O_1253,N_9120,N_9396);
xor UO_1254 (O_1254,N_9854,N_9736);
and UO_1255 (O_1255,N_9889,N_9928);
or UO_1256 (O_1256,N_9532,N_9390);
and UO_1257 (O_1257,N_9084,N_9639);
or UO_1258 (O_1258,N_9827,N_9517);
nand UO_1259 (O_1259,N_9135,N_9613);
nor UO_1260 (O_1260,N_9310,N_9921);
nand UO_1261 (O_1261,N_9949,N_9123);
nand UO_1262 (O_1262,N_9558,N_9414);
xor UO_1263 (O_1263,N_9153,N_9840);
and UO_1264 (O_1264,N_9327,N_9975);
xnor UO_1265 (O_1265,N_9679,N_9045);
nor UO_1266 (O_1266,N_9787,N_9194);
or UO_1267 (O_1267,N_9149,N_9249);
nor UO_1268 (O_1268,N_9294,N_9920);
and UO_1269 (O_1269,N_9289,N_9237);
nor UO_1270 (O_1270,N_9849,N_9544);
and UO_1271 (O_1271,N_9481,N_9037);
or UO_1272 (O_1272,N_9320,N_9178);
and UO_1273 (O_1273,N_9305,N_9719);
xor UO_1274 (O_1274,N_9623,N_9755);
xor UO_1275 (O_1275,N_9997,N_9877);
nor UO_1276 (O_1276,N_9643,N_9508);
nand UO_1277 (O_1277,N_9784,N_9780);
nor UO_1278 (O_1278,N_9071,N_9153);
or UO_1279 (O_1279,N_9145,N_9240);
or UO_1280 (O_1280,N_9842,N_9961);
and UO_1281 (O_1281,N_9594,N_9499);
nand UO_1282 (O_1282,N_9774,N_9421);
nor UO_1283 (O_1283,N_9335,N_9396);
and UO_1284 (O_1284,N_9849,N_9443);
xor UO_1285 (O_1285,N_9399,N_9376);
and UO_1286 (O_1286,N_9820,N_9078);
xor UO_1287 (O_1287,N_9860,N_9275);
nand UO_1288 (O_1288,N_9711,N_9099);
or UO_1289 (O_1289,N_9466,N_9427);
nor UO_1290 (O_1290,N_9605,N_9943);
nor UO_1291 (O_1291,N_9805,N_9885);
and UO_1292 (O_1292,N_9334,N_9305);
nand UO_1293 (O_1293,N_9318,N_9717);
nor UO_1294 (O_1294,N_9027,N_9224);
or UO_1295 (O_1295,N_9495,N_9143);
or UO_1296 (O_1296,N_9913,N_9012);
or UO_1297 (O_1297,N_9259,N_9405);
nand UO_1298 (O_1298,N_9428,N_9960);
nor UO_1299 (O_1299,N_9206,N_9958);
nor UO_1300 (O_1300,N_9690,N_9887);
or UO_1301 (O_1301,N_9616,N_9116);
and UO_1302 (O_1302,N_9772,N_9675);
or UO_1303 (O_1303,N_9227,N_9363);
or UO_1304 (O_1304,N_9984,N_9189);
and UO_1305 (O_1305,N_9389,N_9188);
xnor UO_1306 (O_1306,N_9585,N_9545);
or UO_1307 (O_1307,N_9331,N_9442);
nor UO_1308 (O_1308,N_9856,N_9434);
nor UO_1309 (O_1309,N_9456,N_9564);
nor UO_1310 (O_1310,N_9033,N_9087);
xor UO_1311 (O_1311,N_9130,N_9371);
or UO_1312 (O_1312,N_9890,N_9856);
xnor UO_1313 (O_1313,N_9337,N_9195);
or UO_1314 (O_1314,N_9049,N_9497);
and UO_1315 (O_1315,N_9369,N_9559);
or UO_1316 (O_1316,N_9627,N_9781);
and UO_1317 (O_1317,N_9328,N_9216);
nor UO_1318 (O_1318,N_9642,N_9102);
nor UO_1319 (O_1319,N_9064,N_9335);
or UO_1320 (O_1320,N_9648,N_9079);
and UO_1321 (O_1321,N_9326,N_9960);
xor UO_1322 (O_1322,N_9404,N_9887);
or UO_1323 (O_1323,N_9803,N_9229);
xor UO_1324 (O_1324,N_9016,N_9431);
or UO_1325 (O_1325,N_9522,N_9214);
nand UO_1326 (O_1326,N_9489,N_9914);
or UO_1327 (O_1327,N_9265,N_9638);
nand UO_1328 (O_1328,N_9714,N_9472);
or UO_1329 (O_1329,N_9815,N_9444);
and UO_1330 (O_1330,N_9610,N_9201);
and UO_1331 (O_1331,N_9268,N_9913);
nand UO_1332 (O_1332,N_9533,N_9613);
xnor UO_1333 (O_1333,N_9935,N_9148);
nand UO_1334 (O_1334,N_9039,N_9197);
and UO_1335 (O_1335,N_9752,N_9119);
xor UO_1336 (O_1336,N_9305,N_9356);
nand UO_1337 (O_1337,N_9165,N_9228);
nand UO_1338 (O_1338,N_9408,N_9988);
nand UO_1339 (O_1339,N_9057,N_9790);
and UO_1340 (O_1340,N_9385,N_9842);
nand UO_1341 (O_1341,N_9323,N_9838);
or UO_1342 (O_1342,N_9945,N_9468);
and UO_1343 (O_1343,N_9932,N_9513);
nor UO_1344 (O_1344,N_9918,N_9956);
nor UO_1345 (O_1345,N_9196,N_9793);
or UO_1346 (O_1346,N_9686,N_9984);
xnor UO_1347 (O_1347,N_9535,N_9658);
nand UO_1348 (O_1348,N_9203,N_9334);
or UO_1349 (O_1349,N_9853,N_9165);
xnor UO_1350 (O_1350,N_9130,N_9318);
nor UO_1351 (O_1351,N_9938,N_9734);
nor UO_1352 (O_1352,N_9016,N_9893);
or UO_1353 (O_1353,N_9783,N_9723);
nor UO_1354 (O_1354,N_9870,N_9072);
nor UO_1355 (O_1355,N_9130,N_9114);
and UO_1356 (O_1356,N_9877,N_9881);
nand UO_1357 (O_1357,N_9531,N_9095);
or UO_1358 (O_1358,N_9191,N_9105);
or UO_1359 (O_1359,N_9504,N_9263);
nand UO_1360 (O_1360,N_9377,N_9195);
or UO_1361 (O_1361,N_9733,N_9259);
nor UO_1362 (O_1362,N_9367,N_9392);
nor UO_1363 (O_1363,N_9051,N_9922);
and UO_1364 (O_1364,N_9851,N_9980);
xnor UO_1365 (O_1365,N_9857,N_9397);
and UO_1366 (O_1366,N_9568,N_9363);
nand UO_1367 (O_1367,N_9340,N_9382);
nand UO_1368 (O_1368,N_9990,N_9576);
or UO_1369 (O_1369,N_9623,N_9786);
nor UO_1370 (O_1370,N_9073,N_9389);
nand UO_1371 (O_1371,N_9084,N_9397);
xor UO_1372 (O_1372,N_9302,N_9398);
nand UO_1373 (O_1373,N_9600,N_9124);
xnor UO_1374 (O_1374,N_9459,N_9304);
xor UO_1375 (O_1375,N_9889,N_9702);
nor UO_1376 (O_1376,N_9571,N_9013);
and UO_1377 (O_1377,N_9458,N_9536);
nand UO_1378 (O_1378,N_9060,N_9079);
and UO_1379 (O_1379,N_9218,N_9244);
and UO_1380 (O_1380,N_9048,N_9846);
nor UO_1381 (O_1381,N_9246,N_9205);
nor UO_1382 (O_1382,N_9571,N_9848);
nor UO_1383 (O_1383,N_9788,N_9659);
and UO_1384 (O_1384,N_9738,N_9852);
nand UO_1385 (O_1385,N_9364,N_9570);
nor UO_1386 (O_1386,N_9934,N_9821);
nor UO_1387 (O_1387,N_9926,N_9259);
and UO_1388 (O_1388,N_9136,N_9801);
nor UO_1389 (O_1389,N_9274,N_9588);
nor UO_1390 (O_1390,N_9246,N_9683);
xnor UO_1391 (O_1391,N_9241,N_9950);
or UO_1392 (O_1392,N_9726,N_9382);
nor UO_1393 (O_1393,N_9269,N_9032);
or UO_1394 (O_1394,N_9631,N_9159);
nor UO_1395 (O_1395,N_9915,N_9507);
nor UO_1396 (O_1396,N_9089,N_9109);
or UO_1397 (O_1397,N_9657,N_9608);
and UO_1398 (O_1398,N_9508,N_9995);
xnor UO_1399 (O_1399,N_9890,N_9351);
nand UO_1400 (O_1400,N_9068,N_9099);
nand UO_1401 (O_1401,N_9134,N_9235);
and UO_1402 (O_1402,N_9144,N_9526);
xnor UO_1403 (O_1403,N_9203,N_9251);
nor UO_1404 (O_1404,N_9582,N_9553);
nand UO_1405 (O_1405,N_9418,N_9293);
nand UO_1406 (O_1406,N_9604,N_9551);
nor UO_1407 (O_1407,N_9219,N_9817);
nand UO_1408 (O_1408,N_9572,N_9767);
nor UO_1409 (O_1409,N_9737,N_9861);
nor UO_1410 (O_1410,N_9304,N_9462);
xnor UO_1411 (O_1411,N_9369,N_9947);
nand UO_1412 (O_1412,N_9272,N_9252);
and UO_1413 (O_1413,N_9494,N_9877);
or UO_1414 (O_1414,N_9441,N_9105);
nand UO_1415 (O_1415,N_9814,N_9407);
or UO_1416 (O_1416,N_9435,N_9335);
nand UO_1417 (O_1417,N_9719,N_9832);
xor UO_1418 (O_1418,N_9652,N_9079);
xnor UO_1419 (O_1419,N_9706,N_9485);
nor UO_1420 (O_1420,N_9037,N_9964);
nand UO_1421 (O_1421,N_9662,N_9644);
and UO_1422 (O_1422,N_9125,N_9641);
nor UO_1423 (O_1423,N_9923,N_9446);
or UO_1424 (O_1424,N_9651,N_9578);
nand UO_1425 (O_1425,N_9703,N_9137);
or UO_1426 (O_1426,N_9121,N_9792);
or UO_1427 (O_1427,N_9002,N_9770);
xnor UO_1428 (O_1428,N_9411,N_9030);
or UO_1429 (O_1429,N_9816,N_9033);
or UO_1430 (O_1430,N_9806,N_9075);
nand UO_1431 (O_1431,N_9663,N_9522);
or UO_1432 (O_1432,N_9654,N_9814);
and UO_1433 (O_1433,N_9579,N_9761);
or UO_1434 (O_1434,N_9537,N_9810);
or UO_1435 (O_1435,N_9421,N_9337);
nor UO_1436 (O_1436,N_9330,N_9088);
or UO_1437 (O_1437,N_9588,N_9190);
nor UO_1438 (O_1438,N_9516,N_9807);
xor UO_1439 (O_1439,N_9628,N_9232);
xor UO_1440 (O_1440,N_9255,N_9159);
and UO_1441 (O_1441,N_9361,N_9248);
xor UO_1442 (O_1442,N_9571,N_9103);
and UO_1443 (O_1443,N_9638,N_9890);
nor UO_1444 (O_1444,N_9849,N_9700);
and UO_1445 (O_1445,N_9637,N_9460);
nand UO_1446 (O_1446,N_9678,N_9992);
nand UO_1447 (O_1447,N_9570,N_9417);
nor UO_1448 (O_1448,N_9370,N_9352);
nor UO_1449 (O_1449,N_9759,N_9373);
or UO_1450 (O_1450,N_9417,N_9938);
or UO_1451 (O_1451,N_9457,N_9600);
nor UO_1452 (O_1452,N_9903,N_9045);
nor UO_1453 (O_1453,N_9485,N_9365);
or UO_1454 (O_1454,N_9454,N_9400);
and UO_1455 (O_1455,N_9868,N_9865);
nand UO_1456 (O_1456,N_9002,N_9453);
or UO_1457 (O_1457,N_9344,N_9867);
or UO_1458 (O_1458,N_9716,N_9128);
and UO_1459 (O_1459,N_9261,N_9616);
nor UO_1460 (O_1460,N_9652,N_9279);
nand UO_1461 (O_1461,N_9780,N_9941);
nand UO_1462 (O_1462,N_9781,N_9174);
nor UO_1463 (O_1463,N_9985,N_9538);
xnor UO_1464 (O_1464,N_9190,N_9523);
nor UO_1465 (O_1465,N_9380,N_9767);
or UO_1466 (O_1466,N_9235,N_9356);
nand UO_1467 (O_1467,N_9954,N_9960);
nand UO_1468 (O_1468,N_9682,N_9994);
and UO_1469 (O_1469,N_9561,N_9492);
or UO_1470 (O_1470,N_9123,N_9066);
or UO_1471 (O_1471,N_9988,N_9459);
and UO_1472 (O_1472,N_9141,N_9218);
nand UO_1473 (O_1473,N_9615,N_9922);
and UO_1474 (O_1474,N_9878,N_9521);
nand UO_1475 (O_1475,N_9372,N_9755);
xnor UO_1476 (O_1476,N_9321,N_9004);
and UO_1477 (O_1477,N_9270,N_9498);
nor UO_1478 (O_1478,N_9768,N_9412);
nor UO_1479 (O_1479,N_9405,N_9102);
and UO_1480 (O_1480,N_9607,N_9062);
nand UO_1481 (O_1481,N_9767,N_9022);
xnor UO_1482 (O_1482,N_9433,N_9179);
or UO_1483 (O_1483,N_9838,N_9216);
xor UO_1484 (O_1484,N_9356,N_9788);
xnor UO_1485 (O_1485,N_9831,N_9858);
and UO_1486 (O_1486,N_9623,N_9297);
nand UO_1487 (O_1487,N_9133,N_9995);
xnor UO_1488 (O_1488,N_9859,N_9545);
nand UO_1489 (O_1489,N_9371,N_9224);
and UO_1490 (O_1490,N_9932,N_9087);
or UO_1491 (O_1491,N_9812,N_9168);
and UO_1492 (O_1492,N_9326,N_9877);
xor UO_1493 (O_1493,N_9872,N_9785);
xnor UO_1494 (O_1494,N_9709,N_9556);
nand UO_1495 (O_1495,N_9628,N_9958);
xnor UO_1496 (O_1496,N_9563,N_9816);
and UO_1497 (O_1497,N_9977,N_9232);
nor UO_1498 (O_1498,N_9277,N_9767);
xnor UO_1499 (O_1499,N_9359,N_9460);
endmodule