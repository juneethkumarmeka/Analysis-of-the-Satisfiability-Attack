module basic_3000_30000_3500_10_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_1939,In_1688);
xnor U1 (N_1,In_1025,In_612);
and U2 (N_2,In_2722,In_52);
and U3 (N_3,In_1525,In_2428);
or U4 (N_4,In_341,In_68);
or U5 (N_5,In_727,In_2996);
xnor U6 (N_6,In_2660,In_2066);
nor U7 (N_7,In_1529,In_1030);
xnor U8 (N_8,In_951,In_2739);
nor U9 (N_9,In_243,In_1217);
and U10 (N_10,In_1651,In_1458);
and U11 (N_11,In_2619,In_639);
or U12 (N_12,In_1763,In_2122);
and U13 (N_13,In_1463,In_495);
and U14 (N_14,In_1656,In_366);
nand U15 (N_15,In_787,In_1068);
nand U16 (N_16,In_93,In_784);
nor U17 (N_17,In_1003,In_633);
and U18 (N_18,In_2152,In_1330);
xnor U19 (N_19,In_1565,In_1409);
or U20 (N_20,In_851,In_172);
xnor U21 (N_21,In_1846,In_1363);
nand U22 (N_22,In_2933,In_979);
and U23 (N_23,In_2541,In_21);
nor U24 (N_24,In_1119,In_585);
or U25 (N_25,In_34,In_2671);
and U26 (N_26,In_2178,In_2772);
nor U27 (N_27,In_1252,In_1956);
xor U28 (N_28,In_2733,In_2507);
and U29 (N_29,In_2738,In_872);
nor U30 (N_30,In_2506,In_1289);
or U31 (N_31,In_1157,In_1934);
xnor U32 (N_32,In_1608,In_967);
xor U33 (N_33,In_2342,In_2862);
or U34 (N_34,In_1537,In_819);
nor U35 (N_35,In_1876,In_2576);
nor U36 (N_36,In_316,In_2447);
or U37 (N_37,In_565,In_2692);
and U38 (N_38,In_2670,In_652);
and U39 (N_39,In_1914,In_2972);
xor U40 (N_40,In_922,In_328);
nand U41 (N_41,In_1977,In_168);
xnor U42 (N_42,In_25,In_2238);
or U43 (N_43,In_1169,In_392);
nand U44 (N_44,In_1309,In_2821);
and U45 (N_45,In_467,In_2638);
and U46 (N_46,In_1239,In_1307);
and U47 (N_47,In_996,In_379);
nor U48 (N_48,In_2715,In_2640);
nand U49 (N_49,In_337,In_55);
nor U50 (N_50,In_444,In_2899);
nand U51 (N_51,In_1667,In_715);
or U52 (N_52,In_1556,In_1898);
nand U53 (N_53,In_1933,In_1559);
and U54 (N_54,In_1474,In_696);
nor U55 (N_55,In_14,In_2809);
or U56 (N_56,In_2091,In_2557);
nor U57 (N_57,In_2269,In_1641);
or U58 (N_58,In_2040,In_1418);
or U59 (N_59,In_1820,In_892);
and U60 (N_60,In_2317,In_2486);
nand U61 (N_61,In_1261,In_2526);
xor U62 (N_62,In_2031,In_649);
and U63 (N_63,In_188,In_788);
and U64 (N_64,In_2811,In_1685);
xor U65 (N_65,In_2748,In_1508);
nand U66 (N_66,In_192,In_2088);
and U67 (N_67,In_1633,In_1298);
nand U68 (N_68,In_1429,In_2525);
or U69 (N_69,In_2184,In_2490);
xnor U70 (N_70,In_213,In_1316);
xor U71 (N_71,In_2661,In_1387);
or U72 (N_72,In_704,In_1327);
nor U73 (N_73,In_609,In_1493);
and U74 (N_74,In_1832,In_1069);
xnor U75 (N_75,In_669,In_2052);
xnor U76 (N_76,In_57,In_2193);
nor U77 (N_77,In_2650,In_296);
or U78 (N_78,In_1897,In_738);
nor U79 (N_79,In_2014,In_1737);
xnor U80 (N_80,In_474,In_2888);
and U81 (N_81,In_1008,In_1658);
nor U82 (N_82,In_91,In_1669);
xor U83 (N_83,In_2844,In_1645);
and U84 (N_84,In_1142,In_613);
nor U85 (N_85,In_2243,In_2310);
nor U86 (N_86,In_1097,In_2832);
nor U87 (N_87,In_1968,In_1657);
nor U88 (N_88,In_1627,In_147);
nand U89 (N_89,In_1332,In_2968);
xnor U90 (N_90,In_1014,In_1432);
xor U91 (N_91,In_961,In_1713);
nor U92 (N_92,In_1166,In_1890);
xnor U93 (N_93,In_2104,In_1719);
xor U94 (N_94,In_969,In_809);
nand U95 (N_95,In_126,In_70);
or U96 (N_96,In_2339,In_638);
or U97 (N_97,In_1718,In_112);
or U98 (N_98,In_1563,In_754);
and U99 (N_99,In_2927,In_252);
and U100 (N_100,In_2582,In_975);
and U101 (N_101,In_1882,In_1450);
nor U102 (N_102,In_1400,In_1866);
xnor U103 (N_103,In_582,In_1365);
nand U104 (N_104,In_596,In_1297);
and U105 (N_105,In_373,In_2118);
or U106 (N_106,In_2792,In_2964);
or U107 (N_107,In_1185,In_463);
and U108 (N_108,In_1466,In_2390);
nand U109 (N_109,In_1736,In_166);
xnor U110 (N_110,In_1510,In_1195);
and U111 (N_111,In_1597,In_2286);
xor U112 (N_112,In_1457,In_2227);
and U113 (N_113,In_1990,In_960);
and U114 (N_114,In_2075,In_1946);
and U115 (N_115,In_229,In_2094);
xnor U116 (N_116,In_2699,In_939);
xor U117 (N_117,In_823,In_1740);
nor U118 (N_118,In_778,In_1112);
or U119 (N_119,In_2553,In_2041);
and U120 (N_120,In_2319,In_2986);
or U121 (N_121,In_2536,In_2190);
and U122 (N_122,In_2298,In_496);
and U123 (N_123,In_482,In_2765);
and U124 (N_124,In_1237,In_2998);
nor U125 (N_125,In_2300,In_390);
nand U126 (N_126,In_2420,In_553);
xor U127 (N_127,In_1912,In_2658);
or U128 (N_128,In_2157,In_1935);
and U129 (N_129,In_121,In_2177);
xor U130 (N_130,In_362,In_2645);
and U131 (N_131,In_154,In_2908);
xor U132 (N_132,In_2201,In_2039);
nor U133 (N_133,In_817,In_1838);
nor U134 (N_134,In_483,In_2835);
xor U135 (N_135,In_1588,In_1285);
or U136 (N_136,In_1984,In_792);
xnor U137 (N_137,In_814,In_1147);
or U138 (N_138,In_916,In_2247);
and U139 (N_139,In_2433,In_1481);
nor U140 (N_140,In_1753,In_1581);
nand U141 (N_141,In_400,In_2199);
and U142 (N_142,In_48,In_1377);
nor U143 (N_143,In_2381,In_2947);
xor U144 (N_144,In_458,In_679);
or U145 (N_145,In_2338,In_689);
nand U146 (N_146,In_2641,In_1374);
nand U147 (N_147,In_730,In_2105);
and U148 (N_148,In_271,In_2124);
nand U149 (N_149,In_2939,In_2234);
xnor U150 (N_150,In_2022,In_569);
nand U151 (N_151,In_2736,In_1706);
nand U152 (N_152,In_2489,In_2814);
or U153 (N_153,In_2538,In_163);
xor U154 (N_154,In_557,In_2782);
nor U155 (N_155,In_1089,In_2050);
and U156 (N_156,In_1773,In_937);
nand U157 (N_157,In_1471,In_1498);
xnor U158 (N_158,In_2878,In_1501);
nand U159 (N_159,In_2130,In_1206);
xor U160 (N_160,In_1945,In_773);
xnor U161 (N_161,In_140,In_1333);
nor U162 (N_162,In_2728,In_2027);
nor U163 (N_163,In_842,In_2614);
xor U164 (N_164,In_1547,In_1200);
or U165 (N_165,In_1507,In_2980);
or U166 (N_166,In_2801,In_1057);
or U167 (N_167,In_1433,In_64);
xnor U168 (N_168,In_303,In_1007);
or U169 (N_169,In_957,In_2587);
nor U170 (N_170,In_1861,In_333);
nand U171 (N_171,In_374,In_102);
xnor U172 (N_172,In_554,In_1385);
and U173 (N_173,In_1328,In_1545);
nand U174 (N_174,In_2076,In_1262);
or U175 (N_175,In_436,In_1682);
xnor U176 (N_176,In_220,In_528);
and U177 (N_177,In_254,In_830);
xor U178 (N_178,In_912,In_2200);
and U179 (N_179,In_1465,In_348);
and U180 (N_180,In_2643,In_2720);
and U181 (N_181,In_2713,In_1350);
xor U182 (N_182,In_340,In_2404);
or U183 (N_183,In_1275,In_1910);
nor U184 (N_184,In_1870,In_1610);
nand U185 (N_185,In_505,In_1175);
and U186 (N_186,In_2848,In_875);
nand U187 (N_187,In_850,In_2176);
nor U188 (N_188,In_1437,In_2037);
and U189 (N_189,In_2858,In_802);
xnor U190 (N_190,In_1542,In_1128);
and U191 (N_191,In_591,In_2465);
and U192 (N_192,In_277,In_1416);
and U193 (N_193,In_2999,In_29);
nor U194 (N_194,In_1534,In_2818);
nor U195 (N_195,In_712,In_1360);
or U196 (N_196,In_424,In_1145);
and U197 (N_197,In_865,In_991);
nand U198 (N_198,In_2329,In_201);
or U199 (N_199,In_867,In_2611);
xnor U200 (N_200,In_2916,In_143);
or U201 (N_201,In_428,In_107);
and U202 (N_202,In_309,In_2563);
nand U203 (N_203,In_401,In_2551);
xor U204 (N_204,In_2846,In_2002);
xor U205 (N_205,In_2254,In_96);
nor U206 (N_206,In_2235,In_1406);
xor U207 (N_207,In_748,In_906);
nand U208 (N_208,In_510,In_191);
xnor U209 (N_209,In_2546,In_2241);
nand U210 (N_210,In_1562,In_2861);
nor U211 (N_211,In_2875,In_2886);
and U212 (N_212,In_1911,In_903);
nand U213 (N_213,In_2470,In_2029);
nand U214 (N_214,In_1830,In_283);
xor U215 (N_215,In_2758,In_2753);
or U216 (N_216,In_1967,In_1511);
and U217 (N_217,In_2940,In_2911);
nor U218 (N_218,In_2552,In_186);
xor U219 (N_219,In_2555,In_464);
nand U220 (N_220,In_786,In_2478);
nor U221 (N_221,In_425,In_2706);
and U222 (N_222,In_2141,In_1249);
or U223 (N_223,In_816,In_1628);
xnor U224 (N_224,In_1908,In_1954);
and U225 (N_225,In_2543,In_2994);
xor U226 (N_226,In_1174,In_2891);
nand U227 (N_227,In_2828,In_1615);
nand U228 (N_228,In_326,In_776);
or U229 (N_229,In_1010,In_964);
nand U230 (N_230,In_2539,In_16);
xnor U231 (N_231,In_2085,In_2293);
and U232 (N_232,In_1248,In_62);
nor U233 (N_233,In_406,In_1517);
and U234 (N_234,In_1447,In_677);
nor U235 (N_235,In_1806,In_1855);
nand U236 (N_236,In_2098,In_455);
nand U237 (N_237,In_196,In_329);
nand U238 (N_238,In_1282,In_4);
and U239 (N_239,In_1819,In_935);
xnor U240 (N_240,In_2600,In_1013);
nand U241 (N_241,In_1835,In_1674);
xnor U242 (N_242,In_2082,In_448);
or U243 (N_243,In_2630,In_2982);
nand U244 (N_244,In_1579,In_1136);
nand U245 (N_245,In_821,In_2790);
xor U246 (N_246,In_993,In_2522);
xnor U247 (N_247,In_1788,In_2570);
nand U248 (N_248,In_2497,In_1616);
xnor U249 (N_249,In_176,In_1428);
and U250 (N_250,In_2496,In_255);
and U251 (N_251,In_1050,In_80);
xor U252 (N_252,In_2977,In_688);
xnor U253 (N_253,In_2174,In_1865);
or U254 (N_254,In_2359,In_918);
and U255 (N_255,In_459,In_2416);
xor U256 (N_256,In_1514,In_2573);
nor U257 (N_257,In_159,In_2784);
nor U258 (N_258,In_394,In_2492);
or U259 (N_259,In_76,In_1344);
nor U260 (N_260,In_881,In_2033);
and U261 (N_261,In_952,In_1555);
or U262 (N_262,In_828,In_1549);
nor U263 (N_263,In_1390,In_116);
nand U264 (N_264,In_1825,In_1770);
or U265 (N_265,In_1162,In_2625);
nand U266 (N_266,In_260,In_2482);
and U267 (N_267,In_2501,In_2687);
and U268 (N_268,In_1994,In_2912);
nor U269 (N_269,In_295,In_1840);
and U270 (N_270,In_71,In_1741);
nand U271 (N_271,In_2139,In_1461);
or U272 (N_272,In_1294,In_2441);
nand U273 (N_273,In_477,In_2314);
or U274 (N_274,In_2766,In_2328);
nor U275 (N_275,In_1280,In_2019);
xor U276 (N_276,In_1302,In_2866);
nor U277 (N_277,In_1623,In_2213);
or U278 (N_278,In_2867,In_2363);
xor U279 (N_279,In_2915,In_1696);
nor U280 (N_280,In_1611,In_938);
nand U281 (N_281,In_1270,In_1495);
or U282 (N_282,In_2936,In_217);
nand U283 (N_283,In_1448,In_2787);
or U284 (N_284,In_485,In_1075);
or U285 (N_285,In_1171,In_240);
xor U286 (N_286,In_1973,In_2684);
nor U287 (N_287,In_1422,In_1520);
xor U288 (N_288,In_2353,In_2921);
or U289 (N_289,In_134,In_1342);
and U290 (N_290,In_1196,In_2869);
or U291 (N_291,In_1178,In_2385);
nor U292 (N_292,In_1619,In_1454);
nor U293 (N_293,In_281,In_2392);
nor U294 (N_294,In_607,In_1675);
nand U295 (N_295,In_685,In_54);
xnor U296 (N_296,In_2112,In_962);
and U297 (N_297,In_2966,In_454);
and U298 (N_298,In_1004,In_1205);
xor U299 (N_299,In_1922,In_783);
nand U300 (N_300,In_2150,In_123);
nand U301 (N_301,In_1681,In_396);
and U302 (N_302,In_2841,In_2877);
and U303 (N_303,In_1412,In_2705);
nor U304 (N_304,In_1937,In_1612);
and U305 (N_305,In_620,In_2907);
xnor U306 (N_306,In_2704,In_1634);
and U307 (N_307,In_2820,In_1444);
nand U308 (N_308,In_301,In_1101);
or U309 (N_309,In_2457,In_2698);
or U310 (N_310,In_2799,In_2905);
or U311 (N_311,In_1218,In_2920);
nor U312 (N_312,In_987,In_2580);
and U313 (N_313,In_339,In_835);
and U314 (N_314,In_731,In_1293);
and U315 (N_315,In_1276,In_1841);
and U316 (N_316,In_2356,In_2454);
nor U317 (N_317,In_642,In_1163);
nor U318 (N_318,In_1626,In_2581);
xor U319 (N_319,In_2599,In_2718);
or U320 (N_320,In_1067,In_775);
xor U321 (N_321,In_1426,In_195);
and U322 (N_322,In_1022,In_2396);
xor U323 (N_323,In_1601,In_799);
and U324 (N_324,In_59,In_291);
xnor U325 (N_325,In_793,In_930);
and U326 (N_326,In_429,In_367);
or U327 (N_327,In_2413,In_65);
nand U328 (N_328,In_1644,In_1228);
nand U329 (N_329,In_1519,In_1655);
nor U330 (N_330,In_101,In_921);
or U331 (N_331,In_2185,In_2004);
xnor U332 (N_332,In_494,In_846);
xor U333 (N_333,In_1345,In_353);
nor U334 (N_334,In_752,In_2579);
or U335 (N_335,In_1900,In_1703);
nor U336 (N_336,In_469,In_1234);
nand U337 (N_337,In_2086,In_1769);
and U338 (N_338,In_2802,In_1561);
nor U339 (N_339,In_1269,In_2012);
and U340 (N_340,In_2726,In_1358);
nand U341 (N_341,In_1575,In_162);
or U342 (N_342,In_1460,In_2565);
nor U343 (N_343,In_2252,In_2596);
xor U344 (N_344,In_99,In_2932);
nand U345 (N_345,In_409,In_2471);
and U346 (N_346,In_1931,In_2341);
and U347 (N_347,In_1240,In_2078);
or U348 (N_348,In_2776,In_393);
nor U349 (N_349,In_313,In_882);
xor U350 (N_350,In_125,In_2475);
or U351 (N_351,In_1528,In_2276);
nand U352 (N_352,In_1981,In_1009);
nand U353 (N_353,In_2265,In_659);
xnor U354 (N_354,In_692,In_1993);
or U355 (N_355,In_2610,In_1739);
nor U356 (N_356,In_1420,In_1326);
xnor U357 (N_357,In_1180,In_334);
xnor U358 (N_358,In_114,In_1410);
nor U359 (N_359,In_2226,In_2446);
nand U360 (N_360,In_431,In_796);
nor U361 (N_361,In_173,In_1791);
and U362 (N_362,In_770,In_2080);
or U363 (N_363,In_2863,In_760);
or U364 (N_364,In_2663,In_1662);
nor U365 (N_365,In_1164,In_1782);
or U366 (N_366,In_2384,In_1860);
or U367 (N_367,In_780,In_288);
xor U368 (N_368,In_2332,In_1723);
xor U369 (N_369,In_2026,In_2271);
nor U370 (N_370,In_2079,In_322);
or U371 (N_371,In_656,In_2134);
nand U372 (N_372,In_174,In_1539);
or U373 (N_373,In_1607,In_2438);
nor U374 (N_374,In_263,In_2347);
nand U375 (N_375,In_1296,In_2791);
or U376 (N_376,In_1076,In_1661);
nor U377 (N_377,In_115,In_2096);
or U378 (N_378,In_578,In_3);
xnor U379 (N_379,In_269,In_108);
xor U380 (N_380,In_1571,In_88);
nor U381 (N_381,In_994,In_2623);
nor U382 (N_382,In_858,In_516);
nor U383 (N_383,In_1807,In_2230);
nand U384 (N_384,In_2043,In_1490);
nor U385 (N_385,In_1181,In_878);
or U386 (N_386,In_488,In_437);
nor U387 (N_387,In_2400,In_2974);
or U388 (N_388,In_1038,In_315);
nor U389 (N_389,In_1268,In_910);
nor U390 (N_390,In_1334,In_2188);
or U391 (N_391,In_1045,In_210);
or U392 (N_392,In_1710,In_1417);
nor U393 (N_393,In_2196,In_2087);
nor U394 (N_394,In_2380,In_2387);
nand U395 (N_395,In_2402,In_2852);
and U396 (N_396,In_2215,In_2516);
nor U397 (N_397,In_2405,In_2263);
nand U398 (N_398,In_2559,In_2398);
nor U399 (N_399,In_2827,In_502);
or U400 (N_400,In_1382,In_2280);
and U401 (N_401,In_519,In_800);
and U402 (N_402,In_2352,In_2111);
nand U403 (N_403,In_2153,In_1589);
or U404 (N_404,In_1021,In_1541);
or U405 (N_405,In_83,In_2969);
or U406 (N_406,In_310,In_1857);
or U407 (N_407,In_757,In_1856);
xnor U408 (N_408,In_2755,In_531);
or U409 (N_409,In_1227,In_2311);
nand U410 (N_410,In_2132,In_1489);
and U411 (N_411,In_1484,In_2011);
nand U412 (N_412,In_657,In_2255);
and U413 (N_413,In_1256,In_2373);
xnor U414 (N_414,In_130,In_1639);
nor U415 (N_415,In_2953,In_2742);
nand U416 (N_416,In_1585,In_2952);
nand U417 (N_417,In_2805,In_1082);
or U418 (N_418,In_2935,In_1734);
nor U419 (N_419,In_2549,In_1810);
or U420 (N_420,In_1877,In_1780);
xor U421 (N_421,In_695,In_476);
and U422 (N_422,In_518,In_2880);
nand U423 (N_423,In_1324,In_1138);
nor U424 (N_424,In_1436,In_265);
nand U425 (N_425,In_874,In_1431);
xnor U426 (N_426,In_2922,In_2369);
nor U427 (N_427,In_2180,In_282);
nand U428 (N_428,In_1957,In_1847);
nor U429 (N_429,In_1532,In_2288);
nand U430 (N_430,In_2236,In_1636);
nor U431 (N_431,In_28,In_2147);
nand U432 (N_432,In_2597,In_1137);
or U433 (N_433,In_703,In_1586);
nand U434 (N_434,In_661,In_2700);
and U435 (N_435,In_204,In_1808);
and U436 (N_436,In_1812,In_2943);
nand U437 (N_437,In_1516,In_873);
and U438 (N_438,In_1574,In_2509);
or U439 (N_439,In_2125,In_909);
xor U440 (N_440,In_1843,In_1873);
or U441 (N_441,In_626,In_2449);
and U442 (N_442,In_811,In_1331);
and U443 (N_443,In_901,In_2895);
and U444 (N_444,In_2556,In_1944);
nor U445 (N_445,In_2198,In_2307);
nor U446 (N_446,In_1972,In_1060);
xor U447 (N_447,In_415,In_2006);
nor U448 (N_448,In_699,In_2146);
and U449 (N_449,In_2696,In_87);
and U450 (N_450,In_2128,In_1915);
nor U451 (N_451,In_2393,In_1051);
nand U452 (N_452,In_2309,In_2762);
nor U453 (N_453,In_2204,In_237);
nor U454 (N_454,In_1566,In_2017);
nand U455 (N_455,In_1952,In_1242);
nand U456 (N_456,In_1290,In_2868);
and U457 (N_457,In_1800,In_2429);
nand U458 (N_458,In_2788,In_561);
nand U459 (N_459,In_462,In_1462);
and U460 (N_460,In_2183,In_1043);
and U461 (N_461,In_785,In_2464);
nand U462 (N_462,In_250,In_129);
or U463 (N_463,In_1872,In_1434);
nor U464 (N_464,In_79,In_53);
or U465 (N_465,In_297,In_2383);
and U466 (N_466,In_427,In_2833);
or U467 (N_467,In_1833,In_526);
xor U468 (N_468,In_1692,In_1621);
and U469 (N_469,In_1907,In_1700);
xor U470 (N_470,In_2847,In_2695);
xnor U471 (N_471,In_149,In_2481);
nor U472 (N_472,In_2217,In_122);
or U473 (N_473,In_1613,In_1322);
nand U474 (N_474,In_2030,In_2535);
nand U475 (N_475,In_1047,In_1362);
nand U476 (N_476,In_289,In_349);
xnor U477 (N_477,In_1165,In_1092);
and U478 (N_478,In_2750,In_2681);
xor U479 (N_479,In_258,In_1208);
and U480 (N_480,In_503,In_2930);
or U481 (N_481,In_2926,In_2637);
nor U482 (N_482,In_2620,In_1314);
nor U483 (N_483,In_1499,In_398);
nor U484 (N_484,In_2773,In_1243);
nor U485 (N_485,In_1504,In_2519);
xnor U486 (N_486,In_199,In_1062);
and U487 (N_487,In_2914,In_1384);
nor U488 (N_488,In_801,In_2160);
nor U489 (N_489,In_152,In_2896);
nand U490 (N_490,In_643,In_959);
and U491 (N_491,In_128,In_2137);
and U492 (N_492,In_151,In_1347);
or U493 (N_493,In_997,In_2547);
and U494 (N_494,In_2499,In_1824);
nor U495 (N_495,In_1582,In_610);
or U496 (N_496,In_2389,In_625);
xnor U497 (N_497,In_2068,In_1874);
and U498 (N_498,In_2770,In_2382);
xor U499 (N_499,In_2440,In_2355);
nor U500 (N_500,In_691,In_559);
and U501 (N_501,In_2010,In_1222);
xor U502 (N_502,In_1727,In_1829);
xor U503 (N_503,In_1839,In_1997);
xor U504 (N_504,In_728,In_2919);
nor U505 (N_505,In_1609,In_2114);
or U506 (N_506,In_2524,In_751);
or U507 (N_507,In_897,In_1368);
or U508 (N_508,In_1353,In_2095);
or U509 (N_509,In_2343,In_848);
or U510 (N_510,In_532,In_617);
xnor U511 (N_511,In_1690,In_759);
xnor U512 (N_512,In_1966,In_713);
and U513 (N_513,In_798,In_2657);
and U514 (N_514,In_2368,In_223);
and U515 (N_515,In_2437,In_1054);
nand U516 (N_516,In_1652,In_2377);
xnor U517 (N_517,In_1926,In_347);
and U518 (N_518,In_2768,In_234);
and U519 (N_519,In_2444,In_2194);
nand U520 (N_520,In_2839,In_219);
nor U521 (N_521,In_2606,In_2156);
nor U522 (N_522,In_806,In_546);
nor U523 (N_523,In_131,In_2469);
xor U524 (N_524,In_2604,In_774);
xnor U525 (N_525,In_667,In_36);
and U526 (N_526,In_998,In_222);
nor U527 (N_527,In_1969,In_2305);
nor U528 (N_528,In_733,In_640);
nor U529 (N_529,In_779,In_646);
nand U530 (N_530,In_2432,In_2609);
nand U531 (N_531,In_480,In_43);
nor U532 (N_532,In_2505,In_847);
nor U533 (N_533,In_1711,In_844);
or U534 (N_534,In_1291,In_33);
xnor U535 (N_535,In_389,In_2775);
nand U536 (N_536,In_913,In_2729);
and U537 (N_537,In_820,In_2436);
nor U538 (N_538,In_305,In_580);
and U539 (N_539,In_2583,In_1049);
or U540 (N_540,In_2879,In_1213);
nand U541 (N_541,In_272,In_1407);
nor U542 (N_542,In_750,In_2060);
nor U543 (N_543,In_1886,In_1959);
or U544 (N_544,In_1265,In_38);
and U545 (N_545,In_898,In_1073);
nand U546 (N_546,In_2067,In_631);
nand U547 (N_547,In_259,In_2540);
or U548 (N_548,In_2817,In_1435);
or U549 (N_549,In_1446,In_724);
and U550 (N_550,In_1445,In_1127);
or U551 (N_551,In_2162,In_672);
nor U552 (N_552,In_1339,In_2003);
nor U553 (N_553,In_104,In_1392);
or U554 (N_554,In_2677,In_1721);
xor U555 (N_555,In_629,In_1475);
nor U556 (N_556,In_1982,In_1918);
or U557 (N_557,In_1456,In_1975);
or U558 (N_558,In_914,In_791);
nand U559 (N_559,In_10,In_2714);
and U560 (N_560,In_189,In_244);
and U561 (N_561,In_1088,In_61);
nor U562 (N_562,In_1887,In_746);
nor U563 (N_563,In_323,In_1625);
nor U564 (N_564,In_419,In_1123);
xor U565 (N_565,In_1849,In_2688);
nor U566 (N_566,In_1033,In_1733);
or U567 (N_567,In_233,In_2533);
nor U568 (N_568,In_2511,In_2351);
nor U569 (N_569,In_293,In_1452);
xor U570 (N_570,In_1006,In_1863);
nand U571 (N_571,In_11,In_1821);
xnor U572 (N_572,In_988,In_2732);
or U573 (N_573,In_1424,In_2498);
or U574 (N_574,In_1978,In_2090);
nor U575 (N_575,In_1176,In_211);
nor U576 (N_576,In_2774,In_1179);
xor U577 (N_577,In_529,In_1002);
nor U578 (N_578,In_829,In_622);
xnor U579 (N_579,In_2744,In_2316);
or U580 (N_580,In_701,In_1151);
and U581 (N_581,In_2965,In_2143);
nor U582 (N_582,In_2544,In_2297);
or U583 (N_583,In_2617,In_2070);
and U584 (N_584,In_161,In_2047);
xnor U585 (N_585,In_551,In_575);
xor U586 (N_586,In_744,In_2906);
nand U587 (N_587,In_2036,In_2894);
and U588 (N_588,In_212,In_635);
or U589 (N_589,In_2169,In_1987);
and U590 (N_590,In_1671,In_1593);
and U591 (N_591,In_680,In_1543);
nor U592 (N_592,In_2508,In_944);
nor U593 (N_593,In_1845,In_2159);
xor U594 (N_594,In_249,In_264);
nand U595 (N_595,In_2530,In_584);
xor U596 (N_596,In_1683,In_1746);
and U597 (N_597,In_2431,In_2595);
or U598 (N_598,In_1913,In_369);
or U599 (N_599,In_853,In_2371);
and U600 (N_600,In_1190,In_2745);
nor U601 (N_601,In_2675,In_2290);
xnor U602 (N_602,In_611,In_84);
nand U603 (N_603,In_955,In_1184);
or U604 (N_604,In_1816,In_683);
and U605 (N_605,In_2394,In_1235);
or U606 (N_606,In_2636,In_2283);
or U607 (N_607,In_1509,In_2166);
nor U608 (N_608,In_226,In_2819);
nor U609 (N_609,In_2206,In_1225);
and U610 (N_610,In_1283,In_852);
xor U611 (N_611,In_558,In_2910);
nor U612 (N_612,In_662,In_717);
nand U613 (N_613,In_2616,In_280);
xor U614 (N_614,In_202,In_117);
nor U615 (N_615,In_2992,In_682);
nand U616 (N_616,In_971,In_2365);
nand U617 (N_617,In_1263,In_342);
or U618 (N_618,In_1879,In_137);
nand U619 (N_619,In_2257,In_634);
nand U620 (N_620,In_1771,In_1895);
or U621 (N_621,In_552,In_378);
nor U622 (N_622,In_2115,In_2948);
xnor U623 (N_623,In_2218,In_1798);
and U624 (N_624,In_178,In_1480);
xnor U625 (N_625,In_2534,In_1790);
or U626 (N_626,In_1958,In_522);
xnor U627 (N_627,In_1538,In_2691);
xnor U628 (N_628,In_2256,In_513);
xnor U629 (N_629,In_499,In_207);
and U630 (N_630,In_2284,In_1451);
or U631 (N_631,In_1858,In_1526);
or U632 (N_632,In_2399,In_1844);
xor U633 (N_633,In_1354,In_2119);
xnor U634 (N_634,In_1366,In_2264);
nor U635 (N_635,In_615,In_2051);
nand U636 (N_636,In_1469,In_302);
xor U637 (N_637,In_402,In_676);
and U638 (N_638,In_769,In_737);
and U639 (N_639,In_1287,In_1310);
xor U640 (N_640,In_2192,In_862);
nand U641 (N_641,In_2326,In_1513);
nand U642 (N_642,In_2512,In_2673);
nor U643 (N_643,In_1230,In_236);
and U644 (N_644,In_410,In_452);
or U645 (N_645,In_2484,In_1074);
xnor U646 (N_646,In_2191,In_37);
xor U647 (N_647,In_2308,In_741);
nor U648 (N_648,In_268,In_1916);
xnor U649 (N_649,In_2120,In_535);
xor U650 (N_650,In_60,In_1961);
and U651 (N_651,In_1284,In_537);
nand U652 (N_652,In_637,In_2973);
nand U653 (N_653,In_1531,In_2842);
nand U654 (N_654,In_1735,In_1319);
nand U655 (N_655,In_2995,In_2375);
and U656 (N_656,In_2292,In_2142);
or U657 (N_657,In_2584,In_2796);
and U658 (N_658,In_148,In_2967);
and U659 (N_659,In_225,In_1722);
or U660 (N_660,In_2427,In_19);
nand U661 (N_661,In_2334,In_753);
nor U662 (N_662,In_139,In_2335);
and U663 (N_663,In_2322,In_2652);
nand U664 (N_664,In_1815,In_1321);
xnor U665 (N_665,In_456,In_376);
nor U666 (N_666,In_2406,In_965);
nand U667 (N_667,In_2572,In_435);
or U668 (N_668,In_2391,In_1094);
nand U669 (N_669,In_550,In_2344);
nor U670 (N_670,In_2741,In_896);
xor U671 (N_671,In_1580,In_2884);
or U672 (N_672,In_67,In_2165);
and U673 (N_673,In_1090,In_1881);
nand U674 (N_674,In_2321,In_2330);
xnor U675 (N_675,In_2195,In_274);
and U676 (N_676,In_1246,In_1459);
xnor U677 (N_677,In_97,In_1963);
xor U678 (N_678,In_1415,In_136);
or U679 (N_679,In_90,In_387);
nor U680 (N_680,In_833,In_1095);
nand U681 (N_681,In_2889,In_146);
and U682 (N_682,In_2461,In_2229);
xnor U683 (N_683,In_15,In_1325);
nor U684 (N_684,In_2487,In_999);
nor U685 (N_685,In_257,In_1726);
nor U686 (N_686,In_628,In_2532);
or U687 (N_687,In_797,In_890);
nor U688 (N_688,In_1399,In_2361);
or U689 (N_689,In_838,In_2740);
nor U690 (N_690,In_193,In_1427);
or U691 (N_691,In_1640,In_650);
nor U692 (N_692,In_894,In_2354);
xnor U693 (N_693,In_2567,In_399);
nand U694 (N_694,In_1197,In_1998);
and U695 (N_695,In_2598,In_2900);
xnor U696 (N_696,In_423,In_2483);
and U697 (N_697,In_1383,In_1241);
nor U698 (N_698,In_1107,In_2529);
and U699 (N_699,In_1056,In_1453);
xnor U700 (N_700,In_1425,In_2350);
or U701 (N_701,In_1139,In_1204);
nor U702 (N_702,In_2209,In_1730);
nor U703 (N_703,In_1691,In_1869);
nor U704 (N_704,In_205,In_1058);
xor U705 (N_705,In_1889,In_2345);
and U706 (N_706,In_2395,In_31);
nand U707 (N_707,In_2261,In_1943);
nand U708 (N_708,In_855,In_356);
and U709 (N_709,In_782,In_138);
nand U710 (N_710,In_1629,In_2591);
or U711 (N_711,In_215,In_2561);
nor U712 (N_712,In_899,In_1605);
nor U713 (N_713,In_238,In_2158);
or U714 (N_714,In_2931,In_2800);
xnor U715 (N_715,In_981,In_1814);
xor U716 (N_716,In_2707,In_1182);
xor U717 (N_717,In_2665,In_2608);
nor U718 (N_718,In_671,In_1079);
and U719 (N_719,In_2928,In_911);
nor U720 (N_720,In_2131,In_1352);
nor U721 (N_721,In_2145,In_1920);
nand U722 (N_722,In_1346,In_42);
nand U723 (N_723,In_336,In_2463);
nand U724 (N_724,In_1747,In_1694);
and U725 (N_725,In_2024,In_2938);
or U726 (N_726,In_636,In_1369);
nand U727 (N_727,In_2756,In_2577);
nand U728 (N_728,In_756,In_1828);
nand U729 (N_729,In_1557,In_2548);
and U730 (N_730,In_1,In_1255);
and U731 (N_731,In_230,In_716);
xor U732 (N_732,In_2138,In_2108);
and U733 (N_733,In_194,In_812);
and U734 (N_734,In_135,In_2806);
nand U735 (N_735,In_2074,In_1084);
and U736 (N_736,In_2855,In_2632);
nand U737 (N_737,In_2523,In_1708);
nand U738 (N_738,In_404,In_2423);
or U739 (N_739,In_1797,In_2831);
nor U740 (N_740,In_1238,In_2747);
or U741 (N_741,In_2262,In_2709);
nor U742 (N_742,In_1536,In_1596);
xor U743 (N_743,In_1443,In_411);
and U744 (N_744,In_2813,In_2282);
or U745 (N_745,In_2743,In_1606);
nand U746 (N_746,In_1642,In_2890);
nand U747 (N_747,In_2077,In_2843);
or U748 (N_748,In_2578,In_360);
xnor U749 (N_749,In_722,In_218);
and U750 (N_750,In_2148,In_902);
xnor U751 (N_751,In_1756,In_1160);
xor U752 (N_752,In_2270,In_2459);
xor U753 (N_753,In_538,In_1893);
xnor U754 (N_754,In_941,In_397);
nand U755 (N_755,In_372,In_1187);
and U756 (N_756,In_973,In_1570);
or U757 (N_757,In_2521,In_624);
and U758 (N_758,In_831,In_2537);
xnor U759 (N_759,In_414,In_2593);
nor U760 (N_760,In_2942,In_1019);
or U761 (N_761,In_266,In_1758);
and U762 (N_762,In_2731,In_1892);
and U763 (N_763,In_276,In_472);
xnor U764 (N_764,In_1672,In_2000);
nand U765 (N_765,In_1745,In_245);
or U766 (N_766,In_1535,In_1524);
and U767 (N_767,In_1106,In_693);
or U768 (N_768,In_2976,In_1192);
or U769 (N_769,In_1087,In_946);
nand U770 (N_770,In_2378,In_2277);
xnor U771 (N_771,In_2474,In_2205);
and U772 (N_772,In_1936,In_686);
or U773 (N_773,In_1965,In_742);
nand U774 (N_774,In_1751,In_2648);
nand U775 (N_775,In_2055,In_1716);
nand U776 (N_776,In_164,In_893);
nor U777 (N_777,In_1341,In_2793);
nor U778 (N_778,In_1505,In_1386);
or U779 (N_779,In_2686,In_2214);
nand U780 (N_780,In_541,In_1795);
nand U781 (N_781,In_2850,In_2988);
xor U782 (N_782,In_763,In_2767);
nor U783 (N_783,In_2434,In_834);
xor U784 (N_784,In_2421,In_1476);
nor U785 (N_785,In_1349,In_2769);
xor U786 (N_786,In_1401,In_2545);
nor U787 (N_787,In_2028,In_2161);
and U788 (N_788,In_1085,In_1523);
or U789 (N_789,In_461,In_936);
nand U790 (N_790,In_2812,In_2237);
nand U791 (N_791,In_972,In_2937);
nand U792 (N_792,In_359,In_109);
xor U793 (N_793,In_486,In_1303);
and U794 (N_794,In_465,In_2210);
xor U795 (N_795,In_1759,In_17);
nand U796 (N_796,In_119,In_1247);
or U797 (N_797,In_1552,In_1620);
nand U798 (N_798,In_2981,In_2592);
or U799 (N_799,In_2245,In_963);
nor U800 (N_800,In_20,In_767);
xnor U801 (N_801,In_2984,In_1704);
or U802 (N_802,In_545,In_627);
nand U803 (N_803,In_1064,In_113);
and U804 (N_804,In_1676,In_1116);
xor U805 (N_805,In_27,In_2009);
or U806 (N_806,In_2422,In_484);
nand U807 (N_807,In_1768,In_2397);
or U808 (N_808,In_2304,In_2107);
nor U809 (N_809,In_1315,In_562);
xor U810 (N_810,In_2944,In_1953);
and U811 (N_811,In_100,In_2452);
or U812 (N_812,In_434,In_2168);
nand U813 (N_813,In_888,In_2123);
nand U814 (N_814,In_2171,In_2018);
nand U815 (N_815,In_2913,In_1300);
xor U816 (N_816,In_2840,In_1650);
nor U817 (N_817,In_1102,In_1705);
and U818 (N_818,In_2978,In_2451);
xnor U819 (N_819,In_1938,In_1648);
xnor U820 (N_820,In_579,In_2289);
nor U821 (N_821,In_1518,In_2320);
or U822 (N_822,In_1188,In_1279);
and U823 (N_823,In_433,In_714);
or U824 (N_824,In_1260,In_1109);
and U825 (N_825,In_180,In_2189);
and U826 (N_826,In_2676,In_1891);
and U827 (N_827,In_794,In_1158);
or U828 (N_828,In_885,In_1697);
nand U829 (N_829,In_2035,In_698);
nor U830 (N_830,In_790,In_1438);
and U831 (N_831,In_1482,In_1103);
and U832 (N_832,In_2430,In_1132);
or U833 (N_833,In_1712,In_2960);
xnor U834 (N_834,In_2568,In_2062);
and U835 (N_835,In_150,In_1080);
nand U836 (N_836,In_772,In_1440);
xor U837 (N_837,In_1389,In_1485);
or U838 (N_838,In_1478,In_308);
nand U839 (N_839,In_1971,In_1631);
or U840 (N_840,In_1862,In_765);
xnor U841 (N_841,In_1836,In_2048);
or U842 (N_842,In_449,In_1168);
xor U843 (N_843,In_1851,In_1005);
or U844 (N_844,In_1483,In_616);
nor U845 (N_845,In_2367,In_2737);
and U846 (N_846,In_1903,In_94);
and U847 (N_847,In_2991,In_2987);
or U848 (N_848,In_1811,In_92);
and U849 (N_849,In_227,In_1680);
or U850 (N_850,In_1053,In_413);
or U851 (N_851,In_1391,In_74);
and U852 (N_852,In_542,In_2531);
nand U853 (N_853,In_498,In_224);
xnor U854 (N_854,In_1198,In_2173);
xnor U855 (N_855,In_808,In_2871);
nand U856 (N_856,In_602,In_256);
nand U857 (N_857,In_2719,In_2685);
or U858 (N_858,In_1029,In_889);
nand U859 (N_859,In_710,In_2615);
xnor U860 (N_860,In_576,In_1380);
xnor U861 (N_861,In_2789,In_1193);
nand U862 (N_862,In_73,In_1226);
or U863 (N_863,In_895,In_1755);
and U864 (N_864,In_1414,In_1630);
nor U865 (N_865,In_795,In_1818);
xnor U866 (N_866,In_2045,In_655);
or U867 (N_867,In_324,In_664);
and U868 (N_868,In_72,In_1591);
or U869 (N_869,In_355,In_1996);
or U870 (N_870,In_45,In_942);
nor U871 (N_871,In_2154,In_2918);
or U872 (N_872,In_1161,In_2295);
or U873 (N_873,In_1637,In_1036);
nand U874 (N_874,In_2175,In_534);
nor U875 (N_875,In_2622,In_1024);
nand U876 (N_876,In_2962,In_2435);
nand U877 (N_877,In_1379,In_2049);
or U878 (N_878,In_2126,In_2975);
and U879 (N_879,In_1766,In_702);
xnor U880 (N_880,In_338,In_1376);
xor U881 (N_881,In_931,In_1398);
nand U882 (N_882,In_98,In_2655);
xnor U883 (N_883,In_2934,In_1267);
and U884 (N_884,In_2233,In_983);
nor U885 (N_885,In_198,In_666);
nand U886 (N_886,In_1813,In_451);
and U887 (N_887,In_1207,In_1202);
nor U888 (N_888,In_1281,In_9);
or U889 (N_889,In_2410,In_687);
nand U890 (N_890,In_1155,In_2757);
xnor U891 (N_891,In_2097,In_1744);
xnor U892 (N_892,In_2340,In_2560);
and U893 (N_893,In_1149,In_567);
nor U894 (N_894,In_26,In_2362);
or U895 (N_895,In_507,In_1131);
xor U896 (N_896,In_568,In_442);
nand U897 (N_897,In_739,In_2197);
or U898 (N_898,In_1550,In_253);
or U899 (N_899,In_1473,In_877);
xnor U900 (N_900,In_346,In_2823);
nor U901 (N_901,In_1527,In_2333);
xnor U902 (N_902,In_2220,In_2);
or U903 (N_903,In_1752,In_2260);
xor U904 (N_904,In_1643,In_1304);
nand U905 (N_905,In_352,In_2510);
xnor U906 (N_906,In_694,In_758);
nor U907 (N_907,In_2830,In_841);
xnor U908 (N_908,In_2388,In_420);
or U909 (N_909,In_1496,In_723);
or U910 (N_910,In_1779,In_593);
or U911 (N_911,In_1831,In_82);
and U912 (N_912,In_2357,In_958);
and U913 (N_913,In_2301,In_923);
nand U914 (N_914,In_2959,In_1317);
nand U915 (N_915,In_1826,In_311);
nand U916 (N_916,In_1299,In_2955);
nand U917 (N_917,In_2187,In_275);
or U918 (N_918,In_2654,In_2259);
or U919 (N_919,In_2708,In_1793);
nor U920 (N_920,In_2634,In_2172);
nor U921 (N_921,In_1351,In_5);
xor U922 (N_922,In_1141,In_325);
and U923 (N_923,In_548,In_859);
nor U924 (N_924,In_285,In_1037);
or U925 (N_925,In_1598,In_645);
nor U926 (N_926,In_2710,In_2336);
nand U927 (N_927,In_2179,In_2364);
xnor U928 (N_928,In_2412,In_1822);
nor U929 (N_929,In_2221,In_803);
or U930 (N_930,In_2472,In_1673);
or U931 (N_931,In_500,In_665);
nand U932 (N_932,In_1540,In_2642);
or U933 (N_933,In_2407,In_976);
nor U934 (N_934,In_549,In_1679);
and U935 (N_935,In_1320,In_990);
xor U936 (N_936,In_307,In_1787);
and U937 (N_937,In_1318,In_1337);
nand U938 (N_938,In_2588,In_1834);
nor U939 (N_939,In_1728,In_1678);
and U940 (N_940,In_1129,In_2971);
nor U941 (N_941,In_2223,In_1273);
and U942 (N_942,In_1521,In_1063);
xnor U943 (N_943,In_2275,In_520);
and U944 (N_944,In_706,In_1731);
nor U945 (N_945,In_1699,In_966);
and U946 (N_946,In_745,In_304);
or U947 (N_947,In_284,In_2712);
xor U948 (N_948,In_487,In_2222);
nand U949 (N_949,In_124,In_1803);
nor U950 (N_950,In_2759,In_2059);
nand U951 (N_951,In_2202,In_1487);
or U952 (N_952,In_1622,In_1590);
nor U953 (N_953,In_2735,In_886);
and U954 (N_954,In_1336,In_1494);
xor U955 (N_955,In_2701,In_2925);
nor U956 (N_956,In_1932,In_479);
and U957 (N_957,In_2564,In_165);
and U958 (N_958,In_1709,In_2574);
nand U959 (N_959,In_674,In_361);
xor U960 (N_960,In_1717,In_1167);
nor U961 (N_961,In_491,In_968);
nor U962 (N_962,In_2442,In_1272);
or U963 (N_963,In_2337,In_641);
nor U964 (N_964,In_1701,In_2659);
xnor U965 (N_965,In_1323,In_1083);
nand U966 (N_966,In_1775,In_1477);
nor U967 (N_967,In_2403,In_1044);
xnor U968 (N_968,In_185,In_630);
and U969 (N_969,In_2989,In_920);
nand U970 (N_970,In_319,In_2780);
xor U971 (N_971,In_1065,In_290);
nor U972 (N_972,In_1404,In_2808);
and U973 (N_973,In_1852,In_441);
nor U974 (N_974,In_1986,In_2089);
or U975 (N_975,In_777,In_1052);
or U976 (N_976,In_2749,In_648);
and U977 (N_977,In_351,In_1077);
xnor U978 (N_978,In_1419,In_2666);
nor U979 (N_979,In_2291,In_2303);
or U980 (N_980,In_2348,In_2527);
xnor U981 (N_981,In_417,In_2825);
xnor U982 (N_982,In_466,In_2504);
or U983 (N_983,In_1236,In_2414);
nor U984 (N_984,In_2954,In_570);
or U985 (N_985,In_332,In_2456);
or U986 (N_986,In_954,In_2864);
xnor U987 (N_987,In_934,In_2647);
nor U988 (N_988,In_900,In_725);
or U989 (N_989,In_1761,In_1729);
and U990 (N_990,In_1357,In_543);
nand U991 (N_991,In_388,In_1854);
nand U992 (N_992,In_2990,In_2917);
or U993 (N_993,In_950,In_232);
nor U994 (N_994,In_46,In_1689);
nor U995 (N_995,In_2099,In_370);
nor U996 (N_996,In_445,In_1781);
nor U997 (N_997,In_1760,In_572);
and U998 (N_998,In_619,In_887);
and U999 (N_999,In_460,In_18);
or U1000 (N_1000,In_647,In_403);
or U1001 (N_1001,In_2725,In_504);
nand U1002 (N_1002,In_2278,In_1784);
nor U1003 (N_1003,In_2013,In_1546);
xnor U1004 (N_1004,In_1301,In_1714);
and U1005 (N_1005,In_1663,In_1587);
nor U1006 (N_1006,In_1576,In_2092);
nor U1007 (N_1007,In_382,In_294);
and U1008 (N_1008,In_317,In_2607);
nor U1009 (N_1009,In_2409,In_1486);
or U1010 (N_1010,In_1951,In_1104);
or U1011 (N_1011,In_1604,In_1940);
and U1012 (N_1012,In_0,In_517);
xnor U1013 (N_1013,In_23,In_105);
and U1014 (N_1014,In_2445,In_471);
or U1015 (N_1015,In_720,In_2327);
xor U1016 (N_1016,In_344,In_943);
or U1017 (N_1017,In_2690,In_589);
and U1018 (N_1018,In_1724,In_2061);
nor U1019 (N_1019,In_2116,In_1148);
nand U1020 (N_1020,In_1809,In_2881);
nand U1021 (N_1021,In_1928,In_2667);
and U1022 (N_1022,In_481,In_891);
nand U1023 (N_1023,In_1295,In_2121);
xor U1024 (N_1024,In_1765,In_1229);
and U1025 (N_1025,In_1100,In_815);
nand U1026 (N_1026,In_2904,In_864);
or U1027 (N_1027,In_2476,In_670);
xor U1028 (N_1028,In_2985,In_350);
nor U1029 (N_1029,In_1070,In_184);
nor U1030 (N_1030,In_1789,In_412);
xor U1031 (N_1031,In_2253,In_267);
xnor U1032 (N_1032,In_1560,In_2957);
or U1033 (N_1033,In_1027,In_880);
and U1034 (N_1034,In_868,In_39);
or U1035 (N_1035,In_2312,In_127);
and U1036 (N_1036,In_1837,In_2164);
nor U1037 (N_1037,In_2149,In_1396);
xnor U1038 (N_1038,In_1902,In_1976);
nor U1039 (N_1039,In_571,In_145);
or U1040 (N_1040,In_335,In_2015);
or U1041 (N_1041,In_1776,In_1343);
nand U1042 (N_1042,In_1153,In_1011);
xor U1043 (N_1043,In_2207,In_30);
nor U1044 (N_1044,In_377,In_120);
xor U1045 (N_1045,In_533,In_755);
or U1046 (N_1046,In_948,In_1664);
nand U1047 (N_1047,In_2151,In_2859);
and U1048 (N_1048,In_2008,In_1548);
or U1049 (N_1049,In_588,In_1649);
nand U1050 (N_1050,In_2856,In_2628);
nor U1051 (N_1051,In_1194,In_945);
xor U1052 (N_1052,In_870,In_932);
and U1053 (N_1053,In_364,In_2639);
xnor U1054 (N_1054,In_1687,In_1442);
nor U1055 (N_1055,In_1804,In_1388);
and U1056 (N_1056,In_1258,In_2672);
or U1057 (N_1057,In_735,In_863);
xnor U1058 (N_1058,In_1842,In_590);
and U1059 (N_1059,In_1170,In_1884);
nand U1060 (N_1060,In_1553,In_2181);
nor U1061 (N_1061,In_2644,In_1371);
and U1062 (N_1062,In_544,In_1373);
or U1063 (N_1063,In_1868,In_577);
nor U1064 (N_1064,In_197,In_343);
nor U1065 (N_1065,In_1785,In_1983);
xnor U1066 (N_1066,In_719,In_2025);
nor U1067 (N_1067,In_597,In_2951);
nor U1068 (N_1068,In_2246,In_879);
nor U1069 (N_1069,In_644,In_673);
and U1070 (N_1070,In_2621,In_1707);
or U1071 (N_1071,In_2415,In_2211);
xor U1072 (N_1072,In_2760,In_1962);
and U1073 (N_1073,In_1313,In_1124);
nand U1074 (N_1074,In_675,In_1774);
nor U1075 (N_1075,In_2268,In_2612);
xor U1076 (N_1076,In_2794,In_157);
xnor U1077 (N_1077,In_273,In_2834);
and U1078 (N_1078,In_2946,In_1923);
xor U1079 (N_1079,In_375,In_2876);
or U1080 (N_1080,In_2084,In_586);
nor U1081 (N_1081,In_2318,In_1883);
nor U1082 (N_1082,In_2462,In_155);
xor U1083 (N_1083,In_2212,In_1375);
nor U1084 (N_1084,In_1034,In_1059);
or U1085 (N_1085,In_2618,In_357);
xnor U1086 (N_1086,In_2669,In_2678);
and U1087 (N_1087,In_749,In_2244);
nor U1088 (N_1088,In_1947,In_2815);
or U1089 (N_1089,In_56,In_2779);
and U1090 (N_1090,In_2542,In_1578);
nor U1091 (N_1091,In_50,In_1232);
xor U1092 (N_1092,In_805,In_1850);
nand U1093 (N_1093,In_354,In_1397);
nand U1094 (N_1094,In_1061,In_1602);
nor U1095 (N_1095,In_2069,In_632);
or U1096 (N_1096,In_2810,In_77);
nor U1097 (N_1097,In_1479,In_2129);
or U1098 (N_1098,In_525,In_1305);
nand U1099 (N_1099,In_726,In_1564);
nand U1100 (N_1100,In_1039,In_418);
xor U1101 (N_1101,In_2562,In_2273);
nor U1102 (N_1102,In_1668,In_1277);
or U1103 (N_1103,In_707,In_2674);
nor U1104 (N_1104,In_1381,In_1595);
nand U1105 (N_1105,In_1492,In_103);
nand U1106 (N_1106,In_766,In_555);
and U1107 (N_1107,In_1117,In_560);
xnor U1108 (N_1108,In_771,In_2979);
xor U1109 (N_1109,In_1017,In_1172);
nand U1110 (N_1110,In_1992,In_511);
and U1111 (N_1111,In_1402,In_2208);
nand U1112 (N_1112,In_1684,In_1231);
and U1113 (N_1113,In_181,In_658);
xnor U1114 (N_1114,In_1817,In_2063);
or U1115 (N_1115,In_86,In_1964);
xor U1116 (N_1116,In_2956,In_214);
nor U1117 (N_1117,In_1927,In_2656);
xnor U1118 (N_1118,In_1491,In_2924);
and U1119 (N_1119,In_953,In_2683);
xnor U1120 (N_1120,In_2071,In_2064);
nor U1121 (N_1121,In_530,In_299);
xnor U1122 (N_1122,In_473,In_1150);
nand U1123 (N_1123,In_709,In_175);
and U1124 (N_1124,In_1698,In_747);
nor U1125 (N_1125,In_2133,In_2909);
nand U1126 (N_1126,In_1211,In_2057);
nor U1127 (N_1127,In_1251,In_919);
xnor U1128 (N_1128,In_2418,In_2851);
xor U1129 (N_1129,In_475,In_1646);
and U1130 (N_1130,In_563,In_1464);
nor U1131 (N_1131,In_2331,In_884);
and U1132 (N_1132,In_2016,In_2571);
nand U1133 (N_1133,In_2439,In_247);
nand U1134 (N_1134,In_2923,In_804);
or U1135 (N_1135,In_2225,In_1635);
nor U1136 (N_1136,In_447,In_1224);
or U1137 (N_1137,In_1500,In_978);
xor U1138 (N_1138,In_974,In_980);
and U1139 (N_1139,In_248,In_2624);
nor U1140 (N_1140,In_1764,In_242);
or U1141 (N_1141,In_2468,In_439);
nor U1142 (N_1142,In_1754,In_241);
xnor U1143 (N_1143,In_2679,In_2020);
and U1144 (N_1144,In_2272,In_1257);
xor U1145 (N_1145,In_2324,In_2822);
nand U1146 (N_1146,In_430,In_1012);
nor U1147 (N_1147,In_915,In_603);
or U1148 (N_1148,In_2945,In_566);
and U1149 (N_1149,In_2170,In_1921);
or U1150 (N_1150,In_1031,In_1220);
xnor U1151 (N_1151,In_2251,In_391);
nand U1152 (N_1152,In_1894,In_1653);
xor U1153 (N_1153,In_2258,In_1530);
xnor U1154 (N_1154,In_2680,In_604);
and U1155 (N_1155,In_668,In_708);
nand U1156 (N_1156,In_1120,In_2724);
nor U1157 (N_1157,In_2109,In_1488);
nor U1158 (N_1158,In_1183,In_2585);
xnor U1159 (N_1159,In_262,In_1749);
or U1160 (N_1160,In_940,In_1048);
nor U1161 (N_1161,In_1133,In_2882);
nor U1162 (N_1162,In_1567,In_1467);
nand U1163 (N_1163,In_789,In_1177);
nand U1164 (N_1164,In_2366,In_2372);
xnor U1165 (N_1165,In_1020,In_2717);
or U1166 (N_1166,In_684,In_85);
and U1167 (N_1167,In_2058,In_2155);
nand U1168 (N_1168,In_1219,In_331);
nor U1169 (N_1169,In_933,In_2941);
nor U1170 (N_1170,In_2101,In_1583);
and U1171 (N_1171,In_2550,In_2786);
and U1172 (N_1172,In_574,In_1859);
and U1173 (N_1173,In_1554,In_206);
xor U1174 (N_1174,In_1154,In_1144);
xnor U1175 (N_1175,In_171,In_1802);
or U1176 (N_1176,In_492,In_239);
or U1177 (N_1177,In_1960,In_2520);
or U1178 (N_1178,In_1018,In_408);
or U1179 (N_1179,In_2044,In_2467);
or U1180 (N_1180,In_2664,In_929);
and U1181 (N_1181,In_883,In_1201);
nor U1182 (N_1182,In_2495,In_1042);
and U1183 (N_1183,In_1506,In_599);
and U1184 (N_1184,In_2837,In_2514);
nand U1185 (N_1185,In_827,In_1203);
or U1186 (N_1186,In_2182,In_1312);
xor U1187 (N_1187,In_2752,In_365);
nand U1188 (N_1188,In_2781,In_2450);
and U1189 (N_1189,In_183,In_2723);
and U1190 (N_1190,In_1878,In_1905);
nand U1191 (N_1191,In_287,In_1599);
or U1192 (N_1192,In_1600,In_1497);
and U1193 (N_1193,In_605,In_1670);
or U1194 (N_1194,In_1040,In_924);
nand U1195 (N_1195,In_2635,In_2702);
nand U1196 (N_1196,In_2824,In_824);
or U1197 (N_1197,In_1191,In_2771);
nor U1198 (N_1198,In_2216,In_2997);
and U1199 (N_1199,In_2949,In_527);
and U1200 (N_1200,In_836,In_2764);
nand U1201 (N_1201,In_142,In_318);
or U1202 (N_1202,In_167,In_1214);
or U1203 (N_1203,In_1974,In_1853);
and U1204 (N_1204,In_2488,In_2046);
and U1205 (N_1205,In_2281,In_1110);
nor U1206 (N_1206,In_1778,In_1189);
xnor U1207 (N_1207,In_866,In_2081);
and U1208 (N_1208,In_2460,In_2479);
nor U1209 (N_1209,In_1210,In_501);
or U1210 (N_1210,In_187,In_2021);
nand U1211 (N_1211,In_2466,In_2266);
or U1212 (N_1212,In_2727,In_2626);
nor U1213 (N_1213,In_2167,In_1801);
nor U1214 (N_1214,In_1522,In_2746);
nand U1215 (N_1215,In_2065,In_2853);
nor U1216 (N_1216,In_732,In_2558);
xor U1217 (N_1217,In_407,In_2711);
nor U1218 (N_1218,In_718,In_89);
xor U1219 (N_1219,In_1786,In_2032);
or U1220 (N_1220,In_1502,In_592);
xor U1221 (N_1221,In_2503,In_2513);
and U1222 (N_1222,In_2426,In_66);
and U1223 (N_1223,In_1783,In_2007);
or U1224 (N_1224,In_2590,In_2603);
xnor U1225 (N_1225,In_539,In_1173);
nor U1226 (N_1226,In_6,In_1001);
nor U1227 (N_1227,In_246,In_1792);
nand U1228 (N_1228,In_2299,In_869);
xor U1229 (N_1229,In_1134,In_1618);
nor U1230 (N_1230,In_1259,In_1989);
and U1231 (N_1231,In_2042,In_2325);
and U1232 (N_1232,In_2963,In_1584);
nor U1233 (N_1233,In_2902,In_736);
or U1234 (N_1234,In_813,In_614);
nor U1235 (N_1235,In_1991,In_306);
and U1236 (N_1236,In_1864,In_1274);
nand U1237 (N_1237,In_2502,In_705);
nor U1238 (N_1238,In_106,In_2517);
xor U1239 (N_1239,In_1455,In_2425);
and U1240 (N_1240,In_2417,In_132);
xor U1241 (N_1241,In_2897,In_1904);
or U1242 (N_1242,In_1742,In_1750);
nor U1243 (N_1243,In_231,In_1105);
or U1244 (N_1244,In_1421,In_78);
nand U1245 (N_1245,In_1949,In_2370);
xnor U1246 (N_1246,In_1686,In_1253);
or U1247 (N_1247,In_2477,In_1732);
or U1248 (N_1248,In_2721,In_1338);
nor U1249 (N_1249,In_1695,In_2267);
nand U1250 (N_1250,In_2870,In_182);
and U1251 (N_1251,In_7,In_2613);
xor U1252 (N_1252,In_2751,In_818);
xnor U1253 (N_1253,In_2306,In_807);
xnor U1254 (N_1254,In_1403,In_298);
xor U1255 (N_1255,In_540,In_1757);
xor U1256 (N_1256,In_216,In_110);
and U1257 (N_1257,In_598,In_2034);
xor U1258 (N_1258,In_2528,In_2401);
xor U1259 (N_1259,In_2798,In_2424);
and U1260 (N_1260,In_1919,In_345);
nor U1261 (N_1261,In_697,In_2493);
or U1262 (N_1262,In_1125,In_1901);
nor U1263 (N_1263,In_1925,In_1875);
nand U1264 (N_1264,In_446,In_2250);
or U1265 (N_1265,In_1594,In_221);
xnor U1266 (N_1266,In_1186,In_13);
or U1267 (N_1267,In_156,In_740);
nor U1268 (N_1268,In_556,In_1378);
or U1269 (N_1269,In_2023,In_729);
and U1270 (N_1270,In_2374,In_1308);
nor U1271 (N_1271,In_1221,In_200);
nand U1272 (N_1272,In_1909,In_1212);
or U1273 (N_1273,In_2285,In_453);
xnor U1274 (N_1274,In_2693,In_1244);
or U1275 (N_1275,In_2958,In_2054);
and U1276 (N_1276,In_2860,In_1405);
or U1277 (N_1277,In_1693,In_2804);
nor U1278 (N_1278,In_1888,In_2554);
nor U1279 (N_1279,In_384,In_2689);
nand U1280 (N_1280,In_58,In_810);
or U1281 (N_1281,In_2605,In_1233);
or U1282 (N_1282,In_2485,In_2763);
or U1283 (N_1283,In_312,In_153);
nor U1284 (N_1284,In_1603,In_1016);
or U1285 (N_1285,In_405,In_1970);
xnor U1286 (N_1286,In_371,In_2038);
or U1287 (N_1287,In_1942,In_1720);
xnor U1288 (N_1288,In_1924,In_1096);
nor U1289 (N_1289,In_1999,In_1880);
xnor U1290 (N_1290,In_1430,In_2083);
nand U1291 (N_1291,In_1355,In_279);
xnor U1292 (N_1292,In_1367,In_1470);
nor U1293 (N_1293,In_623,In_1329);
nor U1294 (N_1294,In_41,In_1715);
or U1295 (N_1295,In_2716,In_2829);
or U1296 (N_1296,In_1028,In_1762);
xnor U1297 (N_1297,In_781,In_1093);
nor U1298 (N_1298,In_2113,In_69);
nor U1299 (N_1299,In_1748,In_2100);
nand U1300 (N_1300,In_1055,In_608);
nand U1301 (N_1301,In_2386,In_547);
nor U1302 (N_1302,In_1472,In_1423);
or U1303 (N_1303,In_1135,In_2135);
nor U1304 (N_1304,In_2929,In_2072);
nor U1305 (N_1305,In_1335,In_1512);
nor U1306 (N_1306,In_2631,In_2455);
nand U1307 (N_1307,In_144,In_2443);
nand U1308 (N_1308,In_327,In_947);
and U1309 (N_1309,In_1108,In_2883);
and U1310 (N_1310,In_2816,In_2629);
nor U1311 (N_1311,In_2358,In_1411);
nor U1312 (N_1312,In_1000,In_2346);
nand U1313 (N_1313,In_383,In_443);
xor U1314 (N_1314,In_1738,In_581);
or U1315 (N_1315,In_653,In_2248);
xor U1316 (N_1316,In_2001,In_1140);
nor U1317 (N_1317,In_1796,In_594);
nor U1318 (N_1318,In_314,In_2419);
xor U1319 (N_1319,In_1533,In_209);
xor U1320 (N_1320,In_1647,In_977);
nand U1321 (N_1321,In_44,In_158);
nor U1322 (N_1322,In_2950,In_925);
or U1323 (N_1323,In_1638,In_2872);
xor U1324 (N_1324,In_1264,In_762);
nor U1325 (N_1325,In_986,In_251);
and U1326 (N_1326,In_1867,In_1215);
nand U1327 (N_1327,In_690,In_358);
and U1328 (N_1328,In_1032,In_856);
nor U1329 (N_1329,In_2569,In_2649);
or U1330 (N_1330,In_1078,In_300);
xor U1331 (N_1331,In_2313,In_170);
and U1332 (N_1332,In_1617,In_330);
nor U1333 (N_1333,In_663,In_1772);
xnor U1334 (N_1334,In_141,In_1146);
or U1335 (N_1335,In_2993,In_743);
or U1336 (N_1336,In_2239,In_1408);
xnor U1337 (N_1337,In_2836,In_654);
nand U1338 (N_1338,In_514,In_1286);
or U1339 (N_1339,In_2127,In_1568);
or U1340 (N_1340,In_2797,In_1624);
xor U1341 (N_1341,In_2785,In_1086);
and U1342 (N_1342,In_1394,In_1081);
or U1343 (N_1343,In_2232,In_927);
or U1344 (N_1344,In_1823,In_1725);
or U1345 (N_1345,In_1468,In_2473);
nand U1346 (N_1346,In_509,In_2224);
nor U1347 (N_1347,In_2491,In_2231);
xor U1348 (N_1348,In_270,In_47);
and U1349 (N_1349,In_849,In_512);
nand U1350 (N_1350,In_506,In_1098);
and U1351 (N_1351,In_905,In_843);
or U1352 (N_1352,In_2826,In_2242);
and U1353 (N_1353,In_2887,In_2287);
nand U1354 (N_1354,In_904,In_1159);
nor U1355 (N_1355,In_1980,In_2349);
and U1356 (N_1356,In_660,In_621);
or U1357 (N_1357,In_764,In_2296);
and U1358 (N_1358,In_1794,In_1046);
xnor U1359 (N_1359,In_1250,In_2651);
and U1360 (N_1360,In_1666,In_1979);
and U1361 (N_1361,In_1348,In_618);
and U1362 (N_1362,In_2703,In_2633);
nand U1363 (N_1363,In_133,In_926);
nand U1364 (N_1364,In_1364,In_1573);
xor U1365 (N_1365,In_1370,In_1449);
nor U1366 (N_1366,In_1126,In_380);
nor U1367 (N_1367,In_261,In_2518);
nor U1368 (N_1368,In_2807,In_949);
nand U1369 (N_1369,In_208,In_681);
and U1370 (N_1370,In_907,In_1306);
xnor U1371 (N_1371,In_845,In_595);
nand U1372 (N_1372,In_606,In_1361);
xor U1373 (N_1373,In_734,In_985);
xor U1374 (N_1374,In_2144,In_470);
nor U1375 (N_1375,In_228,In_2961);
or U1376 (N_1376,In_416,In_2376);
xor U1377 (N_1377,In_721,In_2575);
nand U1378 (N_1378,In_2274,In_497);
and U1379 (N_1379,In_1805,In_2885);
nor U1380 (N_1380,In_2778,In_2453);
xnor U1381 (N_1381,In_1930,In_421);
and U1382 (N_1382,In_457,In_1111);
and U1383 (N_1383,In_1929,In_2379);
nor U1384 (N_1384,In_2117,In_871);
xor U1385 (N_1385,In_536,In_1896);
nand U1386 (N_1386,In_1311,In_524);
nor U1387 (N_1387,In_118,In_1041);
nand U1388 (N_1388,In_278,In_1659);
or U1389 (N_1389,In_2106,In_2662);
nor U1390 (N_1390,In_1071,In_450);
nand U1391 (N_1391,In_2697,In_179);
xor U1392 (N_1392,In_2730,In_1395);
xor U1393 (N_1393,In_1278,In_1917);
and U1394 (N_1394,In_190,In_51);
and U1395 (N_1395,In_2601,In_2857);
or U1396 (N_1396,In_2294,In_2865);
or U1397 (N_1397,In_1551,In_2873);
and U1398 (N_1398,In_1955,In_2360);
nand U1399 (N_1399,In_2480,In_490);
xor U1400 (N_1400,In_1356,In_75);
or U1401 (N_1401,In_1767,In_368);
or U1402 (N_1402,In_468,In_2734);
or U1403 (N_1403,In_2627,In_1677);
and U1404 (N_1404,In_711,In_857);
or U1405 (N_1405,In_761,In_2323);
nand U1406 (N_1406,In_1372,In_363);
and U1407 (N_1407,In_2892,In_2602);
xnor U1408 (N_1408,In_2682,In_320);
xnor U1409 (N_1409,In_2302,In_678);
nand U1410 (N_1410,In_440,In_2102);
xnor U1411 (N_1411,In_395,In_426);
xor U1412 (N_1412,In_508,In_1777);
nand U1413 (N_1413,In_1985,In_2893);
nor U1414 (N_1414,In_111,In_1130);
nor U1415 (N_1415,In_2140,In_1871);
or U1416 (N_1416,In_2315,In_1216);
or U1417 (N_1417,In_1439,In_95);
nor U1418 (N_1418,In_1906,In_1015);
nand U1419 (N_1419,In_928,In_1114);
nand U1420 (N_1420,In_1569,In_2777);
xnor U1421 (N_1421,In_81,In_2053);
or U1422 (N_1422,In_2566,In_1156);
xor U1423 (N_1423,In_385,In_1292);
or U1424 (N_1424,In_1503,In_63);
or U1425 (N_1425,In_1393,In_1143);
nor U1426 (N_1426,In_1091,In_1702);
and U1427 (N_1427,In_970,In_1632);
nand U1428 (N_1428,In_1122,In_321);
or U1429 (N_1429,In_1254,In_235);
and U1430 (N_1430,In_1066,In_908);
nand U1431 (N_1431,In_2056,In_1515);
nand U1432 (N_1432,In_651,In_992);
or U1433 (N_1433,In_1266,In_601);
xor U1434 (N_1434,In_587,In_1660);
nand U1435 (N_1435,In_1072,In_1948);
nand U1436 (N_1436,In_1035,In_583);
or U1437 (N_1437,In_2983,In_1413);
xor U1438 (N_1438,In_2515,In_203);
or U1439 (N_1439,In_2668,In_32);
and U1440 (N_1440,In_2754,In_493);
nand U1441 (N_1441,In_2279,In_2073);
and U1442 (N_1442,In_2845,In_1245);
and U1443 (N_1443,In_1544,In_2500);
nor U1444 (N_1444,In_1223,In_1099);
or U1445 (N_1445,In_2458,In_1950);
and U1446 (N_1446,In_12,In_2005);
and U1447 (N_1447,In_2874,In_861);
nand U1448 (N_1448,In_177,In_2903);
or U1449 (N_1449,In_2646,In_22);
xor U1450 (N_1450,In_2219,In_2970);
nor U1451 (N_1451,In_2163,In_1899);
xnor U1452 (N_1452,In_2849,In_2901);
or U1453 (N_1453,In_2448,In_286);
nor U1454 (N_1454,In_2594,In_982);
nor U1455 (N_1455,In_40,In_49);
xnor U1456 (N_1456,In_2803,In_2898);
and U1457 (N_1457,In_2838,In_832);
and U1458 (N_1458,In_1885,In_1827);
and U1459 (N_1459,In_1577,In_422);
and U1460 (N_1460,In_2694,In_2136);
and U1461 (N_1461,In_523,In_1023);
and U1462 (N_1462,In_2186,In_854);
xor U1463 (N_1463,In_2761,In_432);
and U1464 (N_1464,In_837,In_1848);
xor U1465 (N_1465,In_169,In_564);
nand U1466 (N_1466,In_438,In_1572);
xor U1467 (N_1467,In_2586,In_2854);
nor U1468 (N_1468,In_489,In_840);
nand U1469 (N_1469,In_2103,In_1988);
nand U1470 (N_1470,In_2203,In_2093);
xnor U1471 (N_1471,In_1995,In_2411);
and U1472 (N_1472,In_1665,In_822);
xnor U1473 (N_1473,In_1026,In_515);
nor U1474 (N_1474,In_1199,In_1614);
nand U1475 (N_1475,In_292,In_2589);
or U1476 (N_1476,In_2653,In_24);
nor U1477 (N_1477,In_2408,In_478);
xor U1478 (N_1478,In_8,In_1359);
nand U1479 (N_1479,In_876,In_2783);
or U1480 (N_1480,In_839,In_2110);
nand U1481 (N_1481,In_825,In_35);
xor U1482 (N_1482,In_984,In_1340);
nor U1483 (N_1483,In_1799,In_700);
and U1484 (N_1484,In_1592,In_989);
and U1485 (N_1485,In_381,In_826);
nand U1486 (N_1486,In_1288,In_2494);
nand U1487 (N_1487,In_1152,In_573);
and U1488 (N_1488,In_917,In_2795);
and U1489 (N_1489,In_1121,In_1743);
nand U1490 (N_1490,In_600,In_2228);
and U1491 (N_1491,In_2249,In_956);
and U1492 (N_1492,In_768,In_1941);
xor U1493 (N_1493,In_1654,In_1271);
and U1494 (N_1494,In_995,In_521);
and U1495 (N_1495,In_1441,In_1209);
nor U1496 (N_1496,In_1118,In_2240);
nand U1497 (N_1497,In_386,In_860);
or U1498 (N_1498,In_1558,In_160);
nor U1499 (N_1499,In_1113,In_1115);
and U1500 (N_1500,In_2401,In_580);
or U1501 (N_1501,In_435,In_2334);
nand U1502 (N_1502,In_2007,In_460);
nor U1503 (N_1503,In_83,In_1218);
nor U1504 (N_1504,In_2878,In_374);
xnor U1505 (N_1505,In_759,In_1991);
and U1506 (N_1506,In_2228,In_2607);
or U1507 (N_1507,In_2667,In_1717);
xor U1508 (N_1508,In_1176,In_1109);
nor U1509 (N_1509,In_2022,In_1516);
xor U1510 (N_1510,In_296,In_1973);
or U1511 (N_1511,In_2907,In_2015);
or U1512 (N_1512,In_260,In_168);
nand U1513 (N_1513,In_2873,In_2514);
and U1514 (N_1514,In_260,In_2926);
nor U1515 (N_1515,In_2577,In_728);
nand U1516 (N_1516,In_2084,In_2310);
nor U1517 (N_1517,In_1620,In_2814);
nor U1518 (N_1518,In_2970,In_1088);
or U1519 (N_1519,In_772,In_1554);
nand U1520 (N_1520,In_1729,In_662);
nand U1521 (N_1521,In_1691,In_1593);
nand U1522 (N_1522,In_2241,In_2612);
and U1523 (N_1523,In_825,In_1301);
xor U1524 (N_1524,In_2108,In_472);
xnor U1525 (N_1525,In_2638,In_36);
nor U1526 (N_1526,In_581,In_2124);
nor U1527 (N_1527,In_537,In_2078);
xor U1528 (N_1528,In_564,In_1276);
xnor U1529 (N_1529,In_2579,In_2542);
xor U1530 (N_1530,In_2522,In_468);
nand U1531 (N_1531,In_2551,In_557);
and U1532 (N_1532,In_2980,In_2669);
nand U1533 (N_1533,In_2363,In_2287);
xor U1534 (N_1534,In_2861,In_2075);
nand U1535 (N_1535,In_856,In_2619);
nor U1536 (N_1536,In_1218,In_1497);
nor U1537 (N_1537,In_1425,In_1966);
xor U1538 (N_1538,In_2787,In_946);
nand U1539 (N_1539,In_2361,In_2648);
or U1540 (N_1540,In_2209,In_1645);
or U1541 (N_1541,In_829,In_2677);
xnor U1542 (N_1542,In_2369,In_1026);
nand U1543 (N_1543,In_643,In_2952);
or U1544 (N_1544,In_1454,In_2618);
nand U1545 (N_1545,In_246,In_1225);
nand U1546 (N_1546,In_885,In_2990);
or U1547 (N_1547,In_565,In_542);
nand U1548 (N_1548,In_1386,In_1978);
or U1549 (N_1549,In_203,In_1716);
and U1550 (N_1550,In_2316,In_768);
or U1551 (N_1551,In_1078,In_259);
xnor U1552 (N_1552,In_891,In_101);
or U1553 (N_1553,In_2128,In_46);
nor U1554 (N_1554,In_2156,In_2492);
xor U1555 (N_1555,In_449,In_2405);
xor U1556 (N_1556,In_1306,In_258);
or U1557 (N_1557,In_1987,In_2889);
nor U1558 (N_1558,In_2994,In_1726);
nor U1559 (N_1559,In_1596,In_545);
nand U1560 (N_1560,In_377,In_2669);
xor U1561 (N_1561,In_1040,In_1405);
xor U1562 (N_1562,In_2400,In_1282);
xor U1563 (N_1563,In_732,In_1291);
nand U1564 (N_1564,In_632,In_2202);
or U1565 (N_1565,In_2957,In_1116);
and U1566 (N_1566,In_495,In_266);
nor U1567 (N_1567,In_913,In_302);
or U1568 (N_1568,In_491,In_2217);
or U1569 (N_1569,In_951,In_2137);
nand U1570 (N_1570,In_1674,In_1002);
nor U1571 (N_1571,In_2568,In_984);
and U1572 (N_1572,In_577,In_2971);
or U1573 (N_1573,In_2159,In_2203);
nand U1574 (N_1574,In_478,In_757);
xor U1575 (N_1575,In_2283,In_982);
xor U1576 (N_1576,In_477,In_1416);
xnor U1577 (N_1577,In_16,In_682);
xnor U1578 (N_1578,In_2176,In_627);
and U1579 (N_1579,In_2144,In_1409);
xnor U1580 (N_1580,In_987,In_504);
xnor U1581 (N_1581,In_2910,In_1415);
nand U1582 (N_1582,In_2103,In_104);
xnor U1583 (N_1583,In_811,In_1580);
nand U1584 (N_1584,In_739,In_2680);
nand U1585 (N_1585,In_2618,In_1911);
nor U1586 (N_1586,In_2540,In_527);
nor U1587 (N_1587,In_2966,In_23);
nor U1588 (N_1588,In_2982,In_1129);
and U1589 (N_1589,In_260,In_2239);
nand U1590 (N_1590,In_847,In_182);
xor U1591 (N_1591,In_275,In_215);
nor U1592 (N_1592,In_1611,In_763);
nand U1593 (N_1593,In_632,In_1960);
or U1594 (N_1594,In_554,In_2837);
nand U1595 (N_1595,In_1876,In_1953);
nor U1596 (N_1596,In_1426,In_1041);
and U1597 (N_1597,In_66,In_2874);
xor U1598 (N_1598,In_372,In_2167);
and U1599 (N_1599,In_78,In_1128);
and U1600 (N_1600,In_374,In_919);
nor U1601 (N_1601,In_2099,In_1792);
nor U1602 (N_1602,In_2417,In_2876);
or U1603 (N_1603,In_2680,In_1293);
and U1604 (N_1604,In_2089,In_1488);
and U1605 (N_1605,In_344,In_1358);
or U1606 (N_1606,In_2140,In_2774);
nand U1607 (N_1607,In_1076,In_380);
and U1608 (N_1608,In_2216,In_1410);
or U1609 (N_1609,In_2911,In_2637);
nand U1610 (N_1610,In_1280,In_2600);
nand U1611 (N_1611,In_2846,In_1623);
or U1612 (N_1612,In_1640,In_771);
nor U1613 (N_1613,In_855,In_380);
or U1614 (N_1614,In_1190,In_126);
xnor U1615 (N_1615,In_1415,In_688);
nor U1616 (N_1616,In_1367,In_342);
or U1617 (N_1617,In_1798,In_2958);
or U1618 (N_1618,In_2968,In_880);
or U1619 (N_1619,In_2734,In_2984);
or U1620 (N_1620,In_812,In_686);
or U1621 (N_1621,In_431,In_1779);
nor U1622 (N_1622,In_2688,In_462);
or U1623 (N_1623,In_1944,In_1347);
or U1624 (N_1624,In_1574,In_2796);
nor U1625 (N_1625,In_1860,In_784);
xnor U1626 (N_1626,In_1932,In_2733);
nand U1627 (N_1627,In_203,In_2828);
nor U1628 (N_1628,In_1605,In_1600);
and U1629 (N_1629,In_2790,In_917);
nor U1630 (N_1630,In_1122,In_1653);
and U1631 (N_1631,In_1642,In_1261);
nand U1632 (N_1632,In_1153,In_1583);
or U1633 (N_1633,In_1321,In_1081);
nor U1634 (N_1634,In_2970,In_2271);
nand U1635 (N_1635,In_1438,In_2996);
nand U1636 (N_1636,In_1802,In_1857);
or U1637 (N_1637,In_2564,In_2186);
and U1638 (N_1638,In_1205,In_890);
xor U1639 (N_1639,In_2914,In_971);
or U1640 (N_1640,In_982,In_828);
nor U1641 (N_1641,In_2310,In_984);
nand U1642 (N_1642,In_554,In_2671);
nand U1643 (N_1643,In_2373,In_2867);
nor U1644 (N_1644,In_115,In_2189);
nor U1645 (N_1645,In_1024,In_272);
xor U1646 (N_1646,In_2057,In_1386);
nand U1647 (N_1647,In_1420,In_2365);
or U1648 (N_1648,In_2615,In_1076);
and U1649 (N_1649,In_917,In_2214);
xnor U1650 (N_1650,In_1992,In_1347);
xor U1651 (N_1651,In_2428,In_2808);
xnor U1652 (N_1652,In_1883,In_1638);
or U1653 (N_1653,In_940,In_1978);
xor U1654 (N_1654,In_847,In_750);
nor U1655 (N_1655,In_2108,In_528);
nand U1656 (N_1656,In_1521,In_1613);
nand U1657 (N_1657,In_1081,In_2528);
nand U1658 (N_1658,In_573,In_1151);
xor U1659 (N_1659,In_771,In_893);
xnor U1660 (N_1660,In_93,In_2826);
nor U1661 (N_1661,In_139,In_845);
and U1662 (N_1662,In_979,In_1664);
nand U1663 (N_1663,In_2226,In_2602);
or U1664 (N_1664,In_786,In_2613);
xor U1665 (N_1665,In_1522,In_1374);
and U1666 (N_1666,In_2168,In_2464);
nand U1667 (N_1667,In_2207,In_1846);
nor U1668 (N_1668,In_1829,In_469);
or U1669 (N_1669,In_286,In_2230);
xnor U1670 (N_1670,In_1211,In_1304);
and U1671 (N_1671,In_877,In_2259);
or U1672 (N_1672,In_567,In_90);
nor U1673 (N_1673,In_303,In_618);
and U1674 (N_1674,In_1201,In_660);
nand U1675 (N_1675,In_1236,In_301);
nor U1676 (N_1676,In_2507,In_2519);
and U1677 (N_1677,In_969,In_1853);
nand U1678 (N_1678,In_1634,In_1889);
or U1679 (N_1679,In_589,In_2646);
nand U1680 (N_1680,In_1294,In_392);
nor U1681 (N_1681,In_669,In_310);
and U1682 (N_1682,In_2551,In_348);
xnor U1683 (N_1683,In_897,In_1862);
xor U1684 (N_1684,In_2718,In_540);
or U1685 (N_1685,In_1498,In_2766);
nand U1686 (N_1686,In_984,In_1611);
nor U1687 (N_1687,In_1159,In_602);
xnor U1688 (N_1688,In_1451,In_2245);
nor U1689 (N_1689,In_1200,In_1317);
or U1690 (N_1690,In_1204,In_2365);
xnor U1691 (N_1691,In_2269,In_1705);
and U1692 (N_1692,In_1993,In_442);
xor U1693 (N_1693,In_13,In_1724);
or U1694 (N_1694,In_679,In_2264);
nor U1695 (N_1695,In_1422,In_455);
nor U1696 (N_1696,In_2640,In_1054);
nor U1697 (N_1697,In_1730,In_2247);
or U1698 (N_1698,In_1145,In_1126);
nor U1699 (N_1699,In_1573,In_633);
nand U1700 (N_1700,In_773,In_540);
nand U1701 (N_1701,In_1893,In_608);
nor U1702 (N_1702,In_2847,In_2669);
nor U1703 (N_1703,In_2947,In_178);
and U1704 (N_1704,In_44,In_1571);
nand U1705 (N_1705,In_2856,In_2108);
nor U1706 (N_1706,In_2949,In_1026);
and U1707 (N_1707,In_792,In_842);
nor U1708 (N_1708,In_233,In_2077);
xor U1709 (N_1709,In_1201,In_1408);
nand U1710 (N_1710,In_1989,In_2626);
and U1711 (N_1711,In_2384,In_1849);
xnor U1712 (N_1712,In_1447,In_1755);
xnor U1713 (N_1713,In_1599,In_182);
and U1714 (N_1714,In_2716,In_400);
xnor U1715 (N_1715,In_2499,In_2564);
xor U1716 (N_1716,In_2301,In_2253);
and U1717 (N_1717,In_772,In_411);
nand U1718 (N_1718,In_348,In_385);
nor U1719 (N_1719,In_2758,In_2823);
nor U1720 (N_1720,In_1471,In_1745);
xnor U1721 (N_1721,In_1048,In_2224);
xor U1722 (N_1722,In_1388,In_924);
xnor U1723 (N_1723,In_2125,In_1473);
nor U1724 (N_1724,In_1473,In_460);
nor U1725 (N_1725,In_2734,In_2588);
or U1726 (N_1726,In_2610,In_2125);
or U1727 (N_1727,In_2225,In_930);
nor U1728 (N_1728,In_1530,In_1533);
xor U1729 (N_1729,In_1009,In_1002);
or U1730 (N_1730,In_938,In_1116);
or U1731 (N_1731,In_2810,In_2520);
nand U1732 (N_1732,In_435,In_2259);
xnor U1733 (N_1733,In_983,In_212);
and U1734 (N_1734,In_1162,In_2471);
xor U1735 (N_1735,In_2727,In_1600);
xor U1736 (N_1736,In_174,In_2605);
nor U1737 (N_1737,In_2728,In_1386);
or U1738 (N_1738,In_458,In_2898);
and U1739 (N_1739,In_2018,In_823);
and U1740 (N_1740,In_1875,In_1967);
nand U1741 (N_1741,In_2568,In_1685);
xor U1742 (N_1742,In_336,In_980);
xnor U1743 (N_1743,In_557,In_1738);
nor U1744 (N_1744,In_2637,In_281);
or U1745 (N_1745,In_840,In_366);
xor U1746 (N_1746,In_2216,In_2952);
xnor U1747 (N_1747,In_562,In_1246);
nor U1748 (N_1748,In_1200,In_773);
and U1749 (N_1749,In_897,In_1225);
nand U1750 (N_1750,In_6,In_1548);
xnor U1751 (N_1751,In_1051,In_160);
nor U1752 (N_1752,In_1020,In_2523);
xor U1753 (N_1753,In_944,In_2840);
xnor U1754 (N_1754,In_1753,In_2969);
or U1755 (N_1755,In_2746,In_1817);
or U1756 (N_1756,In_1750,In_2742);
and U1757 (N_1757,In_425,In_372);
and U1758 (N_1758,In_754,In_1329);
nand U1759 (N_1759,In_365,In_2908);
nor U1760 (N_1760,In_967,In_1817);
and U1761 (N_1761,In_2557,In_505);
xnor U1762 (N_1762,In_589,In_1139);
and U1763 (N_1763,In_670,In_1574);
and U1764 (N_1764,In_752,In_2177);
xnor U1765 (N_1765,In_2747,In_687);
and U1766 (N_1766,In_2121,In_1660);
nand U1767 (N_1767,In_1828,In_1490);
and U1768 (N_1768,In_916,In_1108);
nand U1769 (N_1769,In_1440,In_323);
and U1770 (N_1770,In_1383,In_2325);
or U1771 (N_1771,In_150,In_1486);
or U1772 (N_1772,In_2024,In_1248);
nor U1773 (N_1773,In_2263,In_1860);
nand U1774 (N_1774,In_2731,In_1247);
xnor U1775 (N_1775,In_623,In_2556);
xor U1776 (N_1776,In_2778,In_650);
nand U1777 (N_1777,In_2872,In_2195);
and U1778 (N_1778,In_1409,In_2161);
nand U1779 (N_1779,In_2820,In_2623);
or U1780 (N_1780,In_1754,In_696);
nor U1781 (N_1781,In_209,In_1725);
nand U1782 (N_1782,In_294,In_1316);
or U1783 (N_1783,In_574,In_1625);
or U1784 (N_1784,In_2506,In_609);
xor U1785 (N_1785,In_1808,In_1955);
xnor U1786 (N_1786,In_2072,In_1744);
and U1787 (N_1787,In_1822,In_1937);
or U1788 (N_1788,In_1328,In_1996);
nor U1789 (N_1789,In_567,In_2177);
nand U1790 (N_1790,In_448,In_531);
nand U1791 (N_1791,In_329,In_535);
nand U1792 (N_1792,In_2119,In_552);
or U1793 (N_1793,In_521,In_1361);
xnor U1794 (N_1794,In_2741,In_169);
xnor U1795 (N_1795,In_423,In_2355);
xnor U1796 (N_1796,In_2783,In_8);
or U1797 (N_1797,In_1435,In_2021);
nand U1798 (N_1798,In_2076,In_2376);
nor U1799 (N_1799,In_2443,In_2863);
and U1800 (N_1800,In_2016,In_34);
and U1801 (N_1801,In_171,In_2563);
nor U1802 (N_1802,In_576,In_251);
or U1803 (N_1803,In_1359,In_374);
xnor U1804 (N_1804,In_77,In_1489);
and U1805 (N_1805,In_1627,In_2121);
or U1806 (N_1806,In_1689,In_627);
nand U1807 (N_1807,In_2673,In_948);
xnor U1808 (N_1808,In_1644,In_2451);
nor U1809 (N_1809,In_1974,In_1198);
nor U1810 (N_1810,In_1656,In_2907);
xnor U1811 (N_1811,In_1363,In_1791);
or U1812 (N_1812,In_2284,In_1851);
or U1813 (N_1813,In_636,In_2437);
nor U1814 (N_1814,In_319,In_2896);
xnor U1815 (N_1815,In_956,In_2894);
or U1816 (N_1816,In_1008,In_1099);
and U1817 (N_1817,In_2011,In_1779);
and U1818 (N_1818,In_171,In_206);
nand U1819 (N_1819,In_2144,In_2058);
and U1820 (N_1820,In_409,In_574);
xnor U1821 (N_1821,In_673,In_1275);
nor U1822 (N_1822,In_2057,In_1354);
nor U1823 (N_1823,In_2256,In_1647);
nand U1824 (N_1824,In_998,In_1790);
and U1825 (N_1825,In_1807,In_2940);
nand U1826 (N_1826,In_993,In_1190);
and U1827 (N_1827,In_995,In_515);
and U1828 (N_1828,In_1,In_156);
and U1829 (N_1829,In_1973,In_1263);
or U1830 (N_1830,In_857,In_1186);
nor U1831 (N_1831,In_1302,In_1598);
xnor U1832 (N_1832,In_2506,In_1344);
xnor U1833 (N_1833,In_1478,In_418);
nor U1834 (N_1834,In_677,In_1810);
and U1835 (N_1835,In_1728,In_2218);
xnor U1836 (N_1836,In_1514,In_558);
or U1837 (N_1837,In_1435,In_1581);
xnor U1838 (N_1838,In_2528,In_1606);
and U1839 (N_1839,In_2999,In_2632);
nand U1840 (N_1840,In_881,In_60);
xor U1841 (N_1841,In_1622,In_2215);
xor U1842 (N_1842,In_860,In_2113);
or U1843 (N_1843,In_2085,In_1107);
nand U1844 (N_1844,In_772,In_911);
xor U1845 (N_1845,In_1193,In_603);
or U1846 (N_1846,In_449,In_272);
xnor U1847 (N_1847,In_1496,In_1272);
nor U1848 (N_1848,In_376,In_1805);
or U1849 (N_1849,In_972,In_739);
nand U1850 (N_1850,In_1228,In_586);
xor U1851 (N_1851,In_372,In_2045);
nor U1852 (N_1852,In_180,In_1600);
nor U1853 (N_1853,In_712,In_2201);
and U1854 (N_1854,In_1254,In_1818);
xnor U1855 (N_1855,In_1034,In_536);
or U1856 (N_1856,In_2585,In_1096);
or U1857 (N_1857,In_1372,In_770);
nor U1858 (N_1858,In_2630,In_1284);
nor U1859 (N_1859,In_703,In_2118);
nand U1860 (N_1860,In_1023,In_2641);
xnor U1861 (N_1861,In_2522,In_1213);
nor U1862 (N_1862,In_1889,In_2497);
or U1863 (N_1863,In_1025,In_2293);
nand U1864 (N_1864,In_1965,In_537);
xor U1865 (N_1865,In_1769,In_1882);
and U1866 (N_1866,In_1643,In_464);
nand U1867 (N_1867,In_58,In_2133);
xnor U1868 (N_1868,In_623,In_332);
nand U1869 (N_1869,In_2227,In_382);
or U1870 (N_1870,In_38,In_2134);
nor U1871 (N_1871,In_1359,In_2619);
and U1872 (N_1872,In_806,In_2877);
nor U1873 (N_1873,In_261,In_286);
and U1874 (N_1874,In_1691,In_1033);
and U1875 (N_1875,In_1347,In_1257);
nand U1876 (N_1876,In_150,In_2878);
nor U1877 (N_1877,In_1681,In_2958);
nor U1878 (N_1878,In_1552,In_186);
nor U1879 (N_1879,In_428,In_482);
nand U1880 (N_1880,In_1101,In_2388);
nor U1881 (N_1881,In_549,In_977);
and U1882 (N_1882,In_2366,In_1154);
or U1883 (N_1883,In_2481,In_846);
and U1884 (N_1884,In_732,In_2585);
xnor U1885 (N_1885,In_1014,In_558);
and U1886 (N_1886,In_2231,In_1913);
nor U1887 (N_1887,In_1148,In_296);
nor U1888 (N_1888,In_175,In_2733);
nand U1889 (N_1889,In_84,In_815);
and U1890 (N_1890,In_2376,In_449);
and U1891 (N_1891,In_2052,In_625);
or U1892 (N_1892,In_2590,In_2618);
xnor U1893 (N_1893,In_1426,In_2199);
and U1894 (N_1894,In_2528,In_1232);
xor U1895 (N_1895,In_162,In_1414);
nand U1896 (N_1896,In_1519,In_555);
nor U1897 (N_1897,In_560,In_923);
nor U1898 (N_1898,In_332,In_119);
nand U1899 (N_1899,In_195,In_2938);
or U1900 (N_1900,In_2165,In_893);
nor U1901 (N_1901,In_633,In_390);
nor U1902 (N_1902,In_464,In_156);
nor U1903 (N_1903,In_2601,In_720);
xnor U1904 (N_1904,In_1312,In_747);
xnor U1905 (N_1905,In_403,In_1169);
and U1906 (N_1906,In_709,In_749);
and U1907 (N_1907,In_2429,In_1716);
nor U1908 (N_1908,In_1092,In_242);
nand U1909 (N_1909,In_402,In_1521);
nor U1910 (N_1910,In_855,In_619);
and U1911 (N_1911,In_412,In_709);
nand U1912 (N_1912,In_1559,In_878);
and U1913 (N_1913,In_775,In_2428);
nor U1914 (N_1914,In_2689,In_2666);
nand U1915 (N_1915,In_1768,In_2704);
nor U1916 (N_1916,In_685,In_547);
or U1917 (N_1917,In_2805,In_2210);
or U1918 (N_1918,In_426,In_213);
or U1919 (N_1919,In_2360,In_2825);
nor U1920 (N_1920,In_1261,In_374);
nand U1921 (N_1921,In_1571,In_2554);
nor U1922 (N_1922,In_2929,In_1865);
and U1923 (N_1923,In_2478,In_2706);
nand U1924 (N_1924,In_628,In_1680);
xor U1925 (N_1925,In_2692,In_1747);
or U1926 (N_1926,In_2385,In_423);
or U1927 (N_1927,In_484,In_1989);
xnor U1928 (N_1928,In_1104,In_396);
nand U1929 (N_1929,In_2410,In_2720);
and U1930 (N_1930,In_2791,In_730);
nor U1931 (N_1931,In_2781,In_1805);
or U1932 (N_1932,In_516,In_674);
nand U1933 (N_1933,In_2658,In_1599);
xor U1934 (N_1934,In_1068,In_1198);
and U1935 (N_1935,In_2350,In_212);
nor U1936 (N_1936,In_1318,In_179);
xnor U1937 (N_1937,In_2352,In_1085);
nand U1938 (N_1938,In_691,In_588);
and U1939 (N_1939,In_1005,In_2090);
xor U1940 (N_1940,In_203,In_1094);
nand U1941 (N_1941,In_257,In_2709);
nand U1942 (N_1942,In_2920,In_1038);
nor U1943 (N_1943,In_1287,In_2004);
nor U1944 (N_1944,In_1764,In_57);
nand U1945 (N_1945,In_2797,In_1675);
and U1946 (N_1946,In_1730,In_711);
nor U1947 (N_1947,In_965,In_2533);
nand U1948 (N_1948,In_2964,In_992);
nand U1949 (N_1949,In_2359,In_1981);
and U1950 (N_1950,In_380,In_1679);
and U1951 (N_1951,In_1954,In_990);
nand U1952 (N_1952,In_451,In_2838);
or U1953 (N_1953,In_2069,In_1104);
or U1954 (N_1954,In_2229,In_1194);
nand U1955 (N_1955,In_702,In_1571);
or U1956 (N_1956,In_2584,In_601);
and U1957 (N_1957,In_2170,In_406);
and U1958 (N_1958,In_176,In_368);
or U1959 (N_1959,In_2719,In_739);
nand U1960 (N_1960,In_2311,In_412);
nor U1961 (N_1961,In_1118,In_1266);
nor U1962 (N_1962,In_1634,In_2305);
and U1963 (N_1963,In_2421,In_2354);
nor U1964 (N_1964,In_809,In_1262);
nor U1965 (N_1965,In_2455,In_1257);
and U1966 (N_1966,In_96,In_42);
or U1967 (N_1967,In_1724,In_1848);
nand U1968 (N_1968,In_668,In_1276);
nor U1969 (N_1969,In_2130,In_192);
nand U1970 (N_1970,In_1620,In_1082);
and U1971 (N_1971,In_2201,In_922);
xor U1972 (N_1972,In_2486,In_2795);
nand U1973 (N_1973,In_292,In_2142);
or U1974 (N_1974,In_2349,In_1567);
nand U1975 (N_1975,In_1179,In_724);
xnor U1976 (N_1976,In_1402,In_894);
or U1977 (N_1977,In_2214,In_2579);
and U1978 (N_1978,In_214,In_2297);
nand U1979 (N_1979,In_1233,In_299);
nor U1980 (N_1980,In_1630,In_677);
and U1981 (N_1981,In_2586,In_2379);
nand U1982 (N_1982,In_2505,In_2188);
nand U1983 (N_1983,In_2128,In_2901);
nand U1984 (N_1984,In_2591,In_1938);
and U1985 (N_1985,In_434,In_187);
or U1986 (N_1986,In_2051,In_193);
and U1987 (N_1987,In_2029,In_33);
and U1988 (N_1988,In_2167,In_2277);
nand U1989 (N_1989,In_2685,In_200);
xor U1990 (N_1990,In_793,In_2787);
nand U1991 (N_1991,In_521,In_695);
nand U1992 (N_1992,In_2210,In_2547);
nor U1993 (N_1993,In_2534,In_1272);
nand U1994 (N_1994,In_1682,In_2725);
nor U1995 (N_1995,In_2473,In_2814);
and U1996 (N_1996,In_2831,In_954);
nand U1997 (N_1997,In_1798,In_1929);
and U1998 (N_1998,In_789,In_1864);
nor U1999 (N_1999,In_2719,In_351);
nor U2000 (N_2000,In_1457,In_2914);
nand U2001 (N_2001,In_1412,In_2990);
nand U2002 (N_2002,In_148,In_819);
nor U2003 (N_2003,In_2285,In_2082);
and U2004 (N_2004,In_2345,In_498);
or U2005 (N_2005,In_1875,In_937);
nand U2006 (N_2006,In_1915,In_1977);
xor U2007 (N_2007,In_360,In_2815);
nor U2008 (N_2008,In_1740,In_2707);
nor U2009 (N_2009,In_1867,In_1336);
nand U2010 (N_2010,In_1371,In_870);
nand U2011 (N_2011,In_2987,In_1539);
and U2012 (N_2012,In_65,In_1883);
and U2013 (N_2013,In_1760,In_2483);
nor U2014 (N_2014,In_2163,In_2948);
xnor U2015 (N_2015,In_1303,In_1720);
xor U2016 (N_2016,In_9,In_1062);
nor U2017 (N_2017,In_453,In_1433);
xor U2018 (N_2018,In_17,In_875);
nand U2019 (N_2019,In_1013,In_342);
or U2020 (N_2020,In_992,In_2157);
xor U2021 (N_2021,In_2973,In_806);
xnor U2022 (N_2022,In_2941,In_2201);
nor U2023 (N_2023,In_1673,In_2684);
nand U2024 (N_2024,In_2066,In_279);
nand U2025 (N_2025,In_1163,In_2564);
and U2026 (N_2026,In_1520,In_383);
or U2027 (N_2027,In_1663,In_932);
or U2028 (N_2028,In_2321,In_2422);
and U2029 (N_2029,In_1643,In_1712);
or U2030 (N_2030,In_2708,In_178);
and U2031 (N_2031,In_1356,In_1073);
or U2032 (N_2032,In_2840,In_2851);
nor U2033 (N_2033,In_1312,In_1929);
xor U2034 (N_2034,In_971,In_1009);
or U2035 (N_2035,In_957,In_1710);
nor U2036 (N_2036,In_2544,In_1236);
and U2037 (N_2037,In_1159,In_1268);
nor U2038 (N_2038,In_1181,In_2293);
xor U2039 (N_2039,In_1387,In_117);
xor U2040 (N_2040,In_494,In_564);
xnor U2041 (N_2041,In_263,In_329);
nand U2042 (N_2042,In_2782,In_895);
xnor U2043 (N_2043,In_741,In_311);
nand U2044 (N_2044,In_1465,In_1910);
xnor U2045 (N_2045,In_2317,In_1322);
and U2046 (N_2046,In_2801,In_1521);
nand U2047 (N_2047,In_113,In_75);
and U2048 (N_2048,In_2514,In_2513);
and U2049 (N_2049,In_1637,In_1942);
and U2050 (N_2050,In_2339,In_162);
nand U2051 (N_2051,In_72,In_1232);
nor U2052 (N_2052,In_1105,In_2912);
and U2053 (N_2053,In_785,In_1220);
nand U2054 (N_2054,In_2446,In_404);
xor U2055 (N_2055,In_2711,In_2815);
nand U2056 (N_2056,In_1629,In_2823);
or U2057 (N_2057,In_1952,In_1824);
xor U2058 (N_2058,In_2729,In_2833);
nand U2059 (N_2059,In_1643,In_2989);
nor U2060 (N_2060,In_618,In_241);
nand U2061 (N_2061,In_2231,In_1647);
or U2062 (N_2062,In_2179,In_597);
xor U2063 (N_2063,In_2436,In_267);
xor U2064 (N_2064,In_1746,In_2090);
or U2065 (N_2065,In_2684,In_2376);
nand U2066 (N_2066,In_490,In_2552);
xnor U2067 (N_2067,In_1892,In_2139);
or U2068 (N_2068,In_1147,In_126);
xnor U2069 (N_2069,In_1522,In_2988);
nand U2070 (N_2070,In_26,In_1451);
or U2071 (N_2071,In_1244,In_747);
nand U2072 (N_2072,In_2826,In_1602);
nand U2073 (N_2073,In_2080,In_1271);
and U2074 (N_2074,In_1599,In_1755);
xor U2075 (N_2075,In_2575,In_1619);
and U2076 (N_2076,In_1771,In_2744);
nor U2077 (N_2077,In_626,In_199);
nand U2078 (N_2078,In_2133,In_634);
and U2079 (N_2079,In_2260,In_137);
nor U2080 (N_2080,In_1610,In_1907);
and U2081 (N_2081,In_1328,In_1912);
or U2082 (N_2082,In_440,In_2992);
xor U2083 (N_2083,In_1454,In_146);
or U2084 (N_2084,In_995,In_2323);
xnor U2085 (N_2085,In_393,In_1415);
nor U2086 (N_2086,In_775,In_346);
xor U2087 (N_2087,In_1949,In_1041);
nor U2088 (N_2088,In_804,In_456);
xor U2089 (N_2089,In_715,In_1957);
or U2090 (N_2090,In_2281,In_2434);
and U2091 (N_2091,In_158,In_1008);
xor U2092 (N_2092,In_2461,In_582);
nor U2093 (N_2093,In_1735,In_2756);
nor U2094 (N_2094,In_2911,In_2223);
and U2095 (N_2095,In_308,In_2524);
xor U2096 (N_2096,In_2847,In_576);
nor U2097 (N_2097,In_1477,In_583);
nor U2098 (N_2098,In_290,In_1470);
nor U2099 (N_2099,In_1899,In_802);
and U2100 (N_2100,In_1546,In_1703);
xor U2101 (N_2101,In_2599,In_2659);
and U2102 (N_2102,In_2258,In_2662);
and U2103 (N_2103,In_210,In_2576);
nand U2104 (N_2104,In_1001,In_2045);
or U2105 (N_2105,In_609,In_2927);
and U2106 (N_2106,In_1304,In_1635);
nor U2107 (N_2107,In_2645,In_2738);
xnor U2108 (N_2108,In_1717,In_2757);
nor U2109 (N_2109,In_56,In_179);
nand U2110 (N_2110,In_482,In_2344);
or U2111 (N_2111,In_442,In_1328);
or U2112 (N_2112,In_2027,In_2660);
nor U2113 (N_2113,In_2439,In_2132);
and U2114 (N_2114,In_954,In_1431);
nand U2115 (N_2115,In_1310,In_1764);
and U2116 (N_2116,In_1041,In_94);
nor U2117 (N_2117,In_2253,In_2340);
or U2118 (N_2118,In_2761,In_132);
xnor U2119 (N_2119,In_2676,In_2186);
nand U2120 (N_2120,In_731,In_1039);
or U2121 (N_2121,In_1748,In_1896);
or U2122 (N_2122,In_685,In_268);
nand U2123 (N_2123,In_1519,In_149);
and U2124 (N_2124,In_2806,In_693);
nor U2125 (N_2125,In_1817,In_2723);
or U2126 (N_2126,In_382,In_1731);
nand U2127 (N_2127,In_862,In_2726);
xnor U2128 (N_2128,In_320,In_2843);
xor U2129 (N_2129,In_1985,In_1242);
xnor U2130 (N_2130,In_22,In_2126);
or U2131 (N_2131,In_1364,In_314);
or U2132 (N_2132,In_2330,In_1576);
and U2133 (N_2133,In_2207,In_2151);
and U2134 (N_2134,In_2024,In_2049);
nand U2135 (N_2135,In_672,In_173);
nor U2136 (N_2136,In_89,In_1039);
and U2137 (N_2137,In_2842,In_2846);
xor U2138 (N_2138,In_1012,In_2009);
and U2139 (N_2139,In_694,In_992);
nand U2140 (N_2140,In_2708,In_393);
xor U2141 (N_2141,In_1889,In_933);
or U2142 (N_2142,In_1266,In_1553);
or U2143 (N_2143,In_1469,In_2218);
xnor U2144 (N_2144,In_205,In_2497);
nand U2145 (N_2145,In_1175,In_1607);
xor U2146 (N_2146,In_1870,In_932);
nor U2147 (N_2147,In_1407,In_1362);
or U2148 (N_2148,In_1975,In_2738);
or U2149 (N_2149,In_530,In_1165);
nand U2150 (N_2150,In_21,In_596);
or U2151 (N_2151,In_1036,In_2306);
and U2152 (N_2152,In_2740,In_1216);
and U2153 (N_2153,In_410,In_357);
xor U2154 (N_2154,In_698,In_1474);
or U2155 (N_2155,In_286,In_963);
nor U2156 (N_2156,In_2745,In_1235);
xnor U2157 (N_2157,In_2326,In_1498);
and U2158 (N_2158,In_1292,In_2232);
nand U2159 (N_2159,In_1940,In_1244);
nor U2160 (N_2160,In_2777,In_398);
and U2161 (N_2161,In_449,In_1813);
and U2162 (N_2162,In_2016,In_48);
nand U2163 (N_2163,In_251,In_2126);
or U2164 (N_2164,In_2198,In_194);
or U2165 (N_2165,In_136,In_663);
nor U2166 (N_2166,In_2514,In_1319);
xnor U2167 (N_2167,In_268,In_2116);
or U2168 (N_2168,In_2968,In_2043);
or U2169 (N_2169,In_1947,In_2295);
or U2170 (N_2170,In_2743,In_576);
xor U2171 (N_2171,In_2284,In_1530);
xnor U2172 (N_2172,In_2723,In_2936);
nand U2173 (N_2173,In_2533,In_553);
xnor U2174 (N_2174,In_365,In_2125);
or U2175 (N_2175,In_185,In_1545);
nor U2176 (N_2176,In_1063,In_2568);
or U2177 (N_2177,In_461,In_621);
and U2178 (N_2178,In_188,In_117);
xor U2179 (N_2179,In_1780,In_856);
nor U2180 (N_2180,In_1,In_1738);
nand U2181 (N_2181,In_208,In_2198);
nand U2182 (N_2182,In_470,In_2216);
or U2183 (N_2183,In_2361,In_112);
nand U2184 (N_2184,In_617,In_77);
xnor U2185 (N_2185,In_1013,In_1903);
nand U2186 (N_2186,In_447,In_2945);
nand U2187 (N_2187,In_1023,In_443);
xor U2188 (N_2188,In_2115,In_470);
nor U2189 (N_2189,In_1809,In_2653);
nand U2190 (N_2190,In_2785,In_887);
nand U2191 (N_2191,In_547,In_1860);
or U2192 (N_2192,In_800,In_2833);
or U2193 (N_2193,In_581,In_2396);
xnor U2194 (N_2194,In_2336,In_1528);
nand U2195 (N_2195,In_2990,In_2379);
nand U2196 (N_2196,In_2259,In_966);
nor U2197 (N_2197,In_2061,In_2630);
and U2198 (N_2198,In_1611,In_596);
xor U2199 (N_2199,In_386,In_494);
or U2200 (N_2200,In_603,In_617);
and U2201 (N_2201,In_65,In_736);
xnor U2202 (N_2202,In_2566,In_620);
xor U2203 (N_2203,In_775,In_1183);
and U2204 (N_2204,In_1877,In_915);
nor U2205 (N_2205,In_2018,In_1137);
xor U2206 (N_2206,In_196,In_2064);
or U2207 (N_2207,In_862,In_2824);
xnor U2208 (N_2208,In_1422,In_1536);
nor U2209 (N_2209,In_2134,In_674);
or U2210 (N_2210,In_2531,In_821);
xnor U2211 (N_2211,In_2839,In_262);
or U2212 (N_2212,In_1321,In_2548);
and U2213 (N_2213,In_2968,In_1677);
or U2214 (N_2214,In_901,In_1051);
xor U2215 (N_2215,In_184,In_1936);
nor U2216 (N_2216,In_1755,In_1062);
nor U2217 (N_2217,In_55,In_2262);
or U2218 (N_2218,In_1450,In_1700);
xor U2219 (N_2219,In_2145,In_633);
and U2220 (N_2220,In_451,In_2723);
or U2221 (N_2221,In_2875,In_2482);
nor U2222 (N_2222,In_2634,In_530);
xnor U2223 (N_2223,In_2591,In_1977);
nor U2224 (N_2224,In_1166,In_1203);
and U2225 (N_2225,In_2731,In_808);
nand U2226 (N_2226,In_2876,In_2155);
nor U2227 (N_2227,In_2772,In_2830);
xnor U2228 (N_2228,In_2502,In_1061);
or U2229 (N_2229,In_1067,In_1427);
nor U2230 (N_2230,In_1291,In_184);
nor U2231 (N_2231,In_1992,In_996);
nor U2232 (N_2232,In_1873,In_1621);
xnor U2233 (N_2233,In_2211,In_1083);
xor U2234 (N_2234,In_155,In_173);
xor U2235 (N_2235,In_392,In_1103);
nand U2236 (N_2236,In_2711,In_1014);
nand U2237 (N_2237,In_1818,In_395);
nand U2238 (N_2238,In_1347,In_1530);
and U2239 (N_2239,In_2314,In_1424);
nor U2240 (N_2240,In_400,In_2010);
nor U2241 (N_2241,In_258,In_2234);
nand U2242 (N_2242,In_1439,In_1793);
and U2243 (N_2243,In_127,In_1893);
nor U2244 (N_2244,In_1826,In_2486);
and U2245 (N_2245,In_2529,In_1023);
xor U2246 (N_2246,In_2969,In_2788);
nand U2247 (N_2247,In_1118,In_2603);
and U2248 (N_2248,In_67,In_454);
xnor U2249 (N_2249,In_2905,In_2867);
nand U2250 (N_2250,In_1004,In_673);
or U2251 (N_2251,In_2839,In_1550);
and U2252 (N_2252,In_2984,In_2019);
nand U2253 (N_2253,In_1403,In_301);
and U2254 (N_2254,In_320,In_2914);
or U2255 (N_2255,In_504,In_1333);
nor U2256 (N_2256,In_1307,In_348);
or U2257 (N_2257,In_1048,In_1215);
nand U2258 (N_2258,In_2592,In_769);
nand U2259 (N_2259,In_2505,In_1669);
xnor U2260 (N_2260,In_480,In_2302);
nand U2261 (N_2261,In_970,In_597);
nor U2262 (N_2262,In_2700,In_1713);
or U2263 (N_2263,In_1998,In_117);
xnor U2264 (N_2264,In_2412,In_2936);
nand U2265 (N_2265,In_1547,In_566);
and U2266 (N_2266,In_936,In_802);
xnor U2267 (N_2267,In_2772,In_1044);
and U2268 (N_2268,In_246,In_2235);
and U2269 (N_2269,In_1706,In_520);
nand U2270 (N_2270,In_488,In_2421);
nand U2271 (N_2271,In_2297,In_169);
nor U2272 (N_2272,In_2310,In_2490);
xor U2273 (N_2273,In_678,In_638);
and U2274 (N_2274,In_76,In_970);
xor U2275 (N_2275,In_1630,In_445);
nand U2276 (N_2276,In_1902,In_1047);
or U2277 (N_2277,In_2898,In_2310);
xnor U2278 (N_2278,In_2191,In_1417);
nor U2279 (N_2279,In_1087,In_1233);
and U2280 (N_2280,In_323,In_1808);
and U2281 (N_2281,In_2661,In_2419);
and U2282 (N_2282,In_1235,In_2367);
nor U2283 (N_2283,In_1214,In_2213);
or U2284 (N_2284,In_2277,In_1708);
or U2285 (N_2285,In_429,In_228);
or U2286 (N_2286,In_744,In_631);
and U2287 (N_2287,In_563,In_1821);
nor U2288 (N_2288,In_2840,In_2789);
nor U2289 (N_2289,In_111,In_2817);
or U2290 (N_2290,In_1264,In_729);
or U2291 (N_2291,In_699,In_1044);
nor U2292 (N_2292,In_474,In_2231);
nand U2293 (N_2293,In_342,In_1204);
and U2294 (N_2294,In_691,In_2197);
nor U2295 (N_2295,In_90,In_741);
and U2296 (N_2296,In_2420,In_673);
or U2297 (N_2297,In_1114,In_384);
or U2298 (N_2298,In_2171,In_1161);
or U2299 (N_2299,In_230,In_1090);
xnor U2300 (N_2300,In_2895,In_2282);
nor U2301 (N_2301,In_578,In_1951);
nor U2302 (N_2302,In_2864,In_499);
nor U2303 (N_2303,In_2367,In_1694);
nor U2304 (N_2304,In_1762,In_645);
and U2305 (N_2305,In_733,In_666);
nand U2306 (N_2306,In_1755,In_1958);
nand U2307 (N_2307,In_2205,In_216);
and U2308 (N_2308,In_1122,In_928);
nand U2309 (N_2309,In_734,In_2114);
nor U2310 (N_2310,In_780,In_2428);
or U2311 (N_2311,In_652,In_2475);
xnor U2312 (N_2312,In_806,In_2858);
xor U2313 (N_2313,In_2929,In_322);
nand U2314 (N_2314,In_2144,In_1766);
and U2315 (N_2315,In_2266,In_2243);
or U2316 (N_2316,In_995,In_1970);
nor U2317 (N_2317,In_2171,In_2295);
or U2318 (N_2318,In_57,In_2463);
nor U2319 (N_2319,In_2191,In_2583);
nand U2320 (N_2320,In_61,In_2847);
xnor U2321 (N_2321,In_267,In_2239);
or U2322 (N_2322,In_306,In_468);
or U2323 (N_2323,In_315,In_1626);
nand U2324 (N_2324,In_132,In_2931);
nand U2325 (N_2325,In_2093,In_2031);
or U2326 (N_2326,In_2851,In_2419);
or U2327 (N_2327,In_1638,In_599);
nor U2328 (N_2328,In_171,In_101);
xnor U2329 (N_2329,In_1855,In_2229);
xnor U2330 (N_2330,In_879,In_2488);
or U2331 (N_2331,In_1736,In_1360);
nor U2332 (N_2332,In_425,In_2828);
nand U2333 (N_2333,In_1528,In_530);
nor U2334 (N_2334,In_900,In_1702);
xor U2335 (N_2335,In_1248,In_465);
nor U2336 (N_2336,In_1835,In_1926);
nor U2337 (N_2337,In_1169,In_878);
nand U2338 (N_2338,In_1655,In_1988);
nor U2339 (N_2339,In_561,In_2576);
and U2340 (N_2340,In_647,In_2137);
and U2341 (N_2341,In_1708,In_1466);
nor U2342 (N_2342,In_1806,In_2924);
or U2343 (N_2343,In_671,In_794);
and U2344 (N_2344,In_1663,In_1810);
nor U2345 (N_2345,In_1773,In_1284);
and U2346 (N_2346,In_630,In_283);
or U2347 (N_2347,In_2536,In_2607);
or U2348 (N_2348,In_2648,In_2921);
nand U2349 (N_2349,In_875,In_359);
or U2350 (N_2350,In_1814,In_1231);
nand U2351 (N_2351,In_899,In_314);
nand U2352 (N_2352,In_646,In_1606);
nand U2353 (N_2353,In_2547,In_94);
nor U2354 (N_2354,In_1233,In_740);
and U2355 (N_2355,In_534,In_1840);
nand U2356 (N_2356,In_78,In_1687);
xor U2357 (N_2357,In_2167,In_427);
and U2358 (N_2358,In_2715,In_1343);
xnor U2359 (N_2359,In_796,In_2827);
xnor U2360 (N_2360,In_2584,In_2630);
nand U2361 (N_2361,In_2587,In_2930);
and U2362 (N_2362,In_2529,In_225);
and U2363 (N_2363,In_430,In_77);
and U2364 (N_2364,In_2631,In_1651);
and U2365 (N_2365,In_1008,In_2235);
nand U2366 (N_2366,In_926,In_2733);
and U2367 (N_2367,In_243,In_2204);
and U2368 (N_2368,In_2540,In_654);
xnor U2369 (N_2369,In_1442,In_1232);
nor U2370 (N_2370,In_753,In_1842);
nand U2371 (N_2371,In_2862,In_1742);
nor U2372 (N_2372,In_1179,In_2336);
nand U2373 (N_2373,In_2536,In_556);
nand U2374 (N_2374,In_2554,In_717);
or U2375 (N_2375,In_2692,In_1471);
or U2376 (N_2376,In_1029,In_196);
and U2377 (N_2377,In_2831,In_2386);
xnor U2378 (N_2378,In_611,In_2902);
nand U2379 (N_2379,In_2676,In_1209);
nor U2380 (N_2380,In_2981,In_1144);
or U2381 (N_2381,In_1918,In_2543);
nor U2382 (N_2382,In_2496,In_2026);
and U2383 (N_2383,In_2429,In_1324);
nor U2384 (N_2384,In_1784,In_2422);
and U2385 (N_2385,In_873,In_1881);
or U2386 (N_2386,In_1537,In_1130);
nor U2387 (N_2387,In_429,In_2258);
or U2388 (N_2388,In_103,In_264);
and U2389 (N_2389,In_795,In_2055);
nor U2390 (N_2390,In_1485,In_2442);
nand U2391 (N_2391,In_1296,In_385);
xor U2392 (N_2392,In_1001,In_2116);
xnor U2393 (N_2393,In_2032,In_2597);
xor U2394 (N_2394,In_764,In_2658);
nor U2395 (N_2395,In_478,In_712);
xnor U2396 (N_2396,In_472,In_867);
and U2397 (N_2397,In_1166,In_1576);
nor U2398 (N_2398,In_2078,In_787);
or U2399 (N_2399,In_1687,In_48);
xnor U2400 (N_2400,In_982,In_912);
and U2401 (N_2401,In_252,In_2829);
or U2402 (N_2402,In_1926,In_2161);
and U2403 (N_2403,In_2398,In_815);
nand U2404 (N_2404,In_1497,In_216);
and U2405 (N_2405,In_295,In_1149);
and U2406 (N_2406,In_476,In_1678);
or U2407 (N_2407,In_25,In_2685);
nand U2408 (N_2408,In_2374,In_6);
nor U2409 (N_2409,In_1231,In_1639);
xor U2410 (N_2410,In_655,In_1319);
xor U2411 (N_2411,In_2276,In_2211);
nor U2412 (N_2412,In_2412,In_225);
xnor U2413 (N_2413,In_833,In_977);
nand U2414 (N_2414,In_177,In_202);
and U2415 (N_2415,In_1098,In_1017);
and U2416 (N_2416,In_559,In_2325);
xor U2417 (N_2417,In_1649,In_1700);
nand U2418 (N_2418,In_2930,In_2837);
and U2419 (N_2419,In_684,In_929);
or U2420 (N_2420,In_2184,In_655);
xnor U2421 (N_2421,In_879,In_2623);
xor U2422 (N_2422,In_772,In_492);
and U2423 (N_2423,In_55,In_397);
and U2424 (N_2424,In_1038,In_2478);
nor U2425 (N_2425,In_358,In_2497);
xor U2426 (N_2426,In_1401,In_2553);
or U2427 (N_2427,In_2147,In_2349);
or U2428 (N_2428,In_806,In_941);
or U2429 (N_2429,In_1777,In_1687);
and U2430 (N_2430,In_2435,In_225);
or U2431 (N_2431,In_259,In_2536);
xor U2432 (N_2432,In_1178,In_596);
nand U2433 (N_2433,In_1709,In_2015);
nor U2434 (N_2434,In_731,In_2286);
nor U2435 (N_2435,In_1301,In_2272);
xor U2436 (N_2436,In_2958,In_2798);
nand U2437 (N_2437,In_2714,In_1075);
nor U2438 (N_2438,In_1375,In_1931);
or U2439 (N_2439,In_231,In_1172);
and U2440 (N_2440,In_2414,In_1159);
nand U2441 (N_2441,In_334,In_51);
nor U2442 (N_2442,In_1095,In_2833);
and U2443 (N_2443,In_2743,In_1259);
nand U2444 (N_2444,In_603,In_2619);
nor U2445 (N_2445,In_2477,In_2376);
and U2446 (N_2446,In_2665,In_1992);
xor U2447 (N_2447,In_1073,In_1925);
nand U2448 (N_2448,In_145,In_31);
and U2449 (N_2449,In_1381,In_2275);
or U2450 (N_2450,In_2891,In_775);
nand U2451 (N_2451,In_2327,In_2819);
nand U2452 (N_2452,In_106,In_1166);
and U2453 (N_2453,In_2685,In_2085);
and U2454 (N_2454,In_234,In_1184);
or U2455 (N_2455,In_1662,In_1184);
nand U2456 (N_2456,In_45,In_290);
and U2457 (N_2457,In_861,In_2689);
nand U2458 (N_2458,In_1433,In_2660);
and U2459 (N_2459,In_2418,In_1709);
nor U2460 (N_2460,In_1643,In_271);
nor U2461 (N_2461,In_1728,In_2073);
or U2462 (N_2462,In_1430,In_2641);
nand U2463 (N_2463,In_865,In_546);
nand U2464 (N_2464,In_232,In_278);
xor U2465 (N_2465,In_1285,In_2906);
xor U2466 (N_2466,In_2473,In_2624);
nor U2467 (N_2467,In_2366,In_1832);
or U2468 (N_2468,In_2562,In_2285);
nand U2469 (N_2469,In_1069,In_2138);
nor U2470 (N_2470,In_1193,In_2148);
nand U2471 (N_2471,In_1463,In_1174);
nand U2472 (N_2472,In_1979,In_2264);
and U2473 (N_2473,In_444,In_393);
nor U2474 (N_2474,In_1843,In_555);
xor U2475 (N_2475,In_2828,In_2110);
or U2476 (N_2476,In_449,In_2835);
or U2477 (N_2477,In_764,In_2491);
nand U2478 (N_2478,In_2463,In_682);
xor U2479 (N_2479,In_1878,In_2933);
nor U2480 (N_2480,In_2184,In_1348);
nor U2481 (N_2481,In_536,In_1549);
and U2482 (N_2482,In_142,In_2632);
nor U2483 (N_2483,In_2963,In_2169);
xnor U2484 (N_2484,In_223,In_1269);
nor U2485 (N_2485,In_1539,In_341);
nand U2486 (N_2486,In_1764,In_2017);
xnor U2487 (N_2487,In_841,In_689);
xor U2488 (N_2488,In_2880,In_2221);
xor U2489 (N_2489,In_1752,In_2825);
nand U2490 (N_2490,In_2735,In_528);
nand U2491 (N_2491,In_872,In_2227);
nand U2492 (N_2492,In_2691,In_1339);
and U2493 (N_2493,In_306,In_507);
nor U2494 (N_2494,In_1965,In_2347);
and U2495 (N_2495,In_1165,In_838);
or U2496 (N_2496,In_1938,In_2859);
or U2497 (N_2497,In_1729,In_2838);
nand U2498 (N_2498,In_2207,In_479);
nor U2499 (N_2499,In_1372,In_825);
xnor U2500 (N_2500,In_1711,In_1262);
or U2501 (N_2501,In_849,In_1298);
nand U2502 (N_2502,In_1874,In_1123);
nand U2503 (N_2503,In_1013,In_159);
nor U2504 (N_2504,In_267,In_1559);
nor U2505 (N_2505,In_830,In_715);
or U2506 (N_2506,In_2848,In_1495);
or U2507 (N_2507,In_42,In_2125);
nor U2508 (N_2508,In_640,In_2369);
or U2509 (N_2509,In_2459,In_587);
and U2510 (N_2510,In_623,In_2345);
nor U2511 (N_2511,In_2610,In_2078);
nand U2512 (N_2512,In_364,In_2629);
and U2513 (N_2513,In_2781,In_2971);
or U2514 (N_2514,In_2110,In_473);
and U2515 (N_2515,In_153,In_1600);
nor U2516 (N_2516,In_2122,In_1906);
xor U2517 (N_2517,In_4,In_1429);
and U2518 (N_2518,In_1307,In_797);
or U2519 (N_2519,In_157,In_1737);
and U2520 (N_2520,In_939,In_931);
xnor U2521 (N_2521,In_251,In_2027);
nand U2522 (N_2522,In_1453,In_1566);
nand U2523 (N_2523,In_2788,In_992);
xnor U2524 (N_2524,In_1662,In_873);
xor U2525 (N_2525,In_2275,In_1445);
or U2526 (N_2526,In_203,In_2902);
nand U2527 (N_2527,In_1556,In_1288);
xnor U2528 (N_2528,In_1452,In_1321);
or U2529 (N_2529,In_757,In_592);
xor U2530 (N_2530,In_1091,In_1717);
nand U2531 (N_2531,In_1474,In_1363);
and U2532 (N_2532,In_2300,In_2149);
or U2533 (N_2533,In_233,In_2498);
and U2534 (N_2534,In_2577,In_1809);
or U2535 (N_2535,In_2723,In_2736);
or U2536 (N_2536,In_2073,In_2298);
nand U2537 (N_2537,In_345,In_909);
and U2538 (N_2538,In_167,In_627);
xor U2539 (N_2539,In_342,In_1041);
nor U2540 (N_2540,In_2175,In_2010);
nand U2541 (N_2541,In_2013,In_2868);
nand U2542 (N_2542,In_1726,In_1909);
and U2543 (N_2543,In_1438,In_2544);
xnor U2544 (N_2544,In_515,In_271);
nor U2545 (N_2545,In_1814,In_1396);
nor U2546 (N_2546,In_1778,In_1904);
nand U2547 (N_2547,In_273,In_324);
nor U2548 (N_2548,In_2901,In_1076);
nor U2549 (N_2549,In_2171,In_1462);
nor U2550 (N_2550,In_351,In_1423);
nor U2551 (N_2551,In_434,In_1554);
or U2552 (N_2552,In_1823,In_2192);
xor U2553 (N_2553,In_691,In_2988);
xor U2554 (N_2554,In_1812,In_762);
and U2555 (N_2555,In_1539,In_2183);
or U2556 (N_2556,In_1284,In_2349);
or U2557 (N_2557,In_2433,In_2929);
or U2558 (N_2558,In_1532,In_202);
nor U2559 (N_2559,In_2471,In_252);
or U2560 (N_2560,In_952,In_1324);
nand U2561 (N_2561,In_585,In_283);
nand U2562 (N_2562,In_2580,In_821);
nor U2563 (N_2563,In_2385,In_2408);
or U2564 (N_2564,In_1036,In_2250);
xnor U2565 (N_2565,In_155,In_707);
xnor U2566 (N_2566,In_244,In_1761);
nand U2567 (N_2567,In_1887,In_2349);
nand U2568 (N_2568,In_1595,In_1244);
and U2569 (N_2569,In_1873,In_2343);
nor U2570 (N_2570,In_1680,In_94);
or U2571 (N_2571,In_408,In_1701);
nand U2572 (N_2572,In_6,In_1122);
nand U2573 (N_2573,In_2146,In_2260);
nor U2574 (N_2574,In_107,In_2200);
nor U2575 (N_2575,In_1248,In_2721);
xnor U2576 (N_2576,In_1930,In_498);
nand U2577 (N_2577,In_1087,In_2195);
xnor U2578 (N_2578,In_2133,In_1936);
or U2579 (N_2579,In_1361,In_1932);
nand U2580 (N_2580,In_20,In_1910);
nor U2581 (N_2581,In_1701,In_944);
nand U2582 (N_2582,In_2694,In_922);
and U2583 (N_2583,In_1011,In_1373);
nor U2584 (N_2584,In_1704,In_1414);
nor U2585 (N_2585,In_970,In_2527);
and U2586 (N_2586,In_2535,In_2373);
nand U2587 (N_2587,In_1708,In_37);
nor U2588 (N_2588,In_1245,In_1431);
nor U2589 (N_2589,In_1278,In_788);
nand U2590 (N_2590,In_2747,In_294);
nand U2591 (N_2591,In_2309,In_562);
nor U2592 (N_2592,In_2264,In_1438);
nand U2593 (N_2593,In_329,In_1187);
nor U2594 (N_2594,In_1220,In_1094);
or U2595 (N_2595,In_1417,In_2857);
or U2596 (N_2596,In_2302,In_1487);
xor U2597 (N_2597,In_1347,In_1976);
nor U2598 (N_2598,In_2429,In_1067);
nor U2599 (N_2599,In_621,In_1091);
and U2600 (N_2600,In_2296,In_2343);
and U2601 (N_2601,In_0,In_536);
xnor U2602 (N_2602,In_2023,In_387);
or U2603 (N_2603,In_1617,In_2466);
xnor U2604 (N_2604,In_2612,In_99);
and U2605 (N_2605,In_2084,In_2993);
xor U2606 (N_2606,In_1549,In_2065);
nand U2607 (N_2607,In_548,In_287);
and U2608 (N_2608,In_2673,In_2731);
nor U2609 (N_2609,In_2583,In_1379);
or U2610 (N_2610,In_1993,In_1221);
xor U2611 (N_2611,In_438,In_1448);
nor U2612 (N_2612,In_613,In_1598);
nand U2613 (N_2613,In_2524,In_1738);
and U2614 (N_2614,In_1818,In_367);
xnor U2615 (N_2615,In_756,In_1445);
xor U2616 (N_2616,In_515,In_2473);
nor U2617 (N_2617,In_78,In_183);
or U2618 (N_2618,In_1762,In_2906);
xnor U2619 (N_2619,In_1193,In_2802);
nand U2620 (N_2620,In_2188,In_1412);
nor U2621 (N_2621,In_2994,In_2933);
nor U2622 (N_2622,In_2283,In_2325);
and U2623 (N_2623,In_2769,In_1115);
nand U2624 (N_2624,In_176,In_666);
nor U2625 (N_2625,In_1959,In_2177);
and U2626 (N_2626,In_1954,In_2142);
nand U2627 (N_2627,In_2887,In_2284);
xor U2628 (N_2628,In_579,In_582);
or U2629 (N_2629,In_791,In_2275);
and U2630 (N_2630,In_381,In_1534);
and U2631 (N_2631,In_2644,In_557);
nor U2632 (N_2632,In_2733,In_1018);
nor U2633 (N_2633,In_2002,In_2731);
xnor U2634 (N_2634,In_59,In_2620);
and U2635 (N_2635,In_16,In_1173);
or U2636 (N_2636,In_1073,In_2232);
nand U2637 (N_2637,In_2072,In_783);
nand U2638 (N_2638,In_1818,In_811);
nand U2639 (N_2639,In_294,In_1262);
nor U2640 (N_2640,In_1568,In_1533);
or U2641 (N_2641,In_2214,In_1151);
xnor U2642 (N_2642,In_620,In_1214);
nor U2643 (N_2643,In_1404,In_801);
and U2644 (N_2644,In_2300,In_161);
and U2645 (N_2645,In_1678,In_626);
nand U2646 (N_2646,In_2548,In_867);
nand U2647 (N_2647,In_751,In_2793);
xnor U2648 (N_2648,In_703,In_56);
xnor U2649 (N_2649,In_2020,In_1438);
nor U2650 (N_2650,In_2449,In_217);
nor U2651 (N_2651,In_1461,In_1981);
nor U2652 (N_2652,In_102,In_14);
nand U2653 (N_2653,In_487,In_783);
nand U2654 (N_2654,In_175,In_1172);
nand U2655 (N_2655,In_125,In_2007);
or U2656 (N_2656,In_2663,In_1211);
nor U2657 (N_2657,In_410,In_836);
or U2658 (N_2658,In_375,In_1798);
nor U2659 (N_2659,In_981,In_2612);
xor U2660 (N_2660,In_2644,In_2604);
xnor U2661 (N_2661,In_574,In_541);
nor U2662 (N_2662,In_1803,In_859);
nor U2663 (N_2663,In_1915,In_981);
nand U2664 (N_2664,In_2007,In_2899);
and U2665 (N_2665,In_1442,In_1580);
and U2666 (N_2666,In_102,In_1778);
or U2667 (N_2667,In_2139,In_2165);
and U2668 (N_2668,In_2845,In_1061);
or U2669 (N_2669,In_493,In_1661);
nor U2670 (N_2670,In_713,In_1291);
nor U2671 (N_2671,In_1797,In_1266);
and U2672 (N_2672,In_720,In_1696);
nor U2673 (N_2673,In_1007,In_737);
or U2674 (N_2674,In_2746,In_948);
nand U2675 (N_2675,In_1856,In_2372);
nand U2676 (N_2676,In_1326,In_943);
and U2677 (N_2677,In_1978,In_2171);
or U2678 (N_2678,In_146,In_1205);
nor U2679 (N_2679,In_912,In_45);
or U2680 (N_2680,In_93,In_2367);
and U2681 (N_2681,In_2763,In_1572);
xnor U2682 (N_2682,In_208,In_2373);
or U2683 (N_2683,In_2386,In_2765);
xnor U2684 (N_2684,In_2678,In_2079);
nand U2685 (N_2685,In_1371,In_2563);
nand U2686 (N_2686,In_666,In_1760);
nor U2687 (N_2687,In_2770,In_438);
xor U2688 (N_2688,In_1419,In_84);
nor U2689 (N_2689,In_2843,In_2574);
nand U2690 (N_2690,In_382,In_1994);
or U2691 (N_2691,In_2675,In_456);
and U2692 (N_2692,In_1361,In_1913);
nand U2693 (N_2693,In_1748,In_176);
xnor U2694 (N_2694,In_1369,In_938);
or U2695 (N_2695,In_1586,In_2509);
xor U2696 (N_2696,In_2115,In_2697);
nand U2697 (N_2697,In_2421,In_2266);
xnor U2698 (N_2698,In_1762,In_2775);
or U2699 (N_2699,In_1992,In_2792);
nand U2700 (N_2700,In_927,In_1279);
or U2701 (N_2701,In_2124,In_321);
xor U2702 (N_2702,In_2479,In_827);
nand U2703 (N_2703,In_2802,In_1852);
nor U2704 (N_2704,In_691,In_2630);
or U2705 (N_2705,In_2226,In_1171);
xnor U2706 (N_2706,In_470,In_136);
xnor U2707 (N_2707,In_2415,In_1056);
nor U2708 (N_2708,In_793,In_2243);
nor U2709 (N_2709,In_2742,In_312);
and U2710 (N_2710,In_1770,In_679);
and U2711 (N_2711,In_2599,In_1594);
nor U2712 (N_2712,In_1186,In_302);
nor U2713 (N_2713,In_1061,In_524);
and U2714 (N_2714,In_2528,In_2760);
and U2715 (N_2715,In_764,In_945);
nor U2716 (N_2716,In_2106,In_1842);
and U2717 (N_2717,In_2316,In_474);
or U2718 (N_2718,In_2749,In_389);
nand U2719 (N_2719,In_2452,In_940);
nand U2720 (N_2720,In_2870,In_253);
xnor U2721 (N_2721,In_1230,In_474);
xnor U2722 (N_2722,In_1424,In_283);
and U2723 (N_2723,In_2106,In_1780);
nor U2724 (N_2724,In_1204,In_1330);
nor U2725 (N_2725,In_32,In_2290);
and U2726 (N_2726,In_2419,In_2414);
or U2727 (N_2727,In_1458,In_2770);
xnor U2728 (N_2728,In_719,In_747);
or U2729 (N_2729,In_190,In_1355);
nand U2730 (N_2730,In_2070,In_1505);
or U2731 (N_2731,In_2403,In_1185);
or U2732 (N_2732,In_1183,In_2968);
xor U2733 (N_2733,In_1110,In_1875);
nor U2734 (N_2734,In_1359,In_2061);
or U2735 (N_2735,In_2789,In_2468);
xor U2736 (N_2736,In_188,In_992);
nand U2737 (N_2737,In_1458,In_2611);
xor U2738 (N_2738,In_2222,In_2205);
and U2739 (N_2739,In_569,In_794);
nand U2740 (N_2740,In_140,In_926);
or U2741 (N_2741,In_174,In_1488);
and U2742 (N_2742,In_1765,In_1134);
or U2743 (N_2743,In_2098,In_2437);
nor U2744 (N_2744,In_40,In_1392);
nand U2745 (N_2745,In_1958,In_2458);
and U2746 (N_2746,In_1397,In_570);
nand U2747 (N_2747,In_2130,In_1919);
nand U2748 (N_2748,In_2657,In_1211);
nor U2749 (N_2749,In_2999,In_217);
nor U2750 (N_2750,In_2253,In_1807);
or U2751 (N_2751,In_2138,In_1979);
or U2752 (N_2752,In_1710,In_1796);
nor U2753 (N_2753,In_2229,In_1932);
nor U2754 (N_2754,In_345,In_790);
or U2755 (N_2755,In_1592,In_971);
and U2756 (N_2756,In_243,In_2314);
and U2757 (N_2757,In_2548,In_213);
nor U2758 (N_2758,In_180,In_338);
and U2759 (N_2759,In_2641,In_2649);
and U2760 (N_2760,In_675,In_2415);
nor U2761 (N_2761,In_1891,In_1526);
and U2762 (N_2762,In_2471,In_2093);
xor U2763 (N_2763,In_219,In_297);
xnor U2764 (N_2764,In_951,In_932);
xnor U2765 (N_2765,In_2986,In_889);
nand U2766 (N_2766,In_342,In_2237);
xor U2767 (N_2767,In_1614,In_2802);
and U2768 (N_2768,In_1608,In_935);
nand U2769 (N_2769,In_2140,In_653);
and U2770 (N_2770,In_659,In_899);
or U2771 (N_2771,In_1501,In_1514);
nor U2772 (N_2772,In_2685,In_1005);
xor U2773 (N_2773,In_786,In_2210);
or U2774 (N_2774,In_188,In_494);
and U2775 (N_2775,In_1545,In_2927);
xnor U2776 (N_2776,In_1581,In_355);
and U2777 (N_2777,In_2107,In_2659);
nand U2778 (N_2778,In_531,In_2262);
nand U2779 (N_2779,In_1930,In_2909);
nand U2780 (N_2780,In_2527,In_674);
nand U2781 (N_2781,In_897,In_401);
or U2782 (N_2782,In_1539,In_2608);
nor U2783 (N_2783,In_398,In_1308);
nand U2784 (N_2784,In_561,In_1345);
or U2785 (N_2785,In_1363,In_2906);
and U2786 (N_2786,In_2780,In_2157);
nand U2787 (N_2787,In_805,In_2037);
and U2788 (N_2788,In_2957,In_2197);
nand U2789 (N_2789,In_2726,In_1705);
xnor U2790 (N_2790,In_2415,In_2273);
xnor U2791 (N_2791,In_1956,In_2792);
or U2792 (N_2792,In_1933,In_1829);
or U2793 (N_2793,In_1937,In_2430);
nand U2794 (N_2794,In_292,In_184);
and U2795 (N_2795,In_1333,In_2837);
or U2796 (N_2796,In_1195,In_126);
xnor U2797 (N_2797,In_1147,In_800);
or U2798 (N_2798,In_1458,In_873);
or U2799 (N_2799,In_1431,In_2704);
nand U2800 (N_2800,In_2670,In_127);
and U2801 (N_2801,In_1907,In_2084);
nor U2802 (N_2802,In_254,In_1375);
and U2803 (N_2803,In_1139,In_2376);
and U2804 (N_2804,In_1729,In_1085);
xor U2805 (N_2805,In_1349,In_479);
nand U2806 (N_2806,In_2934,In_1321);
or U2807 (N_2807,In_2673,In_718);
or U2808 (N_2808,In_2483,In_2526);
nand U2809 (N_2809,In_2771,In_1395);
or U2810 (N_2810,In_349,In_229);
nor U2811 (N_2811,In_2357,In_1243);
nor U2812 (N_2812,In_2242,In_11);
xor U2813 (N_2813,In_325,In_526);
or U2814 (N_2814,In_2880,In_1395);
or U2815 (N_2815,In_1018,In_877);
nand U2816 (N_2816,In_1953,In_1911);
xnor U2817 (N_2817,In_923,In_2756);
xnor U2818 (N_2818,In_1774,In_601);
or U2819 (N_2819,In_1108,In_1049);
nor U2820 (N_2820,In_2761,In_477);
or U2821 (N_2821,In_1600,In_1494);
and U2822 (N_2822,In_1765,In_2101);
and U2823 (N_2823,In_1625,In_2439);
or U2824 (N_2824,In_369,In_1748);
and U2825 (N_2825,In_2664,In_1175);
and U2826 (N_2826,In_2773,In_1211);
nand U2827 (N_2827,In_2697,In_1511);
or U2828 (N_2828,In_1124,In_483);
nor U2829 (N_2829,In_2530,In_1246);
nor U2830 (N_2830,In_537,In_1746);
nor U2831 (N_2831,In_1423,In_1159);
or U2832 (N_2832,In_1348,In_1028);
or U2833 (N_2833,In_1788,In_1655);
nand U2834 (N_2834,In_2207,In_1881);
and U2835 (N_2835,In_2164,In_1710);
xnor U2836 (N_2836,In_2766,In_2192);
or U2837 (N_2837,In_2064,In_146);
nor U2838 (N_2838,In_2996,In_2573);
nand U2839 (N_2839,In_2130,In_1656);
or U2840 (N_2840,In_1183,In_1943);
or U2841 (N_2841,In_512,In_1426);
and U2842 (N_2842,In_2645,In_1795);
xor U2843 (N_2843,In_640,In_793);
nand U2844 (N_2844,In_2834,In_1832);
nand U2845 (N_2845,In_1224,In_1444);
and U2846 (N_2846,In_2528,In_526);
and U2847 (N_2847,In_2226,In_1492);
xnor U2848 (N_2848,In_2519,In_145);
xor U2849 (N_2849,In_1118,In_1802);
nor U2850 (N_2850,In_2123,In_1133);
or U2851 (N_2851,In_704,In_2694);
or U2852 (N_2852,In_315,In_581);
xnor U2853 (N_2853,In_1881,In_2197);
or U2854 (N_2854,In_2889,In_941);
nor U2855 (N_2855,In_1142,In_2398);
nor U2856 (N_2856,In_2878,In_968);
and U2857 (N_2857,In_2795,In_2688);
and U2858 (N_2858,In_2656,In_1979);
nand U2859 (N_2859,In_577,In_2328);
xor U2860 (N_2860,In_37,In_1767);
or U2861 (N_2861,In_724,In_596);
and U2862 (N_2862,In_2510,In_1723);
nor U2863 (N_2863,In_359,In_720);
xnor U2864 (N_2864,In_403,In_2416);
or U2865 (N_2865,In_292,In_1928);
nand U2866 (N_2866,In_1957,In_2258);
xor U2867 (N_2867,In_110,In_386);
and U2868 (N_2868,In_726,In_1956);
nand U2869 (N_2869,In_2410,In_1999);
xor U2870 (N_2870,In_2101,In_371);
nand U2871 (N_2871,In_813,In_815);
nor U2872 (N_2872,In_1771,In_2686);
xnor U2873 (N_2873,In_2247,In_2529);
and U2874 (N_2874,In_1817,In_2674);
xnor U2875 (N_2875,In_639,In_1612);
xor U2876 (N_2876,In_1827,In_957);
xnor U2877 (N_2877,In_1169,In_1082);
and U2878 (N_2878,In_2569,In_1116);
nand U2879 (N_2879,In_2965,In_864);
xor U2880 (N_2880,In_2485,In_223);
or U2881 (N_2881,In_954,In_2333);
xor U2882 (N_2882,In_1516,In_1615);
nor U2883 (N_2883,In_1296,In_2847);
nor U2884 (N_2884,In_2278,In_46);
and U2885 (N_2885,In_142,In_2804);
and U2886 (N_2886,In_2397,In_2332);
xnor U2887 (N_2887,In_2478,In_1261);
nor U2888 (N_2888,In_2714,In_2000);
nor U2889 (N_2889,In_2814,In_1663);
nor U2890 (N_2890,In_132,In_1765);
xnor U2891 (N_2891,In_278,In_973);
and U2892 (N_2892,In_50,In_2203);
nand U2893 (N_2893,In_2572,In_1535);
or U2894 (N_2894,In_2002,In_1794);
or U2895 (N_2895,In_603,In_2405);
or U2896 (N_2896,In_1779,In_1536);
or U2897 (N_2897,In_2927,In_2671);
and U2898 (N_2898,In_973,In_267);
or U2899 (N_2899,In_1471,In_647);
xnor U2900 (N_2900,In_2466,In_1057);
nand U2901 (N_2901,In_653,In_2339);
nor U2902 (N_2902,In_591,In_2770);
nand U2903 (N_2903,In_561,In_1146);
nor U2904 (N_2904,In_832,In_1695);
nor U2905 (N_2905,In_875,In_2196);
nand U2906 (N_2906,In_1445,In_342);
xor U2907 (N_2907,In_1669,In_1424);
and U2908 (N_2908,In_676,In_1853);
and U2909 (N_2909,In_446,In_1);
xor U2910 (N_2910,In_561,In_1989);
nand U2911 (N_2911,In_2689,In_2368);
nor U2912 (N_2912,In_1735,In_1723);
nor U2913 (N_2913,In_1571,In_1082);
or U2914 (N_2914,In_1836,In_1227);
nor U2915 (N_2915,In_977,In_1364);
xnor U2916 (N_2916,In_2989,In_2573);
nand U2917 (N_2917,In_381,In_2862);
nor U2918 (N_2918,In_1807,In_2074);
xor U2919 (N_2919,In_2490,In_1183);
nor U2920 (N_2920,In_1438,In_2649);
nand U2921 (N_2921,In_829,In_2756);
and U2922 (N_2922,In_2657,In_817);
xnor U2923 (N_2923,In_1157,In_232);
nor U2924 (N_2924,In_2791,In_601);
and U2925 (N_2925,In_1708,In_2706);
xnor U2926 (N_2926,In_1319,In_1571);
xor U2927 (N_2927,In_1651,In_2029);
and U2928 (N_2928,In_849,In_2558);
nand U2929 (N_2929,In_1801,In_886);
nand U2930 (N_2930,In_2123,In_1356);
nor U2931 (N_2931,In_1415,In_1417);
and U2932 (N_2932,In_2472,In_2690);
nand U2933 (N_2933,In_1549,In_1433);
and U2934 (N_2934,In_1256,In_418);
and U2935 (N_2935,In_577,In_1497);
xnor U2936 (N_2936,In_874,In_2906);
or U2937 (N_2937,In_2097,In_2872);
nor U2938 (N_2938,In_2860,In_223);
nand U2939 (N_2939,In_746,In_1671);
nor U2940 (N_2940,In_1843,In_2140);
xor U2941 (N_2941,In_1291,In_2379);
xor U2942 (N_2942,In_2363,In_2249);
nand U2943 (N_2943,In_18,In_259);
nand U2944 (N_2944,In_637,In_551);
or U2945 (N_2945,In_171,In_1668);
nor U2946 (N_2946,In_1696,In_2233);
xnor U2947 (N_2947,In_1939,In_1778);
and U2948 (N_2948,In_663,In_280);
xor U2949 (N_2949,In_2671,In_461);
or U2950 (N_2950,In_2797,In_2384);
xnor U2951 (N_2951,In_1149,In_932);
nor U2952 (N_2952,In_1417,In_2391);
or U2953 (N_2953,In_1585,In_2955);
and U2954 (N_2954,In_1668,In_2679);
nor U2955 (N_2955,In_1862,In_363);
nand U2956 (N_2956,In_198,In_2976);
xnor U2957 (N_2957,In_927,In_2570);
xnor U2958 (N_2958,In_2807,In_2359);
and U2959 (N_2959,In_887,In_2237);
nor U2960 (N_2960,In_1185,In_971);
nand U2961 (N_2961,In_704,In_1852);
xor U2962 (N_2962,In_2119,In_150);
and U2963 (N_2963,In_434,In_2573);
or U2964 (N_2964,In_1508,In_2322);
nor U2965 (N_2965,In_2641,In_1972);
nand U2966 (N_2966,In_1968,In_2411);
nand U2967 (N_2967,In_868,In_1887);
or U2968 (N_2968,In_2648,In_2952);
nor U2969 (N_2969,In_2211,In_815);
nor U2970 (N_2970,In_1814,In_273);
nand U2971 (N_2971,In_807,In_2688);
and U2972 (N_2972,In_44,In_2261);
nor U2973 (N_2973,In_897,In_326);
xor U2974 (N_2974,In_386,In_159);
xor U2975 (N_2975,In_2687,In_1631);
or U2976 (N_2976,In_494,In_967);
nand U2977 (N_2977,In_285,In_2737);
xnor U2978 (N_2978,In_1920,In_2780);
nand U2979 (N_2979,In_307,In_1221);
xnor U2980 (N_2980,In_41,In_2331);
and U2981 (N_2981,In_2991,In_939);
or U2982 (N_2982,In_1598,In_2476);
nand U2983 (N_2983,In_2061,In_1349);
and U2984 (N_2984,In_692,In_720);
and U2985 (N_2985,In_2688,In_1780);
nand U2986 (N_2986,In_348,In_2307);
and U2987 (N_2987,In_1526,In_1819);
nand U2988 (N_2988,In_1086,In_1123);
nor U2989 (N_2989,In_374,In_954);
or U2990 (N_2990,In_2462,In_2617);
and U2991 (N_2991,In_1380,In_1866);
xnor U2992 (N_2992,In_1041,In_1304);
nand U2993 (N_2993,In_2619,In_174);
xnor U2994 (N_2994,In_267,In_679);
and U2995 (N_2995,In_302,In_2754);
nor U2996 (N_2996,In_397,In_2516);
and U2997 (N_2997,In_1704,In_781);
nand U2998 (N_2998,In_530,In_1555);
xnor U2999 (N_2999,In_1354,In_754);
xnor U3000 (N_3000,N_618,N_613);
or U3001 (N_3001,N_1683,N_2449);
xnor U3002 (N_3002,N_2128,N_1898);
nand U3003 (N_3003,N_2303,N_1818);
nand U3004 (N_3004,N_2656,N_2079);
xnor U3005 (N_3005,N_1038,N_1511);
nor U3006 (N_3006,N_1870,N_1045);
or U3007 (N_3007,N_1638,N_201);
and U3008 (N_3008,N_1396,N_2609);
or U3009 (N_3009,N_2693,N_1285);
and U3010 (N_3010,N_973,N_2274);
nor U3011 (N_3011,N_2617,N_2942);
or U3012 (N_3012,N_635,N_1086);
or U3013 (N_3013,N_1208,N_1163);
or U3014 (N_3014,N_2275,N_196);
and U3015 (N_3015,N_2721,N_2711);
nand U3016 (N_3016,N_284,N_1185);
nand U3017 (N_3017,N_655,N_2227);
and U3018 (N_3018,N_473,N_1212);
xor U3019 (N_3019,N_865,N_1798);
nor U3020 (N_3020,N_1630,N_1657);
nand U3021 (N_3021,N_146,N_1747);
or U3022 (N_3022,N_104,N_598);
and U3023 (N_3023,N_647,N_2608);
nand U3024 (N_3024,N_519,N_288);
nand U3025 (N_3025,N_1131,N_2252);
nor U3026 (N_3026,N_2030,N_282);
or U3027 (N_3027,N_1112,N_2395);
or U3028 (N_3028,N_2806,N_2421);
xor U3029 (N_3029,N_2097,N_814);
xor U3030 (N_3030,N_1335,N_315);
and U3031 (N_3031,N_2394,N_553);
nand U3032 (N_3032,N_2329,N_1850);
nand U3033 (N_3033,N_2888,N_1017);
nand U3034 (N_3034,N_596,N_1559);
and U3035 (N_3035,N_2927,N_1840);
and U3036 (N_3036,N_2546,N_960);
xnor U3037 (N_3037,N_1391,N_513);
and U3038 (N_3038,N_1243,N_2971);
nor U3039 (N_3039,N_1398,N_795);
xor U3040 (N_3040,N_2054,N_7);
xor U3041 (N_3041,N_2382,N_2388);
nor U3042 (N_3042,N_2095,N_2920);
xnor U3043 (N_3043,N_692,N_2034);
nand U3044 (N_3044,N_1861,N_2710);
nor U3045 (N_3045,N_211,N_788);
nand U3046 (N_3046,N_2154,N_1283);
nor U3047 (N_3047,N_2177,N_538);
nand U3048 (N_3048,N_730,N_10);
and U3049 (N_3049,N_1535,N_1634);
and U3050 (N_3050,N_1232,N_564);
or U3051 (N_3051,N_2381,N_2293);
and U3052 (N_3052,N_1351,N_593);
nand U3053 (N_3053,N_2183,N_1292);
nand U3054 (N_3054,N_2135,N_653);
xor U3055 (N_3055,N_911,N_1701);
and U3056 (N_3056,N_2073,N_509);
nand U3057 (N_3057,N_2545,N_1831);
or U3058 (N_3058,N_2323,N_2651);
xnor U3059 (N_3059,N_1375,N_1011);
nand U3060 (N_3060,N_1247,N_1200);
nand U3061 (N_3061,N_1712,N_2782);
nand U3062 (N_3062,N_1382,N_1151);
nor U3063 (N_3063,N_505,N_2318);
xor U3064 (N_3064,N_1482,N_1230);
xnor U3065 (N_3065,N_1126,N_1052);
xor U3066 (N_3066,N_1751,N_1893);
and U3067 (N_3067,N_2064,N_1580);
or U3068 (N_3068,N_1955,N_2846);
and U3069 (N_3069,N_2899,N_1682);
and U3070 (N_3070,N_2083,N_1229);
and U3071 (N_3071,N_169,N_714);
or U3072 (N_3072,N_1841,N_1012);
nor U3073 (N_3073,N_2103,N_890);
and U3074 (N_3074,N_417,N_1311);
and U3075 (N_3075,N_1463,N_1871);
nor U3076 (N_3076,N_2560,N_851);
nand U3077 (N_3077,N_457,N_2251);
nand U3078 (N_3078,N_1291,N_834);
xor U3079 (N_3079,N_486,N_1828);
nor U3080 (N_3080,N_2984,N_2526);
nand U3081 (N_3081,N_1259,N_1079);
xor U3082 (N_3082,N_265,N_2758);
and U3083 (N_3083,N_250,N_2533);
nand U3084 (N_3084,N_2088,N_1958);
nor U3085 (N_3085,N_2870,N_280);
nor U3086 (N_3086,N_344,N_249);
or U3087 (N_3087,N_2894,N_1813);
nor U3088 (N_3088,N_309,N_1743);
nor U3089 (N_3089,N_1596,N_1923);
nand U3090 (N_3090,N_1250,N_2581);
or U3091 (N_3091,N_1436,N_1280);
and U3092 (N_3092,N_1526,N_1117);
xor U3093 (N_3093,N_2454,N_1114);
xnor U3094 (N_3094,N_212,N_2049);
or U3095 (N_3095,N_2547,N_88);
nor U3096 (N_3096,N_2618,N_1177);
or U3097 (N_3097,N_245,N_337);
nor U3098 (N_3098,N_2360,N_439);
or U3099 (N_3099,N_2181,N_1680);
nand U3100 (N_3100,N_1799,N_218);
xor U3101 (N_3101,N_790,N_2881);
nand U3102 (N_3102,N_979,N_1951);
nor U3103 (N_3103,N_1289,N_2859);
or U3104 (N_3104,N_1990,N_1084);
xnor U3105 (N_3105,N_1889,N_2593);
nor U3106 (N_3106,N_900,N_237);
nor U3107 (N_3107,N_213,N_1197);
and U3108 (N_3108,N_2427,N_1365);
nor U3109 (N_3109,N_651,N_2025);
nand U3110 (N_3110,N_909,N_1171);
nand U3111 (N_3111,N_1096,N_1353);
or U3112 (N_3112,N_2925,N_451);
or U3113 (N_3113,N_2633,N_1306);
nor U3114 (N_3114,N_2489,N_643);
nor U3115 (N_3115,N_1338,N_2813);
nor U3116 (N_3116,N_2759,N_2310);
nor U3117 (N_3117,N_2418,N_312);
and U3118 (N_3118,N_474,N_1183);
nand U3119 (N_3119,N_970,N_2524);
xnor U3120 (N_3120,N_2212,N_722);
xor U3121 (N_3121,N_2527,N_84);
xnor U3122 (N_3122,N_2776,N_2567);
or U3123 (N_3123,N_1920,N_567);
nand U3124 (N_3124,N_1692,N_784);
xnor U3125 (N_3125,N_206,N_2313);
xor U3126 (N_3126,N_132,N_2562);
or U3127 (N_3127,N_1932,N_2820);
nor U3128 (N_3128,N_1325,N_2111);
or U3129 (N_3129,N_159,N_1716);
or U3130 (N_3130,N_264,N_881);
nand U3131 (N_3131,N_1749,N_2844);
or U3132 (N_3132,N_1481,N_2739);
xnor U3133 (N_3133,N_1155,N_1035);
nor U3134 (N_3134,N_310,N_1459);
nand U3135 (N_3135,N_2218,N_378);
or U3136 (N_3136,N_403,N_1890);
nor U3137 (N_3137,N_1165,N_1094);
and U3138 (N_3138,N_397,N_1811);
or U3139 (N_3139,N_414,N_1272);
or U3140 (N_3140,N_2078,N_607);
nand U3141 (N_3141,N_2260,N_2744);
xnor U3142 (N_3142,N_991,N_1862);
and U3143 (N_3143,N_1395,N_1315);
and U3144 (N_3144,N_2455,N_605);
and U3145 (N_3145,N_919,N_2041);
or U3146 (N_3146,N_1191,N_989);
xor U3147 (N_3147,N_2791,N_227);
and U3148 (N_3148,N_1333,N_696);
and U3149 (N_3149,N_2235,N_1342);
xor U3150 (N_3150,N_1872,N_2878);
or U3151 (N_3151,N_1550,N_1790);
or U3152 (N_3152,N_1627,N_1852);
or U3153 (N_3153,N_2977,N_420);
nor U3154 (N_3154,N_2377,N_1153);
xnor U3155 (N_3155,N_1699,N_268);
and U3156 (N_3156,N_2805,N_606);
nor U3157 (N_3157,N_1110,N_1604);
and U3158 (N_3158,N_976,N_1842);
nor U3159 (N_3159,N_828,N_2902);
and U3160 (N_3160,N_1271,N_2043);
or U3161 (N_3161,N_2462,N_1089);
xnor U3162 (N_3162,N_841,N_1521);
nor U3163 (N_3163,N_2819,N_982);
nor U3164 (N_3164,N_359,N_93);
nand U3165 (N_3165,N_117,N_1873);
or U3166 (N_3166,N_2114,N_2331);
xor U3167 (N_3167,N_1132,N_236);
xor U3168 (N_3168,N_511,N_2362);
or U3169 (N_3169,N_2788,N_332);
and U3170 (N_3170,N_2966,N_1694);
nand U3171 (N_3171,N_1928,N_675);
or U3172 (N_3172,N_2487,N_2874);
nor U3173 (N_3173,N_2369,N_929);
nand U3174 (N_3174,N_2745,N_2399);
nand U3175 (N_3175,N_2688,N_543);
or U3176 (N_3176,N_2847,N_1443);
nand U3177 (N_3177,N_1288,N_1925);
or U3178 (N_3178,N_2021,N_2764);
nor U3179 (N_3179,N_1663,N_2226);
or U3180 (N_3180,N_578,N_827);
nand U3181 (N_3181,N_1732,N_380);
nor U3182 (N_3182,N_2386,N_2340);
and U3183 (N_3183,N_2809,N_2150);
nand U3184 (N_3184,N_1464,N_56);
xnor U3185 (N_3185,N_1374,N_1092);
and U3186 (N_3186,N_1565,N_2476);
or U3187 (N_3187,N_2867,N_224);
or U3188 (N_3188,N_782,N_2855);
nor U3189 (N_3189,N_410,N_2722);
or U3190 (N_3190,N_1048,N_835);
xor U3191 (N_3191,N_2193,N_1239);
nor U3192 (N_3192,N_2409,N_1192);
and U3193 (N_3193,N_274,N_1509);
and U3194 (N_3194,N_1707,N_1008);
xor U3195 (N_3195,N_489,N_114);
or U3196 (N_3196,N_456,N_2981);
xor U3197 (N_3197,N_1392,N_604);
and U3198 (N_3198,N_2929,N_2675);
nor U3199 (N_3199,N_1344,N_512);
or U3200 (N_3200,N_2339,N_516);
nor U3201 (N_3201,N_1804,N_16);
nand U3202 (N_3202,N_2668,N_2970);
nor U3203 (N_3203,N_487,N_92);
xor U3204 (N_3204,N_1941,N_1753);
nand U3205 (N_3205,N_1543,N_1942);
nor U3206 (N_3206,N_183,N_2793);
nor U3207 (N_3207,N_2044,N_2324);
nor U3208 (N_3208,N_2731,N_1792);
or U3209 (N_3209,N_147,N_818);
nor U3210 (N_3210,N_2067,N_444);
and U3211 (N_3211,N_1324,N_1300);
xnor U3212 (N_3212,N_2936,N_2900);
nor U3213 (N_3213,N_734,N_2238);
and U3214 (N_3214,N_2792,N_2385);
nand U3215 (N_3215,N_1584,N_2886);
xnor U3216 (N_3216,N_1039,N_317);
nand U3217 (N_3217,N_2954,N_2575);
xnor U3218 (N_3218,N_287,N_1940);
and U3219 (N_3219,N_27,N_2190);
nand U3220 (N_3220,N_770,N_1);
nor U3221 (N_3221,N_51,N_1713);
nor U3222 (N_3222,N_849,N_1946);
or U3223 (N_3223,N_488,N_2845);
xor U3224 (N_3224,N_2007,N_242);
xor U3225 (N_3225,N_703,N_2915);
or U3226 (N_3226,N_2279,N_768);
or U3227 (N_3227,N_2600,N_258);
nand U3228 (N_3228,N_627,N_994);
nor U3229 (N_3229,N_1190,N_2692);
nor U3230 (N_3230,N_2938,N_2176);
xor U3231 (N_3231,N_1671,N_2830);
xor U3232 (N_3232,N_2558,N_176);
nand U3233 (N_3233,N_1181,N_1589);
or U3234 (N_3234,N_531,N_1164);
nor U3235 (N_3235,N_2850,N_353);
xnor U3236 (N_3236,N_2532,N_608);
xor U3237 (N_3237,N_1036,N_1485);
or U3238 (N_3238,N_142,N_1040);
nor U3239 (N_3239,N_244,N_1461);
xnor U3240 (N_3240,N_1269,N_2771);
xnor U3241 (N_3241,N_2725,N_2415);
or U3242 (N_3242,N_2501,N_2093);
xor U3243 (N_3243,N_2167,N_2948);
or U3244 (N_3244,N_1410,N_1927);
nor U3245 (N_3245,N_826,N_921);
or U3246 (N_3246,N_289,N_990);
xnor U3247 (N_3247,N_2307,N_501);
nand U3248 (N_3248,N_1858,N_2991);
and U3249 (N_3249,N_100,N_2282);
nor U3250 (N_3250,N_2854,N_1211);
nor U3251 (N_3251,N_1266,N_431);
nand U3252 (N_3252,N_465,N_1879);
xor U3253 (N_3253,N_1726,N_1445);
and U3254 (N_3254,N_586,N_2736);
or U3255 (N_3255,N_1607,N_185);
nand U3256 (N_3256,N_637,N_755);
nand U3257 (N_3257,N_1063,N_803);
nand U3258 (N_3258,N_573,N_1343);
xor U3259 (N_3259,N_95,N_898);
nor U3260 (N_3260,N_326,N_189);
nor U3261 (N_3261,N_1938,N_2082);
and U3262 (N_3262,N_968,N_1023);
nand U3263 (N_3263,N_1235,N_880);
xor U3264 (N_3264,N_467,N_1959);
xnor U3265 (N_3265,N_219,N_1622);
nand U3266 (N_3266,N_706,N_1275);
nand U3267 (N_3267,N_1406,N_1866);
xor U3268 (N_3268,N_2468,N_188);
nor U3269 (N_3269,N_2892,N_1198);
nand U3270 (N_3270,N_2139,N_2852);
nand U3271 (N_3271,N_2264,N_1549);
and U3272 (N_3272,N_2255,N_937);
and U3273 (N_3273,N_2960,N_666);
nor U3274 (N_3274,N_216,N_978);
or U3275 (N_3275,N_1058,N_2875);
nor U3276 (N_3276,N_1644,N_1625);
xor U3277 (N_3277,N_1546,N_2365);
xnor U3278 (N_3278,N_912,N_1299);
and U3279 (N_3279,N_1782,N_1006);
or U3280 (N_3280,N_1093,N_1158);
nand U3281 (N_3281,N_1655,N_2134);
nand U3282 (N_3282,N_293,N_707);
xnor U3283 (N_3283,N_2587,N_1195);
xnor U3284 (N_3284,N_705,N_2730);
nand U3285 (N_3285,N_1601,N_773);
nor U3286 (N_3286,N_2146,N_1515);
or U3287 (N_3287,N_1797,N_740);
and U3288 (N_3288,N_552,N_471);
nor U3289 (N_3289,N_339,N_1085);
and U3290 (N_3290,N_603,N_1213);
nor U3291 (N_3291,N_1993,N_589);
nand U3292 (N_3292,N_2104,N_2180);
nor U3293 (N_3293,N_744,N_157);
nand U3294 (N_3294,N_2997,N_428);
xor U3295 (N_3295,N_599,N_334);
xor U3296 (N_3296,N_1472,N_934);
nand U3297 (N_3297,N_786,N_616);
and U3298 (N_3298,N_2924,N_1106);
nor U3299 (N_3299,N_2287,N_65);
nand U3300 (N_3300,N_1218,N_861);
and U3301 (N_3301,N_2351,N_2375);
and U3302 (N_3302,N_759,N_1290);
nand U3303 (N_3303,N_1390,N_2374);
or U3304 (N_3304,N_348,N_633);
nand U3305 (N_3305,N_1369,N_761);
xor U3306 (N_3306,N_2160,N_2799);
and U3307 (N_3307,N_2471,N_71);
nor U3308 (N_3308,N_2363,N_2357);
xor U3309 (N_3309,N_376,N_971);
and U3310 (N_3310,N_2740,N_1669);
nand U3311 (N_3311,N_2230,N_1678);
or U3312 (N_3312,N_813,N_430);
nand U3313 (N_3313,N_1567,N_1857);
and U3314 (N_3314,N_229,N_948);
and U3315 (N_3315,N_2045,N_645);
nor U3316 (N_3316,N_1014,N_1834);
xnor U3317 (N_3317,N_402,N_1175);
nand U3318 (N_3318,N_2371,N_847);
nand U3319 (N_3319,N_2572,N_2958);
xnor U3320 (N_3320,N_2963,N_1182);
nand U3321 (N_3321,N_873,N_590);
and U3322 (N_3322,N_98,N_720);
nor U3323 (N_3323,N_2039,N_2108);
nand U3324 (N_3324,N_1825,N_82);
nand U3325 (N_3325,N_278,N_1952);
nor U3326 (N_3326,N_1675,N_178);
nor U3327 (N_3327,N_1849,N_1796);
nand U3328 (N_3328,N_2098,N_2219);
nand U3329 (N_3329,N_314,N_1145);
nor U3330 (N_3330,N_1735,N_1066);
nand U3331 (N_3331,N_498,N_2102);
nand U3332 (N_3332,N_2130,N_1730);
nor U3333 (N_3333,N_2465,N_230);
xnor U3334 (N_3334,N_427,N_2939);
xnor U3335 (N_3335,N_660,N_1108);
nand U3336 (N_3336,N_652,N_2636);
and U3337 (N_3337,N_1746,N_2342);
or U3338 (N_3338,N_1294,N_1314);
nand U3339 (N_3339,N_2109,N_1892);
and U3340 (N_3340,N_2895,N_366);
xnor U3341 (N_3341,N_2442,N_2283);
nor U3342 (N_3342,N_195,N_279);
or U3343 (N_3343,N_850,N_1332);
nand U3344 (N_3344,N_2602,N_2590);
nor U3345 (N_3345,N_2346,N_611);
xor U3346 (N_3346,N_1775,N_601);
or U3347 (N_3347,N_999,N_492);
and U3348 (N_3348,N_2531,N_2300);
and U3349 (N_3349,N_2594,N_2836);
and U3350 (N_3350,N_1400,N_2483);
and U3351 (N_3351,N_1708,N_2988);
and U3352 (N_3352,N_1994,N_2129);
nor U3353 (N_3353,N_2818,N_385);
xor U3354 (N_3354,N_566,N_483);
or U3355 (N_3355,N_685,N_2952);
nor U3356 (N_3356,N_535,N_1965);
and U3357 (N_3357,N_2554,N_412);
or U3358 (N_3358,N_650,N_231);
or U3359 (N_3359,N_1885,N_1317);
and U3360 (N_3360,N_1878,N_832);
and U3361 (N_3361,N_819,N_2519);
nor U3362 (N_3362,N_316,N_1733);
nand U3363 (N_3363,N_2017,N_610);
xor U3364 (N_3364,N_2068,N_1556);
and U3365 (N_3365,N_1054,N_710);
xnor U3366 (N_3366,N_2299,N_554);
nor U3367 (N_3367,N_1523,N_1992);
nor U3368 (N_3368,N_892,N_1805);
and U3369 (N_3369,N_2807,N_2302);
and U3370 (N_3370,N_1217,N_1656);
nor U3371 (N_3371,N_411,N_1019);
nand U3372 (N_3372,N_1128,N_2136);
and U3373 (N_3373,N_1296,N_1659);
nand U3374 (N_3374,N_557,N_2639);
xor U3375 (N_3375,N_2917,N_1109);
nor U3376 (N_3376,N_154,N_2588);
or U3377 (N_3377,N_2426,N_1847);
xor U3378 (N_3378,N_2267,N_331);
and U3379 (N_3379,N_184,N_47);
or U3380 (N_3380,N_9,N_1863);
nand U3381 (N_3381,N_2945,N_2046);
and U3382 (N_3382,N_2990,N_20);
xor U3383 (N_3383,N_2448,N_950);
nor U3384 (N_3384,N_1407,N_1253);
nand U3385 (N_3385,N_2292,N_321);
xor U3386 (N_3386,N_1937,N_2980);
and U3387 (N_3387,N_433,N_2628);
nor U3388 (N_3388,N_2509,N_194);
xnor U3389 (N_3389,N_1537,N_1484);
xnor U3390 (N_3390,N_1608,N_2055);
xnor U3391 (N_3391,N_255,N_2690);
nand U3392 (N_3392,N_83,N_2934);
nand U3393 (N_3393,N_109,N_1767);
xnor U3394 (N_3394,N_2401,N_156);
nand U3395 (N_3395,N_2500,N_676);
or U3396 (N_3396,N_2978,N_1320);
or U3397 (N_3397,N_1826,N_877);
nand U3398 (N_3398,N_1121,N_1224);
nand U3399 (N_3399,N_2753,N_266);
xor U3400 (N_3400,N_2192,N_1843);
nor U3401 (N_3401,N_327,N_700);
or U3402 (N_3402,N_1424,N_1452);
nor U3403 (N_3403,N_1024,N_1427);
nor U3404 (N_3404,N_401,N_137);
nor U3405 (N_3405,N_384,N_1677);
and U3406 (N_3406,N_1493,N_1667);
nor U3407 (N_3407,N_563,N_1950);
nand U3408 (N_3408,N_199,N_358);
nand U3409 (N_3409,N_285,N_895);
nor U3410 (N_3410,N_2992,N_2175);
xnor U3411 (N_3411,N_240,N_1136);
or U3412 (N_3412,N_1724,N_2796);
and U3413 (N_3413,N_1676,N_2277);
and U3414 (N_3414,N_1104,N_526);
nor U3415 (N_3415,N_2622,N_935);
or U3416 (N_3416,N_259,N_152);
and U3417 (N_3417,N_1022,N_924);
and U3418 (N_3418,N_517,N_1557);
and U3419 (N_3419,N_2271,N_2151);
and U3420 (N_3420,N_1803,N_2148);
nand U3421 (N_3421,N_1711,N_2557);
or U3422 (N_3422,N_2775,N_2967);
nand U3423 (N_3423,N_872,N_271);
nand U3424 (N_3424,N_391,N_329);
or U3425 (N_3425,N_1491,N_130);
nand U3426 (N_3426,N_942,N_1379);
nor U3427 (N_3427,N_1100,N_1293);
xor U3428 (N_3428,N_179,N_2170);
xnor U3429 (N_3429,N_2657,N_1623);
xor U3430 (N_3430,N_2076,N_1168);
nor U3431 (N_3431,N_2539,N_2512);
and U3432 (N_3432,N_1483,N_2795);
xor U3433 (N_3433,N_1912,N_2478);
nand U3434 (N_3434,N_1610,N_1929);
or U3435 (N_3435,N_2406,N_1430);
nor U3436 (N_3436,N_1897,N_712);
or U3437 (N_3437,N_134,N_2420);
nor U3438 (N_3438,N_985,N_1738);
and U3439 (N_3439,N_1078,N_779);
xor U3440 (N_3440,N_263,N_139);
and U3441 (N_3441,N_1575,N_736);
xnor U3442 (N_3442,N_17,N_1702);
nor U3443 (N_3443,N_787,N_899);
xnor U3444 (N_3444,N_732,N_737);
or U3445 (N_3445,N_1416,N_558);
and U3446 (N_3446,N_241,N_629);
and U3447 (N_3447,N_772,N_115);
nand U3448 (N_3448,N_1116,N_2432);
or U3449 (N_3449,N_2889,N_1144);
nand U3450 (N_3450,N_1836,N_2451);
xor U3451 (N_3451,N_1974,N_1073);
xor U3452 (N_3452,N_129,N_182);
and U3453 (N_3453,N_1868,N_1612);
nand U3454 (N_3454,N_2215,N_76);
nor U3455 (N_3455,N_580,N_1532);
xnor U3456 (N_3456,N_682,N_717);
nor U3457 (N_3457,N_2695,N_1323);
nor U3458 (N_3458,N_1460,N_1624);
xnor U3459 (N_3459,N_2762,N_2872);
nor U3460 (N_3460,N_187,N_2194);
or U3461 (N_3461,N_1635,N_1563);
nor U3462 (N_3462,N_2428,N_2290);
nor U3463 (N_3463,N_1513,N_571);
nor U3464 (N_3464,N_582,N_2564);
xor U3465 (N_3465,N_2376,N_515);
xor U3466 (N_3466,N_2140,N_1997);
or U3467 (N_3467,N_728,N_1529);
or U3468 (N_3468,N_2770,N_1152);
nand U3469 (N_3469,N_2325,N_1984);
nor U3470 (N_3470,N_2514,N_50);
nor U3471 (N_3471,N_848,N_754);
nor U3472 (N_3472,N_998,N_2957);
nand U3473 (N_3473,N_1772,N_2332);
and U3474 (N_3474,N_1069,N_1361);
xor U3475 (N_3475,N_1238,N_2172);
xnor U3476 (N_3476,N_2520,N_72);
or U3477 (N_3477,N_260,N_1322);
nor U3478 (N_3478,N_2220,N_933);
xnor U3479 (N_3479,N_177,N_1639);
nor U3480 (N_3480,N_1824,N_1422);
or U3481 (N_3481,N_1367,N_2295);
nor U3482 (N_3482,N_2660,N_1387);
nand U3483 (N_3483,N_1789,N_2918);
or U3484 (N_3484,N_1651,N_2502);
or U3485 (N_3485,N_302,N_407);
or U3486 (N_3486,N_1935,N_2666);
or U3487 (N_3487,N_2490,N_2281);
xor U3488 (N_3488,N_1835,N_63);
and U3489 (N_3489,N_1966,N_12);
nor U3490 (N_3490,N_2051,N_2569);
xor U3491 (N_3491,N_5,N_1970);
and U3492 (N_3492,N_1267,N_2998);
xor U3493 (N_3493,N_1770,N_2595);
and U3494 (N_3494,N_447,N_2833);
and U3495 (N_3495,N_2585,N_1853);
xor U3496 (N_3496,N_2372,N_1083);
or U3497 (N_3497,N_1302,N_1473);
xnor U3498 (N_3498,N_1492,N_1989);
nor U3499 (N_3499,N_1995,N_860);
xor U3500 (N_3500,N_2396,N_1855);
nand U3501 (N_3501,N_2497,N_1160);
or U3502 (N_3502,N_1781,N_941);
nor U3503 (N_3503,N_1248,N_1530);
or U3504 (N_3504,N_657,N_1978);
nor U3505 (N_3505,N_2826,N_2133);
nor U3506 (N_3506,N_539,N_2541);
nand U3507 (N_3507,N_2367,N_2306);
or U3508 (N_3508,N_2841,N_2842);
and U3509 (N_3509,N_1233,N_1902);
nand U3510 (N_3510,N_1258,N_352);
xor U3511 (N_3511,N_172,N_2118);
or U3512 (N_3512,N_716,N_2837);
nand U3513 (N_3513,N_1064,N_2115);
xnor U3514 (N_3514,N_1756,N_2384);
nand U3515 (N_3515,N_1748,N_1552);
or U3516 (N_3516,N_1246,N_1007);
nor U3517 (N_3517,N_2752,N_2024);
xor U3518 (N_3518,N_1193,N_1640);
and U3519 (N_3519,N_541,N_785);
nand U3520 (N_3520,N_1357,N_2142);
nor U3521 (N_3521,N_386,N_2817);
or U3522 (N_3522,N_1633,N_1488);
xnor U3523 (N_3523,N_955,N_2494);
and U3524 (N_3524,N_94,N_494);
and U3525 (N_3525,N_1519,N_1318);
or U3526 (N_3526,N_253,N_837);
and U3527 (N_3527,N_220,N_1752);
nand U3528 (N_3528,N_254,N_160);
nor U3529 (N_3529,N_1423,N_520);
nand U3530 (N_3530,N_421,N_1996);
nor U3531 (N_3531,N_2326,N_443);
nor U3532 (N_3532,N_2534,N_550);
or U3533 (N_3533,N_1880,N_1316);
nand U3534 (N_3534,N_1417,N_2050);
and U3535 (N_3535,N_2607,N_965);
and U3536 (N_3536,N_342,N_2366);
xnor U3537 (N_3537,N_2297,N_2015);
nand U3538 (N_3538,N_2968,N_663);
or U3539 (N_3539,N_2492,N_2005);
xor U3540 (N_3540,N_2256,N_1705);
nand U3541 (N_3541,N_1458,N_656);
and U3542 (N_3542,N_90,N_409);
xnor U3543 (N_3543,N_1154,N_2446);
nor U3544 (N_3544,N_1717,N_993);
nand U3545 (N_3545,N_1173,N_1860);
and U3546 (N_3546,N_748,N_2137);
nand U3547 (N_3547,N_640,N_778);
xnor U3548 (N_3548,N_86,N_1146);
xor U3549 (N_3549,N_2540,N_2670);
nand U3550 (N_3550,N_757,N_405);
and U3551 (N_3551,N_1282,N_1157);
and U3552 (N_3552,N_1762,N_1138);
and U3553 (N_3553,N_345,N_355);
nor U3554 (N_3554,N_168,N_79);
nand U3555 (N_3555,N_31,N_1788);
and U3556 (N_3556,N_674,N_171);
or U3557 (N_3557,N_1801,N_1516);
xor U3558 (N_3558,N_448,N_936);
nor U3559 (N_3559,N_1397,N_689);
or U3560 (N_3560,N_1303,N_536);
or U3561 (N_3561,N_1021,N_2729);
nor U3562 (N_3562,N_2597,N_493);
xor U3563 (N_3563,N_762,N_1388);
and U3564 (N_3564,N_2620,N_1060);
or U3565 (N_3565,N_2159,N_2291);
nand U3566 (N_3566,N_1479,N_588);
and U3567 (N_3567,N_1586,N_2596);
xnor U3568 (N_3568,N_1273,N_2341);
or U3569 (N_3569,N_441,N_261);
xnor U3570 (N_3570,N_2570,N_1947);
or U3571 (N_3571,N_1499,N_2223);
nor U3572 (N_3572,N_42,N_2815);
and U3573 (N_3573,N_1189,N_2858);
and U3574 (N_3574,N_2249,N_2132);
nand U3575 (N_3575,N_2683,N_752);
and U3576 (N_3576,N_2345,N_1170);
nor U3577 (N_3577,N_1757,N_2955);
nand U3578 (N_3578,N_2767,N_709);
or U3579 (N_3579,N_1780,N_549);
and U3580 (N_3580,N_504,N_624);
and U3581 (N_3581,N_46,N_434);
or U3582 (N_3582,N_662,N_2787);
xnor U3583 (N_3583,N_592,N_1527);
and U3584 (N_3584,N_1418,N_208);
and U3585 (N_3585,N_2453,N_2839);
or U3586 (N_3586,N_1687,N_1637);
and U3587 (N_3587,N_575,N_869);
and U3588 (N_3588,N_2654,N_789);
or U3589 (N_3589,N_2348,N_2586);
and U3590 (N_3590,N_478,N_823);
and U3591 (N_3591,N_659,N_2090);
nor U3592 (N_3592,N_1105,N_2152);
xor U3593 (N_3593,N_1609,N_1502);
and U3594 (N_3594,N_1226,N_298);
and U3595 (N_3595,N_133,N_817);
nor U3596 (N_3596,N_1648,N_2245);
nand U3597 (N_3597,N_2940,N_1668);
or U3598 (N_3598,N_1072,N_140);
nand U3599 (N_3599,N_2835,N_2714);
nand U3600 (N_3600,N_2943,N_2517);
or U3601 (N_3601,N_699,N_1281);
and U3602 (N_3602,N_1133,N_2643);
or U3603 (N_3603,N_2548,N_767);
or U3604 (N_3604,N_1821,N_144);
and U3605 (N_3605,N_969,N_2209);
nor U3606 (N_3606,N_87,N_2080);
nand U3607 (N_3607,N_1823,N_798);
nor U3608 (N_3608,N_1444,N_307);
nand U3609 (N_3609,N_2822,N_1228);
nor U3610 (N_3610,N_874,N_1184);
xor U3611 (N_3611,N_186,N_2);
nor U3612 (N_3612,N_2308,N_2677);
nand U3613 (N_3613,N_123,N_1734);
nor U3614 (N_3614,N_1360,N_1896);
nand U3615 (N_3615,N_1750,N_927);
and U3616 (N_3616,N_547,N_811);
nor U3617 (N_3617,N_594,N_472);
and U3618 (N_3618,N_2613,N_2624);
or U3619 (N_3619,N_2006,N_1859);
xnor U3620 (N_3620,N_2110,N_2551);
and U3621 (N_3621,N_746,N_617);
xor U3622 (N_3622,N_1924,N_2259);
xor U3623 (N_3623,N_2923,N_806);
or U3624 (N_3624,N_749,N_143);
and U3625 (N_3625,N_2012,N_1237);
nor U3626 (N_3626,N_2258,N_103);
xor U3627 (N_3627,N_2700,N_2379);
xnor U3628 (N_3628,N_791,N_1451);
nor U3629 (N_3629,N_2425,N_2026);
nor U3630 (N_3630,N_1373,N_792);
and U3631 (N_3631,N_1783,N_2278);
nand U3632 (N_3632,N_1141,N_701);
xnor U3633 (N_3633,N_1298,N_1486);
or U3634 (N_3634,N_2515,N_2244);
and U3635 (N_3635,N_1845,N_2699);
nand U3636 (N_3636,N_2909,N_1759);
xor U3637 (N_3637,N_688,N_2014);
and U3638 (N_3638,N_1501,N_119);
nand U3639 (N_3639,N_1431,N_1554);
and U3640 (N_3640,N_2222,N_256);
xor U3641 (N_3641,N_437,N_2649);
or U3642 (N_3642,N_209,N_2993);
nand U3643 (N_3643,N_323,N_2623);
nor U3644 (N_3644,N_61,N_2705);
and U3645 (N_3645,N_1227,N_574);
xnor U3646 (N_3646,N_2774,N_1960);
xnor U3647 (N_3647,N_1030,N_67);
xnor U3648 (N_3648,N_226,N_2937);
and U3649 (N_3649,N_1454,N_2724);
and U3650 (N_3650,N_41,N_2565);
nor U3651 (N_3651,N_1327,N_923);
and U3652 (N_3652,N_1415,N_313);
nor U3653 (N_3653,N_1383,N_1450);
or U3654 (N_3654,N_1786,N_429);
and U3655 (N_3655,N_432,N_1771);
nand U3656 (N_3656,N_844,N_243);
nor U3657 (N_3657,N_579,N_1029);
nor U3658 (N_3658,N_48,N_2472);
and U3659 (N_3659,N_1404,N_297);
or U3660 (N_3660,N_360,N_2459);
and U3661 (N_3661,N_1090,N_1916);
and U3662 (N_3662,N_75,N_394);
or U3663 (N_3663,N_1650,N_1037);
nor U3664 (N_3664,N_695,N_555);
xor U3665 (N_3665,N_887,N_2615);
xnor U3666 (N_3666,N_780,N_2694);
and U3667 (N_3667,N_1882,N_161);
and U3668 (N_3668,N_151,N_1221);
nand U3669 (N_3669,N_1573,N_2122);
xor U3670 (N_3670,N_1047,N_1205);
xor U3671 (N_3671,N_529,N_1065);
nor U3672 (N_3672,N_2435,N_551);
nor U3673 (N_3673,N_1009,N_2200);
or U3674 (N_3674,N_1536,N_1854);
nand U3675 (N_3675,N_1891,N_2491);
and U3676 (N_3676,N_106,N_2276);
or U3677 (N_3677,N_1976,N_131);
nand U3678 (N_3678,N_193,N_2640);
and U3679 (N_3679,N_324,N_2231);
or U3680 (N_3680,N_591,N_1652);
nand U3681 (N_3681,N_49,N_597);
and U3682 (N_3682,N_1779,N_2444);
nor U3683 (N_3683,N_2380,N_476);
xnor U3684 (N_3684,N_1741,N_2480);
or U3685 (N_3685,N_621,N_2921);
xor U3686 (N_3686,N_2383,N_1522);
xnor U3687 (N_3687,N_836,N_742);
or U3688 (N_3688,N_2070,N_856);
nand U3689 (N_3689,N_1010,N_1056);
or U3690 (N_3690,N_980,N_1545);
or U3691 (N_3691,N_1886,N_2266);
nand U3692 (N_3692,N_6,N_932);
nor U3693 (N_3693,N_2035,N_387);
xor U3694 (N_3694,N_170,N_2240);
nor U3695 (N_3695,N_931,N_1956);
and U3696 (N_3696,N_1362,N_68);
and U3697 (N_3697,N_382,N_2648);
and U3698 (N_3698,N_2447,N_2241);
nand U3699 (N_3699,N_1600,N_2317);
and U3700 (N_3700,N_2156,N_868);
nor U3701 (N_3701,N_1059,N_1883);
and U3702 (N_3702,N_2641,N_1611);
and U3703 (N_3703,N_1948,N_296);
or U3704 (N_3704,N_24,N_1649);
and U3705 (N_3705,N_1528,N_2904);
and U3706 (N_3706,N_884,N_2864);
nand U3707 (N_3707,N_2434,N_896);
nand U3708 (N_3708,N_1368,N_1219);
nor U3709 (N_3709,N_1700,N_1939);
nand U3710 (N_3710,N_158,N_821);
and U3711 (N_3711,N_548,N_997);
nand U3712 (N_3712,N_1926,N_947);
and U3713 (N_3713,N_1986,N_1744);
xor U3714 (N_3714,N_2164,N_415);
nand U3715 (N_3715,N_620,N_2284);
and U3716 (N_3716,N_691,N_1251);
and U3717 (N_3717,N_37,N_1643);
xnor U3718 (N_3718,N_667,N_502);
nor U3719 (N_3719,N_1225,N_364);
and U3720 (N_3720,N_1358,N_1874);
xor U3721 (N_3721,N_2311,N_815);
or U3722 (N_3722,N_2020,N_2625);
xnor U3723 (N_3723,N_167,N_2696);
xor U3724 (N_3724,N_30,N_2985);
nand U3725 (N_3725,N_413,N_1615);
xnor U3726 (N_3726,N_1349,N_619);
and U3727 (N_3727,N_500,N_2672);
xor U3728 (N_3728,N_2094,N_1135);
nor U3729 (N_3729,N_404,N_1405);
nand U3730 (N_3730,N_918,N_1118);
nand U3731 (N_3731,N_2481,N_1802);
or U3732 (N_3732,N_1626,N_719);
or U3733 (N_3733,N_708,N_1525);
or U3734 (N_3734,N_745,N_1564);
xor U3735 (N_3735,N_2583,N_1242);
nor U3736 (N_3736,N_2392,N_73);
and U3737 (N_3737,N_1220,N_2373);
and U3738 (N_3738,N_2301,N_1437);
nand U3739 (N_3739,N_854,N_2405);
or U3740 (N_3740,N_2664,N_1673);
nor U3741 (N_3741,N_2911,N_765);
xor U3742 (N_3742,N_1810,N_2935);
nand U3743 (N_3743,N_1727,N_917);
and U3744 (N_3744,N_2702,N_1595);
and U3745 (N_3745,N_1731,N_2023);
nand U3746 (N_3746,N_1166,N_2033);
xnor U3747 (N_3747,N_642,N_888);
and U3748 (N_3748,N_2439,N_66);
or U3749 (N_3749,N_2823,N_1124);
nand U3750 (N_3750,N_913,N_654);
nand U3751 (N_3751,N_2635,N_2349);
xnor U3752 (N_3752,N_2113,N_1149);
nor U3753 (N_3753,N_389,N_215);
or U3754 (N_3754,N_2052,N_2612);
nor U3755 (N_3755,N_1773,N_294);
xnor U3756 (N_3756,N_1354,N_1470);
xor U3757 (N_3757,N_2578,N_2105);
and U3758 (N_3758,N_1646,N_1245);
nand U3759 (N_3759,N_2715,N_2069);
or U3760 (N_3760,N_1378,N_622);
and U3761 (N_3761,N_248,N_544);
nand U3762 (N_3762,N_252,N_2994);
nand U3763 (N_3763,N_1541,N_2004);
nand U3764 (N_3764,N_1684,N_1204);
and U3765 (N_3765,N_2060,N_2463);
nand U3766 (N_3766,N_2131,N_2333);
nor U3767 (N_3767,N_799,N_1568);
nor U3768 (N_3768,N_1355,N_2370);
nor U3769 (N_3769,N_0,N_2450);
or U3770 (N_3770,N_863,N_1508);
or U3771 (N_3771,N_595,N_1352);
nor U3772 (N_3772,N_174,N_203);
or U3773 (N_3773,N_2018,N_1922);
or U3774 (N_3774,N_1531,N_1745);
or U3775 (N_3775,N_680,N_80);
nand U3776 (N_3776,N_2860,N_615);
nand U3777 (N_3777,N_2829,N_392);
nand U3778 (N_3778,N_2125,N_2165);
nor U3779 (N_3779,N_2458,N_1370);
nor U3780 (N_3780,N_756,N_897);
and U3781 (N_3781,N_915,N_1384);
and U3782 (N_3782,N_2124,N_623);
and U3783 (N_3783,N_2591,N_1261);
and U3784 (N_3784,N_1787,N_1572);
or U3785 (N_3785,N_1256,N_375);
nor U3786 (N_3786,N_2042,N_1766);
nor U3787 (N_3787,N_1867,N_949);
and U3788 (N_3788,N_963,N_122);
xnor U3789 (N_3789,N_1975,N_223);
and U3790 (N_3790,N_295,N_2568);
xnor U3791 (N_3791,N_198,N_2645);
nand U3792 (N_3792,N_2577,N_2734);
nand U3793 (N_3793,N_2601,N_2429);
nand U3794 (N_3794,N_2972,N_630);
nor U3795 (N_3795,N_2975,N_395);
nor U3796 (N_3796,N_2422,N_2584);
or U3797 (N_3797,N_238,N_1278);
or U3798 (N_3798,N_1919,N_2356);
or U3799 (N_3799,N_524,N_239);
nor U3800 (N_3800,N_2808,N_107);
xor U3801 (N_3801,N_800,N_1098);
xor U3802 (N_3802,N_959,N_2644);
nor U3803 (N_3803,N_1915,N_57);
and U3804 (N_3804,N_871,N_996);
nand U3805 (N_3805,N_1421,N_235);
nor U3806 (N_3806,N_1453,N_1091);
xnor U3807 (N_3807,N_2288,N_2681);
nor U3808 (N_3808,N_2669,N_570);
nor U3809 (N_3809,N_1562,N_290);
and U3810 (N_3810,N_1179,N_2474);
or U3811 (N_3811,N_1268,N_2289);
nand U3812 (N_3812,N_2661,N_866);
and U3813 (N_3813,N_1016,N_2535);
nor U3814 (N_3814,N_1911,N_269);
and U3815 (N_3815,N_833,N_2243);
nand U3816 (N_3816,N_1968,N_1257);
nor U3817 (N_3817,N_763,N_1547);
and U3818 (N_3818,N_1725,N_2470);
nor U3819 (N_3819,N_2812,N_2720);
xor U3820 (N_3820,N_1440,N_2387);
and U3821 (N_3821,N_987,N_124);
nand U3822 (N_3822,N_232,N_766);
xnor U3823 (N_3823,N_304,N_1201);
and U3824 (N_3824,N_277,N_2684);
and U3825 (N_3825,N_338,N_565);
or U3826 (N_3826,N_723,N_2355);
nor U3827 (N_3827,N_210,N_1737);
or U3828 (N_3828,N_251,N_2789);
nor U3829 (N_3829,N_1321,N_1113);
or U3830 (N_3830,N_2814,N_2336);
nand U3831 (N_3831,N_1973,N_1703);
or U3832 (N_3832,N_891,N_2343);
and U3833 (N_3833,N_2072,N_59);
nor U3834 (N_3834,N_2321,N_69);
nand U3835 (N_3835,N_2233,N_459);
nor U3836 (N_3836,N_769,N_1495);
or U3837 (N_3837,N_2604,N_2188);
nand U3838 (N_3838,N_638,N_1814);
or U3839 (N_3839,N_484,N_2178);
or U3840 (N_3840,N_1999,N_2868);
nor U3841 (N_3841,N_1642,N_2801);
xnor U3842 (N_3842,N_1087,N_2338);
nor U3843 (N_3843,N_1982,N_2265);
and U3844 (N_3844,N_1308,N_225);
xor U3845 (N_3845,N_1051,N_2931);
nand U3846 (N_3846,N_1533,N_1002);
nor U3847 (N_3847,N_2707,N_191);
xnor U3848 (N_3848,N_1222,N_602);
nor U3849 (N_3849,N_2579,N_2016);
or U3850 (N_3850,N_2257,N_2573);
and U3851 (N_3851,N_2726,N_830);
nor U3852 (N_3852,N_1830,N_2441);
or U3853 (N_3853,N_2411,N_2058);
and U3854 (N_3854,N_1270,N_1964);
nand U3855 (N_3855,N_2221,N_1988);
nand U3856 (N_3856,N_1561,N_1714);
nand U3857 (N_3857,N_396,N_853);
xor U3858 (N_3858,N_1918,N_1760);
nor U3859 (N_3859,N_2203,N_1754);
xor U3860 (N_3860,N_21,N_2905);
nor U3861 (N_3861,N_1660,N_2437);
or U3862 (N_3862,N_2718,N_2704);
nand U3863 (N_3863,N_661,N_308);
xor U3864 (N_3864,N_1028,N_2682);
nor U3865 (N_3865,N_322,N_1244);
or U3866 (N_3866,N_797,N_2913);
xnor U3867 (N_3867,N_388,N_283);
xor U3868 (N_3868,N_774,N_956);
nand U3869 (N_3869,N_2486,N_1776);
or U3870 (N_3870,N_2756,N_52);
nor U3871 (N_3871,N_1462,N_2616);
nor U3872 (N_3872,N_1709,N_2538);
nand U3873 (N_3873,N_2542,N_776);
nand U3874 (N_3874,N_2101,N_2141);
and U3875 (N_3875,N_665,N_1088);
or U3876 (N_3876,N_2698,N_1785);
nand U3877 (N_3877,N_1456,N_2208);
nor U3878 (N_3878,N_77,N_2467);
or U3879 (N_3879,N_452,N_1070);
xor U3880 (N_3880,N_2627,N_423);
nand U3881 (N_3881,N_2402,N_1050);
and U3882 (N_3882,N_958,N_1930);
xnor U3883 (N_3883,N_1632,N_246);
nor U3884 (N_3884,N_1875,N_1159);
and U3885 (N_3885,N_330,N_2946);
xnor U3886 (N_3886,N_542,N_1540);
or U3887 (N_3887,N_1480,N_2523);
xor U3888 (N_3888,N_197,N_2469);
nand U3889 (N_3889,N_257,N_121);
and U3890 (N_3890,N_2314,N_2757);
nand U3891 (N_3891,N_2335,N_687);
and U3892 (N_3892,N_1122,N_1506);
nor U3893 (N_3893,N_1829,N_23);
or U3894 (N_3894,N_1758,N_2712);
and U3895 (N_3895,N_1005,N_2184);
or U3896 (N_3896,N_2769,N_1425);
and U3897 (N_3897,N_986,N_272);
and U3898 (N_3898,N_1401,N_118);
nand U3899 (N_3899,N_2202,N_1475);
xnor U3900 (N_3900,N_858,N_2513);
nor U3901 (N_3901,N_2168,N_2610);
nand U3902 (N_3902,N_2761,N_2827);
xnor U3903 (N_3903,N_1619,N_2479);
and U3904 (N_3904,N_1653,N_200);
xnor U3905 (N_3905,N_2040,N_1765);
nand U3906 (N_3906,N_2979,N_1150);
and U3907 (N_3907,N_2433,N_1658);
nand U3908 (N_3908,N_1076,N_2848);
nor U3909 (N_3909,N_816,N_1688);
or U3910 (N_3910,N_1241,N_2143);
nor U3911 (N_3911,N_2516,N_862);
or U3912 (N_3912,N_1962,N_729);
and U3913 (N_3913,N_22,N_1081);
or U3914 (N_3914,N_1945,N_867);
xor U3915 (N_3915,N_1027,N_318);
nand U3916 (N_3916,N_1887,N_2272);
and U3917 (N_3917,N_377,N_801);
or U3918 (N_3918,N_1180,N_2191);
nor U3919 (N_3919,N_1793,N_634);
and U3920 (N_3920,N_2008,N_2543);
nand U3921 (N_3921,N_1449,N_534);
nand U3922 (N_3922,N_664,N_1520);
or U3923 (N_3923,N_1933,N_2280);
nor U3924 (N_3924,N_1364,N_2001);
or U3925 (N_3925,N_1025,N_1304);
xnor U3926 (N_3926,N_2334,N_2127);
and U3927 (N_3927,N_1689,N_1372);
nand U3928 (N_3928,N_2987,N_562);
xnor U3929 (N_3929,N_2161,N_1551);
nand U3930 (N_3930,N_15,N_946);
nand U3931 (N_3931,N_2907,N_406);
nor U3932 (N_3932,N_2075,N_1274);
and U3933 (N_3933,N_1478,N_1822);
nor U3934 (N_3934,N_306,N_741);
or U3935 (N_3935,N_1172,N_1305);
and U3936 (N_3936,N_521,N_299);
or U3937 (N_3937,N_1628,N_1812);
nand U3938 (N_3938,N_1500,N_1359);
or U3939 (N_3939,N_2368,N_2327);
nor U3940 (N_3940,N_2507,N_2803);
or U3941 (N_3941,N_43,N_794);
nor U3942 (N_3942,N_1820,N_507);
nor U3943 (N_3943,N_305,N_2831);
nand U3944 (N_3944,N_1380,N_2582);
nand U3945 (N_3945,N_2510,N_2621);
and U3946 (N_3946,N_2659,N_1123);
or U3947 (N_3947,N_2667,N_2897);
and U3948 (N_3948,N_2772,N_475);
nand U3949 (N_3949,N_2354,N_2751);
nor U3950 (N_3950,N_1510,N_2413);
nor U3951 (N_3951,N_1957,N_1954);
xor U3952 (N_3952,N_2309,N_398);
or U3953 (N_3953,N_2187,N_2646);
and U3954 (N_3954,N_1216,N_2353);
nor U3955 (N_3955,N_35,N_954);
nor U3956 (N_3956,N_952,N_981);
nand U3957 (N_3957,N_1507,N_2922);
nand U3958 (N_3958,N_381,N_1080);
and U3959 (N_3959,N_2614,N_1240);
or U3960 (N_3960,N_2746,N_904);
xor U3961 (N_3961,N_1377,N_374);
nor U3962 (N_3962,N_1587,N_920);
xor U3963 (N_3963,N_1548,N_346);
or U3964 (N_3964,N_2217,N_2430);
xnor U3965 (N_3965,N_2996,N_628);
or U3966 (N_3966,N_852,N_426);
or U3967 (N_3967,N_2989,N_2766);
nand U3968 (N_3968,N_1330,N_468);
nor U3969 (N_3969,N_286,N_1363);
nand U3970 (N_3970,N_2862,N_2556);
or U3971 (N_3971,N_2890,N_2906);
nor U3972 (N_3972,N_2207,N_2009);
xnor U3973 (N_3973,N_135,N_2100);
and U3974 (N_3974,N_102,N_1504);
nand U3975 (N_3975,N_1465,N_2914);
or U3976 (N_3976,N_2250,N_2246);
nor U3977 (N_3977,N_2877,N_303);
xnor U3978 (N_3978,N_97,N_1739);
nand U3979 (N_3979,N_1877,N_2697);
nor U3980 (N_3980,N_2269,N_2022);
xnor U3981 (N_3981,N_60,N_626);
nor U3982 (N_3982,N_2783,N_1769);
or U3983 (N_3983,N_943,N_906);
xnor U3984 (N_3984,N_751,N_2262);
and U3985 (N_3985,N_1539,N_907);
xnor U3986 (N_3986,N_684,N_715);
xor U3987 (N_3987,N_805,N_416);
nand U3988 (N_3988,N_2832,N_2630);
or U3989 (N_3989,N_1371,N_506);
or U3990 (N_3990,N_967,N_2961);
or U3991 (N_3991,N_974,N_2663);
and U3992 (N_3992,N_2571,N_2908);
or U3993 (N_3993,N_480,N_205);
nor U3994 (N_3994,N_1284,N_1721);
nand U3995 (N_3995,N_2206,N_1001);
or U3996 (N_3996,N_2210,N_2748);
nand U3997 (N_3997,N_273,N_1917);
nor U3998 (N_3998,N_1057,N_1129);
and U3999 (N_3999,N_2391,N_914);
or U4000 (N_4000,N_735,N_1602);
nand U4001 (N_4001,N_1015,N_1341);
xor U4002 (N_4002,N_1967,N_2525);
nand U4003 (N_4003,N_1778,N_2950);
and U4004 (N_4004,N_1583,N_2631);
nand U4005 (N_4005,N_864,N_1385);
nor U4006 (N_4006,N_1441,N_966);
xnor U4007 (N_4007,N_479,N_1295);
and U4008 (N_4008,N_2511,N_1206);
xnor U4009 (N_4009,N_2153,N_2197);
and U4010 (N_4010,N_1983,N_1187);
nor U4011 (N_4011,N_422,N_1590);
or U4012 (N_4012,N_2408,N_368);
nor U4013 (N_4013,N_2797,N_2973);
nand U4014 (N_4014,N_2933,N_1366);
and U4015 (N_4015,N_1252,N_173);
nor U4016 (N_4016,N_1287,N_870);
nand U4017 (N_4017,N_690,N_2798);
nand U4018 (N_4018,N_2851,N_1265);
and U4019 (N_4019,N_1592,N_449);
or U4020 (N_4020,N_1971,N_2493);
and U4021 (N_4021,N_28,N_2747);
and U4022 (N_4022,N_1411,N_1542);
nand U4023 (N_4023,N_367,N_2949);
nand U4024 (N_4024,N_2884,N_440);
xnor U4025 (N_4025,N_89,N_783);
or U4026 (N_4026,N_698,N_2031);
nor U4027 (N_4027,N_1931,N_495);
xor U4028 (N_4028,N_1231,N_793);
nor U4029 (N_4029,N_1432,N_2201);
or U4030 (N_4030,N_175,N_166);
and U4031 (N_4031,N_408,N_972);
nor U4032 (N_4032,N_163,N_2056);
nand U4033 (N_4033,N_425,N_1044);
or U4034 (N_4034,N_1581,N_281);
and U4035 (N_4035,N_2028,N_1018);
xnor U4036 (N_4036,N_2347,N_1807);
xnor U4037 (N_4037,N_587,N_522);
nor U4038 (N_4038,N_1518,N_2322);
xor U4039 (N_4039,N_1695,N_2121);
or U4040 (N_4040,N_2626,N_560);
xor U4041 (N_4041,N_111,N_1839);
nor U4042 (N_4042,N_1605,N_1162);
nand U4043 (N_4043,N_393,N_2589);
or U4044 (N_4044,N_1936,N_753);
or U4045 (N_4045,N_957,N_2119);
and U4046 (N_4046,N_930,N_1672);
nor U4047 (N_4047,N_1426,N_53);
nand U4048 (N_4048,N_481,N_34);
nor U4049 (N_4049,N_390,N_1899);
and U4050 (N_4050,N_491,N_2986);
nand U4051 (N_4051,N_1742,N_2816);
nor U4052 (N_4052,N_845,N_2473);
or U4053 (N_4053,N_1597,N_825);
and U4054 (N_4054,N_1621,N_2969);
xor U4055 (N_4055,N_2599,N_2225);
and U4056 (N_4056,N_1409,N_686);
nor U4057 (N_4057,N_2419,N_2117);
nor U4058 (N_4058,N_2898,N_2743);
xnor U4059 (N_4059,N_683,N_1194);
xor U4060 (N_4060,N_2741,N_886);
and U4061 (N_4061,N_1210,N_2828);
nand U4062 (N_4062,N_372,N_532);
or U4063 (N_4063,N_672,N_1497);
and U4064 (N_4064,N_2000,N_2605);
xnor U4065 (N_4065,N_2760,N_1137);
xor U4066 (N_4066,N_2066,N_922);
xnor U4067 (N_4067,N_2983,N_1865);
and U4068 (N_4068,N_528,N_2503);
nor U4069 (N_4069,N_1053,N_583);
nand U4070 (N_4070,N_1176,N_1661);
nor U4071 (N_4071,N_2619,N_2800);
nand U4072 (N_4072,N_2559,N_1077);
and U4073 (N_4073,N_2062,N_1466);
and U4074 (N_4074,N_497,N_1041);
nor U4075 (N_4075,N_938,N_2719);
and U4076 (N_4076,N_681,N_2825);
nor U4077 (N_4077,N_1286,N_632);
xnor U4078 (N_4078,N_879,N_984);
xnor U4079 (N_4079,N_2786,N_36);
or U4080 (N_4080,N_831,N_2261);
or U4081 (N_4081,N_55,N_2737);
and U4082 (N_4082,N_379,N_370);
nand U4083 (N_4083,N_325,N_267);
and U4084 (N_4084,N_228,N_1972);
nand U4085 (N_4085,N_1262,N_1209);
and U4086 (N_4086,N_2755,N_2157);
nand U4087 (N_4087,N_951,N_2237);
and U4088 (N_4088,N_916,N_1856);
or U4089 (N_4089,N_2423,N_1768);
nor U4090 (N_4090,N_2777,N_508);
xnor U4091 (N_4091,N_1276,N_2561);
nand U4092 (N_4092,N_2834,N_112);
xnor U4093 (N_4093,N_2930,N_351);
xnor U4094 (N_4094,N_2328,N_2678);
and U4095 (N_4095,N_569,N_2508);
nor U4096 (N_4096,N_2903,N_221);
xnor U4097 (N_4097,N_702,N_726);
nand U4098 (N_4098,N_2506,N_1851);
xnor U4099 (N_4099,N_2861,N_99);
nand U4100 (N_4100,N_669,N_1234);
nand U4101 (N_4101,N_438,N_1101);
nand U4102 (N_4102,N_125,N_2765);
xor U4103 (N_4103,N_2685,N_2606);
xor U4104 (N_4104,N_145,N_1903);
nor U4105 (N_4105,N_2204,N_883);
nor U4106 (N_4106,N_1614,N_1827);
nand U4107 (N_4107,N_190,N_2263);
xor U4108 (N_4108,N_2749,N_1277);
nor U4109 (N_4109,N_859,N_1654);
or U4110 (N_4110,N_1062,N_2163);
or U4111 (N_4111,N_2364,N_2866);
nor U4112 (N_4112,N_460,N_202);
xnor U4113 (N_4113,N_1991,N_758);
nor U4114 (N_4114,N_1477,N_648);
or U4115 (N_4115,N_1806,N_1571);
or U4116 (N_4116,N_1553,N_1977);
nand U4117 (N_4117,N_1674,N_1876);
nor U4118 (N_4118,N_2294,N_1249);
nor U4119 (N_4119,N_2144,N_455);
and U4120 (N_4120,N_1312,N_673);
and U4121 (N_4121,N_458,N_2099);
xor U4122 (N_4122,N_2498,N_2671);
and U4123 (N_4123,N_1585,N_760);
nand U4124 (N_4124,N_1848,N_2662);
nor U4125 (N_4125,N_545,N_807);
nand U4126 (N_4126,N_2598,N_400);
nor U4127 (N_4127,N_2708,N_1987);
or U4128 (N_4128,N_2304,N_44);
xor U4129 (N_4129,N_964,N_1538);
nor U4130 (N_4130,N_2754,N_461);
xnor U4131 (N_4131,N_2563,N_2063);
or U4132 (N_4132,N_885,N_496);
xnor U4133 (N_4133,N_1904,N_1119);
nor U4134 (N_4134,N_2185,N_424);
or U4135 (N_4135,N_453,N_1348);
nor U4136 (N_4136,N_1419,N_1347);
or U4137 (N_4137,N_2424,N_1718);
nor U4138 (N_4138,N_462,N_2778);
or U4139 (N_4139,N_2431,N_2790);
nor U4140 (N_4140,N_2232,N_1618);
or U4141 (N_4141,N_446,N_14);
xor U4142 (N_4142,N_1186,N_527);
nor U4143 (N_4143,N_568,N_2716);
xnor U4144 (N_4144,N_2653,N_503);
or U4145 (N_4145,N_2216,N_2723);
or U4146 (N_4146,N_1514,N_2891);
xor U4147 (N_4147,N_2869,N_609);
or U4148 (N_4148,N_2253,N_1844);
and U4149 (N_4149,N_2205,N_29);
nor U4150 (N_4150,N_1517,N_2224);
nand U4151 (N_4151,N_369,N_373);
or U4152 (N_4152,N_631,N_2239);
xnor U4153 (N_4153,N_340,N_1833);
or U4154 (N_4154,N_270,N_1979);
and U4155 (N_4155,N_2611,N_2013);
and U4156 (N_4156,N_2061,N_2123);
or U4157 (N_4157,N_2750,N_988);
xor U4158 (N_4158,N_2537,N_1082);
nor U4159 (N_4159,N_1914,N_1264);
nor U4160 (N_4160,N_2947,N_1722);
and U4161 (N_4161,N_671,N_2995);
or U4162 (N_4162,N_2896,N_2149);
nand U4163 (N_4163,N_2477,N_127);
nand U4164 (N_4164,N_1255,N_2549);
and U4165 (N_4165,N_810,N_2213);
nand U4166 (N_4166,N_2319,N_2484);
xor U4167 (N_4167,N_418,N_1706);
and U4168 (N_4168,N_1263,N_1512);
or U4169 (N_4169,N_1846,N_1838);
nand U4170 (N_4170,N_1905,N_721);
nor U4171 (N_4171,N_1588,N_2174);
nand U4172 (N_4172,N_944,N_585);
nor U4173 (N_4173,N_2865,N_2555);
xor U4174 (N_4174,N_2461,N_1043);
nor U4175 (N_4175,N_1107,N_1389);
nand U4176 (N_4176,N_1334,N_1909);
or U4177 (N_4177,N_1004,N_2691);
and U4178 (N_4178,N_546,N_561);
and U4179 (N_4179,N_658,N_165);
xnor U4180 (N_4180,N_1075,N_908);
and U4181 (N_4181,N_2074,N_1386);
nand U4182 (N_4182,N_1662,N_1808);
nor U4183 (N_4183,N_2475,N_2112);
nand U4184 (N_4184,N_2378,N_2466);
xnor U4185 (N_4185,N_1963,N_1900);
nand U4186 (N_4186,N_1534,N_2529);
xor U4187 (N_4187,N_1420,N_1115);
nor U4188 (N_4188,N_96,N_2087);
xor U4189 (N_4189,N_1794,N_2182);
or U4190 (N_4190,N_2680,N_2417);
nand U4191 (N_4191,N_953,N_533);
and U4192 (N_4192,N_2162,N_905);
xor U4193 (N_4193,N_1665,N_2496);
xor U4194 (N_4194,N_181,N_153);
xnor U4195 (N_4195,N_361,N_1148);
nand U4196 (N_4196,N_1307,N_1907);
nand U4197 (N_4197,N_2962,N_2768);
and U4198 (N_4198,N_1346,N_1816);
and U4199 (N_4199,N_1215,N_1034);
nor U4200 (N_4200,N_1620,N_2229);
nand U4201 (N_4201,N_2687,N_1457);
xnor U4202 (N_4202,N_2999,N_2665);
xor U4203 (N_4203,N_677,N_2982);
xnor U4204 (N_4204,N_1447,N_2390);
nand U4205 (N_4205,N_1729,N_2504);
xnor U4206 (N_4206,N_2002,N_1832);
nor U4207 (N_4207,N_1207,N_2553);
and U4208 (N_4208,N_514,N_1412);
nand U4209 (N_4209,N_1403,N_2780);
nor U4210 (N_4210,N_1301,N_2838);
nor U4211 (N_4211,N_1690,N_2941);
nor U4212 (N_4212,N_2344,N_2518);
or U4213 (N_4213,N_2145,N_1774);
and U4214 (N_4214,N_436,N_2811);
nand U4215 (N_4215,N_2629,N_2732);
nor U4216 (N_4216,N_926,N_2096);
and U4217 (N_4217,N_136,N_2676);
or U4218 (N_4218,N_4,N_204);
and U4219 (N_4219,N_808,N_1579);
nand U4220 (N_4220,N_2916,N_2944);
nor U4221 (N_4221,N_2528,N_13);
or U4222 (N_4222,N_523,N_1438);
xnor U4223 (N_4223,N_463,N_2019);
or U4224 (N_4224,N_105,N_2404);
xnor U4225 (N_4225,N_764,N_2195);
and U4226 (N_4226,N_192,N_625);
nand U4227 (N_4227,N_572,N_694);
nand U4228 (N_4228,N_1697,N_1487);
or U4229 (N_4229,N_2038,N_1864);
or U4230 (N_4230,N_1042,N_646);
and U4231 (N_4231,N_1439,N_2285);
xnor U4232 (N_4232,N_2091,N_1795);
nand U4233 (N_4233,N_925,N_1467);
xnor U4234 (N_4234,N_2717,N_2910);
nor U4235 (N_4235,N_2010,N_2166);
xor U4236 (N_4236,N_2863,N_2550);
and U4237 (N_4237,N_842,N_108);
nand U4238 (N_4238,N_1196,N_1279);
and U4239 (N_4239,N_442,N_1381);
xnor U4240 (N_4240,N_2171,N_2521);
nand U4241 (N_4241,N_2316,N_739);
nor U4242 (N_4242,N_530,N_809);
and U4243 (N_4243,N_383,N_1723);
or U4244 (N_4244,N_1740,N_1728);
xnor U4245 (N_4245,N_2956,N_2147);
nand U4246 (N_4246,N_2389,N_2880);
nand U4247 (N_4247,N_1067,N_2397);
xor U4248 (N_4248,N_2727,N_1297);
and U4249 (N_4249,N_1576,N_2773);
or U4250 (N_4250,N_1339,N_1313);
nand U4251 (N_4251,N_2882,N_1710);
xor U4252 (N_4252,N_1869,N_180);
xor U4253 (N_4253,N_2495,N_2138);
xor U4254 (N_4254,N_2298,N_477);
or U4255 (N_4255,N_1429,N_2709);
and U4256 (N_4256,N_1496,N_2873);
xor U4257 (N_4257,N_1033,N_2053);
xnor U4258 (N_4258,N_1819,N_829);
nor U4259 (N_4259,N_1594,N_1095);
xnor U4260 (N_4260,N_2436,N_1953);
and U4261 (N_4261,N_1664,N_1329);
and U4262 (N_4262,N_644,N_435);
nor U4263 (N_4263,N_365,N_945);
or U4264 (N_4264,N_1448,N_363);
or U4265 (N_4265,N_2312,N_839);
xnor U4266 (N_4266,N_1906,N_1336);
or U4267 (N_4267,N_333,N_2544);
xnor U4268 (N_4268,N_2642,N_1111);
xnor U4269 (N_4269,N_1026,N_45);
or U4270 (N_4270,N_1139,N_1202);
xnor U4271 (N_4271,N_581,N_2320);
and U4272 (N_4272,N_113,N_1761);
xor U4273 (N_4273,N_2457,N_1895);
nand U4274 (N_4274,N_556,N_2879);
nor U4275 (N_4275,N_747,N_1631);
xnor U4276 (N_4276,N_1681,N_2638);
xnor U4277 (N_4277,N_939,N_1350);
or U4278 (N_4278,N_81,N_1174);
or U4279 (N_4279,N_1178,N_2358);
and U4280 (N_4280,N_1884,N_335);
xnor U4281 (N_4281,N_975,N_903);
nand U4282 (N_4282,N_2802,N_1809);
nor U4283 (N_4283,N_1784,N_2029);
nand U4284 (N_4284,N_2959,N_2876);
nand U4285 (N_4285,N_1641,N_1985);
or U4286 (N_4286,N_855,N_1061);
nor U4287 (N_4287,N_1837,N_1921);
or U4288 (N_4288,N_1943,N_1980);
xor U4289 (N_4289,N_2804,N_2887);
and U4290 (N_4290,N_445,N_311);
nor U4291 (N_4291,N_777,N_19);
nor U4292 (N_4292,N_1910,N_485);
nor U4293 (N_4293,N_1720,N_2414);
xor U4294 (N_4294,N_275,N_2416);
nor U4295 (N_4295,N_70,N_1399);
nand U4296 (N_4296,N_2912,N_1309);
nor U4297 (N_4297,N_1393,N_2733);
and U4298 (N_4298,N_2305,N_91);
and U4299 (N_4299,N_2037,N_354);
nand U4300 (N_4300,N_1558,N_357);
nand U4301 (N_4301,N_894,N_1476);
nor U4302 (N_4302,N_341,N_2234);
nor U4303 (N_4303,N_1199,N_300);
nor U4304 (N_4304,N_2738,N_2673);
nand U4305 (N_4305,N_1161,N_1591);
or U4306 (N_4306,N_2440,N_110);
xor U4307 (N_4307,N_2893,N_2840);
or U4308 (N_4308,N_1691,N_328);
or U4309 (N_4309,N_2107,N_39);
nor U4310 (N_4310,N_2393,N_2781);
xnor U4311 (N_4311,N_2116,N_2270);
nand U4312 (N_4312,N_2065,N_262);
xor U4313 (N_4313,N_2632,N_1127);
nand U4314 (N_4314,N_38,N_2155);
nand U4315 (N_4315,N_1147,N_2106);
and U4316 (N_4316,N_1188,N_64);
or U4317 (N_4317,N_470,N_1578);
nand U4318 (N_4318,N_636,N_697);
xnor U4319 (N_4319,N_2843,N_2186);
and U4320 (N_4320,N_2964,N_577);
nand U4321 (N_4321,N_2919,N_1755);
nor U4322 (N_4322,N_2499,N_454);
xor U4323 (N_4323,N_2011,N_1260);
nand U4324 (N_4324,N_822,N_1490);
and U4325 (N_4325,N_2350,N_1603);
or U4326 (N_4326,N_1908,N_2713);
and U4327 (N_4327,N_1434,N_1049);
xnor U4328 (N_4328,N_713,N_343);
xnor U4329 (N_4329,N_1577,N_1326);
xnor U4330 (N_4330,N_2871,N_2603);
nand U4331 (N_4331,N_138,N_559);
nor U4332 (N_4332,N_490,N_1203);
xnor U4333 (N_4333,N_2810,N_1345);
and U4334 (N_4334,N_1791,N_1428);
and U4335 (N_4335,N_962,N_2647);
xnor U4336 (N_4336,N_2456,N_2928);
and U4337 (N_4337,N_1394,N_450);
or U4338 (N_4338,N_2403,N_1032);
and U4339 (N_4339,N_2974,N_2398);
or U4340 (N_4340,N_995,N_2443);
or U4341 (N_4341,N_2965,N_2785);
and U4342 (N_4342,N_1593,N_1328);
nor U4343 (N_4343,N_1647,N_518);
nand U4344 (N_4344,N_234,N_2169);
nand U4345 (N_4345,N_78,N_2784);
and U4346 (N_4346,N_1961,N_2228);
nand U4347 (N_4347,N_668,N_2976);
nand U4348 (N_4348,N_940,N_1310);
or U4349 (N_4349,N_1102,N_2779);
nor U4350 (N_4350,N_1815,N_2126);
xor U4351 (N_4351,N_2077,N_2236);
nor U4352 (N_4352,N_1055,N_2742);
or U4353 (N_4353,N_1598,N_2652);
and U4354 (N_4354,N_750,N_2179);
and U4355 (N_4355,N_1670,N_857);
xnor U4356 (N_4356,N_466,N_2085);
nor U4357 (N_4357,N_1142,N_26);
nand U4358 (N_4358,N_2158,N_18);
and U4359 (N_4359,N_2003,N_2189);
nor U4360 (N_4360,N_843,N_291);
nor U4361 (N_4361,N_2445,N_2580);
xor U4362 (N_4362,N_2932,N_1442);
xor U4363 (N_4363,N_1524,N_525);
xor U4364 (N_4364,N_1998,N_875);
and U4365 (N_4365,N_40,N_983);
and U4366 (N_4366,N_2198,N_2057);
xnor U4367 (N_4367,N_2679,N_482);
xor U4368 (N_4368,N_1455,N_25);
nor U4369 (N_4369,N_2689,N_2242);
xor U4370 (N_4370,N_1331,N_1031);
nand U4371 (N_4371,N_2214,N_292);
xnor U4372 (N_4372,N_2901,N_2047);
xnor U4373 (N_4373,N_928,N_2488);
nand U4374 (N_4374,N_2821,N_2400);
xnor U4375 (N_4375,N_600,N_207);
nor U4376 (N_4376,N_336,N_679);
and U4377 (N_4377,N_2273,N_1446);
nand U4378 (N_4378,N_1214,N_2092);
and U4379 (N_4379,N_74,N_1969);
nand U4380 (N_4380,N_2059,N_356);
nand U4381 (N_4381,N_1715,N_233);
and U4382 (N_4382,N_2120,N_901);
nor U4383 (N_4383,N_2566,N_1140);
or U4384 (N_4384,N_2703,N_910);
and U4385 (N_4385,N_1736,N_1223);
nor U4386 (N_4386,N_1616,N_419);
or U4387 (N_4387,N_846,N_2853);
xor U4388 (N_4388,N_1881,N_2701);
or U4389 (N_4389,N_1636,N_8);
nand U4390 (N_4390,N_678,N_1000);
nand U4391 (N_4391,N_1894,N_670);
nand U4392 (N_4392,N_876,N_2885);
nor U4393 (N_4393,N_1169,N_1433);
xor U4394 (N_4394,N_1582,N_2576);
and U4395 (N_4395,N_349,N_2286);
nand U4396 (N_4396,N_2552,N_2926);
and U4397 (N_4397,N_2211,N_2574);
xnor U4398 (N_4398,N_1817,N_2081);
or U4399 (N_4399,N_2407,N_693);
nand U4400 (N_4400,N_1071,N_1337);
xor U4401 (N_4401,N_1435,N_1693);
nor U4402 (N_4402,N_576,N_148);
xnor U4403 (N_4403,N_2536,N_612);
nand U4404 (N_4404,N_1719,N_33);
and U4405 (N_4405,N_738,N_2315);
xnor U4406 (N_4406,N_731,N_1698);
or U4407 (N_4407,N_1981,N_1103);
xor U4408 (N_4408,N_771,N_1340);
and U4409 (N_4409,N_824,N_1503);
nand U4410 (N_4410,N_1402,N_1003);
and U4411 (N_4411,N_2735,N_58);
and U4412 (N_4412,N_1560,N_320);
or U4413 (N_4413,N_2027,N_882);
and U4414 (N_4414,N_2359,N_1020);
and U4415 (N_4415,N_2248,N_961);
nor U4416 (N_4416,N_1613,N_2464);
and U4417 (N_4417,N_2036,N_1666);
nand U4418 (N_4418,N_2071,N_2634);
or U4419 (N_4419,N_1489,N_1414);
nor U4420 (N_4420,N_2485,N_85);
xor U4421 (N_4421,N_1156,N_155);
nor U4422 (N_4422,N_1413,N_614);
xnor U4423 (N_4423,N_2658,N_1606);
and U4424 (N_4424,N_1901,N_128);
xnor U4425 (N_4425,N_1944,N_1074);
nor U4426 (N_4426,N_2592,N_537);
or U4427 (N_4427,N_11,N_2953);
and U4428 (N_4428,N_704,N_1913);
nand U4429 (N_4429,N_2084,N_2505);
nand U4430 (N_4430,N_775,N_1888);
xnor U4431 (N_4431,N_727,N_247);
xnor U4432 (N_4432,N_162,N_1125);
and U4433 (N_4433,N_1685,N_2460);
nor U4434 (N_4434,N_1468,N_1570);
and U4435 (N_4435,N_2254,N_1574);
nand U4436 (N_4436,N_1134,N_62);
nor U4437 (N_4437,N_893,N_469);
or U4438 (N_4438,N_540,N_164);
xor U4439 (N_4439,N_838,N_2352);
xor U4440 (N_4440,N_1679,N_499);
nor U4441 (N_4441,N_2412,N_149);
xnor U4442 (N_4442,N_2686,N_2032);
and U4443 (N_4443,N_1236,N_141);
nor U4444 (N_4444,N_217,N_2856);
nand U4445 (N_4445,N_1319,N_820);
nor U4446 (N_4446,N_2763,N_711);
nand U4447 (N_4447,N_802,N_2794);
or U4448 (N_4448,N_902,N_32);
or U4449 (N_4449,N_116,N_2637);
nor U4450 (N_4450,N_1013,N_724);
or U4451 (N_4451,N_362,N_2089);
xnor U4452 (N_4452,N_1764,N_1763);
and U4453 (N_4453,N_1130,N_2530);
and U4454 (N_4454,N_1800,N_1505);
xnor U4455 (N_4455,N_371,N_399);
xor U4456 (N_4456,N_1376,N_1555);
nand U4457 (N_4457,N_584,N_1566);
nor U4458 (N_4458,N_812,N_2196);
and U4459 (N_4459,N_1167,N_2674);
nand U4460 (N_4460,N_2330,N_2482);
and U4461 (N_4461,N_878,N_2268);
nor U4462 (N_4462,N_3,N_1949);
nand U4463 (N_4463,N_1777,N_1120);
nand U4464 (N_4464,N_1569,N_743);
nand U4465 (N_4465,N_1686,N_1704);
nand U4466 (N_4466,N_2296,N_2824);
or U4467 (N_4467,N_725,N_2857);
nor U4468 (N_4468,N_1469,N_649);
or U4469 (N_4469,N_2438,N_1099);
nand U4470 (N_4470,N_2361,N_347);
nand U4471 (N_4471,N_214,N_101);
xor U4472 (N_4472,N_840,N_1474);
nor U4473 (N_4473,N_2706,N_1046);
or U4474 (N_4474,N_1097,N_276);
xnor U4475 (N_4475,N_1471,N_2522);
xor U4476 (N_4476,N_2728,N_796);
xor U4477 (N_4477,N_781,N_2849);
xnor U4478 (N_4478,N_1645,N_2199);
or U4479 (N_4479,N_2247,N_1068);
or U4480 (N_4480,N_54,N_2173);
xnor U4481 (N_4481,N_350,N_733);
nand U4482 (N_4482,N_639,N_804);
and U4483 (N_4483,N_1696,N_992);
nor U4484 (N_4484,N_1629,N_319);
nor U4485 (N_4485,N_1617,N_1143);
nand U4486 (N_4486,N_1599,N_2951);
or U4487 (N_4487,N_2883,N_1498);
xor U4488 (N_4488,N_641,N_1408);
or U4489 (N_4489,N_510,N_977);
nor U4490 (N_4490,N_1356,N_150);
or U4491 (N_4491,N_1934,N_1544);
nand U4492 (N_4492,N_2452,N_1254);
or U4493 (N_4493,N_222,N_120);
or U4494 (N_4494,N_2337,N_2086);
xnor U4495 (N_4495,N_889,N_2655);
xor U4496 (N_4496,N_2650,N_1494);
or U4497 (N_4497,N_301,N_2048);
nand U4498 (N_4498,N_2410,N_126);
nand U4499 (N_4499,N_464,N_718);
nor U4500 (N_4500,N_1365,N_2519);
nand U4501 (N_4501,N_1074,N_2475);
and U4502 (N_4502,N_2999,N_2760);
xnor U4503 (N_4503,N_1540,N_599);
or U4504 (N_4504,N_1708,N_1893);
and U4505 (N_4505,N_21,N_688);
nor U4506 (N_4506,N_2816,N_102);
nor U4507 (N_4507,N_379,N_2708);
and U4508 (N_4508,N_284,N_364);
nor U4509 (N_4509,N_909,N_269);
nand U4510 (N_4510,N_511,N_423);
xnor U4511 (N_4511,N_1250,N_847);
xnor U4512 (N_4512,N_791,N_1452);
nor U4513 (N_4513,N_1684,N_1402);
nor U4514 (N_4514,N_2402,N_2246);
xnor U4515 (N_4515,N_2014,N_925);
or U4516 (N_4516,N_203,N_535);
xnor U4517 (N_4517,N_2568,N_1395);
and U4518 (N_4518,N_2417,N_651);
or U4519 (N_4519,N_310,N_2880);
nand U4520 (N_4520,N_675,N_2643);
xnor U4521 (N_4521,N_2592,N_15);
and U4522 (N_4522,N_76,N_765);
or U4523 (N_4523,N_459,N_1744);
and U4524 (N_4524,N_2262,N_2402);
xnor U4525 (N_4525,N_1443,N_1841);
nand U4526 (N_4526,N_1850,N_876);
nor U4527 (N_4527,N_1373,N_1885);
nor U4528 (N_4528,N_1046,N_2609);
nand U4529 (N_4529,N_758,N_1755);
nor U4530 (N_4530,N_2099,N_2855);
and U4531 (N_4531,N_18,N_770);
nor U4532 (N_4532,N_2752,N_1010);
or U4533 (N_4533,N_2840,N_1245);
nand U4534 (N_4534,N_1650,N_277);
or U4535 (N_4535,N_1260,N_964);
and U4536 (N_4536,N_1237,N_2336);
and U4537 (N_4537,N_2615,N_23);
nand U4538 (N_4538,N_391,N_1540);
or U4539 (N_4539,N_239,N_2290);
or U4540 (N_4540,N_2761,N_2476);
nor U4541 (N_4541,N_1140,N_1907);
nand U4542 (N_4542,N_2545,N_2503);
nand U4543 (N_4543,N_1771,N_192);
and U4544 (N_4544,N_1557,N_1742);
or U4545 (N_4545,N_47,N_2990);
nand U4546 (N_4546,N_2119,N_1522);
or U4547 (N_4547,N_610,N_371);
nor U4548 (N_4548,N_2109,N_1260);
nand U4549 (N_4549,N_2090,N_98);
or U4550 (N_4550,N_2676,N_1762);
nand U4551 (N_4551,N_2456,N_2179);
and U4552 (N_4552,N_172,N_2403);
nor U4553 (N_4553,N_496,N_1970);
or U4554 (N_4554,N_1655,N_1865);
nand U4555 (N_4555,N_1779,N_2169);
xor U4556 (N_4556,N_687,N_785);
or U4557 (N_4557,N_1280,N_2128);
xor U4558 (N_4558,N_1705,N_692);
and U4559 (N_4559,N_930,N_1664);
and U4560 (N_4560,N_2261,N_2796);
xor U4561 (N_4561,N_496,N_898);
xnor U4562 (N_4562,N_428,N_963);
or U4563 (N_4563,N_1059,N_1029);
nand U4564 (N_4564,N_156,N_2612);
xor U4565 (N_4565,N_1857,N_2297);
or U4566 (N_4566,N_549,N_2073);
nand U4567 (N_4567,N_672,N_2055);
nor U4568 (N_4568,N_1260,N_2794);
nor U4569 (N_4569,N_2059,N_527);
nand U4570 (N_4570,N_39,N_2913);
nand U4571 (N_4571,N_1211,N_2569);
and U4572 (N_4572,N_580,N_2121);
xor U4573 (N_4573,N_158,N_437);
nor U4574 (N_4574,N_1125,N_1844);
and U4575 (N_4575,N_2494,N_2872);
or U4576 (N_4576,N_2996,N_2245);
nor U4577 (N_4577,N_1448,N_2528);
nand U4578 (N_4578,N_1843,N_35);
or U4579 (N_4579,N_77,N_2171);
and U4580 (N_4580,N_1919,N_2346);
xor U4581 (N_4581,N_2805,N_2895);
and U4582 (N_4582,N_1852,N_2765);
or U4583 (N_4583,N_2218,N_451);
nor U4584 (N_4584,N_2419,N_2030);
nand U4585 (N_4585,N_2615,N_2667);
nor U4586 (N_4586,N_2404,N_524);
xor U4587 (N_4587,N_2702,N_313);
and U4588 (N_4588,N_1092,N_1322);
and U4589 (N_4589,N_1477,N_483);
and U4590 (N_4590,N_318,N_1214);
nor U4591 (N_4591,N_1272,N_1147);
or U4592 (N_4592,N_2703,N_1689);
nand U4593 (N_4593,N_2825,N_710);
nor U4594 (N_4594,N_2456,N_1087);
and U4595 (N_4595,N_2958,N_2740);
nand U4596 (N_4596,N_1249,N_2008);
xor U4597 (N_4597,N_1201,N_446);
and U4598 (N_4598,N_2290,N_1812);
nand U4599 (N_4599,N_2829,N_2697);
and U4600 (N_4600,N_732,N_2822);
and U4601 (N_4601,N_294,N_1506);
nand U4602 (N_4602,N_2309,N_969);
and U4603 (N_4603,N_1299,N_2458);
xor U4604 (N_4604,N_2105,N_1020);
and U4605 (N_4605,N_2108,N_1250);
nor U4606 (N_4606,N_1040,N_878);
nand U4607 (N_4607,N_2554,N_136);
nor U4608 (N_4608,N_63,N_1475);
nand U4609 (N_4609,N_734,N_2791);
xor U4610 (N_4610,N_60,N_425);
nor U4611 (N_4611,N_1235,N_1574);
nand U4612 (N_4612,N_179,N_491);
nand U4613 (N_4613,N_2713,N_218);
nand U4614 (N_4614,N_2876,N_2069);
and U4615 (N_4615,N_1226,N_331);
nor U4616 (N_4616,N_595,N_870);
or U4617 (N_4617,N_1001,N_2977);
xnor U4618 (N_4618,N_890,N_1615);
xnor U4619 (N_4619,N_2524,N_275);
or U4620 (N_4620,N_418,N_147);
and U4621 (N_4621,N_212,N_2887);
nand U4622 (N_4622,N_2309,N_1644);
xor U4623 (N_4623,N_701,N_247);
and U4624 (N_4624,N_823,N_2624);
xnor U4625 (N_4625,N_1645,N_92);
nor U4626 (N_4626,N_66,N_1750);
nand U4627 (N_4627,N_2849,N_1721);
xnor U4628 (N_4628,N_256,N_1258);
or U4629 (N_4629,N_2876,N_2191);
xnor U4630 (N_4630,N_135,N_2045);
xor U4631 (N_4631,N_204,N_1315);
nor U4632 (N_4632,N_2641,N_1375);
nor U4633 (N_4633,N_1373,N_2624);
xor U4634 (N_4634,N_2690,N_2971);
nor U4635 (N_4635,N_1575,N_878);
xor U4636 (N_4636,N_2097,N_2944);
or U4637 (N_4637,N_1481,N_2299);
or U4638 (N_4638,N_1858,N_288);
or U4639 (N_4639,N_935,N_245);
xor U4640 (N_4640,N_1656,N_1464);
xnor U4641 (N_4641,N_742,N_2124);
nor U4642 (N_4642,N_1276,N_69);
nor U4643 (N_4643,N_2087,N_412);
nor U4644 (N_4644,N_2336,N_1876);
and U4645 (N_4645,N_2908,N_1766);
xnor U4646 (N_4646,N_2469,N_69);
nor U4647 (N_4647,N_1489,N_385);
and U4648 (N_4648,N_773,N_243);
and U4649 (N_4649,N_2748,N_1769);
xnor U4650 (N_4650,N_2173,N_2922);
or U4651 (N_4651,N_718,N_1796);
or U4652 (N_4652,N_1757,N_1229);
nand U4653 (N_4653,N_1467,N_248);
xor U4654 (N_4654,N_2681,N_536);
and U4655 (N_4655,N_18,N_2311);
nor U4656 (N_4656,N_1557,N_1921);
and U4657 (N_4657,N_832,N_2720);
nand U4658 (N_4658,N_1684,N_414);
and U4659 (N_4659,N_1443,N_2104);
xnor U4660 (N_4660,N_1546,N_2414);
nor U4661 (N_4661,N_2260,N_1817);
nor U4662 (N_4662,N_2298,N_58);
nand U4663 (N_4663,N_2543,N_1889);
or U4664 (N_4664,N_1468,N_1547);
nand U4665 (N_4665,N_1159,N_2999);
or U4666 (N_4666,N_2089,N_1088);
nor U4667 (N_4667,N_2367,N_1596);
and U4668 (N_4668,N_2851,N_781);
xnor U4669 (N_4669,N_539,N_1150);
nand U4670 (N_4670,N_1714,N_1180);
and U4671 (N_4671,N_835,N_617);
or U4672 (N_4672,N_2362,N_1202);
nor U4673 (N_4673,N_1291,N_2559);
xnor U4674 (N_4674,N_596,N_2971);
and U4675 (N_4675,N_430,N_1295);
and U4676 (N_4676,N_1261,N_927);
and U4677 (N_4677,N_1307,N_2558);
nand U4678 (N_4678,N_1721,N_624);
nor U4679 (N_4679,N_2251,N_263);
nor U4680 (N_4680,N_2418,N_1767);
nand U4681 (N_4681,N_743,N_2830);
or U4682 (N_4682,N_575,N_532);
nor U4683 (N_4683,N_716,N_1149);
xnor U4684 (N_4684,N_2067,N_824);
nor U4685 (N_4685,N_685,N_797);
nand U4686 (N_4686,N_2965,N_2132);
nor U4687 (N_4687,N_1041,N_150);
or U4688 (N_4688,N_2798,N_2887);
or U4689 (N_4689,N_1960,N_1143);
or U4690 (N_4690,N_543,N_2747);
and U4691 (N_4691,N_392,N_2453);
xor U4692 (N_4692,N_2251,N_2121);
nand U4693 (N_4693,N_766,N_2908);
or U4694 (N_4694,N_2835,N_1498);
nor U4695 (N_4695,N_1518,N_834);
nor U4696 (N_4696,N_1182,N_2085);
nor U4697 (N_4697,N_1772,N_2491);
or U4698 (N_4698,N_348,N_49);
and U4699 (N_4699,N_309,N_282);
nand U4700 (N_4700,N_2928,N_2317);
nor U4701 (N_4701,N_2702,N_622);
xor U4702 (N_4702,N_1868,N_1298);
nor U4703 (N_4703,N_2426,N_163);
or U4704 (N_4704,N_1066,N_851);
or U4705 (N_4705,N_1238,N_1268);
xnor U4706 (N_4706,N_332,N_311);
and U4707 (N_4707,N_769,N_1455);
and U4708 (N_4708,N_637,N_1297);
and U4709 (N_4709,N_2295,N_1601);
and U4710 (N_4710,N_425,N_1912);
and U4711 (N_4711,N_2113,N_1397);
or U4712 (N_4712,N_542,N_2387);
and U4713 (N_4713,N_2828,N_58);
and U4714 (N_4714,N_1361,N_1383);
or U4715 (N_4715,N_2883,N_2148);
and U4716 (N_4716,N_397,N_2026);
and U4717 (N_4717,N_1852,N_2938);
nor U4718 (N_4718,N_486,N_1683);
nor U4719 (N_4719,N_1666,N_1453);
or U4720 (N_4720,N_347,N_2353);
nand U4721 (N_4721,N_2782,N_2534);
and U4722 (N_4722,N_861,N_1790);
nor U4723 (N_4723,N_1650,N_1076);
xnor U4724 (N_4724,N_1048,N_442);
xor U4725 (N_4725,N_2410,N_1094);
nor U4726 (N_4726,N_1603,N_2120);
xor U4727 (N_4727,N_165,N_841);
and U4728 (N_4728,N_2942,N_466);
and U4729 (N_4729,N_2765,N_805);
nand U4730 (N_4730,N_2842,N_1091);
xnor U4731 (N_4731,N_1720,N_1290);
or U4732 (N_4732,N_26,N_1091);
or U4733 (N_4733,N_1155,N_1339);
xor U4734 (N_4734,N_1558,N_2870);
and U4735 (N_4735,N_344,N_2994);
or U4736 (N_4736,N_1246,N_1012);
or U4737 (N_4737,N_1267,N_1689);
and U4738 (N_4738,N_576,N_629);
xnor U4739 (N_4739,N_2323,N_2414);
nand U4740 (N_4740,N_623,N_1073);
xor U4741 (N_4741,N_2051,N_851);
or U4742 (N_4742,N_578,N_184);
xor U4743 (N_4743,N_2334,N_2414);
nor U4744 (N_4744,N_208,N_1258);
nand U4745 (N_4745,N_2189,N_508);
and U4746 (N_4746,N_2663,N_426);
xor U4747 (N_4747,N_449,N_1896);
or U4748 (N_4748,N_625,N_238);
and U4749 (N_4749,N_172,N_1787);
and U4750 (N_4750,N_1336,N_1123);
or U4751 (N_4751,N_2463,N_797);
nand U4752 (N_4752,N_2045,N_2264);
nand U4753 (N_4753,N_1638,N_2931);
nand U4754 (N_4754,N_1282,N_2253);
nor U4755 (N_4755,N_1372,N_180);
and U4756 (N_4756,N_2053,N_438);
nor U4757 (N_4757,N_1945,N_2482);
nor U4758 (N_4758,N_67,N_1291);
xor U4759 (N_4759,N_185,N_2696);
xnor U4760 (N_4760,N_926,N_758);
or U4761 (N_4761,N_2646,N_2418);
and U4762 (N_4762,N_311,N_2098);
or U4763 (N_4763,N_1059,N_1451);
xor U4764 (N_4764,N_98,N_2919);
or U4765 (N_4765,N_1097,N_1557);
or U4766 (N_4766,N_1873,N_2914);
xnor U4767 (N_4767,N_1087,N_126);
nand U4768 (N_4768,N_601,N_771);
and U4769 (N_4769,N_1737,N_2477);
xnor U4770 (N_4770,N_1970,N_2855);
xnor U4771 (N_4771,N_685,N_2810);
xor U4772 (N_4772,N_749,N_1556);
or U4773 (N_4773,N_1663,N_2829);
and U4774 (N_4774,N_1902,N_703);
and U4775 (N_4775,N_1049,N_161);
xor U4776 (N_4776,N_1362,N_1192);
nor U4777 (N_4777,N_2785,N_353);
xnor U4778 (N_4778,N_1892,N_414);
nand U4779 (N_4779,N_2530,N_1440);
nand U4780 (N_4780,N_417,N_2758);
or U4781 (N_4781,N_59,N_2266);
and U4782 (N_4782,N_2554,N_2757);
and U4783 (N_4783,N_2867,N_2475);
nand U4784 (N_4784,N_91,N_118);
xnor U4785 (N_4785,N_1384,N_10);
or U4786 (N_4786,N_1671,N_2200);
and U4787 (N_4787,N_2344,N_489);
and U4788 (N_4788,N_1459,N_1492);
nor U4789 (N_4789,N_2294,N_840);
xnor U4790 (N_4790,N_2145,N_2872);
and U4791 (N_4791,N_2121,N_2318);
nand U4792 (N_4792,N_1343,N_2697);
and U4793 (N_4793,N_1068,N_2554);
or U4794 (N_4794,N_939,N_2262);
and U4795 (N_4795,N_1830,N_2668);
and U4796 (N_4796,N_2274,N_1212);
nor U4797 (N_4797,N_2948,N_1398);
or U4798 (N_4798,N_2221,N_819);
and U4799 (N_4799,N_440,N_1156);
nor U4800 (N_4800,N_18,N_1326);
nor U4801 (N_4801,N_942,N_2166);
xor U4802 (N_4802,N_1049,N_353);
xnor U4803 (N_4803,N_537,N_806);
nor U4804 (N_4804,N_1981,N_366);
nand U4805 (N_4805,N_1968,N_1088);
and U4806 (N_4806,N_1782,N_1217);
nor U4807 (N_4807,N_712,N_973);
xnor U4808 (N_4808,N_767,N_2071);
nor U4809 (N_4809,N_1070,N_2941);
nor U4810 (N_4810,N_1833,N_2368);
xor U4811 (N_4811,N_2857,N_1581);
nor U4812 (N_4812,N_2461,N_2866);
nor U4813 (N_4813,N_2972,N_742);
or U4814 (N_4814,N_2798,N_549);
nor U4815 (N_4815,N_735,N_44);
and U4816 (N_4816,N_1448,N_1619);
and U4817 (N_4817,N_2349,N_2242);
nand U4818 (N_4818,N_223,N_2310);
nor U4819 (N_4819,N_361,N_1969);
xor U4820 (N_4820,N_342,N_1118);
nand U4821 (N_4821,N_290,N_2177);
xnor U4822 (N_4822,N_21,N_2484);
nand U4823 (N_4823,N_1496,N_1309);
xnor U4824 (N_4824,N_754,N_1344);
or U4825 (N_4825,N_2264,N_900);
nor U4826 (N_4826,N_2933,N_1543);
xor U4827 (N_4827,N_635,N_291);
nand U4828 (N_4828,N_1623,N_1311);
and U4829 (N_4829,N_2847,N_925);
xnor U4830 (N_4830,N_1921,N_432);
nor U4831 (N_4831,N_2698,N_1285);
nand U4832 (N_4832,N_1766,N_2590);
nor U4833 (N_4833,N_350,N_1850);
nand U4834 (N_4834,N_2570,N_1055);
and U4835 (N_4835,N_775,N_1995);
xnor U4836 (N_4836,N_954,N_1687);
and U4837 (N_4837,N_1863,N_2654);
and U4838 (N_4838,N_2909,N_298);
xor U4839 (N_4839,N_2986,N_478);
and U4840 (N_4840,N_398,N_2551);
nor U4841 (N_4841,N_2521,N_960);
nand U4842 (N_4842,N_2994,N_1039);
or U4843 (N_4843,N_2851,N_2760);
or U4844 (N_4844,N_86,N_1795);
or U4845 (N_4845,N_1434,N_180);
and U4846 (N_4846,N_1059,N_2161);
or U4847 (N_4847,N_1956,N_2061);
xor U4848 (N_4848,N_1834,N_59);
nand U4849 (N_4849,N_2451,N_1579);
nor U4850 (N_4850,N_2159,N_2776);
and U4851 (N_4851,N_2179,N_1804);
nand U4852 (N_4852,N_356,N_1148);
and U4853 (N_4853,N_2076,N_2815);
nor U4854 (N_4854,N_2181,N_623);
and U4855 (N_4855,N_1083,N_2287);
nand U4856 (N_4856,N_1152,N_1171);
nand U4857 (N_4857,N_268,N_1451);
nand U4858 (N_4858,N_2172,N_837);
and U4859 (N_4859,N_1682,N_293);
or U4860 (N_4860,N_2386,N_499);
and U4861 (N_4861,N_2501,N_858);
xor U4862 (N_4862,N_475,N_769);
xor U4863 (N_4863,N_1061,N_504);
nand U4864 (N_4864,N_264,N_2867);
nor U4865 (N_4865,N_765,N_2637);
xnor U4866 (N_4866,N_2549,N_2073);
and U4867 (N_4867,N_2010,N_2000);
xnor U4868 (N_4868,N_1022,N_1145);
or U4869 (N_4869,N_1176,N_2929);
nand U4870 (N_4870,N_26,N_1463);
and U4871 (N_4871,N_1468,N_2162);
nand U4872 (N_4872,N_2454,N_982);
nand U4873 (N_4873,N_2601,N_2921);
nand U4874 (N_4874,N_774,N_2892);
and U4875 (N_4875,N_2856,N_1727);
nand U4876 (N_4876,N_2001,N_2303);
and U4877 (N_4877,N_291,N_197);
xor U4878 (N_4878,N_1792,N_1759);
xnor U4879 (N_4879,N_2252,N_2434);
nand U4880 (N_4880,N_1236,N_1187);
xor U4881 (N_4881,N_2923,N_1013);
or U4882 (N_4882,N_5,N_1444);
or U4883 (N_4883,N_2385,N_645);
or U4884 (N_4884,N_2015,N_1968);
nand U4885 (N_4885,N_464,N_1245);
or U4886 (N_4886,N_1897,N_347);
nor U4887 (N_4887,N_2269,N_1823);
nor U4888 (N_4888,N_1954,N_1145);
nand U4889 (N_4889,N_112,N_867);
and U4890 (N_4890,N_345,N_756);
nor U4891 (N_4891,N_952,N_2532);
or U4892 (N_4892,N_2442,N_517);
nand U4893 (N_4893,N_538,N_169);
nand U4894 (N_4894,N_402,N_996);
nand U4895 (N_4895,N_1655,N_992);
xor U4896 (N_4896,N_250,N_2746);
xor U4897 (N_4897,N_2483,N_1476);
xor U4898 (N_4898,N_1939,N_2652);
and U4899 (N_4899,N_2355,N_2198);
or U4900 (N_4900,N_1258,N_614);
xnor U4901 (N_4901,N_2158,N_341);
or U4902 (N_4902,N_450,N_248);
nand U4903 (N_4903,N_2270,N_1049);
or U4904 (N_4904,N_2274,N_2871);
nor U4905 (N_4905,N_2397,N_2648);
and U4906 (N_4906,N_1610,N_1241);
and U4907 (N_4907,N_1131,N_577);
and U4908 (N_4908,N_1301,N_247);
nand U4909 (N_4909,N_2045,N_364);
xor U4910 (N_4910,N_890,N_1741);
xor U4911 (N_4911,N_1797,N_1943);
xnor U4912 (N_4912,N_1963,N_2163);
nand U4913 (N_4913,N_2450,N_2571);
or U4914 (N_4914,N_334,N_2135);
or U4915 (N_4915,N_1181,N_2260);
or U4916 (N_4916,N_1793,N_903);
or U4917 (N_4917,N_1330,N_244);
xnor U4918 (N_4918,N_1389,N_1921);
nand U4919 (N_4919,N_2154,N_86);
or U4920 (N_4920,N_1533,N_2409);
and U4921 (N_4921,N_1088,N_2109);
nor U4922 (N_4922,N_1468,N_669);
nor U4923 (N_4923,N_1094,N_2568);
nand U4924 (N_4924,N_1420,N_1101);
nand U4925 (N_4925,N_2795,N_2806);
or U4926 (N_4926,N_890,N_1112);
nor U4927 (N_4927,N_2923,N_2804);
or U4928 (N_4928,N_2621,N_1603);
or U4929 (N_4929,N_2660,N_2261);
xor U4930 (N_4930,N_2820,N_2985);
or U4931 (N_4931,N_506,N_949);
and U4932 (N_4932,N_1777,N_2848);
or U4933 (N_4933,N_2340,N_823);
or U4934 (N_4934,N_57,N_743);
nand U4935 (N_4935,N_2797,N_2621);
nor U4936 (N_4936,N_2362,N_2427);
nor U4937 (N_4937,N_2630,N_2612);
nor U4938 (N_4938,N_768,N_1690);
and U4939 (N_4939,N_1517,N_2027);
nand U4940 (N_4940,N_722,N_299);
nand U4941 (N_4941,N_1330,N_634);
and U4942 (N_4942,N_660,N_1060);
or U4943 (N_4943,N_748,N_2411);
and U4944 (N_4944,N_2347,N_379);
nand U4945 (N_4945,N_2377,N_768);
nand U4946 (N_4946,N_1446,N_592);
xnor U4947 (N_4947,N_2042,N_1485);
or U4948 (N_4948,N_2505,N_1105);
nor U4949 (N_4949,N_2044,N_2022);
and U4950 (N_4950,N_16,N_1625);
nor U4951 (N_4951,N_166,N_2165);
or U4952 (N_4952,N_2517,N_2116);
nand U4953 (N_4953,N_1068,N_873);
and U4954 (N_4954,N_2730,N_539);
xnor U4955 (N_4955,N_179,N_145);
and U4956 (N_4956,N_1766,N_1131);
and U4957 (N_4957,N_94,N_2445);
and U4958 (N_4958,N_118,N_2539);
and U4959 (N_4959,N_1623,N_2741);
xnor U4960 (N_4960,N_1726,N_1590);
xnor U4961 (N_4961,N_1738,N_759);
nand U4962 (N_4962,N_1266,N_2990);
and U4963 (N_4963,N_11,N_2644);
xor U4964 (N_4964,N_1615,N_2557);
and U4965 (N_4965,N_208,N_2067);
nand U4966 (N_4966,N_1841,N_730);
nor U4967 (N_4967,N_2165,N_1167);
or U4968 (N_4968,N_1004,N_1102);
or U4969 (N_4969,N_2242,N_148);
nand U4970 (N_4970,N_2471,N_21);
xor U4971 (N_4971,N_1297,N_779);
xnor U4972 (N_4972,N_1858,N_2052);
or U4973 (N_4973,N_1123,N_364);
and U4974 (N_4974,N_2278,N_1150);
nand U4975 (N_4975,N_153,N_410);
nand U4976 (N_4976,N_2921,N_2975);
or U4977 (N_4977,N_707,N_2319);
nor U4978 (N_4978,N_658,N_1538);
xnor U4979 (N_4979,N_861,N_1384);
xnor U4980 (N_4980,N_772,N_1053);
nor U4981 (N_4981,N_290,N_2789);
nand U4982 (N_4982,N_1447,N_1282);
nor U4983 (N_4983,N_404,N_1615);
and U4984 (N_4984,N_1463,N_1277);
xor U4985 (N_4985,N_568,N_2554);
nor U4986 (N_4986,N_2667,N_486);
and U4987 (N_4987,N_1755,N_1669);
and U4988 (N_4988,N_1074,N_1922);
xnor U4989 (N_4989,N_1442,N_844);
xor U4990 (N_4990,N_1134,N_2575);
nand U4991 (N_4991,N_1110,N_2252);
and U4992 (N_4992,N_2140,N_1290);
xor U4993 (N_4993,N_82,N_1557);
or U4994 (N_4994,N_2358,N_2627);
nor U4995 (N_4995,N_1609,N_2120);
xor U4996 (N_4996,N_1837,N_1442);
or U4997 (N_4997,N_1092,N_881);
xnor U4998 (N_4998,N_2923,N_374);
and U4999 (N_4999,N_478,N_999);
nand U5000 (N_5000,N_777,N_1252);
or U5001 (N_5001,N_1617,N_234);
xor U5002 (N_5002,N_941,N_618);
nor U5003 (N_5003,N_678,N_2152);
or U5004 (N_5004,N_2605,N_2591);
nand U5005 (N_5005,N_2023,N_174);
xor U5006 (N_5006,N_2873,N_2973);
and U5007 (N_5007,N_1412,N_1647);
nor U5008 (N_5008,N_489,N_2390);
and U5009 (N_5009,N_1461,N_2362);
nand U5010 (N_5010,N_730,N_1089);
nor U5011 (N_5011,N_220,N_1087);
nor U5012 (N_5012,N_2153,N_1522);
nand U5013 (N_5013,N_2790,N_2147);
nor U5014 (N_5014,N_842,N_1157);
nand U5015 (N_5015,N_2328,N_1787);
nand U5016 (N_5016,N_1155,N_2010);
nor U5017 (N_5017,N_2355,N_445);
nand U5018 (N_5018,N_2673,N_2174);
and U5019 (N_5019,N_831,N_68);
or U5020 (N_5020,N_2443,N_1036);
nand U5021 (N_5021,N_2373,N_188);
nor U5022 (N_5022,N_477,N_2840);
nor U5023 (N_5023,N_1800,N_1762);
nand U5024 (N_5024,N_1699,N_2275);
xnor U5025 (N_5025,N_2776,N_845);
xnor U5026 (N_5026,N_370,N_724);
nand U5027 (N_5027,N_2836,N_2624);
xor U5028 (N_5028,N_2892,N_1951);
xnor U5029 (N_5029,N_2397,N_664);
nand U5030 (N_5030,N_592,N_2772);
nor U5031 (N_5031,N_1770,N_1538);
xnor U5032 (N_5032,N_2661,N_1033);
nand U5033 (N_5033,N_1096,N_2107);
xnor U5034 (N_5034,N_1740,N_2356);
or U5035 (N_5035,N_2541,N_33);
xnor U5036 (N_5036,N_956,N_2447);
or U5037 (N_5037,N_1763,N_2037);
nand U5038 (N_5038,N_964,N_1229);
or U5039 (N_5039,N_63,N_1955);
nor U5040 (N_5040,N_2965,N_573);
and U5041 (N_5041,N_1315,N_2711);
nor U5042 (N_5042,N_2904,N_358);
nor U5043 (N_5043,N_2758,N_2567);
nand U5044 (N_5044,N_1161,N_1664);
or U5045 (N_5045,N_2110,N_2698);
xnor U5046 (N_5046,N_2258,N_1770);
or U5047 (N_5047,N_2637,N_1683);
nand U5048 (N_5048,N_1920,N_710);
nand U5049 (N_5049,N_947,N_2321);
and U5050 (N_5050,N_251,N_1354);
nand U5051 (N_5051,N_1458,N_2569);
or U5052 (N_5052,N_1433,N_609);
nand U5053 (N_5053,N_1457,N_909);
xnor U5054 (N_5054,N_703,N_770);
and U5055 (N_5055,N_2138,N_2977);
or U5056 (N_5056,N_826,N_2159);
nand U5057 (N_5057,N_2597,N_134);
or U5058 (N_5058,N_954,N_202);
nor U5059 (N_5059,N_1387,N_2550);
nor U5060 (N_5060,N_1082,N_69);
xor U5061 (N_5061,N_2924,N_935);
or U5062 (N_5062,N_1577,N_920);
xnor U5063 (N_5063,N_1078,N_2748);
nor U5064 (N_5064,N_337,N_1367);
xor U5065 (N_5065,N_465,N_1718);
nor U5066 (N_5066,N_885,N_2190);
nand U5067 (N_5067,N_924,N_1482);
nor U5068 (N_5068,N_215,N_554);
nand U5069 (N_5069,N_1072,N_1006);
nand U5070 (N_5070,N_2040,N_484);
nor U5071 (N_5071,N_2410,N_1393);
nor U5072 (N_5072,N_980,N_191);
and U5073 (N_5073,N_1022,N_1059);
nand U5074 (N_5074,N_2397,N_2354);
nor U5075 (N_5075,N_2348,N_2198);
nor U5076 (N_5076,N_2465,N_1697);
and U5077 (N_5077,N_335,N_2282);
xnor U5078 (N_5078,N_2629,N_1513);
nor U5079 (N_5079,N_2707,N_520);
and U5080 (N_5080,N_434,N_1);
nand U5081 (N_5081,N_2862,N_1451);
and U5082 (N_5082,N_237,N_987);
or U5083 (N_5083,N_1681,N_1286);
and U5084 (N_5084,N_2003,N_2191);
nor U5085 (N_5085,N_997,N_943);
xnor U5086 (N_5086,N_1971,N_2341);
and U5087 (N_5087,N_1103,N_552);
or U5088 (N_5088,N_1349,N_577);
and U5089 (N_5089,N_2486,N_33);
and U5090 (N_5090,N_2710,N_2884);
xnor U5091 (N_5091,N_1337,N_2160);
or U5092 (N_5092,N_1214,N_2228);
or U5093 (N_5093,N_2591,N_2822);
nand U5094 (N_5094,N_2128,N_1085);
xor U5095 (N_5095,N_1487,N_896);
nand U5096 (N_5096,N_1377,N_360);
or U5097 (N_5097,N_1304,N_1595);
nor U5098 (N_5098,N_1020,N_1719);
nor U5099 (N_5099,N_2258,N_1810);
and U5100 (N_5100,N_759,N_163);
nand U5101 (N_5101,N_1489,N_2580);
nand U5102 (N_5102,N_2126,N_1223);
or U5103 (N_5103,N_969,N_354);
nand U5104 (N_5104,N_1674,N_463);
nor U5105 (N_5105,N_1611,N_701);
xnor U5106 (N_5106,N_1627,N_53);
nand U5107 (N_5107,N_1235,N_548);
nor U5108 (N_5108,N_2549,N_2095);
or U5109 (N_5109,N_1975,N_847);
nand U5110 (N_5110,N_662,N_1379);
or U5111 (N_5111,N_2137,N_1930);
xnor U5112 (N_5112,N_2921,N_1115);
nand U5113 (N_5113,N_950,N_2259);
xnor U5114 (N_5114,N_414,N_1484);
xnor U5115 (N_5115,N_2854,N_2521);
nand U5116 (N_5116,N_2065,N_2137);
or U5117 (N_5117,N_1090,N_2309);
or U5118 (N_5118,N_1105,N_2474);
nor U5119 (N_5119,N_1045,N_693);
and U5120 (N_5120,N_1471,N_1800);
xnor U5121 (N_5121,N_647,N_1800);
nor U5122 (N_5122,N_2231,N_2689);
nor U5123 (N_5123,N_1035,N_2951);
nand U5124 (N_5124,N_59,N_851);
and U5125 (N_5125,N_624,N_2338);
nand U5126 (N_5126,N_2931,N_1896);
nand U5127 (N_5127,N_636,N_2510);
xnor U5128 (N_5128,N_2292,N_1344);
xor U5129 (N_5129,N_1234,N_2063);
or U5130 (N_5130,N_1688,N_2866);
nor U5131 (N_5131,N_439,N_1284);
or U5132 (N_5132,N_94,N_1063);
or U5133 (N_5133,N_1769,N_1624);
xnor U5134 (N_5134,N_1553,N_375);
xnor U5135 (N_5135,N_2486,N_2729);
and U5136 (N_5136,N_1411,N_2233);
and U5137 (N_5137,N_802,N_391);
xnor U5138 (N_5138,N_1643,N_2404);
or U5139 (N_5139,N_1925,N_2173);
and U5140 (N_5140,N_2929,N_2325);
nor U5141 (N_5141,N_1101,N_1253);
or U5142 (N_5142,N_2057,N_1811);
nor U5143 (N_5143,N_2813,N_1216);
nand U5144 (N_5144,N_595,N_744);
and U5145 (N_5145,N_1849,N_2872);
and U5146 (N_5146,N_144,N_1639);
and U5147 (N_5147,N_1490,N_1039);
or U5148 (N_5148,N_149,N_48);
and U5149 (N_5149,N_1086,N_1336);
nor U5150 (N_5150,N_2540,N_454);
nand U5151 (N_5151,N_1376,N_646);
and U5152 (N_5152,N_817,N_1770);
or U5153 (N_5153,N_1706,N_527);
or U5154 (N_5154,N_1295,N_542);
xor U5155 (N_5155,N_1149,N_1246);
nor U5156 (N_5156,N_2206,N_677);
nor U5157 (N_5157,N_174,N_2960);
xor U5158 (N_5158,N_2155,N_2497);
xnor U5159 (N_5159,N_383,N_953);
nand U5160 (N_5160,N_1987,N_1859);
xor U5161 (N_5161,N_152,N_5);
nor U5162 (N_5162,N_419,N_509);
xor U5163 (N_5163,N_681,N_676);
xor U5164 (N_5164,N_1625,N_2980);
or U5165 (N_5165,N_1065,N_1746);
and U5166 (N_5166,N_1277,N_2679);
nor U5167 (N_5167,N_1804,N_2386);
or U5168 (N_5168,N_1947,N_1103);
nor U5169 (N_5169,N_536,N_369);
nor U5170 (N_5170,N_2046,N_105);
nand U5171 (N_5171,N_92,N_2914);
nand U5172 (N_5172,N_1467,N_1263);
and U5173 (N_5173,N_939,N_630);
or U5174 (N_5174,N_2471,N_811);
nor U5175 (N_5175,N_212,N_1530);
and U5176 (N_5176,N_1785,N_324);
and U5177 (N_5177,N_2602,N_353);
or U5178 (N_5178,N_2058,N_2117);
and U5179 (N_5179,N_532,N_236);
nor U5180 (N_5180,N_2526,N_794);
and U5181 (N_5181,N_1366,N_2944);
xnor U5182 (N_5182,N_1560,N_529);
nand U5183 (N_5183,N_2110,N_2548);
or U5184 (N_5184,N_2796,N_2689);
xor U5185 (N_5185,N_598,N_1561);
and U5186 (N_5186,N_613,N_387);
xnor U5187 (N_5187,N_2330,N_2874);
nand U5188 (N_5188,N_199,N_2733);
nor U5189 (N_5189,N_557,N_150);
or U5190 (N_5190,N_2251,N_2466);
and U5191 (N_5191,N_2882,N_908);
nor U5192 (N_5192,N_1935,N_2145);
and U5193 (N_5193,N_69,N_2029);
nor U5194 (N_5194,N_301,N_151);
and U5195 (N_5195,N_152,N_1059);
or U5196 (N_5196,N_2488,N_1635);
and U5197 (N_5197,N_1362,N_1749);
or U5198 (N_5198,N_2143,N_1858);
or U5199 (N_5199,N_1634,N_1880);
nor U5200 (N_5200,N_2591,N_1295);
nor U5201 (N_5201,N_2956,N_943);
nor U5202 (N_5202,N_1910,N_1163);
xnor U5203 (N_5203,N_1677,N_335);
nor U5204 (N_5204,N_1271,N_1811);
nor U5205 (N_5205,N_318,N_1926);
and U5206 (N_5206,N_96,N_193);
nor U5207 (N_5207,N_1198,N_1143);
and U5208 (N_5208,N_2772,N_2307);
or U5209 (N_5209,N_60,N_2148);
and U5210 (N_5210,N_646,N_692);
xor U5211 (N_5211,N_2809,N_2393);
or U5212 (N_5212,N_889,N_1161);
and U5213 (N_5213,N_498,N_2647);
xor U5214 (N_5214,N_2923,N_633);
nor U5215 (N_5215,N_2480,N_2063);
or U5216 (N_5216,N_987,N_1731);
or U5217 (N_5217,N_883,N_2485);
and U5218 (N_5218,N_2645,N_1522);
and U5219 (N_5219,N_172,N_873);
and U5220 (N_5220,N_2906,N_659);
nand U5221 (N_5221,N_2276,N_1547);
and U5222 (N_5222,N_195,N_1404);
nor U5223 (N_5223,N_498,N_1926);
or U5224 (N_5224,N_266,N_2792);
nand U5225 (N_5225,N_1120,N_2438);
or U5226 (N_5226,N_180,N_1066);
and U5227 (N_5227,N_1896,N_2023);
xor U5228 (N_5228,N_919,N_1188);
or U5229 (N_5229,N_2872,N_585);
xnor U5230 (N_5230,N_2089,N_1412);
and U5231 (N_5231,N_1471,N_2509);
xnor U5232 (N_5232,N_2377,N_2630);
nor U5233 (N_5233,N_2457,N_1064);
nand U5234 (N_5234,N_643,N_175);
xor U5235 (N_5235,N_2349,N_407);
and U5236 (N_5236,N_2891,N_273);
nand U5237 (N_5237,N_2055,N_1999);
or U5238 (N_5238,N_2912,N_266);
nand U5239 (N_5239,N_1161,N_1393);
and U5240 (N_5240,N_2434,N_1559);
nor U5241 (N_5241,N_1301,N_1539);
or U5242 (N_5242,N_2576,N_705);
nor U5243 (N_5243,N_2329,N_1022);
nor U5244 (N_5244,N_1580,N_1948);
nor U5245 (N_5245,N_1918,N_1256);
and U5246 (N_5246,N_2837,N_2472);
and U5247 (N_5247,N_2072,N_632);
xnor U5248 (N_5248,N_2484,N_461);
xnor U5249 (N_5249,N_224,N_2902);
or U5250 (N_5250,N_2801,N_2570);
nor U5251 (N_5251,N_375,N_440);
nor U5252 (N_5252,N_1580,N_1901);
or U5253 (N_5253,N_2251,N_2174);
nand U5254 (N_5254,N_1428,N_1884);
or U5255 (N_5255,N_879,N_1391);
and U5256 (N_5256,N_1776,N_2590);
or U5257 (N_5257,N_1079,N_389);
and U5258 (N_5258,N_240,N_1023);
and U5259 (N_5259,N_1017,N_1481);
nand U5260 (N_5260,N_1156,N_546);
nor U5261 (N_5261,N_94,N_1920);
nor U5262 (N_5262,N_2019,N_500);
nand U5263 (N_5263,N_122,N_828);
nor U5264 (N_5264,N_276,N_1325);
nand U5265 (N_5265,N_1374,N_1613);
nand U5266 (N_5266,N_181,N_2867);
nand U5267 (N_5267,N_1823,N_2299);
xnor U5268 (N_5268,N_1373,N_2617);
nor U5269 (N_5269,N_2266,N_2952);
nand U5270 (N_5270,N_2448,N_2456);
and U5271 (N_5271,N_1430,N_1737);
nand U5272 (N_5272,N_316,N_1229);
or U5273 (N_5273,N_2001,N_774);
nor U5274 (N_5274,N_607,N_1027);
nor U5275 (N_5275,N_1186,N_703);
nor U5276 (N_5276,N_441,N_1682);
nand U5277 (N_5277,N_2344,N_1765);
or U5278 (N_5278,N_883,N_718);
or U5279 (N_5279,N_1486,N_539);
nor U5280 (N_5280,N_2375,N_2590);
nand U5281 (N_5281,N_903,N_2723);
nand U5282 (N_5282,N_1678,N_496);
nand U5283 (N_5283,N_974,N_471);
or U5284 (N_5284,N_885,N_2439);
and U5285 (N_5285,N_7,N_1241);
or U5286 (N_5286,N_1665,N_33);
xor U5287 (N_5287,N_2290,N_1046);
nor U5288 (N_5288,N_249,N_1769);
nand U5289 (N_5289,N_2365,N_2419);
and U5290 (N_5290,N_1440,N_1449);
nor U5291 (N_5291,N_2747,N_2911);
nor U5292 (N_5292,N_2482,N_672);
or U5293 (N_5293,N_2767,N_1172);
and U5294 (N_5294,N_1273,N_940);
and U5295 (N_5295,N_1515,N_599);
or U5296 (N_5296,N_1763,N_2869);
and U5297 (N_5297,N_2986,N_2282);
nand U5298 (N_5298,N_2144,N_1564);
nand U5299 (N_5299,N_2893,N_2385);
and U5300 (N_5300,N_2517,N_2392);
and U5301 (N_5301,N_2494,N_694);
xor U5302 (N_5302,N_1657,N_2689);
nand U5303 (N_5303,N_463,N_50);
xnor U5304 (N_5304,N_211,N_1542);
xor U5305 (N_5305,N_12,N_1408);
nand U5306 (N_5306,N_751,N_182);
nand U5307 (N_5307,N_1534,N_568);
and U5308 (N_5308,N_1101,N_401);
nand U5309 (N_5309,N_2760,N_2748);
xnor U5310 (N_5310,N_1196,N_2395);
nand U5311 (N_5311,N_2313,N_356);
nand U5312 (N_5312,N_2883,N_2924);
and U5313 (N_5313,N_1283,N_2740);
nor U5314 (N_5314,N_751,N_1684);
and U5315 (N_5315,N_1351,N_1750);
xnor U5316 (N_5316,N_2345,N_2846);
nor U5317 (N_5317,N_2535,N_10);
nand U5318 (N_5318,N_689,N_32);
nor U5319 (N_5319,N_1443,N_1465);
or U5320 (N_5320,N_2070,N_2416);
or U5321 (N_5321,N_2950,N_2096);
nor U5322 (N_5322,N_2489,N_1461);
or U5323 (N_5323,N_2178,N_2377);
and U5324 (N_5324,N_240,N_802);
and U5325 (N_5325,N_859,N_792);
xor U5326 (N_5326,N_60,N_75);
and U5327 (N_5327,N_2676,N_1630);
or U5328 (N_5328,N_2043,N_1666);
or U5329 (N_5329,N_2971,N_239);
nand U5330 (N_5330,N_2617,N_1157);
or U5331 (N_5331,N_250,N_764);
nor U5332 (N_5332,N_1912,N_1555);
nor U5333 (N_5333,N_1738,N_566);
xor U5334 (N_5334,N_1783,N_305);
nand U5335 (N_5335,N_2530,N_547);
xor U5336 (N_5336,N_2506,N_1200);
or U5337 (N_5337,N_2152,N_950);
xnor U5338 (N_5338,N_1968,N_1894);
nor U5339 (N_5339,N_975,N_172);
nand U5340 (N_5340,N_178,N_2823);
nand U5341 (N_5341,N_940,N_78);
nand U5342 (N_5342,N_1613,N_1280);
or U5343 (N_5343,N_2121,N_644);
and U5344 (N_5344,N_2386,N_1299);
nand U5345 (N_5345,N_2865,N_2894);
nand U5346 (N_5346,N_1602,N_2156);
xnor U5347 (N_5347,N_436,N_1785);
and U5348 (N_5348,N_2186,N_77);
and U5349 (N_5349,N_1072,N_415);
xnor U5350 (N_5350,N_190,N_2501);
nor U5351 (N_5351,N_511,N_1887);
or U5352 (N_5352,N_1902,N_2435);
xnor U5353 (N_5353,N_1850,N_2904);
nand U5354 (N_5354,N_1903,N_2484);
and U5355 (N_5355,N_2460,N_2311);
and U5356 (N_5356,N_46,N_1326);
nand U5357 (N_5357,N_1503,N_1654);
and U5358 (N_5358,N_1189,N_1786);
and U5359 (N_5359,N_2652,N_1773);
nor U5360 (N_5360,N_271,N_667);
nor U5361 (N_5361,N_2530,N_1434);
or U5362 (N_5362,N_1922,N_1317);
nand U5363 (N_5363,N_243,N_2431);
xor U5364 (N_5364,N_1211,N_1180);
nor U5365 (N_5365,N_1620,N_2129);
nor U5366 (N_5366,N_457,N_842);
xnor U5367 (N_5367,N_1389,N_2548);
and U5368 (N_5368,N_407,N_2869);
nand U5369 (N_5369,N_2684,N_2030);
nand U5370 (N_5370,N_2008,N_160);
nor U5371 (N_5371,N_1767,N_65);
xor U5372 (N_5372,N_2676,N_418);
nor U5373 (N_5373,N_2123,N_1161);
nand U5374 (N_5374,N_82,N_1124);
nor U5375 (N_5375,N_1449,N_1234);
or U5376 (N_5376,N_981,N_262);
xnor U5377 (N_5377,N_2262,N_820);
nor U5378 (N_5378,N_2702,N_1124);
or U5379 (N_5379,N_714,N_2281);
nor U5380 (N_5380,N_2026,N_1436);
and U5381 (N_5381,N_139,N_876);
xnor U5382 (N_5382,N_980,N_1459);
and U5383 (N_5383,N_1327,N_321);
or U5384 (N_5384,N_257,N_2633);
xnor U5385 (N_5385,N_1516,N_1004);
nor U5386 (N_5386,N_1590,N_2110);
nand U5387 (N_5387,N_286,N_1284);
or U5388 (N_5388,N_1732,N_2801);
and U5389 (N_5389,N_2486,N_751);
nand U5390 (N_5390,N_665,N_654);
nand U5391 (N_5391,N_2779,N_2555);
xor U5392 (N_5392,N_1364,N_2540);
and U5393 (N_5393,N_1613,N_782);
or U5394 (N_5394,N_1063,N_461);
xor U5395 (N_5395,N_2772,N_2286);
xnor U5396 (N_5396,N_2433,N_2574);
xor U5397 (N_5397,N_1266,N_396);
xor U5398 (N_5398,N_581,N_932);
nand U5399 (N_5399,N_2515,N_2402);
nor U5400 (N_5400,N_243,N_2075);
xnor U5401 (N_5401,N_2855,N_1829);
or U5402 (N_5402,N_2362,N_2721);
or U5403 (N_5403,N_2690,N_379);
and U5404 (N_5404,N_2454,N_129);
nand U5405 (N_5405,N_1756,N_1562);
and U5406 (N_5406,N_241,N_11);
or U5407 (N_5407,N_1057,N_1753);
xor U5408 (N_5408,N_1860,N_2888);
nor U5409 (N_5409,N_1088,N_2630);
xor U5410 (N_5410,N_2950,N_2061);
nand U5411 (N_5411,N_675,N_34);
or U5412 (N_5412,N_851,N_1057);
nor U5413 (N_5413,N_1216,N_2027);
and U5414 (N_5414,N_1256,N_1546);
xor U5415 (N_5415,N_1152,N_2235);
nor U5416 (N_5416,N_1526,N_1533);
xnor U5417 (N_5417,N_2472,N_413);
or U5418 (N_5418,N_421,N_79);
nand U5419 (N_5419,N_1820,N_211);
xor U5420 (N_5420,N_1195,N_1805);
nand U5421 (N_5421,N_1945,N_1461);
nor U5422 (N_5422,N_161,N_439);
xor U5423 (N_5423,N_961,N_279);
nor U5424 (N_5424,N_2736,N_1643);
and U5425 (N_5425,N_269,N_2276);
nand U5426 (N_5426,N_135,N_1510);
xnor U5427 (N_5427,N_95,N_180);
nor U5428 (N_5428,N_1120,N_2779);
xor U5429 (N_5429,N_2168,N_359);
and U5430 (N_5430,N_515,N_141);
nor U5431 (N_5431,N_2732,N_1800);
or U5432 (N_5432,N_1676,N_2617);
or U5433 (N_5433,N_1214,N_2972);
or U5434 (N_5434,N_446,N_2058);
nand U5435 (N_5435,N_1869,N_2492);
or U5436 (N_5436,N_1666,N_155);
and U5437 (N_5437,N_2389,N_1888);
and U5438 (N_5438,N_1470,N_695);
nand U5439 (N_5439,N_1061,N_1173);
or U5440 (N_5440,N_2561,N_2745);
nor U5441 (N_5441,N_2358,N_2046);
xor U5442 (N_5442,N_77,N_573);
nand U5443 (N_5443,N_392,N_1541);
or U5444 (N_5444,N_1216,N_2774);
nand U5445 (N_5445,N_1803,N_1243);
or U5446 (N_5446,N_2755,N_1530);
or U5447 (N_5447,N_1215,N_1872);
nand U5448 (N_5448,N_1111,N_1180);
or U5449 (N_5449,N_214,N_849);
nor U5450 (N_5450,N_1714,N_2284);
nor U5451 (N_5451,N_1809,N_2833);
or U5452 (N_5452,N_693,N_28);
nand U5453 (N_5453,N_961,N_80);
nor U5454 (N_5454,N_166,N_2606);
or U5455 (N_5455,N_2500,N_413);
and U5456 (N_5456,N_908,N_1330);
or U5457 (N_5457,N_2116,N_821);
xnor U5458 (N_5458,N_310,N_956);
and U5459 (N_5459,N_1526,N_1713);
xor U5460 (N_5460,N_1639,N_637);
xnor U5461 (N_5461,N_2950,N_1308);
and U5462 (N_5462,N_1634,N_1580);
xor U5463 (N_5463,N_406,N_2470);
nor U5464 (N_5464,N_2155,N_1103);
and U5465 (N_5465,N_994,N_143);
nor U5466 (N_5466,N_1884,N_2713);
nand U5467 (N_5467,N_2877,N_1743);
nand U5468 (N_5468,N_2007,N_1057);
nand U5469 (N_5469,N_2733,N_940);
xor U5470 (N_5470,N_1413,N_779);
nor U5471 (N_5471,N_2753,N_393);
xor U5472 (N_5472,N_742,N_293);
nand U5473 (N_5473,N_1168,N_1511);
nand U5474 (N_5474,N_2004,N_147);
nor U5475 (N_5475,N_2165,N_336);
nor U5476 (N_5476,N_745,N_2116);
nor U5477 (N_5477,N_142,N_2426);
and U5478 (N_5478,N_1409,N_2796);
and U5479 (N_5479,N_664,N_546);
nor U5480 (N_5480,N_2592,N_1834);
or U5481 (N_5481,N_2566,N_2448);
or U5482 (N_5482,N_2361,N_1744);
xnor U5483 (N_5483,N_2069,N_2812);
and U5484 (N_5484,N_1622,N_685);
nor U5485 (N_5485,N_2463,N_1586);
or U5486 (N_5486,N_21,N_562);
nand U5487 (N_5487,N_2715,N_2209);
nand U5488 (N_5488,N_2685,N_1438);
xnor U5489 (N_5489,N_2908,N_321);
xor U5490 (N_5490,N_1874,N_2339);
or U5491 (N_5491,N_2135,N_2925);
and U5492 (N_5492,N_1490,N_667);
and U5493 (N_5493,N_2081,N_2547);
and U5494 (N_5494,N_2948,N_2390);
nand U5495 (N_5495,N_1871,N_1587);
or U5496 (N_5496,N_789,N_91);
or U5497 (N_5497,N_1761,N_599);
and U5498 (N_5498,N_1248,N_2208);
or U5499 (N_5499,N_881,N_1680);
xnor U5500 (N_5500,N_799,N_2666);
xor U5501 (N_5501,N_2983,N_1883);
nand U5502 (N_5502,N_1059,N_2814);
nor U5503 (N_5503,N_1756,N_1804);
and U5504 (N_5504,N_2246,N_1602);
nand U5505 (N_5505,N_496,N_2570);
or U5506 (N_5506,N_455,N_1352);
or U5507 (N_5507,N_2383,N_1210);
or U5508 (N_5508,N_844,N_157);
xnor U5509 (N_5509,N_2320,N_2511);
xor U5510 (N_5510,N_1465,N_2958);
or U5511 (N_5511,N_2395,N_562);
nand U5512 (N_5512,N_1585,N_1874);
nor U5513 (N_5513,N_18,N_2372);
and U5514 (N_5514,N_1445,N_2273);
and U5515 (N_5515,N_2997,N_2559);
nand U5516 (N_5516,N_2952,N_2323);
xnor U5517 (N_5517,N_2543,N_323);
or U5518 (N_5518,N_813,N_2693);
nand U5519 (N_5519,N_2676,N_2843);
nor U5520 (N_5520,N_2202,N_1121);
nor U5521 (N_5521,N_2562,N_2943);
or U5522 (N_5522,N_2936,N_2623);
nor U5523 (N_5523,N_2838,N_1369);
nand U5524 (N_5524,N_2655,N_2386);
and U5525 (N_5525,N_312,N_768);
and U5526 (N_5526,N_2264,N_2818);
xor U5527 (N_5527,N_1594,N_2576);
nor U5528 (N_5528,N_1176,N_1876);
or U5529 (N_5529,N_2661,N_1397);
xnor U5530 (N_5530,N_1471,N_1297);
nor U5531 (N_5531,N_1213,N_27);
xnor U5532 (N_5532,N_245,N_2446);
nor U5533 (N_5533,N_2692,N_2042);
and U5534 (N_5534,N_93,N_1373);
nand U5535 (N_5535,N_952,N_1170);
nor U5536 (N_5536,N_2219,N_229);
or U5537 (N_5537,N_2880,N_478);
nor U5538 (N_5538,N_1955,N_2441);
and U5539 (N_5539,N_1937,N_293);
or U5540 (N_5540,N_2622,N_1513);
or U5541 (N_5541,N_2977,N_1839);
and U5542 (N_5542,N_487,N_1028);
xor U5543 (N_5543,N_1049,N_122);
nand U5544 (N_5544,N_57,N_1313);
nand U5545 (N_5545,N_1899,N_1012);
xor U5546 (N_5546,N_475,N_1348);
nand U5547 (N_5547,N_332,N_1509);
nor U5548 (N_5548,N_443,N_1941);
nand U5549 (N_5549,N_2161,N_1517);
xor U5550 (N_5550,N_1668,N_2507);
and U5551 (N_5551,N_1876,N_2977);
and U5552 (N_5552,N_1804,N_659);
xnor U5553 (N_5553,N_2833,N_1614);
and U5554 (N_5554,N_1919,N_943);
xnor U5555 (N_5555,N_1353,N_549);
or U5556 (N_5556,N_2922,N_2780);
nand U5557 (N_5557,N_1496,N_1050);
xnor U5558 (N_5558,N_2529,N_837);
nand U5559 (N_5559,N_2761,N_244);
and U5560 (N_5560,N_2140,N_230);
and U5561 (N_5561,N_1490,N_148);
and U5562 (N_5562,N_444,N_2415);
and U5563 (N_5563,N_400,N_291);
and U5564 (N_5564,N_1688,N_1841);
and U5565 (N_5565,N_2478,N_362);
or U5566 (N_5566,N_322,N_2680);
nor U5567 (N_5567,N_2151,N_2604);
or U5568 (N_5568,N_786,N_1690);
nor U5569 (N_5569,N_1352,N_351);
nor U5570 (N_5570,N_513,N_1235);
or U5571 (N_5571,N_2983,N_1618);
nor U5572 (N_5572,N_848,N_606);
nor U5573 (N_5573,N_1719,N_1221);
nor U5574 (N_5574,N_1697,N_2838);
or U5575 (N_5575,N_84,N_2737);
xor U5576 (N_5576,N_1091,N_1492);
and U5577 (N_5577,N_1214,N_2537);
xnor U5578 (N_5578,N_1779,N_713);
and U5579 (N_5579,N_825,N_57);
xor U5580 (N_5580,N_1419,N_1737);
nand U5581 (N_5581,N_1574,N_2199);
and U5582 (N_5582,N_2339,N_822);
nand U5583 (N_5583,N_2285,N_2869);
nor U5584 (N_5584,N_1382,N_200);
nor U5585 (N_5585,N_2075,N_1148);
or U5586 (N_5586,N_2734,N_2905);
and U5587 (N_5587,N_2355,N_2371);
nor U5588 (N_5588,N_2699,N_2141);
or U5589 (N_5589,N_185,N_2592);
nor U5590 (N_5590,N_2978,N_2384);
and U5591 (N_5591,N_1691,N_2700);
nand U5592 (N_5592,N_2374,N_2670);
or U5593 (N_5593,N_2703,N_1813);
xnor U5594 (N_5594,N_2688,N_2578);
nand U5595 (N_5595,N_1252,N_101);
nand U5596 (N_5596,N_396,N_1472);
nand U5597 (N_5597,N_2754,N_2403);
and U5598 (N_5598,N_935,N_2747);
nor U5599 (N_5599,N_1969,N_2001);
or U5600 (N_5600,N_2759,N_1339);
and U5601 (N_5601,N_1075,N_781);
xnor U5602 (N_5602,N_2852,N_1964);
nor U5603 (N_5603,N_2315,N_979);
nand U5604 (N_5604,N_1694,N_2659);
nor U5605 (N_5605,N_2322,N_970);
nand U5606 (N_5606,N_2588,N_2711);
nand U5607 (N_5607,N_1271,N_311);
xor U5608 (N_5608,N_395,N_1722);
and U5609 (N_5609,N_2218,N_1987);
nand U5610 (N_5610,N_1945,N_844);
xor U5611 (N_5611,N_2960,N_737);
xor U5612 (N_5612,N_2357,N_555);
and U5613 (N_5613,N_285,N_2006);
or U5614 (N_5614,N_1018,N_1165);
and U5615 (N_5615,N_1722,N_747);
xor U5616 (N_5616,N_65,N_2380);
and U5617 (N_5617,N_353,N_283);
nor U5618 (N_5618,N_1973,N_2779);
and U5619 (N_5619,N_2470,N_2774);
nand U5620 (N_5620,N_1933,N_1913);
nand U5621 (N_5621,N_2830,N_2006);
nor U5622 (N_5622,N_1653,N_1820);
or U5623 (N_5623,N_1691,N_542);
nor U5624 (N_5624,N_2674,N_1173);
nor U5625 (N_5625,N_2085,N_2974);
and U5626 (N_5626,N_397,N_2356);
xnor U5627 (N_5627,N_2906,N_2761);
nor U5628 (N_5628,N_1185,N_2204);
nand U5629 (N_5629,N_1889,N_1302);
nor U5630 (N_5630,N_763,N_2646);
xnor U5631 (N_5631,N_993,N_173);
xnor U5632 (N_5632,N_2211,N_1218);
nand U5633 (N_5633,N_113,N_943);
xnor U5634 (N_5634,N_662,N_781);
and U5635 (N_5635,N_330,N_970);
xor U5636 (N_5636,N_2199,N_135);
xnor U5637 (N_5637,N_2361,N_1564);
and U5638 (N_5638,N_944,N_96);
or U5639 (N_5639,N_1696,N_1272);
and U5640 (N_5640,N_2650,N_2864);
or U5641 (N_5641,N_726,N_2221);
nand U5642 (N_5642,N_474,N_524);
and U5643 (N_5643,N_2678,N_2285);
nor U5644 (N_5644,N_1289,N_613);
nor U5645 (N_5645,N_2615,N_1999);
or U5646 (N_5646,N_360,N_2352);
xnor U5647 (N_5647,N_388,N_2863);
xor U5648 (N_5648,N_2669,N_829);
or U5649 (N_5649,N_2506,N_1483);
and U5650 (N_5650,N_1649,N_1960);
and U5651 (N_5651,N_1082,N_1709);
nor U5652 (N_5652,N_1321,N_982);
and U5653 (N_5653,N_2523,N_1701);
nand U5654 (N_5654,N_898,N_174);
xor U5655 (N_5655,N_1547,N_990);
xor U5656 (N_5656,N_494,N_1572);
nand U5657 (N_5657,N_2275,N_2400);
nor U5658 (N_5658,N_1449,N_1177);
nand U5659 (N_5659,N_1280,N_2429);
nand U5660 (N_5660,N_2929,N_454);
and U5661 (N_5661,N_812,N_2214);
xor U5662 (N_5662,N_590,N_2941);
nor U5663 (N_5663,N_670,N_182);
xnor U5664 (N_5664,N_2277,N_2505);
nor U5665 (N_5665,N_29,N_355);
xnor U5666 (N_5666,N_209,N_1966);
nand U5667 (N_5667,N_2855,N_602);
xor U5668 (N_5668,N_1193,N_2448);
and U5669 (N_5669,N_1562,N_2888);
and U5670 (N_5670,N_2321,N_1199);
xor U5671 (N_5671,N_2866,N_230);
nor U5672 (N_5672,N_2810,N_709);
and U5673 (N_5673,N_2469,N_1287);
nor U5674 (N_5674,N_2023,N_192);
xnor U5675 (N_5675,N_323,N_2876);
nor U5676 (N_5676,N_1223,N_1292);
nand U5677 (N_5677,N_2448,N_2052);
nand U5678 (N_5678,N_1905,N_1231);
xor U5679 (N_5679,N_2762,N_264);
and U5680 (N_5680,N_1674,N_1660);
and U5681 (N_5681,N_1247,N_1668);
xor U5682 (N_5682,N_1393,N_2337);
and U5683 (N_5683,N_2368,N_295);
nand U5684 (N_5684,N_2435,N_2280);
and U5685 (N_5685,N_264,N_1251);
nor U5686 (N_5686,N_466,N_1236);
nor U5687 (N_5687,N_1013,N_2588);
and U5688 (N_5688,N_1444,N_1925);
and U5689 (N_5689,N_2266,N_224);
and U5690 (N_5690,N_1923,N_2835);
or U5691 (N_5691,N_1969,N_113);
xnor U5692 (N_5692,N_404,N_209);
nor U5693 (N_5693,N_2714,N_2623);
xnor U5694 (N_5694,N_2040,N_1395);
and U5695 (N_5695,N_1647,N_117);
and U5696 (N_5696,N_909,N_1045);
xor U5697 (N_5697,N_1144,N_1979);
nor U5698 (N_5698,N_1055,N_2942);
nor U5699 (N_5699,N_267,N_2561);
nand U5700 (N_5700,N_1748,N_2062);
nand U5701 (N_5701,N_1557,N_534);
and U5702 (N_5702,N_2325,N_2580);
nor U5703 (N_5703,N_2246,N_2104);
or U5704 (N_5704,N_1269,N_919);
xnor U5705 (N_5705,N_2528,N_1245);
or U5706 (N_5706,N_1448,N_535);
nand U5707 (N_5707,N_2047,N_1284);
nand U5708 (N_5708,N_2879,N_2440);
nor U5709 (N_5709,N_2051,N_1433);
or U5710 (N_5710,N_893,N_2138);
or U5711 (N_5711,N_300,N_2675);
and U5712 (N_5712,N_2276,N_1369);
or U5713 (N_5713,N_2713,N_1440);
nor U5714 (N_5714,N_2951,N_1085);
nor U5715 (N_5715,N_1164,N_2893);
and U5716 (N_5716,N_2619,N_1285);
or U5717 (N_5717,N_570,N_1366);
or U5718 (N_5718,N_189,N_555);
nand U5719 (N_5719,N_898,N_2996);
xnor U5720 (N_5720,N_2175,N_929);
or U5721 (N_5721,N_142,N_1387);
or U5722 (N_5722,N_2673,N_872);
nand U5723 (N_5723,N_1333,N_208);
nor U5724 (N_5724,N_1723,N_2730);
nand U5725 (N_5725,N_278,N_1454);
and U5726 (N_5726,N_2486,N_1754);
or U5727 (N_5727,N_1922,N_983);
or U5728 (N_5728,N_1350,N_300);
or U5729 (N_5729,N_701,N_2908);
and U5730 (N_5730,N_1299,N_167);
nor U5731 (N_5731,N_1660,N_2083);
nor U5732 (N_5732,N_240,N_876);
nor U5733 (N_5733,N_458,N_559);
and U5734 (N_5734,N_2686,N_1452);
and U5735 (N_5735,N_2656,N_2233);
or U5736 (N_5736,N_1672,N_1979);
or U5737 (N_5737,N_357,N_808);
or U5738 (N_5738,N_454,N_1367);
nor U5739 (N_5739,N_1181,N_2130);
nand U5740 (N_5740,N_319,N_1961);
or U5741 (N_5741,N_2521,N_512);
or U5742 (N_5742,N_2715,N_884);
nand U5743 (N_5743,N_741,N_641);
xnor U5744 (N_5744,N_1074,N_1763);
nand U5745 (N_5745,N_2880,N_1584);
nand U5746 (N_5746,N_2404,N_1886);
or U5747 (N_5747,N_1088,N_576);
nand U5748 (N_5748,N_197,N_1092);
nand U5749 (N_5749,N_1729,N_2325);
nor U5750 (N_5750,N_422,N_847);
and U5751 (N_5751,N_2417,N_1650);
or U5752 (N_5752,N_462,N_2114);
nand U5753 (N_5753,N_2035,N_327);
xnor U5754 (N_5754,N_2187,N_729);
nand U5755 (N_5755,N_1424,N_129);
xor U5756 (N_5756,N_2190,N_1074);
nand U5757 (N_5757,N_1098,N_2752);
and U5758 (N_5758,N_1633,N_2191);
xor U5759 (N_5759,N_2401,N_599);
xor U5760 (N_5760,N_1781,N_895);
xor U5761 (N_5761,N_2085,N_1284);
xor U5762 (N_5762,N_2748,N_1530);
and U5763 (N_5763,N_1646,N_2172);
nor U5764 (N_5764,N_439,N_2751);
or U5765 (N_5765,N_956,N_1516);
and U5766 (N_5766,N_1931,N_1569);
and U5767 (N_5767,N_2822,N_2195);
xor U5768 (N_5768,N_869,N_1492);
xnor U5769 (N_5769,N_478,N_1856);
and U5770 (N_5770,N_2653,N_2906);
and U5771 (N_5771,N_2836,N_1238);
or U5772 (N_5772,N_1075,N_417);
nand U5773 (N_5773,N_616,N_1378);
and U5774 (N_5774,N_2796,N_1391);
nor U5775 (N_5775,N_2588,N_635);
and U5776 (N_5776,N_1971,N_1964);
nor U5777 (N_5777,N_2550,N_189);
xnor U5778 (N_5778,N_558,N_345);
or U5779 (N_5779,N_1749,N_1853);
or U5780 (N_5780,N_2992,N_1395);
and U5781 (N_5781,N_1653,N_551);
or U5782 (N_5782,N_1017,N_830);
nor U5783 (N_5783,N_157,N_79);
nand U5784 (N_5784,N_544,N_2542);
or U5785 (N_5785,N_2767,N_601);
nand U5786 (N_5786,N_2333,N_765);
xor U5787 (N_5787,N_2366,N_904);
nand U5788 (N_5788,N_1552,N_539);
or U5789 (N_5789,N_213,N_1341);
nand U5790 (N_5790,N_1288,N_1088);
nand U5791 (N_5791,N_1347,N_2906);
nor U5792 (N_5792,N_653,N_1008);
nand U5793 (N_5793,N_2349,N_1102);
xnor U5794 (N_5794,N_2584,N_959);
xor U5795 (N_5795,N_2709,N_41);
or U5796 (N_5796,N_1117,N_701);
and U5797 (N_5797,N_928,N_275);
and U5798 (N_5798,N_185,N_1563);
nor U5799 (N_5799,N_2256,N_347);
xor U5800 (N_5800,N_2044,N_2148);
and U5801 (N_5801,N_1889,N_2036);
and U5802 (N_5802,N_457,N_1939);
and U5803 (N_5803,N_1234,N_603);
nor U5804 (N_5804,N_1600,N_2801);
or U5805 (N_5805,N_1570,N_1091);
nor U5806 (N_5806,N_874,N_14);
nor U5807 (N_5807,N_584,N_2468);
or U5808 (N_5808,N_1743,N_2545);
xnor U5809 (N_5809,N_2345,N_281);
and U5810 (N_5810,N_430,N_2657);
nand U5811 (N_5811,N_632,N_1698);
and U5812 (N_5812,N_547,N_2985);
and U5813 (N_5813,N_876,N_2578);
xor U5814 (N_5814,N_1853,N_34);
nand U5815 (N_5815,N_2227,N_816);
xor U5816 (N_5816,N_45,N_1920);
nand U5817 (N_5817,N_1785,N_1750);
or U5818 (N_5818,N_1082,N_923);
and U5819 (N_5819,N_1742,N_1390);
xor U5820 (N_5820,N_11,N_2650);
nor U5821 (N_5821,N_920,N_1239);
and U5822 (N_5822,N_1885,N_184);
xor U5823 (N_5823,N_984,N_1780);
nor U5824 (N_5824,N_1893,N_1976);
xnor U5825 (N_5825,N_1338,N_2462);
nor U5826 (N_5826,N_2525,N_1882);
nor U5827 (N_5827,N_1674,N_229);
and U5828 (N_5828,N_1586,N_453);
and U5829 (N_5829,N_2911,N_1001);
nor U5830 (N_5830,N_1853,N_504);
and U5831 (N_5831,N_995,N_291);
nor U5832 (N_5832,N_718,N_2471);
xnor U5833 (N_5833,N_2095,N_1195);
xor U5834 (N_5834,N_1777,N_2613);
nand U5835 (N_5835,N_1283,N_1873);
nor U5836 (N_5836,N_2028,N_1573);
nor U5837 (N_5837,N_229,N_71);
and U5838 (N_5838,N_1111,N_2671);
or U5839 (N_5839,N_2253,N_2879);
nand U5840 (N_5840,N_410,N_937);
xnor U5841 (N_5841,N_485,N_1578);
nor U5842 (N_5842,N_2607,N_2803);
or U5843 (N_5843,N_1435,N_2926);
nor U5844 (N_5844,N_2969,N_992);
nor U5845 (N_5845,N_2934,N_1962);
or U5846 (N_5846,N_133,N_458);
or U5847 (N_5847,N_2371,N_1128);
xnor U5848 (N_5848,N_1284,N_2860);
nand U5849 (N_5849,N_2822,N_1777);
xor U5850 (N_5850,N_1013,N_453);
or U5851 (N_5851,N_987,N_2716);
and U5852 (N_5852,N_866,N_2016);
nor U5853 (N_5853,N_451,N_2042);
nand U5854 (N_5854,N_1492,N_535);
xnor U5855 (N_5855,N_1127,N_0);
xnor U5856 (N_5856,N_2816,N_178);
xor U5857 (N_5857,N_1039,N_1235);
nor U5858 (N_5858,N_1403,N_2830);
and U5859 (N_5859,N_2459,N_814);
or U5860 (N_5860,N_1672,N_470);
and U5861 (N_5861,N_1967,N_1512);
and U5862 (N_5862,N_1025,N_1820);
xnor U5863 (N_5863,N_1136,N_2025);
and U5864 (N_5864,N_2248,N_2534);
and U5865 (N_5865,N_994,N_1447);
or U5866 (N_5866,N_1476,N_1148);
nor U5867 (N_5867,N_2106,N_737);
nand U5868 (N_5868,N_267,N_299);
and U5869 (N_5869,N_1659,N_590);
xor U5870 (N_5870,N_1811,N_1117);
and U5871 (N_5871,N_214,N_984);
nand U5872 (N_5872,N_2937,N_1926);
xor U5873 (N_5873,N_586,N_368);
or U5874 (N_5874,N_1801,N_312);
nor U5875 (N_5875,N_382,N_1690);
nand U5876 (N_5876,N_1282,N_2882);
or U5877 (N_5877,N_2136,N_323);
and U5878 (N_5878,N_1683,N_493);
nor U5879 (N_5879,N_2894,N_1488);
and U5880 (N_5880,N_771,N_266);
nand U5881 (N_5881,N_650,N_2712);
nand U5882 (N_5882,N_1824,N_446);
xor U5883 (N_5883,N_242,N_2044);
or U5884 (N_5884,N_430,N_816);
or U5885 (N_5885,N_1696,N_2661);
xnor U5886 (N_5886,N_1345,N_419);
xor U5887 (N_5887,N_37,N_1283);
or U5888 (N_5888,N_440,N_2828);
nor U5889 (N_5889,N_956,N_1959);
nor U5890 (N_5890,N_1425,N_675);
nand U5891 (N_5891,N_981,N_2204);
xnor U5892 (N_5892,N_2106,N_1891);
nand U5893 (N_5893,N_2090,N_1795);
nand U5894 (N_5894,N_2829,N_2273);
nand U5895 (N_5895,N_870,N_2102);
or U5896 (N_5896,N_214,N_2850);
nor U5897 (N_5897,N_1509,N_2696);
or U5898 (N_5898,N_2283,N_724);
nor U5899 (N_5899,N_963,N_298);
nand U5900 (N_5900,N_1320,N_1261);
nor U5901 (N_5901,N_268,N_2561);
xor U5902 (N_5902,N_2319,N_2048);
nor U5903 (N_5903,N_766,N_1819);
and U5904 (N_5904,N_527,N_1404);
and U5905 (N_5905,N_2888,N_833);
nor U5906 (N_5906,N_2791,N_1621);
and U5907 (N_5907,N_1990,N_1789);
or U5908 (N_5908,N_266,N_2254);
nor U5909 (N_5909,N_1461,N_668);
xnor U5910 (N_5910,N_23,N_2463);
and U5911 (N_5911,N_2057,N_527);
nand U5912 (N_5912,N_2616,N_2232);
or U5913 (N_5913,N_2783,N_2983);
xor U5914 (N_5914,N_1145,N_2133);
nor U5915 (N_5915,N_886,N_1843);
nand U5916 (N_5916,N_353,N_1909);
nand U5917 (N_5917,N_1819,N_2904);
and U5918 (N_5918,N_970,N_2292);
or U5919 (N_5919,N_858,N_1682);
nor U5920 (N_5920,N_1529,N_366);
nor U5921 (N_5921,N_1397,N_584);
xnor U5922 (N_5922,N_2794,N_1166);
or U5923 (N_5923,N_1407,N_1095);
nand U5924 (N_5924,N_2640,N_1940);
and U5925 (N_5925,N_1565,N_2459);
nor U5926 (N_5926,N_680,N_1061);
nand U5927 (N_5927,N_410,N_1636);
xnor U5928 (N_5928,N_1281,N_2864);
xnor U5929 (N_5929,N_1370,N_2009);
xor U5930 (N_5930,N_1293,N_1749);
and U5931 (N_5931,N_2353,N_736);
nor U5932 (N_5932,N_1726,N_1512);
nand U5933 (N_5933,N_107,N_2469);
xnor U5934 (N_5934,N_2628,N_1328);
nor U5935 (N_5935,N_1593,N_1238);
or U5936 (N_5936,N_1258,N_271);
xnor U5937 (N_5937,N_1299,N_420);
nor U5938 (N_5938,N_68,N_543);
nand U5939 (N_5939,N_1605,N_2951);
nand U5940 (N_5940,N_2956,N_2004);
or U5941 (N_5941,N_1420,N_310);
nand U5942 (N_5942,N_528,N_1842);
or U5943 (N_5943,N_1422,N_1591);
xnor U5944 (N_5944,N_556,N_60);
nor U5945 (N_5945,N_360,N_752);
nand U5946 (N_5946,N_1395,N_1604);
nand U5947 (N_5947,N_1348,N_2370);
nor U5948 (N_5948,N_526,N_1697);
and U5949 (N_5949,N_2760,N_2553);
or U5950 (N_5950,N_1727,N_1145);
nand U5951 (N_5951,N_2941,N_1921);
and U5952 (N_5952,N_261,N_1898);
xnor U5953 (N_5953,N_313,N_786);
nand U5954 (N_5954,N_1109,N_1562);
nand U5955 (N_5955,N_1658,N_2613);
nand U5956 (N_5956,N_1343,N_2815);
or U5957 (N_5957,N_964,N_2113);
xnor U5958 (N_5958,N_2319,N_2346);
and U5959 (N_5959,N_2899,N_31);
and U5960 (N_5960,N_811,N_1954);
and U5961 (N_5961,N_2970,N_1941);
xnor U5962 (N_5962,N_866,N_2385);
nand U5963 (N_5963,N_1934,N_1778);
and U5964 (N_5964,N_2256,N_1790);
nand U5965 (N_5965,N_992,N_672);
and U5966 (N_5966,N_660,N_2522);
nor U5967 (N_5967,N_1135,N_244);
and U5968 (N_5968,N_1411,N_313);
and U5969 (N_5969,N_2020,N_2285);
xnor U5970 (N_5970,N_55,N_1119);
and U5971 (N_5971,N_2588,N_1996);
xnor U5972 (N_5972,N_82,N_60);
xor U5973 (N_5973,N_2993,N_473);
nand U5974 (N_5974,N_1584,N_582);
and U5975 (N_5975,N_2004,N_988);
xnor U5976 (N_5976,N_175,N_195);
nor U5977 (N_5977,N_2768,N_984);
and U5978 (N_5978,N_2696,N_705);
and U5979 (N_5979,N_758,N_2928);
and U5980 (N_5980,N_51,N_2827);
and U5981 (N_5981,N_2768,N_2839);
nor U5982 (N_5982,N_1076,N_1834);
or U5983 (N_5983,N_2145,N_1812);
or U5984 (N_5984,N_2916,N_159);
nand U5985 (N_5985,N_1990,N_2564);
nand U5986 (N_5986,N_1355,N_408);
or U5987 (N_5987,N_863,N_2989);
and U5988 (N_5988,N_2199,N_399);
and U5989 (N_5989,N_193,N_2921);
xor U5990 (N_5990,N_1011,N_788);
or U5991 (N_5991,N_2445,N_1602);
or U5992 (N_5992,N_639,N_587);
nor U5993 (N_5993,N_2826,N_664);
nand U5994 (N_5994,N_1941,N_800);
and U5995 (N_5995,N_2939,N_194);
nand U5996 (N_5996,N_767,N_714);
nor U5997 (N_5997,N_2358,N_359);
and U5998 (N_5998,N_2882,N_2191);
nor U5999 (N_5999,N_1426,N_858);
xnor U6000 (N_6000,N_5073,N_3352);
or U6001 (N_6001,N_4284,N_3620);
nor U6002 (N_6002,N_3051,N_3408);
xor U6003 (N_6003,N_5920,N_4438);
or U6004 (N_6004,N_4901,N_3237);
nand U6005 (N_6005,N_5468,N_4541);
and U6006 (N_6006,N_5118,N_4013);
or U6007 (N_6007,N_5200,N_3245);
xor U6008 (N_6008,N_4372,N_3359);
nor U6009 (N_6009,N_5836,N_5159);
or U6010 (N_6010,N_4976,N_5615);
and U6011 (N_6011,N_4293,N_3785);
nor U6012 (N_6012,N_5804,N_4998);
xnor U6013 (N_6013,N_5488,N_3626);
nor U6014 (N_6014,N_4895,N_4965);
and U6015 (N_6015,N_5373,N_3697);
and U6016 (N_6016,N_5524,N_5346);
nor U6017 (N_6017,N_3947,N_4913);
and U6018 (N_6018,N_4511,N_5393);
and U6019 (N_6019,N_4548,N_3740);
xor U6020 (N_6020,N_5193,N_5039);
xnor U6021 (N_6021,N_5639,N_5873);
and U6022 (N_6022,N_4409,N_5883);
nor U6023 (N_6023,N_5376,N_4297);
nand U6024 (N_6024,N_3759,N_3341);
or U6025 (N_6025,N_5948,N_5640);
xor U6026 (N_6026,N_5495,N_4498);
nand U6027 (N_6027,N_3707,N_5568);
xor U6028 (N_6028,N_5945,N_5909);
or U6029 (N_6029,N_5380,N_5561);
or U6030 (N_6030,N_3095,N_5983);
or U6031 (N_6031,N_4380,N_3046);
nand U6032 (N_6032,N_5294,N_4116);
or U6033 (N_6033,N_4620,N_4054);
and U6034 (N_6034,N_3519,N_3601);
or U6035 (N_6035,N_4042,N_3239);
and U6036 (N_6036,N_4786,N_3331);
xnor U6037 (N_6037,N_3528,N_5835);
nand U6038 (N_6038,N_5768,N_5086);
and U6039 (N_6039,N_5274,N_4279);
xnor U6040 (N_6040,N_3869,N_3549);
and U6041 (N_6041,N_3579,N_3985);
xor U6042 (N_6042,N_3884,N_4303);
and U6043 (N_6043,N_4450,N_3992);
xnor U6044 (N_6044,N_3373,N_3060);
and U6045 (N_6045,N_4322,N_3290);
nor U6046 (N_6046,N_4345,N_3039);
and U6047 (N_6047,N_5046,N_5537);
and U6048 (N_6048,N_4684,N_5175);
xor U6049 (N_6049,N_4257,N_5272);
nand U6050 (N_6050,N_5656,N_4654);
and U6051 (N_6051,N_4236,N_4416);
nand U6052 (N_6052,N_4018,N_3205);
or U6053 (N_6053,N_4449,N_3372);
and U6054 (N_6054,N_4627,N_5044);
or U6055 (N_6055,N_3847,N_4275);
xor U6056 (N_6056,N_3763,N_4085);
nor U6057 (N_6057,N_5192,N_3996);
nand U6058 (N_6058,N_4102,N_3030);
or U6059 (N_6059,N_5383,N_4748);
xnor U6060 (N_6060,N_4983,N_3649);
or U6061 (N_6061,N_4943,N_4609);
or U6062 (N_6062,N_3045,N_5223);
or U6063 (N_6063,N_5788,N_5989);
and U6064 (N_6064,N_4166,N_4785);
and U6065 (N_6065,N_4183,N_5459);
xor U6066 (N_6066,N_5312,N_5542);
or U6067 (N_6067,N_4945,N_5300);
nand U6068 (N_6068,N_4958,N_3991);
xor U6069 (N_6069,N_3930,N_3210);
nor U6070 (N_6070,N_3508,N_3221);
or U6071 (N_6071,N_5752,N_4132);
xor U6072 (N_6072,N_5152,N_4235);
and U6073 (N_6073,N_4766,N_3833);
and U6074 (N_6074,N_3881,N_3880);
or U6075 (N_6075,N_5766,N_3470);
or U6076 (N_6076,N_3185,N_3106);
nand U6077 (N_6077,N_5941,N_3075);
and U6078 (N_6078,N_4792,N_3453);
and U6079 (N_6079,N_3204,N_5924);
nand U6080 (N_6080,N_5437,N_3107);
xor U6081 (N_6081,N_5614,N_4872);
or U6082 (N_6082,N_5314,N_4103);
and U6083 (N_6083,N_5151,N_4064);
and U6084 (N_6084,N_4725,N_5647);
xor U6085 (N_6085,N_5458,N_4544);
and U6086 (N_6086,N_5114,N_4014);
or U6087 (N_6087,N_4364,N_4573);
nor U6088 (N_6088,N_3547,N_5605);
and U6089 (N_6089,N_5792,N_4542);
and U6090 (N_6090,N_5101,N_5699);
xor U6091 (N_6091,N_5517,N_3003);
or U6092 (N_6092,N_3456,N_3268);
xnor U6093 (N_6093,N_3187,N_5023);
and U6094 (N_6094,N_3958,N_4815);
nand U6095 (N_6095,N_4986,N_4262);
nor U6096 (N_6096,N_5663,N_4837);
xnor U6097 (N_6097,N_5331,N_3180);
xor U6098 (N_6098,N_3317,N_3443);
or U6099 (N_6099,N_4436,N_5692);
and U6100 (N_6100,N_5953,N_4090);
or U6101 (N_6101,N_5230,N_5181);
or U6102 (N_6102,N_3417,N_5037);
xor U6103 (N_6103,N_5739,N_3010);
and U6104 (N_6104,N_4879,N_4862);
and U6105 (N_6105,N_4520,N_4070);
nand U6106 (N_6106,N_4291,N_3640);
nand U6107 (N_6107,N_4462,N_4509);
and U6108 (N_6108,N_4617,N_4966);
or U6109 (N_6109,N_5578,N_4367);
nor U6110 (N_6110,N_5079,N_3156);
nor U6111 (N_6111,N_3061,N_5560);
and U6112 (N_6112,N_5403,N_5619);
nor U6113 (N_6113,N_3147,N_3751);
nor U6114 (N_6114,N_5877,N_4636);
xor U6115 (N_6115,N_3770,N_4399);
nor U6116 (N_6116,N_3575,N_4497);
and U6117 (N_6117,N_3391,N_4144);
and U6118 (N_6118,N_4747,N_5706);
and U6119 (N_6119,N_5474,N_3594);
and U6120 (N_6120,N_5102,N_3335);
nor U6121 (N_6121,N_4063,N_4594);
and U6122 (N_6122,N_3843,N_3986);
and U6123 (N_6123,N_4124,N_3701);
nor U6124 (N_6124,N_4948,N_4935);
nand U6125 (N_6125,N_4782,N_3232);
and U6126 (N_6126,N_4962,N_4820);
xnor U6127 (N_6127,N_3710,N_3980);
xor U6128 (N_6128,N_5203,N_4570);
nand U6129 (N_6129,N_4665,N_3236);
and U6130 (N_6130,N_3186,N_4767);
nand U6131 (N_6131,N_3089,N_4553);
nand U6132 (N_6132,N_3747,N_5604);
nand U6133 (N_6133,N_4027,N_3734);
xor U6134 (N_6134,N_5533,N_4863);
xnor U6135 (N_6135,N_3840,N_5472);
nor U6136 (N_6136,N_3494,N_4675);
xnor U6137 (N_6137,N_4406,N_5617);
or U6138 (N_6138,N_4930,N_3586);
nor U6139 (N_6139,N_5007,N_5315);
and U6140 (N_6140,N_4667,N_3550);
nor U6141 (N_6141,N_5187,N_5477);
or U6142 (N_6142,N_5498,N_5387);
and U6143 (N_6143,N_5245,N_3954);
xor U6144 (N_6144,N_4316,N_5496);
nand U6145 (N_6145,N_5600,N_3536);
and U6146 (N_6146,N_4836,N_5796);
nor U6147 (N_6147,N_5462,N_4181);
or U6148 (N_6148,N_3149,N_4196);
nand U6149 (N_6149,N_3423,N_3824);
nor U6150 (N_6150,N_5642,N_5427);
and U6151 (N_6151,N_5370,N_3484);
nand U6152 (N_6152,N_5136,N_3800);
and U6153 (N_6153,N_5157,N_5842);
and U6154 (N_6154,N_3603,N_4469);
xor U6155 (N_6155,N_5287,N_4970);
nor U6156 (N_6156,N_5292,N_4692);
xnor U6157 (N_6157,N_4067,N_5205);
nand U6158 (N_6158,N_5077,N_3587);
nor U6159 (N_6159,N_3110,N_5407);
and U6160 (N_6160,N_5405,N_5504);
and U6161 (N_6161,N_4877,N_5662);
or U6162 (N_6162,N_5807,N_5497);
and U6163 (N_6163,N_3977,N_3076);
nor U6164 (N_6164,N_3247,N_3224);
nor U6165 (N_6165,N_5142,N_4414);
or U6166 (N_6166,N_3686,N_5627);
nor U6167 (N_6167,N_4957,N_3428);
xnor U6168 (N_6168,N_3452,N_5534);
or U6169 (N_6169,N_5961,N_3019);
xnor U6170 (N_6170,N_4152,N_5938);
nor U6171 (N_6171,N_3856,N_4677);
nor U6172 (N_6172,N_3558,N_3486);
and U6173 (N_6173,N_4404,N_4022);
xor U6174 (N_6174,N_4900,N_3404);
and U6175 (N_6175,N_5912,N_4269);
and U6176 (N_6176,N_5813,N_4905);
or U6177 (N_6177,N_4602,N_4478);
nor U6178 (N_6178,N_5893,N_4489);
nand U6179 (N_6179,N_3338,N_3875);
or U6180 (N_6180,N_4752,N_5279);
or U6181 (N_6181,N_5651,N_4659);
and U6182 (N_6182,N_3078,N_4390);
nand U6183 (N_6183,N_4306,N_5762);
or U6184 (N_6184,N_5124,N_5671);
xor U6185 (N_6185,N_5799,N_5816);
nand U6186 (N_6186,N_5456,N_3094);
nor U6187 (N_6187,N_4025,N_4530);
nand U6188 (N_6188,N_3301,N_4107);
and U6189 (N_6189,N_5969,N_3031);
and U6190 (N_6190,N_5153,N_5234);
or U6191 (N_6191,N_3731,N_4113);
or U6192 (N_6192,N_5525,N_5362);
nor U6193 (N_6193,N_4314,N_4330);
and U6194 (N_6194,N_3882,N_5580);
and U6195 (N_6195,N_5271,N_4337);
xnor U6196 (N_6196,N_3292,N_3804);
nor U6197 (N_6197,N_4444,N_4247);
nand U6198 (N_6198,N_3316,N_3278);
nand U6199 (N_6199,N_5252,N_4225);
and U6200 (N_6200,N_4805,N_3709);
nand U6201 (N_6201,N_4835,N_4685);
or U6202 (N_6202,N_4268,N_4410);
nand U6203 (N_6203,N_4202,N_4033);
nor U6204 (N_6204,N_3899,N_4683);
or U6205 (N_6205,N_5658,N_5839);
nor U6206 (N_6206,N_5539,N_3406);
and U6207 (N_6207,N_5997,N_3819);
xor U6208 (N_6208,N_3325,N_4179);
nor U6209 (N_6209,N_5216,N_5782);
or U6210 (N_6210,N_3636,N_5821);
xnor U6211 (N_6211,N_3023,N_5531);
nor U6212 (N_6212,N_3801,N_4177);
or U6213 (N_6213,N_4535,N_4673);
nor U6214 (N_6214,N_3664,N_4439);
nand U6215 (N_6215,N_4645,N_5161);
or U6216 (N_6216,N_5618,N_3546);
nand U6217 (N_6217,N_3018,N_5991);
and U6218 (N_6218,N_4583,N_4080);
xor U6219 (N_6219,N_5475,N_3157);
nand U6220 (N_6220,N_3438,N_3191);
nand U6221 (N_6221,N_3643,N_5527);
xnor U6222 (N_6222,N_3002,N_3016);
nand U6223 (N_6223,N_5235,N_5392);
xnor U6224 (N_6224,N_5061,N_3449);
or U6225 (N_6225,N_4007,N_3355);
nand U6226 (N_6226,N_4593,N_5625);
nand U6227 (N_6227,N_3468,N_4119);
nand U6228 (N_6228,N_5590,N_5484);
or U6229 (N_6229,N_3296,N_4058);
nand U6230 (N_6230,N_3291,N_3534);
xor U6231 (N_6231,N_5691,N_5278);
and U6232 (N_6232,N_4256,N_4759);
nand U6233 (N_6233,N_4203,N_3678);
nor U6234 (N_6234,N_3950,N_3207);
and U6235 (N_6235,N_5931,N_3451);
nand U6236 (N_6236,N_5188,N_5648);
or U6237 (N_6237,N_5875,N_3313);
nand U6238 (N_6238,N_3118,N_3457);
or U6239 (N_6239,N_5176,N_3483);
nor U6240 (N_6240,N_4971,N_5812);
and U6241 (N_6241,N_3320,N_4440);
nor U6242 (N_6242,N_4849,N_4607);
xor U6243 (N_6243,N_4916,N_3615);
nand U6244 (N_6244,N_5958,N_4569);
and U6245 (N_6245,N_3112,N_5646);
nand U6246 (N_6246,N_3065,N_5431);
nor U6247 (N_6247,N_3403,N_5838);
xor U6248 (N_6248,N_5038,N_5017);
or U6249 (N_6249,N_4694,N_4138);
xnor U6250 (N_6250,N_3786,N_5322);
nor U6251 (N_6251,N_5112,N_5927);
nand U6252 (N_6252,N_5825,N_4017);
nand U6253 (N_6253,N_5872,N_4960);
nand U6254 (N_6254,N_4549,N_4892);
xor U6255 (N_6255,N_3396,N_4338);
and U6256 (N_6256,N_3848,N_4407);
nor U6257 (N_6257,N_5045,N_3746);
nand U6258 (N_6258,N_3211,N_5256);
or U6259 (N_6259,N_3934,N_5012);
nand U6260 (N_6260,N_3101,N_3995);
and U6261 (N_6261,N_5638,N_5361);
nor U6262 (N_6262,N_5858,N_5607);
nand U6263 (N_6263,N_4969,N_4245);
nand U6264 (N_6264,N_3253,N_5328);
nor U6265 (N_6265,N_3412,N_4205);
or U6266 (N_6266,N_5928,N_3755);
or U6267 (N_6267,N_3913,N_3151);
nor U6268 (N_6268,N_4655,N_4742);
and U6269 (N_6269,N_5404,N_5180);
or U6270 (N_6270,N_5819,N_4105);
or U6271 (N_6271,N_4369,N_4799);
nand U6272 (N_6272,N_4526,N_3527);
xnor U6273 (N_6273,N_4072,N_4461);
and U6274 (N_6274,N_5913,N_5158);
nand U6275 (N_6275,N_3197,N_4046);
and U6276 (N_6276,N_3498,N_4674);
nand U6277 (N_6277,N_3038,N_4158);
nor U6278 (N_6278,N_5069,N_4903);
nor U6279 (N_6279,N_5528,N_4790);
nor U6280 (N_6280,N_5682,N_3572);
or U6281 (N_6281,N_3036,N_3700);
and U6282 (N_6282,N_3582,N_5727);
or U6283 (N_6283,N_4887,N_3892);
nand U6284 (N_6284,N_5464,N_3681);
xnor U6285 (N_6285,N_4512,N_3748);
and U6286 (N_6286,N_3784,N_3853);
xnor U6287 (N_6287,N_5417,N_3074);
nor U6288 (N_6288,N_4884,N_4395);
nand U6289 (N_6289,N_4130,N_4422);
and U6290 (N_6290,N_5240,N_4405);
nand U6291 (N_6291,N_4878,N_3596);
and U6292 (N_6292,N_4506,N_4468);
or U6293 (N_6293,N_4755,N_3032);
nand U6294 (N_6294,N_4104,N_3104);
or U6295 (N_6295,N_3024,N_4988);
or U6296 (N_6296,N_5492,N_4949);
and U6297 (N_6297,N_4953,N_4231);
xnor U6298 (N_6298,N_4811,N_3281);
xor U6299 (N_6299,N_4596,N_5641);
nor U6300 (N_6300,N_3657,N_4274);
nor U6301 (N_6301,N_3310,N_5447);
nor U6302 (N_6302,N_4324,N_4289);
nor U6303 (N_6303,N_4176,N_3192);
or U6304 (N_6304,N_3612,N_5402);
nand U6305 (N_6305,N_5441,N_4037);
xnor U6306 (N_6306,N_4795,N_5676);
and U6307 (N_6307,N_5206,N_4097);
or U6308 (N_6308,N_5080,N_3822);
xnor U6309 (N_6309,N_3165,N_4501);
and U6310 (N_6310,N_4827,N_3960);
nor U6311 (N_6311,N_3295,N_3783);
and U6312 (N_6312,N_5649,N_4198);
or U6313 (N_6313,N_5967,N_5643);
and U6314 (N_6314,N_3602,N_5954);
or U6315 (N_6315,N_4313,N_4554);
xnor U6316 (N_6316,N_3902,N_4224);
nor U6317 (N_6317,N_3863,N_5702);
nand U6318 (N_6318,N_5384,N_3390);
and U6319 (N_6319,N_5522,N_4030);
xor U6320 (N_6320,N_5942,N_3234);
nor U6321 (N_6321,N_3490,N_4540);
nand U6322 (N_6322,N_4999,N_5144);
nand U6323 (N_6323,N_5532,N_4494);
nor U6324 (N_6324,N_4215,N_5876);
or U6325 (N_6325,N_3047,N_3727);
nor U6326 (N_6326,N_4516,N_4719);
nor U6327 (N_6327,N_5668,N_4121);
nor U6328 (N_6328,N_4031,N_5805);
xnor U6329 (N_6329,N_4629,N_3266);
nor U6330 (N_6330,N_5921,N_4458);
or U6331 (N_6331,N_4239,N_3179);
or U6332 (N_6332,N_4273,N_3589);
nor U6333 (N_6333,N_3922,N_5587);
nor U6334 (N_6334,N_4959,N_4349);
nand U6335 (N_6335,N_4601,N_4180);
or U6336 (N_6336,N_3702,N_5479);
nor U6337 (N_6337,N_5556,N_4632);
nand U6338 (N_6338,N_3982,N_5394);
or U6339 (N_6339,N_3148,N_5898);
nor U6340 (N_6340,N_3834,N_4034);
nand U6341 (N_6341,N_3956,N_3936);
and U6342 (N_6342,N_3441,N_4652);
nand U6343 (N_6343,N_3063,N_4242);
nor U6344 (N_6344,N_5520,N_3427);
or U6345 (N_6345,N_3668,N_3172);
and U6346 (N_6346,N_5994,N_5555);
or U6347 (N_6347,N_5806,N_3749);
and U6348 (N_6348,N_4760,N_3979);
and U6349 (N_6349,N_4928,N_4550);
xnor U6350 (N_6350,N_5139,N_4984);
nor U6351 (N_6351,N_4477,N_4933);
or U6352 (N_6352,N_3425,N_5963);
nor U6353 (N_6353,N_4266,N_5845);
xor U6354 (N_6354,N_5189,N_5490);
and U6355 (N_6355,N_3113,N_5451);
nand U6356 (N_6356,N_5117,N_5264);
nand U6357 (N_6357,N_5540,N_3916);
or U6358 (N_6358,N_4049,N_5878);
xor U6359 (N_6359,N_5770,N_3208);
xnor U6360 (N_6360,N_4388,N_3041);
nand U6361 (N_6361,N_4157,N_4931);
or U6362 (N_6362,N_3369,N_5209);
nand U6363 (N_6363,N_4211,N_4006);
and U6364 (N_6364,N_4163,N_4137);
nand U6365 (N_6365,N_4623,N_3908);
xnor U6366 (N_6366,N_5977,N_4408);
or U6367 (N_6367,N_3017,N_5436);
and U6368 (N_6368,N_5422,N_4889);
xor U6369 (N_6369,N_4897,N_5065);
or U6370 (N_6370,N_3272,N_5814);
or U6371 (N_6371,N_5514,N_4092);
xor U6372 (N_6372,N_4704,N_3007);
nor U6373 (N_6373,N_5946,N_5390);
and U6374 (N_6374,N_4243,N_3931);
and U6375 (N_6375,N_5843,N_4234);
nor U6376 (N_6376,N_4834,N_4226);
xor U6377 (N_6377,N_3628,N_3103);
nand U6378 (N_6378,N_3915,N_5107);
and U6379 (N_6379,N_5013,N_5062);
and U6380 (N_6380,N_4078,N_5182);
xnor U6381 (N_6381,N_4964,N_3919);
nor U6382 (N_6382,N_4083,N_3816);
xor U6383 (N_6383,N_4634,N_4093);
or U6384 (N_6384,N_4740,N_3791);
nand U6385 (N_6385,N_4465,N_3001);
nand U6386 (N_6386,N_5460,N_4723);
and U6387 (N_6387,N_4145,N_5529);
or U6388 (N_6388,N_4383,N_3326);
or U6389 (N_6389,N_3170,N_3924);
and U6390 (N_6390,N_5134,N_4387);
xnor U6391 (N_6391,N_5184,N_5866);
nand U6392 (N_6392,N_4429,N_5071);
nand U6393 (N_6393,N_5267,N_5583);
and U6394 (N_6394,N_3263,N_3070);
nor U6395 (N_6395,N_4304,N_4587);
nand U6396 (N_6396,N_4076,N_3242);
or U6397 (N_6397,N_4902,N_4951);
nand U6398 (N_6398,N_5712,N_4802);
nand U6399 (N_6399,N_3651,N_5521);
nor U6400 (N_6400,N_5434,N_3943);
nor U6401 (N_6401,N_3855,N_5650);
or U6402 (N_6402,N_3466,N_5844);
and U6403 (N_6403,N_3903,N_5338);
or U6404 (N_6404,N_3767,N_4908);
or U6405 (N_6405,N_5756,N_4323);
and U6406 (N_6406,N_4051,N_5754);
and U6407 (N_6407,N_5341,N_4420);
and U6408 (N_6408,N_3136,N_5775);
or U6409 (N_6409,N_3507,N_3781);
xor U6410 (N_6410,N_5409,N_3006);
and U6411 (N_6411,N_5541,N_4442);
or U6412 (N_6412,N_5690,N_4010);
or U6413 (N_6413,N_3190,N_4564);
and U6414 (N_6414,N_4963,N_5289);
or U6415 (N_6415,N_4567,N_5760);
xnor U6416 (N_6416,N_3214,N_5137);
xnor U6417 (N_6417,N_5675,N_3225);
nor U6418 (N_6418,N_5949,N_3079);
xnor U6419 (N_6419,N_5115,N_4170);
or U6420 (N_6420,N_5143,N_5667);
and U6421 (N_6421,N_4578,N_3715);
nand U6422 (N_6422,N_3968,N_5075);
or U6423 (N_6423,N_5904,N_4821);
nor U6424 (N_6424,N_4187,N_5466);
or U6425 (N_6425,N_3322,N_4074);
nor U6426 (N_6426,N_3358,N_3203);
nand U6427 (N_6427,N_5979,N_5244);
nor U6428 (N_6428,N_3220,N_4808);
nand U6429 (N_6429,N_3200,N_4362);
xor U6430 (N_6430,N_3111,N_3917);
or U6431 (N_6431,N_3393,N_5592);
nand U6432 (N_6432,N_4689,N_4475);
xor U6433 (N_6433,N_3872,N_4508);
nor U6434 (N_6434,N_4996,N_4890);
xor U6435 (N_6435,N_4730,N_5558);
and U6436 (N_6436,N_3551,N_4668);
or U6437 (N_6437,N_5616,N_4381);
xnor U6438 (N_6438,N_5793,N_5377);
nand U6439 (N_6439,N_5902,N_5040);
xnor U6440 (N_6440,N_4956,N_5598);
nor U6441 (N_6441,N_4700,N_5713);
or U6442 (N_6442,N_5703,N_4947);
or U6443 (N_6443,N_4411,N_5396);
and U6444 (N_6444,N_4112,N_5442);
nand U6445 (N_6445,N_4237,N_4894);
or U6446 (N_6446,N_4087,N_3108);
and U6447 (N_6447,N_3472,N_4041);
xnor U6448 (N_6448,N_3436,N_5930);
xor U6449 (N_6449,N_4114,N_4864);
xnor U6450 (N_6450,N_5631,N_5119);
xnor U6451 (N_6451,N_3100,N_3067);
or U6452 (N_6452,N_3037,N_5781);
or U6453 (N_6453,N_3841,N_5571);
nor U6454 (N_6454,N_4705,N_3548);
xnor U6455 (N_6455,N_4218,N_5848);
or U6456 (N_6456,N_4117,N_5608);
nor U6457 (N_6457,N_3416,N_4100);
nor U6458 (N_6458,N_4208,N_5000);
xor U6459 (N_6459,N_3518,N_5601);
or U6460 (N_6460,N_3512,N_3769);
xor U6461 (N_6461,N_5030,N_5779);
nor U6462 (N_6462,N_3418,N_4670);
nand U6463 (N_6463,N_5185,N_5413);
and U6464 (N_6464,N_3084,N_3474);
and U6465 (N_6465,N_5014,N_5988);
nand U6466 (N_6466,N_5741,N_4443);
and U6467 (N_6467,N_4662,N_5365);
xor U6468 (N_6468,N_3162,N_5829);
nor U6469 (N_6469,N_5318,N_5258);
nand U6470 (N_6470,N_4246,N_3836);
nand U6471 (N_6471,N_4459,N_4733);
or U6472 (N_6472,N_4360,N_3228);
and U6473 (N_6473,N_4728,N_3181);
or U6474 (N_6474,N_3144,N_5585);
xnor U6475 (N_6475,N_5678,N_4784);
nand U6476 (N_6476,N_3666,N_3267);
xor U6477 (N_6477,N_3957,N_3249);
nor U6478 (N_6478,N_5333,N_4818);
nor U6479 (N_6479,N_5074,N_3570);
nand U6480 (N_6480,N_5432,N_3539);
xnor U6481 (N_6481,N_5262,N_3500);
and U6482 (N_6482,N_3175,N_4914);
nand U6483 (N_6483,N_3631,N_3085);
xnor U6484 (N_6484,N_5374,N_4467);
xnor U6485 (N_6485,N_4630,N_4804);
or U6486 (N_6486,N_5603,N_3794);
nand U6487 (N_6487,N_3565,N_3661);
nand U6488 (N_6488,N_5636,N_5265);
nor U6489 (N_6489,N_5281,N_4371);
nand U6490 (N_6490,N_4826,N_3497);
or U6491 (N_6491,N_4968,N_3034);
nand U6492 (N_6492,N_5550,N_5826);
or U6493 (N_6493,N_5769,N_3944);
nor U6494 (N_6494,N_3566,N_3901);
nand U6495 (N_6495,N_5502,N_5697);
xnor U6496 (N_6496,N_4355,N_5305);
or U6497 (N_6497,N_4529,N_4403);
nor U6498 (N_6498,N_5146,N_4590);
nor U6499 (N_6499,N_3167,N_5553);
or U6500 (N_6500,N_5049,N_5063);
nor U6501 (N_6501,N_5131,N_4745);
and U6502 (N_6502,N_3904,N_5709);
nor U6503 (N_6503,N_4536,N_5421);
or U6504 (N_6504,N_3998,N_3387);
and U6505 (N_6505,N_5364,N_3860);
nor U6506 (N_6506,N_3685,N_5299);
xor U6507 (N_6507,N_4643,N_5693);
nor U6508 (N_6508,N_3694,N_5950);
nand U6509 (N_6509,N_4612,N_3910);
nand U6510 (N_6510,N_5728,N_5068);
and U6511 (N_6511,N_5784,N_5113);
xnor U6512 (N_6512,N_3202,N_5059);
or U6513 (N_6513,N_4946,N_3758);
nor U6514 (N_6514,N_5724,N_5174);
or U6515 (N_6515,N_3049,N_5066);
xnor U6516 (N_6516,N_5211,N_4184);
nor U6517 (N_6517,N_3849,N_3015);
or U6518 (N_6518,N_3057,N_3231);
nand U6519 (N_6519,N_4796,N_3496);
xnor U6520 (N_6520,N_3655,N_3343);
nor U6521 (N_6521,N_4057,N_3102);
and U6522 (N_6522,N_3690,N_3845);
xnor U6523 (N_6523,N_3544,N_4800);
nand U6524 (N_6524,N_3614,N_5672);
or U6525 (N_6525,N_4173,N_5551);
or U6526 (N_6526,N_3832,N_4357);
or U6527 (N_6527,N_3611,N_4389);
or U6528 (N_6528,N_3091,N_3271);
nor U6529 (N_6529,N_5135,N_3595);
nand U6530 (N_6530,N_4265,N_5500);
or U6531 (N_6531,N_5242,N_5797);
xor U6532 (N_6532,N_3096,N_3305);
nor U6533 (N_6533,N_5406,N_4418);
or U6534 (N_6534,N_3618,N_5172);
nand U6535 (N_6535,N_4190,N_5298);
nand U6536 (N_6536,N_3773,N_5395);
xor U6537 (N_6537,N_4712,N_3487);
or U6538 (N_6538,N_4695,N_4744);
and U6539 (N_6539,N_5019,N_5029);
nand U6540 (N_6540,N_3725,N_4891);
nand U6541 (N_6541,N_3262,N_5116);
nor U6542 (N_6542,N_3932,N_4146);
or U6543 (N_6543,N_3409,N_5738);
nand U6544 (N_6544,N_5864,N_5818);
and U6545 (N_6545,N_4451,N_4004);
nand U6546 (N_6546,N_3571,N_4286);
nand U6547 (N_6547,N_3921,N_5778);
nand U6548 (N_6548,N_5681,N_5508);
nor U6549 (N_6549,N_3376,N_4545);
and U6550 (N_6550,N_4702,N_5461);
xnor U6551 (N_6551,N_4504,N_5018);
xnor U6552 (N_6552,N_3647,N_5218);
xnor U6553 (N_6553,N_5236,N_4869);
nand U6554 (N_6554,N_3460,N_5670);
or U6555 (N_6555,N_3196,N_4731);
and U6556 (N_6556,N_3703,N_4774);
and U6557 (N_6557,N_3173,N_3644);
nand U6558 (N_6558,N_5347,N_4206);
or U6559 (N_6559,N_3117,N_4071);
nor U6560 (N_6560,N_3795,N_5133);
nor U6561 (N_6561,N_3780,N_4868);
nor U6562 (N_6562,N_3233,N_4794);
xnor U6563 (N_6563,N_5710,N_4729);
nand U6564 (N_6564,N_3432,N_4164);
or U6565 (N_6565,N_5493,N_3386);
nand U6566 (N_6566,N_4756,N_3392);
nor U6567 (N_6567,N_3625,N_5170);
nor U6568 (N_6568,N_3227,N_4264);
nand U6569 (N_6569,N_4336,N_3098);
and U6570 (N_6570,N_3777,N_4688);
nand U6571 (N_6571,N_5789,N_3064);
nand U6572 (N_6572,N_5820,N_5567);
xnor U6573 (N_6573,N_5195,N_3068);
xnor U6574 (N_6574,N_5856,N_5263);
xnor U6575 (N_6575,N_3624,N_3887);
nor U6576 (N_6576,N_4954,N_5357);
nand U6577 (N_6577,N_5048,N_3776);
nand U6578 (N_6578,N_4650,N_3820);
xor U6579 (N_6579,N_3653,N_5290);
nand U6580 (N_6580,N_4035,N_3733);
xnor U6581 (N_6581,N_4860,N_4793);
nand U6582 (N_6582,N_5226,N_3974);
or U6583 (N_6583,N_3435,N_4576);
or U6584 (N_6584,N_3194,N_3708);
or U6585 (N_6585,N_5968,N_4679);
and U6586 (N_6586,N_4479,N_4079);
nand U6587 (N_6587,N_3265,N_4277);
nor U6588 (N_6588,N_5773,N_5076);
xor U6589 (N_6589,N_3382,N_4492);
and U6590 (N_6590,N_5197,N_4505);
and U6591 (N_6591,N_3013,N_5090);
or U6592 (N_6592,N_4292,N_3479);
nor U6593 (N_6593,N_3364,N_5901);
and U6594 (N_6594,N_5121,N_3677);
nand U6595 (N_6595,N_4151,N_5725);
or U6596 (N_6596,N_3782,N_5885);
nor U6597 (N_6597,N_3370,N_3984);
and U6598 (N_6598,N_4481,N_3318);
nand U6599 (N_6599,N_4538,N_4191);
or U6600 (N_6600,N_3246,N_3803);
and U6601 (N_6601,N_4437,N_4642);
nand U6602 (N_6602,N_4178,N_3206);
xnor U6603 (N_6603,N_3183,N_3375);
xor U6604 (N_6604,N_3909,N_4379);
nor U6605 (N_6605,N_3599,N_3555);
nor U6606 (N_6606,N_4865,N_4348);
nor U6607 (N_6607,N_5148,N_4207);
or U6608 (N_6608,N_3878,N_5111);
and U6609 (N_6609,N_4354,N_3059);
nor U6610 (N_6610,N_3394,N_3461);
nor U6611 (N_6611,N_3588,N_5729);
nand U6612 (N_6612,N_3632,N_4561);
nand U6613 (N_6613,N_3867,N_3025);
nand U6614 (N_6614,N_4749,N_3948);
xor U6615 (N_6615,N_5060,N_5483);
and U6616 (N_6616,N_5323,N_5750);
and U6617 (N_6617,N_3426,N_4859);
xnor U6618 (N_6618,N_3699,N_5088);
xnor U6619 (N_6619,N_3961,N_3126);
nand U6620 (N_6620,N_4626,N_4344);
nor U6621 (N_6621,N_4391,N_4343);
nor U6622 (N_6622,N_5957,N_3040);
nand U6623 (N_6623,N_4171,N_3439);
and U6624 (N_6624,N_5548,N_4011);
or U6625 (N_6625,N_3941,N_5926);
nand U6626 (N_6626,N_3240,N_4882);
nand U6627 (N_6627,N_3116,N_3215);
or U6628 (N_6628,N_4474,N_3768);
nand U6629 (N_6629,N_4373,N_4640);
and U6630 (N_6630,N_5922,N_4932);
and U6631 (N_6631,N_4143,N_4664);
and U6632 (N_6632,N_5164,N_3385);
and U6633 (N_6633,N_3489,N_3750);
and U6634 (N_6634,N_4310,N_5002);
and U6635 (N_6635,N_5378,N_4193);
or U6636 (N_6636,N_5327,N_4555);
xor U6637 (N_6637,N_5385,N_5433);
or U6638 (N_6638,N_5330,N_3398);
nand U6639 (N_6639,N_4923,N_4994);
nand U6640 (N_6640,N_5399,N_3520);
and U6641 (N_6641,N_3714,N_3877);
nand U6642 (N_6642,N_5266,N_5943);
or U6643 (N_6643,N_3303,N_4096);
nand U6644 (N_6644,N_3168,N_4830);
nor U6645 (N_6645,N_4798,N_4927);
nor U6646 (N_6646,N_5194,N_3923);
and U6647 (N_6647,N_5740,N_5808);
nand U6648 (N_6648,N_3261,N_3821);
nor U6649 (N_6649,N_4577,N_3082);
nand U6650 (N_6650,N_4531,N_3735);
and U6651 (N_6651,N_5526,N_5576);
nor U6652 (N_6652,N_5356,N_3955);
and U6653 (N_6653,N_4129,N_5450);
or U6654 (N_6654,N_4084,N_4280);
xor U6655 (N_6655,N_3669,N_3560);
or U6656 (N_6656,N_4513,N_5232);
nand U6657 (N_6657,N_5247,N_4761);
and U6658 (N_6658,N_5610,N_3308);
or U6659 (N_6659,N_5219,N_4240);
nor U6660 (N_6660,N_3650,N_4746);
or U6661 (N_6661,N_3545,N_4591);
or U6662 (N_6662,N_5032,N_4618);
xnor U6663 (N_6663,N_4906,N_3792);
and U6664 (N_6664,N_3810,N_5078);
nor U6665 (N_6665,N_5091,N_5515);
nor U6666 (N_6666,N_5612,N_4711);
nand U6667 (N_6667,N_4082,N_4221);
or U6668 (N_6668,N_4753,N_5414);
or U6669 (N_6669,N_4981,N_4055);
or U6670 (N_6670,N_3361,N_3455);
and U6671 (N_6671,N_3297,N_4839);
or U6672 (N_6672,N_3083,N_5273);
nor U6673 (N_6673,N_3159,N_5410);
nand U6674 (N_6674,N_3811,N_5476);
xnor U6675 (N_6675,N_4886,N_5606);
xnor U6676 (N_6676,N_3021,N_4866);
nor U6677 (N_6677,N_3526,N_5332);
and U6678 (N_6678,N_3964,N_4047);
xnor U6679 (N_6679,N_4077,N_5653);
or U6680 (N_6680,N_4809,N_3516);
and U6681 (N_6681,N_4168,N_4880);
or U6682 (N_6682,N_3248,N_4775);
nor U6683 (N_6683,N_3377,N_5923);
xnor U6684 (N_6684,N_4036,N_4413);
xor U6685 (N_6685,N_5714,N_5987);
and U6686 (N_6686,N_3951,N_3395);
and U6687 (N_6687,N_3446,N_4515);
nor U6688 (N_6688,N_4366,N_3689);
and U6689 (N_6689,N_4227,N_5722);
xor U6690 (N_6690,N_3022,N_5123);
and U6691 (N_6691,N_3090,N_4421);
nand U6692 (N_6692,N_5511,N_4086);
nand U6693 (N_6693,N_4991,N_4934);
nor U6694 (N_6694,N_3491,N_5106);
or U6695 (N_6695,N_3737,N_5250);
xor U6696 (N_6696,N_3713,N_4534);
and U6697 (N_6697,N_5828,N_5711);
or U6698 (N_6698,N_4326,N_3704);
nand U6699 (N_6699,N_3552,N_5516);
xor U6700 (N_6700,N_5006,N_4311);
nor U6701 (N_6701,N_5140,N_4715);
or U6702 (N_6702,N_3854,N_5369);
and U6703 (N_6703,N_5851,N_3837);
nand U6704 (N_6704,N_3099,N_5594);
or U6705 (N_6705,N_4175,N_4023);
xor U6706 (N_6706,N_3692,N_4724);
xor U6707 (N_6707,N_3005,N_5755);
nand U6708 (N_6708,N_4812,N_4238);
xnor U6709 (N_6709,N_4350,N_3056);
nor U6710 (N_6710,N_5443,N_3633);
nor U6711 (N_6711,N_5798,N_4741);
nor U6712 (N_6712,N_4299,N_4294);
or U6713 (N_6713,N_5344,N_3563);
nor U6714 (N_6714,N_3627,N_4363);
xnor U6715 (N_6715,N_5398,N_3482);
or U6716 (N_6716,N_5939,N_5880);
nand U6717 (N_6717,N_3299,N_4929);
or U6718 (N_6718,N_3971,N_4558);
xor U6719 (N_6719,N_3351,N_3155);
nand U6720 (N_6720,N_3311,N_4920);
nand U6721 (N_6721,N_3334,N_4423);
nand U6722 (N_6722,N_5687,N_3093);
nor U6723 (N_6723,N_5884,N_4915);
xor U6724 (N_6724,N_4669,N_5042);
or U6725 (N_6725,N_3166,N_3097);
nand U6726 (N_6726,N_5214,N_4514);
or U6727 (N_6727,N_5751,N_3133);
nand U6728 (N_6728,N_5507,N_5577);
xor U6729 (N_6729,N_3282,N_3275);
xor U6730 (N_6730,N_3728,N_5489);
xnor U6731 (N_6731,N_4867,N_4631);
and U6732 (N_6732,N_3121,N_5891);
or U6733 (N_6733,N_3639,N_5020);
and U6734 (N_6734,N_3254,N_4822);
and U6735 (N_6735,N_5620,N_4039);
and U6736 (N_6736,N_5467,N_4126);
nand U6737 (N_6737,N_5634,N_4169);
or U6738 (N_6738,N_3621,N_5734);
or U6739 (N_6739,N_5419,N_3893);
and U6740 (N_6740,N_5291,N_3846);
nor U6741 (N_6741,N_4320,N_5261);
or U6742 (N_6742,N_5564,N_5276);
and U6743 (N_6743,N_4150,N_3028);
xnor U6744 (N_6744,N_5629,N_3092);
nand U6745 (N_6745,N_5122,N_3635);
nand U6746 (N_6746,N_4572,N_3537);
nand U6747 (N_6747,N_3020,N_4743);
nand U6748 (N_6748,N_3255,N_4167);
nand U6749 (N_6749,N_5491,N_4331);
nor U6750 (N_6750,N_4697,N_5721);
and U6751 (N_6751,N_4690,N_4628);
xor U6752 (N_6752,N_4123,N_5254);
or U6753 (N_6753,N_5105,N_5695);
nand U6754 (N_6754,N_4833,N_3434);
or U6755 (N_6755,N_5270,N_5081);
xnor U6756 (N_6756,N_3676,N_4228);
nand U6757 (N_6757,N_3340,N_3542);
or U6758 (N_6758,N_5847,N_5098);
and U6759 (N_6759,N_5982,N_4604);
and U6760 (N_6760,N_4789,N_4517);
nor U6761 (N_6761,N_5128,N_5763);
nor U6762 (N_6762,N_3865,N_3421);
nor U6763 (N_6763,N_3711,N_4044);
xnor U6764 (N_6764,N_5882,N_3929);
nand U6765 (N_6765,N_4875,N_3503);
nand U6766 (N_6766,N_3345,N_4625);
nand U6767 (N_6767,N_4658,N_3920);
nor U6768 (N_6768,N_5008,N_4648);
xnor U6769 (N_6769,N_5621,N_3789);
nand U6770 (N_6770,N_5538,N_4287);
xnor U6771 (N_6771,N_5368,N_4989);
or U6772 (N_6772,N_3798,N_3209);
and U6773 (N_6773,N_4525,N_3087);
nor U6774 (N_6774,N_4524,N_4276);
and U6775 (N_6775,N_3667,N_5355);
and U6776 (N_6776,N_3431,N_5391);
nand U6777 (N_6777,N_3222,N_4135);
nand U6778 (N_6778,N_3086,N_3815);
nand U6779 (N_6779,N_4290,N_4776);
xnor U6780 (N_6780,N_4059,N_4824);
and U6781 (N_6781,N_5809,N_4703);
or U6782 (N_6782,N_3764,N_5554);
nand U6783 (N_6783,N_4456,N_3280);
or U6784 (N_6784,N_4980,N_4871);
nand U6785 (N_6785,N_5351,N_4339);
or U6786 (N_6786,N_3480,N_5664);
or U6787 (N_6787,N_3577,N_3182);
or U6788 (N_6788,N_5852,N_3928);
nand U6789 (N_6789,N_3029,N_4850);
xor U6790 (N_6790,N_3742,N_4616);
xor U6791 (N_6791,N_4463,N_3557);
nor U6792 (N_6792,N_4825,N_5802);
nand U6793 (N_6793,N_5846,N_5449);
and U6794 (N_6794,N_3976,N_4419);
xnor U6795 (N_6795,N_5623,N_3732);
and U6796 (N_6796,N_4806,N_5633);
and U6797 (N_6797,N_4696,N_4919);
and U6798 (N_6798,N_4881,N_3738);
nand U6799 (N_6799,N_5085,N_3495);
nand U6800 (N_6800,N_5874,N_5833);
nor U6801 (N_6801,N_4283,N_4854);
xor U6802 (N_6802,N_5613,N_3808);
nor U6803 (N_6803,N_5233,N_5221);
nand U6804 (N_6804,N_5742,N_5309);
or U6805 (N_6805,N_5004,N_5335);
or U6806 (N_6806,N_5530,N_5326);
nor U6807 (N_6807,N_4847,N_3598);
nor U6808 (N_6808,N_3994,N_4910);
xnor U6809 (N_6809,N_4319,N_5446);
nor U6810 (N_6810,N_4883,N_5104);
or U6811 (N_6811,N_4156,N_5337);
and U6812 (N_6812,N_4120,N_3511);
and U6813 (N_6813,N_3900,N_4832);
nor U6814 (N_6814,N_4750,N_5053);
xor U6815 (N_6815,N_4917,N_4401);
and U6816 (N_6816,N_3477,N_5810);
xnor U6817 (N_6817,N_5645,N_5215);
nor U6818 (N_6818,N_5321,N_5665);
xnor U6819 (N_6819,N_4335,N_3772);
xnor U6820 (N_6820,N_4499,N_4029);
or U6821 (N_6821,N_5720,N_4220);
nand U6822 (N_6822,N_3890,N_3720);
xnor U6823 (N_6823,N_3978,N_3153);
nand U6824 (N_6824,N_5765,N_5138);
nand U6825 (N_6825,N_5795,N_4699);
and U6826 (N_6826,N_3745,N_4639);
nor U6827 (N_6827,N_4737,N_3970);
and U6828 (N_6828,N_3868,N_3062);
xnor U6829 (N_6829,N_3809,N_3609);
or U6830 (N_6830,N_4638,N_5800);
or U6831 (N_6831,N_3270,N_3216);
or U6832 (N_6832,N_4000,N_5509);
xor U6833 (N_6833,N_3357,N_4936);
xor U6834 (N_6834,N_3736,N_5196);
xnor U6835 (N_6835,N_5881,N_4562);
nor U6836 (N_6836,N_3109,N_4194);
and U6837 (N_6837,N_4209,N_3321);
xnor U6838 (N_6838,N_3139,N_5787);
xor U6839 (N_6839,N_5372,N_3706);
nor U6840 (N_6840,N_4975,N_4950);
or U6841 (N_6841,N_3378,N_3473);
and U6842 (N_6842,N_4995,N_4285);
and U6843 (N_6843,N_4375,N_5444);
nand U6844 (N_6844,N_3363,N_4197);
nor U6845 (N_6845,N_4003,N_5036);
nor U6846 (N_6846,N_5198,N_5546);
and U6847 (N_6847,N_5794,N_3026);
nor U6848 (N_6848,N_5562,N_3642);
nand U6849 (N_6849,N_3693,N_5126);
nor U6850 (N_6850,N_5169,N_3217);
or U6851 (N_6851,N_5109,N_4773);
xor U6852 (N_6852,N_5204,N_4329);
nand U6853 (N_6853,N_4460,N_5595);
nor U6854 (N_6854,N_3679,N_3504);
nor U6855 (N_6855,N_3330,N_4125);
xor U6856 (N_6856,N_5339,N_3226);
and U6857 (N_6857,N_3879,N_3743);
and U6858 (N_6858,N_3492,N_3790);
xor U6859 (N_6859,N_3817,N_5870);
or U6860 (N_6860,N_3184,N_3405);
or U6861 (N_6861,N_3212,N_3871);
xor U6862 (N_6862,N_3674,N_4457);
nand U6863 (N_6863,N_5992,N_5937);
or U6864 (N_6864,N_4053,N_3499);
xor U6865 (N_6865,N_3629,N_3825);
nand U6866 (N_6866,N_5743,N_3543);
or U6867 (N_6867,N_4267,N_3161);
nand U6868 (N_6868,N_5096,N_4312);
or U6869 (N_6869,N_3283,N_5353);
nor U6870 (N_6870,N_5757,N_5424);
and U6871 (N_6871,N_5911,N_5593);
and U6872 (N_6872,N_4201,N_4552);
and U6873 (N_6873,N_3407,N_4606);
or U6874 (N_6874,N_5892,N_4533);
xnor U6875 (N_6875,N_5785,N_5544);
nor U6876 (N_6876,N_5589,N_3533);
nor U6877 (N_6877,N_3329,N_3638);
and U6878 (N_6878,N_3114,N_3235);
nor U6879 (N_6879,N_4671,N_4281);
or U6880 (N_6880,N_4551,N_3488);
and U6881 (N_6881,N_4217,N_4309);
nand U6882 (N_6882,N_3388,N_4720);
and U6883 (N_6883,N_4635,N_4482);
xnor U6884 (N_6884,N_5761,N_3420);
nand U6885 (N_6885,N_3665,N_4359);
and U6886 (N_6886,N_5054,N_4140);
xnor U6887 (N_6887,N_3384,N_3866);
nor U6888 (N_6888,N_4816,N_4870);
nor U6889 (N_6889,N_4547,N_4500);
or U6890 (N_6890,N_4765,N_5861);
or U6891 (N_6891,N_5317,N_5293);
or U6892 (N_6892,N_4200,N_5167);
xor U6893 (N_6893,N_5637,N_5125);
or U6894 (N_6894,N_5871,N_3284);
nand U6895 (N_6895,N_3371,N_5849);
xor U6896 (N_6896,N_5862,N_5831);
nor U6897 (N_6897,N_3838,N_3027);
and U6898 (N_6898,N_5243,N_5730);
nor U6899 (N_6899,N_5001,N_3722);
and U6900 (N_6900,N_3478,N_3273);
nand U6901 (N_6901,N_5565,N_5343);
and U6902 (N_6902,N_3712,N_3138);
or U6903 (N_6903,N_4653,N_3933);
or U6904 (N_6904,N_3894,N_4614);
or U6905 (N_6905,N_5910,N_3716);
or U6906 (N_6906,N_4672,N_3959);
nor U6907 (N_6907,N_4813,N_5915);
xor U6908 (N_6908,N_3323,N_4258);
or U6909 (N_6909,N_3829,N_5469);
and U6910 (N_6910,N_3874,N_4898);
and U6911 (N_6911,N_3152,N_3481);
nand U6912 (N_6912,N_5412,N_4873);
or U6913 (N_6913,N_5723,N_3033);
nand U6914 (N_6914,N_3356,N_4840);
nor U6915 (N_6915,N_3411,N_4213);
nand U6916 (N_6916,N_4115,N_5349);
and U6917 (N_6917,N_5890,N_3580);
nor U6918 (N_6918,N_5716,N_4066);
or U6919 (N_6919,N_5644,N_5868);
nor U6920 (N_6920,N_4251,N_3753);
nor U6921 (N_6921,N_3073,N_3999);
or U6922 (N_6922,N_5336,N_3171);
nand U6923 (N_6923,N_3454,N_5371);
nor U6924 (N_6924,N_4772,N_3433);
nand U6925 (N_6925,N_3515,N_4990);
nor U6926 (N_6926,N_5984,N_4038);
and U6927 (N_6927,N_3128,N_3043);
xor U6928 (N_6928,N_5701,N_4108);
and U6929 (N_6929,N_4754,N_5853);
nand U6930 (N_6930,N_3008,N_5827);
or U6931 (N_6931,N_3458,N_5916);
and U6932 (N_6932,N_4791,N_3368);
nor U6933 (N_6933,N_3256,N_4714);
and U6934 (N_6934,N_5070,N_5905);
nor U6935 (N_6935,N_3997,N_5154);
xnor U6936 (N_6936,N_3044,N_3058);
xor U6937 (N_6937,N_3353,N_3119);
nor U6938 (N_6938,N_5918,N_3319);
nor U6939 (N_6939,N_5869,N_4938);
nor U6940 (N_6940,N_3906,N_5425);
and U6941 (N_6941,N_4361,N_5962);
nand U6942 (N_6942,N_3442,N_5009);
nand U6943 (N_6943,N_3938,N_3646);
nand U6944 (N_6944,N_5655,N_3293);
nand U6945 (N_6945,N_5632,N_5110);
and U6946 (N_6946,N_5306,N_5944);
xor U6947 (N_6947,N_3600,N_5732);
nor U6948 (N_6948,N_5748,N_5438);
and U6949 (N_6949,N_3953,N_4611);
or U6950 (N_6950,N_4353,N_5708);
nor U6951 (N_6951,N_4009,N_4334);
nand U6952 (N_6952,N_5626,N_3410);
or U6953 (N_6953,N_4298,N_4649);
or U6954 (N_6954,N_4657,N_3654);
nor U6955 (N_6955,N_3721,N_4376);
xor U6956 (N_6956,N_5239,N_4435);
and U6957 (N_6957,N_5581,N_4212);
or U6958 (N_6958,N_4751,N_5165);
xor U6959 (N_6959,N_4032,N_5047);
nand U6960 (N_6960,N_3055,N_5932);
xnor U6961 (N_6961,N_5016,N_5470);
nand U6962 (N_6962,N_3306,N_3945);
nand U6963 (N_6963,N_5082,N_4446);
nor U6964 (N_6964,N_5791,N_5933);
nor U6965 (N_6965,N_3641,N_5191);
nand U6966 (N_6966,N_4781,N_4595);
xnor U6967 (N_6967,N_3949,N_3199);
and U6968 (N_6968,N_3726,N_3591);
nand U6969 (N_6969,N_5964,N_3052);
xor U6970 (N_6970,N_3911,N_4182);
xnor U6971 (N_6971,N_5698,N_5249);
or U6972 (N_6972,N_4222,N_3012);
and U6973 (N_6973,N_4939,N_3198);
nand U6974 (N_6974,N_4528,N_5213);
xor U6975 (N_6975,N_4296,N_4430);
and U6976 (N_6976,N_3444,N_5127);
or U6977 (N_6977,N_4325,N_4819);
or U6978 (N_6978,N_4651,N_5834);
xor U6979 (N_6979,N_3367,N_4328);
and U6980 (N_6980,N_3169,N_4400);
xnor U6981 (N_6981,N_5817,N_4374);
nand U6982 (N_6982,N_5260,N_5974);
nand U6983 (N_6983,N_5440,N_5900);
nor U6984 (N_6984,N_4368,N_4165);
xnor U6985 (N_6985,N_3687,N_3990);
nand U6986 (N_6986,N_5609,N_4710);
and U6987 (N_6987,N_4148,N_4843);
or U6988 (N_6988,N_5952,N_4678);
xnor U6989 (N_6989,N_4188,N_3009);
nand U6990 (N_6990,N_4621,N_3827);
or U6991 (N_6991,N_5366,N_4028);
nand U6992 (N_6992,N_5083,N_5285);
or U6993 (N_6993,N_5028,N_5611);
or U6994 (N_6994,N_4622,N_3870);
nor U6995 (N_6995,N_4838,N_5141);
nand U6996 (N_6996,N_5859,N_5976);
or U6997 (N_6997,N_5574,N_3260);
xnor U6998 (N_6998,N_4043,N_3381);
nand U6999 (N_6999,N_4997,N_4768);
nand U7000 (N_7000,N_5749,N_3342);
and U7001 (N_7001,N_4263,N_5375);
nand U7002 (N_7002,N_3145,N_5034);
and U7003 (N_7003,N_4153,N_5487);
xnor U7004 (N_7004,N_3510,N_5940);
and U7005 (N_7005,N_5579,N_5925);
xor U7006 (N_7006,N_5178,N_4024);
and U7007 (N_7007,N_5026,N_5549);
nand U7008 (N_7008,N_5283,N_5767);
or U7009 (N_7009,N_3839,N_5280);
or U7010 (N_7010,N_5622,N_5552);
xor U7011 (N_7011,N_4282,N_4942);
and U7012 (N_7012,N_3574,N_4270);
nand U7013 (N_7013,N_4346,N_3502);
xnor U7014 (N_7014,N_3775,N_5201);
nor U7015 (N_7015,N_5998,N_4317);
xnor U7016 (N_7016,N_5227,N_3556);
xor U7017 (N_7017,N_3137,N_4641);
nor U7018 (N_7018,N_5093,N_4924);
nand U7019 (N_7019,N_4412,N_5929);
or U7020 (N_7020,N_4801,N_5679);
and U7021 (N_7021,N_4858,N_4844);
xor U7022 (N_7022,N_5241,N_3347);
or U7023 (N_7023,N_4483,N_3279);
and U7024 (N_7024,N_3286,N_4052);
or U7025 (N_7025,N_5947,N_5886);
or U7026 (N_7026,N_5277,N_3160);
and U7027 (N_7027,N_5428,N_3897);
nand U7028 (N_7028,N_4091,N_5035);
or U7029 (N_7029,N_4216,N_4518);
and U7030 (N_7030,N_5887,N_5010);
nand U7031 (N_7031,N_5628,N_3429);
and U7032 (N_7032,N_4861,N_4613);
xnor U7033 (N_7033,N_3914,N_4977);
nand U7034 (N_7034,N_3573,N_5841);
nand U7035 (N_7035,N_5811,N_4386);
nor U7036 (N_7036,N_4803,N_3942);
nand U7037 (N_7037,N_3688,N_3778);
or U7038 (N_7038,N_5744,N_3440);
or U7039 (N_7039,N_4396,N_3797);
or U7040 (N_7040,N_3876,N_3071);
or U7041 (N_7041,N_5423,N_3562);
nor U7042 (N_7042,N_5207,N_4445);
nor U7043 (N_7043,N_5224,N_3088);
xnor U7044 (N_7044,N_3905,N_3223);
xor U7045 (N_7045,N_3349,N_5031);
xnor U7046 (N_7046,N_3813,N_5238);
or U7047 (N_7047,N_5786,N_3852);
nor U7048 (N_7048,N_3766,N_4523);
or U7049 (N_7049,N_4810,N_5731);
nand U7050 (N_7050,N_5824,N_4432);
nand U7051 (N_7051,N_4073,N_5051);
or U7052 (N_7052,N_5726,N_4447);
and U7053 (N_7053,N_4565,N_3383);
xnor U7054 (N_7054,N_5830,N_3535);
xnor U7055 (N_7055,N_4060,N_5599);
nand U7056 (N_7056,N_3229,N_3584);
nor U7057 (N_7057,N_5951,N_3475);
or U7058 (N_7058,N_4056,N_3973);
nor U7059 (N_7059,N_5041,N_5771);
or U7060 (N_7060,N_5584,N_4582);
or U7061 (N_7061,N_4415,N_4691);
xnor U7062 (N_7062,N_3366,N_3672);
nor U7063 (N_7063,N_4855,N_3077);
xnor U7064 (N_7064,N_4876,N_4002);
nor U7065 (N_7065,N_4490,N_5397);
and U7066 (N_7066,N_5415,N_3105);
nor U7067 (N_7067,N_3812,N_5166);
nand U7068 (N_7068,N_3593,N_3327);
xor U7069 (N_7069,N_5094,N_5304);
xor U7070 (N_7070,N_3501,N_3150);
nand U7071 (N_7071,N_5056,N_4788);
xor U7072 (N_7072,N_3135,N_4259);
and U7073 (N_7073,N_4993,N_4315);
nor U7074 (N_7074,N_4972,N_4358);
and U7075 (N_7075,N_5251,N_4519);
nand U7076 (N_7076,N_5465,N_5168);
nor U7077 (N_7077,N_4471,N_5360);
and U7078 (N_7078,N_4393,N_3493);
nor U7079 (N_7079,N_5043,N_3787);
or U7080 (N_7080,N_3553,N_5156);
xnor U7081 (N_7081,N_4147,N_3585);
or U7082 (N_7082,N_4098,N_3509);
nor U7083 (N_7083,N_5055,N_4189);
and U7084 (N_7084,N_3201,N_5536);
or U7085 (N_7085,N_4510,N_4718);
or U7086 (N_7086,N_3467,N_4122);
xnor U7087 (N_7087,N_4394,N_3774);
nor U7088 (N_7088,N_4701,N_3886);
or U7089 (N_7089,N_5401,N_3907);
and U7090 (N_7090,N_3130,N_3656);
nor U7091 (N_7091,N_4223,N_5503);
nor U7092 (N_7092,N_5832,N_5733);
or U7093 (N_7093,N_4706,N_4161);
and U7094 (N_7094,N_4563,N_4543);
nand U7095 (N_7095,N_5097,N_3752);
and U7096 (N_7096,N_3122,N_5050);
nor U7097 (N_7097,N_3658,N_3606);
or U7098 (N_7098,N_4941,N_3963);
nand U7099 (N_7099,N_4425,N_4893);
nor U7100 (N_7100,N_5903,N_5478);
nand U7101 (N_7101,N_5022,N_3723);
nand U7102 (N_7102,N_4503,N_3437);
or U7103 (N_7103,N_3673,N_5700);
xnor U7104 (N_7104,N_4398,N_4089);
or U7105 (N_7105,N_3538,N_5359);
nand U7106 (N_7106,N_3967,N_5745);
xnor U7107 (N_7107,N_5358,N_4579);
or U7108 (N_7108,N_5416,N_3719);
nand U7109 (N_7109,N_4660,N_4127);
or U7110 (N_7110,N_4857,N_3131);
or U7111 (N_7111,N_4377,N_3788);
nand U7112 (N_7112,N_5774,N_5092);
or U7113 (N_7113,N_5736,N_5319);
xnor U7114 (N_7114,N_3525,N_3754);
nand U7115 (N_7115,N_5535,N_3885);
or U7116 (N_7116,N_4979,N_5400);
nor U7117 (N_7117,N_4592,N_4434);
xor U7118 (N_7118,N_3309,N_5980);
xnor U7119 (N_7119,N_5978,N_3760);
or U7120 (N_7120,N_4911,N_3660);
nand U7121 (N_7121,N_5324,N_4476);
xor U7122 (N_7122,N_4260,N_4738);
nor U7123 (N_7123,N_5473,N_5860);
xor U7124 (N_7124,N_3344,N_4402);
or U7125 (N_7125,N_5889,N_5624);
nand U7126 (N_7126,N_4341,N_3300);
or U7127 (N_7127,N_3541,N_5652);
xnor U7128 (N_7128,N_5677,N_5269);
nand U7129 (N_7129,N_5559,N_3277);
nor U7130 (N_7130,N_5659,N_4502);
nand U7131 (N_7131,N_4633,N_3861);
nand U7132 (N_7132,N_4252,N_5955);
nand U7133 (N_7133,N_3337,N_3969);
nand U7134 (N_7134,N_5635,N_5435);
nand U7135 (N_7135,N_4068,N_5705);
xnor U7136 (N_7136,N_4585,N_3054);
or U7137 (N_7137,N_3659,N_5308);
nand U7138 (N_7138,N_5505,N_3380);
nor U7139 (N_7139,N_3630,N_4713);
nor U7140 (N_7140,N_3989,N_3761);
or U7141 (N_7141,N_4874,N_4455);
and U7142 (N_7142,N_3981,N_4656);
or U7143 (N_7143,N_5388,N_3756);
nand U7144 (N_7144,N_3140,N_4352);
and U7145 (N_7145,N_5199,N_4040);
nand U7146 (N_7146,N_3251,N_4382);
xnor U7147 (N_7147,N_5780,N_5381);
and U7148 (N_7148,N_3379,N_5448);
nor U7149 (N_7149,N_5569,N_5975);
or U7150 (N_7150,N_3424,N_5689);
or U7151 (N_7151,N_4134,N_3524);
and U7152 (N_7152,N_5855,N_3529);
and U7153 (N_7153,N_4433,N_3818);
xor U7154 (N_7154,N_3864,N_5259);
nand U7155 (N_7155,N_5523,N_4985);
xnor U7156 (N_7156,N_3218,N_4687);
nor U7157 (N_7157,N_4118,N_4940);
and U7158 (N_7158,N_3250,N_4333);
nor U7159 (N_7159,N_5363,N_4955);
nor U7160 (N_7160,N_4271,N_3274);
and U7161 (N_7161,N_4347,N_3195);
and U7162 (N_7162,N_4532,N_3129);
nor U7163 (N_7163,N_4600,N_4162);
nand U7164 (N_7164,N_5688,N_5208);
and U7165 (N_7165,N_5217,N_4186);
or U7166 (N_7166,N_3806,N_5747);
xor U7167 (N_7167,N_3946,N_3312);
nor U7168 (N_7168,N_3120,N_4452);
xnor U7169 (N_7169,N_3485,N_4647);
nand U7170 (N_7170,N_5145,N_3622);
nor U7171 (N_7171,N_4829,N_5822);
nor U7172 (N_7172,N_5325,N_5801);
xnor U7173 (N_7173,N_3578,N_4142);
or U7174 (N_7174,N_3530,N_5572);
nand U7175 (N_7175,N_3289,N_4769);
nand U7176 (N_7176,N_4356,N_5857);
or U7177 (N_7177,N_4557,N_4539);
nand U7178 (N_7178,N_4770,N_4787);
nand U7179 (N_7179,N_5850,N_3972);
or U7180 (N_7180,N_5320,N_4427);
nor U7181 (N_7181,N_4278,N_4160);
and U7182 (N_7182,N_4466,N_5777);
xnor U7183 (N_7183,N_4581,N_3134);
nand U7184 (N_7184,N_5420,N_3430);
nor U7185 (N_7185,N_5919,N_3189);
and U7186 (N_7186,N_4605,N_5310);
nand U7187 (N_7187,N_3662,N_5345);
nand U7188 (N_7188,N_4973,N_4288);
or U7189 (N_7189,N_4537,N_4619);
and U7190 (N_7190,N_3605,N_3581);
nor U7191 (N_7191,N_3402,N_3675);
nor U7192 (N_7192,N_4764,N_5753);
xor U7193 (N_7193,N_5455,N_3315);
or U7194 (N_7194,N_3831,N_4608);
nand U7195 (N_7195,N_3828,N_4992);
nor U7196 (N_7196,N_3414,N_5313);
or U7197 (N_7197,N_3464,N_5630);
nand U7198 (N_7198,N_4110,N_3583);
or U7199 (N_7199,N_3123,N_3360);
and U7200 (N_7200,N_5588,N_4448);
nand U7201 (N_7201,N_4707,N_5879);
nand U7202 (N_7202,N_5985,N_3862);
or U7203 (N_7203,N_5959,N_4726);
xor U7204 (N_7204,N_4340,N_5057);
xor U7205 (N_7205,N_3988,N_3844);
xor U7206 (N_7206,N_3604,N_5907);
and U7207 (N_7207,N_3389,N_5960);
nor U7208 (N_7208,N_3912,N_3506);
or U7209 (N_7209,N_4480,N_4722);
nor U7210 (N_7210,N_4088,N_3993);
nor U7211 (N_7211,N_4099,N_5237);
and U7212 (N_7212,N_5382,N_4885);
and U7213 (N_7213,N_5275,N_4841);
or U7214 (N_7214,N_4856,N_3698);
nor U7215 (N_7215,N_3035,N_4610);
xor U7216 (N_7216,N_4580,N_4918);
nand U7217 (N_7217,N_3952,N_4185);
xor U7218 (N_7218,N_4464,N_4069);
xnor U7219 (N_7219,N_4454,N_5229);
and U7220 (N_7220,N_5408,N_5707);
nor U7221 (N_7221,N_3374,N_3648);
or U7222 (N_7222,N_5303,N_5683);
nand U7223 (N_7223,N_5186,N_4210);
nor U7224 (N_7224,N_4081,N_3154);
nor U7225 (N_7225,N_4342,N_3568);
and U7226 (N_7226,N_4244,N_5288);
and U7227 (N_7227,N_5563,N_5596);
and U7228 (N_7228,N_5100,N_5494);
and U7229 (N_7229,N_3178,N_5840);
nand U7230 (N_7230,N_5602,N_5257);
nand U7231 (N_7231,N_3324,N_4644);
nand U7232 (N_7232,N_3463,N_5255);
nand U7233 (N_7233,N_5268,N_4780);
nor U7234 (N_7234,N_5228,N_4807);
nor U7235 (N_7235,N_3966,N_5445);
or U7236 (N_7236,N_5297,N_5759);
or U7237 (N_7237,N_4762,N_4172);
nand U7238 (N_7238,N_3011,N_5301);
nor U7239 (N_7239,N_4131,N_5573);
nor U7240 (N_7240,N_4261,N_4851);
and U7241 (N_7241,N_4589,N_3314);
nand U7242 (N_7242,N_5863,N_3124);
xnor U7243 (N_7243,N_4397,N_3695);
nand U7244 (N_7244,N_4922,N_5512);
nand U7245 (N_7245,N_4961,N_5481);
xnor U7246 (N_7246,N_3569,N_5718);
nand U7247 (N_7247,N_3132,N_5463);
and U7248 (N_7248,N_3146,N_4384);
or U7249 (N_7249,N_3142,N_5518);
and U7250 (N_7250,N_3287,N_5072);
nand U7251 (N_7251,N_3447,N_4507);
nor U7252 (N_7252,N_5547,N_5704);
xnor U7253 (N_7253,N_4473,N_4721);
xor U7254 (N_7254,N_3851,N_4307);
xor U7255 (N_7255,N_5386,N_3252);
and U7256 (N_7256,N_3081,N_3895);
nor U7257 (N_7257,N_3066,N_4907);
or U7258 (N_7258,N_4491,N_5680);
and U7259 (N_7259,N_5246,N_4727);
xnor U7260 (N_7260,N_5783,N_3683);
nand U7261 (N_7261,N_5971,N_3741);
and U7262 (N_7262,N_5177,N_3610);
nor U7263 (N_7263,N_3796,N_5222);
nand U7264 (N_7264,N_3983,N_4637);
and U7265 (N_7265,N_5914,N_4556);
and U7266 (N_7266,N_5179,N_5973);
nor U7267 (N_7267,N_3188,N_3399);
or U7268 (N_7268,N_5426,N_5906);
and U7269 (N_7269,N_5990,N_4229);
nor U7270 (N_7270,N_4598,N_4739);
nor U7271 (N_7271,N_3304,N_3663);
xnor U7272 (N_7272,N_3799,N_5519);
xor U7273 (N_7273,N_4075,N_3164);
and U7274 (N_7274,N_5897,N_3561);
and U7275 (N_7275,N_4527,N_3645);
or U7276 (N_7276,N_5087,N_5696);
and U7277 (N_7277,N_5253,N_3965);
nor U7278 (N_7278,N_4174,N_4230);
and U7279 (N_7279,N_3670,N_5815);
xnor U7280 (N_7280,N_5854,N_5865);
or U7281 (N_7281,N_5970,N_3465);
nand U7282 (N_7282,N_3684,N_4888);
and U7283 (N_7283,N_5543,N_3918);
or U7284 (N_7284,N_3354,N_4012);
nor U7285 (N_7285,N_5248,N_3350);
nand U7286 (N_7286,N_3241,N_5099);
or U7287 (N_7287,N_3298,N_5981);
and U7288 (N_7288,N_4912,N_3857);
and U7289 (N_7289,N_4428,N_3926);
and U7290 (N_7290,N_4351,N_4308);
nor U7291 (N_7291,N_3805,N_4571);
nor U7292 (N_7292,N_4814,N_4301);
nand U7293 (N_7293,N_5302,N_4909);
nand U7294 (N_7294,N_5296,N_3540);
nand U7295 (N_7295,N_5888,N_4693);
or U7296 (N_7296,N_4484,N_4823);
or U7297 (N_7297,N_4615,N_3532);
nand U7298 (N_7298,N_5666,N_4599);
and U7299 (N_7299,N_4021,N_5510);
nor U7300 (N_7300,N_4921,N_4470);
and U7301 (N_7301,N_3592,N_4094);
xor U7302 (N_7302,N_4522,N_5120);
nand U7303 (N_7303,N_4952,N_3705);
nand U7304 (N_7304,N_4453,N_5776);
and U7305 (N_7305,N_5064,N_3765);
and U7306 (N_7306,N_3940,N_5027);
nor U7307 (N_7307,N_3163,N_3288);
and U7308 (N_7308,N_3830,N_3462);
and U7309 (N_7309,N_5501,N_4682);
xnor U7310 (N_7310,N_3935,N_4139);
or U7311 (N_7311,N_4141,N_3193);
nor U7312 (N_7312,N_4521,N_3696);
nand U7313 (N_7313,N_4332,N_3823);
nor U7314 (N_7314,N_3858,N_5894);
nor U7315 (N_7315,N_4925,N_5674);
and U7316 (N_7316,N_4295,N_5454);
or U7317 (N_7317,N_5597,N_3744);
nor U7318 (N_7318,N_4392,N_3779);
or U7319 (N_7319,N_3505,N_3307);
xnor U7320 (N_7320,N_4248,N_4698);
nand U7321 (N_7321,N_5570,N_3939);
nand U7322 (N_7322,N_3590,N_5163);
nor U7323 (N_7323,N_4488,N_3471);
xnor U7324 (N_7324,N_5899,N_5758);
and U7325 (N_7325,N_5282,N_5486);
nor U7326 (N_7326,N_3413,N_3365);
or U7327 (N_7327,N_3339,N_5746);
nor U7328 (N_7328,N_5411,N_5586);
xnor U7329 (N_7329,N_3513,N_3762);
nor U7330 (N_7330,N_4663,N_3522);
or U7331 (N_7331,N_5686,N_5654);
nand U7332 (N_7332,N_3757,N_5340);
xor U7333 (N_7333,N_5295,N_3927);
and U7334 (N_7334,N_5095,N_5350);
nor U7335 (N_7335,N_5661,N_5591);
and U7336 (N_7336,N_5965,N_5803);
nand U7337 (N_7337,N_5513,N_5024);
xnor U7338 (N_7338,N_3244,N_4597);
nor U7339 (N_7339,N_3080,N_5286);
xor U7340 (N_7340,N_3793,N_4255);
xor U7341 (N_7341,N_5329,N_3069);
and U7342 (N_7342,N_4015,N_5284);
or U7343 (N_7343,N_5717,N_3177);
nand U7344 (N_7344,N_4370,N_4431);
nor U7345 (N_7345,N_3276,N_5956);
nand U7346 (N_7346,N_3294,N_4757);
and U7347 (N_7347,N_5575,N_5150);
nand U7348 (N_7348,N_3014,N_4926);
xnor U7349 (N_7349,N_5011,N_4586);
nor U7350 (N_7350,N_3243,N_3873);
xor U7351 (N_7351,N_4159,N_3445);
or U7352 (N_7352,N_3637,N_4219);
nand U7353 (N_7353,N_4566,N_5452);
and U7354 (N_7354,N_3564,N_4546);
and U7355 (N_7355,N_3174,N_4417);
and U7356 (N_7356,N_3514,N_3567);
nand U7357 (N_7357,N_5089,N_5190);
nand U7358 (N_7358,N_3450,N_3476);
nand U7359 (N_7359,N_5457,N_3531);
and U7360 (N_7360,N_4853,N_4111);
and U7361 (N_7361,N_5986,N_4318);
and U7362 (N_7362,N_4568,N_4681);
or U7363 (N_7363,N_5162,N_4732);
nand U7364 (N_7364,N_3937,N_4676);
nor U7365 (N_7365,N_3680,N_4365);
nor U7366 (N_7366,N_4574,N_5735);
nand U7367 (N_7367,N_3691,N_4199);
nor U7368 (N_7368,N_3554,N_5934);
nor U7369 (N_7369,N_5129,N_4214);
and U7370 (N_7370,N_4896,N_4061);
and U7371 (N_7371,N_3608,N_3346);
or U7372 (N_7372,N_3718,N_4192);
and U7373 (N_7373,N_4904,N_5379);
nand U7374 (N_7374,N_4026,N_3617);
nor U7375 (N_7375,N_3415,N_3143);
or U7376 (N_7376,N_3826,N_3925);
or U7377 (N_7377,N_3422,N_4777);
and U7378 (N_7378,N_4204,N_4426);
nor U7379 (N_7379,N_5737,N_5171);
or U7380 (N_7380,N_3898,N_4560);
nor U7381 (N_7381,N_4327,N_5908);
and U7382 (N_7382,N_3459,N_5966);
nor U7383 (N_7383,N_5348,N_5935);
or U7384 (N_7384,N_4302,N_5130);
and U7385 (N_7385,N_3814,N_5506);
and U7386 (N_7386,N_3724,N_5005);
and U7387 (N_7387,N_5694,N_5160);
nand U7388 (N_7388,N_4974,N_3682);
xor U7389 (N_7389,N_5499,N_4305);
nor U7390 (N_7390,N_5895,N_5225);
and U7391 (N_7391,N_3619,N_5685);
or U7392 (N_7392,N_3883,N_5837);
xor U7393 (N_7393,N_5482,N_3889);
nor U7394 (N_7394,N_3328,N_4797);
nand U7395 (N_7395,N_3652,N_5657);
or U7396 (N_7396,N_3717,N_5673);
and U7397 (N_7397,N_3671,N_4763);
nor U7398 (N_7398,N_5715,N_4584);
xor U7399 (N_7399,N_5896,N_4708);
nor U7400 (N_7400,N_3238,N_5996);
and U7401 (N_7401,N_5764,N_4136);
xnor U7402 (N_7402,N_5210,N_4852);
nand U7403 (N_7403,N_4232,N_3739);
and U7404 (N_7404,N_4001,N_3613);
nand U7405 (N_7405,N_3333,N_4495);
and U7406 (N_7406,N_3053,N_3336);
and U7407 (N_7407,N_5557,N_3807);
and U7408 (N_7408,N_3302,N_3469);
and U7409 (N_7409,N_5052,N_4734);
nor U7410 (N_7410,N_5936,N_3213);
xnor U7411 (N_7411,N_4050,N_4778);
nand U7412 (N_7412,N_4062,N_5790);
nand U7413 (N_7413,N_3269,N_5003);
nor U7414 (N_7414,N_3176,N_5202);
nand U7415 (N_7415,N_3975,N_5485);
or U7416 (N_7416,N_3521,N_3517);
nand U7417 (N_7417,N_5429,N_4128);
nor U7418 (N_7418,N_3257,N_5582);
nand U7419 (N_7419,N_4588,N_3896);
or U7420 (N_7420,N_3397,N_4424);
nand U7421 (N_7421,N_4065,N_3230);
or U7422 (N_7422,N_5058,N_4646);
xor U7423 (N_7423,N_5025,N_4771);
or U7424 (N_7424,N_5999,N_5545);
xnor U7425 (N_7425,N_4736,N_4106);
and U7426 (N_7426,N_5772,N_5471);
and U7427 (N_7427,N_4019,N_4624);
nand U7428 (N_7428,N_4559,N_3400);
xor U7429 (N_7429,N_3850,N_4967);
or U7430 (N_7430,N_4666,N_4016);
nor U7431 (N_7431,N_4385,N_5316);
nor U7432 (N_7432,N_4845,N_4109);
or U7433 (N_7433,N_5147,N_5212);
or U7434 (N_7434,N_4716,N_5669);
or U7435 (N_7435,N_4321,N_5993);
and U7436 (N_7436,N_4154,N_3962);
and U7437 (N_7437,N_5480,N_5033);
nand U7438 (N_7438,N_3259,N_5684);
xnor U7439 (N_7439,N_4493,N_4095);
or U7440 (N_7440,N_5307,N_4846);
and U7441 (N_7441,N_3842,N_4686);
and U7442 (N_7442,N_4241,N_5103);
and U7443 (N_7443,N_4978,N_3050);
xnor U7444 (N_7444,N_4779,N_5084);
xor U7445 (N_7445,N_3348,N_5823);
nand U7446 (N_7446,N_5021,N_4254);
nand U7447 (N_7447,N_4944,N_3419);
nor U7448 (N_7448,N_3127,N_3042);
nand U7449 (N_7449,N_5917,N_5342);
xnor U7450 (N_7450,N_3616,N_3888);
or U7451 (N_7451,N_5352,N_4472);
and U7452 (N_7452,N_4020,N_3000);
and U7453 (N_7453,N_5367,N_3264);
xor U7454 (N_7454,N_3158,N_5867);
nand U7455 (N_7455,N_3891,N_3362);
or U7456 (N_7456,N_3401,N_4575);
nand U7457 (N_7457,N_4195,N_5719);
nor U7458 (N_7458,N_4982,N_4758);
nand U7459 (N_7459,N_4008,N_3771);
nand U7460 (N_7460,N_3730,N_3141);
or U7461 (N_7461,N_3859,N_4603);
nand U7462 (N_7462,N_5108,N_4661);
nand U7463 (N_7463,N_4848,N_5220);
or U7464 (N_7464,N_4485,N_5173);
nand U7465 (N_7465,N_4496,N_4817);
nor U7466 (N_7466,N_4045,N_3332);
xnor U7467 (N_7467,N_4486,N_3448);
nor U7468 (N_7468,N_4899,N_3125);
or U7469 (N_7469,N_5418,N_4253);
or U7470 (N_7470,N_3219,N_3835);
xnor U7471 (N_7471,N_3634,N_4249);
xor U7472 (N_7472,N_5972,N_5453);
xnor U7473 (N_7473,N_5389,N_4155);
xnor U7474 (N_7474,N_5334,N_5231);
and U7475 (N_7475,N_4272,N_5149);
and U7476 (N_7476,N_5183,N_5311);
nand U7477 (N_7477,N_4101,N_3004);
nand U7478 (N_7478,N_4842,N_4937);
or U7479 (N_7479,N_4441,N_5566);
nand U7480 (N_7480,N_4378,N_3559);
and U7481 (N_7481,N_4680,N_5995);
xnor U7482 (N_7482,N_4735,N_3285);
nand U7483 (N_7483,N_4487,N_4709);
xnor U7484 (N_7484,N_4250,N_4233);
and U7485 (N_7485,N_3072,N_5067);
and U7486 (N_7486,N_4783,N_4133);
nand U7487 (N_7487,N_3048,N_3523);
nor U7488 (N_7488,N_5015,N_5155);
nand U7489 (N_7489,N_4005,N_3576);
and U7490 (N_7490,N_4300,N_4149);
xnor U7491 (N_7491,N_3623,N_5439);
nand U7492 (N_7492,N_5660,N_4828);
nor U7493 (N_7493,N_4717,N_3597);
xor U7494 (N_7494,N_4831,N_3258);
nor U7495 (N_7495,N_5354,N_5430);
nand U7496 (N_7496,N_4048,N_3115);
or U7497 (N_7497,N_3987,N_3607);
or U7498 (N_7498,N_3729,N_5132);
xnor U7499 (N_7499,N_4987,N_3802);
nand U7500 (N_7500,N_5286,N_4988);
xor U7501 (N_7501,N_3856,N_5249);
and U7502 (N_7502,N_5135,N_5587);
nand U7503 (N_7503,N_5746,N_5869);
xnor U7504 (N_7504,N_3432,N_4656);
and U7505 (N_7505,N_3375,N_4458);
nor U7506 (N_7506,N_3944,N_3614);
or U7507 (N_7507,N_5458,N_4066);
or U7508 (N_7508,N_3159,N_4622);
xnor U7509 (N_7509,N_4886,N_5281);
nor U7510 (N_7510,N_3091,N_5319);
xnor U7511 (N_7511,N_5618,N_5183);
and U7512 (N_7512,N_4607,N_4814);
nand U7513 (N_7513,N_3898,N_3861);
nand U7514 (N_7514,N_3592,N_5369);
nor U7515 (N_7515,N_4400,N_4918);
nand U7516 (N_7516,N_5314,N_3933);
xor U7517 (N_7517,N_3002,N_5564);
xnor U7518 (N_7518,N_4096,N_4719);
nand U7519 (N_7519,N_5152,N_4364);
and U7520 (N_7520,N_3391,N_4437);
nor U7521 (N_7521,N_3052,N_3898);
nor U7522 (N_7522,N_4403,N_3859);
nand U7523 (N_7523,N_4280,N_4510);
nor U7524 (N_7524,N_3388,N_4876);
or U7525 (N_7525,N_5878,N_3781);
nand U7526 (N_7526,N_3736,N_5819);
and U7527 (N_7527,N_3933,N_5243);
nand U7528 (N_7528,N_4582,N_5220);
nand U7529 (N_7529,N_5323,N_4269);
and U7530 (N_7530,N_3072,N_5391);
or U7531 (N_7531,N_4016,N_3922);
or U7532 (N_7532,N_5035,N_4515);
nor U7533 (N_7533,N_4572,N_5298);
nand U7534 (N_7534,N_3492,N_5102);
nor U7535 (N_7535,N_4165,N_5833);
nor U7536 (N_7536,N_5149,N_4401);
and U7537 (N_7537,N_4437,N_4292);
xnor U7538 (N_7538,N_4272,N_3227);
nor U7539 (N_7539,N_5807,N_4102);
nand U7540 (N_7540,N_5250,N_3885);
xnor U7541 (N_7541,N_5699,N_4509);
nand U7542 (N_7542,N_4900,N_4738);
or U7543 (N_7543,N_4536,N_5663);
xor U7544 (N_7544,N_4097,N_4923);
or U7545 (N_7545,N_5550,N_5036);
nor U7546 (N_7546,N_5444,N_4387);
xor U7547 (N_7547,N_3021,N_3322);
nand U7548 (N_7548,N_4305,N_4621);
or U7549 (N_7549,N_4661,N_4523);
nand U7550 (N_7550,N_3705,N_4304);
xnor U7551 (N_7551,N_4854,N_5238);
or U7552 (N_7552,N_3670,N_4856);
nand U7553 (N_7553,N_3359,N_5169);
nor U7554 (N_7554,N_4202,N_4304);
or U7555 (N_7555,N_3394,N_3398);
nand U7556 (N_7556,N_3744,N_3962);
nor U7557 (N_7557,N_3739,N_5188);
or U7558 (N_7558,N_5270,N_5137);
xnor U7559 (N_7559,N_3492,N_4258);
xor U7560 (N_7560,N_4825,N_3890);
xnor U7561 (N_7561,N_5560,N_5352);
nand U7562 (N_7562,N_3016,N_4893);
nor U7563 (N_7563,N_4616,N_5392);
nor U7564 (N_7564,N_5475,N_4945);
nand U7565 (N_7565,N_5761,N_3761);
and U7566 (N_7566,N_5148,N_3340);
nand U7567 (N_7567,N_3445,N_3530);
nor U7568 (N_7568,N_4395,N_4328);
nand U7569 (N_7569,N_3752,N_4945);
nand U7570 (N_7570,N_4919,N_3696);
nand U7571 (N_7571,N_5118,N_3576);
and U7572 (N_7572,N_3432,N_5939);
nand U7573 (N_7573,N_4027,N_4573);
or U7574 (N_7574,N_3946,N_3231);
or U7575 (N_7575,N_4116,N_4088);
and U7576 (N_7576,N_4547,N_4183);
and U7577 (N_7577,N_4150,N_4379);
and U7578 (N_7578,N_5284,N_5480);
nor U7579 (N_7579,N_4732,N_5373);
and U7580 (N_7580,N_4190,N_5357);
nor U7581 (N_7581,N_5283,N_5851);
xnor U7582 (N_7582,N_5422,N_3758);
nand U7583 (N_7583,N_3334,N_5594);
xnor U7584 (N_7584,N_5478,N_3704);
nand U7585 (N_7585,N_5927,N_3717);
and U7586 (N_7586,N_3571,N_5997);
or U7587 (N_7587,N_3529,N_4699);
nor U7588 (N_7588,N_4720,N_4291);
nor U7589 (N_7589,N_4195,N_5474);
nand U7590 (N_7590,N_4891,N_3343);
nor U7591 (N_7591,N_3824,N_5067);
nor U7592 (N_7592,N_4968,N_4680);
nor U7593 (N_7593,N_5732,N_3123);
nand U7594 (N_7594,N_4327,N_5788);
nor U7595 (N_7595,N_3859,N_5820);
nand U7596 (N_7596,N_3562,N_4373);
xnor U7597 (N_7597,N_4493,N_4711);
nor U7598 (N_7598,N_5278,N_3637);
nor U7599 (N_7599,N_3348,N_4272);
nor U7600 (N_7600,N_4419,N_3589);
or U7601 (N_7601,N_5249,N_4146);
nor U7602 (N_7602,N_3948,N_4213);
xor U7603 (N_7603,N_4333,N_5454);
xnor U7604 (N_7604,N_5229,N_3281);
and U7605 (N_7605,N_4999,N_3736);
nor U7606 (N_7606,N_3792,N_3874);
xor U7607 (N_7607,N_4488,N_3796);
and U7608 (N_7608,N_4337,N_5641);
nor U7609 (N_7609,N_3168,N_5615);
xor U7610 (N_7610,N_5146,N_4849);
xnor U7611 (N_7611,N_3476,N_5304);
nor U7612 (N_7612,N_3782,N_4743);
xnor U7613 (N_7613,N_3149,N_3609);
nor U7614 (N_7614,N_3345,N_5358);
nor U7615 (N_7615,N_3189,N_4748);
nand U7616 (N_7616,N_5353,N_5628);
or U7617 (N_7617,N_4799,N_4037);
or U7618 (N_7618,N_4429,N_5562);
nand U7619 (N_7619,N_5783,N_4276);
or U7620 (N_7620,N_3470,N_4641);
or U7621 (N_7621,N_5122,N_4720);
or U7622 (N_7622,N_3266,N_5302);
xor U7623 (N_7623,N_5345,N_3314);
and U7624 (N_7624,N_4901,N_3083);
or U7625 (N_7625,N_5877,N_4115);
nand U7626 (N_7626,N_4260,N_4650);
or U7627 (N_7627,N_3173,N_5578);
and U7628 (N_7628,N_5446,N_3775);
nor U7629 (N_7629,N_4671,N_5556);
nor U7630 (N_7630,N_4151,N_5884);
nand U7631 (N_7631,N_5482,N_3737);
nor U7632 (N_7632,N_5963,N_5784);
nand U7633 (N_7633,N_4791,N_5938);
nand U7634 (N_7634,N_5530,N_5869);
nand U7635 (N_7635,N_4697,N_3043);
or U7636 (N_7636,N_5920,N_3943);
nand U7637 (N_7637,N_3505,N_5907);
xor U7638 (N_7638,N_4453,N_3832);
and U7639 (N_7639,N_3631,N_4765);
nor U7640 (N_7640,N_3258,N_3059);
and U7641 (N_7641,N_5933,N_5328);
nand U7642 (N_7642,N_4732,N_5459);
or U7643 (N_7643,N_5390,N_5077);
or U7644 (N_7644,N_3304,N_5590);
or U7645 (N_7645,N_4648,N_3348);
and U7646 (N_7646,N_5176,N_3401);
nand U7647 (N_7647,N_5972,N_5599);
and U7648 (N_7648,N_3230,N_3270);
and U7649 (N_7649,N_4231,N_3605);
or U7650 (N_7650,N_4474,N_3588);
nand U7651 (N_7651,N_3605,N_3736);
nand U7652 (N_7652,N_5171,N_4841);
nor U7653 (N_7653,N_4356,N_3681);
xor U7654 (N_7654,N_5902,N_4223);
xnor U7655 (N_7655,N_5036,N_4860);
or U7656 (N_7656,N_5840,N_3674);
nand U7657 (N_7657,N_5595,N_4104);
xor U7658 (N_7658,N_3679,N_4907);
or U7659 (N_7659,N_3539,N_4600);
and U7660 (N_7660,N_5000,N_4840);
or U7661 (N_7661,N_3455,N_5580);
and U7662 (N_7662,N_3817,N_3093);
or U7663 (N_7663,N_4131,N_5416);
and U7664 (N_7664,N_3506,N_4232);
nor U7665 (N_7665,N_3173,N_5562);
or U7666 (N_7666,N_5319,N_5265);
nor U7667 (N_7667,N_5158,N_3008);
and U7668 (N_7668,N_5989,N_3832);
and U7669 (N_7669,N_4754,N_4916);
nand U7670 (N_7670,N_3805,N_3154);
xnor U7671 (N_7671,N_3936,N_5682);
or U7672 (N_7672,N_4518,N_5405);
nand U7673 (N_7673,N_4661,N_3583);
and U7674 (N_7674,N_3654,N_4014);
and U7675 (N_7675,N_4406,N_3145);
xnor U7676 (N_7676,N_4398,N_5356);
and U7677 (N_7677,N_4606,N_3345);
or U7678 (N_7678,N_4308,N_3631);
or U7679 (N_7679,N_3844,N_5458);
nand U7680 (N_7680,N_5224,N_5840);
or U7681 (N_7681,N_4522,N_3808);
nor U7682 (N_7682,N_4814,N_3807);
nand U7683 (N_7683,N_3470,N_5860);
nor U7684 (N_7684,N_3689,N_4844);
and U7685 (N_7685,N_4834,N_5160);
and U7686 (N_7686,N_3585,N_3724);
or U7687 (N_7687,N_4344,N_5906);
or U7688 (N_7688,N_3128,N_5219);
or U7689 (N_7689,N_4526,N_3881);
xnor U7690 (N_7690,N_5167,N_3479);
and U7691 (N_7691,N_4197,N_5482);
nor U7692 (N_7692,N_3252,N_5085);
xor U7693 (N_7693,N_3968,N_3651);
or U7694 (N_7694,N_5728,N_3516);
nor U7695 (N_7695,N_4577,N_3042);
nor U7696 (N_7696,N_5054,N_4627);
nand U7697 (N_7697,N_3231,N_3780);
or U7698 (N_7698,N_3809,N_5757);
xnor U7699 (N_7699,N_5149,N_5103);
or U7700 (N_7700,N_5490,N_3637);
and U7701 (N_7701,N_3616,N_4794);
nor U7702 (N_7702,N_5070,N_5281);
and U7703 (N_7703,N_3341,N_5578);
nand U7704 (N_7704,N_3326,N_3681);
nand U7705 (N_7705,N_5491,N_5205);
xor U7706 (N_7706,N_3392,N_5254);
and U7707 (N_7707,N_4378,N_4934);
and U7708 (N_7708,N_3374,N_4396);
nand U7709 (N_7709,N_4805,N_4516);
or U7710 (N_7710,N_3907,N_4053);
and U7711 (N_7711,N_3700,N_5603);
and U7712 (N_7712,N_4039,N_5202);
xnor U7713 (N_7713,N_3647,N_5140);
and U7714 (N_7714,N_3487,N_5253);
and U7715 (N_7715,N_5439,N_3011);
nor U7716 (N_7716,N_4551,N_5141);
and U7717 (N_7717,N_3681,N_3514);
nand U7718 (N_7718,N_4727,N_4876);
nand U7719 (N_7719,N_5407,N_3148);
nand U7720 (N_7720,N_5439,N_5367);
or U7721 (N_7721,N_4840,N_5666);
nor U7722 (N_7722,N_5014,N_3948);
nand U7723 (N_7723,N_4031,N_3999);
xnor U7724 (N_7724,N_5965,N_5138);
xnor U7725 (N_7725,N_3481,N_3668);
or U7726 (N_7726,N_4304,N_4699);
nand U7727 (N_7727,N_4323,N_5213);
and U7728 (N_7728,N_4406,N_3614);
nor U7729 (N_7729,N_5557,N_4643);
nand U7730 (N_7730,N_4889,N_3511);
and U7731 (N_7731,N_3023,N_3811);
xnor U7732 (N_7732,N_3555,N_4462);
or U7733 (N_7733,N_3218,N_3970);
or U7734 (N_7734,N_5185,N_4205);
and U7735 (N_7735,N_3904,N_5147);
or U7736 (N_7736,N_3284,N_5362);
or U7737 (N_7737,N_5692,N_4908);
or U7738 (N_7738,N_5630,N_3236);
and U7739 (N_7739,N_5014,N_4268);
nor U7740 (N_7740,N_3307,N_3386);
xor U7741 (N_7741,N_5480,N_5114);
nor U7742 (N_7742,N_5833,N_3949);
and U7743 (N_7743,N_4928,N_5710);
nor U7744 (N_7744,N_3524,N_4945);
and U7745 (N_7745,N_5945,N_5660);
and U7746 (N_7746,N_4514,N_3422);
and U7747 (N_7747,N_5398,N_3146);
xor U7748 (N_7748,N_4763,N_4873);
or U7749 (N_7749,N_5653,N_4903);
and U7750 (N_7750,N_4250,N_3548);
or U7751 (N_7751,N_5765,N_5651);
and U7752 (N_7752,N_5390,N_4934);
nand U7753 (N_7753,N_5947,N_3004);
nand U7754 (N_7754,N_4848,N_5251);
nor U7755 (N_7755,N_5839,N_3033);
nand U7756 (N_7756,N_5859,N_3157);
xnor U7757 (N_7757,N_4677,N_4137);
nor U7758 (N_7758,N_4171,N_3616);
and U7759 (N_7759,N_4632,N_4866);
nor U7760 (N_7760,N_3431,N_3106);
and U7761 (N_7761,N_3962,N_5586);
xnor U7762 (N_7762,N_5466,N_3427);
and U7763 (N_7763,N_3880,N_5554);
or U7764 (N_7764,N_4418,N_3112);
nand U7765 (N_7765,N_5679,N_3228);
nor U7766 (N_7766,N_5972,N_5283);
and U7767 (N_7767,N_4909,N_3703);
nor U7768 (N_7768,N_4171,N_3274);
or U7769 (N_7769,N_3241,N_4110);
nor U7770 (N_7770,N_3771,N_5809);
nor U7771 (N_7771,N_3002,N_4493);
nand U7772 (N_7772,N_4155,N_3390);
nor U7773 (N_7773,N_5437,N_5773);
nor U7774 (N_7774,N_5967,N_3559);
xnor U7775 (N_7775,N_5705,N_5610);
nand U7776 (N_7776,N_5382,N_5675);
nand U7777 (N_7777,N_5183,N_5295);
xor U7778 (N_7778,N_5497,N_3380);
nor U7779 (N_7779,N_5089,N_3954);
nor U7780 (N_7780,N_4194,N_5714);
nand U7781 (N_7781,N_4525,N_5663);
and U7782 (N_7782,N_5822,N_3897);
or U7783 (N_7783,N_5906,N_5213);
nor U7784 (N_7784,N_3547,N_4785);
xor U7785 (N_7785,N_4596,N_5086);
and U7786 (N_7786,N_3409,N_3934);
xnor U7787 (N_7787,N_5916,N_4805);
nor U7788 (N_7788,N_3890,N_4631);
nor U7789 (N_7789,N_4584,N_5226);
nor U7790 (N_7790,N_3232,N_4033);
xnor U7791 (N_7791,N_5280,N_5389);
nand U7792 (N_7792,N_4384,N_3013);
or U7793 (N_7793,N_5510,N_5787);
or U7794 (N_7794,N_3452,N_4265);
nand U7795 (N_7795,N_5100,N_5782);
or U7796 (N_7796,N_3620,N_3084);
nor U7797 (N_7797,N_4888,N_4108);
or U7798 (N_7798,N_5826,N_5997);
nor U7799 (N_7799,N_5022,N_5462);
xnor U7800 (N_7800,N_5505,N_5657);
or U7801 (N_7801,N_3704,N_3321);
and U7802 (N_7802,N_4837,N_3695);
and U7803 (N_7803,N_5565,N_5721);
or U7804 (N_7804,N_3098,N_4539);
xor U7805 (N_7805,N_5316,N_4970);
nor U7806 (N_7806,N_5643,N_3502);
or U7807 (N_7807,N_5138,N_5538);
or U7808 (N_7808,N_3129,N_4075);
nand U7809 (N_7809,N_5569,N_4362);
and U7810 (N_7810,N_5791,N_5530);
nand U7811 (N_7811,N_3093,N_5833);
and U7812 (N_7812,N_5560,N_4617);
and U7813 (N_7813,N_4725,N_5396);
xor U7814 (N_7814,N_3847,N_5873);
xor U7815 (N_7815,N_3910,N_4741);
xor U7816 (N_7816,N_3656,N_3945);
nor U7817 (N_7817,N_3519,N_3488);
nand U7818 (N_7818,N_3855,N_3836);
nand U7819 (N_7819,N_4588,N_3411);
nand U7820 (N_7820,N_5859,N_3968);
nor U7821 (N_7821,N_4485,N_5342);
xnor U7822 (N_7822,N_5322,N_4251);
nand U7823 (N_7823,N_4702,N_4994);
nor U7824 (N_7824,N_4198,N_4404);
or U7825 (N_7825,N_3387,N_4070);
xor U7826 (N_7826,N_3550,N_4673);
nor U7827 (N_7827,N_3843,N_5231);
or U7828 (N_7828,N_5150,N_4266);
nand U7829 (N_7829,N_3143,N_4914);
xor U7830 (N_7830,N_5362,N_4141);
nor U7831 (N_7831,N_5591,N_5795);
xor U7832 (N_7832,N_3443,N_3153);
xnor U7833 (N_7833,N_5748,N_4249);
nand U7834 (N_7834,N_5705,N_5571);
or U7835 (N_7835,N_5254,N_4186);
and U7836 (N_7836,N_3252,N_4886);
nor U7837 (N_7837,N_5297,N_4404);
nand U7838 (N_7838,N_5789,N_5552);
or U7839 (N_7839,N_4343,N_3006);
nand U7840 (N_7840,N_5707,N_5712);
nand U7841 (N_7841,N_4870,N_5969);
nand U7842 (N_7842,N_4999,N_3147);
xnor U7843 (N_7843,N_5734,N_3015);
nor U7844 (N_7844,N_3842,N_3492);
and U7845 (N_7845,N_3293,N_3261);
nor U7846 (N_7846,N_3714,N_5344);
and U7847 (N_7847,N_5291,N_4997);
nor U7848 (N_7848,N_5733,N_4599);
xnor U7849 (N_7849,N_5352,N_5599);
nor U7850 (N_7850,N_5367,N_4509);
and U7851 (N_7851,N_5134,N_5670);
xor U7852 (N_7852,N_4245,N_4432);
or U7853 (N_7853,N_5856,N_5213);
nor U7854 (N_7854,N_4735,N_3365);
nand U7855 (N_7855,N_5376,N_3820);
xor U7856 (N_7856,N_4007,N_5601);
and U7857 (N_7857,N_5801,N_5610);
nor U7858 (N_7858,N_3642,N_5939);
and U7859 (N_7859,N_3641,N_5185);
or U7860 (N_7860,N_4389,N_3663);
nor U7861 (N_7861,N_5452,N_5274);
and U7862 (N_7862,N_3365,N_5728);
and U7863 (N_7863,N_4791,N_5129);
nor U7864 (N_7864,N_5805,N_3417);
nand U7865 (N_7865,N_3848,N_4478);
nor U7866 (N_7866,N_3446,N_5195);
nand U7867 (N_7867,N_3634,N_3240);
and U7868 (N_7868,N_5530,N_5735);
nor U7869 (N_7869,N_3054,N_3525);
xor U7870 (N_7870,N_3739,N_4277);
nand U7871 (N_7871,N_3971,N_4718);
nor U7872 (N_7872,N_5065,N_3741);
nand U7873 (N_7873,N_3591,N_5230);
nand U7874 (N_7874,N_5911,N_5955);
nand U7875 (N_7875,N_5412,N_3389);
xor U7876 (N_7876,N_3025,N_5106);
nand U7877 (N_7877,N_4391,N_5941);
nand U7878 (N_7878,N_4869,N_5088);
nand U7879 (N_7879,N_3296,N_3611);
nor U7880 (N_7880,N_4900,N_4578);
and U7881 (N_7881,N_4711,N_4307);
nand U7882 (N_7882,N_5314,N_5445);
xnor U7883 (N_7883,N_4767,N_3939);
xor U7884 (N_7884,N_4882,N_5857);
nor U7885 (N_7885,N_4560,N_3825);
nand U7886 (N_7886,N_4199,N_3378);
xor U7887 (N_7887,N_5841,N_5695);
nor U7888 (N_7888,N_3338,N_4184);
or U7889 (N_7889,N_3495,N_3473);
nor U7890 (N_7890,N_4819,N_4541);
nand U7891 (N_7891,N_5512,N_4513);
nand U7892 (N_7892,N_4007,N_5497);
and U7893 (N_7893,N_5541,N_4391);
and U7894 (N_7894,N_5005,N_5173);
nor U7895 (N_7895,N_3871,N_4608);
nor U7896 (N_7896,N_3865,N_5246);
and U7897 (N_7897,N_3937,N_3832);
nand U7898 (N_7898,N_3196,N_5320);
nand U7899 (N_7899,N_5837,N_5045);
xnor U7900 (N_7900,N_4068,N_5717);
nor U7901 (N_7901,N_4020,N_4843);
or U7902 (N_7902,N_4961,N_3941);
xor U7903 (N_7903,N_5613,N_4293);
xnor U7904 (N_7904,N_5848,N_4264);
or U7905 (N_7905,N_4596,N_5930);
nor U7906 (N_7906,N_5636,N_5052);
xor U7907 (N_7907,N_5323,N_5423);
nor U7908 (N_7908,N_3346,N_3152);
and U7909 (N_7909,N_5899,N_3269);
nor U7910 (N_7910,N_3518,N_3411);
or U7911 (N_7911,N_4841,N_3384);
and U7912 (N_7912,N_4597,N_4536);
or U7913 (N_7913,N_5349,N_4675);
nand U7914 (N_7914,N_4444,N_3207);
xnor U7915 (N_7915,N_3757,N_4138);
nor U7916 (N_7916,N_3655,N_5772);
xor U7917 (N_7917,N_4927,N_3385);
or U7918 (N_7918,N_3103,N_5138);
nand U7919 (N_7919,N_5041,N_3873);
xor U7920 (N_7920,N_5890,N_4290);
or U7921 (N_7921,N_5489,N_4978);
nor U7922 (N_7922,N_4073,N_3147);
xnor U7923 (N_7923,N_3791,N_3916);
or U7924 (N_7924,N_3158,N_4083);
nor U7925 (N_7925,N_5312,N_3437);
nor U7926 (N_7926,N_5485,N_5615);
xor U7927 (N_7927,N_4202,N_4749);
and U7928 (N_7928,N_3168,N_4602);
or U7929 (N_7929,N_4553,N_3054);
nand U7930 (N_7930,N_3367,N_4648);
or U7931 (N_7931,N_3490,N_5612);
or U7932 (N_7932,N_4804,N_4591);
or U7933 (N_7933,N_5875,N_5933);
and U7934 (N_7934,N_3811,N_4538);
nor U7935 (N_7935,N_4579,N_4407);
xor U7936 (N_7936,N_5704,N_3510);
and U7937 (N_7937,N_4636,N_3882);
or U7938 (N_7938,N_5458,N_4388);
or U7939 (N_7939,N_5338,N_4135);
xnor U7940 (N_7940,N_3144,N_3055);
xor U7941 (N_7941,N_3146,N_3201);
nand U7942 (N_7942,N_4495,N_5433);
nand U7943 (N_7943,N_4303,N_5346);
and U7944 (N_7944,N_3196,N_5576);
and U7945 (N_7945,N_5619,N_5448);
nor U7946 (N_7946,N_3357,N_5640);
nand U7947 (N_7947,N_3984,N_4870);
or U7948 (N_7948,N_4339,N_5103);
nor U7949 (N_7949,N_4064,N_5999);
and U7950 (N_7950,N_3089,N_5790);
xnor U7951 (N_7951,N_4660,N_4166);
and U7952 (N_7952,N_3489,N_4233);
xnor U7953 (N_7953,N_4470,N_3004);
xor U7954 (N_7954,N_4960,N_5203);
and U7955 (N_7955,N_5195,N_5223);
and U7956 (N_7956,N_5596,N_3381);
nor U7957 (N_7957,N_3871,N_5280);
and U7958 (N_7958,N_4481,N_5493);
and U7959 (N_7959,N_4602,N_3727);
and U7960 (N_7960,N_5999,N_4781);
and U7961 (N_7961,N_3372,N_3655);
and U7962 (N_7962,N_5692,N_3347);
or U7963 (N_7963,N_4710,N_4157);
or U7964 (N_7964,N_3276,N_4215);
xor U7965 (N_7965,N_4570,N_4006);
xnor U7966 (N_7966,N_3989,N_4536);
nor U7967 (N_7967,N_4874,N_5435);
nor U7968 (N_7968,N_4863,N_3268);
nor U7969 (N_7969,N_3543,N_5714);
and U7970 (N_7970,N_5966,N_5133);
or U7971 (N_7971,N_4805,N_5175);
xor U7972 (N_7972,N_4966,N_3904);
and U7973 (N_7973,N_5936,N_5402);
and U7974 (N_7974,N_5755,N_4168);
and U7975 (N_7975,N_4104,N_5967);
or U7976 (N_7976,N_3235,N_4975);
and U7977 (N_7977,N_3840,N_4852);
nand U7978 (N_7978,N_5623,N_4914);
nor U7979 (N_7979,N_3398,N_3375);
nand U7980 (N_7980,N_3162,N_4174);
nor U7981 (N_7981,N_4134,N_5477);
or U7982 (N_7982,N_4156,N_3570);
xnor U7983 (N_7983,N_5104,N_3410);
and U7984 (N_7984,N_5223,N_3537);
nor U7985 (N_7985,N_4727,N_5561);
nand U7986 (N_7986,N_5677,N_5160);
xnor U7987 (N_7987,N_5164,N_5605);
nand U7988 (N_7988,N_4760,N_4553);
and U7989 (N_7989,N_5071,N_3243);
nand U7990 (N_7990,N_5523,N_4019);
or U7991 (N_7991,N_5079,N_3960);
and U7992 (N_7992,N_5329,N_5912);
nor U7993 (N_7993,N_5137,N_5184);
and U7994 (N_7994,N_3086,N_4632);
or U7995 (N_7995,N_4620,N_3401);
nand U7996 (N_7996,N_4646,N_3212);
xor U7997 (N_7997,N_4697,N_4761);
nor U7998 (N_7998,N_5349,N_4141);
xnor U7999 (N_7999,N_4598,N_5832);
nor U8000 (N_8000,N_5096,N_3538);
xnor U8001 (N_8001,N_5419,N_5997);
nor U8002 (N_8002,N_3594,N_5000);
xnor U8003 (N_8003,N_5271,N_3584);
and U8004 (N_8004,N_4933,N_4532);
xnor U8005 (N_8005,N_4544,N_4598);
nand U8006 (N_8006,N_5761,N_3709);
nand U8007 (N_8007,N_4279,N_5801);
xor U8008 (N_8008,N_3859,N_3733);
nor U8009 (N_8009,N_4460,N_5497);
or U8010 (N_8010,N_5174,N_5116);
nor U8011 (N_8011,N_5152,N_3063);
xnor U8012 (N_8012,N_4132,N_4728);
xnor U8013 (N_8013,N_4655,N_5005);
xor U8014 (N_8014,N_5891,N_5950);
nand U8015 (N_8015,N_3538,N_3233);
nor U8016 (N_8016,N_4531,N_5905);
or U8017 (N_8017,N_4711,N_5201);
nand U8018 (N_8018,N_4498,N_3320);
or U8019 (N_8019,N_4836,N_3948);
xnor U8020 (N_8020,N_5233,N_4409);
and U8021 (N_8021,N_5241,N_3894);
nor U8022 (N_8022,N_4344,N_5078);
and U8023 (N_8023,N_4456,N_4051);
or U8024 (N_8024,N_3221,N_5871);
nor U8025 (N_8025,N_3132,N_3930);
and U8026 (N_8026,N_5666,N_5865);
and U8027 (N_8027,N_3996,N_5888);
nor U8028 (N_8028,N_3331,N_4008);
nor U8029 (N_8029,N_3611,N_3865);
nor U8030 (N_8030,N_3072,N_5208);
nand U8031 (N_8031,N_4933,N_4362);
nor U8032 (N_8032,N_4232,N_5971);
nor U8033 (N_8033,N_3929,N_3361);
and U8034 (N_8034,N_3979,N_3658);
xor U8035 (N_8035,N_3083,N_4032);
nand U8036 (N_8036,N_5275,N_5040);
nor U8037 (N_8037,N_3087,N_3584);
nor U8038 (N_8038,N_5021,N_3305);
nor U8039 (N_8039,N_5658,N_4127);
nand U8040 (N_8040,N_3504,N_3075);
nand U8041 (N_8041,N_3772,N_4139);
nand U8042 (N_8042,N_4510,N_5475);
or U8043 (N_8043,N_4582,N_3936);
nand U8044 (N_8044,N_4506,N_4719);
and U8045 (N_8045,N_5659,N_3972);
nor U8046 (N_8046,N_3318,N_5253);
nand U8047 (N_8047,N_3439,N_4005);
nor U8048 (N_8048,N_3012,N_5503);
or U8049 (N_8049,N_5883,N_4694);
nor U8050 (N_8050,N_4736,N_3675);
xor U8051 (N_8051,N_4382,N_3586);
or U8052 (N_8052,N_5854,N_5288);
or U8053 (N_8053,N_3989,N_3073);
xnor U8054 (N_8054,N_4466,N_4436);
nor U8055 (N_8055,N_5357,N_5034);
or U8056 (N_8056,N_4635,N_3431);
nand U8057 (N_8057,N_5634,N_3324);
and U8058 (N_8058,N_5938,N_4861);
and U8059 (N_8059,N_5617,N_3763);
nor U8060 (N_8060,N_4091,N_4007);
or U8061 (N_8061,N_4969,N_3619);
or U8062 (N_8062,N_3048,N_5832);
xor U8063 (N_8063,N_5767,N_3647);
xor U8064 (N_8064,N_4466,N_3629);
xor U8065 (N_8065,N_4804,N_4138);
and U8066 (N_8066,N_3102,N_5620);
or U8067 (N_8067,N_3560,N_3183);
and U8068 (N_8068,N_4648,N_5577);
nand U8069 (N_8069,N_3015,N_4630);
nand U8070 (N_8070,N_5770,N_5028);
xor U8071 (N_8071,N_3988,N_4407);
xnor U8072 (N_8072,N_5237,N_4507);
and U8073 (N_8073,N_3493,N_5965);
nor U8074 (N_8074,N_4545,N_5312);
xnor U8075 (N_8075,N_4549,N_5424);
xnor U8076 (N_8076,N_4994,N_3537);
nand U8077 (N_8077,N_4032,N_3484);
and U8078 (N_8078,N_3897,N_5142);
or U8079 (N_8079,N_3124,N_5016);
or U8080 (N_8080,N_5776,N_3718);
or U8081 (N_8081,N_5706,N_5456);
xor U8082 (N_8082,N_4169,N_5097);
nand U8083 (N_8083,N_4428,N_5164);
nand U8084 (N_8084,N_5005,N_4519);
nand U8085 (N_8085,N_5792,N_5292);
or U8086 (N_8086,N_4252,N_3366);
or U8087 (N_8087,N_5066,N_4988);
and U8088 (N_8088,N_3111,N_5887);
xor U8089 (N_8089,N_5339,N_3172);
and U8090 (N_8090,N_5666,N_5783);
nand U8091 (N_8091,N_5598,N_4692);
nand U8092 (N_8092,N_5235,N_5832);
and U8093 (N_8093,N_3218,N_4837);
and U8094 (N_8094,N_3991,N_4314);
xor U8095 (N_8095,N_3803,N_4233);
or U8096 (N_8096,N_5925,N_3804);
xor U8097 (N_8097,N_5669,N_3465);
or U8098 (N_8098,N_3833,N_3607);
or U8099 (N_8099,N_3151,N_3154);
xor U8100 (N_8100,N_3227,N_4402);
xnor U8101 (N_8101,N_4499,N_5271);
and U8102 (N_8102,N_3338,N_5249);
nor U8103 (N_8103,N_4337,N_5035);
nor U8104 (N_8104,N_4022,N_3325);
and U8105 (N_8105,N_3894,N_5086);
xor U8106 (N_8106,N_4129,N_4501);
or U8107 (N_8107,N_3966,N_3299);
or U8108 (N_8108,N_5295,N_5953);
nand U8109 (N_8109,N_4279,N_3045);
or U8110 (N_8110,N_5711,N_5725);
xor U8111 (N_8111,N_4788,N_5732);
nor U8112 (N_8112,N_3650,N_5739);
or U8113 (N_8113,N_3117,N_4377);
nand U8114 (N_8114,N_4834,N_4525);
xnor U8115 (N_8115,N_4051,N_3338);
or U8116 (N_8116,N_3040,N_3435);
and U8117 (N_8117,N_5700,N_3630);
xor U8118 (N_8118,N_4220,N_4365);
xor U8119 (N_8119,N_3226,N_5307);
nor U8120 (N_8120,N_3530,N_3392);
and U8121 (N_8121,N_4988,N_4420);
and U8122 (N_8122,N_3493,N_3974);
and U8123 (N_8123,N_4218,N_4648);
xnor U8124 (N_8124,N_4975,N_3872);
and U8125 (N_8125,N_4862,N_3412);
and U8126 (N_8126,N_4903,N_3774);
or U8127 (N_8127,N_5516,N_5213);
and U8128 (N_8128,N_3341,N_3009);
nor U8129 (N_8129,N_5773,N_3398);
nor U8130 (N_8130,N_3802,N_4755);
nor U8131 (N_8131,N_5766,N_4680);
nand U8132 (N_8132,N_4873,N_4396);
xor U8133 (N_8133,N_5418,N_3891);
nand U8134 (N_8134,N_3979,N_3143);
xor U8135 (N_8135,N_3913,N_3012);
xnor U8136 (N_8136,N_4340,N_3405);
xor U8137 (N_8137,N_5750,N_4491);
nor U8138 (N_8138,N_3128,N_5780);
xor U8139 (N_8139,N_3479,N_4421);
xor U8140 (N_8140,N_5506,N_3635);
and U8141 (N_8141,N_3435,N_4854);
nor U8142 (N_8142,N_5091,N_4243);
nand U8143 (N_8143,N_4644,N_5595);
and U8144 (N_8144,N_5213,N_5525);
xor U8145 (N_8145,N_3478,N_5545);
xnor U8146 (N_8146,N_5859,N_5360);
xor U8147 (N_8147,N_4206,N_3952);
nand U8148 (N_8148,N_3747,N_4787);
and U8149 (N_8149,N_5912,N_4789);
xor U8150 (N_8150,N_3458,N_5285);
nand U8151 (N_8151,N_5433,N_4986);
nor U8152 (N_8152,N_4369,N_3124);
or U8153 (N_8153,N_4445,N_5377);
or U8154 (N_8154,N_4369,N_5136);
nand U8155 (N_8155,N_3113,N_5279);
nand U8156 (N_8156,N_3767,N_5001);
nand U8157 (N_8157,N_4046,N_5957);
or U8158 (N_8158,N_4432,N_4989);
or U8159 (N_8159,N_5475,N_3720);
or U8160 (N_8160,N_3155,N_4507);
xnor U8161 (N_8161,N_4007,N_4545);
nand U8162 (N_8162,N_3464,N_5345);
or U8163 (N_8163,N_4127,N_4826);
xnor U8164 (N_8164,N_5422,N_5673);
and U8165 (N_8165,N_5549,N_3866);
and U8166 (N_8166,N_3146,N_5045);
nand U8167 (N_8167,N_4602,N_4523);
nor U8168 (N_8168,N_3034,N_5905);
nor U8169 (N_8169,N_5256,N_5068);
nand U8170 (N_8170,N_4370,N_3751);
and U8171 (N_8171,N_3113,N_4056);
and U8172 (N_8172,N_5487,N_3963);
nor U8173 (N_8173,N_3764,N_4206);
xor U8174 (N_8174,N_4210,N_4363);
nand U8175 (N_8175,N_3327,N_3386);
xor U8176 (N_8176,N_4880,N_5481);
nand U8177 (N_8177,N_4475,N_5899);
or U8178 (N_8178,N_3462,N_5890);
nand U8179 (N_8179,N_5633,N_3790);
and U8180 (N_8180,N_4866,N_3810);
xnor U8181 (N_8181,N_4614,N_3175);
and U8182 (N_8182,N_4708,N_3576);
or U8183 (N_8183,N_4644,N_3208);
xnor U8184 (N_8184,N_3378,N_4790);
nor U8185 (N_8185,N_5020,N_5511);
nand U8186 (N_8186,N_3166,N_4381);
or U8187 (N_8187,N_5242,N_3336);
nand U8188 (N_8188,N_5454,N_3188);
nor U8189 (N_8189,N_3468,N_3045);
or U8190 (N_8190,N_4115,N_4400);
or U8191 (N_8191,N_4267,N_3764);
and U8192 (N_8192,N_5771,N_4483);
or U8193 (N_8193,N_5942,N_5050);
and U8194 (N_8194,N_4067,N_5277);
and U8195 (N_8195,N_3000,N_4363);
or U8196 (N_8196,N_3782,N_5483);
or U8197 (N_8197,N_5706,N_3655);
or U8198 (N_8198,N_4154,N_3488);
nor U8199 (N_8199,N_5976,N_5407);
and U8200 (N_8200,N_5289,N_5714);
and U8201 (N_8201,N_3702,N_4689);
nand U8202 (N_8202,N_3991,N_3019);
and U8203 (N_8203,N_3067,N_4750);
xnor U8204 (N_8204,N_3457,N_3689);
and U8205 (N_8205,N_5199,N_3276);
or U8206 (N_8206,N_4282,N_4162);
xor U8207 (N_8207,N_5458,N_4435);
nor U8208 (N_8208,N_4456,N_5852);
nand U8209 (N_8209,N_5919,N_3534);
and U8210 (N_8210,N_5608,N_5251);
nand U8211 (N_8211,N_5566,N_4439);
and U8212 (N_8212,N_3101,N_4155);
nand U8213 (N_8213,N_5483,N_3491);
or U8214 (N_8214,N_5737,N_3222);
and U8215 (N_8215,N_4986,N_5475);
xnor U8216 (N_8216,N_5482,N_5405);
xnor U8217 (N_8217,N_4343,N_3249);
and U8218 (N_8218,N_4965,N_3717);
xor U8219 (N_8219,N_4663,N_5460);
nand U8220 (N_8220,N_5307,N_4491);
or U8221 (N_8221,N_3751,N_4564);
nor U8222 (N_8222,N_4042,N_3274);
xor U8223 (N_8223,N_3807,N_5340);
and U8224 (N_8224,N_4327,N_3132);
or U8225 (N_8225,N_4893,N_5753);
or U8226 (N_8226,N_5037,N_5032);
and U8227 (N_8227,N_5574,N_3689);
or U8228 (N_8228,N_4735,N_5031);
xnor U8229 (N_8229,N_3399,N_3482);
nand U8230 (N_8230,N_3145,N_5355);
nor U8231 (N_8231,N_4534,N_3839);
xnor U8232 (N_8232,N_5631,N_5467);
xor U8233 (N_8233,N_4115,N_5138);
or U8234 (N_8234,N_3963,N_3642);
xor U8235 (N_8235,N_4538,N_3304);
and U8236 (N_8236,N_5070,N_3975);
or U8237 (N_8237,N_3671,N_5642);
or U8238 (N_8238,N_5849,N_4894);
nand U8239 (N_8239,N_5215,N_4755);
nor U8240 (N_8240,N_3656,N_3620);
nand U8241 (N_8241,N_3562,N_5925);
nand U8242 (N_8242,N_3257,N_4094);
and U8243 (N_8243,N_5293,N_4582);
or U8244 (N_8244,N_5893,N_4548);
or U8245 (N_8245,N_5007,N_3518);
and U8246 (N_8246,N_4240,N_3350);
nand U8247 (N_8247,N_3201,N_5337);
or U8248 (N_8248,N_5136,N_5636);
and U8249 (N_8249,N_5224,N_5136);
and U8250 (N_8250,N_5059,N_4150);
nand U8251 (N_8251,N_5229,N_4099);
or U8252 (N_8252,N_5648,N_3913);
or U8253 (N_8253,N_3166,N_5043);
nand U8254 (N_8254,N_4853,N_4552);
nor U8255 (N_8255,N_3109,N_5459);
and U8256 (N_8256,N_5429,N_4881);
or U8257 (N_8257,N_3866,N_4816);
and U8258 (N_8258,N_4899,N_5416);
or U8259 (N_8259,N_5825,N_4034);
or U8260 (N_8260,N_4280,N_3061);
and U8261 (N_8261,N_3376,N_5023);
xnor U8262 (N_8262,N_3235,N_5701);
nand U8263 (N_8263,N_3446,N_5814);
and U8264 (N_8264,N_4204,N_3926);
nor U8265 (N_8265,N_5477,N_4902);
and U8266 (N_8266,N_4029,N_5901);
nor U8267 (N_8267,N_4503,N_5092);
nor U8268 (N_8268,N_5870,N_4834);
or U8269 (N_8269,N_5202,N_4542);
and U8270 (N_8270,N_3401,N_4510);
and U8271 (N_8271,N_5116,N_3521);
or U8272 (N_8272,N_3205,N_4682);
xor U8273 (N_8273,N_5747,N_4966);
and U8274 (N_8274,N_3550,N_4163);
and U8275 (N_8275,N_3580,N_4926);
and U8276 (N_8276,N_5460,N_3584);
and U8277 (N_8277,N_5267,N_4891);
xnor U8278 (N_8278,N_4660,N_4920);
nand U8279 (N_8279,N_3908,N_3539);
nand U8280 (N_8280,N_4548,N_5447);
nand U8281 (N_8281,N_5666,N_4682);
nor U8282 (N_8282,N_4509,N_3786);
xor U8283 (N_8283,N_5570,N_5569);
nor U8284 (N_8284,N_4467,N_4689);
nor U8285 (N_8285,N_3137,N_3305);
xor U8286 (N_8286,N_3263,N_4580);
xnor U8287 (N_8287,N_3191,N_5231);
or U8288 (N_8288,N_4580,N_4983);
or U8289 (N_8289,N_4255,N_5653);
nor U8290 (N_8290,N_5551,N_5081);
nand U8291 (N_8291,N_3355,N_4429);
and U8292 (N_8292,N_5679,N_4503);
nor U8293 (N_8293,N_3771,N_3871);
or U8294 (N_8294,N_5162,N_4057);
xor U8295 (N_8295,N_3698,N_3148);
nor U8296 (N_8296,N_3621,N_3313);
and U8297 (N_8297,N_5304,N_4839);
xnor U8298 (N_8298,N_5999,N_5510);
and U8299 (N_8299,N_5412,N_4423);
xor U8300 (N_8300,N_5526,N_3493);
nor U8301 (N_8301,N_4450,N_3968);
and U8302 (N_8302,N_3707,N_5271);
or U8303 (N_8303,N_3567,N_4992);
or U8304 (N_8304,N_3780,N_4537);
xnor U8305 (N_8305,N_4930,N_4154);
xor U8306 (N_8306,N_3601,N_4336);
and U8307 (N_8307,N_4702,N_5413);
xor U8308 (N_8308,N_5123,N_5140);
or U8309 (N_8309,N_5669,N_4256);
xor U8310 (N_8310,N_4834,N_4689);
nor U8311 (N_8311,N_5047,N_5768);
and U8312 (N_8312,N_5793,N_5206);
nand U8313 (N_8313,N_3213,N_3537);
nor U8314 (N_8314,N_3591,N_4088);
xor U8315 (N_8315,N_4455,N_5248);
and U8316 (N_8316,N_3020,N_5271);
or U8317 (N_8317,N_4994,N_5237);
xor U8318 (N_8318,N_3229,N_4213);
xnor U8319 (N_8319,N_3194,N_3677);
and U8320 (N_8320,N_4333,N_5069);
or U8321 (N_8321,N_4945,N_3736);
or U8322 (N_8322,N_5321,N_3051);
or U8323 (N_8323,N_3755,N_3607);
nor U8324 (N_8324,N_5839,N_3663);
or U8325 (N_8325,N_5370,N_3237);
nand U8326 (N_8326,N_5704,N_4278);
or U8327 (N_8327,N_4162,N_4305);
or U8328 (N_8328,N_5121,N_5233);
nand U8329 (N_8329,N_3437,N_3286);
or U8330 (N_8330,N_5453,N_3887);
nand U8331 (N_8331,N_4476,N_4397);
xor U8332 (N_8332,N_4930,N_3126);
nor U8333 (N_8333,N_5394,N_4506);
or U8334 (N_8334,N_4953,N_5007);
and U8335 (N_8335,N_5432,N_5599);
or U8336 (N_8336,N_4109,N_5063);
nand U8337 (N_8337,N_4315,N_4829);
nand U8338 (N_8338,N_5748,N_3942);
xor U8339 (N_8339,N_4576,N_4392);
and U8340 (N_8340,N_3601,N_4723);
and U8341 (N_8341,N_3113,N_5688);
or U8342 (N_8342,N_4258,N_4764);
and U8343 (N_8343,N_3149,N_5427);
nor U8344 (N_8344,N_3280,N_3721);
or U8345 (N_8345,N_4093,N_5424);
nor U8346 (N_8346,N_3180,N_5126);
or U8347 (N_8347,N_4654,N_3417);
nand U8348 (N_8348,N_3413,N_3042);
nor U8349 (N_8349,N_3600,N_4273);
or U8350 (N_8350,N_4731,N_3596);
nor U8351 (N_8351,N_4893,N_5588);
nor U8352 (N_8352,N_3690,N_5609);
or U8353 (N_8353,N_4031,N_5798);
nand U8354 (N_8354,N_5264,N_5615);
xor U8355 (N_8355,N_5939,N_5140);
nor U8356 (N_8356,N_5333,N_4459);
nor U8357 (N_8357,N_5965,N_5973);
nand U8358 (N_8358,N_4867,N_5152);
xor U8359 (N_8359,N_5398,N_5311);
xor U8360 (N_8360,N_3172,N_3579);
and U8361 (N_8361,N_3525,N_5833);
xor U8362 (N_8362,N_3901,N_5069);
xor U8363 (N_8363,N_5403,N_5747);
nor U8364 (N_8364,N_3326,N_3958);
nor U8365 (N_8365,N_5971,N_4917);
or U8366 (N_8366,N_3764,N_5635);
nand U8367 (N_8367,N_5839,N_3763);
or U8368 (N_8368,N_4940,N_5238);
xnor U8369 (N_8369,N_4230,N_3015);
nand U8370 (N_8370,N_3099,N_5633);
nand U8371 (N_8371,N_4597,N_5788);
nand U8372 (N_8372,N_4467,N_4015);
or U8373 (N_8373,N_5351,N_3453);
or U8374 (N_8374,N_3387,N_5229);
nand U8375 (N_8375,N_4194,N_5608);
or U8376 (N_8376,N_5266,N_5729);
nor U8377 (N_8377,N_4656,N_5630);
and U8378 (N_8378,N_3923,N_4589);
nor U8379 (N_8379,N_4669,N_4590);
nor U8380 (N_8380,N_4509,N_5119);
and U8381 (N_8381,N_5100,N_5089);
or U8382 (N_8382,N_3315,N_5433);
nand U8383 (N_8383,N_3219,N_4133);
nand U8384 (N_8384,N_3151,N_4337);
nand U8385 (N_8385,N_3216,N_3311);
nor U8386 (N_8386,N_5439,N_3609);
nand U8387 (N_8387,N_5114,N_4305);
nor U8388 (N_8388,N_4419,N_4680);
xnor U8389 (N_8389,N_4014,N_5212);
nor U8390 (N_8390,N_3928,N_5665);
nor U8391 (N_8391,N_4940,N_5410);
and U8392 (N_8392,N_3384,N_4071);
or U8393 (N_8393,N_3205,N_4902);
nand U8394 (N_8394,N_5112,N_3429);
xor U8395 (N_8395,N_5786,N_4693);
or U8396 (N_8396,N_3069,N_4633);
and U8397 (N_8397,N_5255,N_3134);
nand U8398 (N_8398,N_5251,N_5520);
or U8399 (N_8399,N_3070,N_5753);
nor U8400 (N_8400,N_5870,N_4910);
nand U8401 (N_8401,N_5253,N_4162);
xor U8402 (N_8402,N_3535,N_3343);
and U8403 (N_8403,N_3097,N_3995);
and U8404 (N_8404,N_4322,N_3447);
or U8405 (N_8405,N_3656,N_4177);
or U8406 (N_8406,N_4760,N_5843);
or U8407 (N_8407,N_4664,N_3410);
nand U8408 (N_8408,N_5124,N_5950);
or U8409 (N_8409,N_4666,N_4917);
or U8410 (N_8410,N_5842,N_5674);
nand U8411 (N_8411,N_4666,N_3772);
or U8412 (N_8412,N_5529,N_4460);
or U8413 (N_8413,N_4477,N_5672);
nor U8414 (N_8414,N_3376,N_5859);
nand U8415 (N_8415,N_4492,N_4852);
and U8416 (N_8416,N_5329,N_3082);
nor U8417 (N_8417,N_5658,N_4390);
and U8418 (N_8418,N_5150,N_4023);
nor U8419 (N_8419,N_5771,N_3955);
xnor U8420 (N_8420,N_3576,N_4694);
or U8421 (N_8421,N_4934,N_3261);
nand U8422 (N_8422,N_3014,N_4470);
xor U8423 (N_8423,N_4376,N_3189);
nor U8424 (N_8424,N_3454,N_4290);
nor U8425 (N_8425,N_4216,N_5834);
nor U8426 (N_8426,N_5388,N_5547);
nor U8427 (N_8427,N_4813,N_4790);
and U8428 (N_8428,N_3125,N_3883);
or U8429 (N_8429,N_5257,N_3418);
nor U8430 (N_8430,N_3221,N_3765);
nand U8431 (N_8431,N_5742,N_4727);
nand U8432 (N_8432,N_3167,N_4880);
and U8433 (N_8433,N_5231,N_5801);
or U8434 (N_8434,N_5688,N_3649);
and U8435 (N_8435,N_4966,N_5578);
nor U8436 (N_8436,N_3664,N_3831);
xor U8437 (N_8437,N_4871,N_4909);
nand U8438 (N_8438,N_3428,N_3523);
nand U8439 (N_8439,N_3232,N_5045);
and U8440 (N_8440,N_4207,N_3212);
xnor U8441 (N_8441,N_5253,N_5954);
and U8442 (N_8442,N_5402,N_4182);
and U8443 (N_8443,N_4126,N_5909);
xor U8444 (N_8444,N_5996,N_4319);
xor U8445 (N_8445,N_4262,N_3753);
and U8446 (N_8446,N_3324,N_5143);
xnor U8447 (N_8447,N_4007,N_3119);
nor U8448 (N_8448,N_4390,N_3641);
nor U8449 (N_8449,N_5641,N_5934);
xnor U8450 (N_8450,N_3105,N_3045);
nor U8451 (N_8451,N_3778,N_4907);
or U8452 (N_8452,N_5389,N_5796);
nand U8453 (N_8453,N_5393,N_5865);
nand U8454 (N_8454,N_3553,N_4125);
or U8455 (N_8455,N_4887,N_5629);
xnor U8456 (N_8456,N_3914,N_3743);
or U8457 (N_8457,N_5599,N_4813);
xor U8458 (N_8458,N_5934,N_4727);
nor U8459 (N_8459,N_5026,N_4881);
or U8460 (N_8460,N_3567,N_4688);
or U8461 (N_8461,N_3972,N_4151);
and U8462 (N_8462,N_4165,N_5618);
and U8463 (N_8463,N_5418,N_4251);
and U8464 (N_8464,N_5752,N_3240);
nand U8465 (N_8465,N_3285,N_3474);
nand U8466 (N_8466,N_5775,N_5874);
nand U8467 (N_8467,N_5647,N_5898);
xnor U8468 (N_8468,N_4121,N_4455);
xor U8469 (N_8469,N_3265,N_3819);
nor U8470 (N_8470,N_3259,N_4628);
nor U8471 (N_8471,N_5664,N_5512);
nand U8472 (N_8472,N_5711,N_4399);
nand U8473 (N_8473,N_5598,N_5186);
nand U8474 (N_8474,N_4120,N_4569);
xor U8475 (N_8475,N_3374,N_3046);
nand U8476 (N_8476,N_5624,N_4354);
and U8477 (N_8477,N_5911,N_4023);
nand U8478 (N_8478,N_3063,N_3700);
and U8479 (N_8479,N_4051,N_4965);
xor U8480 (N_8480,N_3700,N_3070);
nor U8481 (N_8481,N_4638,N_3699);
xor U8482 (N_8482,N_3837,N_3408);
xor U8483 (N_8483,N_5876,N_4111);
or U8484 (N_8484,N_5534,N_3249);
nand U8485 (N_8485,N_5966,N_4620);
and U8486 (N_8486,N_4723,N_4354);
nand U8487 (N_8487,N_3839,N_5661);
and U8488 (N_8488,N_3939,N_4274);
and U8489 (N_8489,N_5972,N_4467);
xor U8490 (N_8490,N_4413,N_5158);
nor U8491 (N_8491,N_5380,N_5080);
nand U8492 (N_8492,N_3390,N_4413);
nor U8493 (N_8493,N_3066,N_3953);
and U8494 (N_8494,N_5966,N_4243);
xor U8495 (N_8495,N_3181,N_4855);
nand U8496 (N_8496,N_3300,N_5589);
or U8497 (N_8497,N_5336,N_5572);
or U8498 (N_8498,N_5783,N_4527);
or U8499 (N_8499,N_4013,N_4673);
xnor U8500 (N_8500,N_4088,N_4472);
nor U8501 (N_8501,N_5297,N_3170);
nor U8502 (N_8502,N_5937,N_5474);
or U8503 (N_8503,N_4117,N_5636);
xor U8504 (N_8504,N_3217,N_5639);
nor U8505 (N_8505,N_5877,N_4010);
xor U8506 (N_8506,N_4396,N_4564);
nand U8507 (N_8507,N_3532,N_5014);
or U8508 (N_8508,N_3150,N_3577);
nor U8509 (N_8509,N_5791,N_5043);
and U8510 (N_8510,N_5521,N_4817);
and U8511 (N_8511,N_3095,N_3532);
nor U8512 (N_8512,N_4121,N_3640);
or U8513 (N_8513,N_3381,N_5417);
xor U8514 (N_8514,N_4067,N_3067);
or U8515 (N_8515,N_5019,N_3545);
or U8516 (N_8516,N_4663,N_5417);
and U8517 (N_8517,N_3682,N_4921);
and U8518 (N_8518,N_3890,N_5572);
nand U8519 (N_8519,N_3051,N_4381);
nor U8520 (N_8520,N_4507,N_5020);
or U8521 (N_8521,N_3465,N_5419);
and U8522 (N_8522,N_4372,N_5631);
nand U8523 (N_8523,N_3871,N_4019);
or U8524 (N_8524,N_4734,N_5634);
and U8525 (N_8525,N_3522,N_5407);
xnor U8526 (N_8526,N_3124,N_3535);
or U8527 (N_8527,N_5848,N_3328);
nor U8528 (N_8528,N_4296,N_5304);
nand U8529 (N_8529,N_4959,N_3459);
and U8530 (N_8530,N_3175,N_5654);
nand U8531 (N_8531,N_3071,N_4395);
xor U8532 (N_8532,N_5600,N_3421);
and U8533 (N_8533,N_4335,N_5752);
nand U8534 (N_8534,N_5716,N_4086);
nor U8535 (N_8535,N_5411,N_3862);
nand U8536 (N_8536,N_5950,N_5670);
nand U8537 (N_8537,N_5866,N_5678);
xnor U8538 (N_8538,N_5142,N_3216);
nand U8539 (N_8539,N_5013,N_4375);
or U8540 (N_8540,N_4283,N_5681);
xnor U8541 (N_8541,N_3617,N_4435);
xnor U8542 (N_8542,N_4397,N_5248);
and U8543 (N_8543,N_4193,N_4194);
nor U8544 (N_8544,N_4665,N_3645);
xor U8545 (N_8545,N_5069,N_4505);
and U8546 (N_8546,N_5092,N_3243);
nand U8547 (N_8547,N_5843,N_4903);
and U8548 (N_8548,N_4010,N_4966);
and U8549 (N_8549,N_4399,N_5401);
and U8550 (N_8550,N_5048,N_4979);
and U8551 (N_8551,N_3704,N_3921);
or U8552 (N_8552,N_5295,N_4525);
xnor U8553 (N_8553,N_4978,N_4449);
nand U8554 (N_8554,N_3839,N_3196);
nor U8555 (N_8555,N_3726,N_5972);
nand U8556 (N_8556,N_5136,N_3082);
and U8557 (N_8557,N_4214,N_3192);
and U8558 (N_8558,N_3376,N_5696);
and U8559 (N_8559,N_4746,N_3223);
or U8560 (N_8560,N_3370,N_4152);
and U8561 (N_8561,N_4155,N_3458);
nor U8562 (N_8562,N_4813,N_5093);
xnor U8563 (N_8563,N_4381,N_4797);
nand U8564 (N_8564,N_5201,N_3603);
nor U8565 (N_8565,N_5982,N_4215);
or U8566 (N_8566,N_5487,N_3490);
and U8567 (N_8567,N_5511,N_4245);
or U8568 (N_8568,N_3726,N_3376);
and U8569 (N_8569,N_3441,N_5289);
nor U8570 (N_8570,N_4144,N_4977);
or U8571 (N_8571,N_4638,N_4152);
and U8572 (N_8572,N_5510,N_5781);
nor U8573 (N_8573,N_3625,N_3930);
nand U8574 (N_8574,N_3749,N_4718);
or U8575 (N_8575,N_5655,N_4707);
nand U8576 (N_8576,N_4636,N_4227);
and U8577 (N_8577,N_5919,N_4244);
nor U8578 (N_8578,N_3210,N_4512);
nand U8579 (N_8579,N_4803,N_3180);
nor U8580 (N_8580,N_4284,N_3634);
xnor U8581 (N_8581,N_3001,N_5570);
xnor U8582 (N_8582,N_5257,N_4636);
or U8583 (N_8583,N_5622,N_3627);
and U8584 (N_8584,N_5300,N_3536);
or U8585 (N_8585,N_4615,N_4765);
nand U8586 (N_8586,N_3716,N_3845);
nand U8587 (N_8587,N_4298,N_4651);
nor U8588 (N_8588,N_5136,N_5761);
and U8589 (N_8589,N_3718,N_4091);
nor U8590 (N_8590,N_4425,N_4765);
nor U8591 (N_8591,N_4451,N_3922);
xnor U8592 (N_8592,N_4348,N_4622);
or U8593 (N_8593,N_3626,N_5159);
nand U8594 (N_8594,N_4139,N_4871);
xnor U8595 (N_8595,N_3534,N_4983);
nand U8596 (N_8596,N_3392,N_5223);
xor U8597 (N_8597,N_5762,N_4459);
nor U8598 (N_8598,N_4979,N_3053);
or U8599 (N_8599,N_4480,N_3281);
nor U8600 (N_8600,N_3082,N_3181);
and U8601 (N_8601,N_5381,N_4077);
and U8602 (N_8602,N_5204,N_4723);
xor U8603 (N_8603,N_4110,N_4593);
and U8604 (N_8604,N_4091,N_4895);
and U8605 (N_8605,N_5663,N_3645);
xor U8606 (N_8606,N_5934,N_3485);
nor U8607 (N_8607,N_4525,N_4277);
and U8608 (N_8608,N_3285,N_4666);
nor U8609 (N_8609,N_4979,N_3745);
or U8610 (N_8610,N_3397,N_4893);
or U8611 (N_8611,N_4691,N_4219);
nor U8612 (N_8612,N_3719,N_3549);
and U8613 (N_8613,N_3262,N_5756);
nand U8614 (N_8614,N_5302,N_4769);
or U8615 (N_8615,N_3334,N_4829);
xor U8616 (N_8616,N_4512,N_5493);
xnor U8617 (N_8617,N_5206,N_4175);
nor U8618 (N_8618,N_5609,N_3153);
nor U8619 (N_8619,N_4872,N_5689);
nor U8620 (N_8620,N_5377,N_3755);
nand U8621 (N_8621,N_3602,N_3017);
xor U8622 (N_8622,N_5680,N_3620);
and U8623 (N_8623,N_4140,N_5175);
and U8624 (N_8624,N_4160,N_5785);
xnor U8625 (N_8625,N_3949,N_5214);
xnor U8626 (N_8626,N_5365,N_5636);
xor U8627 (N_8627,N_3715,N_5199);
or U8628 (N_8628,N_4993,N_4367);
or U8629 (N_8629,N_4425,N_4154);
and U8630 (N_8630,N_5712,N_4156);
nand U8631 (N_8631,N_3380,N_4457);
and U8632 (N_8632,N_3829,N_3008);
nand U8633 (N_8633,N_4626,N_4430);
nor U8634 (N_8634,N_5335,N_5185);
nand U8635 (N_8635,N_5742,N_4730);
xnor U8636 (N_8636,N_5181,N_4012);
nand U8637 (N_8637,N_3687,N_5889);
nor U8638 (N_8638,N_3228,N_4418);
or U8639 (N_8639,N_4667,N_3461);
nand U8640 (N_8640,N_4830,N_4491);
or U8641 (N_8641,N_5402,N_5307);
xor U8642 (N_8642,N_3039,N_4825);
nand U8643 (N_8643,N_5202,N_5325);
nand U8644 (N_8644,N_5072,N_3336);
xnor U8645 (N_8645,N_5600,N_5952);
nand U8646 (N_8646,N_4334,N_5676);
nor U8647 (N_8647,N_5381,N_4441);
nand U8648 (N_8648,N_5258,N_3238);
nand U8649 (N_8649,N_4315,N_3361);
xnor U8650 (N_8650,N_5983,N_5633);
or U8651 (N_8651,N_3041,N_5453);
xor U8652 (N_8652,N_4133,N_3065);
nor U8653 (N_8653,N_5880,N_5020);
or U8654 (N_8654,N_3114,N_5445);
xnor U8655 (N_8655,N_4051,N_4585);
or U8656 (N_8656,N_3253,N_3900);
nor U8657 (N_8657,N_3654,N_4482);
nand U8658 (N_8658,N_4066,N_5312);
nand U8659 (N_8659,N_3814,N_5871);
and U8660 (N_8660,N_4194,N_3790);
xor U8661 (N_8661,N_3567,N_5258);
and U8662 (N_8662,N_3414,N_4145);
nor U8663 (N_8663,N_4816,N_5786);
nor U8664 (N_8664,N_3638,N_5304);
nand U8665 (N_8665,N_3697,N_4375);
and U8666 (N_8666,N_4451,N_4770);
nor U8667 (N_8667,N_3236,N_3463);
and U8668 (N_8668,N_5718,N_5607);
and U8669 (N_8669,N_5582,N_5688);
nand U8670 (N_8670,N_5212,N_3739);
or U8671 (N_8671,N_3574,N_3499);
nor U8672 (N_8672,N_4745,N_4084);
nor U8673 (N_8673,N_3515,N_5017);
xor U8674 (N_8674,N_4181,N_5256);
or U8675 (N_8675,N_5734,N_3377);
or U8676 (N_8676,N_3932,N_3411);
nor U8677 (N_8677,N_4777,N_4754);
nand U8678 (N_8678,N_4090,N_3288);
and U8679 (N_8679,N_4800,N_4553);
xnor U8680 (N_8680,N_5134,N_3701);
nand U8681 (N_8681,N_4678,N_4004);
nand U8682 (N_8682,N_5078,N_5111);
and U8683 (N_8683,N_3442,N_3807);
and U8684 (N_8684,N_4114,N_3298);
nand U8685 (N_8685,N_3664,N_5824);
xor U8686 (N_8686,N_4482,N_3182);
nor U8687 (N_8687,N_3555,N_3409);
nor U8688 (N_8688,N_5256,N_5306);
nand U8689 (N_8689,N_4111,N_4535);
and U8690 (N_8690,N_3124,N_3262);
nand U8691 (N_8691,N_3250,N_4430);
nand U8692 (N_8692,N_4652,N_3542);
nor U8693 (N_8693,N_3413,N_4807);
nand U8694 (N_8694,N_4203,N_5897);
or U8695 (N_8695,N_3681,N_4467);
nor U8696 (N_8696,N_5241,N_5770);
or U8697 (N_8697,N_3470,N_3211);
and U8698 (N_8698,N_4206,N_3506);
nor U8699 (N_8699,N_5720,N_3526);
nand U8700 (N_8700,N_3159,N_5386);
and U8701 (N_8701,N_5531,N_5349);
xor U8702 (N_8702,N_3337,N_3138);
nand U8703 (N_8703,N_3857,N_5169);
nand U8704 (N_8704,N_5389,N_4633);
nand U8705 (N_8705,N_3794,N_4972);
xor U8706 (N_8706,N_4511,N_3231);
nor U8707 (N_8707,N_5546,N_5745);
nor U8708 (N_8708,N_3926,N_3091);
nor U8709 (N_8709,N_3399,N_5045);
and U8710 (N_8710,N_4872,N_3400);
nand U8711 (N_8711,N_3913,N_3478);
nand U8712 (N_8712,N_5745,N_5685);
xor U8713 (N_8713,N_5866,N_3277);
or U8714 (N_8714,N_3908,N_5786);
nor U8715 (N_8715,N_3255,N_5688);
or U8716 (N_8716,N_3538,N_4953);
and U8717 (N_8717,N_4740,N_3957);
and U8718 (N_8718,N_3776,N_5461);
or U8719 (N_8719,N_4695,N_3093);
and U8720 (N_8720,N_5407,N_5463);
and U8721 (N_8721,N_4465,N_3902);
nand U8722 (N_8722,N_3995,N_3399);
xnor U8723 (N_8723,N_3135,N_4192);
nand U8724 (N_8724,N_4647,N_5069);
nand U8725 (N_8725,N_4713,N_3647);
and U8726 (N_8726,N_4189,N_4828);
nor U8727 (N_8727,N_3071,N_3565);
nor U8728 (N_8728,N_3450,N_4813);
xnor U8729 (N_8729,N_4988,N_5975);
xor U8730 (N_8730,N_4800,N_4781);
xnor U8731 (N_8731,N_3722,N_4802);
nand U8732 (N_8732,N_4796,N_4857);
and U8733 (N_8733,N_5538,N_4202);
nor U8734 (N_8734,N_4211,N_5260);
xnor U8735 (N_8735,N_4786,N_4410);
nor U8736 (N_8736,N_5724,N_4947);
and U8737 (N_8737,N_4370,N_3733);
and U8738 (N_8738,N_3390,N_5195);
nand U8739 (N_8739,N_5868,N_4922);
or U8740 (N_8740,N_3014,N_4315);
nor U8741 (N_8741,N_4130,N_3123);
xor U8742 (N_8742,N_3412,N_5752);
and U8743 (N_8743,N_3511,N_3453);
nor U8744 (N_8744,N_3245,N_4805);
and U8745 (N_8745,N_5471,N_5680);
nand U8746 (N_8746,N_3441,N_3484);
and U8747 (N_8747,N_5760,N_3430);
or U8748 (N_8748,N_4907,N_4167);
xnor U8749 (N_8749,N_3772,N_5279);
or U8750 (N_8750,N_4896,N_5862);
or U8751 (N_8751,N_5797,N_5800);
and U8752 (N_8752,N_3281,N_5921);
and U8753 (N_8753,N_5986,N_3517);
or U8754 (N_8754,N_3258,N_3103);
nor U8755 (N_8755,N_5293,N_4117);
or U8756 (N_8756,N_5548,N_5563);
or U8757 (N_8757,N_4545,N_3687);
and U8758 (N_8758,N_5056,N_3091);
nand U8759 (N_8759,N_4706,N_5274);
and U8760 (N_8760,N_3531,N_4329);
nor U8761 (N_8761,N_5817,N_4757);
and U8762 (N_8762,N_3946,N_4515);
xnor U8763 (N_8763,N_3075,N_5166);
nand U8764 (N_8764,N_5490,N_3165);
or U8765 (N_8765,N_5415,N_3688);
and U8766 (N_8766,N_5656,N_3352);
or U8767 (N_8767,N_5970,N_5129);
xnor U8768 (N_8768,N_3405,N_5210);
and U8769 (N_8769,N_4643,N_4498);
and U8770 (N_8770,N_4470,N_5265);
nor U8771 (N_8771,N_5701,N_4142);
nor U8772 (N_8772,N_3689,N_3003);
nand U8773 (N_8773,N_4998,N_5245);
or U8774 (N_8774,N_5468,N_5789);
nand U8775 (N_8775,N_5097,N_3290);
or U8776 (N_8776,N_3451,N_3180);
nand U8777 (N_8777,N_4549,N_3670);
or U8778 (N_8778,N_3021,N_3943);
nand U8779 (N_8779,N_3439,N_3916);
xor U8780 (N_8780,N_5937,N_3626);
and U8781 (N_8781,N_4393,N_4233);
or U8782 (N_8782,N_4623,N_3206);
nand U8783 (N_8783,N_4076,N_3740);
nor U8784 (N_8784,N_3981,N_4786);
xor U8785 (N_8785,N_3122,N_3318);
or U8786 (N_8786,N_4305,N_4859);
and U8787 (N_8787,N_3411,N_4680);
nor U8788 (N_8788,N_5942,N_5006);
nand U8789 (N_8789,N_4119,N_4816);
or U8790 (N_8790,N_3334,N_4310);
or U8791 (N_8791,N_4768,N_5488);
nor U8792 (N_8792,N_5219,N_5853);
and U8793 (N_8793,N_5440,N_3206);
xor U8794 (N_8794,N_5499,N_5809);
xor U8795 (N_8795,N_4929,N_4893);
and U8796 (N_8796,N_4885,N_4189);
nand U8797 (N_8797,N_4727,N_4908);
and U8798 (N_8798,N_3827,N_4041);
or U8799 (N_8799,N_4849,N_4716);
or U8800 (N_8800,N_4743,N_3937);
and U8801 (N_8801,N_4600,N_5167);
xor U8802 (N_8802,N_3403,N_5951);
or U8803 (N_8803,N_3738,N_5690);
or U8804 (N_8804,N_5532,N_4876);
nand U8805 (N_8805,N_5485,N_3658);
or U8806 (N_8806,N_4014,N_4522);
and U8807 (N_8807,N_5460,N_5519);
nand U8808 (N_8808,N_5982,N_3677);
nor U8809 (N_8809,N_3278,N_5810);
nand U8810 (N_8810,N_4326,N_4244);
and U8811 (N_8811,N_4646,N_4742);
or U8812 (N_8812,N_5651,N_3793);
or U8813 (N_8813,N_4061,N_3427);
or U8814 (N_8814,N_5594,N_5892);
xor U8815 (N_8815,N_4803,N_4455);
xnor U8816 (N_8816,N_3864,N_3527);
or U8817 (N_8817,N_5925,N_4744);
nor U8818 (N_8818,N_5171,N_3010);
nor U8819 (N_8819,N_4691,N_3507);
xor U8820 (N_8820,N_3021,N_4544);
or U8821 (N_8821,N_5621,N_3378);
xnor U8822 (N_8822,N_3964,N_5829);
nand U8823 (N_8823,N_4535,N_3866);
and U8824 (N_8824,N_3400,N_5851);
or U8825 (N_8825,N_4967,N_3021);
or U8826 (N_8826,N_4266,N_5197);
and U8827 (N_8827,N_3285,N_4973);
nor U8828 (N_8828,N_5776,N_3290);
or U8829 (N_8829,N_4766,N_4945);
and U8830 (N_8830,N_4675,N_3487);
and U8831 (N_8831,N_3320,N_4625);
or U8832 (N_8832,N_3996,N_4191);
xnor U8833 (N_8833,N_5578,N_4529);
xor U8834 (N_8834,N_4830,N_5002);
nor U8835 (N_8835,N_4762,N_4016);
xor U8836 (N_8836,N_5849,N_4848);
or U8837 (N_8837,N_3417,N_3528);
nor U8838 (N_8838,N_3769,N_5775);
nand U8839 (N_8839,N_5550,N_5324);
or U8840 (N_8840,N_4930,N_3098);
or U8841 (N_8841,N_4238,N_3023);
nor U8842 (N_8842,N_3241,N_4663);
nor U8843 (N_8843,N_5029,N_3472);
nor U8844 (N_8844,N_3389,N_5084);
or U8845 (N_8845,N_5303,N_3825);
and U8846 (N_8846,N_3568,N_4537);
nor U8847 (N_8847,N_5491,N_4955);
nand U8848 (N_8848,N_4965,N_3218);
and U8849 (N_8849,N_4771,N_3149);
or U8850 (N_8850,N_3986,N_5576);
nand U8851 (N_8851,N_4644,N_5260);
nor U8852 (N_8852,N_4460,N_5964);
and U8853 (N_8853,N_4066,N_3336);
and U8854 (N_8854,N_3031,N_4184);
and U8855 (N_8855,N_5524,N_5688);
nand U8856 (N_8856,N_4743,N_4562);
and U8857 (N_8857,N_4831,N_3795);
nor U8858 (N_8858,N_5493,N_5448);
nand U8859 (N_8859,N_5660,N_3832);
and U8860 (N_8860,N_5293,N_3112);
or U8861 (N_8861,N_5504,N_4947);
nand U8862 (N_8862,N_3806,N_4189);
and U8863 (N_8863,N_5397,N_3073);
and U8864 (N_8864,N_4329,N_4388);
nand U8865 (N_8865,N_4934,N_4881);
xnor U8866 (N_8866,N_5667,N_5693);
xnor U8867 (N_8867,N_4159,N_3929);
nand U8868 (N_8868,N_5073,N_5587);
and U8869 (N_8869,N_3015,N_3143);
or U8870 (N_8870,N_4427,N_5799);
and U8871 (N_8871,N_4143,N_3617);
nand U8872 (N_8872,N_5053,N_5407);
xor U8873 (N_8873,N_4147,N_3686);
nor U8874 (N_8874,N_4508,N_5202);
nor U8875 (N_8875,N_3132,N_4025);
nor U8876 (N_8876,N_5013,N_4816);
xor U8877 (N_8877,N_3359,N_3633);
or U8878 (N_8878,N_4439,N_5769);
or U8879 (N_8879,N_3889,N_3905);
or U8880 (N_8880,N_4465,N_5296);
nor U8881 (N_8881,N_5479,N_3547);
nor U8882 (N_8882,N_5688,N_4617);
xor U8883 (N_8883,N_3362,N_5752);
and U8884 (N_8884,N_5727,N_4739);
xor U8885 (N_8885,N_3911,N_5198);
nand U8886 (N_8886,N_4504,N_4805);
nor U8887 (N_8887,N_4673,N_4973);
and U8888 (N_8888,N_4443,N_4845);
nor U8889 (N_8889,N_5680,N_4005);
nand U8890 (N_8890,N_4582,N_5028);
xor U8891 (N_8891,N_4547,N_5259);
nor U8892 (N_8892,N_5607,N_4066);
or U8893 (N_8893,N_5098,N_5341);
or U8894 (N_8894,N_5323,N_4572);
or U8895 (N_8895,N_4742,N_4509);
or U8896 (N_8896,N_4380,N_3297);
or U8897 (N_8897,N_3767,N_5981);
or U8898 (N_8898,N_4944,N_3907);
or U8899 (N_8899,N_5229,N_5933);
or U8900 (N_8900,N_5624,N_3735);
nand U8901 (N_8901,N_4322,N_3645);
nand U8902 (N_8902,N_5631,N_5905);
and U8903 (N_8903,N_5187,N_4983);
and U8904 (N_8904,N_4387,N_4996);
nor U8905 (N_8905,N_3273,N_4863);
and U8906 (N_8906,N_4578,N_5826);
nand U8907 (N_8907,N_4605,N_4831);
xor U8908 (N_8908,N_4028,N_4245);
nand U8909 (N_8909,N_4501,N_4391);
or U8910 (N_8910,N_5973,N_4158);
or U8911 (N_8911,N_3854,N_5522);
nand U8912 (N_8912,N_5710,N_5707);
nand U8913 (N_8913,N_3549,N_4763);
or U8914 (N_8914,N_4368,N_3315);
and U8915 (N_8915,N_3517,N_5691);
or U8916 (N_8916,N_5599,N_5812);
or U8917 (N_8917,N_3042,N_3520);
xnor U8918 (N_8918,N_4388,N_4633);
nor U8919 (N_8919,N_4569,N_5816);
or U8920 (N_8920,N_3797,N_3223);
nor U8921 (N_8921,N_4786,N_3730);
nand U8922 (N_8922,N_4473,N_3509);
nand U8923 (N_8923,N_5820,N_5253);
nand U8924 (N_8924,N_3009,N_5104);
and U8925 (N_8925,N_5031,N_3608);
xor U8926 (N_8926,N_5147,N_5327);
and U8927 (N_8927,N_3928,N_3965);
and U8928 (N_8928,N_3699,N_3495);
nand U8929 (N_8929,N_3894,N_5810);
and U8930 (N_8930,N_3028,N_3370);
nand U8931 (N_8931,N_3894,N_4076);
nor U8932 (N_8932,N_3673,N_5857);
nor U8933 (N_8933,N_5074,N_4324);
nor U8934 (N_8934,N_5392,N_4331);
and U8935 (N_8935,N_4564,N_5932);
nand U8936 (N_8936,N_5316,N_5768);
nand U8937 (N_8937,N_5353,N_4220);
or U8938 (N_8938,N_5449,N_5259);
and U8939 (N_8939,N_4641,N_4851);
and U8940 (N_8940,N_5032,N_4123);
nor U8941 (N_8941,N_4613,N_4530);
and U8942 (N_8942,N_3848,N_4712);
and U8943 (N_8943,N_3019,N_4384);
nor U8944 (N_8944,N_5873,N_4590);
xor U8945 (N_8945,N_4737,N_5643);
or U8946 (N_8946,N_3006,N_5195);
nand U8947 (N_8947,N_5084,N_4346);
xnor U8948 (N_8948,N_4077,N_4252);
or U8949 (N_8949,N_4327,N_4107);
xnor U8950 (N_8950,N_3946,N_5005);
xnor U8951 (N_8951,N_5105,N_3756);
or U8952 (N_8952,N_3332,N_5133);
and U8953 (N_8953,N_5124,N_3539);
xnor U8954 (N_8954,N_5631,N_4688);
xnor U8955 (N_8955,N_4681,N_3314);
nand U8956 (N_8956,N_5654,N_5002);
nor U8957 (N_8957,N_5493,N_3763);
and U8958 (N_8958,N_5539,N_5311);
nor U8959 (N_8959,N_3219,N_4036);
nand U8960 (N_8960,N_3470,N_5631);
xor U8961 (N_8961,N_3517,N_4384);
nor U8962 (N_8962,N_5590,N_4283);
xnor U8963 (N_8963,N_3374,N_3107);
xor U8964 (N_8964,N_4763,N_5972);
nand U8965 (N_8965,N_5014,N_3753);
nor U8966 (N_8966,N_5939,N_4676);
xor U8967 (N_8967,N_3451,N_3814);
and U8968 (N_8968,N_3658,N_5476);
nand U8969 (N_8969,N_4139,N_4759);
or U8970 (N_8970,N_3830,N_5216);
or U8971 (N_8971,N_4335,N_3514);
and U8972 (N_8972,N_5995,N_5031);
nor U8973 (N_8973,N_4452,N_4755);
xor U8974 (N_8974,N_4203,N_5176);
or U8975 (N_8975,N_4001,N_4536);
nand U8976 (N_8976,N_4447,N_4492);
xor U8977 (N_8977,N_4916,N_4847);
nor U8978 (N_8978,N_3743,N_5536);
and U8979 (N_8979,N_5299,N_5256);
or U8980 (N_8980,N_4594,N_3022);
nor U8981 (N_8981,N_4607,N_3715);
and U8982 (N_8982,N_4426,N_4851);
nor U8983 (N_8983,N_3134,N_5295);
nand U8984 (N_8984,N_3779,N_3741);
xnor U8985 (N_8985,N_3147,N_3774);
and U8986 (N_8986,N_3088,N_4359);
or U8987 (N_8987,N_3995,N_5323);
xor U8988 (N_8988,N_3775,N_3363);
nand U8989 (N_8989,N_4617,N_3453);
nand U8990 (N_8990,N_4102,N_3949);
nand U8991 (N_8991,N_4821,N_5498);
and U8992 (N_8992,N_4620,N_4372);
nor U8993 (N_8993,N_4648,N_4163);
and U8994 (N_8994,N_5602,N_5841);
xnor U8995 (N_8995,N_4781,N_5198);
xor U8996 (N_8996,N_5403,N_3856);
nor U8997 (N_8997,N_3996,N_4499);
xor U8998 (N_8998,N_5072,N_3035);
and U8999 (N_8999,N_3228,N_4347);
or U9000 (N_9000,N_7856,N_7839);
nand U9001 (N_9001,N_7690,N_7428);
xnor U9002 (N_9002,N_7957,N_6816);
nand U9003 (N_9003,N_6315,N_6591);
xnor U9004 (N_9004,N_7866,N_6686);
nor U9005 (N_9005,N_8154,N_6020);
or U9006 (N_9006,N_6067,N_7554);
and U9007 (N_9007,N_7951,N_7697);
nor U9008 (N_9008,N_8530,N_7001);
xnor U9009 (N_9009,N_6465,N_6423);
nand U9010 (N_9010,N_7847,N_7923);
or U9011 (N_9011,N_7802,N_6030);
nor U9012 (N_9012,N_8397,N_6204);
or U9013 (N_9013,N_7787,N_8691);
and U9014 (N_9014,N_6333,N_7713);
nand U9015 (N_9015,N_6434,N_8762);
xnor U9016 (N_9016,N_7340,N_6502);
nand U9017 (N_9017,N_8953,N_7973);
nor U9018 (N_9018,N_8703,N_7635);
nor U9019 (N_9019,N_6092,N_7005);
or U9020 (N_9020,N_8045,N_8727);
nor U9021 (N_9021,N_7263,N_8574);
and U9022 (N_9022,N_6191,N_8428);
and U9023 (N_9023,N_8495,N_8377);
xor U9024 (N_9024,N_8635,N_6342);
or U9025 (N_9025,N_8618,N_7834);
or U9026 (N_9026,N_7492,N_8331);
xor U9027 (N_9027,N_8255,N_7541);
nand U9028 (N_9028,N_6751,N_6582);
nand U9029 (N_9029,N_8003,N_7682);
nand U9030 (N_9030,N_8219,N_6226);
and U9031 (N_9031,N_6606,N_7711);
and U9032 (N_9032,N_7507,N_6113);
or U9033 (N_9033,N_6167,N_6171);
nor U9034 (N_9034,N_6773,N_6593);
or U9035 (N_9035,N_7646,N_6600);
xnor U9036 (N_9036,N_7396,N_8900);
and U9037 (N_9037,N_7833,N_6868);
or U9038 (N_9038,N_8764,N_7377);
or U9039 (N_9039,N_8141,N_6481);
and U9040 (N_9040,N_6199,N_7485);
and U9041 (N_9041,N_6185,N_6636);
and U9042 (N_9042,N_6879,N_8493);
xnor U9043 (N_9043,N_7247,N_7110);
xnor U9044 (N_9044,N_7088,N_8018);
or U9045 (N_9045,N_7175,N_6206);
nand U9046 (N_9046,N_8786,N_6234);
or U9047 (N_9047,N_8015,N_7859);
and U9048 (N_9048,N_7550,N_6224);
and U9049 (N_9049,N_7022,N_7292);
nand U9050 (N_9050,N_8292,N_6190);
nor U9051 (N_9051,N_6564,N_6466);
or U9052 (N_9052,N_8956,N_7035);
or U9053 (N_9053,N_6691,N_6344);
or U9054 (N_9054,N_8127,N_7013);
nand U9055 (N_9055,N_8627,N_6918);
xnor U9056 (N_9056,N_6876,N_6601);
and U9057 (N_9057,N_6986,N_7685);
or U9058 (N_9058,N_7388,N_6425);
or U9059 (N_9059,N_8676,N_7553);
xnor U9060 (N_9060,N_7749,N_7286);
and U9061 (N_9061,N_8481,N_7364);
or U9062 (N_9062,N_6827,N_7478);
nand U9063 (N_9063,N_6880,N_7440);
nand U9064 (N_9064,N_7234,N_7501);
and U9065 (N_9065,N_6468,N_8624);
xor U9066 (N_9066,N_6676,N_7895);
xnor U9067 (N_9067,N_8091,N_6475);
nand U9068 (N_9068,N_6808,N_8130);
or U9069 (N_9069,N_7048,N_6872);
nor U9070 (N_9070,N_8022,N_8920);
or U9071 (N_9071,N_6367,N_8487);
nor U9072 (N_9072,N_7722,N_6631);
xnor U9073 (N_9073,N_7611,N_7066);
xnor U9074 (N_9074,N_6650,N_6172);
nand U9075 (N_9075,N_6145,N_7824);
or U9076 (N_9076,N_7223,N_8419);
nand U9077 (N_9077,N_7023,N_8573);
xor U9078 (N_9078,N_7097,N_6705);
nor U9079 (N_9079,N_6835,N_7257);
nand U9080 (N_9080,N_8374,N_6613);
xnor U9081 (N_9081,N_8284,N_8478);
or U9082 (N_9082,N_6850,N_6871);
nor U9083 (N_9083,N_8551,N_6043);
xor U9084 (N_9084,N_7952,N_7532);
nand U9085 (N_9085,N_8083,N_8375);
nor U9086 (N_9086,N_6073,N_7886);
nor U9087 (N_9087,N_6942,N_8979);
xor U9088 (N_9088,N_6058,N_7304);
nand U9089 (N_9089,N_7917,N_7433);
nor U9090 (N_9090,N_6543,N_8500);
xnor U9091 (N_9091,N_7903,N_6565);
xnor U9092 (N_9092,N_8547,N_8895);
xnor U9093 (N_9093,N_7766,N_7430);
and U9094 (N_9094,N_8062,N_8224);
xnor U9095 (N_9095,N_6015,N_7876);
and U9096 (N_9096,N_7363,N_8776);
nand U9097 (N_9097,N_7865,N_7931);
or U9098 (N_9098,N_7870,N_6744);
xor U9099 (N_9099,N_8008,N_7042);
xnor U9100 (N_9100,N_7046,N_7618);
or U9101 (N_9101,N_6122,N_8823);
nor U9102 (N_9102,N_7450,N_7318);
nor U9103 (N_9103,N_8090,N_6347);
nor U9104 (N_9104,N_8166,N_7301);
nor U9105 (N_9105,N_8978,N_7344);
xnor U9106 (N_9106,N_7813,N_7379);
nand U9107 (N_9107,N_7965,N_6080);
and U9108 (N_9108,N_7881,N_8741);
or U9109 (N_9109,N_7493,N_6138);
and U9110 (N_9110,N_8537,N_8151);
and U9111 (N_9111,N_7176,N_6904);
nand U9112 (N_9112,N_7626,N_6895);
xor U9113 (N_9113,N_6027,N_6694);
and U9114 (N_9114,N_8153,N_7087);
nand U9115 (N_9115,N_6970,N_8519);
nand U9116 (N_9116,N_8173,N_7103);
and U9117 (N_9117,N_6523,N_7768);
or U9118 (N_9118,N_6651,N_8039);
and U9119 (N_9119,N_8633,N_8730);
or U9120 (N_9120,N_7648,N_8840);
nand U9121 (N_9121,N_6075,N_8156);
nand U9122 (N_9122,N_7303,N_8801);
nand U9123 (N_9123,N_7845,N_8886);
xor U9124 (N_9124,N_8448,N_7309);
and U9125 (N_9125,N_7921,N_8854);
and U9126 (N_9126,N_7323,N_6007);
nand U9127 (N_9127,N_8975,N_8929);
nand U9128 (N_9128,N_8174,N_8833);
and U9129 (N_9129,N_7556,N_7663);
nand U9130 (N_9130,N_7276,N_7267);
or U9131 (N_9131,N_6897,N_7579);
nand U9132 (N_9132,N_6361,N_8079);
nor U9133 (N_9133,N_6304,N_7704);
nand U9134 (N_9134,N_8287,N_8928);
nor U9135 (N_9135,N_6718,N_6503);
nand U9136 (N_9136,N_6045,N_6737);
or U9137 (N_9137,N_6758,N_7255);
nor U9138 (N_9138,N_6196,N_7157);
nor U9139 (N_9139,N_6499,N_6783);
and U9140 (N_9140,N_7819,N_7893);
nand U9141 (N_9141,N_8588,N_7037);
and U9142 (N_9142,N_6979,N_6252);
and U9143 (N_9143,N_6143,N_8451);
nor U9144 (N_9144,N_7278,N_7185);
nor U9145 (N_9145,N_8390,N_6464);
nand U9146 (N_9146,N_8641,N_8334);
nand U9147 (N_9147,N_8602,N_8693);
and U9148 (N_9148,N_6653,N_8414);
or U9149 (N_9149,N_7021,N_8778);
nand U9150 (N_9150,N_6507,N_8494);
nand U9151 (N_9151,N_8791,N_7708);
nor U9152 (N_9152,N_6921,N_8328);
nand U9153 (N_9153,N_7641,N_8903);
nor U9154 (N_9154,N_6585,N_6800);
nor U9155 (N_9155,N_7566,N_7788);
xor U9156 (N_9156,N_8545,N_7140);
nor U9157 (N_9157,N_6748,N_7622);
and U9158 (N_9158,N_7426,N_6662);
or U9159 (N_9159,N_6767,N_6928);
xnor U9160 (N_9160,N_8252,N_6449);
and U9161 (N_9161,N_8430,N_6011);
nor U9162 (N_9162,N_6525,N_8695);
nor U9163 (N_9163,N_8209,N_7745);
nand U9164 (N_9164,N_6671,N_6726);
and U9165 (N_9165,N_7806,N_7130);
or U9166 (N_9166,N_6697,N_8059);
xnor U9167 (N_9167,N_8054,N_7068);
and U9168 (N_9168,N_8068,N_6262);
and U9169 (N_9169,N_6055,N_8866);
and U9170 (N_9170,N_7112,N_7432);
or U9171 (N_9171,N_6513,N_7131);
and U9172 (N_9172,N_6088,N_7366);
xnor U9173 (N_9173,N_8132,N_7996);
xor U9174 (N_9174,N_6109,N_7974);
nand U9175 (N_9175,N_6340,N_8733);
and U9176 (N_9176,N_6780,N_8459);
xor U9177 (N_9177,N_8055,N_8101);
xnor U9178 (N_9178,N_6991,N_8014);
nand U9179 (N_9179,N_7853,N_8009);
and U9180 (N_9180,N_8491,N_7864);
nor U9181 (N_9181,N_8612,N_6424);
nand U9182 (N_9182,N_8615,N_6687);
nand U9183 (N_9183,N_6642,N_6992);
nand U9184 (N_9184,N_8197,N_7762);
or U9185 (N_9185,N_8653,N_6711);
xnor U9186 (N_9186,N_8657,N_8844);
xor U9187 (N_9187,N_6188,N_6064);
xor U9188 (N_9188,N_6978,N_7907);
nand U9189 (N_9189,N_7533,N_6397);
xnor U9190 (N_9190,N_6715,N_8282);
and U9191 (N_9191,N_6965,N_7683);
or U9192 (N_9192,N_8097,N_7198);
nand U9193 (N_9193,N_8885,N_6273);
nor U9194 (N_9194,N_8926,N_8195);
xnor U9195 (N_9195,N_8152,N_6387);
nor U9196 (N_9196,N_7457,N_7446);
or U9197 (N_9197,N_8623,N_7522);
and U9198 (N_9198,N_8095,N_8011);
nor U9199 (N_9199,N_8598,N_6455);
or U9200 (N_9200,N_8000,N_6032);
nor U9201 (N_9201,N_7291,N_6328);
nand U9202 (N_9202,N_8146,N_8276);
nand U9203 (N_9203,N_6858,N_8590);
nor U9204 (N_9204,N_8768,N_7427);
and U9205 (N_9205,N_8632,N_7577);
or U9206 (N_9206,N_8348,N_7030);
or U9207 (N_9207,N_7144,N_6669);
and U9208 (N_9208,N_7837,N_8852);
or U9209 (N_9209,N_8382,N_8061);
and U9210 (N_9210,N_6542,N_8483);
or U9211 (N_9211,N_7961,N_7410);
nor U9212 (N_9212,N_8629,N_8706);
and U9213 (N_9213,N_6268,N_6104);
and U9214 (N_9214,N_8820,N_6442);
or U9215 (N_9215,N_8444,N_6903);
nor U9216 (N_9216,N_8467,N_7898);
and U9217 (N_9217,N_6799,N_6739);
and U9218 (N_9218,N_8666,N_7193);
or U9219 (N_9219,N_6278,N_6009);
xor U9220 (N_9220,N_6153,N_7225);
nand U9221 (N_9221,N_6418,N_6017);
xor U9222 (N_9222,N_6555,N_6364);
nand U9223 (N_9223,N_7380,N_7435);
nor U9224 (N_9224,N_8177,N_6626);
or U9225 (N_9225,N_7095,N_8119);
nand U9226 (N_9226,N_8933,N_6356);
xor U9227 (N_9227,N_8476,N_6812);
xor U9228 (N_9228,N_7238,N_8589);
and U9229 (N_9229,N_6628,N_6137);
or U9230 (N_9230,N_6862,N_6955);
xor U9231 (N_9231,N_7592,N_6474);
and U9232 (N_9232,N_6777,N_8032);
and U9233 (N_9233,N_6989,N_7997);
xor U9234 (N_9234,N_6205,N_6453);
xnor U9235 (N_9235,N_6702,N_8980);
or U9236 (N_9236,N_8231,N_6237);
nand U9237 (N_9237,N_8725,N_6335);
and U9238 (N_9238,N_6139,N_8535);
nand U9239 (N_9239,N_7591,N_7976);
and U9240 (N_9240,N_7424,N_6522);
or U9241 (N_9241,N_8363,N_8115);
nand U9242 (N_9242,N_7699,N_6864);
xnor U9243 (N_9243,N_6443,N_7456);
or U9244 (N_9244,N_7496,N_6240);
xnor U9245 (N_9245,N_6810,N_7521);
nand U9246 (N_9246,N_7063,N_6209);
and U9247 (N_9247,N_6791,N_6225);
and U9248 (N_9248,N_8549,N_8966);
nor U9249 (N_9249,N_6785,N_6487);
xnor U9250 (N_9250,N_8896,N_7906);
nand U9251 (N_9251,N_8202,N_7986);
or U9252 (N_9252,N_8527,N_8668);
nor U9253 (N_9253,N_6458,N_7673);
nand U9254 (N_9254,N_8138,N_6359);
or U9255 (N_9255,N_8290,N_8437);
xnor U9256 (N_9256,N_7347,N_8396);
and U9257 (N_9257,N_8184,N_7777);
xnor U9258 (N_9258,N_7888,N_7154);
xor U9259 (N_9259,N_8626,N_7720);
and U9260 (N_9260,N_6415,N_6648);
xor U9261 (N_9261,N_6736,N_7273);
nor U9262 (N_9262,N_7733,N_6042);
nor U9263 (N_9263,N_7992,N_8826);
xnor U9264 (N_9264,N_7275,N_6127);
nor U9265 (N_9265,N_8771,N_6231);
nand U9266 (N_9266,N_8423,N_7786);
and U9267 (N_9267,N_8557,N_7718);
and U9268 (N_9268,N_8908,N_7111);
and U9269 (N_9269,N_7395,N_7100);
or U9270 (N_9270,N_8824,N_8572);
nor U9271 (N_9271,N_6692,N_6269);
nor U9272 (N_9272,N_6065,N_8073);
and U9273 (N_9273,N_6511,N_7387);
xnor U9274 (N_9274,N_8690,N_7354);
and U9275 (N_9275,N_8973,N_7561);
and U9276 (N_9276,N_8313,N_7989);
xnor U9277 (N_9277,N_6257,N_7190);
nor U9278 (N_9278,N_8389,N_7171);
nand U9279 (N_9279,N_6118,N_7345);
nor U9280 (N_9280,N_6771,N_7638);
nand U9281 (N_9281,N_8378,N_6454);
nor U9282 (N_9282,N_7288,N_7857);
nor U9283 (N_9283,N_8967,N_8385);
xnor U9284 (N_9284,N_6912,N_7196);
xnor U9285 (N_9285,N_6002,N_6050);
nand U9286 (N_9286,N_6625,N_8575);
xnor U9287 (N_9287,N_7772,N_7164);
xor U9288 (N_9288,N_6324,N_7880);
nor U9289 (N_9289,N_7399,N_8244);
and U9290 (N_9290,N_7464,N_8497);
or U9291 (N_9291,N_6312,N_7631);
nand U9292 (N_9292,N_7400,N_7576);
or U9293 (N_9293,N_7734,N_6663);
xor U9294 (N_9294,N_6132,N_6515);
and U9295 (N_9295,N_8314,N_7513);
or U9296 (N_9296,N_6670,N_8964);
nor U9297 (N_9297,N_7873,N_6099);
nor U9298 (N_9298,N_7723,N_8888);
nand U9299 (N_9299,N_8064,N_8944);
nand U9300 (N_9300,N_6878,N_6162);
xor U9301 (N_9301,N_8458,N_6557);
and U9302 (N_9302,N_6158,N_8354);
nor U9303 (N_9303,N_6301,N_7069);
nor U9304 (N_9304,N_7589,N_7072);
and U9305 (N_9305,N_7445,N_8369);
nand U9306 (N_9306,N_7544,N_6016);
and U9307 (N_9307,N_6980,N_8664);
and U9308 (N_9308,N_7167,N_7927);
and U9309 (N_9309,N_8832,N_6313);
nor U9310 (N_9310,N_6570,N_8634);
nand U9311 (N_9311,N_7114,N_6260);
or U9312 (N_9312,N_8991,N_8404);
nor U9313 (N_9313,N_7872,N_8552);
or U9314 (N_9314,N_6426,N_6953);
or U9315 (N_9315,N_8279,N_7245);
and U9316 (N_9316,N_7536,N_6221);
nand U9317 (N_9317,N_8422,N_8889);
xnor U9318 (N_9318,N_6552,N_6111);
or U9319 (N_9319,N_7331,N_7517);
and U9320 (N_9320,N_6629,N_8431);
nor U9321 (N_9321,N_6594,N_6411);
or U9322 (N_9322,N_6000,N_8591);
or U9323 (N_9323,N_7148,N_6738);
or U9324 (N_9324,N_6633,N_7503);
nand U9325 (N_9325,N_8140,N_6379);
nand U9326 (N_9326,N_7179,N_7601);
or U9327 (N_9327,N_8894,N_6500);
nor U9328 (N_9328,N_6828,N_7629);
xnor U9329 (N_9329,N_6235,N_8230);
nand U9330 (N_9330,N_7346,N_7914);
and U9331 (N_9331,N_6866,N_6971);
xnor U9332 (N_9332,N_6077,N_7919);
nor U9333 (N_9333,N_6721,N_6517);
nand U9334 (N_9334,N_7827,N_7143);
or U9335 (N_9335,N_7706,N_6709);
nor U9336 (N_9336,N_7365,N_6968);
xnor U9337 (N_9337,N_6433,N_7102);
or U9338 (N_9338,N_7260,N_6504);
xnor U9339 (N_9339,N_7531,N_7017);
xnor U9340 (N_9340,N_8904,N_6090);
and U9341 (N_9341,N_8857,N_8781);
xor U9342 (N_9342,N_7836,N_7341);
or U9343 (N_9343,N_6100,N_8344);
and U9344 (N_9344,N_6657,N_6762);
xor U9345 (N_9345,N_7644,N_6383);
nand U9346 (N_9346,N_7221,N_6526);
and U9347 (N_9347,N_8872,N_8723);
and U9348 (N_9348,N_7324,N_7352);
or U9349 (N_9349,N_6887,N_7737);
xnor U9350 (N_9350,N_8912,N_8106);
xor U9351 (N_9351,N_6822,N_6553);
nand U9352 (N_9352,N_7280,N_8718);
nand U9353 (N_9353,N_8319,N_8324);
nand U9354 (N_9354,N_8553,N_8793);
nor U9355 (N_9355,N_6031,N_7594);
or U9356 (N_9356,N_8168,N_7476);
or U9357 (N_9357,N_6976,N_8020);
xnor U9358 (N_9358,N_8372,N_7082);
and U9359 (N_9359,N_8858,N_7712);
nand U9360 (N_9360,N_8272,N_6796);
or U9361 (N_9361,N_8098,N_7142);
nor U9362 (N_9362,N_6619,N_8205);
xnor U9363 (N_9363,N_6326,N_8782);
and U9364 (N_9364,N_7538,N_7816);
or U9365 (N_9365,N_6298,N_7943);
xnor U9366 (N_9366,N_7851,N_7359);
and U9367 (N_9367,N_8651,N_7200);
xor U9368 (N_9368,N_6168,N_6070);
nor U9369 (N_9369,N_7739,N_6919);
and U9370 (N_9370,N_6062,N_7617);
xnor U9371 (N_9371,N_8248,N_8931);
or U9372 (N_9372,N_7272,N_6926);
nor U9373 (N_9373,N_7606,N_6322);
xnor U9374 (N_9374,N_7401,N_6414);
xnor U9375 (N_9375,N_7206,N_7560);
or U9376 (N_9376,N_7707,N_6284);
nor U9377 (N_9377,N_7133,N_6392);
and U9378 (N_9378,N_7823,N_7939);
or U9379 (N_9379,N_6314,N_6643);
or U9380 (N_9380,N_7877,N_6134);
or U9381 (N_9381,N_8442,N_8253);
or U9382 (N_9382,N_6166,N_8439);
and U9383 (N_9383,N_6461,N_7728);
and U9384 (N_9384,N_6181,N_7709);
and U9385 (N_9385,N_8142,N_7242);
nor U9386 (N_9386,N_6130,N_7466);
or U9387 (N_9387,N_7209,N_6469);
or U9388 (N_9388,N_7306,N_7858);
xnor U9389 (N_9389,N_8460,N_8189);
nand U9390 (N_9390,N_6374,N_7826);
nand U9391 (N_9391,N_7960,N_6627);
and U9392 (N_9392,N_7376,N_7894);
and U9393 (N_9393,N_6365,N_8835);
xor U9394 (N_9394,N_8673,N_6877);
or U9395 (N_9395,N_8760,N_8601);
and U9396 (N_9396,N_8679,N_8688);
or U9397 (N_9397,N_8913,N_8465);
nor U9398 (N_9398,N_7458,N_7878);
or U9399 (N_9399,N_6659,N_6700);
and U9400 (N_9400,N_8479,N_7925);
nor U9401 (N_9401,N_6982,N_8941);
nand U9402 (N_9402,N_8120,N_8084);
and U9403 (N_9403,N_8171,N_8860);
or U9404 (N_9404,N_7724,N_7451);
nor U9405 (N_9405,N_6894,N_8906);
and U9406 (N_9406,N_7564,N_7192);
or U9407 (N_9407,N_7049,N_6655);
nor U9408 (N_9408,N_8897,N_7669);
xor U9409 (N_9409,N_6925,N_6041);
nand U9410 (N_9410,N_7372,N_6784);
nand U9411 (N_9411,N_7811,N_8383);
or U9412 (N_9412,N_7163,N_7809);
and U9413 (N_9413,N_8147,N_6837);
and U9414 (N_9414,N_8016,N_6490);
and U9415 (N_9415,N_6095,N_8600);
xnor U9416 (N_9416,N_6867,N_6615);
nor U9417 (N_9417,N_6961,N_7414);
and U9418 (N_9418,N_7980,N_8105);
nand U9419 (N_9419,N_6439,N_8874);
or U9420 (N_9420,N_7639,N_7295);
nor U9421 (N_9421,N_6714,N_7890);
xnor U9422 (N_9422,N_6610,N_7310);
or U9423 (N_9423,N_6579,N_8568);
xnor U9424 (N_9424,N_6561,N_8167);
or U9425 (N_9425,N_6178,N_7123);
xnor U9426 (N_9426,N_7094,N_7357);
or U9427 (N_9427,N_6775,N_7080);
and U9428 (N_9428,N_6875,N_8243);
or U9429 (N_9429,N_8110,N_8997);
or U9430 (N_9430,N_7854,N_7239);
or U9431 (N_9431,N_8124,N_8373);
nand U9432 (N_9432,N_8092,N_8655);
nor U9433 (N_9433,N_6819,N_6580);
or U9434 (N_9434,N_7370,N_7573);
or U9435 (N_9435,N_6200,N_7012);
nor U9436 (N_9436,N_7759,N_8560);
xnor U9437 (N_9437,N_6456,N_8939);
xnor U9438 (N_9438,N_7381,N_8339);
nand U9439 (N_9439,N_7738,N_6958);
and U9440 (N_9440,N_7735,N_7028);
xor U9441 (N_9441,N_6232,N_8299);
nand U9442 (N_9442,N_6477,N_7882);
or U9443 (N_9443,N_6352,N_7804);
xnor U9444 (N_9444,N_6985,N_7071);
or U9445 (N_9445,N_6803,N_6369);
nand U9446 (N_9446,N_7570,N_6505);
xnor U9447 (N_9447,N_6512,N_7236);
and U9448 (N_9448,N_6381,N_8402);
nand U9449 (N_9449,N_8914,N_8058);
xor U9450 (N_9450,N_7009,N_7180);
or U9451 (N_9451,N_6734,N_6267);
xnor U9452 (N_9452,N_7096,N_8204);
nand U9453 (N_9453,N_7948,N_8183);
xnor U9454 (N_9454,N_7373,N_7434);
xnor U9455 (N_9455,N_8780,N_8454);
nand U9456 (N_9456,N_8955,N_6366);
nor U9457 (N_9457,N_7632,N_7855);
nor U9458 (N_9458,N_8995,N_8795);
xnor U9459 (N_9459,N_8395,N_6782);
or U9460 (N_9460,N_6214,N_7059);
or U9461 (N_9461,N_6963,N_8546);
nand U9462 (N_9462,N_7835,N_8300);
xnor U9463 (N_9463,N_8845,N_7256);
xor U9464 (N_9464,N_6938,N_6845);
nand U9465 (N_9465,N_7916,N_7398);
xor U9466 (N_9466,N_8265,N_7060);
or U9467 (N_9467,N_8355,N_6789);
or U9468 (N_9468,N_7983,N_8471);
nand U9469 (N_9469,N_7885,N_7731);
xor U9470 (N_9470,N_7934,N_7355);
and U9471 (N_9471,N_6436,N_8511);
nor U9472 (N_9472,N_7993,N_6853);
xor U9473 (N_9473,N_8747,N_8398);
nand U9474 (N_9474,N_7829,N_6576);
or U9475 (N_9475,N_6219,N_8685);
or U9476 (N_9476,N_8994,N_6899);
or U9477 (N_9477,N_6933,N_7329);
or U9478 (N_9478,N_8880,N_6757);
or U9479 (N_9479,N_8522,N_8486);
xnor U9480 (N_9480,N_7208,N_8697);
xor U9481 (N_9481,N_8357,N_8320);
nor U9482 (N_9482,N_6173,N_7808);
and U9483 (N_9483,N_6222,N_7092);
nand U9484 (N_9484,N_7681,N_7266);
nor U9485 (N_9485,N_8485,N_7901);
xor U9486 (N_9486,N_6759,N_8607);
and U9487 (N_9487,N_7844,N_8686);
xor U9488 (N_9488,N_8133,N_7313);
nor U9489 (N_9489,N_6203,N_8744);
nor U9490 (N_9490,N_6620,N_6578);
nand U9491 (N_9491,N_7867,N_6612);
nand U9492 (N_9492,N_6212,N_6447);
and U9493 (N_9493,N_7757,N_6401);
and U9494 (N_9494,N_8859,N_8785);
and U9495 (N_9495,N_7812,N_6688);
and U9496 (N_9496,N_6975,N_6901);
xor U9497 (N_9497,N_7480,N_8558);
xor U9498 (N_9498,N_7231,N_8427);
and U9499 (N_9499,N_7019,N_7403);
or U9500 (N_9500,N_6572,N_7038);
nor U9501 (N_9501,N_6695,N_6107);
and U9502 (N_9502,N_6331,N_6683);
nor U9503 (N_9503,N_8873,N_7086);
or U9504 (N_9504,N_6054,N_7074);
xnor U9505 (N_9505,N_8989,N_7004);
nand U9506 (N_9506,N_6696,N_8802);
nor U9507 (N_9507,N_7525,N_6717);
nor U9508 (N_9508,N_7540,N_6851);
nor U9509 (N_9509,N_8525,N_8915);
nand U9510 (N_9510,N_8950,N_8724);
and U9511 (N_9511,N_8490,N_8069);
nand U9512 (N_9512,N_7688,N_8108);
nor U9513 (N_9513,N_6623,N_7694);
or U9514 (N_9514,N_7375,N_8176);
nor U9515 (N_9515,N_8644,N_6826);
and U9516 (N_9516,N_8192,N_6972);
nand U9517 (N_9517,N_6531,N_6797);
and U9518 (N_9518,N_6760,N_8254);
and U9519 (N_9519,N_7431,N_6962);
nor U9520 (N_9520,N_8608,N_7698);
and U9521 (N_9521,N_7454,N_8751);
or U9522 (N_9522,N_6622,N_7298);
nand U9523 (N_9523,N_7563,N_6472);
nand U9524 (N_9524,N_6892,N_7990);
nand U9525 (N_9525,N_7505,N_8850);
or U9526 (N_9526,N_6292,N_6201);
or U9527 (N_9527,N_7582,N_6544);
nand U9528 (N_9528,N_8433,N_8298);
nor U9529 (N_9529,N_7293,N_7546);
and U9530 (N_9530,N_8839,N_8529);
and U9531 (N_9531,N_8214,N_7169);
nor U9532 (N_9532,N_7653,N_8512);
xnor U9533 (N_9533,N_8709,N_7797);
nand U9534 (N_9534,N_6951,N_6459);
xor U9535 (N_9535,N_8816,N_6927);
or U9536 (N_9536,N_8466,N_6289);
xnor U9537 (N_9537,N_8893,N_7002);
nor U9538 (N_9538,N_7453,N_6479);
or U9539 (N_9539,N_6860,N_7442);
nor U9540 (N_9540,N_8707,N_8501);
nor U9541 (N_9541,N_8238,N_6699);
and U9542 (N_9542,N_8463,N_6993);
and U9543 (N_9543,N_6730,N_8837);
and U9544 (N_9544,N_7572,N_6940);
nand U9545 (N_9545,N_6830,N_8998);
xnor U9546 (N_9546,N_6108,N_7736);
nor U9547 (N_9547,N_7268,N_8712);
and U9548 (N_9548,N_8242,N_8620);
nand U9549 (N_9549,N_8853,N_6605);
and U9550 (N_9550,N_8232,N_7774);
and U9551 (N_9551,N_8905,N_7029);
nor U9552 (N_9552,N_6501,N_8870);
xnor U9553 (N_9553,N_8452,N_8808);
nand U9554 (N_9554,N_8200,N_6995);
nand U9555 (N_9555,N_7258,N_8364);
or U9556 (N_9556,N_6838,N_6834);
and U9557 (N_9557,N_8401,N_6338);
nand U9558 (N_9558,N_8756,N_6150);
nand U9559 (N_9559,N_7748,N_7506);
and U9560 (N_9560,N_6913,N_6563);
nor U9561 (N_9561,N_8281,N_7008);
xnor U9562 (N_9562,N_8213,N_6774);
nor U9563 (N_9563,N_8477,N_6920);
nand U9564 (N_9564,N_7312,N_8155);
nor U9565 (N_9565,N_7991,N_7620);
or U9566 (N_9566,N_8233,N_7184);
nor U9567 (N_9567,N_7944,N_6341);
xor U9568 (N_9568,N_6362,N_6484);
and U9569 (N_9569,N_6489,N_6568);
and U9570 (N_9570,N_7207,N_8416);
or U9571 (N_9571,N_8273,N_8569);
and U9572 (N_9572,N_6457,N_6567);
nor U9573 (N_9573,N_6840,N_7640);
xor U9574 (N_9574,N_6616,N_8125);
xnor U9575 (N_9575,N_8502,N_7228);
or U9576 (N_9576,N_7186,N_8052);
and U9577 (N_9577,N_6677,N_7448);
and U9578 (N_9578,N_7122,N_8473);
and U9579 (N_9579,N_8783,N_6528);
xnor U9580 (N_9580,N_8732,N_6410);
nor U9581 (N_9581,N_7443,N_7789);
and U9582 (N_9582,N_6176,N_8267);
nand U9583 (N_9583,N_8643,N_8221);
nor U9584 (N_9584,N_6184,N_6794);
nor U9585 (N_9585,N_8484,N_6779);
xor U9586 (N_9586,N_7539,N_7840);
and U9587 (N_9587,N_8654,N_6417);
or U9588 (N_9588,N_8687,N_8028);
and U9589 (N_9589,N_8236,N_8207);
or U9590 (N_9590,N_7999,N_6242);
or U9591 (N_9591,N_8963,N_8985);
nand U9592 (N_9592,N_7597,N_8322);
or U9593 (N_9593,N_8285,N_6019);
or U9594 (N_9594,N_7281,N_8367);
and U9595 (N_9595,N_8611,N_8102);
xor U9596 (N_9596,N_6355,N_8631);
nand U9597 (N_9597,N_7756,N_6083);
nor U9598 (N_9598,N_6710,N_8086);
nor U9599 (N_9599,N_6558,N_6536);
and U9600 (N_9600,N_6101,N_7106);
or U9601 (N_9601,N_7710,N_7165);
or U9602 (N_9602,N_7821,N_8761);
nand U9603 (N_9603,N_6516,N_6882);
and U9604 (N_9604,N_8610,N_6022);
or U9605 (N_9605,N_8800,N_6082);
xor U9606 (N_9606,N_8114,N_6087);
nor U9607 (N_9607,N_6679,N_7499);
and U9608 (N_9608,N_7526,N_8379);
or U9609 (N_9609,N_6157,N_8464);
nand U9610 (N_9610,N_8260,N_6427);
and U9611 (N_9611,N_7025,N_8675);
xor U9612 (N_9612,N_8834,N_7213);
xnor U9613 (N_9613,N_7040,N_8050);
nand U9614 (N_9614,N_8033,N_6805);
or U9615 (N_9615,N_6518,N_7128);
and U9616 (N_9616,N_6916,N_8038);
or U9617 (N_9617,N_7385,N_7585);
or U9618 (N_9618,N_8739,N_6350);
xnor U9619 (N_9619,N_6251,N_8619);
xor U9620 (N_9620,N_6949,N_6317);
nor U9621 (N_9621,N_7216,N_8936);
and U9622 (N_9622,N_8294,N_7803);
xor U9623 (N_9623,N_6519,N_8954);
and U9624 (N_9624,N_8093,N_7394);
or U9625 (N_9625,N_8291,N_7590);
nor U9626 (N_9626,N_6375,N_6534);
xnor U9627 (N_9627,N_8907,N_7181);
nor U9628 (N_9628,N_6272,N_7481);
nor U9629 (N_9629,N_7891,N_6193);
and U9630 (N_9630,N_8270,N_6884);
nor U9631 (N_9631,N_6360,N_7284);
nand U9632 (N_9632,N_7070,N_6363);
xnor U9633 (N_9633,N_6069,N_6889);
xnor U9634 (N_9634,N_7875,N_6549);
nor U9635 (N_9635,N_6227,N_7316);
or U9636 (N_9636,N_7447,N_8335);
xnor U9637 (N_9637,N_7145,N_6413);
and U9638 (N_9638,N_6310,N_6318);
xnor U9639 (N_9639,N_7959,N_6208);
or U9640 (N_9640,N_8436,N_8455);
nand U9641 (N_9641,N_6254,N_6216);
or U9642 (N_9642,N_7751,N_7243);
and U9643 (N_9643,N_7730,N_6311);
and U9644 (N_9644,N_8883,N_7792);
nor U9645 (N_9645,N_7514,N_8717);
or U9646 (N_9646,N_7510,N_6321);
xnor U9647 (N_9647,N_6435,N_6028);
nand U9648 (N_9648,N_7018,N_8082);
nor U9649 (N_9649,N_6404,N_8999);
and U9650 (N_9650,N_6776,N_7495);
and U9651 (N_9651,N_6377,N_6422);
or U9652 (N_9652,N_8506,N_6735);
and U9653 (N_9653,N_7988,N_7660);
nor U9654 (N_9654,N_7034,N_6983);
nor U9655 (N_9655,N_6403,N_6674);
or U9656 (N_9656,N_7197,N_6907);
xnor U9657 (N_9657,N_6136,N_8342);
and U9658 (N_9658,N_7386,N_8597);
and U9659 (N_9659,N_7319,N_7850);
xor U9660 (N_9660,N_6247,N_6498);
nor U9661 (N_9661,N_8450,N_6228);
and U9662 (N_9662,N_8658,N_6640);
nand U9663 (N_9663,N_8187,N_7863);
and U9664 (N_9664,N_6451,N_6026);
or U9665 (N_9665,N_8228,N_7985);
nor U9666 (N_9666,N_8945,N_7714);
xor U9667 (N_9667,N_8391,N_6164);
or U9668 (N_9668,N_6658,N_6051);
xnor U9669 (N_9669,N_8663,N_7408);
or U9670 (N_9670,N_7199,N_6546);
or U9671 (N_9671,N_8149,N_8469);
or U9672 (N_9672,N_7537,N_7261);
xnor U9673 (N_9673,N_7475,N_8592);
and U9674 (N_9674,N_7308,N_7972);
nor U9675 (N_9675,N_7543,N_8215);
nand U9676 (N_9676,N_7814,N_8135);
nor U9677 (N_9677,N_7073,N_7670);
xnor U9678 (N_9678,N_6068,N_8520);
and U9679 (N_9679,N_7441,N_6142);
or U9680 (N_9680,N_6004,N_7614);
xnor U9681 (N_9681,N_6048,N_7652);
or U9682 (N_9682,N_7027,N_6047);
and U9683 (N_9683,N_7116,N_7439);
or U9684 (N_9684,N_6368,N_7998);
nand U9685 (N_9685,N_6821,N_6680);
nor U9686 (N_9686,N_6595,N_8268);
nor U9687 (N_9687,N_6141,N_7107);
xor U9688 (N_9688,N_6727,N_8036);
nand U9689 (N_9689,N_8505,N_8001);
xnor U9690 (N_9690,N_8798,N_7264);
and U9691 (N_9691,N_8350,N_8737);
and U9692 (N_9692,N_6189,N_8424);
nor U9693 (N_9693,N_8562,N_8158);
and U9694 (N_9694,N_8797,N_8013);
or U9695 (N_9695,N_6170,N_6941);
nand U9696 (N_9696,N_6412,N_6330);
and U9697 (N_9697,N_7194,N_7138);
nor U9698 (N_9698,N_6881,N_6059);
xnor U9699 (N_9699,N_6039,N_8407);
nor U9700 (N_9700,N_7799,N_7780);
xor U9701 (N_9701,N_6393,N_8581);
xor U9702 (N_9702,N_8499,N_7423);
and U9703 (N_9703,N_8578,N_8755);
xnor U9704 (N_9704,N_8586,N_7497);
or U9705 (N_9705,N_7527,N_8949);
nand U9706 (N_9706,N_6329,N_8353);
xnor U9707 (N_9707,N_6527,N_6195);
nand U9708 (N_9708,N_7479,N_7053);
nand U9709 (N_9709,N_6180,N_7869);
or U9710 (N_9710,N_6388,N_8148);
and U9711 (N_9711,N_8704,N_8692);
or U9712 (N_9712,N_7062,N_8763);
nor U9713 (N_9713,N_6233,N_6848);
or U9714 (N_9714,N_7815,N_7581);
or U9715 (N_9715,N_8580,N_8745);
xor U9716 (N_9716,N_8729,N_8178);
nand U9717 (N_9717,N_8968,N_7162);
xnor U9718 (N_9718,N_7483,N_6126);
xor U9719 (N_9719,N_8047,N_7259);
and U9720 (N_9720,N_8605,N_7967);
and U9721 (N_9721,N_8042,N_8208);
and U9722 (N_9722,N_8266,N_7674);
xor U9723 (N_9723,N_6554,N_6156);
nand U9724 (N_9724,N_6123,N_7754);
and U9725 (N_9725,N_7463,N_7166);
or U9726 (N_9726,N_6339,N_7604);
and U9727 (N_9727,N_6496,N_8361);
nor U9728 (N_9728,N_7204,N_8769);
and U9729 (N_9729,N_8137,N_6621);
and U9730 (N_9730,N_8081,N_6856);
and U9731 (N_9731,N_8078,N_7567);
nor U9732 (N_9732,N_8743,N_7090);
and U9733 (N_9733,N_7054,N_8338);
nor U9734 (N_9734,N_6450,N_6437);
nor U9735 (N_9735,N_7599,N_6740);
nor U9736 (N_9736,N_7406,N_8972);
nor U9737 (N_9737,N_7338,N_6215);
nand U9738 (N_9738,N_7269,N_6165);
or U9739 (N_9739,N_6587,N_7828);
and U9740 (N_9740,N_8881,N_7218);
nand U9741 (N_9741,N_7417,N_8412);
and U9742 (N_9742,N_6934,N_6550);
and U9743 (N_9743,N_7574,N_8767);
or U9744 (N_9744,N_6046,N_8974);
and U9745 (N_9745,N_8864,N_6745);
xor U9746 (N_9746,N_8384,N_8218);
nand U9747 (N_9747,N_8457,N_7459);
xnor U9748 (N_9748,N_8030,N_6917);
nor U9749 (N_9749,N_7108,N_6732);
nand U9750 (N_9750,N_6706,N_7667);
nand U9751 (N_9751,N_6608,N_8831);
nor U9752 (N_9752,N_8072,N_7796);
xor U9753 (N_9753,N_7545,N_7781);
xor U9754 (N_9754,N_6001,N_7471);
nor U9755 (N_9755,N_8051,N_6332);
and U9756 (N_9756,N_8777,N_7178);
or U9757 (N_9757,N_6539,N_6815);
or U9758 (N_9758,N_8822,N_7956);
nand U9759 (N_9759,N_8309,N_8677);
nor U9760 (N_9760,N_6192,N_6023);
nor U9761 (N_9761,N_8884,N_8587);
or U9762 (N_9762,N_6243,N_8935);
and U9763 (N_9763,N_6533,N_6545);
xnor U9764 (N_9764,N_7470,N_7084);
xnor U9765 (N_9765,N_6371,N_7051);
nor U9766 (N_9766,N_7668,N_7026);
nor U9767 (N_9767,N_8134,N_8821);
nand U9768 (N_9768,N_6287,N_8223);
nor U9769 (N_9769,N_7609,N_6218);
or U9770 (N_9770,N_6859,N_7970);
or U9771 (N_9771,N_8316,N_8418);
and U9772 (N_9772,N_7297,N_8211);
xnor U9773 (N_9773,N_7994,N_8247);
and U9774 (N_9774,N_7515,N_7689);
xor U9775 (N_9775,N_8720,N_8170);
or U9776 (N_9776,N_8898,N_8144);
and U9777 (N_9777,N_7849,N_8836);
xor U9778 (N_9778,N_7677,N_7634);
and U9779 (N_9779,N_8304,N_6293);
nor U9780 (N_9780,N_6654,N_6693);
or U9781 (N_9781,N_6128,N_6390);
and U9782 (N_9782,N_8708,N_8538);
xnor U9783 (N_9783,N_7742,N_6358);
nor U9784 (N_9784,N_8542,N_6084);
or U9785 (N_9785,N_8559,N_6861);
and U9786 (N_9786,N_6729,N_6006);
and U9787 (N_9787,N_8199,N_8417);
or U9788 (N_9788,N_7741,N_8696);
or U9789 (N_9789,N_8012,N_6577);
and U9790 (N_9790,N_6689,N_6597);
nor U9791 (N_9791,N_7700,N_6389);
nor U9792 (N_9792,N_6637,N_7271);
nand U9793 (N_9793,N_8196,N_7779);
nand U9794 (N_9794,N_8163,N_6429);
or U9795 (N_9795,N_6210,N_6036);
nand U9796 (N_9796,N_6105,N_7117);
or U9797 (N_9797,N_8742,N_7465);
nand U9798 (N_9798,N_7922,N_6645);
nor U9799 (N_9799,N_6053,N_8438);
nand U9800 (N_9800,N_6984,N_6223);
and U9801 (N_9801,N_7842,N_6886);
nand U9802 (N_9802,N_8074,N_6044);
xnor U9803 (N_9803,N_8492,N_6506);
nand U9804 (N_9804,N_7085,N_7770);
nand U9805 (N_9805,N_8504,N_7605);
and U9806 (N_9806,N_7884,N_6491);
xnor U9807 (N_9807,N_7384,N_6098);
nand U9808 (N_9808,N_6480,N_7044);
and U9809 (N_9809,N_7691,N_8565);
nor U9810 (N_9810,N_7105,N_7402);
or U9811 (N_9811,N_8443,N_6675);
and U9812 (N_9812,N_8336,N_8277);
nor U9813 (N_9813,N_8891,N_8986);
nor U9814 (N_9814,N_7061,N_7317);
nand U9815 (N_9815,N_7977,N_8188);
and U9816 (N_9816,N_8358,N_6106);
xor U9817 (N_9817,N_8650,N_6960);
or U9818 (N_9818,N_8067,N_8037);
xor U9819 (N_9819,N_8246,N_6731);
or U9820 (N_9820,N_7651,N_8563);
nor U9821 (N_9821,N_8169,N_7055);
nor U9822 (N_9822,N_6589,N_7769);
xnor U9823 (N_9823,N_8104,N_8829);
and U9824 (N_9824,N_8659,N_8694);
xor U9825 (N_9825,N_7444,N_7314);
or U9826 (N_9826,N_7091,N_7868);
or U9827 (N_9827,N_8811,N_6396);
nor U9828 (N_9828,N_6966,N_8113);
and U9829 (N_9829,N_7703,N_7727);
nor U9830 (N_9830,N_7462,N_8726);
or U9831 (N_9831,N_8302,N_8007);
nor U9832 (N_9832,N_8371,N_8337);
and U9833 (N_9833,N_6906,N_8799);
and U9834 (N_9834,N_7717,N_6755);
or U9835 (N_9835,N_7339,N_6307);
or U9836 (N_9836,N_7332,N_8892);
or U9837 (N_9837,N_8689,N_6857);
nor U9838 (N_9838,N_8099,N_7232);
nor U9839 (N_9839,N_6556,N_6685);
and U9840 (N_9840,N_7520,N_6409);
nand U9841 (N_9841,N_8193,N_6066);
nand U9842 (N_9842,N_8510,N_6560);
nand U9843 (N_9843,N_6581,N_6081);
or U9844 (N_9844,N_6652,N_7899);
nand U9845 (N_9845,N_6786,N_7838);
or U9846 (N_9846,N_7136,N_6407);
and U9847 (N_9847,N_7935,N_8131);
xor U9848 (N_9848,N_7079,N_7330);
nor U9849 (N_9849,N_7489,N_6245);
and U9850 (N_9850,N_8326,N_6836);
or U9851 (N_9851,N_7235,N_6566);
nand U9852 (N_9852,N_7729,N_6849);
nand U9853 (N_9853,N_8010,N_6261);
or U9854 (N_9854,N_7549,N_7795);
nand U9855 (N_9855,N_6202,N_7246);
nand U9856 (N_9856,N_8096,N_7661);
nand U9857 (N_9857,N_6712,N_8327);
nand U9858 (N_9858,N_6514,N_7279);
xor U9859 (N_9859,N_6129,N_7202);
or U9860 (N_9860,N_7841,N_8728);
or U9861 (N_9861,N_6987,N_7926);
nand U9862 (N_9862,N_7938,N_7918);
or U9863 (N_9863,N_8004,N_7608);
xnor U9864 (N_9864,N_7360,N_7425);
or U9865 (N_9865,N_8877,N_8669);
xor U9866 (N_9866,N_8305,N_6241);
nand U9867 (N_9867,N_8044,N_7785);
nand U9868 (N_9868,N_7654,N_8100);
xor U9869 (N_9869,N_6431,N_8217);
nor U9870 (N_9870,N_8060,N_6509);
and U9871 (N_9871,N_7602,N_8649);
or U9872 (N_9872,N_7498,N_6323);
and U9873 (N_9873,N_6948,N_6603);
and U9874 (N_9874,N_6258,N_8593);
nor U9875 (N_9875,N_8934,N_8513);
nor U9876 (N_9876,N_6005,N_8609);
nor U9877 (N_9877,N_7065,N_7928);
nand U9878 (N_9878,N_7883,N_7887);
or U9879 (N_9879,N_7153,N_8981);
xor U9880 (N_9880,N_8622,N_7557);
nor U9881 (N_9881,N_8347,N_6299);
and U9882 (N_9882,N_6641,N_7187);
nor U9883 (N_9883,N_8919,N_6996);
nor U9884 (N_9884,N_8988,N_6708);
xor U9885 (N_9885,N_8548,N_6494);
xnor U9886 (N_9886,N_8394,N_6385);
nor U9887 (N_9887,N_6154,N_7438);
xnor U9888 (N_9888,N_6255,N_7057);
and U9889 (N_9889,N_6378,N_8301);
nand U9890 (N_9890,N_6265,N_8159);
nor U9891 (N_9891,N_8351,N_7251);
nor U9892 (N_9892,N_8794,N_8543);
nor U9893 (N_9893,N_8280,N_8043);
nand U9894 (N_9894,N_8080,N_8746);
nand U9895 (N_9895,N_7219,N_6336);
and U9896 (N_9896,N_6306,N_6248);
nand U9897 (N_9897,N_8240,N_8393);
or U9898 (N_9898,N_6551,N_6598);
and U9899 (N_9899,N_6419,N_6666);
nand U9900 (N_9900,N_6152,N_8470);
nor U9901 (N_9901,N_8508,N_8749);
xor U9902 (N_9902,N_7168,N_8034);
xnor U9903 (N_9903,N_6014,N_8924);
xor U9904 (N_9904,N_7361,N_8804);
xnor U9905 (N_9905,N_8088,N_6870);
nand U9906 (N_9906,N_8957,N_7963);
nand U9907 (N_9907,N_8774,N_6754);
or U9908 (N_9908,N_7050,N_8006);
or U9909 (N_9909,N_7784,N_7342);
nand U9910 (N_9910,N_6571,N_8296);
nand U9911 (N_9911,N_7810,N_7351);
and U9912 (N_9912,N_8496,N_7552);
nand U9913 (N_9913,N_6999,N_6441);
or U9914 (N_9914,N_6765,N_8165);
xor U9915 (N_9915,N_8990,N_8498);
xnor U9916 (N_9916,N_8117,N_8890);
and U9917 (N_9917,N_6548,N_7041);
nand U9918 (N_9918,N_7798,N_6772);
xor U9919 (N_9919,N_6703,N_8825);
nand U9920 (N_9920,N_6890,N_7512);
xnor U9921 (N_9921,N_8779,N_7158);
xor U9922 (N_9922,N_7518,N_8323);
and U9923 (N_9923,N_7383,N_8311);
nand U9924 (N_9924,N_8878,N_7418);
xor U9925 (N_9925,N_7964,N_7226);
or U9926 (N_9926,N_7455,N_7349);
or U9927 (N_9927,N_7984,N_6495);
nand U9928 (N_9928,N_8848,N_7978);
nor U9929 (N_9929,N_7832,N_8869);
nor U9930 (N_9930,N_6647,N_6798);
xnor U9931 (N_9931,N_8332,N_7033);
nand U9932 (N_9932,N_6140,N_6024);
nand U9933 (N_9933,N_6308,N_8982);
xor U9934 (N_9934,N_7149,N_8940);
nand U9935 (N_9935,N_7613,N_7516);
xnor U9936 (N_9936,N_7562,N_7064);
or U9937 (N_9937,N_7791,N_8340);
or U9938 (N_9938,N_8532,N_6911);
nor U9939 (N_9939,N_7763,N_8269);
xor U9940 (N_9940,N_7800,N_8842);
nor U9941 (N_9941,N_8180,N_8480);
xor U9942 (N_9942,N_7393,N_7101);
xor U9943 (N_9943,N_8345,N_7740);
and U9944 (N_9944,N_8413,N_8288);
nor U9945 (N_9945,N_6632,N_7203);
and U9946 (N_9946,N_7924,N_6854);
nand U9947 (N_9947,N_7015,N_7860);
and U9948 (N_9948,N_8645,N_6446);
nor U9949 (N_9949,N_6408,N_8946);
and U9950 (N_9950,N_8297,N_7118);
xnor U9951 (N_9951,N_7958,N_8190);
and U9952 (N_9952,N_6584,N_6809);
nand U9953 (N_9953,N_8066,N_7220);
nand U9954 (N_9954,N_6644,N_7776);
or U9955 (N_9955,N_6112,N_7936);
and U9956 (N_9956,N_8325,N_7077);
or U9957 (N_9957,N_6722,N_7024);
xor U9958 (N_9958,N_8161,N_6618);
or U9959 (N_9959,N_8555,N_8803);
nand U9960 (N_9960,N_8065,N_6997);
nand U9961 (N_9961,N_6541,N_8143);
nand U9962 (N_9962,N_6018,N_8408);
and U9963 (N_9963,N_6896,N_6346);
xnor U9964 (N_9964,N_8109,N_7548);
xnor U9965 (N_9965,N_6756,N_7946);
and U9966 (N_9966,N_7230,N_8698);
or U9967 (N_9967,N_8053,N_8932);
xnor U9968 (N_9968,N_8198,N_7535);
and U9969 (N_9969,N_7474,N_7645);
xnor U9970 (N_9970,N_8388,N_7504);
nor U9971 (N_9971,N_8790,N_8111);
nand U9972 (N_9972,N_8754,N_7615);
xor U9973 (N_9973,N_6839,N_8136);
nor U9974 (N_9974,N_6086,N_8841);
or U9975 (N_9975,N_7356,N_6781);
and U9976 (N_9976,N_6183,N_7909);
nor U9977 (N_9977,N_7511,N_6842);
nor U9978 (N_9978,N_8056,N_6818);
and U9979 (N_9979,N_8916,N_8524);
and U9980 (N_9980,N_6071,N_7161);
nand U9981 (N_9981,N_7861,N_7672);
nor U9982 (N_9982,N_7905,N_6974);
and U9983 (N_9983,N_7679,N_6444);
xor U9984 (N_9984,N_7588,N_8910);
xor U9985 (N_9985,N_6286,N_6445);
and U9986 (N_9986,N_6353,N_8812);
or U9987 (N_9987,N_8002,N_6635);
nand U9988 (N_9988,N_8678,N_7637);
xnor U9989 (N_9989,N_8521,N_6649);
nor U9990 (N_9990,N_8237,N_6707);
nand U9991 (N_9991,N_8750,N_7793);
or U9992 (N_9992,N_8515,N_6147);
nand U9993 (N_9993,N_7852,N_8879);
nand U9994 (N_9994,N_8203,N_6296);
nand U9995 (N_9995,N_8164,N_6430);
nand U9996 (N_9996,N_6562,N_7244);
nand U9997 (N_9997,N_6847,N_7932);
nand U9998 (N_9998,N_7382,N_8116);
xor U9999 (N_9999,N_8249,N_6483);
and U10000 (N_10000,N_8614,N_6931);
nand U10001 (N_10001,N_7368,N_7007);
or U10002 (N_10002,N_8029,N_6281);
and U10003 (N_10003,N_7253,N_6063);
xor U10004 (N_10004,N_8818,N_8306);
nor U10005 (N_10005,N_6125,N_6300);
xor U10006 (N_10006,N_6486,N_7047);
xor U10007 (N_10007,N_7189,N_7212);
or U10008 (N_10008,N_7807,N_8503);
xnor U10009 (N_10009,N_8429,N_6833);
and U10010 (N_10010,N_8628,N_7771);
xnor U10011 (N_10011,N_7862,N_8403);
nor U10012 (N_10012,N_8359,N_7612);
nor U10013 (N_10013,N_8531,N_6003);
and U10014 (N_10014,N_6939,N_8843);
and U10015 (N_10015,N_7643,N_7233);
nand U10016 (N_10016,N_6922,N_8862);
or U10017 (N_10017,N_6161,N_6405);
or U10018 (N_10018,N_8026,N_8971);
xnor U10019 (N_10019,N_7392,N_6008);
nor U10020 (N_10020,N_8186,N_7874);
nand U10021 (N_10021,N_6102,N_7083);
or U10022 (N_10022,N_6493,N_8996);
or U10023 (N_10023,N_8461,N_8245);
or U10024 (N_10024,N_8310,N_8182);
or U10025 (N_10025,N_7528,N_8902);
xor U10026 (N_10026,N_8784,N_7598);
nand U10027 (N_10027,N_6097,N_8642);
xor U10028 (N_10028,N_6395,N_8735);
or U10029 (N_10029,N_6908,N_8121);
or U10030 (N_10030,N_8201,N_7321);
or U10031 (N_10031,N_8456,N_8921);
and U10032 (N_10032,N_7205,N_6236);
and U10033 (N_10033,N_7211,N_8923);
and U10034 (N_10034,N_6115,N_8700);
nor U10035 (N_10035,N_7416,N_8415);
xnor U10036 (N_10036,N_8031,N_6547);
or U10037 (N_10037,N_7081,N_7121);
or U10038 (N_10038,N_8258,N_7752);
or U10039 (N_10039,N_7265,N_8716);
nor U10040 (N_10040,N_7437,N_8210);
or U10041 (N_10041,N_7327,N_7947);
xnor U10042 (N_10042,N_6213,N_8475);
nor U10043 (N_10043,N_7981,N_6590);
nand U10044 (N_10044,N_6843,N_8977);
and U10045 (N_10045,N_6952,N_7287);
xor U10046 (N_10046,N_8701,N_7201);
nor U10047 (N_10047,N_7765,N_8867);
or U10048 (N_10048,N_6211,N_7126);
or U10049 (N_10049,N_6678,N_6646);
nor U10050 (N_10050,N_6282,N_6295);
nand U10051 (N_10051,N_7678,N_8817);
xor U10052 (N_10052,N_6482,N_8381);
xor U10053 (N_10053,N_6120,N_8606);
nand U10054 (N_10054,N_6034,N_7519);
and U10055 (N_10055,N_8566,N_8616);
xor U10056 (N_10056,N_7603,N_6661);
and U10057 (N_10057,N_7930,N_8757);
xor U10058 (N_10058,N_8425,N_6037);
nand U10059 (N_10059,N_6470,N_7743);
and U10060 (N_10060,N_8275,N_6865);
and U10061 (N_10061,N_7950,N_6945);
or U10062 (N_10062,N_8257,N_7031);
and U10063 (N_10063,N_6967,N_7995);
or U10064 (N_10064,N_8960,N_7593);
nor U10065 (N_10065,N_7696,N_6753);
xnor U10066 (N_10066,N_7587,N_8992);
nor U10067 (N_10067,N_8289,N_7150);
nand U10068 (N_10068,N_6320,N_7534);
nor U10069 (N_10069,N_8851,N_8868);
nand U10070 (N_10070,N_8122,N_6238);
nor U10071 (N_10071,N_7146,N_8540);
nor U10072 (N_10072,N_6079,N_7362);
xor U10073 (N_10073,N_8671,N_8489);
xor U10074 (N_10074,N_7747,N_6521);
or U10075 (N_10075,N_6667,N_8094);
nand U10076 (N_10076,N_7000,N_7337);
and U10077 (N_10077,N_7805,N_8516);
and U10078 (N_10078,N_7322,N_7610);
and U10079 (N_10079,N_6277,N_8071);
nand U10080 (N_10080,N_8938,N_8646);
nor U10081 (N_10081,N_6795,N_6467);
xnor U10082 (N_10082,N_8579,N_6096);
nand U10083 (N_10083,N_6040,N_7407);
or U10084 (N_10084,N_6698,N_7484);
xor U10085 (N_10085,N_6348,N_6146);
and U10086 (N_10086,N_8775,N_7115);
nor U10087 (N_10087,N_7843,N_7767);
or U10088 (N_10088,N_6763,N_6155);
xor U10089 (N_10089,N_8447,N_7452);
xnor U10090 (N_10090,N_7262,N_6891);
nand U10091 (N_10091,N_6244,N_6485);
nand U10092 (N_10092,N_8162,N_7397);
and U10093 (N_10093,N_7941,N_7551);
xor U10094 (N_10094,N_6029,N_6747);
nor U10095 (N_10095,N_8362,N_6061);
nand U10096 (N_10096,N_6151,N_6915);
nand U10097 (N_10097,N_7159,N_7374);
and U10098 (N_10098,N_8376,N_6998);
or U10099 (N_10099,N_7469,N_8937);
nor U10100 (N_10100,N_6060,N_7982);
nand U10101 (N_10101,N_7155,N_7283);
or U10102 (N_10102,N_8356,N_8262);
xor U10103 (N_10103,N_8386,N_8613);
xnor U10104 (N_10104,N_7825,N_8387);
xnor U10105 (N_10105,N_6376,N_8126);
nand U10106 (N_10106,N_6768,N_6869);
nand U10107 (N_10107,N_6373,N_6914);
nand U10108 (N_10108,N_7229,N_6386);
nor U10109 (N_10109,N_7067,N_6179);
nor U10110 (N_10110,N_8680,N_6959);
and U10111 (N_10111,N_8861,N_7911);
and U10112 (N_10112,N_8160,N_7490);
nand U10113 (N_10113,N_7953,N_6148);
or U10114 (N_10114,N_6160,N_7500);
nand U10115 (N_10115,N_7170,N_6742);
nand U10116 (N_10116,N_8293,N_8400);
and U10117 (N_10117,N_6220,N_8286);
xor U10118 (N_10118,N_7302,N_6969);
or U10119 (N_10119,N_6302,N_8528);
or U10120 (N_10120,N_7623,N_8702);
and U10121 (N_10121,N_8621,N_8123);
and U10122 (N_10122,N_8409,N_6701);
nand U10123 (N_10123,N_7794,N_8329);
nand U10124 (N_10124,N_8636,N_8432);
xnor U10125 (N_10125,N_8406,N_6357);
and U10126 (N_10126,N_8715,N_7848);
xnor U10127 (N_10127,N_7477,N_7353);
nor U10128 (N_10128,N_6690,N_8976);
xor U10129 (N_10129,N_7945,N_6207);
xnor U10130 (N_10130,N_7124,N_7575);
nor U10131 (N_10131,N_6135,N_8089);
xor U10132 (N_10132,N_8399,N_8576);
xnor U10133 (N_10133,N_8315,N_8453);
nand U10134 (N_10134,N_6599,N_8561);
nor U10135 (N_10135,N_7241,N_6824);
or U10136 (N_10136,N_7147,N_8365);
or U10137 (N_10137,N_6749,N_8770);
or U10138 (N_10138,N_6790,N_6420);
and U10139 (N_10139,N_8625,N_8682);
or U10140 (N_10140,N_6752,N_7188);
xor U10141 (N_10141,N_8129,N_7296);
nand U10142 (N_10142,N_7910,N_7045);
or U10143 (N_10143,N_6888,N_8875);
nor U10144 (N_10144,N_6025,N_6288);
nand U10145 (N_10145,N_6033,N_6609);
and U10146 (N_10146,N_7043,N_8719);
xnor U10147 (N_10147,N_7119,N_8321);
nor U10148 (N_10148,N_8899,N_6716);
xor U10149 (N_10149,N_6873,N_7467);
or U10150 (N_10150,N_8250,N_6660);
or U10151 (N_10151,N_8713,N_8308);
xor U10152 (N_10152,N_8849,N_6672);
nand U10153 (N_10153,N_8303,N_7113);
nand U10154 (N_10154,N_8049,N_6131);
nand U10155 (N_10155,N_6817,N_8806);
and U10156 (N_10156,N_7156,N_6831);
xor U10157 (N_10157,N_7940,N_7358);
nand U10158 (N_10158,N_6668,N_7299);
nand U10159 (N_10159,N_6823,N_6778);
xor U10160 (N_10160,N_6520,N_7892);
and U10161 (N_10161,N_8005,N_7715);
xnor U10162 (N_10162,N_6497,N_7343);
xnor U10163 (N_10163,N_7530,N_6421);
nor U10164 (N_10164,N_7987,N_8523);
nor U10165 (N_10165,N_8759,N_7173);
nor U10166 (N_10166,N_6384,N_6923);
xor U10167 (N_10167,N_8766,N_8550);
or U10168 (N_10168,N_8772,N_8128);
nand U10169 (N_10169,N_7915,N_6530);
nor U10170 (N_10170,N_8564,N_8212);
xnor U10171 (N_10171,N_7595,N_8533);
nand U10172 (N_10172,N_6343,N_8421);
xor U10173 (N_10173,N_7818,N_6159);
nor U10174 (N_10174,N_8554,N_7732);
xor U10175 (N_10175,N_7686,N_7624);
nor U10176 (N_10176,N_8665,N_6825);
or U10177 (N_10177,N_7650,N_7962);
and U10178 (N_10178,N_7014,N_6230);
xor U10179 (N_10179,N_8539,N_7954);
and U10180 (N_10180,N_8876,N_6370);
or U10181 (N_10181,N_6400,N_8948);
nand U10182 (N_10182,N_7830,N_7336);
nand U10183 (N_10183,N_8556,N_6149);
xnor U10184 (N_10184,N_7036,N_8863);
xnor U10185 (N_10185,N_6094,N_7222);
and U10186 (N_10186,N_7913,N_6319);
or U10187 (N_10187,N_8674,N_6535);
or U10188 (N_10188,N_8446,N_6586);
nor U10189 (N_10189,N_6728,N_8229);
xor U10190 (N_10190,N_7172,N_7912);
or U10191 (N_10191,N_6524,N_8930);
and U10192 (N_10192,N_7089,N_6883);
and U10193 (N_10193,N_7436,N_8241);
xor U10194 (N_10194,N_6977,N_7801);
nor U10195 (N_10195,N_7773,N_7831);
and U10196 (N_10196,N_8925,N_7902);
xnor U10197 (N_10197,N_8604,N_7449);
nand U10198 (N_10198,N_7240,N_7607);
and U10199 (N_10199,N_8652,N_8488);
or U10200 (N_10200,N_6723,N_7578);
nand U10201 (N_10201,N_8965,N_8341);
or U10202 (N_10202,N_8271,N_8420);
xor U10203 (N_10203,N_8191,N_7820);
nor U10204 (N_10204,N_7461,N_8830);
or U10205 (N_10205,N_8235,N_6399);
xnor U10206 (N_10206,N_8181,N_6844);
and U10207 (N_10207,N_7415,N_6807);
nor U10208 (N_10208,N_7404,N_8961);
xor U10209 (N_10209,N_8035,N_8952);
nor U10210 (N_10210,N_6305,N_7764);
nand U10211 (N_10211,N_6937,N_6085);
and U10212 (N_10212,N_6529,N_6463);
xnor U10213 (N_10213,N_6611,N_7684);
nand U10214 (N_10214,N_8603,N_6279);
xor U10215 (N_10215,N_7141,N_7600);
and U10216 (N_10216,N_6239,N_6943);
or U10217 (N_10217,N_8871,N_6291);
and U10218 (N_10218,N_7778,N_6665);
nor U10219 (N_10219,N_6846,N_7215);
xor U10220 (N_10220,N_7616,N_8278);
and U10221 (N_10221,N_7409,N_8789);
or U10222 (N_10222,N_7132,N_8139);
nor U10223 (N_10223,N_8748,N_8918);
or U10224 (N_10224,N_6787,N_8638);
nor U10225 (N_10225,N_8317,N_7191);
xor U10226 (N_10226,N_6283,N_6124);
nand U10227 (N_10227,N_7120,N_6573);
xnor U10228 (N_10228,N_7078,N_7753);
or U10229 (N_10229,N_7571,N_6398);
nor U10230 (N_10230,N_7350,N_6280);
xor U10231 (N_10231,N_7971,N_6382);
nor U10232 (N_10232,N_8927,N_8585);
nand U10233 (N_10233,N_7473,N_7006);
nor U10234 (N_10234,N_6664,N_6078);
nor U10235 (N_10235,N_7719,N_6885);
and U10236 (N_10236,N_7817,N_6462);
or U10237 (N_10237,N_7003,N_7250);
xor U10238 (N_10238,N_8577,N_7658);
xnor U10239 (N_10239,N_8040,N_8239);
xor U10240 (N_10240,N_8662,N_6440);
or U10241 (N_10241,N_7702,N_6936);
nor U10242 (N_10242,N_7127,N_6950);
or U10243 (N_10243,N_7020,N_8828);
and U10244 (N_10244,N_8942,N_8640);
nand U10245 (N_10245,N_8172,N_6271);
and U10246 (N_10246,N_7625,N_6432);
nor U10247 (N_10247,N_7630,N_7487);
xnor U10248 (N_10248,N_8259,N_7933);
xor U10249 (N_10249,N_6792,N_6334);
nor U10250 (N_10250,N_6290,N_8846);
and U10251 (N_10251,N_8295,N_7482);
and U10252 (N_10252,N_6174,N_7378);
nor U10253 (N_10253,N_7325,N_8814);
or U10254 (N_10254,N_7217,N_6297);
or U10255 (N_10255,N_8107,N_7010);
or U10256 (N_10256,N_8541,N_6617);
and U10257 (N_10257,N_6197,N_8226);
nand U10258 (N_10258,N_6452,N_8349);
nor U10259 (N_10259,N_7134,N_6793);
and U10260 (N_10260,N_8731,N_8534);
nor U10261 (N_10261,N_7627,N_8987);
nor U10262 (N_10262,N_8711,N_6246);
nand U10263 (N_10263,N_8194,N_8445);
nor U10264 (N_10264,N_8787,N_6510);
or U10265 (N_10265,N_6049,N_8057);
nor U10266 (N_10266,N_8017,N_6713);
nand U10267 (N_10267,N_6801,N_6614);
xnor U10268 (N_10268,N_7348,N_7968);
xnor U10269 (N_10269,N_7248,N_7488);
or U10270 (N_10270,N_6091,N_8683);
and U10271 (N_10271,N_8264,N_7413);
and U10272 (N_10272,N_8571,N_6276);
xnor U10273 (N_10273,N_8225,N_6270);
or U10274 (N_10274,N_7583,N_8435);
nor U10275 (N_10275,N_7896,N_6349);
nand U10276 (N_10276,N_6624,N_7676);
nand U10277 (N_10277,N_7655,N_7558);
or U10278 (N_10278,N_6103,N_7565);
and U10279 (N_10279,N_8070,N_6448);
or U10280 (N_10280,N_7846,N_6639);
xor U10281 (N_10281,N_7285,N_6316);
nand U10282 (N_10282,N_6656,N_6957);
and U10283 (N_10283,N_8887,N_7628);
or U10284 (N_10284,N_7214,N_8661);
and U10285 (N_10285,N_8063,N_6538);
nor U10286 (N_10286,N_8865,N_7542);
or U10287 (N_10287,N_8947,N_8076);
or U10288 (N_10288,N_6829,N_8426);
nand U10289 (N_10289,N_8752,N_6719);
nand U10290 (N_10290,N_8922,N_7642);
nand U10291 (N_10291,N_8175,N_7227);
nand U10292 (N_10292,N_6052,N_6406);
xnor U10293 (N_10293,N_8024,N_8805);
nor U10294 (N_10294,N_8714,N_6259);
nor U10295 (N_10295,N_8984,N_6741);
or U10296 (N_10296,N_7889,N_7300);
and U10297 (N_10297,N_6194,N_7649);
nand U10298 (N_10298,N_7695,N_6021);
or U10299 (N_10299,N_8474,N_7195);
xnor U10300 (N_10300,N_6569,N_8959);
or U10301 (N_10301,N_7584,N_7369);
xor U10302 (N_10302,N_8813,N_7908);
or U10303 (N_10303,N_6602,N_8951);
and U10304 (N_10304,N_6575,N_6540);
and U10305 (N_10305,N_7746,N_6559);
or U10306 (N_10306,N_6010,N_8596);
xnor U10307 (N_10307,N_8468,N_6250);
nor U10308 (N_10308,N_8333,N_6820);
nand U10309 (N_10309,N_7705,N_6583);
or U10310 (N_10310,N_6832,N_6725);
or U10311 (N_10311,N_6428,N_7182);
nand U10312 (N_10312,N_8261,N_8075);
nor U10313 (N_10313,N_8150,N_6813);
xor U10314 (N_10314,N_6275,N_7782);
xor U10315 (N_10315,N_8256,N_6607);
nor U10316 (N_10316,N_7761,N_7422);
or U10317 (N_10317,N_7790,N_6402);
xnor U10318 (N_10318,N_7333,N_7502);
and U10319 (N_10319,N_8462,N_7555);
nand U10320 (N_10320,N_6537,N_7725);
nor U10321 (N_10321,N_8765,N_7680);
xnor U10322 (N_10322,N_8796,N_7421);
or U10323 (N_10323,N_7334,N_6263);
or U10324 (N_10324,N_7596,N_7237);
or U10325 (N_10325,N_7580,N_8517);
nand U10326 (N_10326,N_8234,N_8758);
nand U10327 (N_10327,N_7125,N_7758);
nand U10328 (N_10328,N_8103,N_8440);
xnor U10329 (N_10329,N_8216,N_7335);
and U10330 (N_10330,N_8410,N_7254);
nand U10331 (N_10331,N_6988,N_8705);
and U10332 (N_10332,N_7692,N_8307);
and U10333 (N_10333,N_8274,N_7659);
and U10334 (N_10334,N_8567,N_7568);
and U10335 (N_10335,N_8019,N_7547);
xor U10336 (N_10336,N_8380,N_6337);
and U10337 (N_10337,N_6072,N_7109);
or U10338 (N_10338,N_7177,N_6013);
and U10339 (N_10339,N_8346,N_7129);
nand U10340 (N_10340,N_8441,N_7320);
and U10341 (N_10341,N_6056,N_6954);
xnor U10342 (N_10342,N_7326,N_7955);
and U10343 (N_10343,N_7524,N_6114);
or U10344 (N_10344,N_7307,N_6946);
and U10345 (N_10345,N_8856,N_8648);
xor U10346 (N_10346,N_8449,N_8312);
nand U10347 (N_10347,N_8819,N_6932);
and U10348 (N_10348,N_8251,N_6488);
nand U10349 (N_10349,N_7420,N_6806);
nor U10350 (N_10350,N_7871,N_8514);
xnor U10351 (N_10351,N_8838,N_7966);
and U10352 (N_10352,N_8157,N_6852);
nor U10353 (N_10353,N_6746,N_8736);
nand U10354 (N_10354,N_8118,N_7032);
or U10355 (N_10355,N_8901,N_8993);
nor U10356 (N_10356,N_8263,N_6035);
nor U10357 (N_10357,N_7460,N_6119);
nor U10358 (N_10358,N_6327,N_7311);
and U10359 (N_10359,N_8617,N_7949);
and U10360 (N_10360,N_6438,N_7569);
and U10361 (N_10361,N_7904,N_7429);
xor U10362 (N_10362,N_7468,N_7664);
and U10363 (N_10363,N_8570,N_6929);
nor U10364 (N_10364,N_8077,N_6733);
or U10365 (N_10365,N_8507,N_8827);
xor U10366 (N_10366,N_6947,N_6460);
or U10367 (N_10367,N_7058,N_8722);
and U10368 (N_10368,N_6900,N_7508);
nand U10369 (N_10369,N_6471,N_6478);
or U10370 (N_10370,N_8672,N_6673);
nor U10371 (N_10371,N_8206,N_7290);
xor U10372 (N_10372,N_8583,N_7636);
and U10373 (N_10373,N_6274,N_7328);
nor U10374 (N_10374,N_6766,N_6898);
nor U10375 (N_10375,N_6416,N_7647);
nor U10376 (N_10376,N_6910,N_6924);
or U10377 (N_10377,N_8792,N_8594);
xnor U10378 (N_10378,N_6198,N_8179);
nand U10379 (N_10379,N_7305,N_8753);
xor U10380 (N_10380,N_6074,N_6720);
nand U10381 (N_10381,N_6116,N_7139);
nor U10382 (N_10382,N_6217,N_8482);
and U10383 (N_10383,N_6182,N_6681);
or U10384 (N_10384,N_7879,N_6110);
or U10385 (N_10385,N_7412,N_7152);
xor U10386 (N_10386,N_7391,N_6089);
xnor U10387 (N_10387,N_7224,N_6994);
nor U10388 (N_10388,N_8699,N_7371);
nand U10389 (N_10389,N_6345,N_8021);
nor U10390 (N_10390,N_6855,N_7721);
or U10391 (N_10391,N_7289,N_7687);
or U10392 (N_10392,N_8773,N_8411);
xor U10393 (N_10393,N_8283,N_7282);
xor U10394 (N_10394,N_6169,N_8544);
xnor U10395 (N_10395,N_7274,N_6682);
and U10396 (N_10396,N_6264,N_7900);
or U10397 (N_10397,N_7491,N_6905);
nor U10398 (N_10398,N_7716,N_6038);
nand U10399 (N_10399,N_8048,N_7137);
xor U10400 (N_10400,N_7750,N_8970);
nor U10401 (N_10401,N_7760,N_7942);
and U10402 (N_10402,N_8710,N_8318);
and U10403 (N_10403,N_6093,N_8637);
and U10404 (N_10404,N_7701,N_6893);
or U10405 (N_10405,N_6391,N_7160);
nand U10406 (N_10406,N_7075,N_6473);
or U10407 (N_10407,N_7559,N_6638);
xor U10408 (N_10408,N_8185,N_6592);
or U10409 (N_10409,N_7076,N_6964);
nor U10410 (N_10410,N_7586,N_6981);
xnor U10411 (N_10411,N_7920,N_6186);
or U10412 (N_10412,N_7755,N_6372);
and U10413 (N_10413,N_8222,N_7494);
nor U10414 (N_10414,N_6508,N_7183);
nor U10415 (N_10415,N_8392,N_8855);
nor U10416 (N_10416,N_7662,N_6057);
xnor U10417 (N_10417,N_6266,N_6532);
and U10418 (N_10418,N_8368,N_8909);
xnor U10419 (N_10419,N_8911,N_7666);
nor U10420 (N_10420,N_6476,N_7270);
and U10421 (N_10421,N_6133,N_6956);
nand U10422 (N_10422,N_6121,N_6076);
or U10423 (N_10423,N_8962,N_8670);
or U10424 (N_10424,N_8518,N_6935);
xnor U10425 (N_10425,N_6814,N_8734);
nor U10426 (N_10426,N_8882,N_6704);
nand U10427 (N_10427,N_7665,N_7529);
nand U10428 (N_10428,N_7633,N_8807);
and U10429 (N_10429,N_6724,N_6902);
or U10430 (N_10430,N_6930,N_6788);
xor U10431 (N_10431,N_8366,N_8087);
xnor U10432 (N_10432,N_8227,N_6973);
and U10433 (N_10433,N_7039,N_7726);
xor U10434 (N_10434,N_6750,N_6802);
nand U10435 (N_10435,N_8330,N_8584);
nand U10436 (N_10436,N_8738,N_7052);
or U10437 (N_10437,N_6604,N_6804);
and U10438 (N_10438,N_7619,N_6394);
and U10439 (N_10439,N_6294,N_6285);
nor U10440 (N_10440,N_8434,N_7389);
and U10441 (N_10441,N_6492,N_6309);
xor U10442 (N_10442,N_8788,N_8684);
or U10443 (N_10443,N_7979,N_7744);
nand U10444 (N_10444,N_8630,N_7969);
nor U10445 (N_10445,N_8721,N_8472);
nand U10446 (N_10446,N_7104,N_7657);
nor U10447 (N_10447,N_7011,N_8509);
and U10448 (N_10448,N_8025,N_8667);
nor U10449 (N_10449,N_7419,N_6841);
or U10450 (N_10450,N_7405,N_8046);
xnor U10451 (N_10451,N_7671,N_8639);
nor U10452 (N_10452,N_7783,N_7929);
nand U10453 (N_10453,N_6634,N_7693);
and U10454 (N_10454,N_8405,N_8740);
nor U10455 (N_10455,N_8526,N_6187);
nand U10456 (N_10456,N_7509,N_6630);
nand U10457 (N_10457,N_8599,N_7975);
or U10458 (N_10458,N_8681,N_8145);
xor U10459 (N_10459,N_6249,N_6253);
and U10460 (N_10460,N_7775,N_8352);
and U10461 (N_10461,N_6229,N_7675);
nor U10462 (N_10462,N_6990,N_8220);
nor U10463 (N_10463,N_8027,N_8815);
nor U10464 (N_10464,N_8660,N_8656);
nor U10465 (N_10465,N_6684,N_6909);
nor U10466 (N_10466,N_7016,N_7093);
and U10467 (N_10467,N_6012,N_6811);
nor U10468 (N_10468,N_7151,N_8647);
nand U10469 (N_10469,N_6596,N_6588);
or U10470 (N_10470,N_6354,N_6770);
or U10471 (N_10471,N_8810,N_7098);
nor U10472 (N_10472,N_7210,N_6769);
xnor U10473 (N_10473,N_7486,N_8943);
nand U10474 (N_10474,N_8536,N_7897);
xor U10475 (N_10475,N_6944,N_7411);
or U10476 (N_10476,N_7367,N_6303);
nor U10477 (N_10477,N_6574,N_8360);
xor U10478 (N_10478,N_7099,N_7656);
xor U10479 (N_10479,N_6117,N_7056);
nor U10480 (N_10480,N_8370,N_7249);
xnor U10481 (N_10481,N_6863,N_6177);
or U10482 (N_10482,N_7277,N_7135);
or U10483 (N_10483,N_6764,N_6325);
and U10484 (N_10484,N_8343,N_7294);
and U10485 (N_10485,N_6175,N_6163);
xor U10486 (N_10486,N_6743,N_8847);
xnor U10487 (N_10487,N_6761,N_6144);
nor U10488 (N_10488,N_7472,N_6256);
nor U10489 (N_10489,N_8917,N_7523);
or U10490 (N_10490,N_8969,N_7390);
and U10491 (N_10491,N_7621,N_8809);
xnor U10492 (N_10492,N_8085,N_8023);
xor U10493 (N_10493,N_7822,N_8112);
or U10494 (N_10494,N_7252,N_8041);
or U10495 (N_10495,N_6380,N_8595);
nor U10496 (N_10496,N_8958,N_6874);
nand U10497 (N_10497,N_6351,N_7315);
nor U10498 (N_10498,N_7937,N_7174);
or U10499 (N_10499,N_8582,N_8983);
xnor U10500 (N_10500,N_8071,N_8206);
nand U10501 (N_10501,N_6307,N_6557);
nor U10502 (N_10502,N_7740,N_7044);
xor U10503 (N_10503,N_8704,N_6708);
xor U10504 (N_10504,N_7087,N_8013);
or U10505 (N_10505,N_7912,N_8638);
xor U10506 (N_10506,N_8488,N_8351);
or U10507 (N_10507,N_6718,N_6263);
and U10508 (N_10508,N_6244,N_7751);
and U10509 (N_10509,N_7164,N_6714);
xnor U10510 (N_10510,N_6894,N_8493);
or U10511 (N_10511,N_8226,N_7516);
nor U10512 (N_10512,N_8943,N_8363);
or U10513 (N_10513,N_6072,N_7429);
and U10514 (N_10514,N_6013,N_8281);
or U10515 (N_10515,N_7855,N_6064);
xor U10516 (N_10516,N_6085,N_6010);
nor U10517 (N_10517,N_8172,N_7876);
nand U10518 (N_10518,N_6006,N_6051);
or U10519 (N_10519,N_7962,N_8657);
or U10520 (N_10520,N_8914,N_7666);
nor U10521 (N_10521,N_8608,N_6324);
nor U10522 (N_10522,N_6811,N_8706);
and U10523 (N_10523,N_6681,N_6401);
nand U10524 (N_10524,N_6772,N_6370);
xnor U10525 (N_10525,N_6384,N_6929);
or U10526 (N_10526,N_6908,N_8376);
or U10527 (N_10527,N_6633,N_6201);
nand U10528 (N_10528,N_7147,N_6867);
nand U10529 (N_10529,N_8739,N_8043);
nor U10530 (N_10530,N_6763,N_7805);
nand U10531 (N_10531,N_7751,N_8879);
and U10532 (N_10532,N_8719,N_6396);
nor U10533 (N_10533,N_6019,N_7237);
and U10534 (N_10534,N_8107,N_8957);
and U10535 (N_10535,N_7446,N_6460);
or U10536 (N_10536,N_6940,N_7699);
and U10537 (N_10537,N_6676,N_7544);
or U10538 (N_10538,N_6227,N_8455);
and U10539 (N_10539,N_7385,N_8783);
nor U10540 (N_10540,N_6124,N_7628);
or U10541 (N_10541,N_6645,N_7333);
or U10542 (N_10542,N_6992,N_6999);
nand U10543 (N_10543,N_7554,N_8545);
nand U10544 (N_10544,N_6769,N_8949);
and U10545 (N_10545,N_6684,N_6075);
or U10546 (N_10546,N_6170,N_6023);
or U10547 (N_10547,N_7507,N_8331);
xor U10548 (N_10548,N_6142,N_7350);
xor U10549 (N_10549,N_7633,N_7989);
and U10550 (N_10550,N_6615,N_8938);
nand U10551 (N_10551,N_7948,N_8928);
or U10552 (N_10552,N_6670,N_6787);
xor U10553 (N_10553,N_8766,N_6930);
nor U10554 (N_10554,N_7846,N_6782);
nand U10555 (N_10555,N_8036,N_7035);
or U10556 (N_10556,N_6262,N_6220);
or U10557 (N_10557,N_6037,N_7665);
or U10558 (N_10558,N_7579,N_8854);
and U10559 (N_10559,N_6831,N_8240);
and U10560 (N_10560,N_7061,N_6534);
and U10561 (N_10561,N_6647,N_7567);
nor U10562 (N_10562,N_8585,N_7186);
nor U10563 (N_10563,N_7948,N_7342);
or U10564 (N_10564,N_8486,N_6926);
and U10565 (N_10565,N_7216,N_6482);
nand U10566 (N_10566,N_6107,N_6402);
xnor U10567 (N_10567,N_6929,N_6039);
nand U10568 (N_10568,N_7822,N_8278);
and U10569 (N_10569,N_6157,N_6455);
nor U10570 (N_10570,N_6398,N_6186);
and U10571 (N_10571,N_8799,N_7724);
and U10572 (N_10572,N_8080,N_7754);
or U10573 (N_10573,N_6171,N_6418);
or U10574 (N_10574,N_8625,N_7663);
and U10575 (N_10575,N_6395,N_6067);
xor U10576 (N_10576,N_6497,N_6344);
nand U10577 (N_10577,N_6369,N_7852);
or U10578 (N_10578,N_6754,N_7754);
nand U10579 (N_10579,N_8198,N_7983);
xnor U10580 (N_10580,N_8463,N_7925);
nand U10581 (N_10581,N_6994,N_7424);
or U10582 (N_10582,N_7456,N_8842);
and U10583 (N_10583,N_8228,N_7469);
or U10584 (N_10584,N_7585,N_6137);
nand U10585 (N_10585,N_7238,N_8101);
and U10586 (N_10586,N_8412,N_6725);
and U10587 (N_10587,N_6764,N_7827);
or U10588 (N_10588,N_8130,N_8645);
xnor U10589 (N_10589,N_7423,N_6647);
xnor U10590 (N_10590,N_7146,N_7221);
xor U10591 (N_10591,N_7225,N_6802);
and U10592 (N_10592,N_7590,N_7077);
or U10593 (N_10593,N_7888,N_6596);
nor U10594 (N_10594,N_7397,N_6657);
and U10595 (N_10595,N_6784,N_6107);
nand U10596 (N_10596,N_6383,N_8798);
and U10597 (N_10597,N_8009,N_7326);
xnor U10598 (N_10598,N_6137,N_7341);
nand U10599 (N_10599,N_8090,N_6591);
xnor U10600 (N_10600,N_8458,N_7383);
or U10601 (N_10601,N_8880,N_7505);
xnor U10602 (N_10602,N_8963,N_7754);
and U10603 (N_10603,N_6815,N_8082);
nand U10604 (N_10604,N_8293,N_8584);
nand U10605 (N_10605,N_8832,N_8999);
and U10606 (N_10606,N_6925,N_7391);
nand U10607 (N_10607,N_7774,N_7859);
nand U10608 (N_10608,N_6096,N_8422);
or U10609 (N_10609,N_8294,N_6814);
or U10610 (N_10610,N_7958,N_6283);
or U10611 (N_10611,N_6164,N_8946);
nor U10612 (N_10612,N_6814,N_8389);
or U10613 (N_10613,N_8771,N_8777);
or U10614 (N_10614,N_7841,N_7206);
nor U10615 (N_10615,N_8702,N_6682);
nand U10616 (N_10616,N_7022,N_6846);
or U10617 (N_10617,N_8526,N_8789);
xor U10618 (N_10618,N_7589,N_6938);
or U10619 (N_10619,N_6853,N_6732);
nand U10620 (N_10620,N_6519,N_6509);
and U10621 (N_10621,N_8773,N_6453);
or U10622 (N_10622,N_8166,N_7719);
xnor U10623 (N_10623,N_6997,N_6256);
and U10624 (N_10624,N_8958,N_8205);
nor U10625 (N_10625,N_6809,N_8974);
and U10626 (N_10626,N_6828,N_6135);
xnor U10627 (N_10627,N_8725,N_6028);
or U10628 (N_10628,N_7690,N_6565);
nor U10629 (N_10629,N_7655,N_7184);
nor U10630 (N_10630,N_7288,N_8884);
and U10631 (N_10631,N_8616,N_7254);
nand U10632 (N_10632,N_8014,N_8088);
xor U10633 (N_10633,N_8084,N_8495);
nand U10634 (N_10634,N_6728,N_8825);
nor U10635 (N_10635,N_8438,N_7603);
xnor U10636 (N_10636,N_6630,N_8912);
or U10637 (N_10637,N_6084,N_7797);
nor U10638 (N_10638,N_8893,N_6916);
nand U10639 (N_10639,N_7034,N_6015);
nor U10640 (N_10640,N_8676,N_7704);
and U10641 (N_10641,N_8080,N_7004);
xnor U10642 (N_10642,N_6569,N_8044);
or U10643 (N_10643,N_6417,N_7059);
nand U10644 (N_10644,N_7117,N_6524);
and U10645 (N_10645,N_7670,N_8292);
nor U10646 (N_10646,N_8401,N_8458);
and U10647 (N_10647,N_7658,N_6026);
nor U10648 (N_10648,N_6746,N_8002);
and U10649 (N_10649,N_8873,N_7850);
and U10650 (N_10650,N_7589,N_8727);
nor U10651 (N_10651,N_7744,N_7641);
or U10652 (N_10652,N_7737,N_8474);
nand U10653 (N_10653,N_6567,N_6210);
xnor U10654 (N_10654,N_6324,N_7084);
or U10655 (N_10655,N_7929,N_7803);
and U10656 (N_10656,N_8475,N_6555);
and U10657 (N_10657,N_7580,N_8873);
and U10658 (N_10658,N_8737,N_8724);
or U10659 (N_10659,N_8116,N_8248);
xnor U10660 (N_10660,N_8743,N_8935);
nand U10661 (N_10661,N_7838,N_7303);
xor U10662 (N_10662,N_7048,N_7605);
and U10663 (N_10663,N_7302,N_8030);
and U10664 (N_10664,N_7088,N_6710);
and U10665 (N_10665,N_6119,N_8390);
and U10666 (N_10666,N_7331,N_8445);
nor U10667 (N_10667,N_7198,N_6387);
nand U10668 (N_10668,N_8594,N_7882);
nand U10669 (N_10669,N_6545,N_6256);
xor U10670 (N_10670,N_6427,N_7154);
or U10671 (N_10671,N_7006,N_8658);
xnor U10672 (N_10672,N_6529,N_6818);
or U10673 (N_10673,N_6285,N_7482);
nand U10674 (N_10674,N_6212,N_7039);
or U10675 (N_10675,N_7314,N_7310);
and U10676 (N_10676,N_7936,N_8998);
and U10677 (N_10677,N_7603,N_8957);
nor U10678 (N_10678,N_8118,N_7041);
xnor U10679 (N_10679,N_6759,N_6619);
xor U10680 (N_10680,N_8251,N_6838);
nor U10681 (N_10681,N_8347,N_8153);
nor U10682 (N_10682,N_8129,N_8555);
and U10683 (N_10683,N_8188,N_7843);
or U10684 (N_10684,N_7025,N_8511);
xnor U10685 (N_10685,N_7487,N_8931);
nor U10686 (N_10686,N_6109,N_8287);
or U10687 (N_10687,N_7908,N_7396);
nor U10688 (N_10688,N_6272,N_6867);
nand U10689 (N_10689,N_7572,N_7112);
and U10690 (N_10690,N_6862,N_8075);
nand U10691 (N_10691,N_7101,N_6857);
and U10692 (N_10692,N_8626,N_8648);
xnor U10693 (N_10693,N_7503,N_8435);
xnor U10694 (N_10694,N_7577,N_8864);
nor U10695 (N_10695,N_8835,N_6600);
xor U10696 (N_10696,N_8142,N_6603);
xnor U10697 (N_10697,N_8157,N_6314);
nand U10698 (N_10698,N_8954,N_7728);
xnor U10699 (N_10699,N_7416,N_8930);
nand U10700 (N_10700,N_7118,N_8576);
and U10701 (N_10701,N_8712,N_7887);
and U10702 (N_10702,N_7545,N_7724);
nand U10703 (N_10703,N_6869,N_7493);
nor U10704 (N_10704,N_6417,N_6987);
nand U10705 (N_10705,N_7329,N_6225);
nand U10706 (N_10706,N_6815,N_8833);
and U10707 (N_10707,N_8865,N_6276);
xnor U10708 (N_10708,N_6761,N_8505);
or U10709 (N_10709,N_6556,N_6593);
and U10710 (N_10710,N_8916,N_7663);
nand U10711 (N_10711,N_8737,N_8852);
nor U10712 (N_10712,N_8807,N_8860);
or U10713 (N_10713,N_7818,N_8620);
xor U10714 (N_10714,N_6855,N_6913);
and U10715 (N_10715,N_7466,N_7365);
and U10716 (N_10716,N_7001,N_8419);
xor U10717 (N_10717,N_7113,N_8300);
and U10718 (N_10718,N_8901,N_8319);
and U10719 (N_10719,N_7469,N_7364);
nor U10720 (N_10720,N_8535,N_6848);
or U10721 (N_10721,N_6711,N_7411);
nand U10722 (N_10722,N_6334,N_7034);
or U10723 (N_10723,N_7140,N_8436);
nor U10724 (N_10724,N_8248,N_7637);
and U10725 (N_10725,N_7736,N_7974);
nor U10726 (N_10726,N_8035,N_7033);
and U10727 (N_10727,N_8599,N_7883);
and U10728 (N_10728,N_8417,N_6810);
or U10729 (N_10729,N_7359,N_6311);
nand U10730 (N_10730,N_6870,N_7577);
and U10731 (N_10731,N_6027,N_8829);
and U10732 (N_10732,N_7358,N_8069);
and U10733 (N_10733,N_6171,N_7867);
nand U10734 (N_10734,N_6486,N_6034);
nand U10735 (N_10735,N_8905,N_6022);
nor U10736 (N_10736,N_7569,N_6946);
and U10737 (N_10737,N_7064,N_6468);
nor U10738 (N_10738,N_7499,N_7244);
or U10739 (N_10739,N_8789,N_7508);
and U10740 (N_10740,N_7251,N_6151);
xnor U10741 (N_10741,N_8062,N_8154);
or U10742 (N_10742,N_6544,N_7169);
nor U10743 (N_10743,N_6606,N_6447);
or U10744 (N_10744,N_7173,N_8398);
nand U10745 (N_10745,N_6494,N_8251);
and U10746 (N_10746,N_7790,N_6200);
and U10747 (N_10747,N_6786,N_6127);
nand U10748 (N_10748,N_8310,N_8872);
nor U10749 (N_10749,N_8267,N_8948);
nand U10750 (N_10750,N_8054,N_7690);
xnor U10751 (N_10751,N_6278,N_7674);
nor U10752 (N_10752,N_6814,N_7589);
or U10753 (N_10753,N_8654,N_7598);
or U10754 (N_10754,N_7819,N_7089);
nor U10755 (N_10755,N_8012,N_6942);
xor U10756 (N_10756,N_7721,N_8739);
and U10757 (N_10757,N_8202,N_7719);
or U10758 (N_10758,N_6418,N_8615);
and U10759 (N_10759,N_6385,N_6321);
nand U10760 (N_10760,N_6620,N_6148);
and U10761 (N_10761,N_7130,N_7345);
nor U10762 (N_10762,N_6004,N_8406);
nand U10763 (N_10763,N_7784,N_7748);
xor U10764 (N_10764,N_6583,N_8497);
nand U10765 (N_10765,N_8492,N_7505);
and U10766 (N_10766,N_6674,N_8892);
nand U10767 (N_10767,N_7847,N_8403);
and U10768 (N_10768,N_8701,N_8803);
and U10769 (N_10769,N_6717,N_6017);
nand U10770 (N_10770,N_6279,N_6999);
or U10771 (N_10771,N_6049,N_7706);
and U10772 (N_10772,N_7043,N_6024);
and U10773 (N_10773,N_6443,N_7667);
nor U10774 (N_10774,N_7208,N_8369);
nor U10775 (N_10775,N_8053,N_6525);
nand U10776 (N_10776,N_7234,N_7784);
and U10777 (N_10777,N_8507,N_6926);
or U10778 (N_10778,N_7028,N_6964);
or U10779 (N_10779,N_8616,N_7785);
nand U10780 (N_10780,N_6195,N_6587);
nand U10781 (N_10781,N_6727,N_8004);
nand U10782 (N_10782,N_8742,N_8248);
or U10783 (N_10783,N_6271,N_6734);
nand U10784 (N_10784,N_8029,N_6121);
and U10785 (N_10785,N_6817,N_7073);
or U10786 (N_10786,N_8121,N_6363);
nor U10787 (N_10787,N_7674,N_7595);
nor U10788 (N_10788,N_7159,N_6168);
xor U10789 (N_10789,N_8780,N_8717);
or U10790 (N_10790,N_7399,N_7292);
and U10791 (N_10791,N_7949,N_7012);
or U10792 (N_10792,N_8045,N_6663);
or U10793 (N_10793,N_8280,N_8680);
or U10794 (N_10794,N_8079,N_8203);
xnor U10795 (N_10795,N_8079,N_6078);
xnor U10796 (N_10796,N_8795,N_6559);
nand U10797 (N_10797,N_6896,N_8660);
nand U10798 (N_10798,N_7829,N_6334);
xnor U10799 (N_10799,N_8693,N_6122);
nor U10800 (N_10800,N_6840,N_6446);
nand U10801 (N_10801,N_8097,N_7550);
nor U10802 (N_10802,N_8233,N_6424);
and U10803 (N_10803,N_8177,N_8109);
and U10804 (N_10804,N_6242,N_8137);
nand U10805 (N_10805,N_8401,N_8288);
xor U10806 (N_10806,N_8366,N_7628);
nor U10807 (N_10807,N_8371,N_8477);
or U10808 (N_10808,N_6831,N_7574);
or U10809 (N_10809,N_6451,N_7764);
nor U10810 (N_10810,N_6303,N_6291);
or U10811 (N_10811,N_8277,N_6534);
nor U10812 (N_10812,N_8308,N_8467);
and U10813 (N_10813,N_8801,N_8984);
or U10814 (N_10814,N_7040,N_6259);
or U10815 (N_10815,N_8719,N_8674);
or U10816 (N_10816,N_7886,N_6504);
and U10817 (N_10817,N_8875,N_7720);
and U10818 (N_10818,N_6409,N_8524);
and U10819 (N_10819,N_8844,N_6922);
xor U10820 (N_10820,N_7131,N_8550);
nand U10821 (N_10821,N_7033,N_6564);
xnor U10822 (N_10822,N_6294,N_6909);
and U10823 (N_10823,N_6588,N_8016);
nand U10824 (N_10824,N_8731,N_8785);
nor U10825 (N_10825,N_8186,N_7945);
nor U10826 (N_10826,N_6950,N_6992);
xnor U10827 (N_10827,N_7874,N_6012);
xor U10828 (N_10828,N_8340,N_8024);
xnor U10829 (N_10829,N_8476,N_6190);
xnor U10830 (N_10830,N_7493,N_7850);
nor U10831 (N_10831,N_8863,N_8908);
or U10832 (N_10832,N_7763,N_6999);
xnor U10833 (N_10833,N_7492,N_8088);
xor U10834 (N_10834,N_6426,N_8648);
and U10835 (N_10835,N_7436,N_7015);
xor U10836 (N_10836,N_8937,N_6415);
xnor U10837 (N_10837,N_6899,N_6078);
nand U10838 (N_10838,N_6706,N_6040);
and U10839 (N_10839,N_7140,N_7015);
or U10840 (N_10840,N_6111,N_7541);
or U10841 (N_10841,N_6715,N_7830);
nand U10842 (N_10842,N_8339,N_7627);
nand U10843 (N_10843,N_8189,N_8881);
xnor U10844 (N_10844,N_7240,N_7859);
nor U10845 (N_10845,N_8857,N_7176);
xnor U10846 (N_10846,N_7564,N_7176);
or U10847 (N_10847,N_7486,N_7497);
xor U10848 (N_10848,N_7336,N_7565);
and U10849 (N_10849,N_6825,N_7404);
or U10850 (N_10850,N_6666,N_8053);
nand U10851 (N_10851,N_7525,N_8914);
nor U10852 (N_10852,N_6671,N_7631);
and U10853 (N_10853,N_7804,N_7509);
xnor U10854 (N_10854,N_7068,N_8518);
xor U10855 (N_10855,N_7082,N_6166);
nand U10856 (N_10856,N_6603,N_6380);
or U10857 (N_10857,N_8140,N_8740);
or U10858 (N_10858,N_8244,N_6342);
nor U10859 (N_10859,N_6141,N_7889);
nor U10860 (N_10860,N_7055,N_6751);
or U10861 (N_10861,N_8930,N_8943);
and U10862 (N_10862,N_6183,N_8371);
nor U10863 (N_10863,N_7722,N_6459);
nand U10864 (N_10864,N_8052,N_6904);
xnor U10865 (N_10865,N_8544,N_8089);
nor U10866 (N_10866,N_7591,N_6049);
nand U10867 (N_10867,N_8336,N_8621);
nand U10868 (N_10868,N_8152,N_7057);
nor U10869 (N_10869,N_7883,N_7137);
nand U10870 (N_10870,N_8976,N_6894);
nand U10871 (N_10871,N_6581,N_7838);
and U10872 (N_10872,N_7498,N_8451);
nand U10873 (N_10873,N_7664,N_6624);
xnor U10874 (N_10874,N_7567,N_6695);
xnor U10875 (N_10875,N_8411,N_8972);
xnor U10876 (N_10876,N_6464,N_6538);
and U10877 (N_10877,N_8995,N_8434);
nor U10878 (N_10878,N_8739,N_8915);
nand U10879 (N_10879,N_7893,N_7648);
or U10880 (N_10880,N_8552,N_6879);
nand U10881 (N_10881,N_8340,N_7544);
nand U10882 (N_10882,N_8685,N_7397);
and U10883 (N_10883,N_8575,N_7731);
xnor U10884 (N_10884,N_8768,N_7647);
xor U10885 (N_10885,N_6289,N_7624);
xor U10886 (N_10886,N_8816,N_8218);
nor U10887 (N_10887,N_7749,N_8106);
nand U10888 (N_10888,N_6043,N_7616);
or U10889 (N_10889,N_7461,N_6410);
xor U10890 (N_10890,N_7821,N_7306);
xnor U10891 (N_10891,N_7325,N_6656);
xor U10892 (N_10892,N_7428,N_7986);
xor U10893 (N_10893,N_8619,N_8745);
and U10894 (N_10894,N_6090,N_6611);
and U10895 (N_10895,N_8490,N_7540);
nor U10896 (N_10896,N_8421,N_8491);
and U10897 (N_10897,N_8409,N_7645);
or U10898 (N_10898,N_8668,N_8255);
xnor U10899 (N_10899,N_8600,N_8547);
nand U10900 (N_10900,N_8534,N_8270);
nand U10901 (N_10901,N_6853,N_7814);
nand U10902 (N_10902,N_8215,N_8923);
and U10903 (N_10903,N_7351,N_8595);
or U10904 (N_10904,N_7142,N_7942);
and U10905 (N_10905,N_6746,N_6376);
nand U10906 (N_10906,N_6396,N_8492);
nand U10907 (N_10907,N_6208,N_6380);
nor U10908 (N_10908,N_8917,N_8730);
and U10909 (N_10909,N_7486,N_8052);
xor U10910 (N_10910,N_7916,N_7400);
and U10911 (N_10911,N_8956,N_6834);
xor U10912 (N_10912,N_8080,N_8514);
nand U10913 (N_10913,N_6789,N_7127);
and U10914 (N_10914,N_8473,N_8975);
or U10915 (N_10915,N_8073,N_6745);
nand U10916 (N_10916,N_7605,N_6046);
or U10917 (N_10917,N_7902,N_7933);
nand U10918 (N_10918,N_6736,N_7155);
and U10919 (N_10919,N_6514,N_7986);
xor U10920 (N_10920,N_7275,N_6243);
nand U10921 (N_10921,N_6138,N_6002);
nand U10922 (N_10922,N_8263,N_8327);
nand U10923 (N_10923,N_6394,N_7889);
nor U10924 (N_10924,N_7758,N_8896);
or U10925 (N_10925,N_7286,N_8283);
nand U10926 (N_10926,N_6703,N_8329);
xor U10927 (N_10927,N_8128,N_6724);
nor U10928 (N_10928,N_7946,N_7575);
xor U10929 (N_10929,N_8474,N_7858);
or U10930 (N_10930,N_8691,N_8336);
or U10931 (N_10931,N_7603,N_7192);
and U10932 (N_10932,N_7774,N_7552);
or U10933 (N_10933,N_8582,N_8549);
and U10934 (N_10934,N_8655,N_6285);
nand U10935 (N_10935,N_8857,N_8025);
nand U10936 (N_10936,N_7962,N_8785);
and U10937 (N_10937,N_8787,N_7452);
nand U10938 (N_10938,N_6436,N_8851);
nand U10939 (N_10939,N_8070,N_8680);
and U10940 (N_10940,N_7495,N_7147);
or U10941 (N_10941,N_6921,N_6233);
xnor U10942 (N_10942,N_8391,N_7587);
nor U10943 (N_10943,N_8137,N_8701);
xnor U10944 (N_10944,N_7258,N_8525);
nor U10945 (N_10945,N_6582,N_7843);
xnor U10946 (N_10946,N_8672,N_8726);
nand U10947 (N_10947,N_6794,N_8955);
and U10948 (N_10948,N_6324,N_7435);
or U10949 (N_10949,N_6258,N_7029);
nor U10950 (N_10950,N_8216,N_6052);
nor U10951 (N_10951,N_8183,N_7932);
nor U10952 (N_10952,N_8240,N_7292);
nand U10953 (N_10953,N_8108,N_7740);
or U10954 (N_10954,N_8983,N_7019);
nor U10955 (N_10955,N_7760,N_7643);
xnor U10956 (N_10956,N_6340,N_6322);
xnor U10957 (N_10957,N_6763,N_8192);
and U10958 (N_10958,N_8711,N_8811);
and U10959 (N_10959,N_6556,N_7660);
nor U10960 (N_10960,N_6396,N_8939);
or U10961 (N_10961,N_8351,N_8750);
or U10962 (N_10962,N_8872,N_7885);
or U10963 (N_10963,N_8752,N_6710);
nand U10964 (N_10964,N_8021,N_6340);
xor U10965 (N_10965,N_8332,N_8347);
and U10966 (N_10966,N_6603,N_6276);
xor U10967 (N_10967,N_6025,N_8637);
or U10968 (N_10968,N_7768,N_6171);
or U10969 (N_10969,N_6303,N_8307);
and U10970 (N_10970,N_8040,N_6659);
nand U10971 (N_10971,N_6651,N_7242);
or U10972 (N_10972,N_7319,N_8977);
xnor U10973 (N_10973,N_8294,N_8750);
nor U10974 (N_10974,N_6037,N_7831);
xor U10975 (N_10975,N_7330,N_8489);
xnor U10976 (N_10976,N_7974,N_7703);
nand U10977 (N_10977,N_7383,N_6789);
nor U10978 (N_10978,N_7445,N_8605);
or U10979 (N_10979,N_6062,N_8237);
xnor U10980 (N_10980,N_8036,N_6499);
and U10981 (N_10981,N_7308,N_7050);
or U10982 (N_10982,N_7131,N_6553);
and U10983 (N_10983,N_6882,N_8222);
nand U10984 (N_10984,N_6080,N_6166);
and U10985 (N_10985,N_7353,N_8137);
and U10986 (N_10986,N_8116,N_6174);
nand U10987 (N_10987,N_6473,N_6893);
nand U10988 (N_10988,N_7809,N_6340);
and U10989 (N_10989,N_7650,N_8365);
nand U10990 (N_10990,N_8503,N_8528);
and U10991 (N_10991,N_7122,N_8617);
nand U10992 (N_10992,N_8902,N_8282);
nor U10993 (N_10993,N_8884,N_7092);
or U10994 (N_10994,N_6977,N_7377);
xor U10995 (N_10995,N_7936,N_8909);
nor U10996 (N_10996,N_8801,N_8199);
nand U10997 (N_10997,N_7420,N_8000);
nor U10998 (N_10998,N_7584,N_8280);
nand U10999 (N_10999,N_7282,N_7196);
nand U11000 (N_11000,N_8462,N_6188);
or U11001 (N_11001,N_6581,N_6129);
or U11002 (N_11002,N_7443,N_7580);
xnor U11003 (N_11003,N_7656,N_7071);
nand U11004 (N_11004,N_6330,N_6876);
or U11005 (N_11005,N_7710,N_8535);
nand U11006 (N_11006,N_8532,N_8172);
and U11007 (N_11007,N_6029,N_8001);
nor U11008 (N_11008,N_8520,N_8571);
xor U11009 (N_11009,N_7526,N_7061);
or U11010 (N_11010,N_7577,N_8593);
nand U11011 (N_11011,N_6755,N_8543);
and U11012 (N_11012,N_6905,N_8324);
nor U11013 (N_11013,N_8245,N_7149);
xor U11014 (N_11014,N_6700,N_8538);
xnor U11015 (N_11015,N_8121,N_8166);
and U11016 (N_11016,N_8935,N_6238);
and U11017 (N_11017,N_8326,N_8038);
and U11018 (N_11018,N_8276,N_7955);
nor U11019 (N_11019,N_6371,N_6180);
xnor U11020 (N_11020,N_8725,N_6492);
xor U11021 (N_11021,N_8032,N_6929);
and U11022 (N_11022,N_8322,N_8070);
nand U11023 (N_11023,N_7205,N_7440);
nand U11024 (N_11024,N_8360,N_8676);
and U11025 (N_11025,N_7636,N_7402);
nor U11026 (N_11026,N_8951,N_6204);
or U11027 (N_11027,N_7712,N_7463);
or U11028 (N_11028,N_6329,N_6557);
xnor U11029 (N_11029,N_8638,N_8390);
nor U11030 (N_11030,N_8595,N_7304);
or U11031 (N_11031,N_6032,N_6293);
nor U11032 (N_11032,N_7713,N_6208);
and U11033 (N_11033,N_6049,N_7117);
and U11034 (N_11034,N_6861,N_7868);
and U11035 (N_11035,N_8360,N_6081);
nand U11036 (N_11036,N_8651,N_8955);
or U11037 (N_11037,N_6374,N_8309);
xor U11038 (N_11038,N_7518,N_8259);
xor U11039 (N_11039,N_7117,N_8261);
nand U11040 (N_11040,N_6122,N_7820);
xnor U11041 (N_11041,N_6844,N_7714);
nor U11042 (N_11042,N_7888,N_6411);
xor U11043 (N_11043,N_8101,N_7944);
or U11044 (N_11044,N_8433,N_7385);
nand U11045 (N_11045,N_6440,N_6659);
xnor U11046 (N_11046,N_7065,N_8022);
or U11047 (N_11047,N_7026,N_7289);
nor U11048 (N_11048,N_8366,N_7719);
or U11049 (N_11049,N_7261,N_7095);
and U11050 (N_11050,N_7865,N_6551);
xnor U11051 (N_11051,N_7557,N_7995);
or U11052 (N_11052,N_7097,N_6259);
nand U11053 (N_11053,N_7413,N_7544);
nor U11054 (N_11054,N_7562,N_7786);
nor U11055 (N_11055,N_8230,N_8103);
nand U11056 (N_11056,N_8229,N_8286);
xor U11057 (N_11057,N_6581,N_6174);
nor U11058 (N_11058,N_7617,N_6936);
and U11059 (N_11059,N_8281,N_7464);
nor U11060 (N_11060,N_6477,N_7798);
nor U11061 (N_11061,N_7783,N_7325);
nor U11062 (N_11062,N_6852,N_6159);
nor U11063 (N_11063,N_8849,N_8662);
nor U11064 (N_11064,N_7033,N_8944);
nand U11065 (N_11065,N_7551,N_7200);
nor U11066 (N_11066,N_8638,N_7842);
and U11067 (N_11067,N_6138,N_7889);
nand U11068 (N_11068,N_6137,N_6572);
nand U11069 (N_11069,N_6842,N_6760);
or U11070 (N_11070,N_7531,N_7573);
xnor U11071 (N_11071,N_7997,N_8249);
xnor U11072 (N_11072,N_6211,N_6142);
nor U11073 (N_11073,N_6591,N_6065);
nand U11074 (N_11074,N_6064,N_8154);
xor U11075 (N_11075,N_8885,N_7064);
nand U11076 (N_11076,N_7621,N_7678);
nand U11077 (N_11077,N_6294,N_7018);
nand U11078 (N_11078,N_7071,N_8714);
and U11079 (N_11079,N_8407,N_8343);
xnor U11080 (N_11080,N_6563,N_6103);
nand U11081 (N_11081,N_8465,N_8798);
nand U11082 (N_11082,N_6818,N_8330);
or U11083 (N_11083,N_7873,N_6041);
xnor U11084 (N_11084,N_7122,N_6241);
nor U11085 (N_11085,N_7191,N_6682);
and U11086 (N_11086,N_7301,N_7060);
nand U11087 (N_11087,N_6254,N_7977);
or U11088 (N_11088,N_8915,N_6026);
and U11089 (N_11089,N_8989,N_8323);
or U11090 (N_11090,N_6893,N_6541);
or U11091 (N_11091,N_8457,N_7886);
nor U11092 (N_11092,N_6957,N_8090);
nor U11093 (N_11093,N_7570,N_8527);
nand U11094 (N_11094,N_8566,N_6796);
xnor U11095 (N_11095,N_7397,N_8727);
nand U11096 (N_11096,N_6697,N_7765);
nor U11097 (N_11097,N_6189,N_6448);
and U11098 (N_11098,N_7906,N_6455);
xor U11099 (N_11099,N_8654,N_8653);
or U11100 (N_11100,N_7887,N_7689);
nor U11101 (N_11101,N_8985,N_8073);
nor U11102 (N_11102,N_6965,N_7606);
and U11103 (N_11103,N_7091,N_7512);
xor U11104 (N_11104,N_7186,N_7740);
nand U11105 (N_11105,N_8641,N_7714);
xor U11106 (N_11106,N_7233,N_6139);
or U11107 (N_11107,N_7368,N_8212);
or U11108 (N_11108,N_8723,N_8857);
or U11109 (N_11109,N_7249,N_7924);
nor U11110 (N_11110,N_7612,N_7379);
xor U11111 (N_11111,N_6659,N_7378);
xor U11112 (N_11112,N_8038,N_8782);
xor U11113 (N_11113,N_6722,N_7035);
nor U11114 (N_11114,N_6041,N_7649);
nor U11115 (N_11115,N_6424,N_6172);
nor U11116 (N_11116,N_6379,N_7342);
nor U11117 (N_11117,N_6959,N_7818);
xnor U11118 (N_11118,N_7715,N_7116);
xor U11119 (N_11119,N_8513,N_8206);
nor U11120 (N_11120,N_6912,N_8426);
xor U11121 (N_11121,N_8611,N_8939);
nand U11122 (N_11122,N_7755,N_7250);
xnor U11123 (N_11123,N_6239,N_6458);
or U11124 (N_11124,N_6594,N_8745);
xor U11125 (N_11125,N_7663,N_7493);
or U11126 (N_11126,N_7096,N_7786);
nor U11127 (N_11127,N_8935,N_8939);
nand U11128 (N_11128,N_7896,N_8844);
and U11129 (N_11129,N_6368,N_6007);
xor U11130 (N_11130,N_7487,N_8718);
and U11131 (N_11131,N_6268,N_8199);
nor U11132 (N_11132,N_8932,N_6737);
nor U11133 (N_11133,N_6935,N_8446);
and U11134 (N_11134,N_8708,N_8423);
xnor U11135 (N_11135,N_8087,N_8768);
nor U11136 (N_11136,N_7538,N_8504);
and U11137 (N_11137,N_7429,N_6145);
nand U11138 (N_11138,N_7610,N_6317);
nor U11139 (N_11139,N_6481,N_8949);
and U11140 (N_11140,N_6140,N_8694);
or U11141 (N_11141,N_6840,N_7834);
and U11142 (N_11142,N_6110,N_7212);
and U11143 (N_11143,N_7182,N_6575);
nor U11144 (N_11144,N_7411,N_8507);
and U11145 (N_11145,N_8119,N_7963);
or U11146 (N_11146,N_7886,N_7058);
nor U11147 (N_11147,N_8375,N_7897);
nand U11148 (N_11148,N_6750,N_7950);
or U11149 (N_11149,N_7733,N_6278);
and U11150 (N_11150,N_7510,N_8879);
xor U11151 (N_11151,N_8905,N_7581);
nand U11152 (N_11152,N_6728,N_8555);
nor U11153 (N_11153,N_8865,N_8222);
nand U11154 (N_11154,N_8456,N_7075);
nor U11155 (N_11155,N_6703,N_6712);
xnor U11156 (N_11156,N_7021,N_7809);
nand U11157 (N_11157,N_7812,N_8035);
or U11158 (N_11158,N_6501,N_7411);
nor U11159 (N_11159,N_6429,N_8629);
nor U11160 (N_11160,N_6952,N_6315);
or U11161 (N_11161,N_6787,N_8872);
or U11162 (N_11162,N_6455,N_6390);
and U11163 (N_11163,N_8285,N_6560);
xor U11164 (N_11164,N_7020,N_7718);
or U11165 (N_11165,N_6687,N_7007);
nand U11166 (N_11166,N_7144,N_6559);
and U11167 (N_11167,N_8846,N_7089);
and U11168 (N_11168,N_6277,N_8995);
nor U11169 (N_11169,N_6751,N_6249);
and U11170 (N_11170,N_8513,N_8394);
xnor U11171 (N_11171,N_6059,N_7769);
nand U11172 (N_11172,N_6259,N_6792);
xor U11173 (N_11173,N_6390,N_7150);
or U11174 (N_11174,N_8691,N_8740);
and U11175 (N_11175,N_6137,N_6844);
and U11176 (N_11176,N_7485,N_7274);
and U11177 (N_11177,N_6861,N_8684);
xor U11178 (N_11178,N_8738,N_8745);
or U11179 (N_11179,N_8450,N_8688);
nor U11180 (N_11180,N_6019,N_6440);
xor U11181 (N_11181,N_8782,N_7323);
or U11182 (N_11182,N_7115,N_7478);
and U11183 (N_11183,N_8624,N_6647);
nand U11184 (N_11184,N_8176,N_7837);
xnor U11185 (N_11185,N_7331,N_8860);
and U11186 (N_11186,N_8059,N_6704);
nand U11187 (N_11187,N_7350,N_8001);
and U11188 (N_11188,N_7393,N_6367);
xnor U11189 (N_11189,N_6851,N_8744);
or U11190 (N_11190,N_7392,N_8610);
xor U11191 (N_11191,N_8977,N_7058);
nand U11192 (N_11192,N_6939,N_8490);
nand U11193 (N_11193,N_8035,N_8365);
and U11194 (N_11194,N_8020,N_8786);
or U11195 (N_11195,N_7134,N_8459);
and U11196 (N_11196,N_8566,N_8316);
nor U11197 (N_11197,N_8794,N_6879);
nand U11198 (N_11198,N_7503,N_6366);
nand U11199 (N_11199,N_8374,N_8840);
nor U11200 (N_11200,N_6209,N_8695);
or U11201 (N_11201,N_8926,N_6651);
xor U11202 (N_11202,N_8840,N_8168);
or U11203 (N_11203,N_7675,N_7331);
nor U11204 (N_11204,N_7797,N_8337);
xor U11205 (N_11205,N_7329,N_6649);
nand U11206 (N_11206,N_6316,N_6810);
and U11207 (N_11207,N_8584,N_8175);
nor U11208 (N_11208,N_6796,N_7392);
xor U11209 (N_11209,N_8941,N_7410);
and U11210 (N_11210,N_6713,N_6109);
and U11211 (N_11211,N_6696,N_8163);
xnor U11212 (N_11212,N_7928,N_7978);
nand U11213 (N_11213,N_8152,N_7812);
nor U11214 (N_11214,N_8098,N_6797);
nor U11215 (N_11215,N_7914,N_7152);
nand U11216 (N_11216,N_8636,N_6162);
xnor U11217 (N_11217,N_6910,N_6017);
nand U11218 (N_11218,N_6697,N_8449);
and U11219 (N_11219,N_8620,N_7626);
nand U11220 (N_11220,N_7004,N_6464);
and U11221 (N_11221,N_6337,N_7942);
and U11222 (N_11222,N_6787,N_8593);
nand U11223 (N_11223,N_7077,N_6733);
nor U11224 (N_11224,N_8713,N_8315);
or U11225 (N_11225,N_8124,N_8800);
nor U11226 (N_11226,N_6290,N_8658);
nand U11227 (N_11227,N_8976,N_7480);
or U11228 (N_11228,N_7980,N_7415);
and U11229 (N_11229,N_7128,N_7985);
nor U11230 (N_11230,N_8049,N_7178);
xnor U11231 (N_11231,N_6492,N_7789);
nand U11232 (N_11232,N_8906,N_8611);
nand U11233 (N_11233,N_7220,N_8441);
nor U11234 (N_11234,N_7778,N_7174);
and U11235 (N_11235,N_6859,N_8072);
or U11236 (N_11236,N_7256,N_7034);
and U11237 (N_11237,N_8860,N_7792);
xor U11238 (N_11238,N_6521,N_8122);
nor U11239 (N_11239,N_6207,N_8316);
or U11240 (N_11240,N_7995,N_6717);
nor U11241 (N_11241,N_7968,N_6576);
xor U11242 (N_11242,N_6970,N_7536);
nor U11243 (N_11243,N_6286,N_6904);
or U11244 (N_11244,N_8454,N_8611);
and U11245 (N_11245,N_6423,N_7917);
nand U11246 (N_11246,N_7855,N_8682);
or U11247 (N_11247,N_6061,N_8184);
or U11248 (N_11248,N_8099,N_7981);
and U11249 (N_11249,N_6809,N_8652);
xnor U11250 (N_11250,N_6624,N_7168);
nor U11251 (N_11251,N_6201,N_8152);
or U11252 (N_11252,N_8178,N_7977);
nor U11253 (N_11253,N_8174,N_6289);
nor U11254 (N_11254,N_8346,N_6964);
or U11255 (N_11255,N_7855,N_8926);
and U11256 (N_11256,N_7818,N_6825);
or U11257 (N_11257,N_7143,N_6927);
and U11258 (N_11258,N_7015,N_6487);
xnor U11259 (N_11259,N_6003,N_8642);
and U11260 (N_11260,N_6503,N_7262);
xor U11261 (N_11261,N_7053,N_6067);
nor U11262 (N_11262,N_7313,N_7105);
nor U11263 (N_11263,N_8353,N_8600);
and U11264 (N_11264,N_7931,N_6194);
nand U11265 (N_11265,N_8654,N_8836);
xor U11266 (N_11266,N_8998,N_7638);
xor U11267 (N_11267,N_8148,N_7069);
xnor U11268 (N_11268,N_8281,N_8235);
nand U11269 (N_11269,N_7569,N_7395);
nor U11270 (N_11270,N_7632,N_7453);
nand U11271 (N_11271,N_8202,N_6307);
and U11272 (N_11272,N_7268,N_7534);
xor U11273 (N_11273,N_8114,N_6015);
nor U11274 (N_11274,N_7307,N_7640);
or U11275 (N_11275,N_8744,N_6249);
or U11276 (N_11276,N_8155,N_6177);
and U11277 (N_11277,N_6504,N_7773);
nor U11278 (N_11278,N_6579,N_7445);
or U11279 (N_11279,N_8963,N_8597);
nor U11280 (N_11280,N_6166,N_7752);
and U11281 (N_11281,N_8887,N_8471);
nand U11282 (N_11282,N_6456,N_6870);
nor U11283 (N_11283,N_8225,N_7988);
xor U11284 (N_11284,N_7564,N_8060);
or U11285 (N_11285,N_8159,N_8373);
and U11286 (N_11286,N_8110,N_6915);
nand U11287 (N_11287,N_7819,N_8650);
nand U11288 (N_11288,N_8938,N_8054);
or U11289 (N_11289,N_8781,N_7722);
nand U11290 (N_11290,N_6717,N_8979);
and U11291 (N_11291,N_7761,N_8654);
and U11292 (N_11292,N_7910,N_7330);
xor U11293 (N_11293,N_6626,N_7224);
xor U11294 (N_11294,N_7672,N_6827);
and U11295 (N_11295,N_6738,N_7121);
xor U11296 (N_11296,N_6139,N_6184);
and U11297 (N_11297,N_6119,N_7892);
xor U11298 (N_11298,N_6334,N_7357);
or U11299 (N_11299,N_8997,N_6739);
nand U11300 (N_11300,N_7956,N_6321);
nor U11301 (N_11301,N_6035,N_6231);
nand U11302 (N_11302,N_8774,N_7388);
xor U11303 (N_11303,N_8475,N_8603);
nor U11304 (N_11304,N_8368,N_6590);
and U11305 (N_11305,N_8664,N_8592);
and U11306 (N_11306,N_8137,N_7801);
and U11307 (N_11307,N_8995,N_8722);
nand U11308 (N_11308,N_8754,N_8556);
and U11309 (N_11309,N_7231,N_7376);
and U11310 (N_11310,N_6712,N_7207);
nor U11311 (N_11311,N_8668,N_8745);
nor U11312 (N_11312,N_8472,N_7197);
or U11313 (N_11313,N_8394,N_7864);
xor U11314 (N_11314,N_6696,N_6219);
nor U11315 (N_11315,N_8122,N_7502);
nand U11316 (N_11316,N_7124,N_6121);
xnor U11317 (N_11317,N_8377,N_7698);
and U11318 (N_11318,N_7377,N_7544);
and U11319 (N_11319,N_7039,N_7151);
nor U11320 (N_11320,N_6964,N_6893);
nor U11321 (N_11321,N_6971,N_6985);
or U11322 (N_11322,N_7417,N_8619);
or U11323 (N_11323,N_8756,N_7797);
or U11324 (N_11324,N_7205,N_7045);
nand U11325 (N_11325,N_7687,N_8501);
nand U11326 (N_11326,N_6971,N_8431);
nand U11327 (N_11327,N_7280,N_7493);
xnor U11328 (N_11328,N_8147,N_7205);
nor U11329 (N_11329,N_6380,N_6249);
and U11330 (N_11330,N_6619,N_8936);
or U11331 (N_11331,N_8190,N_8894);
nor U11332 (N_11332,N_6132,N_7558);
or U11333 (N_11333,N_7977,N_8594);
xnor U11334 (N_11334,N_8526,N_6595);
nand U11335 (N_11335,N_7102,N_6549);
xor U11336 (N_11336,N_8072,N_8654);
and U11337 (N_11337,N_8921,N_8997);
or U11338 (N_11338,N_6629,N_8876);
nor U11339 (N_11339,N_7826,N_6526);
and U11340 (N_11340,N_7250,N_7302);
xor U11341 (N_11341,N_8385,N_6357);
or U11342 (N_11342,N_6322,N_8292);
xnor U11343 (N_11343,N_8352,N_6246);
nand U11344 (N_11344,N_7262,N_7605);
or U11345 (N_11345,N_6409,N_6317);
nand U11346 (N_11346,N_7780,N_7429);
nand U11347 (N_11347,N_6982,N_7698);
xnor U11348 (N_11348,N_7191,N_7972);
nand U11349 (N_11349,N_6340,N_8560);
or U11350 (N_11350,N_8882,N_7701);
and U11351 (N_11351,N_6986,N_8989);
or U11352 (N_11352,N_6805,N_6262);
and U11353 (N_11353,N_8123,N_6123);
nor U11354 (N_11354,N_6827,N_7765);
nand U11355 (N_11355,N_8205,N_7640);
nor U11356 (N_11356,N_8758,N_6840);
and U11357 (N_11357,N_8449,N_8845);
or U11358 (N_11358,N_8209,N_8784);
xnor U11359 (N_11359,N_7430,N_7164);
or U11360 (N_11360,N_8251,N_7632);
nand U11361 (N_11361,N_8499,N_7249);
or U11362 (N_11362,N_7245,N_6101);
xnor U11363 (N_11363,N_6937,N_8464);
or U11364 (N_11364,N_6866,N_7966);
xor U11365 (N_11365,N_8616,N_8483);
nor U11366 (N_11366,N_8511,N_7787);
and U11367 (N_11367,N_6188,N_7912);
and U11368 (N_11368,N_6152,N_6509);
nor U11369 (N_11369,N_6597,N_8949);
nor U11370 (N_11370,N_8237,N_8789);
and U11371 (N_11371,N_7785,N_7644);
nor U11372 (N_11372,N_8769,N_6108);
nand U11373 (N_11373,N_8366,N_6047);
nand U11374 (N_11374,N_6090,N_7210);
xor U11375 (N_11375,N_6289,N_8987);
xor U11376 (N_11376,N_7159,N_8079);
or U11377 (N_11377,N_8582,N_6444);
nand U11378 (N_11378,N_6128,N_6016);
nor U11379 (N_11379,N_7666,N_6337);
nand U11380 (N_11380,N_6929,N_8226);
nor U11381 (N_11381,N_7209,N_8687);
nand U11382 (N_11382,N_8266,N_6230);
or U11383 (N_11383,N_8789,N_8348);
nand U11384 (N_11384,N_8963,N_7396);
nand U11385 (N_11385,N_7479,N_7804);
nor U11386 (N_11386,N_7848,N_7369);
and U11387 (N_11387,N_7860,N_8736);
and U11388 (N_11388,N_7057,N_8227);
or U11389 (N_11389,N_7913,N_7010);
nand U11390 (N_11390,N_7369,N_7405);
nand U11391 (N_11391,N_6179,N_8285);
or U11392 (N_11392,N_7842,N_6422);
nor U11393 (N_11393,N_7004,N_6376);
or U11394 (N_11394,N_8567,N_6109);
xor U11395 (N_11395,N_7376,N_6503);
nand U11396 (N_11396,N_6665,N_8710);
nor U11397 (N_11397,N_6316,N_7245);
and U11398 (N_11398,N_6005,N_6423);
and U11399 (N_11399,N_6267,N_8593);
xnor U11400 (N_11400,N_6660,N_8434);
and U11401 (N_11401,N_7121,N_8256);
and U11402 (N_11402,N_7389,N_8269);
nand U11403 (N_11403,N_6560,N_6096);
nor U11404 (N_11404,N_8881,N_8706);
nor U11405 (N_11405,N_6506,N_8884);
and U11406 (N_11406,N_7812,N_6460);
or U11407 (N_11407,N_6260,N_8859);
or U11408 (N_11408,N_6785,N_6134);
nor U11409 (N_11409,N_6956,N_7084);
and U11410 (N_11410,N_6227,N_7246);
nor U11411 (N_11411,N_6604,N_8439);
or U11412 (N_11412,N_8573,N_6405);
or U11413 (N_11413,N_6258,N_6577);
or U11414 (N_11414,N_7503,N_8597);
nand U11415 (N_11415,N_6602,N_8218);
nor U11416 (N_11416,N_6613,N_7951);
or U11417 (N_11417,N_6213,N_8134);
xor U11418 (N_11418,N_8957,N_6483);
nor U11419 (N_11419,N_7348,N_6137);
nand U11420 (N_11420,N_8097,N_8425);
and U11421 (N_11421,N_8342,N_6462);
or U11422 (N_11422,N_6734,N_7751);
or U11423 (N_11423,N_6912,N_7779);
nand U11424 (N_11424,N_7357,N_6302);
nand U11425 (N_11425,N_7118,N_6260);
or U11426 (N_11426,N_8941,N_8401);
nand U11427 (N_11427,N_6357,N_6701);
nor U11428 (N_11428,N_8923,N_6379);
nor U11429 (N_11429,N_6406,N_7985);
nand U11430 (N_11430,N_7430,N_8260);
nand U11431 (N_11431,N_6714,N_6475);
xnor U11432 (N_11432,N_7485,N_8181);
nand U11433 (N_11433,N_6264,N_8184);
nand U11434 (N_11434,N_8288,N_8506);
xnor U11435 (N_11435,N_6882,N_7621);
nand U11436 (N_11436,N_7288,N_8890);
nand U11437 (N_11437,N_7528,N_6101);
or U11438 (N_11438,N_7109,N_7553);
xnor U11439 (N_11439,N_8516,N_6261);
nor U11440 (N_11440,N_6505,N_7909);
nand U11441 (N_11441,N_6918,N_8814);
xor U11442 (N_11442,N_8414,N_7672);
or U11443 (N_11443,N_6701,N_7076);
nor U11444 (N_11444,N_7900,N_7543);
and U11445 (N_11445,N_7286,N_8672);
or U11446 (N_11446,N_8710,N_6491);
xor U11447 (N_11447,N_7582,N_8828);
or U11448 (N_11448,N_6290,N_7469);
nand U11449 (N_11449,N_8246,N_8182);
xnor U11450 (N_11450,N_8264,N_6852);
nand U11451 (N_11451,N_8472,N_7782);
nand U11452 (N_11452,N_6182,N_8792);
and U11453 (N_11453,N_7692,N_6278);
or U11454 (N_11454,N_6635,N_6752);
nor U11455 (N_11455,N_7465,N_8856);
xor U11456 (N_11456,N_8869,N_7121);
xor U11457 (N_11457,N_7712,N_6100);
and U11458 (N_11458,N_8426,N_6707);
and U11459 (N_11459,N_8410,N_8064);
or U11460 (N_11460,N_8423,N_6115);
nor U11461 (N_11461,N_8628,N_7707);
or U11462 (N_11462,N_6502,N_7397);
nand U11463 (N_11463,N_8675,N_6709);
or U11464 (N_11464,N_6417,N_7639);
and U11465 (N_11465,N_8863,N_7544);
nor U11466 (N_11466,N_7877,N_7304);
nand U11467 (N_11467,N_7970,N_7399);
xor U11468 (N_11468,N_6695,N_8289);
xor U11469 (N_11469,N_7264,N_6595);
and U11470 (N_11470,N_6000,N_6048);
or U11471 (N_11471,N_7494,N_8382);
nand U11472 (N_11472,N_7248,N_8891);
nor U11473 (N_11473,N_7491,N_8856);
or U11474 (N_11474,N_7056,N_7996);
xor U11475 (N_11475,N_7504,N_7685);
and U11476 (N_11476,N_6413,N_8861);
and U11477 (N_11477,N_7895,N_8326);
and U11478 (N_11478,N_7740,N_8482);
nor U11479 (N_11479,N_6405,N_8658);
nor U11480 (N_11480,N_7476,N_7851);
nand U11481 (N_11481,N_6825,N_8794);
xor U11482 (N_11482,N_8198,N_8091);
xnor U11483 (N_11483,N_6351,N_6465);
or U11484 (N_11484,N_8853,N_8539);
or U11485 (N_11485,N_7839,N_6250);
or U11486 (N_11486,N_8668,N_8070);
xor U11487 (N_11487,N_7363,N_6742);
xor U11488 (N_11488,N_6035,N_7433);
and U11489 (N_11489,N_6751,N_7333);
nor U11490 (N_11490,N_8094,N_6037);
nor U11491 (N_11491,N_6682,N_6047);
nor U11492 (N_11492,N_6362,N_6562);
xnor U11493 (N_11493,N_8446,N_7255);
and U11494 (N_11494,N_6290,N_8385);
and U11495 (N_11495,N_8251,N_6055);
and U11496 (N_11496,N_7781,N_7928);
and U11497 (N_11497,N_8481,N_7316);
nor U11498 (N_11498,N_7093,N_7731);
nor U11499 (N_11499,N_8590,N_8257);
and U11500 (N_11500,N_6667,N_6414);
nor U11501 (N_11501,N_7336,N_7799);
nand U11502 (N_11502,N_7513,N_8695);
nor U11503 (N_11503,N_6600,N_6488);
or U11504 (N_11504,N_7363,N_7764);
and U11505 (N_11505,N_7073,N_6021);
xor U11506 (N_11506,N_8007,N_6625);
and U11507 (N_11507,N_7366,N_7112);
and U11508 (N_11508,N_6371,N_7895);
and U11509 (N_11509,N_6395,N_6157);
or U11510 (N_11510,N_7809,N_7864);
xor U11511 (N_11511,N_6914,N_7721);
xnor U11512 (N_11512,N_7247,N_8706);
nand U11513 (N_11513,N_7633,N_7054);
and U11514 (N_11514,N_6813,N_8393);
and U11515 (N_11515,N_7299,N_6603);
nor U11516 (N_11516,N_7028,N_8221);
nand U11517 (N_11517,N_8507,N_8796);
nand U11518 (N_11518,N_8527,N_8596);
nand U11519 (N_11519,N_6733,N_6197);
nor U11520 (N_11520,N_7250,N_7320);
nor U11521 (N_11521,N_6835,N_7749);
nor U11522 (N_11522,N_7042,N_7356);
or U11523 (N_11523,N_8147,N_7886);
nand U11524 (N_11524,N_6310,N_7681);
xor U11525 (N_11525,N_6261,N_8008);
nand U11526 (N_11526,N_7883,N_8716);
nor U11527 (N_11527,N_7284,N_8930);
nand U11528 (N_11528,N_8313,N_8505);
nand U11529 (N_11529,N_7756,N_8363);
xnor U11530 (N_11530,N_8651,N_6533);
nor U11531 (N_11531,N_8646,N_8922);
or U11532 (N_11532,N_6137,N_7937);
nand U11533 (N_11533,N_6434,N_6443);
and U11534 (N_11534,N_8136,N_8501);
xor U11535 (N_11535,N_6673,N_6770);
nor U11536 (N_11536,N_7151,N_8521);
nor U11537 (N_11537,N_6142,N_8914);
xor U11538 (N_11538,N_8660,N_6769);
or U11539 (N_11539,N_7752,N_7548);
xor U11540 (N_11540,N_6527,N_7705);
nand U11541 (N_11541,N_6069,N_8707);
and U11542 (N_11542,N_7940,N_6010);
nand U11543 (N_11543,N_8663,N_7040);
xor U11544 (N_11544,N_8717,N_6688);
or U11545 (N_11545,N_8349,N_8444);
and U11546 (N_11546,N_6423,N_8471);
xor U11547 (N_11547,N_7085,N_6044);
nor U11548 (N_11548,N_6516,N_6569);
or U11549 (N_11549,N_7590,N_8343);
and U11550 (N_11550,N_8789,N_8693);
and U11551 (N_11551,N_6430,N_6079);
nor U11552 (N_11552,N_6876,N_7878);
and U11553 (N_11553,N_8808,N_8337);
xor U11554 (N_11554,N_7663,N_7999);
nor U11555 (N_11555,N_6402,N_7142);
xnor U11556 (N_11556,N_7797,N_6606);
and U11557 (N_11557,N_7753,N_7890);
xor U11558 (N_11558,N_8610,N_7936);
nand U11559 (N_11559,N_7584,N_8837);
or U11560 (N_11560,N_7373,N_6265);
nand U11561 (N_11561,N_6442,N_8081);
xor U11562 (N_11562,N_8663,N_8344);
xor U11563 (N_11563,N_6277,N_6665);
xnor U11564 (N_11564,N_7018,N_7708);
nor U11565 (N_11565,N_7092,N_7685);
or U11566 (N_11566,N_7650,N_6821);
or U11567 (N_11567,N_7812,N_8902);
or U11568 (N_11568,N_7891,N_8336);
nand U11569 (N_11569,N_8879,N_8955);
or U11570 (N_11570,N_8441,N_6893);
nand U11571 (N_11571,N_6478,N_8712);
nor U11572 (N_11572,N_8843,N_7822);
or U11573 (N_11573,N_6959,N_8512);
xor U11574 (N_11574,N_7073,N_7918);
nor U11575 (N_11575,N_6684,N_8530);
or U11576 (N_11576,N_6771,N_8966);
or U11577 (N_11577,N_8187,N_6749);
xnor U11578 (N_11578,N_8574,N_8692);
nand U11579 (N_11579,N_7182,N_7797);
or U11580 (N_11580,N_8415,N_6267);
nand U11581 (N_11581,N_6199,N_8547);
and U11582 (N_11582,N_8422,N_7390);
nand U11583 (N_11583,N_6007,N_7394);
nand U11584 (N_11584,N_6547,N_7473);
xor U11585 (N_11585,N_8621,N_7082);
xnor U11586 (N_11586,N_8061,N_8870);
nand U11587 (N_11587,N_8060,N_8069);
xor U11588 (N_11588,N_7579,N_7754);
xnor U11589 (N_11589,N_7638,N_6211);
xor U11590 (N_11590,N_7691,N_8688);
nor U11591 (N_11591,N_7403,N_8843);
nor U11592 (N_11592,N_8134,N_8017);
nor U11593 (N_11593,N_8884,N_6648);
nor U11594 (N_11594,N_7594,N_7649);
or U11595 (N_11595,N_8670,N_7301);
xor U11596 (N_11596,N_6131,N_8560);
nand U11597 (N_11597,N_8328,N_8929);
nor U11598 (N_11598,N_6864,N_8052);
and U11599 (N_11599,N_8909,N_8595);
xor U11600 (N_11600,N_6730,N_6854);
nor U11601 (N_11601,N_6745,N_7318);
and U11602 (N_11602,N_6811,N_8318);
xnor U11603 (N_11603,N_7595,N_6224);
nand U11604 (N_11604,N_8617,N_8712);
and U11605 (N_11605,N_8858,N_7945);
or U11606 (N_11606,N_7944,N_7482);
nand U11607 (N_11607,N_6940,N_8914);
or U11608 (N_11608,N_6974,N_7325);
and U11609 (N_11609,N_7134,N_8908);
or U11610 (N_11610,N_7018,N_8780);
or U11611 (N_11611,N_8185,N_6492);
nor U11612 (N_11612,N_8030,N_6761);
and U11613 (N_11613,N_6386,N_7687);
and U11614 (N_11614,N_7353,N_8875);
nand U11615 (N_11615,N_7093,N_6430);
nor U11616 (N_11616,N_7466,N_6532);
and U11617 (N_11617,N_6383,N_7971);
nor U11618 (N_11618,N_6397,N_7321);
or U11619 (N_11619,N_6782,N_8696);
or U11620 (N_11620,N_8718,N_8666);
xnor U11621 (N_11621,N_7501,N_7700);
xor U11622 (N_11622,N_7061,N_6981);
and U11623 (N_11623,N_8578,N_7203);
nor U11624 (N_11624,N_7461,N_7793);
nor U11625 (N_11625,N_6268,N_8152);
and U11626 (N_11626,N_7113,N_6286);
nand U11627 (N_11627,N_6021,N_7086);
nand U11628 (N_11628,N_8530,N_8880);
nor U11629 (N_11629,N_8826,N_8796);
xnor U11630 (N_11630,N_7156,N_6898);
or U11631 (N_11631,N_6269,N_8379);
nor U11632 (N_11632,N_8687,N_6095);
and U11633 (N_11633,N_7171,N_7120);
or U11634 (N_11634,N_7900,N_8583);
xor U11635 (N_11635,N_8058,N_6462);
xnor U11636 (N_11636,N_6378,N_7407);
nor U11637 (N_11637,N_8638,N_7791);
nand U11638 (N_11638,N_7692,N_7429);
xnor U11639 (N_11639,N_7999,N_6721);
nand U11640 (N_11640,N_7454,N_7704);
or U11641 (N_11641,N_8273,N_6355);
or U11642 (N_11642,N_7510,N_7826);
and U11643 (N_11643,N_7651,N_6270);
nand U11644 (N_11644,N_6517,N_8566);
and U11645 (N_11645,N_8849,N_7290);
nor U11646 (N_11646,N_8467,N_6201);
nand U11647 (N_11647,N_7018,N_6477);
xor U11648 (N_11648,N_8216,N_6389);
xnor U11649 (N_11649,N_6111,N_7576);
and U11650 (N_11650,N_8395,N_6514);
xnor U11651 (N_11651,N_6716,N_8496);
nand U11652 (N_11652,N_8908,N_8973);
and U11653 (N_11653,N_6588,N_7760);
and U11654 (N_11654,N_6769,N_6280);
nand U11655 (N_11655,N_7315,N_7738);
or U11656 (N_11656,N_6206,N_6623);
and U11657 (N_11657,N_7452,N_8397);
and U11658 (N_11658,N_7001,N_8247);
nand U11659 (N_11659,N_6191,N_6061);
xor U11660 (N_11660,N_7309,N_8119);
xnor U11661 (N_11661,N_8476,N_7965);
or U11662 (N_11662,N_6045,N_8508);
or U11663 (N_11663,N_6126,N_7826);
xnor U11664 (N_11664,N_7200,N_7918);
nor U11665 (N_11665,N_8884,N_7498);
nor U11666 (N_11666,N_8217,N_8085);
and U11667 (N_11667,N_7242,N_6101);
or U11668 (N_11668,N_8235,N_8495);
and U11669 (N_11669,N_6416,N_8016);
and U11670 (N_11670,N_7685,N_6731);
nand U11671 (N_11671,N_6632,N_7490);
xnor U11672 (N_11672,N_7152,N_8934);
and U11673 (N_11673,N_6798,N_7653);
xnor U11674 (N_11674,N_7858,N_6052);
nand U11675 (N_11675,N_8174,N_6555);
xor U11676 (N_11676,N_8688,N_6100);
and U11677 (N_11677,N_7621,N_7155);
nand U11678 (N_11678,N_6799,N_7079);
and U11679 (N_11679,N_8892,N_7479);
nor U11680 (N_11680,N_6517,N_8253);
xor U11681 (N_11681,N_7690,N_7668);
or U11682 (N_11682,N_6664,N_7144);
xor U11683 (N_11683,N_7057,N_6547);
or U11684 (N_11684,N_8898,N_7492);
and U11685 (N_11685,N_6836,N_7546);
nand U11686 (N_11686,N_8452,N_6613);
xor U11687 (N_11687,N_7473,N_7174);
nor U11688 (N_11688,N_6574,N_7980);
xor U11689 (N_11689,N_8901,N_8523);
or U11690 (N_11690,N_8723,N_7710);
and U11691 (N_11691,N_7318,N_8949);
nand U11692 (N_11692,N_6562,N_8489);
nor U11693 (N_11693,N_7773,N_6491);
xnor U11694 (N_11694,N_8156,N_8775);
or U11695 (N_11695,N_8959,N_6859);
nor U11696 (N_11696,N_8596,N_6270);
xnor U11697 (N_11697,N_7439,N_7350);
xnor U11698 (N_11698,N_7120,N_6669);
and U11699 (N_11699,N_8103,N_7692);
nand U11700 (N_11700,N_7683,N_8761);
and U11701 (N_11701,N_7519,N_8172);
and U11702 (N_11702,N_6099,N_8567);
nand U11703 (N_11703,N_7226,N_6891);
nor U11704 (N_11704,N_7949,N_8178);
and U11705 (N_11705,N_6877,N_6152);
xor U11706 (N_11706,N_8141,N_6205);
nand U11707 (N_11707,N_7362,N_6336);
nand U11708 (N_11708,N_7449,N_7909);
xnor U11709 (N_11709,N_6600,N_7160);
and U11710 (N_11710,N_8569,N_6086);
and U11711 (N_11711,N_6357,N_8542);
or U11712 (N_11712,N_6843,N_7504);
nand U11713 (N_11713,N_6230,N_8338);
nor U11714 (N_11714,N_6061,N_6249);
or U11715 (N_11715,N_8275,N_6425);
and U11716 (N_11716,N_7520,N_8611);
xor U11717 (N_11717,N_6770,N_6479);
and U11718 (N_11718,N_7465,N_8499);
or U11719 (N_11719,N_8158,N_8703);
and U11720 (N_11720,N_8215,N_6134);
or U11721 (N_11721,N_8445,N_6259);
or U11722 (N_11722,N_7277,N_7707);
nand U11723 (N_11723,N_8245,N_6755);
and U11724 (N_11724,N_8808,N_7764);
or U11725 (N_11725,N_8108,N_7535);
and U11726 (N_11726,N_6475,N_8975);
and U11727 (N_11727,N_6934,N_6223);
and U11728 (N_11728,N_8846,N_6765);
or U11729 (N_11729,N_8319,N_7748);
or U11730 (N_11730,N_7251,N_6896);
xor U11731 (N_11731,N_6926,N_7323);
and U11732 (N_11732,N_8029,N_8175);
and U11733 (N_11733,N_8245,N_8204);
xor U11734 (N_11734,N_7648,N_7162);
and U11735 (N_11735,N_7889,N_8352);
nor U11736 (N_11736,N_8597,N_6099);
xnor U11737 (N_11737,N_6444,N_6578);
nand U11738 (N_11738,N_7582,N_8920);
nand U11739 (N_11739,N_6893,N_6833);
nor U11740 (N_11740,N_6129,N_8118);
xor U11741 (N_11741,N_7819,N_8908);
or U11742 (N_11742,N_7382,N_7637);
nor U11743 (N_11743,N_8142,N_7061);
or U11744 (N_11744,N_7024,N_6478);
xor U11745 (N_11745,N_6816,N_6774);
or U11746 (N_11746,N_6720,N_8747);
nor U11747 (N_11747,N_7814,N_8344);
nand U11748 (N_11748,N_8758,N_7050);
xnor U11749 (N_11749,N_8807,N_8468);
and U11750 (N_11750,N_8786,N_8709);
nand U11751 (N_11751,N_6289,N_6541);
nand U11752 (N_11752,N_6796,N_8968);
or U11753 (N_11753,N_6533,N_6500);
nor U11754 (N_11754,N_6075,N_6125);
nand U11755 (N_11755,N_7173,N_8972);
xor U11756 (N_11756,N_8591,N_8490);
or U11757 (N_11757,N_6747,N_8131);
nor U11758 (N_11758,N_7142,N_8940);
or U11759 (N_11759,N_8245,N_8839);
or U11760 (N_11760,N_6352,N_8442);
or U11761 (N_11761,N_6506,N_7550);
xor U11762 (N_11762,N_6032,N_6635);
nor U11763 (N_11763,N_8759,N_8699);
or U11764 (N_11764,N_6454,N_6738);
or U11765 (N_11765,N_8230,N_6341);
nor U11766 (N_11766,N_7421,N_7937);
xor U11767 (N_11767,N_7815,N_8583);
xnor U11768 (N_11768,N_6183,N_7318);
nor U11769 (N_11769,N_7193,N_8411);
or U11770 (N_11770,N_7323,N_8064);
or U11771 (N_11771,N_6589,N_7850);
xor U11772 (N_11772,N_6002,N_7897);
and U11773 (N_11773,N_6500,N_8254);
xnor U11774 (N_11774,N_6794,N_8722);
nor U11775 (N_11775,N_6145,N_7814);
nor U11776 (N_11776,N_6055,N_6504);
nor U11777 (N_11777,N_6929,N_7550);
and U11778 (N_11778,N_7758,N_7796);
or U11779 (N_11779,N_6534,N_8158);
nand U11780 (N_11780,N_8578,N_7596);
and U11781 (N_11781,N_8429,N_8451);
or U11782 (N_11782,N_6104,N_7943);
and U11783 (N_11783,N_8660,N_6491);
and U11784 (N_11784,N_7742,N_6492);
and U11785 (N_11785,N_7666,N_8067);
or U11786 (N_11786,N_8924,N_6919);
xnor U11787 (N_11787,N_8022,N_6679);
and U11788 (N_11788,N_8822,N_6050);
or U11789 (N_11789,N_8973,N_7324);
and U11790 (N_11790,N_6091,N_8097);
xor U11791 (N_11791,N_6982,N_8737);
and U11792 (N_11792,N_6525,N_6728);
and U11793 (N_11793,N_8869,N_7469);
nor U11794 (N_11794,N_8783,N_8630);
xor U11795 (N_11795,N_8704,N_8611);
and U11796 (N_11796,N_6313,N_6703);
xor U11797 (N_11797,N_6545,N_6496);
xnor U11798 (N_11798,N_7580,N_8105);
xor U11799 (N_11799,N_6749,N_6984);
or U11800 (N_11800,N_6108,N_8407);
or U11801 (N_11801,N_6878,N_8609);
xor U11802 (N_11802,N_8805,N_8780);
or U11803 (N_11803,N_6105,N_7240);
and U11804 (N_11804,N_8606,N_6893);
or U11805 (N_11805,N_8213,N_8782);
and U11806 (N_11806,N_6601,N_6623);
or U11807 (N_11807,N_6364,N_6372);
nor U11808 (N_11808,N_6829,N_8669);
xnor U11809 (N_11809,N_7616,N_7780);
nor U11810 (N_11810,N_6877,N_8184);
nand U11811 (N_11811,N_6159,N_6435);
or U11812 (N_11812,N_7671,N_8973);
or U11813 (N_11813,N_7633,N_6870);
xnor U11814 (N_11814,N_8995,N_7991);
or U11815 (N_11815,N_6408,N_6476);
nand U11816 (N_11816,N_7878,N_7067);
xor U11817 (N_11817,N_6334,N_6674);
and U11818 (N_11818,N_8255,N_6678);
or U11819 (N_11819,N_8825,N_6293);
nand U11820 (N_11820,N_7993,N_6909);
or U11821 (N_11821,N_7622,N_7593);
xnor U11822 (N_11822,N_8633,N_7765);
xor U11823 (N_11823,N_6309,N_6567);
and U11824 (N_11824,N_8302,N_6564);
nand U11825 (N_11825,N_6651,N_8832);
nand U11826 (N_11826,N_7776,N_6073);
nor U11827 (N_11827,N_6932,N_8354);
nand U11828 (N_11828,N_6549,N_7207);
nor U11829 (N_11829,N_8898,N_7993);
nand U11830 (N_11830,N_6255,N_7116);
and U11831 (N_11831,N_6374,N_6817);
and U11832 (N_11832,N_8504,N_7386);
and U11833 (N_11833,N_6317,N_8678);
or U11834 (N_11834,N_6336,N_7662);
xnor U11835 (N_11835,N_6274,N_6237);
or U11836 (N_11836,N_8328,N_8055);
nor U11837 (N_11837,N_7782,N_8175);
nand U11838 (N_11838,N_7349,N_6560);
nand U11839 (N_11839,N_8855,N_6234);
nor U11840 (N_11840,N_7292,N_6076);
and U11841 (N_11841,N_8279,N_8910);
and U11842 (N_11842,N_7438,N_6004);
or U11843 (N_11843,N_7079,N_6370);
xor U11844 (N_11844,N_8370,N_7795);
xor U11845 (N_11845,N_7321,N_6665);
nor U11846 (N_11846,N_7435,N_8267);
nand U11847 (N_11847,N_7378,N_8299);
nor U11848 (N_11848,N_8785,N_8987);
and U11849 (N_11849,N_7125,N_6175);
nor U11850 (N_11850,N_6018,N_7723);
nand U11851 (N_11851,N_7110,N_7636);
and U11852 (N_11852,N_6811,N_7359);
nand U11853 (N_11853,N_6093,N_7370);
nand U11854 (N_11854,N_7744,N_7675);
or U11855 (N_11855,N_7167,N_7524);
xor U11856 (N_11856,N_6004,N_7717);
and U11857 (N_11857,N_7566,N_7584);
nand U11858 (N_11858,N_8506,N_6337);
and U11859 (N_11859,N_6824,N_7417);
and U11860 (N_11860,N_7100,N_7332);
nand U11861 (N_11861,N_8018,N_6602);
xor U11862 (N_11862,N_8297,N_8497);
nor U11863 (N_11863,N_7453,N_8958);
and U11864 (N_11864,N_8515,N_8666);
or U11865 (N_11865,N_6749,N_6360);
xnor U11866 (N_11866,N_7979,N_6605);
nor U11867 (N_11867,N_7874,N_6802);
or U11868 (N_11868,N_8827,N_6278);
and U11869 (N_11869,N_7790,N_7486);
xor U11870 (N_11870,N_6902,N_6544);
nor U11871 (N_11871,N_6030,N_8396);
or U11872 (N_11872,N_8302,N_8897);
or U11873 (N_11873,N_6623,N_8038);
and U11874 (N_11874,N_7294,N_8006);
nand U11875 (N_11875,N_7353,N_6768);
and U11876 (N_11876,N_6248,N_6733);
nand U11877 (N_11877,N_6069,N_7807);
xor U11878 (N_11878,N_6155,N_6444);
or U11879 (N_11879,N_8732,N_8537);
or U11880 (N_11880,N_6624,N_7533);
nor U11881 (N_11881,N_6652,N_6299);
nor U11882 (N_11882,N_6771,N_8694);
xnor U11883 (N_11883,N_6328,N_7558);
or U11884 (N_11884,N_7279,N_7135);
nor U11885 (N_11885,N_6873,N_6705);
or U11886 (N_11886,N_7918,N_6021);
xor U11887 (N_11887,N_6136,N_8933);
or U11888 (N_11888,N_8087,N_8193);
or U11889 (N_11889,N_6628,N_7517);
nor U11890 (N_11890,N_7975,N_8093);
nand U11891 (N_11891,N_7424,N_6342);
or U11892 (N_11892,N_8036,N_7474);
xor U11893 (N_11893,N_8176,N_8246);
nor U11894 (N_11894,N_6023,N_8513);
nand U11895 (N_11895,N_8813,N_7989);
nor U11896 (N_11896,N_8070,N_7158);
nor U11897 (N_11897,N_6340,N_6850);
nand U11898 (N_11898,N_8898,N_8755);
or U11899 (N_11899,N_7793,N_8724);
nor U11900 (N_11900,N_8895,N_6724);
nor U11901 (N_11901,N_6755,N_6054);
or U11902 (N_11902,N_6894,N_8966);
nand U11903 (N_11903,N_7162,N_8208);
nand U11904 (N_11904,N_7059,N_7417);
xor U11905 (N_11905,N_7651,N_6853);
and U11906 (N_11906,N_6592,N_6207);
nand U11907 (N_11907,N_6169,N_7519);
nand U11908 (N_11908,N_6541,N_7330);
nor U11909 (N_11909,N_7115,N_8058);
nand U11910 (N_11910,N_6007,N_7180);
nand U11911 (N_11911,N_6539,N_7631);
nor U11912 (N_11912,N_8233,N_6210);
or U11913 (N_11913,N_6060,N_8450);
xnor U11914 (N_11914,N_8667,N_8374);
nor U11915 (N_11915,N_7124,N_6686);
nand U11916 (N_11916,N_8984,N_8920);
or U11917 (N_11917,N_6200,N_7450);
nor U11918 (N_11918,N_6264,N_8254);
and U11919 (N_11919,N_7062,N_6819);
and U11920 (N_11920,N_6352,N_7104);
nand U11921 (N_11921,N_6817,N_8620);
nor U11922 (N_11922,N_7148,N_7498);
nor U11923 (N_11923,N_7101,N_8631);
or U11924 (N_11924,N_7288,N_8464);
xor U11925 (N_11925,N_7355,N_8225);
or U11926 (N_11926,N_6108,N_6901);
xor U11927 (N_11927,N_8298,N_7272);
xor U11928 (N_11928,N_7550,N_7396);
and U11929 (N_11929,N_7870,N_7983);
or U11930 (N_11930,N_7841,N_7826);
or U11931 (N_11931,N_6556,N_7177);
or U11932 (N_11932,N_8062,N_7658);
nor U11933 (N_11933,N_7793,N_8293);
nand U11934 (N_11934,N_7031,N_7903);
nor U11935 (N_11935,N_8698,N_6592);
or U11936 (N_11936,N_7116,N_6123);
nor U11937 (N_11937,N_6560,N_8005);
and U11938 (N_11938,N_7324,N_8609);
nand U11939 (N_11939,N_7038,N_7674);
or U11940 (N_11940,N_8144,N_8496);
nor U11941 (N_11941,N_7351,N_6345);
nand U11942 (N_11942,N_8726,N_8067);
or U11943 (N_11943,N_7719,N_7233);
and U11944 (N_11944,N_8484,N_8630);
nor U11945 (N_11945,N_7087,N_8552);
xnor U11946 (N_11946,N_6973,N_6379);
xnor U11947 (N_11947,N_8347,N_8701);
nand U11948 (N_11948,N_6430,N_7371);
nand U11949 (N_11949,N_7411,N_6424);
nand U11950 (N_11950,N_7308,N_6952);
and U11951 (N_11951,N_8760,N_7804);
nor U11952 (N_11952,N_8790,N_7827);
xnor U11953 (N_11953,N_6534,N_7431);
and U11954 (N_11954,N_8505,N_8600);
xor U11955 (N_11955,N_8776,N_7043);
nand U11956 (N_11956,N_6071,N_6930);
nor U11957 (N_11957,N_8291,N_7052);
or U11958 (N_11958,N_7949,N_8601);
nor U11959 (N_11959,N_7650,N_6301);
nand U11960 (N_11960,N_8250,N_7287);
nand U11961 (N_11961,N_8497,N_8800);
xor U11962 (N_11962,N_6408,N_8831);
xnor U11963 (N_11963,N_6743,N_7829);
nor U11964 (N_11964,N_8831,N_8297);
nand U11965 (N_11965,N_6864,N_6562);
and U11966 (N_11966,N_7944,N_6664);
nor U11967 (N_11967,N_6037,N_8437);
nand U11968 (N_11968,N_8861,N_8613);
nor U11969 (N_11969,N_8649,N_7464);
nor U11970 (N_11970,N_7486,N_8371);
nand U11971 (N_11971,N_8933,N_6566);
or U11972 (N_11972,N_8177,N_7154);
or U11973 (N_11973,N_7322,N_8683);
nor U11974 (N_11974,N_6091,N_8954);
or U11975 (N_11975,N_7695,N_8380);
or U11976 (N_11976,N_7558,N_6166);
xnor U11977 (N_11977,N_7957,N_6492);
and U11978 (N_11978,N_6656,N_6349);
nor U11979 (N_11979,N_6650,N_7214);
or U11980 (N_11980,N_8805,N_7675);
nor U11981 (N_11981,N_6544,N_6411);
and U11982 (N_11982,N_7904,N_7525);
or U11983 (N_11983,N_7030,N_7442);
xor U11984 (N_11984,N_8190,N_7221);
xor U11985 (N_11985,N_7732,N_8508);
or U11986 (N_11986,N_8003,N_6766);
nand U11987 (N_11987,N_6339,N_8120);
xor U11988 (N_11988,N_8527,N_8854);
xnor U11989 (N_11989,N_7314,N_7781);
xor U11990 (N_11990,N_7062,N_6807);
xnor U11991 (N_11991,N_8421,N_8338);
nor U11992 (N_11992,N_7819,N_6502);
xnor U11993 (N_11993,N_6062,N_6016);
or U11994 (N_11994,N_6581,N_8710);
and U11995 (N_11995,N_6262,N_7904);
nor U11996 (N_11996,N_8350,N_8546);
or U11997 (N_11997,N_6349,N_7907);
or U11998 (N_11998,N_8068,N_7948);
xnor U11999 (N_11999,N_7532,N_8964);
nand U12000 (N_12000,N_10021,N_10936);
nand U12001 (N_12001,N_10980,N_11193);
or U12002 (N_12002,N_10134,N_10135);
xnor U12003 (N_12003,N_9697,N_9740);
nor U12004 (N_12004,N_11457,N_10436);
or U12005 (N_12005,N_11238,N_11762);
xnor U12006 (N_12006,N_9722,N_11237);
and U12007 (N_12007,N_11089,N_9715);
nand U12008 (N_12008,N_11392,N_10730);
nand U12009 (N_12009,N_9028,N_9467);
xor U12010 (N_12010,N_10507,N_10771);
nor U12011 (N_12011,N_10117,N_10704);
nor U12012 (N_12012,N_11270,N_9294);
or U12013 (N_12013,N_10431,N_11765);
xnor U12014 (N_12014,N_10623,N_10348);
xnor U12015 (N_12015,N_9012,N_9227);
or U12016 (N_12016,N_11408,N_9631);
or U12017 (N_12017,N_11825,N_10752);
xor U12018 (N_12018,N_10801,N_11917);
nor U12019 (N_12019,N_9373,N_9585);
nor U12020 (N_12020,N_10976,N_10778);
or U12021 (N_12021,N_11766,N_9871);
or U12022 (N_12022,N_9531,N_10889);
nand U12023 (N_12023,N_9301,N_9721);
and U12024 (N_12024,N_9070,N_10399);
xnor U12025 (N_12025,N_11062,N_9716);
xnor U12026 (N_12026,N_10747,N_10813);
xor U12027 (N_12027,N_9802,N_10774);
nor U12028 (N_12028,N_10016,N_11714);
nor U12029 (N_12029,N_9753,N_10896);
nor U12030 (N_12030,N_10960,N_10029);
and U12031 (N_12031,N_10834,N_11891);
and U12032 (N_12032,N_9464,N_10259);
nor U12033 (N_12033,N_11326,N_11311);
or U12034 (N_12034,N_9605,N_9989);
or U12035 (N_12035,N_9002,N_9698);
xnor U12036 (N_12036,N_10908,N_9843);
nand U12037 (N_12037,N_9336,N_11470);
or U12038 (N_12038,N_11110,N_9582);
nor U12039 (N_12039,N_11897,N_11654);
or U12040 (N_12040,N_10123,N_9759);
nor U12041 (N_12041,N_10128,N_10068);
xor U12042 (N_12042,N_10072,N_9797);
nor U12043 (N_12043,N_10334,N_11795);
or U12044 (N_12044,N_9306,N_10411);
xor U12045 (N_12045,N_10052,N_11355);
and U12046 (N_12046,N_9577,N_11087);
xor U12047 (N_12047,N_9397,N_10915);
xnor U12048 (N_12048,N_9986,N_9128);
nand U12049 (N_12049,N_9885,N_10626);
nand U12050 (N_12050,N_9654,N_9090);
nand U12051 (N_12051,N_9075,N_11091);
or U12052 (N_12052,N_11636,N_10639);
xnor U12053 (N_12053,N_10200,N_9601);
and U12054 (N_12054,N_11942,N_11977);
xor U12055 (N_12055,N_9785,N_10794);
and U12056 (N_12056,N_9180,N_11582);
xor U12057 (N_12057,N_9170,N_11450);
or U12058 (N_12058,N_10581,N_11444);
or U12059 (N_12059,N_11442,N_10577);
and U12060 (N_12060,N_9096,N_11514);
and U12061 (N_12061,N_10501,N_10167);
nor U12062 (N_12062,N_11082,N_10853);
or U12063 (N_12063,N_11866,N_11386);
or U12064 (N_12064,N_9746,N_9019);
nand U12065 (N_12065,N_10737,N_11836);
xor U12066 (N_12066,N_11902,N_9513);
nor U12067 (N_12067,N_11036,N_10148);
and U12068 (N_12068,N_9253,N_11877);
or U12069 (N_12069,N_11433,N_10755);
xor U12070 (N_12070,N_11466,N_9825);
nor U12071 (N_12071,N_10879,N_10007);
xor U12072 (N_12072,N_11850,N_9223);
and U12073 (N_12073,N_11286,N_11189);
xor U12074 (N_12074,N_11012,N_9938);
and U12075 (N_12075,N_9678,N_9137);
or U12076 (N_12076,N_11979,N_11710);
nand U12077 (N_12077,N_10653,N_9714);
xnor U12078 (N_12078,N_10972,N_11081);
and U12079 (N_12079,N_9472,N_11031);
nor U12080 (N_12080,N_11078,N_11400);
and U12081 (N_12081,N_11840,N_9144);
nand U12082 (N_12082,N_10209,N_11929);
and U12083 (N_12083,N_9265,N_9092);
nor U12084 (N_12084,N_9813,N_11882);
xnor U12085 (N_12085,N_10579,N_9644);
xor U12086 (N_12086,N_9438,N_11673);
or U12087 (N_12087,N_9165,N_10600);
and U12088 (N_12088,N_11161,N_10696);
and U12089 (N_12089,N_10215,N_10783);
nand U12090 (N_12090,N_10337,N_10598);
and U12091 (N_12091,N_9080,N_9973);
and U12092 (N_12092,N_10358,N_10687);
xnor U12093 (N_12093,N_11742,N_10349);
xnor U12094 (N_12094,N_9828,N_11841);
or U12095 (N_12095,N_10086,N_9668);
nand U12096 (N_12096,N_11758,N_10003);
xnor U12097 (N_12097,N_11941,N_10561);
or U12098 (N_12098,N_10257,N_9819);
xor U12099 (N_12099,N_11733,N_9120);
nor U12100 (N_12100,N_10524,N_10784);
xnor U12101 (N_12101,N_9880,N_11528);
nor U12102 (N_12102,N_10112,N_9728);
or U12103 (N_12103,N_11801,N_10920);
or U12104 (N_12104,N_9937,N_9815);
or U12105 (N_12105,N_11340,N_9894);
or U12106 (N_12106,N_11409,N_9095);
or U12107 (N_12107,N_9172,N_11904);
nand U12108 (N_12108,N_10698,N_11013);
xor U12109 (N_12109,N_11190,N_10519);
nor U12110 (N_12110,N_9914,N_9534);
or U12111 (N_12111,N_9786,N_9672);
xnor U12112 (N_12112,N_9752,N_9013);
and U12113 (N_12113,N_11749,N_11506);
nand U12114 (N_12114,N_10062,N_10728);
nor U12115 (N_12115,N_11982,N_9806);
and U12116 (N_12116,N_11324,N_11318);
nor U12117 (N_12117,N_9805,N_9595);
nor U12118 (N_12118,N_11601,N_9287);
and U12119 (N_12119,N_9097,N_9031);
and U12120 (N_12120,N_10320,N_11132);
or U12121 (N_12121,N_11557,N_10186);
or U12122 (N_12122,N_10464,N_9285);
xor U12123 (N_12123,N_10875,N_9270);
or U12124 (N_12124,N_11684,N_10330);
or U12125 (N_12125,N_10506,N_11754);
xnor U12126 (N_12126,N_10239,N_11205);
or U12127 (N_12127,N_11508,N_10212);
or U12128 (N_12128,N_10660,N_11681);
and U12129 (N_12129,N_10489,N_11786);
xor U12130 (N_12130,N_11389,N_9449);
nand U12131 (N_12131,N_11414,N_10253);
nand U12132 (N_12132,N_11056,N_11246);
nand U12133 (N_12133,N_11332,N_11554);
xor U12134 (N_12134,N_11674,N_10846);
xor U12135 (N_12135,N_11724,N_11160);
nand U12136 (N_12136,N_9182,N_9490);
or U12137 (N_12137,N_10077,N_9380);
xnor U12138 (N_12138,N_10088,N_10594);
xnor U12139 (N_12139,N_9311,N_10495);
or U12140 (N_12140,N_10001,N_10825);
nand U12141 (N_12141,N_11652,N_9007);
and U12142 (N_12142,N_10893,N_10140);
or U12143 (N_12143,N_10485,N_9623);
xnor U12144 (N_12144,N_9011,N_9596);
or U12145 (N_12145,N_11080,N_9291);
nand U12146 (N_12146,N_10986,N_9532);
xnor U12147 (N_12147,N_10706,N_9258);
xor U12148 (N_12148,N_9840,N_9361);
nor U12149 (N_12149,N_10869,N_11425);
xor U12150 (N_12150,N_9071,N_10336);
and U12151 (N_12151,N_9857,N_9737);
or U12152 (N_12152,N_9745,N_9948);
or U12153 (N_12153,N_11910,N_11556);
nor U12154 (N_12154,N_9078,N_9168);
xor U12155 (N_12155,N_11021,N_11104);
or U12156 (N_12156,N_11992,N_10708);
nor U12157 (N_12157,N_11806,N_10517);
or U12158 (N_12158,N_9807,N_11284);
and U12159 (N_12159,N_9742,N_11153);
xor U12160 (N_12160,N_11975,N_10447);
or U12161 (N_12161,N_9956,N_11893);
and U12162 (N_12162,N_10012,N_10030);
xnor U12163 (N_12163,N_9845,N_9498);
or U12164 (N_12164,N_10985,N_10913);
xor U12165 (N_12165,N_11655,N_10087);
and U12166 (N_12166,N_9317,N_11876);
nand U12167 (N_12167,N_10493,N_10681);
nand U12168 (N_12168,N_9407,N_9187);
nand U12169 (N_12169,N_11622,N_10081);
or U12170 (N_12170,N_9391,N_11984);
or U12171 (N_12171,N_9116,N_11227);
xnor U12172 (N_12172,N_9437,N_11404);
xnor U12173 (N_12173,N_10291,N_10786);
nand U12174 (N_12174,N_9283,N_11165);
xnor U12175 (N_12175,N_11810,N_10116);
or U12176 (N_12176,N_9591,N_10544);
nand U12177 (N_12177,N_9401,N_9339);
or U12178 (N_12178,N_9670,N_9417);
xor U12179 (N_12179,N_11211,N_11319);
nand U12180 (N_12180,N_10812,N_10703);
nor U12181 (N_12181,N_11073,N_9976);
and U12182 (N_12182,N_11343,N_10545);
or U12183 (N_12183,N_10763,N_9041);
or U12184 (N_12184,N_10480,N_11843);
and U12185 (N_12185,N_11767,N_10810);
nor U12186 (N_12186,N_9503,N_11633);
or U12187 (N_12187,N_9156,N_11236);
or U12188 (N_12188,N_9827,N_11463);
and U12189 (N_12189,N_9733,N_9206);
xor U12190 (N_12190,N_9318,N_11625);
nand U12191 (N_12191,N_10572,N_9225);
or U12192 (N_12192,N_10638,N_9302);
nand U12193 (N_12193,N_11239,N_11581);
nand U12194 (N_12194,N_10322,N_11264);
nand U12195 (N_12195,N_11271,N_11471);
and U12196 (N_12196,N_11320,N_11456);
xnor U12197 (N_12197,N_11464,N_10731);
xor U12198 (N_12198,N_10033,N_9549);
or U12199 (N_12199,N_9719,N_10028);
nand U12200 (N_12200,N_11645,N_9916);
xor U12201 (N_12201,N_11844,N_9789);
or U12202 (N_12202,N_10292,N_10234);
nand U12203 (N_12203,N_10839,N_9942);
and U12204 (N_12204,N_10655,N_9014);
and U12205 (N_12205,N_10611,N_11865);
and U12206 (N_12206,N_11587,N_9922);
nor U12207 (N_12207,N_10452,N_9061);
or U12208 (N_12208,N_9264,N_10843);
xor U12209 (N_12209,N_11148,N_9091);
xnor U12210 (N_12210,N_11222,N_11546);
and U12211 (N_12211,N_9276,N_11138);
nand U12212 (N_12212,N_9627,N_10175);
or U12213 (N_12213,N_9088,N_11930);
and U12214 (N_12214,N_10329,N_9705);
xnor U12215 (N_12215,N_11512,N_11493);
nand U12216 (N_12216,N_10923,N_11640);
or U12217 (N_12217,N_11194,N_10300);
nand U12218 (N_12218,N_10232,N_9675);
nor U12219 (N_12219,N_9502,N_11668);
or U12220 (N_12220,N_11487,N_11621);
nor U12221 (N_12221,N_9163,N_10897);
nand U12222 (N_12222,N_10224,N_11075);
nor U12223 (N_12223,N_9680,N_9215);
nor U12224 (N_12224,N_11993,N_9337);
and U12225 (N_12225,N_9148,N_10251);
nand U12226 (N_12226,N_10629,N_11229);
nand U12227 (N_12227,N_10083,N_10136);
xnor U12228 (N_12228,N_11037,N_11356);
or U12229 (N_12229,N_10105,N_9383);
xnor U12230 (N_12230,N_11751,N_11994);
or U12231 (N_12231,N_11159,N_11517);
and U12232 (N_12232,N_11925,N_9844);
nand U12233 (N_12233,N_9693,N_10888);
nor U12234 (N_12234,N_10158,N_11116);
nor U12235 (N_12235,N_9134,N_9882);
or U12236 (N_12236,N_9546,N_11792);
xor U12237 (N_12237,N_11443,N_9257);
and U12238 (N_12238,N_11880,N_11798);
nor U12239 (N_12239,N_9114,N_11120);
nand U12240 (N_12240,N_10060,N_11720);
xor U12241 (N_12241,N_11774,N_11848);
nor U12242 (N_12242,N_11963,N_11396);
nand U12243 (N_12243,N_11538,N_9691);
or U12244 (N_12244,N_10332,N_10034);
xor U12245 (N_12245,N_9418,N_10591);
xor U12246 (N_12246,N_9848,N_10394);
and U12247 (N_12247,N_10020,N_11378);
nor U12248 (N_12248,N_9760,N_11357);
and U12249 (N_12249,N_10546,N_10475);
or U12250 (N_12250,N_11564,N_9436);
and U12251 (N_12251,N_9608,N_10126);
nand U12252 (N_12252,N_11136,N_10548);
nor U12253 (N_12253,N_10098,N_11813);
and U12254 (N_12254,N_11938,N_10351);
xnor U12255 (N_12255,N_10631,N_11417);
xor U12256 (N_12256,N_10570,N_10926);
nor U12257 (N_12257,N_9125,N_11723);
nor U12258 (N_12258,N_9996,N_10018);
and U12259 (N_12259,N_10650,N_9330);
xor U12260 (N_12260,N_10002,N_10726);
or U12261 (N_12261,N_11743,N_9564);
nor U12262 (N_12262,N_9739,N_10019);
and U12263 (N_12263,N_11288,N_10318);
nand U12264 (N_12264,N_11192,N_11359);
or U12265 (N_12265,N_10230,N_11651);
nor U12266 (N_12266,N_9385,N_11352);
and U12267 (N_12267,N_9933,N_10804);
nand U12268 (N_12268,N_10191,N_9776);
and U12269 (N_12269,N_11609,N_10701);
nor U12270 (N_12270,N_9348,N_11691);
and U12271 (N_12271,N_11516,N_10335);
nor U12272 (N_12272,N_11446,N_9669);
and U12273 (N_12273,N_9485,N_9695);
nand U12274 (N_12274,N_10961,N_10789);
or U12275 (N_12275,N_11331,N_9247);
or U12276 (N_12276,N_11947,N_9350);
and U12277 (N_12277,N_11029,N_11928);
and U12278 (N_12278,N_10798,N_11501);
and U12279 (N_12279,N_11971,N_10724);
xor U12280 (N_12280,N_9833,N_10564);
nand U12281 (N_12281,N_9602,N_11883);
nand U12282 (N_12282,N_10011,N_11044);
nand U12283 (N_12283,N_10366,N_11335);
and U12284 (N_12284,N_11111,N_9780);
or U12285 (N_12285,N_9646,N_11643);
and U12286 (N_12286,N_9779,N_10067);
nand U12287 (N_12287,N_10064,N_11033);
and U12288 (N_12288,N_9661,N_11230);
nand U12289 (N_12289,N_9934,N_11093);
nor U12290 (N_12290,N_11195,N_10993);
or U12291 (N_12291,N_11669,N_10766);
and U12292 (N_12292,N_10910,N_9682);
nand U12293 (N_12293,N_10237,N_10427);
or U12294 (N_12294,N_9851,N_9015);
nand U12295 (N_12295,N_11771,N_10822);
or U12296 (N_12296,N_11641,N_10848);
and U12297 (N_12297,N_10610,N_11753);
nand U12298 (N_12298,N_11095,N_10947);
nor U12299 (N_12299,N_11967,N_11346);
nor U12300 (N_12300,N_11421,N_9685);
and U12301 (N_12301,N_11043,N_11265);
nor U12302 (N_12302,N_10401,N_10829);
nand U12303 (N_12303,N_9100,N_9769);
nor U12304 (N_12304,N_10663,N_11807);
nand U12305 (N_12305,N_9958,N_10599);
xor U12306 (N_12306,N_10159,N_9947);
xnor U12307 (N_12307,N_10521,N_9898);
and U12308 (N_12308,N_10576,N_9205);
nand U12309 (N_12309,N_10114,N_10141);
nor U12310 (N_12310,N_10757,N_9523);
nand U12311 (N_12311,N_9507,N_10015);
xnor U12312 (N_12312,N_9526,N_11853);
or U12313 (N_12313,N_9190,N_11174);
and U12314 (N_12314,N_10602,N_9950);
xnor U12315 (N_12315,N_9312,N_11997);
or U12316 (N_12316,N_9069,N_10362);
xnor U12317 (N_12317,N_11732,N_9694);
nand U12318 (N_12318,N_11495,N_11634);
and U12319 (N_12319,N_11816,N_11115);
nand U12320 (N_12320,N_11112,N_9706);
nor U12321 (N_12321,N_11234,N_9588);
nand U12322 (N_12322,N_9370,N_9539);
nand U12323 (N_12323,N_10145,N_11197);
nor U12324 (N_12324,N_11933,N_10635);
xor U12325 (N_12325,N_9451,N_9266);
xnor U12326 (N_12326,N_10963,N_10743);
nand U12327 (N_12327,N_10202,N_9943);
nor U12328 (N_12328,N_9701,N_11822);
or U12329 (N_12329,N_10421,N_9505);
nand U12330 (N_12330,N_11348,N_9838);
nor U12331 (N_12331,N_9511,N_10571);
nor U12332 (N_12332,N_11272,N_11418);
or U12333 (N_12333,N_10227,N_9518);
xnor U12334 (N_12334,N_9619,N_11468);
xnor U12335 (N_12335,N_10860,N_9463);
and U12336 (N_12336,N_9560,N_11410);
or U12337 (N_12337,N_10343,N_11076);
and U12338 (N_12338,N_11533,N_9858);
xor U12339 (N_12339,N_11305,N_11750);
nand U12340 (N_12340,N_10820,N_10575);
nor U12341 (N_12341,N_10453,N_11868);
nor U12342 (N_12342,N_9852,N_11047);
xnor U12343 (N_12343,N_9246,N_10551);
and U12344 (N_12344,N_9025,N_11618);
nand U12345 (N_12345,N_11679,N_10612);
and U12346 (N_12346,N_9089,N_10680);
nor U12347 (N_12347,N_10405,N_9136);
nand U12348 (N_12348,N_11066,N_11793);
nor U12349 (N_12349,N_11591,N_9001);
xnor U12350 (N_12350,N_11274,N_10628);
nor U12351 (N_12351,N_10950,N_11469);
nor U12352 (N_12352,N_10206,N_9583);
or U12353 (N_12353,N_9626,N_11596);
nor U12354 (N_12354,N_11858,N_10844);
or U12355 (N_12355,N_10404,N_10768);
nand U12356 (N_12356,N_9191,N_9349);
and U12357 (N_12357,N_10945,N_9030);
or U12358 (N_12358,N_10074,N_10616);
and U12359 (N_12359,N_10473,N_11181);
or U12360 (N_12360,N_9913,N_11358);
xor U12361 (N_12361,N_9024,N_10125);
and U12362 (N_12362,N_11861,N_9643);
and U12363 (N_12363,N_9847,N_9791);
xnor U12364 (N_12364,N_10270,N_11981);
or U12365 (N_12365,N_9767,N_9677);
xnor U12366 (N_12366,N_11524,N_11188);
and U12367 (N_12367,N_9204,N_11064);
or U12368 (N_12368,N_10759,N_10023);
or U12369 (N_12369,N_11615,N_10168);
or U12370 (N_12370,N_10876,N_11809);
or U12371 (N_12371,N_11692,N_9964);
nor U12372 (N_12372,N_10694,N_10949);
xnor U12373 (N_12373,N_9261,N_10688);
nor U12374 (N_12374,N_10723,N_9495);
and U12375 (N_12375,N_11086,N_10177);
or U12376 (N_12376,N_10921,N_9709);
and U12377 (N_12377,N_10739,N_11162);
and U12378 (N_12378,N_9084,N_10668);
nor U12379 (N_12379,N_11206,N_9320);
nor U12380 (N_12380,N_9907,N_9936);
nor U12381 (N_12381,N_11656,N_9198);
or U12382 (N_12382,N_11527,N_10373);
nor U12383 (N_12383,N_9712,N_10981);
nand U12384 (N_12384,N_9782,N_10805);
or U12385 (N_12385,N_10199,N_11040);
xnor U12386 (N_12386,N_10966,N_10043);
or U12387 (N_12387,N_11828,N_11778);
nand U12388 (N_12388,N_10090,N_11350);
nand U12389 (N_12389,N_9057,N_11867);
and U12390 (N_12390,N_11398,N_11739);
xor U12391 (N_12391,N_10832,N_10264);
or U12392 (N_12392,N_10652,N_9130);
nand U12393 (N_12393,N_11143,N_10323);
and U12394 (N_12394,N_11048,N_11505);
or U12395 (N_12395,N_10396,N_11913);
and U12396 (N_12396,N_10118,N_11452);
nor U12397 (N_12397,N_9667,N_9101);
nand U12398 (N_12398,N_10111,N_10543);
or U12399 (N_12399,N_10375,N_10455);
nor U12400 (N_12400,N_11577,N_9972);
and U12401 (N_12401,N_10483,N_9296);
xor U12402 (N_12402,N_9260,N_11662);
or U12403 (N_12403,N_10710,N_11127);
and U12404 (N_12404,N_10228,N_10536);
nor U12405 (N_12405,N_9085,N_9876);
and U12406 (N_12406,N_11440,N_11122);
and U12407 (N_12407,N_11004,N_10540);
nand U12408 (N_12408,N_10356,N_9192);
or U12409 (N_12409,N_11612,N_11509);
xor U12410 (N_12410,N_11874,N_11385);
or U12411 (N_12411,N_10818,N_10044);
or U12412 (N_12412,N_9957,N_11819);
or U12413 (N_12413,N_11650,N_10496);
or U12414 (N_12414,N_9365,N_9637);
nand U12415 (N_12415,N_11360,N_11183);
or U12416 (N_12416,N_9375,N_10925);
and U12417 (N_12417,N_11413,N_10533);
nand U12418 (N_12418,N_11199,N_11383);
and U12419 (N_12419,N_11247,N_10780);
nand U12420 (N_12420,N_10243,N_10578);
xnor U12421 (N_12421,N_11336,N_11071);
nand U12422 (N_12422,N_10390,N_10155);
nand U12423 (N_12423,N_11368,N_10513);
and U12424 (N_12424,N_11186,N_9930);
xnor U12425 (N_12425,N_10718,N_9338);
nand U12426 (N_12426,N_9820,N_9704);
xnor U12427 (N_12427,N_11329,N_11321);
nand U12428 (N_12428,N_9951,N_10425);
nor U12429 (N_12429,N_10894,N_9792);
or U12430 (N_12430,N_11182,N_11627);
nor U12431 (N_12431,N_10903,N_10223);
and U12432 (N_12432,N_9652,N_10659);
and U12433 (N_12433,N_10370,N_10213);
nand U12434 (N_12434,N_9650,N_10194);
nor U12435 (N_12435,N_11969,N_11569);
or U12436 (N_12436,N_9974,N_9415);
nor U12437 (N_12437,N_10583,N_11965);
nand U12438 (N_12438,N_11057,N_9919);
nor U12439 (N_12439,N_10817,N_11576);
or U12440 (N_12440,N_10933,N_11939);
xnor U12441 (N_12441,N_9980,N_9049);
or U12442 (N_12442,N_11688,N_10107);
or U12443 (N_12443,N_10120,N_9141);
and U12444 (N_12444,N_10313,N_10625);
xnor U12445 (N_12445,N_10661,N_9272);
or U12446 (N_12446,N_9881,N_11559);
nor U12447 (N_12447,N_10153,N_11130);
nor U12448 (N_12448,N_11846,N_11046);
nand U12449 (N_12449,N_9911,N_11500);
and U12450 (N_12450,N_10745,N_11697);
or U12451 (N_12451,N_11026,N_9457);
nor U12452 (N_12452,N_9896,N_9662);
nor U12453 (N_12453,N_9404,N_10384);
nand U12454 (N_12454,N_10646,N_10870);
and U12455 (N_12455,N_9887,N_10727);
and U12456 (N_12456,N_11394,N_11515);
or U12457 (N_12457,N_9064,N_9371);
nand U12458 (N_12458,N_10437,N_9132);
and U12459 (N_12459,N_11313,N_11568);
and U12460 (N_12460,N_10884,N_10308);
or U12461 (N_12461,N_9409,N_10285);
or U12462 (N_12462,N_10665,N_10382);
nand U12463 (N_12463,N_11455,N_10053);
or U12464 (N_12464,N_10998,N_10103);
nand U12465 (N_12465,N_10361,N_9750);
or U12466 (N_12466,N_9432,N_9673);
nand U12467 (N_12467,N_9770,N_11873);
or U12468 (N_12468,N_11032,N_11756);
and U12469 (N_12469,N_10826,N_9459);
or U12470 (N_12470,N_9026,N_9105);
or U12471 (N_12471,N_9658,N_10025);
nor U12472 (N_12472,N_9445,N_11261);
nor U12473 (N_12473,N_11334,N_10809);
nand U12474 (N_12474,N_10150,N_10605);
nand U12475 (N_12475,N_10272,N_9452);
xor U12476 (N_12476,N_9181,N_9803);
nor U12477 (N_12477,N_10410,N_9629);
nand U12478 (N_12478,N_11291,N_9736);
and U12479 (N_12479,N_9441,N_9022);
and U12480 (N_12480,N_11241,N_11834);
and U12481 (N_12481,N_11805,N_9959);
or U12482 (N_12482,N_11536,N_10250);
and U12483 (N_12483,N_10099,N_10642);
nand U12484 (N_12484,N_10836,N_9081);
nand U12485 (N_12485,N_9965,N_11168);
xnor U12486 (N_12486,N_11716,N_9506);
nand U12487 (N_12487,N_11968,N_9902);
nor U12488 (N_12488,N_11972,N_9717);
xor U12489 (N_12489,N_11263,N_9488);
nand U12490 (N_12490,N_9589,N_9476);
or U12491 (N_12491,N_9173,N_10038);
nor U12492 (N_12492,N_10248,N_9656);
and U12493 (N_12493,N_11072,N_9633);
xor U12494 (N_12494,N_11233,N_10440);
nand U12495 (N_12495,N_9139,N_9590);
xnor U12496 (N_12496,N_9448,N_10262);
or U12497 (N_12497,N_9891,N_10271);
xor U12498 (N_12498,N_9045,N_11363);
and U12499 (N_12499,N_11737,N_11889);
xnor U12500 (N_12500,N_10758,N_10807);
nor U12501 (N_12501,N_9413,N_10733);
and U12502 (N_12502,N_10208,N_9376);
xnor U12503 (N_12503,N_11049,N_9119);
and U12504 (N_12504,N_11025,N_11314);
and U12505 (N_12505,N_10664,N_10917);
nor U12506 (N_12506,N_10235,N_9360);
nand U12507 (N_12507,N_11124,N_10890);
or U12508 (N_12508,N_11472,N_9671);
nor U12509 (N_12509,N_11718,N_11594);
or U12510 (N_12510,N_11451,N_11502);
or U12511 (N_12511,N_9328,N_11776);
and U12512 (N_12512,N_10838,N_11520);
nand U12513 (N_12513,N_9058,N_9932);
nand U12514 (N_12514,N_9524,N_9610);
xnor U12515 (N_12515,N_11058,N_10218);
xor U12516 (N_12516,N_10472,N_10039);
or U12517 (N_12517,N_9681,N_9278);
and U12518 (N_12518,N_11966,N_11478);
nand U12519 (N_12519,N_11906,N_10845);
xor U12520 (N_12520,N_11054,N_9632);
or U12521 (N_12521,N_11098,N_9405);
nand U12522 (N_12522,N_10907,N_9234);
nor U12523 (N_12523,N_10641,N_9235);
or U12524 (N_12524,N_10924,N_9928);
and U12525 (N_12525,N_10584,N_11403);
and U12526 (N_12526,N_10449,N_10984);
or U12527 (N_12527,N_9411,N_9179);
and U12528 (N_12528,N_11173,N_10788);
nor U12529 (N_12529,N_10299,N_9649);
xnor U12530 (N_12530,N_9766,N_9905);
and U12531 (N_12531,N_11106,N_11172);
xnor U12532 (N_12532,N_10061,N_11084);
nor U12533 (N_12533,N_9940,N_9453);
nand U12534 (N_12534,N_10909,N_9293);
nand U12535 (N_12535,N_11202,N_11099);
xnor U12536 (N_12536,N_11781,N_11665);
and U12537 (N_12537,N_9434,N_11842);
nor U12538 (N_12538,N_9479,N_11550);
nor U12539 (N_12539,N_11983,N_9798);
nor U12540 (N_12540,N_10971,N_10964);
nor U12541 (N_12541,N_11391,N_9810);
nor U12542 (N_12542,N_10415,N_10070);
nor U12543 (N_12543,N_9889,N_10672);
xnor U12544 (N_12544,N_11580,N_9018);
nor U12545 (N_12545,N_10877,N_11296);
nand U12546 (N_12546,N_9177,N_11510);
and U12547 (N_12547,N_11590,N_10138);
nor U12548 (N_12548,N_10066,N_10514);
or U12549 (N_12549,N_9612,N_10245);
and U12550 (N_12550,N_10014,N_9423);
or U12551 (N_12551,N_11375,N_11815);
and U12552 (N_12552,N_11624,N_9210);
nand U12553 (N_12553,N_10376,N_11915);
or U12554 (N_12554,N_11257,N_11584);
nand U12555 (N_12555,N_9273,N_10619);
xnor U12556 (N_12556,N_10770,N_11273);
or U12557 (N_12557,N_9254,N_11845);
or U12558 (N_12558,N_10937,N_9581);
nand U12559 (N_12559,N_10071,N_11905);
xor U12560 (N_12560,N_9545,N_10402);
nor U12561 (N_12561,N_11126,N_10263);
or U12562 (N_12562,N_11214,N_9399);
or U12563 (N_12563,N_10327,N_9628);
xnor U12564 (N_12564,N_10049,N_11921);
xor U12565 (N_12565,N_11006,N_10857);
or U12566 (N_12566,N_11773,N_9222);
or U12567 (N_12567,N_10381,N_11277);
nor U12568 (N_12568,N_11817,N_11337);
nor U12569 (N_12569,N_10442,N_11731);
and U12570 (N_12570,N_9651,N_11041);
nand U12571 (N_12571,N_10772,N_10955);
nand U12572 (N_12572,N_11626,N_10231);
and U12573 (N_12573,N_9150,N_9968);
or U12574 (N_12574,N_9072,N_10725);
and U12575 (N_12575,N_10719,N_10942);
and U12576 (N_12576,N_11871,N_10046);
nand U12577 (N_12577,N_10613,N_10595);
nand U12578 (N_12578,N_10482,N_10531);
nand U12579 (N_12579,N_9006,N_11644);
xnor U12580 (N_12580,N_9931,N_11235);
nand U12581 (N_12581,N_10782,N_11196);
or U12582 (N_12582,N_10360,N_9250);
or U12583 (N_12583,N_10439,N_10525);
xnor U12584 (N_12584,N_9991,N_11678);
nand U12585 (N_12585,N_11281,N_9474);
nand U12586 (N_12586,N_9865,N_11571);
nor U12587 (N_12587,N_11872,N_9720);
and U12588 (N_12588,N_9242,N_9086);
nor U12589 (N_12589,N_11243,N_10448);
xnor U12590 (N_12590,N_11606,N_11912);
nor U12591 (N_12591,N_11477,N_10851);
xnor U12592 (N_12592,N_9038,N_9363);
nand U12593 (N_12593,N_9599,N_10471);
nor U12594 (N_12594,N_11849,N_10684);
nand U12595 (N_12595,N_9550,N_9334);
nor U12596 (N_12596,N_10428,N_10643);
nor U12597 (N_12597,N_9846,N_9307);
nand U12598 (N_12598,N_10147,N_11705);
xor U12599 (N_12599,N_11342,N_11035);
or U12600 (N_12600,N_10741,N_11610);
nand U12601 (N_12601,N_9473,N_10333);
nand U12602 (N_12602,N_10487,N_11831);
nand U12603 (N_12603,N_10065,N_10562);
nor U12604 (N_12604,N_11632,N_9855);
nor U12605 (N_12605,N_9489,N_10386);
or U12606 (N_12606,N_9103,N_11974);
or U12607 (N_12607,N_11447,N_10657);
nor U12608 (N_12608,N_11927,N_10567);
nor U12609 (N_12609,N_11371,N_9184);
or U12610 (N_12610,N_9431,N_9984);
and U12611 (N_12611,N_11407,N_9877);
nor U12612 (N_12612,N_10918,N_10863);
nor U12613 (N_12613,N_10697,N_11646);
nor U12614 (N_12614,N_11002,N_9226);
or U12615 (N_12615,N_9738,N_10178);
nor U12616 (N_12616,N_10144,N_9176);
xor U12617 (N_12617,N_9941,N_10523);
nand U12618 (N_12618,N_9189,N_10840);
nor U12619 (N_12619,N_10604,N_9175);
and U12620 (N_12620,N_11395,N_9239);
and U12621 (N_12621,N_9744,N_9381);
nand U12622 (N_12622,N_10035,N_9939);
or U12623 (N_12623,N_9332,N_11830);
nand U12624 (N_12624,N_10522,N_9726);
and U12625 (N_12625,N_10873,N_9113);
and U12626 (N_12626,N_11207,N_10340);
xnor U12627 (N_12627,N_10849,N_9850);
nand U12628 (N_12628,N_11962,N_9461);
nor U12629 (N_12629,N_11764,N_10944);
nor U12630 (N_12630,N_9430,N_11299);
and U12631 (N_12631,N_10978,N_10406);
nand U12632 (N_12632,N_9945,N_10497);
xnor U12633 (N_12633,N_10282,N_11519);
and U12634 (N_12634,N_9040,N_10904);
nand U12635 (N_12635,N_10097,N_10886);
or U12636 (N_12636,N_9112,N_11886);
nor U12637 (N_12637,N_11154,N_9558);
nand U12638 (N_12638,N_9009,N_10310);
or U12639 (N_12639,N_9603,N_10342);
xor U12640 (N_12640,N_10510,N_10553);
xor U12641 (N_12641,N_10586,N_11824);
or U12642 (N_12642,N_11123,N_10319);
xor U12643 (N_12643,N_10236,N_9893);
nor U12644 (N_12644,N_10720,N_10180);
and U12645 (N_12645,N_10420,N_11973);
nand U12646 (N_12646,N_10968,N_11998);
nand U12647 (N_12647,N_11734,N_11995);
nor U12648 (N_12648,N_9108,N_11061);
or U12649 (N_12649,N_10520,N_10547);
nand U12650 (N_12650,N_10750,N_11525);
nor U12651 (N_12651,N_9224,N_10566);
xor U12652 (N_12652,N_9369,N_10858);
nor U12653 (N_12653,N_10899,N_10871);
or U12654 (N_12654,N_9926,N_11693);
and U12655 (N_12655,N_11366,N_9010);
nand U12656 (N_12656,N_10791,N_9429);
xor U12657 (N_12657,N_10528,N_11957);
or U12658 (N_12658,N_11715,N_11338);
nor U12659 (N_12659,N_9978,N_11940);
or U12660 (N_12660,N_9895,N_10988);
nor U12661 (N_12661,N_9286,N_10005);
nand U12662 (N_12662,N_11784,N_9949);
and U12663 (N_12663,N_9079,N_9483);
nor U12664 (N_12664,N_10769,N_9842);
nand U12665 (N_12665,N_10093,N_9985);
and U12666 (N_12666,N_9878,N_11647);
nor U12667 (N_12667,N_9625,N_9077);
or U12668 (N_12668,N_11381,N_10991);
nand U12669 (N_12669,N_11768,N_9830);
xor U12670 (N_12670,N_11294,N_9703);
xnor U12671 (N_12671,N_10713,N_10537);
nand U12672 (N_12672,N_11266,N_11899);
xnor U12673 (N_12673,N_9207,N_11245);
or U12674 (N_12674,N_9297,N_10363);
and U12675 (N_12675,N_9525,N_10106);
nor U12676 (N_12676,N_10256,N_9519);
or U12677 (N_12677,N_10722,N_11016);
and U12678 (N_12678,N_10042,N_10582);
xnor U12679 (N_12679,N_9347,N_11490);
nor U12680 (N_12680,N_10563,N_10378);
xnor U12681 (N_12681,N_10407,N_9496);
xor U12682 (N_12682,N_9620,N_10339);
or U12683 (N_12683,N_11499,N_10127);
or U12684 (N_12684,N_9357,N_9553);
and U12685 (N_12685,N_9053,N_11620);
or U12686 (N_12686,N_9528,N_10468);
nor U12687 (N_12687,N_10193,N_11323);
xor U12688 (N_12688,N_10795,N_11015);
nand U12689 (N_12689,N_11376,N_10295);
nand U12690 (N_12690,N_11422,N_9068);
xor U12691 (N_12691,N_11936,N_10634);
nor U12692 (N_12692,N_11476,N_10079);
or U12693 (N_12693,N_11419,N_11783);
nor U12694 (N_12694,N_11022,N_9267);
xnor U12695 (N_12695,N_9835,N_11996);
nand U12696 (N_12696,N_9915,N_11438);
or U12697 (N_12697,N_9083,N_10069);
nand U12698 (N_12698,N_9837,N_11757);
xnor U12699 (N_12699,N_9188,N_9870);
nand U12700 (N_12700,N_10989,N_10423);
nand U12701 (N_12701,N_10614,N_10644);
xnor U12702 (N_12702,N_11420,N_11289);
and U12703 (N_12703,N_10190,N_11042);
xnor U12704 (N_12704,N_10430,N_9774);
nor U12705 (N_12705,N_11553,N_9358);
and U12706 (N_12706,N_9289,N_11507);
xnor U12707 (N_12707,N_11800,N_10273);
xor U12708 (N_12708,N_9754,N_11613);
nand U12709 (N_12709,N_10091,N_11638);
or U12710 (N_12710,N_10424,N_9493);
nand U12711 (N_12711,N_10075,N_11797);
and U12712 (N_12712,N_11659,N_9274);
xnor U12713 (N_12713,N_11488,N_11707);
nor U12714 (N_12714,N_9143,N_9194);
or U12715 (N_12715,N_10255,N_10847);
and U12716 (N_12716,N_9248,N_11789);
nor U12717 (N_12717,N_11009,N_10073);
or U12718 (N_12718,N_11726,N_11221);
xor U12719 (N_12719,N_11708,N_11717);
nand U12720 (N_12720,N_10938,N_11050);
xor U12721 (N_12721,N_11804,N_9218);
nand U12722 (N_12722,N_9402,N_9433);
nand U12723 (N_12723,N_9725,N_10973);
nor U12724 (N_12724,N_11696,N_11287);
and U12725 (N_12725,N_10233,N_11108);
nor U12726 (N_12726,N_10247,N_9484);
nand U12727 (N_12727,N_9710,N_9690);
nand U12728 (N_12728,N_11427,N_10096);
nor U12729 (N_12729,N_11178,N_9046);
nor U12730 (N_12730,N_10269,N_11954);
nor U12731 (N_12731,N_9059,N_11275);
and U12732 (N_12732,N_11473,N_11100);
xnor U12733 (N_12733,N_9809,N_10316);
xor U12734 (N_12734,N_10380,N_10306);
or U12735 (N_12735,N_11262,N_11114);
nor U12736 (N_12736,N_9899,N_10293);
nand U12737 (N_12737,N_10184,N_11325);
or U12738 (N_12738,N_10397,N_11608);
and U12739 (N_12739,N_11217,N_10573);
nor U12740 (N_12740,N_9501,N_10841);
nand U12741 (N_12741,N_11907,N_10242);
nor U12742 (N_12742,N_10119,N_9552);
or U12743 (N_12743,N_11269,N_9309);
or U12744 (N_12744,N_9971,N_11529);
xnor U12745 (N_12745,N_10887,N_9153);
nand U12746 (N_12746,N_10865,N_10620);
xnor U12747 (N_12747,N_9034,N_9634);
nor U12748 (N_12748,N_9390,N_9829);
or U12749 (N_12749,N_9853,N_9098);
xor U12750 (N_12750,N_11698,N_11639);
or U12751 (N_12751,N_9480,N_11551);
or U12752 (N_12752,N_11937,N_9065);
and U12753 (N_12753,N_9406,N_10353);
or U12754 (N_12754,N_10717,N_10603);
nor U12755 (N_12755,N_11978,N_10413);
xnor U12756 (N_12756,N_10996,N_11951);
nand U12757 (N_12757,N_9308,N_9110);
nand U12758 (N_12758,N_11847,N_10651);
nand U12759 (N_12759,N_10792,N_10108);
xnor U12760 (N_12760,N_10379,N_11548);
xnor U12761 (N_12761,N_9801,N_10403);
or U12762 (N_12762,N_10345,N_9562);
xor U12763 (N_12763,N_10580,N_10649);
nor U12764 (N_12764,N_9185,N_11676);
xor U12765 (N_12765,N_10314,N_11298);
and U12766 (N_12766,N_9454,N_11467);
nand U12767 (N_12767,N_11256,N_9645);
xor U12768 (N_12768,N_9197,N_11248);
or U12769 (N_12769,N_10746,N_10862);
nand U12770 (N_12770,N_10290,N_10941);
nand U12771 (N_12771,N_10821,N_9211);
or U12772 (N_12772,N_10121,N_11480);
and U12773 (N_12773,N_10214,N_9367);
xor U12774 (N_12774,N_11552,N_10161);
or U12775 (N_12775,N_10762,N_10518);
nor U12776 (N_12776,N_10534,N_9295);
and U12777 (N_12777,N_10085,N_9477);
nor U12778 (N_12778,N_11513,N_9872);
or U12779 (N_12779,N_9621,N_9249);
nor U12780 (N_12780,N_10164,N_9908);
or U12781 (N_12781,N_10975,N_11703);
xor U12782 (N_12782,N_11010,N_10997);
xnor U12783 (N_12783,N_9606,N_11856);
nor U12784 (N_12784,N_10760,N_9657);
nand U12785 (N_12785,N_9952,N_9963);
and U12786 (N_12786,N_10872,N_11101);
nor U12787 (N_12787,N_9243,N_11869);
or U12788 (N_12788,N_11249,N_9160);
xor U12789 (N_12789,N_11614,N_10157);
or U12790 (N_12790,N_11543,N_11881);
nor U12791 (N_12791,N_9142,N_9326);
or U12792 (N_12792,N_10970,N_9000);
xnor U12793 (N_12793,N_9236,N_9281);
and U12794 (N_12794,N_10137,N_9052);
nand U12795 (N_12795,N_9427,N_10051);
or U12796 (N_12796,N_9469,N_9912);
nor U12797 (N_12797,N_11402,N_9574);
xor U12798 (N_12798,N_10478,N_9342);
nor U12799 (N_12799,N_9027,N_10776);
nor U12800 (N_12800,N_10621,N_9664);
or U12801 (N_12801,N_11916,N_11667);
xor U12802 (N_12802,N_10450,N_9062);
nor U12803 (N_12803,N_10900,N_11393);
nor U12804 (N_12804,N_11267,N_9630);
nor U12805 (N_12805,N_9051,N_11770);
xor U12806 (N_12806,N_9310,N_10492);
nor U12807 (N_12807,N_11562,N_11137);
or U12808 (N_12808,N_10317,N_9592);
nor U12809 (N_12809,N_10754,N_9440);
or U12810 (N_12810,N_10675,N_10000);
xor U12811 (N_12811,N_10676,N_9995);
and U12812 (N_12812,N_11170,N_10151);
nor U12813 (N_12813,N_9133,N_10490);
nor U12814 (N_12814,N_10670,N_9886);
and U12815 (N_12815,N_9730,N_11372);
or U12816 (N_12816,N_9252,N_11254);
nand U12817 (N_12817,N_11210,N_10266);
nand U12818 (N_12818,N_11649,N_10852);
nor U12819 (N_12819,N_11901,N_9576);
xor U12820 (N_12820,N_9804,N_10195);
nand U12821 (N_12821,N_10465,N_10174);
nand U12822 (N_12822,N_10979,N_10588);
nand U12823 (N_12823,N_11635,N_11474);
nand U12824 (N_12824,N_10693,N_11839);
or U12825 (N_12825,N_10347,N_9106);
xor U12826 (N_12826,N_10204,N_11598);
nand U12827 (N_12827,N_11069,N_10589);
or U12828 (N_12828,N_10775,N_11361);
nand U12829 (N_12829,N_9784,N_10275);
and U12830 (N_12830,N_9324,N_9008);
or U12831 (N_12831,N_10205,N_11312);
and U12832 (N_12832,N_9530,N_9563);
or U12833 (N_12833,N_10249,N_9676);
or U12834 (N_12834,N_9355,N_9609);
xnor U12835 (N_12835,N_10101,N_9508);
xnor U12836 (N_12836,N_10781,N_9447);
and U12837 (N_12837,N_10802,N_9897);
or U12838 (N_12838,N_10338,N_11709);
nor U12839 (N_12839,N_10677,N_9424);
or U12840 (N_12840,N_11725,N_11118);
nand U12841 (N_12841,N_9396,N_11711);
nor U12842 (N_12842,N_11496,N_9923);
or U12843 (N_12843,N_11736,N_10549);
nor U12844 (N_12844,N_11034,N_11105);
xnor U12845 (N_12845,N_10254,N_10326);
nand U12846 (N_12846,N_10244,N_11769);
nand U12847 (N_12847,N_9783,N_10063);
nor U12848 (N_12848,N_10287,N_9584);
and U12849 (N_12849,N_11944,N_10987);
xnor U12850 (N_12850,N_10284,N_9322);
xor U12851 (N_12851,N_10500,N_10041);
nand U12852 (N_12852,N_9593,N_9359);
or U12853 (N_12853,N_9824,N_11690);
or U12854 (N_12854,N_11007,N_9707);
xor U12855 (N_12855,N_9372,N_9131);
or U12856 (N_12856,N_10277,N_11588);
nor U12857 (N_12857,N_9037,N_10268);
nor U12858 (N_12858,N_11411,N_9600);
nor U12859 (N_12859,N_9492,N_10210);
and U12860 (N_12860,N_9255,N_9987);
xor U12861 (N_12861,N_10711,N_9129);
xnor U12862 (N_12862,N_9123,N_9200);
and U12863 (N_12863,N_9729,N_11573);
xor U12864 (N_12864,N_9512,N_11701);
nand U12865 (N_12865,N_11570,N_11729);
nor U12866 (N_12866,N_11301,N_11497);
xnor U12867 (N_12867,N_11401,N_10458);
or U12868 (N_12868,N_11566,N_9466);
and U12869 (N_12869,N_11459,N_10466);
and U12870 (N_12870,N_9331,N_11018);
nand U12871 (N_12871,N_11706,N_10279);
and U12872 (N_12872,N_10129,N_10438);
and U12873 (N_12873,N_11775,N_11129);
and U12874 (N_12874,N_11878,N_10304);
and U12875 (N_12875,N_9115,N_9960);
xnor U12876 (N_12876,N_10092,N_11680);
xnor U12877 (N_12877,N_10398,N_11117);
and U12878 (N_12878,N_10294,N_9316);
nor U12879 (N_12879,N_10008,N_11107);
and U12880 (N_12880,N_10303,N_10203);
nor U12881 (N_12881,N_9256,N_9554);
and U12882 (N_12882,N_11859,N_11145);
and U12883 (N_12883,N_10796,N_10445);
xnor U12884 (N_12884,N_10977,N_10265);
nor U12885 (N_12885,N_9571,N_9036);
nor U12886 (N_12886,N_11424,N_11240);
and U12887 (N_12887,N_10047,N_10289);
xnor U12888 (N_12888,N_11540,N_9749);
or U12889 (N_12889,N_11539,N_11909);
or U12890 (N_12890,N_10828,N_9416);
nand U12891 (N_12891,N_10967,N_9056);
nand U12892 (N_12892,N_11537,N_10685);
nor U12893 (N_12893,N_11794,N_9708);
nor U12894 (N_12894,N_11700,N_9566);
nor U12895 (N_12895,N_11958,N_9327);
and U12896 (N_12896,N_10352,N_11852);
nor U12897 (N_12897,N_10503,N_9400);
xor U12898 (N_12898,N_10133,N_10433);
and U12899 (N_12899,N_11079,N_9269);
nor U12900 (N_12900,N_10535,N_9573);
nor U12901 (N_12901,N_10124,N_9660);
xor U12902 (N_12902,N_11387,N_10031);
nand U12903 (N_12903,N_11150,N_9787);
or U12904 (N_12904,N_9494,N_9775);
or U12905 (N_12905,N_9305,N_10512);
nor U12906 (N_12906,N_11914,N_9073);
and U12907 (N_12907,N_9579,N_11347);
nand U12908 (N_12908,N_9238,N_9412);
nand U12909 (N_12909,N_9700,N_10806);
nor U12910 (N_12910,N_9859,N_9470);
or U12911 (N_12911,N_10176,N_10491);
or U12912 (N_12912,N_11434,N_9614);
or U12913 (N_12913,N_11479,N_11200);
and U12914 (N_12914,N_9162,N_11415);
or U12915 (N_12915,N_10494,N_9444);
and U12916 (N_12916,N_11349,N_9890);
nand U12917 (N_12917,N_11658,N_11663);
and U12918 (N_12918,N_10412,N_11344);
nand U12919 (N_12919,N_9640,N_10139);
nand U12920 (N_12920,N_11702,N_11695);
xnor U12921 (N_12921,N_11453,N_9988);
nor U12922 (N_12922,N_11999,N_9478);
nand U12923 (N_12923,N_9458,N_10297);
or U12924 (N_12924,N_10891,N_9861);
and U12925 (N_12925,N_11637,N_9903);
xor U12926 (N_12926,N_10171,N_10451);
nor U12927 (N_12927,N_11292,N_9354);
or U12928 (N_12928,N_10615,N_9193);
xor U12929 (N_12929,N_10258,N_11932);
or U12930 (N_12930,N_11005,N_10283);
nand U12931 (N_12931,N_11333,N_11067);
nand U12932 (N_12932,N_11354,N_10609);
nor U12933 (N_12933,N_11209,N_10252);
nand U12934 (N_12934,N_11898,N_9832);
or U12935 (N_12935,N_9228,N_11053);
nand U12936 (N_12936,N_9598,N_9146);
or U12937 (N_12937,N_11212,N_11818);
or U12938 (N_12938,N_10298,N_9966);
or U12939 (N_12939,N_9183,N_11330);
nand U12940 (N_12940,N_11961,N_9126);
xnor U12941 (N_12941,N_10601,N_9970);
nor U12942 (N_12942,N_9393,N_9169);
nor U12943 (N_12943,N_9382,N_10076);
nand U12944 (N_12944,N_9043,N_10182);
or U12945 (N_12945,N_11133,N_10013);
nor U12946 (N_12946,N_10388,N_10409);
xor U12947 (N_12947,N_11790,N_11028);
nor U12948 (N_12948,N_11060,N_11578);
nor U12949 (N_12949,N_9456,N_11367);
nand U12950 (N_12950,N_11522,N_10992);
and U12951 (N_12951,N_9237,N_10751);
xnor U12952 (N_12952,N_9259,N_11602);
nand U12953 (N_12953,N_11310,N_11864);
nor U12954 (N_12954,N_10221,N_11475);
or U12955 (N_12955,N_9929,N_10593);
xor U12956 (N_12956,N_9319,N_9580);
nand U12957 (N_12957,N_10542,N_9395);
xor U12958 (N_12958,N_9946,N_11857);
or U12959 (N_12959,N_11661,N_9121);
and U12960 (N_12960,N_9811,N_10842);
nand U12961 (N_12961,N_9356,N_9067);
xnor U12962 (N_12962,N_9199,N_10800);
xnor U12963 (N_12963,N_9288,N_11829);
nand U12964 (N_12964,N_11436,N_10509);
nand U12965 (N_12965,N_10678,N_9586);
and U12966 (N_12966,N_11426,N_9195);
nand U12967 (N_12967,N_10744,N_11300);
and U12968 (N_12968,N_9692,N_9768);
nand U12969 (N_12969,N_9023,N_9994);
or U12970 (N_12970,N_9298,N_11364);
or U12971 (N_12971,N_9875,N_11027);
and U12972 (N_12972,N_9565,N_9240);
and U12973 (N_12973,N_9758,N_11896);
or U12974 (N_12974,N_10667,N_11863);
xor U12975 (N_12975,N_11445,N_11486);
xnor U12976 (N_12976,N_11180,N_9481);
and U12977 (N_12977,N_10460,N_9161);
or U12978 (N_12978,N_11719,N_10162);
nor U12979 (N_12979,N_10110,N_10859);
nor U12980 (N_12980,N_10797,N_10286);
nand U12981 (N_12981,N_11812,N_9074);
xor U12982 (N_12982,N_9147,N_10369);
and U12983 (N_12983,N_10882,N_11892);
nor U12984 (N_12984,N_10474,N_9426);
nand U12985 (N_12985,N_9491,N_10969);
xnor U12986 (N_12986,N_9066,N_10502);
nor U12987 (N_12987,N_9460,N_11315);
nor U12988 (N_12988,N_9900,N_9547);
or U12989 (N_12989,N_9732,N_9924);
nor U12990 (N_12990,N_10569,N_10477);
xor U12991 (N_12991,N_11399,N_9303);
xnor U12992 (N_12992,N_10196,N_11113);
nand U12993 (N_12993,N_11782,N_9796);
and U12994 (N_12994,N_9487,N_10790);
or U12995 (N_12995,N_10831,N_10592);
and U12996 (N_12996,N_9982,N_10618);
nand U12997 (N_12997,N_9216,N_10341);
and U12998 (N_12998,N_10132,N_9032);
xnor U12999 (N_12999,N_10895,N_9042);
xnor U13000 (N_13000,N_11295,N_10654);
nand U13001 (N_13001,N_11922,N_10624);
nand U13002 (N_13002,N_9333,N_11213);
or U13003 (N_13003,N_10350,N_9826);
xnor U13004 (N_13004,N_10929,N_9642);
or U13005 (N_13005,N_10056,N_10695);
and U13006 (N_13006,N_11074,N_11727);
and U13007 (N_13007,N_9196,N_10156);
xnor U13008 (N_13008,N_10516,N_10527);
and U13009 (N_13009,N_10868,N_9800);
xnor U13010 (N_13010,N_10377,N_10674);
and U13011 (N_13011,N_10389,N_9537);
xor U13012 (N_13012,N_11808,N_10229);
nand U13013 (N_13013,N_10885,N_9377);
or U13014 (N_13014,N_9262,N_11592);
and U13015 (N_13015,N_10994,N_9536);
and U13016 (N_13016,N_11955,N_11097);
xnor U13017 (N_13017,N_10679,N_11019);
nor U13018 (N_13018,N_10359,N_9567);
or U13019 (N_13019,N_9849,N_11134);
or U13020 (N_13020,N_11351,N_9208);
nor U13021 (N_13021,N_11068,N_11139);
or U13022 (N_13022,N_9812,N_10443);
and U13023 (N_13023,N_10160,N_9392);
and U13024 (N_13024,N_11666,N_9860);
and U13025 (N_13025,N_9446,N_11791);
nand U13026 (N_13026,N_9975,N_11088);
nor U13027 (N_13027,N_11014,N_11735);
xor U13028 (N_13028,N_10779,N_9341);
nor U13029 (N_13029,N_11685,N_9482);
nor U13030 (N_13030,N_9428,N_11216);
xnor U13031 (N_13031,N_11946,N_9869);
or U13032 (N_13032,N_11432,N_10686);
xor U13033 (N_13033,N_9425,N_11832);
xor U13034 (N_13034,N_11430,N_10995);
nor U13035 (N_13035,N_10354,N_10656);
xnor U13036 (N_13036,N_11989,N_10426);
nand U13037 (N_13037,N_9268,N_11561);
or U13038 (N_13038,N_9499,N_9304);
nor U13039 (N_13039,N_9384,N_10391);
nand U13040 (N_13040,N_10948,N_9901);
and U13041 (N_13041,N_9731,N_9209);
xor U13042 (N_13042,N_9639,N_11448);
or U13043 (N_13043,N_10707,N_10109);
nand U13044 (N_13044,N_9638,N_9284);
xor U13045 (N_13045,N_9442,N_9005);
nand U13046 (N_13046,N_9152,N_9587);
and U13047 (N_13047,N_11255,N_10716);
and U13048 (N_13048,N_11918,N_9159);
and U13049 (N_13049,N_10419,N_10699);
or U13050 (N_13050,N_10922,N_9683);
nor U13051 (N_13051,N_10732,N_9659);
nand U13052 (N_13052,N_11462,N_10364);
nor U13053 (N_13053,N_9763,N_11481);
nand U13054 (N_13054,N_11406,N_11908);
or U13055 (N_13055,N_10368,N_11631);
or U13056 (N_13056,N_11990,N_9107);
and U13057 (N_13057,N_10735,N_9927);
nor U13058 (N_13058,N_11664,N_9504);
nor U13059 (N_13059,N_11498,N_11788);
nor U13060 (N_13060,N_9748,N_9616);
nand U13061 (N_13061,N_10943,N_11489);
xor U13062 (N_13062,N_11574,N_11491);
xnor U13063 (N_13063,N_9138,N_11599);
nand U13064 (N_13064,N_10276,N_9904);
or U13065 (N_13065,N_11077,N_10422);
nand U13066 (N_13066,N_9953,N_10372);
xnor U13067 (N_13067,N_9727,N_9831);
nand U13068 (N_13068,N_9741,N_11960);
and U13069 (N_13069,N_10080,N_10690);
or U13070 (N_13070,N_9315,N_11541);
and U13071 (N_13071,N_9462,N_11959);
and U13072 (N_13072,N_11565,N_11156);
nand U13073 (N_13073,N_10260,N_9109);
or U13074 (N_13074,N_10939,N_10216);
or U13075 (N_13075,N_10785,N_11435);
xnor U13076 (N_13076,N_11307,N_10824);
nor U13077 (N_13077,N_10736,N_10185);
xor U13078 (N_13078,N_9021,N_11373);
or U13079 (N_13079,N_11465,N_11895);
nor U13080 (N_13080,N_11948,N_10278);
xnor U13081 (N_13081,N_9713,N_11380);
xnor U13082 (N_13082,N_11616,N_10700);
and U13083 (N_13083,N_10881,N_9450);
nor U13084 (N_13084,N_10508,N_10102);
xnor U13085 (N_13085,N_10559,N_9471);
xnor U13086 (N_13086,N_11177,N_9823);
xor U13087 (N_13087,N_9542,N_11039);
or U13088 (N_13088,N_11201,N_9127);
and U13089 (N_13089,N_11653,N_9663);
nand U13090 (N_13090,N_10115,N_9118);
nor U13091 (N_13091,N_10627,N_11772);
nand U13092 (N_13092,N_10058,N_11258);
and U13093 (N_13093,N_10498,N_9686);
nor U13094 (N_13094,N_9854,N_10456);
xnor U13095 (N_13095,N_10878,N_11558);
or U13096 (N_13096,N_9280,N_11523);
and U13097 (N_13097,N_11223,N_9794);
xnor U13098 (N_13098,N_11746,N_11439);
or U13099 (N_13099,N_11980,N_11252);
or U13100 (N_13100,N_9818,N_10666);
nor U13101 (N_13101,N_9003,N_9773);
nor U13102 (N_13102,N_11823,N_11952);
and U13103 (N_13103,N_11826,N_11226);
nor U13104 (N_13104,N_9918,N_9421);
and U13105 (N_13105,N_11339,N_10130);
nand U13106 (N_13106,N_10154,N_11521);
nand U13107 (N_13107,N_10919,N_10911);
xor U13108 (N_13108,N_9999,N_11623);
xnor U13109 (N_13109,N_9743,N_9979);
nand U13110 (N_13110,N_11225,N_10864);
xor U13111 (N_13111,N_10488,N_10022);
xor U13112 (N_13112,N_9551,N_10952);
and U13113 (N_13113,N_10152,N_11950);
xnor U13114 (N_13114,N_11545,N_10931);
nand U13115 (N_13115,N_10669,N_9856);
xor U13116 (N_13116,N_9666,N_11147);
nor U13117 (N_13117,N_10658,N_9340);
nor U13118 (N_13118,N_9655,N_11738);
nand U13119 (N_13119,N_9299,N_9201);
or U13120 (N_13120,N_9527,N_11730);
or U13121 (N_13121,N_10636,N_9862);
xor U13122 (N_13122,N_10765,N_9816);
or U13123 (N_13123,N_10883,N_10240);
xor U13124 (N_13124,N_10172,N_9300);
or U13125 (N_13125,N_10198,N_10146);
and U13126 (N_13126,N_10082,N_11278);
or U13127 (N_13127,N_10874,N_10898);
nand U13128 (N_13128,N_11460,N_9232);
nand U13129 (N_13129,N_9282,N_11316);
or U13130 (N_13130,N_10662,N_9044);
nand U13131 (N_13131,N_10764,N_9535);
and U13132 (N_13132,N_10311,N_11677);
nor U13133 (N_13133,N_10905,N_9468);
nand U13134 (N_13134,N_9841,N_9702);
or U13135 (N_13135,N_9541,N_10026);
and U13136 (N_13136,N_9561,N_11604);
nor U13137 (N_13137,N_10715,N_11377);
nor U13138 (N_13138,N_11763,N_9540);
xnor U13139 (N_13139,N_11128,N_9054);
and U13140 (N_13140,N_11382,N_10866);
or U13141 (N_13141,N_11593,N_11934);
and U13142 (N_13142,N_11379,N_11429);
nand U13143 (N_13143,N_9420,N_10055);
nand U13144 (N_13144,N_9155,N_10084);
and U13145 (N_13145,N_9615,N_9665);
nand U13146 (N_13146,N_9233,N_11423);
nand U13147 (N_13147,N_9569,N_11155);
xnor U13148 (N_13148,N_10365,N_11011);
nor U13149 (N_13149,N_10749,N_11628);
and U13150 (N_13150,N_9788,N_9486);
xnor U13151 (N_13151,N_9935,N_10705);
nor U13152 (N_13152,N_11837,N_11388);
or U13153 (N_13153,N_10301,N_11777);
nand U13154 (N_13154,N_11547,N_11140);
nor U13155 (N_13155,N_10371,N_9368);
nand U13156 (N_13156,N_9977,N_11953);
nand U13157 (N_13157,N_10682,N_10803);
nand U13158 (N_13158,N_11297,N_9171);
nand U13159 (N_13159,N_11671,N_9925);
nand U13160 (N_13160,N_11607,N_11585);
nand U13161 (N_13161,N_10811,N_11660);
nand U13162 (N_13162,N_11492,N_9386);
and U13163 (N_13163,N_9435,N_10045);
xnor U13164 (N_13164,N_9836,N_10374);
xor U13165 (N_13165,N_11141,N_9117);
nand U13166 (N_13166,N_11163,N_11964);
and U13167 (N_13167,N_10630,N_10557);
nand U13168 (N_13168,N_11672,N_11290);
nor U13169 (N_13169,N_11279,N_11535);
nand U13170 (N_13170,N_11956,N_10461);
or U13171 (N_13171,N_9214,N_10532);
xnor U13172 (N_13172,N_11461,N_9004);
nand U13173 (N_13173,N_9039,N_10958);
xor U13174 (N_13174,N_9998,N_9076);
and U13175 (N_13175,N_9538,N_11198);
or U13176 (N_13176,N_9050,N_9521);
nand U13177 (N_13177,N_10740,N_9145);
xnor U13178 (N_13178,N_11985,N_11675);
nor U13179 (N_13179,N_9781,N_11131);
xor U13180 (N_13180,N_10059,N_10315);
xnor U13181 (N_13181,N_10089,N_10683);
and U13182 (N_13182,N_10721,N_9422);
or U13183 (N_13183,N_11070,N_9867);
or U13184 (N_13184,N_11317,N_11532);
nor U13185 (N_13185,N_10607,N_10261);
and U13186 (N_13186,N_11017,N_11555);
nor U13187 (N_13187,N_9230,N_9981);
nand U13188 (N_13188,N_9378,N_9762);
nor U13189 (N_13189,N_11748,N_11870);
nor U13190 (N_13190,N_9244,N_10331);
or U13191 (N_13191,N_11051,N_11293);
xnor U13192 (N_13192,N_11283,N_11428);
nor U13193 (N_13193,N_10201,N_9166);
nor U13194 (N_13194,N_10307,N_10954);
and U13195 (N_13195,N_10689,N_10856);
and U13196 (N_13196,N_11362,N_10094);
nor U13197 (N_13197,N_11184,N_10457);
nor U13198 (N_13198,N_10324,N_10793);
nand U13199 (N_13199,N_11000,N_10906);
nand U13200 (N_13200,N_11683,N_11454);
or U13201 (N_13201,N_9954,N_11722);
nor U13202 (N_13202,N_10940,N_11642);
nor U13203 (N_13203,N_10078,N_9863);
or U13204 (N_13204,N_11589,N_9157);
xor U13205 (N_13205,N_10367,N_11302);
and U13206 (N_13206,N_11987,N_11228);
or U13207 (N_13207,N_9864,N_9455);
or U13208 (N_13208,N_9060,N_11405);
nand U13209 (N_13209,N_11109,N_11682);
nor U13210 (N_13210,N_10632,N_10486);
or U13211 (N_13211,N_11629,N_11384);
xnor U13212 (N_13212,N_10714,N_10280);
or U13213 (N_13213,N_9817,N_11575);
nor U13214 (N_13214,N_11923,N_9016);
nor U13215 (N_13215,N_10241,N_9517);
nand U13216 (N_13216,N_9622,N_9352);
xor U13217 (N_13217,N_11657,N_11862);
nand U13218 (N_13218,N_10383,N_9757);
nand U13219 (N_13219,N_10554,N_9597);
nand U13220 (N_13220,N_11242,N_10009);
and U13221 (N_13221,N_9594,N_9696);
or U13222 (N_13222,N_11704,N_11860);
xnor U13223 (N_13223,N_10169,N_10192);
nor U13224 (N_13224,N_10024,N_9687);
or U13225 (N_13225,N_9343,N_10767);
and U13226 (N_13226,N_11630,N_11579);
xnor U13227 (N_13227,N_9087,N_9220);
or U13228 (N_13228,N_10183,N_9124);
nand U13229 (N_13229,N_10479,N_11970);
nor U13230 (N_13230,N_9275,N_11549);
and U13231 (N_13231,N_9624,N_10346);
or U13232 (N_13232,N_10633,N_10142);
nand U13233 (N_13233,N_10541,N_11686);
or U13234 (N_13234,N_11879,N_9325);
nor U13235 (N_13235,N_11135,N_10463);
nand U13236 (N_13236,N_10321,N_10640);
nand U13237 (N_13237,N_9548,N_11328);
nor U13238 (N_13238,N_10418,N_10459);
nor U13239 (N_13239,N_9520,N_11412);
and U13240 (N_13240,N_10692,N_11309);
nor U13241 (N_13241,N_9883,N_9164);
or U13242 (N_13242,N_10187,N_10504);
or U13243 (N_13243,N_11416,N_11931);
or U13244 (N_13244,N_9111,N_9920);
nand U13245 (N_13245,N_9921,N_9879);
nor U13246 (N_13246,N_11055,N_9992);
xor U13247 (N_13247,N_9509,N_9154);
xor U13248 (N_13248,N_11020,N_9910);
nand U13249 (N_13249,N_10855,N_9636);
nand U13250 (N_13250,N_11083,N_9497);
nor U13251 (N_13251,N_10222,N_11583);
xor U13252 (N_13252,N_10355,N_11851);
and U13253 (N_13253,N_11260,N_10815);
xnor U13254 (N_13254,N_9514,N_10036);
nand U13255 (N_13255,N_9607,N_9419);
nand U13256 (N_13256,N_10550,N_9961);
nor U13257 (N_13257,N_11494,N_9277);
and U13258 (N_13258,N_10596,N_10032);
nor U13259 (N_13259,N_11752,N_11820);
and U13260 (N_13260,N_10469,N_10953);
nor U13261 (N_13261,N_11322,N_10197);
or U13262 (N_13262,N_11157,N_10738);
and U13263 (N_13263,N_9735,N_11215);
and U13264 (N_13264,N_10484,N_11390);
xnor U13265 (N_13265,N_11670,N_10267);
or U13266 (N_13266,N_11166,N_9653);
nand U13267 (N_13267,N_10552,N_11835);
or U13268 (N_13268,N_10238,N_10462);
and U13269 (N_13269,N_11208,N_11250);
xor U13270 (N_13270,N_9604,N_10709);
xor U13271 (N_13271,N_10226,N_9962);
and U13272 (N_13272,N_11504,N_9873);
nand U13273 (N_13273,N_11341,N_10827);
nand U13274 (N_13274,N_10753,N_9990);
nor U13275 (N_13275,N_9533,N_11779);
nor U13276 (N_13276,N_11761,N_11345);
nor U13277 (N_13277,N_11611,N_11218);
nor U13278 (N_13278,N_10928,N_9346);
or U13279 (N_13279,N_11253,N_10296);
xor U13280 (N_13280,N_9839,N_9764);
nor U13281 (N_13281,N_11526,N_9723);
nor U13282 (N_13282,N_10867,N_11276);
nand U13283 (N_13283,N_9556,N_11595);
nand U13284 (N_13284,N_10538,N_10220);
or U13285 (N_13285,N_10742,N_9983);
xnor U13286 (N_13286,N_11431,N_11024);
nor U13287 (N_13287,N_10122,N_10935);
or U13288 (N_13288,N_9388,N_9292);
nand U13289 (N_13289,N_10166,N_11185);
xnor U13290 (N_13290,N_10027,N_11887);
xnor U13291 (N_13291,N_9578,N_11119);
xnor U13292 (N_13292,N_11986,N_9510);
nand U13293 (N_13293,N_10880,N_9335);
or U13294 (N_13294,N_9674,N_9475);
nand U13295 (N_13295,N_11949,N_9684);
nor U13296 (N_13296,N_9955,N_9555);
nor U13297 (N_13297,N_10850,N_10476);
nand U13298 (N_13298,N_11179,N_10305);
xnor U13299 (N_13299,N_11149,N_10143);
nor U13300 (N_13300,N_11796,N_10400);
xnor U13301 (N_13301,N_11511,N_9969);
nor U13302 (N_13302,N_11884,N_9617);
nand U13303 (N_13303,N_10432,N_11280);
xnor U13304 (N_13304,N_10444,N_10511);
and U13305 (N_13305,N_11888,N_9202);
or U13306 (N_13306,N_9734,N_11903);
or U13307 (N_13307,N_11482,N_9868);
nand U13308 (N_13308,N_9351,N_11121);
nor U13309 (N_13309,N_10648,N_11755);
nor U13310 (N_13310,N_11092,N_9167);
nor U13311 (N_13311,N_10054,N_11780);
nand U13312 (N_13312,N_10565,N_9944);
nor U13313 (N_13313,N_11924,N_10912);
or U13314 (N_13314,N_11191,N_11023);
nand U13315 (N_13315,N_11158,N_9771);
nand U13316 (N_13316,N_9967,N_11745);
xor U13317 (N_13317,N_11920,N_9611);
and U13318 (N_13318,N_11885,N_11169);
xor U13319 (N_13319,N_10040,N_10530);
or U13320 (N_13320,N_11353,N_9529);
or U13321 (N_13321,N_10529,N_11619);
and U13322 (N_13322,N_9755,N_10499);
or U13323 (N_13323,N_11821,N_10467);
nor U13324 (N_13324,N_10916,N_9772);
nand U13325 (N_13325,N_11648,N_11572);
nor U13326 (N_13326,N_11744,N_9314);
or U13327 (N_13327,N_9635,N_10983);
or U13328 (N_13328,N_10048,N_10606);
and U13329 (N_13329,N_10830,N_10932);
nor U13330 (N_13330,N_10808,N_10756);
or U13331 (N_13331,N_10934,N_11875);
nor U13332 (N_13332,N_9777,N_10387);
or U13333 (N_13333,N_10211,N_11605);
xor U13334 (N_13334,N_10729,N_11045);
nand U13335 (N_13335,N_9364,N_10288);
nand U13336 (N_13336,N_9410,N_9793);
or U13337 (N_13337,N_10814,N_10163);
and U13338 (N_13338,N_11687,N_9048);
nand U13339 (N_13339,N_9158,N_10207);
nand U13340 (N_13340,N_10702,N_11811);
nand U13341 (N_13341,N_10946,N_10505);
xnor U13342 (N_13342,N_11713,N_10246);
and U13343 (N_13343,N_9099,N_11103);
nand U13344 (N_13344,N_11146,N_10470);
nor U13345 (N_13345,N_10833,N_10957);
nor U13346 (N_13346,N_10057,N_9221);
or U13347 (N_13347,N_11534,N_11203);
nor U13348 (N_13348,N_10004,N_9575);
nor U13349 (N_13349,N_9568,N_10010);
nand U13350 (N_13350,N_10637,N_9029);
and U13351 (N_13351,N_11063,N_9997);
and U13352 (N_13352,N_11503,N_11699);
xnor U13353 (N_13353,N_11721,N_9140);
nand U13354 (N_13354,N_11085,N_9104);
xor U13355 (N_13355,N_10892,N_10385);
and U13356 (N_13356,N_11151,N_11530);
and U13357 (N_13357,N_9082,N_10113);
or U13358 (N_13358,N_9711,N_10927);
xor U13359 (N_13359,N_11560,N_11935);
xnor U13360 (N_13360,N_9439,N_11760);
or U13361 (N_13361,N_9387,N_10481);
nand U13362 (N_13362,N_10597,N_11052);
nor U13363 (N_13363,N_11171,N_10357);
xnor U13364 (N_13364,N_10902,N_11485);
and U13365 (N_13365,N_11458,N_9231);
and U13366 (N_13366,N_10982,N_9017);
or U13367 (N_13367,N_10149,N_9557);
xnor U13368 (N_13368,N_9884,N_9544);
nand U13369 (N_13369,N_10434,N_11144);
nand U13370 (N_13370,N_9917,N_10799);
and U13371 (N_13371,N_9321,N_11926);
xor U13372 (N_13372,N_11803,N_11437);
nor U13373 (N_13373,N_10104,N_11943);
and U13374 (N_13374,N_10100,N_9263);
or U13375 (N_13375,N_9323,N_11304);
nand U13376 (N_13376,N_9795,N_9094);
xor U13377 (N_13377,N_9679,N_10854);
nor U13378 (N_13378,N_9229,N_11059);
and U13379 (N_13379,N_10999,N_9888);
nor U13380 (N_13380,N_9689,N_11563);
xor U13381 (N_13381,N_9641,N_11365);
xnor U13382 (N_13382,N_11833,N_11814);
nor U13383 (N_13383,N_11911,N_9245);
and U13384 (N_13384,N_9892,N_11441);
or U13385 (N_13385,N_10188,N_10181);
xor U13386 (N_13386,N_9648,N_9186);
and U13387 (N_13387,N_10309,N_10556);
nor U13388 (N_13388,N_9761,N_9414);
nand U13389 (N_13389,N_9408,N_11449);
or U13390 (N_13390,N_10417,N_9398);
and U13391 (N_13391,N_10787,N_11303);
and U13392 (N_13392,N_10673,N_10914);
xnor U13393 (N_13393,N_10585,N_11268);
and U13394 (N_13394,N_10312,N_11728);
nand U13395 (N_13395,N_11308,N_10558);
and U13396 (N_13396,N_9389,N_10131);
xnor U13397 (N_13397,N_9747,N_11976);
nand U13398 (N_13398,N_10408,N_9345);
nand U13399 (N_13399,N_11855,N_10761);
nand U13400 (N_13400,N_11003,N_10173);
nor U13401 (N_13401,N_10617,N_9271);
nand U13402 (N_13402,N_9906,N_11600);
and U13403 (N_13403,N_11483,N_11603);
and U13404 (N_13404,N_10645,N_9362);
and U13405 (N_13405,N_11370,N_9516);
xnor U13406 (N_13406,N_10590,N_11597);
nand U13407 (N_13407,N_10568,N_10773);
or U13408 (N_13408,N_10225,N_10956);
nor U13409 (N_13409,N_9822,N_10861);
xor U13410 (N_13410,N_10037,N_9366);
nand U13411 (N_13411,N_11282,N_11102);
xor U13412 (N_13412,N_11164,N_11890);
and U13413 (N_13413,N_10526,N_10930);
nand U13414 (N_13414,N_10006,N_9102);
nor U13415 (N_13415,N_11187,N_10671);
nand U13416 (N_13416,N_10555,N_10179);
and U13417 (N_13417,N_11827,N_11802);
or U13418 (N_13418,N_11204,N_10446);
nor U13419 (N_13419,N_10965,N_9790);
xnor U13420 (N_13420,N_9313,N_9814);
nand U13421 (N_13421,N_10560,N_9020);
xnor U13422 (N_13422,N_9778,N_9799);
nor U13423 (N_13423,N_9353,N_11567);
xor U13424 (N_13424,N_9178,N_9756);
or U13425 (N_13425,N_10217,N_11919);
and U13426 (N_13426,N_9149,N_11544);
nand U13427 (N_13427,N_9063,N_11001);
and U13428 (N_13428,N_10734,N_11142);
and U13429 (N_13429,N_9055,N_11854);
nor U13430 (N_13430,N_9379,N_9559);
xor U13431 (N_13431,N_10819,N_9618);
nor U13432 (N_13432,N_10441,N_9135);
or U13433 (N_13433,N_11787,N_11096);
or U13434 (N_13434,N_10962,N_11220);
or U13435 (N_13435,N_9203,N_11219);
and U13436 (N_13436,N_9724,N_9834);
nand U13437 (N_13437,N_9765,N_11090);
and U13438 (N_13438,N_11065,N_10777);
and U13439 (N_13439,N_9219,N_9212);
xnor U13440 (N_13440,N_10837,N_10392);
xor U13441 (N_13441,N_10393,N_10959);
xnor U13442 (N_13442,N_9035,N_11374);
nand U13443 (N_13443,N_11838,N_11484);
or U13444 (N_13444,N_10454,N_11306);
nand U13445 (N_13445,N_9613,N_11542);
nand U13446 (N_13446,N_11176,N_10990);
nor U13447 (N_13447,N_11785,N_10835);
nor U13448 (N_13448,N_10515,N_9570);
nand U13449 (N_13449,N_11397,N_10974);
and U13450 (N_13450,N_11991,N_10823);
or U13451 (N_13451,N_10325,N_11008);
or U13452 (N_13452,N_11740,N_11167);
and U13453 (N_13453,N_9500,N_9290);
xnor U13454 (N_13454,N_9751,N_10416);
nand U13455 (N_13455,N_10302,N_11518);
or U13456 (N_13456,N_10165,N_9217);
nor U13457 (N_13457,N_9866,N_11125);
xor U13458 (N_13458,N_10647,N_10951);
nor U13459 (N_13459,N_9515,N_9329);
or U13460 (N_13460,N_9213,N_9033);
and U13461 (N_13461,N_9241,N_10219);
nand U13462 (N_13462,N_9122,N_9821);
and U13463 (N_13463,N_9522,N_10344);
and U13464 (N_13464,N_10748,N_10189);
or U13465 (N_13465,N_10328,N_9344);
nand U13466 (N_13466,N_11894,N_9093);
xnor U13467 (N_13467,N_11327,N_10395);
and U13468 (N_13468,N_9403,N_11232);
nor U13469 (N_13469,N_11251,N_11369);
or U13470 (N_13470,N_11617,N_11231);
and U13471 (N_13471,N_11094,N_10274);
xor U13472 (N_13472,N_9909,N_10691);
xnor U13473 (N_13473,N_9465,N_10095);
and U13474 (N_13474,N_11747,N_10017);
xor U13475 (N_13475,N_9543,N_9647);
and U13476 (N_13476,N_9174,N_10816);
xor U13477 (N_13477,N_10712,N_10574);
or U13478 (N_13478,N_9688,N_10901);
or U13479 (N_13479,N_9718,N_11689);
xor U13480 (N_13480,N_9251,N_9808);
and U13481 (N_13481,N_9047,N_10608);
and U13482 (N_13482,N_9699,N_9394);
or U13483 (N_13483,N_9993,N_11030);
and U13484 (N_13484,N_11244,N_11694);
nor U13485 (N_13485,N_11988,N_10587);
nand U13486 (N_13486,N_10170,N_10429);
and U13487 (N_13487,N_10539,N_9279);
xnor U13488 (N_13488,N_11712,N_10414);
nor U13489 (N_13489,N_10435,N_11759);
and U13490 (N_13490,N_11531,N_9374);
or U13491 (N_13491,N_11259,N_11741);
xnor U13492 (N_13492,N_10050,N_11945);
or U13493 (N_13493,N_11175,N_11799);
nand U13494 (N_13494,N_11152,N_11900);
xnor U13495 (N_13495,N_11586,N_9151);
and U13496 (N_13496,N_10622,N_10281);
xnor U13497 (N_13497,N_9572,N_9874);
nand U13498 (N_13498,N_11285,N_11224);
nand U13499 (N_13499,N_11038,N_9443);
and U13500 (N_13500,N_9145,N_11683);
and U13501 (N_13501,N_9301,N_10643);
or U13502 (N_13502,N_9623,N_10740);
nor U13503 (N_13503,N_9783,N_9451);
and U13504 (N_13504,N_11836,N_11246);
nor U13505 (N_13505,N_10946,N_10442);
xnor U13506 (N_13506,N_9693,N_11025);
nor U13507 (N_13507,N_11690,N_10466);
nand U13508 (N_13508,N_11694,N_10265);
xor U13509 (N_13509,N_10751,N_10640);
nor U13510 (N_13510,N_9398,N_9499);
xnor U13511 (N_13511,N_10022,N_9936);
nand U13512 (N_13512,N_9763,N_9712);
or U13513 (N_13513,N_9770,N_10349);
xor U13514 (N_13514,N_10850,N_11748);
xnor U13515 (N_13515,N_11578,N_10245);
xnor U13516 (N_13516,N_11231,N_11413);
and U13517 (N_13517,N_9768,N_10100);
xnor U13518 (N_13518,N_9790,N_10280);
or U13519 (N_13519,N_10089,N_9571);
and U13520 (N_13520,N_9122,N_10479);
nand U13521 (N_13521,N_10237,N_11225);
nand U13522 (N_13522,N_9166,N_11366);
nand U13523 (N_13523,N_10577,N_10215);
or U13524 (N_13524,N_10792,N_10739);
xor U13525 (N_13525,N_10069,N_11997);
nor U13526 (N_13526,N_11636,N_11861);
nor U13527 (N_13527,N_10325,N_9892);
or U13528 (N_13528,N_10815,N_10304);
or U13529 (N_13529,N_9768,N_10899);
nor U13530 (N_13530,N_10555,N_9959);
or U13531 (N_13531,N_11661,N_10938);
nand U13532 (N_13532,N_9061,N_10379);
nand U13533 (N_13533,N_10167,N_9624);
or U13534 (N_13534,N_9720,N_10780);
or U13535 (N_13535,N_11306,N_9531);
nor U13536 (N_13536,N_11804,N_9026);
or U13537 (N_13537,N_11761,N_10782);
nor U13538 (N_13538,N_9421,N_10109);
nand U13539 (N_13539,N_10475,N_9802);
or U13540 (N_13540,N_11813,N_11066);
or U13541 (N_13541,N_9447,N_10669);
nor U13542 (N_13542,N_10606,N_10328);
xnor U13543 (N_13543,N_9217,N_11816);
xnor U13544 (N_13544,N_11302,N_11055);
or U13545 (N_13545,N_10782,N_11016);
nand U13546 (N_13546,N_11114,N_9551);
xor U13547 (N_13547,N_9658,N_11960);
xnor U13548 (N_13548,N_9165,N_10336);
xor U13549 (N_13549,N_10889,N_11468);
and U13550 (N_13550,N_9016,N_11954);
xnor U13551 (N_13551,N_9708,N_11839);
nor U13552 (N_13552,N_10275,N_10255);
nor U13553 (N_13553,N_11920,N_9223);
xor U13554 (N_13554,N_11680,N_10482);
and U13555 (N_13555,N_10539,N_11237);
nand U13556 (N_13556,N_9465,N_9154);
and U13557 (N_13557,N_11012,N_10496);
xnor U13558 (N_13558,N_11172,N_10481);
nor U13559 (N_13559,N_9565,N_11090);
or U13560 (N_13560,N_11691,N_10423);
or U13561 (N_13561,N_11624,N_11499);
or U13562 (N_13562,N_11689,N_9666);
nor U13563 (N_13563,N_10835,N_11297);
nand U13564 (N_13564,N_11586,N_9801);
nand U13565 (N_13565,N_11381,N_11097);
xor U13566 (N_13566,N_11732,N_9301);
xor U13567 (N_13567,N_11457,N_10241);
xor U13568 (N_13568,N_9406,N_10006);
and U13569 (N_13569,N_11275,N_9320);
or U13570 (N_13570,N_10336,N_9417);
nor U13571 (N_13571,N_11938,N_11718);
nand U13572 (N_13572,N_9240,N_10650);
xor U13573 (N_13573,N_11891,N_11499);
nand U13574 (N_13574,N_11923,N_11973);
nor U13575 (N_13575,N_11834,N_9050);
xnor U13576 (N_13576,N_10592,N_11870);
nor U13577 (N_13577,N_10017,N_10649);
xnor U13578 (N_13578,N_9180,N_9068);
nor U13579 (N_13579,N_10919,N_11113);
xor U13580 (N_13580,N_11296,N_10938);
xor U13581 (N_13581,N_10412,N_10472);
nor U13582 (N_13582,N_11188,N_9090);
nor U13583 (N_13583,N_10374,N_9627);
or U13584 (N_13584,N_11928,N_10609);
and U13585 (N_13585,N_11270,N_10063);
nand U13586 (N_13586,N_11178,N_11113);
xor U13587 (N_13587,N_11895,N_9564);
and U13588 (N_13588,N_11735,N_9579);
nor U13589 (N_13589,N_10951,N_11881);
xor U13590 (N_13590,N_10169,N_10937);
and U13591 (N_13591,N_11015,N_10028);
and U13592 (N_13592,N_11104,N_11962);
xor U13593 (N_13593,N_10628,N_10937);
nor U13594 (N_13594,N_9354,N_9136);
and U13595 (N_13595,N_10725,N_11474);
nand U13596 (N_13596,N_11779,N_10788);
nand U13597 (N_13597,N_9455,N_9100);
nor U13598 (N_13598,N_9759,N_10500);
nor U13599 (N_13599,N_9438,N_11849);
nand U13600 (N_13600,N_11351,N_9836);
xnor U13601 (N_13601,N_10777,N_11669);
nand U13602 (N_13602,N_9550,N_10028);
and U13603 (N_13603,N_9373,N_9431);
or U13604 (N_13604,N_9471,N_10870);
or U13605 (N_13605,N_10830,N_10115);
nand U13606 (N_13606,N_11922,N_10074);
xnor U13607 (N_13607,N_9374,N_9117);
or U13608 (N_13608,N_11788,N_9416);
xor U13609 (N_13609,N_10244,N_9709);
nor U13610 (N_13610,N_11409,N_11537);
nand U13611 (N_13611,N_11181,N_10668);
or U13612 (N_13612,N_11959,N_11611);
or U13613 (N_13613,N_11979,N_11218);
xor U13614 (N_13614,N_9076,N_11860);
and U13615 (N_13615,N_9874,N_9812);
xor U13616 (N_13616,N_11547,N_11323);
nor U13617 (N_13617,N_11518,N_10868);
or U13618 (N_13618,N_11724,N_9559);
and U13619 (N_13619,N_11493,N_9652);
and U13620 (N_13620,N_9404,N_9483);
nand U13621 (N_13621,N_10347,N_9884);
nor U13622 (N_13622,N_11248,N_10968);
or U13623 (N_13623,N_10142,N_11931);
xnor U13624 (N_13624,N_9466,N_9254);
nor U13625 (N_13625,N_11714,N_10460);
and U13626 (N_13626,N_10079,N_11487);
or U13627 (N_13627,N_11486,N_11213);
nand U13628 (N_13628,N_9619,N_10434);
nand U13629 (N_13629,N_11049,N_11057);
or U13630 (N_13630,N_11628,N_11668);
xor U13631 (N_13631,N_10571,N_9399);
nor U13632 (N_13632,N_11665,N_10288);
and U13633 (N_13633,N_11514,N_9852);
nand U13634 (N_13634,N_10142,N_10907);
nand U13635 (N_13635,N_9548,N_10677);
and U13636 (N_13636,N_11812,N_9618);
nand U13637 (N_13637,N_10968,N_10190);
and U13638 (N_13638,N_10839,N_9300);
nor U13639 (N_13639,N_9745,N_9954);
and U13640 (N_13640,N_9562,N_11746);
xor U13641 (N_13641,N_11259,N_9993);
or U13642 (N_13642,N_11214,N_9509);
or U13643 (N_13643,N_9920,N_9042);
xnor U13644 (N_13644,N_10925,N_9050);
or U13645 (N_13645,N_11475,N_11300);
nor U13646 (N_13646,N_11833,N_9136);
nor U13647 (N_13647,N_11614,N_11446);
xor U13648 (N_13648,N_9160,N_10943);
and U13649 (N_13649,N_10198,N_9537);
xnor U13650 (N_13650,N_10624,N_10155);
xnor U13651 (N_13651,N_10977,N_11294);
nand U13652 (N_13652,N_11687,N_10664);
nand U13653 (N_13653,N_11877,N_11558);
nand U13654 (N_13654,N_9485,N_9779);
nor U13655 (N_13655,N_10550,N_11595);
nand U13656 (N_13656,N_11299,N_9005);
nand U13657 (N_13657,N_11188,N_11664);
nor U13658 (N_13658,N_9354,N_11961);
and U13659 (N_13659,N_10543,N_11261);
xnor U13660 (N_13660,N_10951,N_9162);
nor U13661 (N_13661,N_10457,N_11990);
nand U13662 (N_13662,N_10080,N_10969);
and U13663 (N_13663,N_10572,N_11362);
and U13664 (N_13664,N_10166,N_9738);
and U13665 (N_13665,N_11307,N_10453);
nand U13666 (N_13666,N_9709,N_11780);
xor U13667 (N_13667,N_9983,N_9230);
and U13668 (N_13668,N_10069,N_10641);
xor U13669 (N_13669,N_9323,N_10416);
xor U13670 (N_13670,N_9931,N_10342);
nand U13671 (N_13671,N_10692,N_9449);
and U13672 (N_13672,N_11410,N_9892);
nor U13673 (N_13673,N_11057,N_11832);
xor U13674 (N_13674,N_9050,N_10628);
nor U13675 (N_13675,N_10467,N_11681);
nand U13676 (N_13676,N_11826,N_11391);
and U13677 (N_13677,N_10761,N_9173);
nor U13678 (N_13678,N_11423,N_10021);
nand U13679 (N_13679,N_9046,N_11713);
nor U13680 (N_13680,N_9673,N_9009);
nand U13681 (N_13681,N_10796,N_11965);
or U13682 (N_13682,N_11443,N_10368);
or U13683 (N_13683,N_10948,N_9581);
nor U13684 (N_13684,N_9163,N_10613);
nor U13685 (N_13685,N_11175,N_10619);
and U13686 (N_13686,N_9797,N_11294);
and U13687 (N_13687,N_9649,N_10431);
xnor U13688 (N_13688,N_11740,N_10921);
xnor U13689 (N_13689,N_9660,N_10976);
and U13690 (N_13690,N_11025,N_11917);
xnor U13691 (N_13691,N_10973,N_10704);
xnor U13692 (N_13692,N_10285,N_11749);
nand U13693 (N_13693,N_9890,N_11158);
nor U13694 (N_13694,N_11440,N_11749);
nand U13695 (N_13695,N_11464,N_11280);
and U13696 (N_13696,N_10345,N_11932);
xor U13697 (N_13697,N_11776,N_10469);
nor U13698 (N_13698,N_9101,N_10547);
nand U13699 (N_13699,N_9060,N_9903);
nand U13700 (N_13700,N_10005,N_10157);
and U13701 (N_13701,N_11225,N_9815);
nor U13702 (N_13702,N_9222,N_10746);
nor U13703 (N_13703,N_11260,N_10786);
and U13704 (N_13704,N_10698,N_9991);
and U13705 (N_13705,N_10597,N_9178);
or U13706 (N_13706,N_10555,N_9541);
nor U13707 (N_13707,N_9175,N_10737);
and U13708 (N_13708,N_10173,N_11095);
or U13709 (N_13709,N_9926,N_11504);
or U13710 (N_13710,N_10359,N_10095);
nor U13711 (N_13711,N_9884,N_11824);
and U13712 (N_13712,N_9645,N_11605);
nand U13713 (N_13713,N_9619,N_10424);
xor U13714 (N_13714,N_10884,N_11246);
nand U13715 (N_13715,N_11959,N_11374);
and U13716 (N_13716,N_10749,N_11551);
and U13717 (N_13717,N_10327,N_11881);
xor U13718 (N_13718,N_11959,N_11995);
xnor U13719 (N_13719,N_11181,N_10755);
and U13720 (N_13720,N_10230,N_9177);
nand U13721 (N_13721,N_9079,N_9735);
nor U13722 (N_13722,N_11184,N_10672);
nor U13723 (N_13723,N_10971,N_10448);
or U13724 (N_13724,N_11278,N_9914);
and U13725 (N_13725,N_11800,N_11071);
or U13726 (N_13726,N_9047,N_10634);
nor U13727 (N_13727,N_10167,N_9234);
nand U13728 (N_13728,N_9331,N_11825);
nand U13729 (N_13729,N_11951,N_9621);
nor U13730 (N_13730,N_9656,N_10008);
and U13731 (N_13731,N_10585,N_10484);
and U13732 (N_13732,N_9412,N_10953);
or U13733 (N_13733,N_9311,N_11187);
nand U13734 (N_13734,N_10117,N_11489);
or U13735 (N_13735,N_11603,N_11701);
or U13736 (N_13736,N_9666,N_11708);
or U13737 (N_13737,N_9918,N_10070);
nor U13738 (N_13738,N_9557,N_10330);
nand U13739 (N_13739,N_10807,N_11119);
nand U13740 (N_13740,N_9370,N_9746);
nor U13741 (N_13741,N_10736,N_10097);
or U13742 (N_13742,N_11298,N_10600);
xnor U13743 (N_13743,N_10422,N_10540);
nand U13744 (N_13744,N_10522,N_11119);
or U13745 (N_13745,N_11667,N_11031);
and U13746 (N_13746,N_9206,N_9550);
xor U13747 (N_13747,N_11276,N_10224);
nand U13748 (N_13748,N_11752,N_11307);
nand U13749 (N_13749,N_9118,N_9468);
or U13750 (N_13750,N_9498,N_11848);
xnor U13751 (N_13751,N_9420,N_10836);
xor U13752 (N_13752,N_11174,N_9069);
or U13753 (N_13753,N_10989,N_10961);
nand U13754 (N_13754,N_11519,N_11562);
nand U13755 (N_13755,N_9241,N_10827);
xnor U13756 (N_13756,N_11735,N_9364);
or U13757 (N_13757,N_9583,N_10323);
xnor U13758 (N_13758,N_10257,N_9095);
or U13759 (N_13759,N_10627,N_9897);
or U13760 (N_13760,N_10401,N_10226);
or U13761 (N_13761,N_10175,N_11387);
and U13762 (N_13762,N_10265,N_9096);
xor U13763 (N_13763,N_11201,N_10794);
nand U13764 (N_13764,N_11676,N_11274);
and U13765 (N_13765,N_11871,N_10673);
xor U13766 (N_13766,N_9262,N_9142);
and U13767 (N_13767,N_9800,N_10451);
xor U13768 (N_13768,N_10632,N_10329);
nor U13769 (N_13769,N_11053,N_10978);
nor U13770 (N_13770,N_10806,N_10997);
and U13771 (N_13771,N_10163,N_9818);
xnor U13772 (N_13772,N_10728,N_11780);
or U13773 (N_13773,N_10720,N_11348);
xnor U13774 (N_13774,N_11120,N_9124);
and U13775 (N_13775,N_10012,N_11698);
nand U13776 (N_13776,N_10336,N_10130);
nand U13777 (N_13777,N_9801,N_9081);
xor U13778 (N_13778,N_9352,N_10741);
and U13779 (N_13779,N_10944,N_11388);
nand U13780 (N_13780,N_10737,N_9318);
and U13781 (N_13781,N_9329,N_9673);
or U13782 (N_13782,N_9307,N_9740);
or U13783 (N_13783,N_9356,N_10598);
and U13784 (N_13784,N_10816,N_10830);
xor U13785 (N_13785,N_9664,N_9356);
or U13786 (N_13786,N_11431,N_9119);
xnor U13787 (N_13787,N_9478,N_10424);
nand U13788 (N_13788,N_11321,N_11311);
nor U13789 (N_13789,N_11768,N_9512);
and U13790 (N_13790,N_10757,N_11396);
nand U13791 (N_13791,N_9530,N_10613);
and U13792 (N_13792,N_11253,N_10635);
nor U13793 (N_13793,N_11401,N_9796);
nor U13794 (N_13794,N_11961,N_11184);
nor U13795 (N_13795,N_11648,N_9397);
nor U13796 (N_13796,N_11278,N_9450);
nand U13797 (N_13797,N_9358,N_9797);
or U13798 (N_13798,N_9511,N_9801);
or U13799 (N_13799,N_9253,N_10093);
and U13800 (N_13800,N_11692,N_11926);
nand U13801 (N_13801,N_10241,N_11787);
xor U13802 (N_13802,N_9205,N_9855);
nor U13803 (N_13803,N_11986,N_11322);
xor U13804 (N_13804,N_9420,N_10966);
xor U13805 (N_13805,N_9176,N_11411);
or U13806 (N_13806,N_9570,N_10429);
xor U13807 (N_13807,N_11864,N_11616);
and U13808 (N_13808,N_11263,N_9740);
nor U13809 (N_13809,N_9127,N_11920);
or U13810 (N_13810,N_10885,N_11425);
nor U13811 (N_13811,N_9365,N_9104);
or U13812 (N_13812,N_10965,N_9721);
nand U13813 (N_13813,N_10983,N_11454);
xnor U13814 (N_13814,N_10384,N_9604);
xnor U13815 (N_13815,N_11602,N_9367);
nand U13816 (N_13816,N_9242,N_9451);
nor U13817 (N_13817,N_10961,N_11562);
nor U13818 (N_13818,N_10709,N_11202);
nor U13819 (N_13819,N_10604,N_11858);
nand U13820 (N_13820,N_10796,N_9401);
or U13821 (N_13821,N_9778,N_10300);
xor U13822 (N_13822,N_11175,N_11871);
and U13823 (N_13823,N_10330,N_11344);
xnor U13824 (N_13824,N_10066,N_10669);
and U13825 (N_13825,N_11100,N_9346);
or U13826 (N_13826,N_9490,N_9223);
nor U13827 (N_13827,N_10084,N_10168);
and U13828 (N_13828,N_11608,N_9389);
or U13829 (N_13829,N_10164,N_11638);
nand U13830 (N_13830,N_11835,N_11778);
or U13831 (N_13831,N_10389,N_10042);
and U13832 (N_13832,N_9032,N_10554);
xor U13833 (N_13833,N_10906,N_11210);
xor U13834 (N_13834,N_9517,N_9062);
nor U13835 (N_13835,N_10951,N_11516);
nand U13836 (N_13836,N_9766,N_9088);
and U13837 (N_13837,N_9912,N_10274);
or U13838 (N_13838,N_9630,N_9719);
nor U13839 (N_13839,N_9045,N_10631);
and U13840 (N_13840,N_10062,N_11856);
or U13841 (N_13841,N_10170,N_9944);
xnor U13842 (N_13842,N_9900,N_9377);
or U13843 (N_13843,N_10094,N_10905);
nand U13844 (N_13844,N_10664,N_9601);
xor U13845 (N_13845,N_11090,N_10101);
xnor U13846 (N_13846,N_11453,N_10963);
nor U13847 (N_13847,N_9547,N_9019);
xnor U13848 (N_13848,N_10985,N_9826);
or U13849 (N_13849,N_10474,N_10827);
or U13850 (N_13850,N_9758,N_9371);
nand U13851 (N_13851,N_9927,N_10243);
or U13852 (N_13852,N_11149,N_10694);
nand U13853 (N_13853,N_10849,N_10349);
xor U13854 (N_13854,N_10866,N_10355);
and U13855 (N_13855,N_9968,N_11866);
or U13856 (N_13856,N_10244,N_11834);
xor U13857 (N_13857,N_9667,N_10521);
nor U13858 (N_13858,N_9169,N_10854);
nor U13859 (N_13859,N_11566,N_9386);
or U13860 (N_13860,N_9354,N_10083);
xnor U13861 (N_13861,N_9882,N_9084);
xor U13862 (N_13862,N_11102,N_11978);
xor U13863 (N_13863,N_11637,N_10807);
or U13864 (N_13864,N_10622,N_11732);
and U13865 (N_13865,N_9254,N_11045);
nand U13866 (N_13866,N_11939,N_10278);
xnor U13867 (N_13867,N_10299,N_10899);
and U13868 (N_13868,N_9597,N_10505);
xor U13869 (N_13869,N_10738,N_11683);
or U13870 (N_13870,N_11542,N_9214);
and U13871 (N_13871,N_9184,N_11409);
nand U13872 (N_13872,N_9148,N_11285);
nor U13873 (N_13873,N_11586,N_11279);
nor U13874 (N_13874,N_11542,N_11563);
xnor U13875 (N_13875,N_11771,N_10222);
and U13876 (N_13876,N_11010,N_9838);
or U13877 (N_13877,N_10236,N_9793);
nor U13878 (N_13878,N_10402,N_9137);
nand U13879 (N_13879,N_10809,N_9904);
nand U13880 (N_13880,N_9140,N_10300);
nand U13881 (N_13881,N_11118,N_9057);
and U13882 (N_13882,N_10686,N_11780);
nor U13883 (N_13883,N_10525,N_10342);
or U13884 (N_13884,N_11976,N_10020);
xnor U13885 (N_13885,N_10794,N_9713);
nor U13886 (N_13886,N_9607,N_10912);
and U13887 (N_13887,N_9788,N_9411);
or U13888 (N_13888,N_11931,N_10861);
or U13889 (N_13889,N_11075,N_11780);
or U13890 (N_13890,N_10688,N_9567);
nor U13891 (N_13891,N_10291,N_11470);
xor U13892 (N_13892,N_10001,N_9093);
nor U13893 (N_13893,N_10498,N_10024);
nor U13894 (N_13894,N_10628,N_9723);
and U13895 (N_13895,N_11572,N_11892);
and U13896 (N_13896,N_9465,N_10967);
nand U13897 (N_13897,N_11691,N_11519);
nor U13898 (N_13898,N_10174,N_9412);
and U13899 (N_13899,N_9686,N_11430);
nor U13900 (N_13900,N_11872,N_11562);
xnor U13901 (N_13901,N_10478,N_10486);
or U13902 (N_13902,N_11389,N_10217);
nand U13903 (N_13903,N_11561,N_11152);
nor U13904 (N_13904,N_10699,N_9235);
nand U13905 (N_13905,N_11298,N_11172);
and U13906 (N_13906,N_11005,N_10337);
or U13907 (N_13907,N_9029,N_11812);
nand U13908 (N_13908,N_9488,N_11827);
nor U13909 (N_13909,N_11173,N_9747);
nand U13910 (N_13910,N_9689,N_9516);
and U13911 (N_13911,N_9014,N_9189);
nor U13912 (N_13912,N_11112,N_9019);
or U13913 (N_13913,N_10596,N_9305);
xor U13914 (N_13914,N_10281,N_11867);
xor U13915 (N_13915,N_9757,N_11008);
xnor U13916 (N_13916,N_10066,N_9961);
or U13917 (N_13917,N_11461,N_10734);
nand U13918 (N_13918,N_11325,N_11609);
and U13919 (N_13919,N_11487,N_10345);
nor U13920 (N_13920,N_9242,N_11756);
nand U13921 (N_13921,N_9702,N_9477);
nor U13922 (N_13922,N_10009,N_9053);
xnor U13923 (N_13923,N_11270,N_9752);
nor U13924 (N_13924,N_10766,N_9707);
xor U13925 (N_13925,N_10763,N_11992);
nor U13926 (N_13926,N_9829,N_10832);
and U13927 (N_13927,N_9620,N_11499);
nor U13928 (N_13928,N_9408,N_10352);
or U13929 (N_13929,N_10354,N_11557);
nor U13930 (N_13930,N_10808,N_10076);
nor U13931 (N_13931,N_9000,N_10458);
and U13932 (N_13932,N_10314,N_10740);
and U13933 (N_13933,N_11088,N_10265);
xnor U13934 (N_13934,N_10046,N_11083);
nand U13935 (N_13935,N_9496,N_10246);
xor U13936 (N_13936,N_10886,N_10226);
nand U13937 (N_13937,N_9340,N_10677);
or U13938 (N_13938,N_10035,N_11681);
nor U13939 (N_13939,N_9125,N_10454);
or U13940 (N_13940,N_9485,N_9997);
or U13941 (N_13941,N_10033,N_9123);
and U13942 (N_13942,N_10792,N_10141);
or U13943 (N_13943,N_11305,N_10184);
xnor U13944 (N_13944,N_10612,N_11524);
xnor U13945 (N_13945,N_9744,N_9656);
nand U13946 (N_13946,N_10863,N_11487);
nand U13947 (N_13947,N_11154,N_11940);
nand U13948 (N_13948,N_10195,N_9366);
nor U13949 (N_13949,N_10342,N_10699);
xnor U13950 (N_13950,N_9138,N_9444);
or U13951 (N_13951,N_11856,N_9766);
xor U13952 (N_13952,N_10936,N_10166);
nor U13953 (N_13953,N_9006,N_10619);
nand U13954 (N_13954,N_11981,N_9383);
xnor U13955 (N_13955,N_9362,N_10393);
nand U13956 (N_13956,N_9734,N_9990);
nand U13957 (N_13957,N_11116,N_9663);
and U13958 (N_13958,N_9146,N_10700);
or U13959 (N_13959,N_9518,N_10378);
or U13960 (N_13960,N_10779,N_11143);
xnor U13961 (N_13961,N_9251,N_9503);
nand U13962 (N_13962,N_10772,N_10649);
or U13963 (N_13963,N_11661,N_10480);
nand U13964 (N_13964,N_9716,N_11912);
or U13965 (N_13965,N_9620,N_10951);
nand U13966 (N_13966,N_10982,N_10187);
xnor U13967 (N_13967,N_9575,N_11088);
and U13968 (N_13968,N_10235,N_10008);
xnor U13969 (N_13969,N_11125,N_9179);
nand U13970 (N_13970,N_10095,N_11907);
and U13971 (N_13971,N_11106,N_9604);
or U13972 (N_13972,N_10973,N_10059);
nor U13973 (N_13973,N_10489,N_10527);
or U13974 (N_13974,N_10506,N_11537);
nand U13975 (N_13975,N_11628,N_9842);
and U13976 (N_13976,N_10615,N_11727);
xor U13977 (N_13977,N_9177,N_10614);
and U13978 (N_13978,N_9064,N_9667);
xor U13979 (N_13979,N_11884,N_10251);
xnor U13980 (N_13980,N_10130,N_11232);
and U13981 (N_13981,N_11712,N_9166);
or U13982 (N_13982,N_9470,N_9080);
nor U13983 (N_13983,N_10594,N_10066);
nand U13984 (N_13984,N_11696,N_11021);
and U13985 (N_13985,N_11981,N_10216);
and U13986 (N_13986,N_10843,N_11974);
and U13987 (N_13987,N_11956,N_11535);
nand U13988 (N_13988,N_10517,N_11945);
or U13989 (N_13989,N_9831,N_11069);
or U13990 (N_13990,N_9081,N_10066);
nor U13991 (N_13991,N_10224,N_10578);
and U13992 (N_13992,N_9947,N_11577);
and U13993 (N_13993,N_10579,N_9619);
xor U13994 (N_13994,N_9223,N_9185);
nand U13995 (N_13995,N_11591,N_10782);
xor U13996 (N_13996,N_9962,N_11555);
or U13997 (N_13997,N_11507,N_11567);
nand U13998 (N_13998,N_11504,N_11062);
and U13999 (N_13999,N_9529,N_11424);
nand U14000 (N_14000,N_9906,N_9828);
nand U14001 (N_14001,N_11324,N_9599);
or U14002 (N_14002,N_10411,N_10971);
xnor U14003 (N_14003,N_9838,N_9666);
nor U14004 (N_14004,N_9804,N_11251);
xor U14005 (N_14005,N_10759,N_10780);
nand U14006 (N_14006,N_9164,N_9549);
xnor U14007 (N_14007,N_10347,N_11209);
or U14008 (N_14008,N_10018,N_10842);
and U14009 (N_14009,N_10407,N_11639);
xnor U14010 (N_14010,N_11683,N_10957);
xnor U14011 (N_14011,N_10807,N_11984);
and U14012 (N_14012,N_10514,N_9279);
and U14013 (N_14013,N_10679,N_10664);
xnor U14014 (N_14014,N_10425,N_10922);
nand U14015 (N_14015,N_9471,N_9230);
nand U14016 (N_14016,N_11674,N_10845);
nand U14017 (N_14017,N_11042,N_11099);
xor U14018 (N_14018,N_9561,N_11121);
xnor U14019 (N_14019,N_11707,N_9232);
or U14020 (N_14020,N_10845,N_11360);
or U14021 (N_14021,N_9641,N_10232);
xor U14022 (N_14022,N_9316,N_10230);
and U14023 (N_14023,N_9011,N_11636);
or U14024 (N_14024,N_10715,N_10985);
nand U14025 (N_14025,N_11706,N_11051);
and U14026 (N_14026,N_10164,N_9644);
or U14027 (N_14027,N_10564,N_10382);
or U14028 (N_14028,N_9188,N_11236);
and U14029 (N_14029,N_10166,N_11222);
or U14030 (N_14030,N_10854,N_10544);
and U14031 (N_14031,N_11928,N_10453);
and U14032 (N_14032,N_9745,N_9305);
nor U14033 (N_14033,N_11521,N_9700);
or U14034 (N_14034,N_10538,N_10385);
nand U14035 (N_14035,N_10052,N_10065);
xor U14036 (N_14036,N_9880,N_10718);
xnor U14037 (N_14037,N_10902,N_9313);
xnor U14038 (N_14038,N_9298,N_9565);
nor U14039 (N_14039,N_9035,N_11767);
and U14040 (N_14040,N_11622,N_11340);
nor U14041 (N_14041,N_11729,N_11826);
nand U14042 (N_14042,N_9170,N_9490);
and U14043 (N_14043,N_9167,N_10515);
xnor U14044 (N_14044,N_11067,N_10521);
nand U14045 (N_14045,N_10185,N_10071);
and U14046 (N_14046,N_11417,N_11750);
nand U14047 (N_14047,N_10179,N_9705);
xnor U14048 (N_14048,N_9150,N_11909);
nor U14049 (N_14049,N_10331,N_9688);
nand U14050 (N_14050,N_10002,N_10676);
or U14051 (N_14051,N_9940,N_10702);
xnor U14052 (N_14052,N_9827,N_11307);
or U14053 (N_14053,N_10430,N_9851);
nor U14054 (N_14054,N_9990,N_9516);
or U14055 (N_14055,N_10921,N_11780);
nor U14056 (N_14056,N_10017,N_9936);
xnor U14057 (N_14057,N_9085,N_9393);
or U14058 (N_14058,N_9632,N_10262);
and U14059 (N_14059,N_9815,N_11847);
nor U14060 (N_14060,N_11781,N_9720);
nand U14061 (N_14061,N_10967,N_11831);
nand U14062 (N_14062,N_9566,N_10633);
nand U14063 (N_14063,N_10036,N_10659);
xnor U14064 (N_14064,N_10200,N_10217);
nor U14065 (N_14065,N_9710,N_10271);
and U14066 (N_14066,N_10235,N_10034);
xor U14067 (N_14067,N_10004,N_10729);
nor U14068 (N_14068,N_10588,N_11101);
nor U14069 (N_14069,N_10566,N_9029);
xor U14070 (N_14070,N_11092,N_9667);
and U14071 (N_14071,N_9700,N_11698);
nand U14072 (N_14072,N_10868,N_11991);
nor U14073 (N_14073,N_11050,N_10003);
xnor U14074 (N_14074,N_10366,N_11164);
and U14075 (N_14075,N_10283,N_9645);
and U14076 (N_14076,N_9042,N_11458);
and U14077 (N_14077,N_10191,N_11317);
nand U14078 (N_14078,N_11918,N_9607);
nand U14079 (N_14079,N_11132,N_9412);
xnor U14080 (N_14080,N_10950,N_10305);
and U14081 (N_14081,N_9405,N_10842);
xnor U14082 (N_14082,N_9907,N_11459);
nor U14083 (N_14083,N_10989,N_11363);
xor U14084 (N_14084,N_11061,N_10088);
or U14085 (N_14085,N_9567,N_9511);
and U14086 (N_14086,N_9246,N_10966);
or U14087 (N_14087,N_10600,N_9933);
xnor U14088 (N_14088,N_11734,N_10384);
or U14089 (N_14089,N_11697,N_11695);
nand U14090 (N_14090,N_9135,N_11555);
and U14091 (N_14091,N_9885,N_9483);
or U14092 (N_14092,N_10580,N_9550);
and U14093 (N_14093,N_9748,N_9272);
nand U14094 (N_14094,N_9762,N_9183);
nand U14095 (N_14095,N_10592,N_10893);
and U14096 (N_14096,N_11469,N_10299);
xor U14097 (N_14097,N_9343,N_9995);
nand U14098 (N_14098,N_11799,N_9057);
xnor U14099 (N_14099,N_11423,N_9042);
nor U14100 (N_14100,N_10147,N_11922);
xnor U14101 (N_14101,N_9906,N_10769);
and U14102 (N_14102,N_9327,N_9590);
or U14103 (N_14103,N_10061,N_9155);
nand U14104 (N_14104,N_10985,N_10403);
and U14105 (N_14105,N_10210,N_9887);
and U14106 (N_14106,N_11411,N_9984);
nor U14107 (N_14107,N_10507,N_11447);
and U14108 (N_14108,N_11233,N_9751);
or U14109 (N_14109,N_10754,N_9951);
nand U14110 (N_14110,N_10104,N_11540);
and U14111 (N_14111,N_10750,N_11368);
and U14112 (N_14112,N_11793,N_9137);
xor U14113 (N_14113,N_11228,N_10564);
nand U14114 (N_14114,N_9252,N_9423);
nand U14115 (N_14115,N_11468,N_9165);
nand U14116 (N_14116,N_11080,N_11254);
nand U14117 (N_14117,N_11912,N_9415);
or U14118 (N_14118,N_9174,N_11448);
xnor U14119 (N_14119,N_9681,N_9479);
nand U14120 (N_14120,N_11640,N_9030);
or U14121 (N_14121,N_10379,N_10705);
or U14122 (N_14122,N_9861,N_11521);
nand U14123 (N_14123,N_11579,N_11076);
nor U14124 (N_14124,N_9934,N_9983);
xnor U14125 (N_14125,N_10483,N_9611);
nand U14126 (N_14126,N_11638,N_10505);
xnor U14127 (N_14127,N_11233,N_9193);
nand U14128 (N_14128,N_9196,N_10410);
nor U14129 (N_14129,N_11778,N_11444);
xor U14130 (N_14130,N_9971,N_9384);
nand U14131 (N_14131,N_10743,N_11589);
or U14132 (N_14132,N_9008,N_9622);
and U14133 (N_14133,N_10643,N_10280);
and U14134 (N_14134,N_10672,N_10889);
nor U14135 (N_14135,N_11855,N_10213);
and U14136 (N_14136,N_11925,N_9760);
and U14137 (N_14137,N_10674,N_10988);
or U14138 (N_14138,N_11211,N_11767);
nand U14139 (N_14139,N_9796,N_10211);
or U14140 (N_14140,N_10586,N_11378);
nor U14141 (N_14141,N_11921,N_11021);
nor U14142 (N_14142,N_9047,N_11498);
nand U14143 (N_14143,N_11752,N_11532);
xor U14144 (N_14144,N_11840,N_10328);
xnor U14145 (N_14145,N_11036,N_10355);
xor U14146 (N_14146,N_11357,N_10879);
nor U14147 (N_14147,N_9324,N_9858);
or U14148 (N_14148,N_11745,N_9740);
xor U14149 (N_14149,N_9027,N_10917);
and U14150 (N_14150,N_11920,N_9716);
xnor U14151 (N_14151,N_10115,N_11527);
or U14152 (N_14152,N_10746,N_9435);
nor U14153 (N_14153,N_11890,N_11756);
nor U14154 (N_14154,N_10254,N_11736);
and U14155 (N_14155,N_11640,N_11031);
and U14156 (N_14156,N_10772,N_10391);
and U14157 (N_14157,N_10543,N_9355);
xnor U14158 (N_14158,N_10361,N_9837);
nand U14159 (N_14159,N_10330,N_9779);
and U14160 (N_14160,N_9712,N_11983);
or U14161 (N_14161,N_11121,N_10969);
or U14162 (N_14162,N_10823,N_9499);
or U14163 (N_14163,N_9485,N_9805);
xnor U14164 (N_14164,N_10110,N_10262);
xor U14165 (N_14165,N_10966,N_9938);
nand U14166 (N_14166,N_10742,N_10079);
or U14167 (N_14167,N_11681,N_10719);
or U14168 (N_14168,N_10743,N_9237);
nand U14169 (N_14169,N_9305,N_9803);
xor U14170 (N_14170,N_9234,N_10739);
nor U14171 (N_14171,N_10741,N_10457);
nand U14172 (N_14172,N_11230,N_11682);
nand U14173 (N_14173,N_9976,N_11521);
and U14174 (N_14174,N_10611,N_9835);
nand U14175 (N_14175,N_11507,N_11154);
nor U14176 (N_14176,N_9876,N_11480);
xor U14177 (N_14177,N_10240,N_10755);
nor U14178 (N_14178,N_9983,N_11345);
xnor U14179 (N_14179,N_11625,N_9436);
or U14180 (N_14180,N_10331,N_9309);
nand U14181 (N_14181,N_9676,N_11522);
nor U14182 (N_14182,N_10247,N_9966);
or U14183 (N_14183,N_10041,N_9904);
and U14184 (N_14184,N_10648,N_9483);
or U14185 (N_14185,N_10372,N_10819);
and U14186 (N_14186,N_9924,N_11076);
nand U14187 (N_14187,N_9386,N_11601);
nor U14188 (N_14188,N_10225,N_11820);
and U14189 (N_14189,N_9773,N_11641);
and U14190 (N_14190,N_10175,N_11638);
nand U14191 (N_14191,N_9159,N_10817);
or U14192 (N_14192,N_11531,N_10806);
nor U14193 (N_14193,N_10391,N_9147);
nor U14194 (N_14194,N_11024,N_11599);
nand U14195 (N_14195,N_9201,N_10617);
xor U14196 (N_14196,N_9347,N_11605);
xor U14197 (N_14197,N_10511,N_9953);
nor U14198 (N_14198,N_11317,N_11341);
or U14199 (N_14199,N_10538,N_10388);
xor U14200 (N_14200,N_9581,N_10334);
xor U14201 (N_14201,N_11869,N_9532);
nand U14202 (N_14202,N_10413,N_9966);
nand U14203 (N_14203,N_9605,N_10033);
nor U14204 (N_14204,N_10274,N_10680);
xor U14205 (N_14205,N_11872,N_11498);
and U14206 (N_14206,N_10404,N_11542);
nor U14207 (N_14207,N_10501,N_11733);
xor U14208 (N_14208,N_11520,N_11122);
nor U14209 (N_14209,N_11336,N_11350);
or U14210 (N_14210,N_11154,N_10753);
or U14211 (N_14211,N_9742,N_10104);
nor U14212 (N_14212,N_10598,N_9319);
xor U14213 (N_14213,N_10228,N_10283);
and U14214 (N_14214,N_11821,N_9916);
nand U14215 (N_14215,N_10217,N_9972);
or U14216 (N_14216,N_10388,N_9362);
xor U14217 (N_14217,N_11355,N_9542);
nor U14218 (N_14218,N_10824,N_10916);
nand U14219 (N_14219,N_9604,N_10267);
and U14220 (N_14220,N_10048,N_11794);
xnor U14221 (N_14221,N_11742,N_10688);
and U14222 (N_14222,N_10825,N_11975);
nand U14223 (N_14223,N_10361,N_11134);
xnor U14224 (N_14224,N_10818,N_9268);
nand U14225 (N_14225,N_11427,N_9390);
xor U14226 (N_14226,N_11734,N_11109);
nor U14227 (N_14227,N_10905,N_11457);
xnor U14228 (N_14228,N_9804,N_11223);
nor U14229 (N_14229,N_11585,N_10168);
nand U14230 (N_14230,N_10539,N_9329);
and U14231 (N_14231,N_11172,N_11557);
nor U14232 (N_14232,N_9020,N_10246);
xor U14233 (N_14233,N_11449,N_10292);
nor U14234 (N_14234,N_9696,N_9674);
nor U14235 (N_14235,N_9952,N_9391);
nand U14236 (N_14236,N_11305,N_10515);
xnor U14237 (N_14237,N_10206,N_9358);
or U14238 (N_14238,N_10626,N_9021);
nor U14239 (N_14239,N_9370,N_9708);
and U14240 (N_14240,N_9426,N_11114);
or U14241 (N_14241,N_10598,N_10637);
nor U14242 (N_14242,N_9825,N_10142);
nor U14243 (N_14243,N_9614,N_9674);
nor U14244 (N_14244,N_9350,N_9459);
nor U14245 (N_14245,N_11694,N_10364);
nand U14246 (N_14246,N_9184,N_9660);
xor U14247 (N_14247,N_10465,N_11401);
and U14248 (N_14248,N_9827,N_11206);
or U14249 (N_14249,N_10927,N_9096);
nand U14250 (N_14250,N_10955,N_9467);
or U14251 (N_14251,N_9865,N_9284);
or U14252 (N_14252,N_11889,N_11455);
and U14253 (N_14253,N_11932,N_9747);
nor U14254 (N_14254,N_10753,N_9626);
nand U14255 (N_14255,N_11007,N_11589);
or U14256 (N_14256,N_10551,N_10393);
or U14257 (N_14257,N_11476,N_11705);
and U14258 (N_14258,N_10166,N_9531);
and U14259 (N_14259,N_10107,N_10661);
xnor U14260 (N_14260,N_11454,N_9778);
and U14261 (N_14261,N_11436,N_9611);
nor U14262 (N_14262,N_11811,N_9458);
nor U14263 (N_14263,N_10110,N_11068);
or U14264 (N_14264,N_9553,N_9117);
and U14265 (N_14265,N_9566,N_9345);
and U14266 (N_14266,N_11666,N_11891);
and U14267 (N_14267,N_11595,N_10873);
nor U14268 (N_14268,N_9965,N_10360);
and U14269 (N_14269,N_9521,N_10821);
nor U14270 (N_14270,N_11570,N_11599);
or U14271 (N_14271,N_11138,N_11695);
or U14272 (N_14272,N_11900,N_9398);
nor U14273 (N_14273,N_10969,N_10852);
xnor U14274 (N_14274,N_9605,N_10142);
nor U14275 (N_14275,N_9644,N_9457);
or U14276 (N_14276,N_11383,N_10543);
nor U14277 (N_14277,N_9688,N_10180);
xnor U14278 (N_14278,N_10560,N_9239);
xor U14279 (N_14279,N_9147,N_10530);
nand U14280 (N_14280,N_11297,N_10968);
or U14281 (N_14281,N_10015,N_10387);
or U14282 (N_14282,N_9997,N_10245);
nand U14283 (N_14283,N_11263,N_11764);
xor U14284 (N_14284,N_9802,N_9702);
xnor U14285 (N_14285,N_10618,N_11056);
and U14286 (N_14286,N_10353,N_10732);
xnor U14287 (N_14287,N_9522,N_11090);
and U14288 (N_14288,N_11669,N_10304);
and U14289 (N_14289,N_9365,N_11068);
xnor U14290 (N_14290,N_11855,N_11471);
nand U14291 (N_14291,N_10845,N_9512);
or U14292 (N_14292,N_11158,N_9851);
or U14293 (N_14293,N_10675,N_11661);
and U14294 (N_14294,N_10610,N_11173);
or U14295 (N_14295,N_11571,N_10838);
and U14296 (N_14296,N_11372,N_10012);
nor U14297 (N_14297,N_9816,N_11286);
nand U14298 (N_14298,N_11518,N_10441);
and U14299 (N_14299,N_10705,N_9559);
xnor U14300 (N_14300,N_11357,N_9763);
and U14301 (N_14301,N_9341,N_11788);
nor U14302 (N_14302,N_10467,N_9905);
nand U14303 (N_14303,N_9740,N_9652);
and U14304 (N_14304,N_10727,N_9007);
nand U14305 (N_14305,N_11975,N_10042);
nand U14306 (N_14306,N_11345,N_9857);
nor U14307 (N_14307,N_10498,N_9625);
nor U14308 (N_14308,N_11308,N_9044);
or U14309 (N_14309,N_10874,N_9489);
and U14310 (N_14310,N_11446,N_11631);
xor U14311 (N_14311,N_9294,N_10274);
nor U14312 (N_14312,N_9501,N_10797);
or U14313 (N_14313,N_11049,N_9980);
nand U14314 (N_14314,N_11636,N_10986);
nor U14315 (N_14315,N_11457,N_9714);
and U14316 (N_14316,N_10359,N_9534);
xnor U14317 (N_14317,N_10176,N_9526);
nand U14318 (N_14318,N_9835,N_10342);
and U14319 (N_14319,N_11509,N_9945);
xor U14320 (N_14320,N_11588,N_9229);
xor U14321 (N_14321,N_11432,N_10780);
nor U14322 (N_14322,N_11725,N_9532);
and U14323 (N_14323,N_9824,N_11971);
and U14324 (N_14324,N_9550,N_9519);
and U14325 (N_14325,N_9678,N_9887);
or U14326 (N_14326,N_10230,N_10018);
or U14327 (N_14327,N_10259,N_9651);
or U14328 (N_14328,N_10144,N_9406);
or U14329 (N_14329,N_11307,N_9723);
xnor U14330 (N_14330,N_10141,N_11472);
and U14331 (N_14331,N_9148,N_9398);
and U14332 (N_14332,N_10685,N_10279);
xnor U14333 (N_14333,N_10276,N_11008);
or U14334 (N_14334,N_10570,N_9887);
or U14335 (N_14335,N_9493,N_9379);
and U14336 (N_14336,N_11006,N_10859);
xnor U14337 (N_14337,N_10853,N_10740);
nor U14338 (N_14338,N_11850,N_9094);
and U14339 (N_14339,N_9319,N_9529);
xnor U14340 (N_14340,N_11045,N_10368);
xor U14341 (N_14341,N_11104,N_10872);
xor U14342 (N_14342,N_10907,N_11414);
or U14343 (N_14343,N_10306,N_11976);
xor U14344 (N_14344,N_10843,N_11695);
or U14345 (N_14345,N_9738,N_9128);
xor U14346 (N_14346,N_10780,N_10882);
nand U14347 (N_14347,N_10237,N_10911);
or U14348 (N_14348,N_10793,N_9452);
and U14349 (N_14349,N_10019,N_9416);
xnor U14350 (N_14350,N_10850,N_11870);
nand U14351 (N_14351,N_10071,N_10326);
and U14352 (N_14352,N_10691,N_10579);
nor U14353 (N_14353,N_10033,N_11545);
or U14354 (N_14354,N_11193,N_9619);
and U14355 (N_14355,N_9777,N_10512);
nor U14356 (N_14356,N_11529,N_11872);
and U14357 (N_14357,N_9009,N_11810);
xor U14358 (N_14358,N_11412,N_9577);
or U14359 (N_14359,N_11012,N_11301);
and U14360 (N_14360,N_11131,N_11066);
nor U14361 (N_14361,N_10973,N_10423);
nand U14362 (N_14362,N_11228,N_9370);
nand U14363 (N_14363,N_10064,N_10112);
xor U14364 (N_14364,N_11363,N_11727);
nor U14365 (N_14365,N_11484,N_11380);
or U14366 (N_14366,N_9812,N_11686);
nor U14367 (N_14367,N_9383,N_11652);
nand U14368 (N_14368,N_9806,N_9192);
nor U14369 (N_14369,N_10729,N_10290);
nor U14370 (N_14370,N_9694,N_10371);
and U14371 (N_14371,N_11713,N_9469);
or U14372 (N_14372,N_10257,N_9880);
nand U14373 (N_14373,N_11774,N_9746);
nor U14374 (N_14374,N_11878,N_10876);
nor U14375 (N_14375,N_10274,N_10861);
nand U14376 (N_14376,N_10737,N_11407);
and U14377 (N_14377,N_10262,N_11033);
nor U14378 (N_14378,N_11873,N_10251);
and U14379 (N_14379,N_11127,N_9465);
nand U14380 (N_14380,N_11770,N_11627);
and U14381 (N_14381,N_9027,N_10109);
nand U14382 (N_14382,N_9025,N_10224);
and U14383 (N_14383,N_10428,N_9973);
nor U14384 (N_14384,N_11635,N_10774);
nor U14385 (N_14385,N_10522,N_9804);
nand U14386 (N_14386,N_10858,N_10820);
nand U14387 (N_14387,N_11209,N_11778);
nor U14388 (N_14388,N_10074,N_9257);
xnor U14389 (N_14389,N_10694,N_9847);
or U14390 (N_14390,N_10940,N_10368);
and U14391 (N_14391,N_9560,N_9145);
xnor U14392 (N_14392,N_9695,N_9005);
nor U14393 (N_14393,N_11664,N_11365);
nand U14394 (N_14394,N_10083,N_10127);
and U14395 (N_14395,N_9060,N_11172);
or U14396 (N_14396,N_10455,N_11675);
nor U14397 (N_14397,N_11144,N_9223);
and U14398 (N_14398,N_11209,N_9027);
xor U14399 (N_14399,N_9946,N_9383);
nand U14400 (N_14400,N_11791,N_11216);
and U14401 (N_14401,N_11052,N_11604);
and U14402 (N_14402,N_9531,N_9846);
nand U14403 (N_14403,N_11430,N_11740);
nor U14404 (N_14404,N_10524,N_11592);
nand U14405 (N_14405,N_11435,N_9764);
xor U14406 (N_14406,N_10683,N_10132);
xnor U14407 (N_14407,N_11927,N_9365);
nand U14408 (N_14408,N_9270,N_10845);
or U14409 (N_14409,N_10601,N_11319);
and U14410 (N_14410,N_11564,N_10021);
nand U14411 (N_14411,N_10190,N_11355);
nor U14412 (N_14412,N_10306,N_11285);
xnor U14413 (N_14413,N_11300,N_11830);
nor U14414 (N_14414,N_10742,N_9952);
xnor U14415 (N_14415,N_9076,N_10707);
xor U14416 (N_14416,N_9924,N_9585);
nand U14417 (N_14417,N_11723,N_10616);
nand U14418 (N_14418,N_10224,N_9351);
nand U14419 (N_14419,N_11656,N_9421);
nor U14420 (N_14420,N_10091,N_11119);
nor U14421 (N_14421,N_11861,N_10431);
xnor U14422 (N_14422,N_9723,N_9679);
xnor U14423 (N_14423,N_9820,N_9124);
and U14424 (N_14424,N_10252,N_9322);
or U14425 (N_14425,N_11008,N_11790);
or U14426 (N_14426,N_11881,N_11279);
and U14427 (N_14427,N_9934,N_9490);
nand U14428 (N_14428,N_10966,N_11770);
or U14429 (N_14429,N_11380,N_11893);
nand U14430 (N_14430,N_9195,N_11196);
xor U14431 (N_14431,N_10154,N_10409);
xor U14432 (N_14432,N_10909,N_10723);
or U14433 (N_14433,N_11476,N_10717);
xor U14434 (N_14434,N_11363,N_9139);
nand U14435 (N_14435,N_9389,N_10858);
nand U14436 (N_14436,N_11305,N_9802);
nand U14437 (N_14437,N_11651,N_9656);
nor U14438 (N_14438,N_9619,N_11911);
xor U14439 (N_14439,N_9693,N_11919);
or U14440 (N_14440,N_11120,N_9568);
nor U14441 (N_14441,N_9588,N_9661);
or U14442 (N_14442,N_9467,N_10516);
and U14443 (N_14443,N_9865,N_10328);
and U14444 (N_14444,N_10305,N_11216);
xor U14445 (N_14445,N_11482,N_11925);
nor U14446 (N_14446,N_10017,N_10117);
nor U14447 (N_14447,N_9294,N_9816);
or U14448 (N_14448,N_10181,N_10992);
or U14449 (N_14449,N_11898,N_9111);
nand U14450 (N_14450,N_11776,N_9861);
nor U14451 (N_14451,N_11579,N_11389);
nand U14452 (N_14452,N_9350,N_11422);
nand U14453 (N_14453,N_9855,N_11421);
nand U14454 (N_14454,N_9574,N_9925);
xnor U14455 (N_14455,N_9773,N_10683);
nand U14456 (N_14456,N_11565,N_9918);
xnor U14457 (N_14457,N_10617,N_11981);
nor U14458 (N_14458,N_9310,N_10496);
or U14459 (N_14459,N_10177,N_11251);
and U14460 (N_14460,N_11257,N_11695);
nor U14461 (N_14461,N_11141,N_10174);
and U14462 (N_14462,N_10541,N_10459);
xnor U14463 (N_14463,N_10349,N_10231);
xnor U14464 (N_14464,N_11727,N_11176);
nor U14465 (N_14465,N_10115,N_10509);
and U14466 (N_14466,N_11252,N_11622);
and U14467 (N_14467,N_9312,N_9411);
or U14468 (N_14468,N_11207,N_10965);
or U14469 (N_14469,N_11021,N_9454);
nand U14470 (N_14470,N_9715,N_11558);
nor U14471 (N_14471,N_9635,N_11948);
or U14472 (N_14472,N_10834,N_10645);
xnor U14473 (N_14473,N_9314,N_9379);
nor U14474 (N_14474,N_11233,N_10395);
xor U14475 (N_14475,N_10623,N_9388);
xor U14476 (N_14476,N_9503,N_11375);
or U14477 (N_14477,N_11264,N_9193);
xnor U14478 (N_14478,N_10711,N_9196);
xor U14479 (N_14479,N_11351,N_10581);
nand U14480 (N_14480,N_10576,N_11449);
and U14481 (N_14481,N_9347,N_11993);
and U14482 (N_14482,N_11829,N_11383);
xnor U14483 (N_14483,N_11236,N_10155);
nor U14484 (N_14484,N_11983,N_11113);
nand U14485 (N_14485,N_11432,N_10481);
nand U14486 (N_14486,N_9731,N_10442);
nor U14487 (N_14487,N_9227,N_9637);
nor U14488 (N_14488,N_10201,N_10942);
nand U14489 (N_14489,N_10910,N_10930);
nor U14490 (N_14490,N_10518,N_9118);
nand U14491 (N_14491,N_11676,N_11045);
nand U14492 (N_14492,N_11203,N_9113);
and U14493 (N_14493,N_10820,N_9176);
nand U14494 (N_14494,N_9811,N_10661);
xor U14495 (N_14495,N_10491,N_9091);
or U14496 (N_14496,N_9278,N_9096);
xnor U14497 (N_14497,N_9214,N_10776);
nand U14498 (N_14498,N_9269,N_9463);
nand U14499 (N_14499,N_9848,N_9140);
nand U14500 (N_14500,N_9472,N_10783);
nor U14501 (N_14501,N_11872,N_9295);
nand U14502 (N_14502,N_10369,N_11417);
and U14503 (N_14503,N_9194,N_9943);
xnor U14504 (N_14504,N_11557,N_11598);
and U14505 (N_14505,N_10049,N_9930);
nor U14506 (N_14506,N_9778,N_11393);
and U14507 (N_14507,N_11450,N_9685);
nor U14508 (N_14508,N_10858,N_9390);
nor U14509 (N_14509,N_9326,N_9877);
xor U14510 (N_14510,N_9860,N_11463);
nand U14511 (N_14511,N_11729,N_10514);
and U14512 (N_14512,N_9977,N_10686);
and U14513 (N_14513,N_10316,N_11379);
or U14514 (N_14514,N_11822,N_11846);
xnor U14515 (N_14515,N_11987,N_9265);
or U14516 (N_14516,N_11202,N_9140);
nand U14517 (N_14517,N_10035,N_9512);
and U14518 (N_14518,N_10604,N_9664);
xnor U14519 (N_14519,N_10722,N_11901);
and U14520 (N_14520,N_9897,N_11282);
nand U14521 (N_14521,N_9405,N_10912);
nand U14522 (N_14522,N_10987,N_10278);
or U14523 (N_14523,N_10145,N_9345);
nor U14524 (N_14524,N_9099,N_10711);
and U14525 (N_14525,N_11353,N_9058);
or U14526 (N_14526,N_10566,N_11989);
or U14527 (N_14527,N_10254,N_11437);
nor U14528 (N_14528,N_9920,N_10939);
xnor U14529 (N_14529,N_11304,N_11003);
or U14530 (N_14530,N_10694,N_11306);
xor U14531 (N_14531,N_9083,N_10089);
xnor U14532 (N_14532,N_11347,N_11139);
and U14533 (N_14533,N_10188,N_9204);
and U14534 (N_14534,N_10800,N_11625);
nand U14535 (N_14535,N_9128,N_10752);
xnor U14536 (N_14536,N_11781,N_11127);
xnor U14537 (N_14537,N_10226,N_11219);
or U14538 (N_14538,N_10559,N_11973);
nand U14539 (N_14539,N_11123,N_10420);
xnor U14540 (N_14540,N_11636,N_11129);
and U14541 (N_14541,N_10322,N_10379);
nand U14542 (N_14542,N_10749,N_11364);
nor U14543 (N_14543,N_10811,N_10356);
nand U14544 (N_14544,N_11961,N_10585);
and U14545 (N_14545,N_9743,N_10691);
and U14546 (N_14546,N_9771,N_11284);
or U14547 (N_14547,N_9713,N_10529);
xor U14548 (N_14548,N_9119,N_9870);
and U14549 (N_14549,N_10973,N_11154);
or U14550 (N_14550,N_11942,N_11688);
xnor U14551 (N_14551,N_9202,N_10892);
or U14552 (N_14552,N_9619,N_9329);
and U14553 (N_14553,N_10717,N_10125);
nand U14554 (N_14554,N_11422,N_11406);
nor U14555 (N_14555,N_10760,N_11429);
or U14556 (N_14556,N_11847,N_10205);
xor U14557 (N_14557,N_11015,N_9640);
xor U14558 (N_14558,N_10222,N_10411);
nand U14559 (N_14559,N_10113,N_11141);
and U14560 (N_14560,N_11089,N_11043);
or U14561 (N_14561,N_10107,N_10042);
nor U14562 (N_14562,N_10546,N_10699);
and U14563 (N_14563,N_11241,N_9789);
and U14564 (N_14564,N_9632,N_9925);
nand U14565 (N_14565,N_11060,N_11479);
nand U14566 (N_14566,N_11081,N_9789);
and U14567 (N_14567,N_10747,N_10347);
or U14568 (N_14568,N_10849,N_11546);
xnor U14569 (N_14569,N_9147,N_10086);
xnor U14570 (N_14570,N_11860,N_10835);
xor U14571 (N_14571,N_9036,N_10490);
nor U14572 (N_14572,N_10139,N_10215);
nor U14573 (N_14573,N_11704,N_9014);
nand U14574 (N_14574,N_9660,N_11998);
nand U14575 (N_14575,N_9893,N_11860);
nor U14576 (N_14576,N_11444,N_11705);
xor U14577 (N_14577,N_10412,N_9866);
or U14578 (N_14578,N_11056,N_9245);
nand U14579 (N_14579,N_11602,N_10477);
nand U14580 (N_14580,N_11901,N_10435);
nor U14581 (N_14581,N_9317,N_9385);
and U14582 (N_14582,N_10144,N_10725);
and U14583 (N_14583,N_9052,N_10102);
and U14584 (N_14584,N_11168,N_9683);
or U14585 (N_14585,N_10960,N_10204);
or U14586 (N_14586,N_9997,N_10592);
xnor U14587 (N_14587,N_11456,N_11005);
xnor U14588 (N_14588,N_10583,N_9242);
nand U14589 (N_14589,N_11398,N_10563);
and U14590 (N_14590,N_11255,N_11624);
and U14591 (N_14591,N_9585,N_11081);
and U14592 (N_14592,N_10346,N_10089);
or U14593 (N_14593,N_9506,N_10826);
nor U14594 (N_14594,N_10828,N_11270);
or U14595 (N_14595,N_9864,N_10612);
xor U14596 (N_14596,N_10021,N_10450);
or U14597 (N_14597,N_10623,N_10539);
nand U14598 (N_14598,N_10543,N_11755);
and U14599 (N_14599,N_10731,N_9403);
or U14600 (N_14600,N_11048,N_11944);
and U14601 (N_14601,N_9509,N_11892);
or U14602 (N_14602,N_10471,N_11366);
or U14603 (N_14603,N_10770,N_9564);
and U14604 (N_14604,N_10496,N_11926);
or U14605 (N_14605,N_11309,N_11742);
nor U14606 (N_14606,N_10497,N_9220);
xnor U14607 (N_14607,N_9917,N_9196);
nor U14608 (N_14608,N_10590,N_9430);
xnor U14609 (N_14609,N_9577,N_11729);
nor U14610 (N_14610,N_10363,N_10580);
xor U14611 (N_14611,N_10214,N_9619);
nor U14612 (N_14612,N_10109,N_10290);
or U14613 (N_14613,N_10534,N_9843);
xor U14614 (N_14614,N_10424,N_10944);
or U14615 (N_14615,N_9162,N_11122);
or U14616 (N_14616,N_10118,N_11951);
and U14617 (N_14617,N_9260,N_10397);
or U14618 (N_14618,N_10184,N_10511);
nand U14619 (N_14619,N_11429,N_11364);
xnor U14620 (N_14620,N_11039,N_9844);
nor U14621 (N_14621,N_10528,N_11324);
nand U14622 (N_14622,N_11186,N_9828);
or U14623 (N_14623,N_10025,N_11769);
xnor U14624 (N_14624,N_11472,N_9505);
xnor U14625 (N_14625,N_9604,N_11249);
or U14626 (N_14626,N_9699,N_10204);
xor U14627 (N_14627,N_9368,N_10254);
or U14628 (N_14628,N_10465,N_9417);
xor U14629 (N_14629,N_10609,N_11767);
nor U14630 (N_14630,N_10684,N_9816);
or U14631 (N_14631,N_11611,N_11403);
nor U14632 (N_14632,N_11673,N_9708);
xnor U14633 (N_14633,N_11133,N_11571);
or U14634 (N_14634,N_11831,N_10209);
and U14635 (N_14635,N_11772,N_10001);
xnor U14636 (N_14636,N_10728,N_9962);
nand U14637 (N_14637,N_9596,N_11575);
nor U14638 (N_14638,N_11244,N_10000);
or U14639 (N_14639,N_10402,N_11597);
nor U14640 (N_14640,N_9950,N_11504);
nand U14641 (N_14641,N_9214,N_11153);
nor U14642 (N_14642,N_11668,N_9130);
nor U14643 (N_14643,N_9196,N_11648);
xnor U14644 (N_14644,N_10337,N_11740);
nand U14645 (N_14645,N_10807,N_9622);
xnor U14646 (N_14646,N_11112,N_10406);
nor U14647 (N_14647,N_11409,N_11791);
or U14648 (N_14648,N_11090,N_11128);
or U14649 (N_14649,N_9164,N_10825);
or U14650 (N_14650,N_11481,N_11965);
nor U14651 (N_14651,N_9410,N_10365);
and U14652 (N_14652,N_11682,N_9206);
nand U14653 (N_14653,N_10354,N_10975);
nor U14654 (N_14654,N_10364,N_10687);
nand U14655 (N_14655,N_11214,N_9096);
xnor U14656 (N_14656,N_9238,N_9183);
nor U14657 (N_14657,N_9751,N_10331);
and U14658 (N_14658,N_9361,N_10598);
xor U14659 (N_14659,N_11938,N_10567);
or U14660 (N_14660,N_10201,N_11731);
nand U14661 (N_14661,N_9180,N_11215);
and U14662 (N_14662,N_11521,N_9800);
nand U14663 (N_14663,N_10977,N_10480);
and U14664 (N_14664,N_9311,N_9618);
nand U14665 (N_14665,N_9292,N_9937);
or U14666 (N_14666,N_9411,N_10237);
and U14667 (N_14667,N_11328,N_10075);
xnor U14668 (N_14668,N_11494,N_10596);
xor U14669 (N_14669,N_9650,N_11562);
and U14670 (N_14670,N_11998,N_9372);
xnor U14671 (N_14671,N_10916,N_11607);
nor U14672 (N_14672,N_11709,N_11508);
xor U14673 (N_14673,N_9309,N_11986);
xnor U14674 (N_14674,N_9366,N_9372);
and U14675 (N_14675,N_9014,N_9052);
and U14676 (N_14676,N_11541,N_11520);
or U14677 (N_14677,N_11683,N_11953);
or U14678 (N_14678,N_11602,N_9812);
or U14679 (N_14679,N_11831,N_11903);
nor U14680 (N_14680,N_11003,N_9535);
xnor U14681 (N_14681,N_9656,N_10363);
and U14682 (N_14682,N_11233,N_11752);
nor U14683 (N_14683,N_11087,N_9190);
and U14684 (N_14684,N_11401,N_9277);
xnor U14685 (N_14685,N_11086,N_9397);
nor U14686 (N_14686,N_11333,N_10920);
or U14687 (N_14687,N_10264,N_10855);
nor U14688 (N_14688,N_10617,N_9715);
nor U14689 (N_14689,N_11839,N_11788);
xnor U14690 (N_14690,N_11630,N_11650);
nor U14691 (N_14691,N_11784,N_10452);
or U14692 (N_14692,N_10700,N_9826);
nand U14693 (N_14693,N_10512,N_11919);
xnor U14694 (N_14694,N_11610,N_11107);
and U14695 (N_14695,N_11115,N_9838);
or U14696 (N_14696,N_9939,N_9168);
or U14697 (N_14697,N_11471,N_10541);
and U14698 (N_14698,N_11038,N_10435);
nand U14699 (N_14699,N_10078,N_11949);
or U14700 (N_14700,N_10731,N_11687);
xnor U14701 (N_14701,N_10852,N_9805);
or U14702 (N_14702,N_10718,N_10305);
and U14703 (N_14703,N_10461,N_10588);
and U14704 (N_14704,N_9354,N_10510);
nand U14705 (N_14705,N_11700,N_10817);
xnor U14706 (N_14706,N_11419,N_10237);
and U14707 (N_14707,N_11309,N_9242);
and U14708 (N_14708,N_9325,N_9463);
and U14709 (N_14709,N_11354,N_9025);
xor U14710 (N_14710,N_10723,N_9466);
nor U14711 (N_14711,N_9493,N_9153);
xor U14712 (N_14712,N_10207,N_9551);
xor U14713 (N_14713,N_9565,N_10185);
and U14714 (N_14714,N_9475,N_9733);
nor U14715 (N_14715,N_11773,N_9234);
nor U14716 (N_14716,N_10975,N_9775);
nor U14717 (N_14717,N_9055,N_10502);
nand U14718 (N_14718,N_11636,N_9995);
nor U14719 (N_14719,N_9034,N_11020);
or U14720 (N_14720,N_11866,N_11912);
xnor U14721 (N_14721,N_10151,N_9443);
nor U14722 (N_14722,N_10119,N_9222);
or U14723 (N_14723,N_11277,N_10072);
nor U14724 (N_14724,N_9527,N_10335);
or U14725 (N_14725,N_10682,N_11321);
xor U14726 (N_14726,N_11781,N_10145);
nand U14727 (N_14727,N_10302,N_10130);
and U14728 (N_14728,N_9740,N_10438);
nor U14729 (N_14729,N_11290,N_11220);
and U14730 (N_14730,N_9831,N_11530);
and U14731 (N_14731,N_10296,N_9933);
or U14732 (N_14732,N_10393,N_10179);
xor U14733 (N_14733,N_10651,N_10285);
nor U14734 (N_14734,N_11934,N_10724);
nand U14735 (N_14735,N_11841,N_10851);
nor U14736 (N_14736,N_11488,N_10358);
xnor U14737 (N_14737,N_11285,N_9565);
nand U14738 (N_14738,N_9832,N_11471);
xor U14739 (N_14739,N_10253,N_10963);
xnor U14740 (N_14740,N_11897,N_10489);
or U14741 (N_14741,N_9456,N_11434);
or U14742 (N_14742,N_9896,N_9904);
xor U14743 (N_14743,N_10561,N_9311);
nor U14744 (N_14744,N_9788,N_9262);
nand U14745 (N_14745,N_11849,N_9249);
or U14746 (N_14746,N_9169,N_11970);
nor U14747 (N_14747,N_11233,N_9705);
nor U14748 (N_14748,N_10883,N_10250);
nor U14749 (N_14749,N_11840,N_9658);
and U14750 (N_14750,N_10847,N_11424);
nand U14751 (N_14751,N_10826,N_11998);
xnor U14752 (N_14752,N_9345,N_11504);
xor U14753 (N_14753,N_10345,N_10038);
nor U14754 (N_14754,N_10047,N_9754);
nor U14755 (N_14755,N_9213,N_9968);
nand U14756 (N_14756,N_9936,N_11084);
nand U14757 (N_14757,N_9780,N_11983);
nor U14758 (N_14758,N_11464,N_11386);
nand U14759 (N_14759,N_10334,N_11591);
and U14760 (N_14760,N_11356,N_10469);
nor U14761 (N_14761,N_11865,N_10066);
nand U14762 (N_14762,N_9560,N_10725);
or U14763 (N_14763,N_10348,N_11918);
nand U14764 (N_14764,N_9661,N_11320);
xor U14765 (N_14765,N_9714,N_9841);
xor U14766 (N_14766,N_9733,N_11537);
or U14767 (N_14767,N_9761,N_10523);
xor U14768 (N_14768,N_9144,N_11907);
or U14769 (N_14769,N_9847,N_10863);
xor U14770 (N_14770,N_9979,N_11171);
nor U14771 (N_14771,N_11724,N_11790);
xnor U14772 (N_14772,N_9584,N_10834);
nor U14773 (N_14773,N_10713,N_11398);
nor U14774 (N_14774,N_9031,N_10443);
and U14775 (N_14775,N_9224,N_10295);
nand U14776 (N_14776,N_10986,N_9879);
xor U14777 (N_14777,N_10700,N_9443);
or U14778 (N_14778,N_10381,N_9574);
or U14779 (N_14779,N_10348,N_9330);
or U14780 (N_14780,N_10513,N_11714);
or U14781 (N_14781,N_10971,N_11705);
or U14782 (N_14782,N_10215,N_11482);
or U14783 (N_14783,N_11391,N_11304);
nand U14784 (N_14784,N_10343,N_11755);
or U14785 (N_14785,N_10269,N_10871);
xor U14786 (N_14786,N_9745,N_9275);
nand U14787 (N_14787,N_11505,N_11331);
or U14788 (N_14788,N_10180,N_11042);
nand U14789 (N_14789,N_10975,N_11762);
or U14790 (N_14790,N_10754,N_11551);
and U14791 (N_14791,N_11907,N_9275);
or U14792 (N_14792,N_9293,N_11373);
or U14793 (N_14793,N_10136,N_11947);
nand U14794 (N_14794,N_9274,N_11576);
xor U14795 (N_14795,N_10965,N_9586);
or U14796 (N_14796,N_10054,N_11023);
and U14797 (N_14797,N_11082,N_11766);
nand U14798 (N_14798,N_9142,N_11943);
and U14799 (N_14799,N_10965,N_11396);
or U14800 (N_14800,N_11738,N_9038);
xnor U14801 (N_14801,N_9757,N_11400);
nand U14802 (N_14802,N_9467,N_9126);
or U14803 (N_14803,N_11154,N_9673);
nand U14804 (N_14804,N_11242,N_9036);
nand U14805 (N_14805,N_11871,N_9510);
nor U14806 (N_14806,N_11580,N_10696);
xor U14807 (N_14807,N_10674,N_11169);
nor U14808 (N_14808,N_10451,N_9934);
nand U14809 (N_14809,N_10630,N_10446);
and U14810 (N_14810,N_9665,N_9988);
or U14811 (N_14811,N_9972,N_11023);
and U14812 (N_14812,N_11685,N_9192);
nand U14813 (N_14813,N_11892,N_9071);
nand U14814 (N_14814,N_11867,N_9661);
nor U14815 (N_14815,N_10886,N_11946);
or U14816 (N_14816,N_9159,N_10269);
and U14817 (N_14817,N_10558,N_9233);
xor U14818 (N_14818,N_9208,N_11814);
nand U14819 (N_14819,N_11752,N_10852);
nand U14820 (N_14820,N_9098,N_10750);
xnor U14821 (N_14821,N_9740,N_10587);
nor U14822 (N_14822,N_9545,N_9823);
xor U14823 (N_14823,N_11002,N_9445);
and U14824 (N_14824,N_11574,N_10987);
nand U14825 (N_14825,N_11766,N_10977);
and U14826 (N_14826,N_11654,N_10362);
or U14827 (N_14827,N_10834,N_9508);
nand U14828 (N_14828,N_10270,N_10347);
nand U14829 (N_14829,N_9286,N_11173);
xor U14830 (N_14830,N_11493,N_10531);
or U14831 (N_14831,N_10276,N_10661);
or U14832 (N_14832,N_9546,N_9974);
nor U14833 (N_14833,N_9901,N_11642);
or U14834 (N_14834,N_10892,N_10302);
xnor U14835 (N_14835,N_10444,N_9868);
xor U14836 (N_14836,N_10376,N_10561);
and U14837 (N_14837,N_10386,N_9426);
or U14838 (N_14838,N_10534,N_9854);
or U14839 (N_14839,N_9784,N_10800);
nand U14840 (N_14840,N_11259,N_11135);
nand U14841 (N_14841,N_9471,N_9830);
or U14842 (N_14842,N_10137,N_11366);
or U14843 (N_14843,N_9959,N_10045);
nand U14844 (N_14844,N_11288,N_11744);
and U14845 (N_14845,N_10345,N_10477);
and U14846 (N_14846,N_11736,N_9410);
and U14847 (N_14847,N_10571,N_9786);
nor U14848 (N_14848,N_10702,N_10989);
nand U14849 (N_14849,N_11991,N_10581);
and U14850 (N_14850,N_9002,N_9099);
nor U14851 (N_14851,N_10677,N_11220);
xnor U14852 (N_14852,N_9106,N_11844);
or U14853 (N_14853,N_10112,N_11031);
xor U14854 (N_14854,N_9391,N_9271);
or U14855 (N_14855,N_10901,N_9954);
and U14856 (N_14856,N_11055,N_9758);
or U14857 (N_14857,N_9970,N_9572);
nor U14858 (N_14858,N_10563,N_11184);
and U14859 (N_14859,N_11590,N_9685);
or U14860 (N_14860,N_10204,N_9875);
xor U14861 (N_14861,N_11473,N_10745);
xnor U14862 (N_14862,N_10322,N_11445);
nor U14863 (N_14863,N_9792,N_11125);
nand U14864 (N_14864,N_11751,N_11018);
and U14865 (N_14865,N_9745,N_10309);
nand U14866 (N_14866,N_11283,N_9496);
or U14867 (N_14867,N_9919,N_9303);
and U14868 (N_14868,N_11716,N_11622);
nor U14869 (N_14869,N_11233,N_9394);
or U14870 (N_14870,N_9727,N_10215);
nor U14871 (N_14871,N_10686,N_9960);
nand U14872 (N_14872,N_9753,N_10157);
nor U14873 (N_14873,N_9854,N_11537);
and U14874 (N_14874,N_9330,N_10019);
nor U14875 (N_14875,N_11192,N_9727);
xnor U14876 (N_14876,N_11166,N_9220);
xnor U14877 (N_14877,N_9644,N_10174);
xor U14878 (N_14878,N_11771,N_9609);
and U14879 (N_14879,N_11490,N_11890);
nand U14880 (N_14880,N_11791,N_10474);
nand U14881 (N_14881,N_11371,N_11977);
nor U14882 (N_14882,N_11106,N_10972);
and U14883 (N_14883,N_11859,N_10837);
or U14884 (N_14884,N_9515,N_9242);
nor U14885 (N_14885,N_11436,N_9200);
and U14886 (N_14886,N_9679,N_9151);
nand U14887 (N_14887,N_10168,N_9209);
or U14888 (N_14888,N_10953,N_10043);
or U14889 (N_14889,N_11464,N_11622);
and U14890 (N_14890,N_9335,N_11596);
nor U14891 (N_14891,N_11457,N_11139);
xor U14892 (N_14892,N_10748,N_11594);
or U14893 (N_14893,N_9106,N_11031);
or U14894 (N_14894,N_10998,N_9477);
nand U14895 (N_14895,N_11278,N_11798);
and U14896 (N_14896,N_10799,N_10482);
or U14897 (N_14897,N_9870,N_10061);
nand U14898 (N_14898,N_11195,N_9874);
nor U14899 (N_14899,N_9357,N_10953);
and U14900 (N_14900,N_11052,N_10670);
nand U14901 (N_14901,N_11883,N_10048);
nor U14902 (N_14902,N_11436,N_11494);
nor U14903 (N_14903,N_11237,N_10988);
xnor U14904 (N_14904,N_9991,N_11750);
xnor U14905 (N_14905,N_9762,N_11485);
xor U14906 (N_14906,N_9144,N_9684);
nand U14907 (N_14907,N_10009,N_9376);
xnor U14908 (N_14908,N_9179,N_10379);
xnor U14909 (N_14909,N_9205,N_11090);
or U14910 (N_14910,N_9256,N_10578);
nor U14911 (N_14911,N_9288,N_11363);
and U14912 (N_14912,N_11080,N_11997);
and U14913 (N_14913,N_11083,N_9310);
and U14914 (N_14914,N_9665,N_10172);
xor U14915 (N_14915,N_9707,N_10686);
nor U14916 (N_14916,N_11196,N_9011);
xor U14917 (N_14917,N_11850,N_9008);
nand U14918 (N_14918,N_10371,N_9541);
or U14919 (N_14919,N_10949,N_10882);
nor U14920 (N_14920,N_10949,N_10774);
and U14921 (N_14921,N_11277,N_11772);
nand U14922 (N_14922,N_10192,N_9401);
nand U14923 (N_14923,N_9380,N_10802);
xor U14924 (N_14924,N_10402,N_11023);
and U14925 (N_14925,N_9471,N_11553);
or U14926 (N_14926,N_9379,N_11265);
and U14927 (N_14927,N_11174,N_10351);
and U14928 (N_14928,N_10846,N_10212);
and U14929 (N_14929,N_10197,N_11466);
or U14930 (N_14930,N_9214,N_9290);
nor U14931 (N_14931,N_11079,N_10255);
nand U14932 (N_14932,N_9571,N_11590);
nand U14933 (N_14933,N_11128,N_10243);
nand U14934 (N_14934,N_10017,N_9012);
nand U14935 (N_14935,N_10642,N_11365);
xnor U14936 (N_14936,N_10824,N_9826);
or U14937 (N_14937,N_10147,N_9988);
or U14938 (N_14938,N_9006,N_11180);
or U14939 (N_14939,N_11476,N_9732);
xor U14940 (N_14940,N_9267,N_9876);
xnor U14941 (N_14941,N_11710,N_10750);
nand U14942 (N_14942,N_9861,N_10111);
nand U14943 (N_14943,N_10507,N_10450);
or U14944 (N_14944,N_10764,N_11906);
nor U14945 (N_14945,N_9970,N_10176);
xnor U14946 (N_14946,N_11418,N_11660);
and U14947 (N_14947,N_10671,N_9360);
or U14948 (N_14948,N_10145,N_9782);
xnor U14949 (N_14949,N_10966,N_11152);
xor U14950 (N_14950,N_10620,N_10071);
and U14951 (N_14951,N_10878,N_9640);
xnor U14952 (N_14952,N_10077,N_10192);
nor U14953 (N_14953,N_11721,N_10665);
nand U14954 (N_14954,N_9460,N_11957);
xnor U14955 (N_14955,N_11452,N_11495);
and U14956 (N_14956,N_10285,N_10444);
or U14957 (N_14957,N_9447,N_10194);
xor U14958 (N_14958,N_11134,N_11612);
and U14959 (N_14959,N_9597,N_11283);
xnor U14960 (N_14960,N_9710,N_10250);
nor U14961 (N_14961,N_11098,N_10501);
nand U14962 (N_14962,N_11495,N_11490);
and U14963 (N_14963,N_9298,N_9142);
and U14964 (N_14964,N_11095,N_10816);
or U14965 (N_14965,N_10842,N_11475);
nor U14966 (N_14966,N_9063,N_11645);
xor U14967 (N_14967,N_11402,N_11365);
nand U14968 (N_14968,N_9891,N_9296);
or U14969 (N_14969,N_10704,N_9015);
nand U14970 (N_14970,N_10263,N_11264);
xor U14971 (N_14971,N_10981,N_11715);
xnor U14972 (N_14972,N_9332,N_9831);
nor U14973 (N_14973,N_9096,N_11682);
xnor U14974 (N_14974,N_9517,N_10001);
or U14975 (N_14975,N_10598,N_10218);
nor U14976 (N_14976,N_10374,N_10518);
or U14977 (N_14977,N_10281,N_10478);
or U14978 (N_14978,N_11864,N_11581);
nand U14979 (N_14979,N_11605,N_11181);
or U14980 (N_14980,N_10501,N_10341);
xnor U14981 (N_14981,N_11506,N_10627);
xnor U14982 (N_14982,N_9611,N_11844);
nand U14983 (N_14983,N_9690,N_9151);
nand U14984 (N_14984,N_9691,N_11859);
xnor U14985 (N_14985,N_9727,N_11415);
or U14986 (N_14986,N_10182,N_10085);
and U14987 (N_14987,N_9686,N_9384);
nand U14988 (N_14988,N_10686,N_10350);
or U14989 (N_14989,N_9513,N_11588);
or U14990 (N_14990,N_9945,N_11301);
xor U14991 (N_14991,N_9188,N_11126);
and U14992 (N_14992,N_10852,N_9154);
xor U14993 (N_14993,N_10255,N_10648);
nand U14994 (N_14994,N_11438,N_11823);
xor U14995 (N_14995,N_11523,N_10105);
nor U14996 (N_14996,N_11353,N_11601);
xnor U14997 (N_14997,N_10221,N_10076);
nor U14998 (N_14998,N_11230,N_11825);
nand U14999 (N_14999,N_10299,N_10684);
and U15000 (N_15000,N_12952,N_12098);
or U15001 (N_15001,N_12322,N_12499);
or U15002 (N_15002,N_14402,N_14475);
or U15003 (N_15003,N_13546,N_13620);
nand U15004 (N_15004,N_13053,N_13954);
xnor U15005 (N_15005,N_13371,N_12054);
nand U15006 (N_15006,N_13678,N_13912);
and U15007 (N_15007,N_13801,N_13779);
nor U15008 (N_15008,N_13504,N_12187);
and U15009 (N_15009,N_14988,N_12540);
or U15010 (N_15010,N_14750,N_13323);
nand U15011 (N_15011,N_12260,N_13332);
xor U15012 (N_15012,N_12692,N_13548);
nand U15013 (N_15013,N_14708,N_14295);
and U15014 (N_15014,N_14860,N_14246);
nor U15015 (N_15015,N_12029,N_14211);
xnor U15016 (N_15016,N_13243,N_14282);
or U15017 (N_15017,N_12996,N_12657);
and U15018 (N_15018,N_13988,N_14081);
nand U15019 (N_15019,N_12658,N_14610);
or U15020 (N_15020,N_13310,N_13203);
nand U15021 (N_15021,N_14560,N_13676);
or U15022 (N_15022,N_13439,N_12326);
nand U15023 (N_15023,N_14118,N_14710);
nand U15024 (N_15024,N_13986,N_14338);
and U15025 (N_15025,N_12794,N_12860);
nand U15026 (N_15026,N_13422,N_12174);
nand U15027 (N_15027,N_12044,N_14464);
xnor U15028 (N_15028,N_12778,N_12505);
xor U15029 (N_15029,N_14827,N_14365);
and U15030 (N_15030,N_13214,N_12739);
or U15031 (N_15031,N_14615,N_12071);
and U15032 (N_15032,N_13916,N_12127);
nor U15033 (N_15033,N_12500,N_14993);
and U15034 (N_15034,N_14408,N_12144);
and U15035 (N_15035,N_12106,N_14740);
nand U15036 (N_15036,N_12353,N_14648);
nor U15037 (N_15037,N_14370,N_14284);
nand U15038 (N_15038,N_14700,N_13931);
xnor U15039 (N_15039,N_14389,N_12443);
nand U15040 (N_15040,N_14042,N_12792);
and U15041 (N_15041,N_12669,N_12817);
and U15042 (N_15042,N_14459,N_12003);
or U15043 (N_15043,N_12628,N_13218);
nand U15044 (N_15044,N_12440,N_14661);
nand U15045 (N_15045,N_14624,N_13345);
or U15046 (N_15046,N_12367,N_14020);
nor U15047 (N_15047,N_14482,N_12747);
or U15048 (N_15048,N_12150,N_13343);
or U15049 (N_15049,N_13478,N_12972);
xnor U15050 (N_15050,N_13339,N_13118);
or U15051 (N_15051,N_12185,N_14314);
nand U15052 (N_15052,N_13408,N_14257);
and U15053 (N_15053,N_13461,N_12093);
xor U15054 (N_15054,N_13087,N_13711);
nor U15055 (N_15055,N_14622,N_12049);
and U15056 (N_15056,N_13274,N_12570);
or U15057 (N_15057,N_14714,N_12284);
or U15058 (N_15058,N_12194,N_12644);
or U15059 (N_15059,N_12230,N_14405);
nand U15060 (N_15060,N_14972,N_12744);
nand U15061 (N_15061,N_14015,N_14256);
nor U15062 (N_15062,N_13945,N_12234);
xor U15063 (N_15063,N_12653,N_14852);
xor U15064 (N_15064,N_12730,N_13248);
or U15065 (N_15065,N_14625,N_12471);
nor U15066 (N_15066,N_12387,N_14356);
and U15067 (N_15067,N_14251,N_12766);
nand U15068 (N_15068,N_13261,N_12982);
and U15069 (N_15069,N_14878,N_14091);
and U15070 (N_15070,N_13024,N_12183);
and U15071 (N_15071,N_14795,N_14749);
xnor U15072 (N_15072,N_12955,N_13498);
nand U15073 (N_15073,N_13455,N_14919);
and U15074 (N_15074,N_13458,N_13199);
xor U15075 (N_15075,N_14302,N_13970);
nand U15076 (N_15076,N_12749,N_13532);
nor U15077 (N_15077,N_14078,N_13657);
xor U15078 (N_15078,N_13895,N_13840);
nor U15079 (N_15079,N_12215,N_13095);
nor U15080 (N_15080,N_13627,N_13204);
and U15081 (N_15081,N_12232,N_13100);
or U15082 (N_15082,N_14016,N_13948);
or U15083 (N_15083,N_14718,N_14004);
and U15084 (N_15084,N_14554,N_14634);
nor U15085 (N_15085,N_12572,N_12961);
and U15086 (N_15086,N_12461,N_14910);
or U15087 (N_15087,N_13534,N_13445);
xnor U15088 (N_15088,N_12268,N_12016);
or U15089 (N_15089,N_14541,N_14641);
or U15090 (N_15090,N_14316,N_14924);
nor U15091 (N_15091,N_12090,N_13847);
or U15092 (N_15092,N_12812,N_12409);
nand U15093 (N_15093,N_12965,N_14744);
nand U15094 (N_15094,N_14715,N_13667);
xor U15095 (N_15095,N_14550,N_14031);
nor U15096 (N_15096,N_12124,N_14328);
xor U15097 (N_15097,N_12686,N_14094);
xor U15098 (N_15098,N_13704,N_13978);
and U15099 (N_15099,N_14990,N_13056);
nand U15100 (N_15100,N_12064,N_12013);
nor U15101 (N_15101,N_12201,N_14638);
or U15102 (N_15102,N_13707,N_14717);
and U15103 (N_15103,N_12608,N_14962);
xor U15104 (N_15104,N_12487,N_13036);
xor U15105 (N_15105,N_14593,N_12231);
xor U15106 (N_15106,N_13415,N_14659);
and U15107 (N_15107,N_12698,N_13104);
or U15108 (N_15108,N_14259,N_13968);
and U15109 (N_15109,N_12298,N_14944);
nor U15110 (N_15110,N_13474,N_13722);
nor U15111 (N_15111,N_12432,N_12709);
and U15112 (N_15112,N_14604,N_14064);
or U15113 (N_15113,N_14479,N_13173);
nand U15114 (N_15114,N_12903,N_14010);
nand U15115 (N_15115,N_14301,N_12844);
nand U15116 (N_15116,N_14269,N_14870);
xor U15117 (N_15117,N_14649,N_14508);
nor U15118 (N_15118,N_12642,N_12280);
nand U15119 (N_15119,N_14174,N_13318);
and U15120 (N_15120,N_12079,N_14556);
xnor U15121 (N_15121,N_13702,N_13975);
and U15122 (N_15122,N_14192,N_14838);
nor U15123 (N_15123,N_14821,N_13511);
or U15124 (N_15124,N_12330,N_12114);
or U15125 (N_15125,N_12905,N_12211);
nand U15126 (N_15126,N_13977,N_14672);
or U15127 (N_15127,N_14453,N_14461);
nand U15128 (N_15128,N_14522,N_13322);
nand U15129 (N_15129,N_13698,N_14986);
and U15130 (N_15130,N_13877,N_12950);
or U15131 (N_15131,N_14431,N_14952);
nor U15132 (N_15132,N_13156,N_14486);
or U15133 (N_15133,N_12179,N_12087);
xor U15134 (N_15134,N_12702,N_14893);
or U15135 (N_15135,N_14800,N_12610);
xor U15136 (N_15136,N_12202,N_13932);
xnor U15137 (N_15137,N_14588,N_13241);
nor U15138 (N_15138,N_13959,N_13418);
nand U15139 (N_15139,N_13183,N_14616);
nor U15140 (N_15140,N_13216,N_12863);
or U15141 (N_15141,N_13842,N_14601);
nor U15142 (N_15142,N_14177,N_12308);
nand U15143 (N_15143,N_13290,N_13784);
nand U15144 (N_15144,N_12160,N_12327);
nand U15145 (N_15145,N_13868,N_12890);
xor U15146 (N_15146,N_13939,N_14983);
and U15147 (N_15147,N_14375,N_14580);
xnor U15148 (N_15148,N_12162,N_13633);
nand U15149 (N_15149,N_12963,N_12303);
xor U15150 (N_15150,N_12395,N_12385);
xor U15151 (N_15151,N_12929,N_13835);
xnor U15152 (N_15152,N_13068,N_13741);
xnor U15153 (N_15153,N_14707,N_13120);
xnor U15154 (N_15154,N_13206,N_12904);
xnor U15155 (N_15155,N_12891,N_14403);
nor U15156 (N_15156,N_13761,N_13757);
and U15157 (N_15157,N_14936,N_12586);
xor U15158 (N_15158,N_14546,N_13855);
xnor U15159 (N_15159,N_12780,N_14327);
nor U15160 (N_15160,N_12544,N_14846);
or U15161 (N_15161,N_14837,N_14653);
nor U15162 (N_15162,N_14500,N_13090);
nand U15163 (N_15163,N_14782,N_14529);
nand U15164 (N_15164,N_13544,N_14680);
nor U15165 (N_15165,N_14501,N_13116);
nand U15166 (N_15166,N_13346,N_12804);
and U15167 (N_15167,N_12997,N_12184);
xor U15168 (N_15168,N_13860,N_12810);
xor U15169 (N_15169,N_12301,N_13136);
nor U15170 (N_15170,N_14263,N_14805);
xnor U15171 (N_15171,N_12641,N_12449);
or U15172 (N_15172,N_14854,N_14527);
nand U15173 (N_15173,N_14466,N_13794);
nor U15174 (N_15174,N_13328,N_13121);
and U15175 (N_15175,N_12828,N_12726);
xor U15176 (N_15176,N_14340,N_14332);
or U15177 (N_15177,N_13688,N_13046);
or U15178 (N_15178,N_12683,N_14571);
xnor U15179 (N_15179,N_13453,N_13683);
and U15180 (N_15180,N_14640,N_12480);
nor U15181 (N_15181,N_14791,N_12085);
and U15182 (N_15182,N_12816,N_13781);
xnor U15183 (N_15183,N_14117,N_14558);
nor U15184 (N_15184,N_13250,N_14669);
nand U15185 (N_15185,N_14404,N_13078);
xnor U15186 (N_15186,N_13712,N_12271);
nor U15187 (N_15187,N_13993,N_12428);
nand U15188 (N_15188,N_13837,N_12012);
nor U15189 (N_15189,N_13485,N_12228);
and U15190 (N_15190,N_13174,N_13251);
nor U15191 (N_15191,N_14047,N_14339);
xor U15192 (N_15192,N_14977,N_14084);
xor U15193 (N_15193,N_12836,N_14916);
xnor U15194 (N_15194,N_13446,N_13198);
nor U15195 (N_15195,N_14543,N_14364);
xnor U15196 (N_15196,N_12645,N_12634);
and U15197 (N_15197,N_12519,N_13872);
or U15198 (N_15198,N_14563,N_12140);
and U15199 (N_15199,N_12244,N_14219);
or U15200 (N_15200,N_12027,N_12694);
xor U15201 (N_15201,N_13226,N_13043);
and U15202 (N_15202,N_12763,N_12306);
and U15203 (N_15203,N_14242,N_14573);
nand U15204 (N_15204,N_12199,N_13867);
and U15205 (N_15205,N_14080,N_12893);
nand U15206 (N_15206,N_12210,N_13486);
or U15207 (N_15207,N_12055,N_12565);
nor U15208 (N_15208,N_12946,N_13002);
xnor U15209 (N_15209,N_12801,N_12486);
xor U15210 (N_15210,N_13184,N_14658);
or U15211 (N_15211,N_12751,N_13933);
nand U15212 (N_15212,N_14807,N_14545);
nor U15213 (N_15213,N_13831,N_14609);
and U15214 (N_15214,N_12907,N_14238);
nor U15215 (N_15215,N_13822,N_12411);
nor U15216 (N_15216,N_13969,N_13473);
xnor U15217 (N_15217,N_13049,N_12916);
nor U15218 (N_15218,N_13890,N_14165);
xor U15219 (N_15219,N_14154,N_12623);
xor U15220 (N_15220,N_12571,N_13144);
nor U15221 (N_15221,N_12897,N_13137);
nor U15222 (N_15222,N_12881,N_13426);
nor U15223 (N_15223,N_14412,N_14937);
nor U15224 (N_15224,N_14141,N_13736);
nor U15225 (N_15225,N_13268,N_13244);
or U15226 (N_15226,N_14022,N_13480);
xnor U15227 (N_15227,N_13744,N_13012);
nor U15228 (N_15228,N_12932,N_13409);
nor U15229 (N_15229,N_12545,N_14864);
and U15230 (N_15230,N_13723,N_13319);
nand U15231 (N_15231,N_13530,N_12771);
nor U15232 (N_15232,N_13283,N_12913);
nor U15233 (N_15233,N_13605,N_13745);
xnor U15234 (N_15234,N_13186,N_12323);
or U15235 (N_15235,N_13812,N_12377);
nand U15236 (N_15236,N_14841,N_12360);
or U15237 (N_15237,N_14665,N_12464);
and U15238 (N_15238,N_13971,N_13070);
xnor U15239 (N_15239,N_12663,N_14419);
and U15240 (N_15240,N_14430,N_13560);
or U15241 (N_15241,N_12439,N_13776);
xor U15242 (N_15242,N_12148,N_14025);
nand U15243 (N_15243,N_14865,N_14243);
or U15244 (N_15244,N_13720,N_14934);
nand U15245 (N_15245,N_13232,N_13569);
and U15246 (N_15246,N_14848,N_12137);
nor U15247 (N_15247,N_14746,N_14682);
or U15248 (N_15248,N_14823,N_14853);
nand U15249 (N_15249,N_14828,N_14191);
nor U15250 (N_15250,N_12261,N_14462);
and U15251 (N_15251,N_13314,N_13879);
and U15252 (N_15252,N_13354,N_12309);
xnor U15253 (N_15253,N_14420,N_12257);
xor U15254 (N_15254,N_12580,N_12563);
xor U15255 (N_15255,N_12962,N_12100);
nand U15256 (N_15256,N_14945,N_13773);
nand U15257 (N_15257,N_12638,N_12442);
or U15258 (N_15258,N_13699,N_12237);
nor U15259 (N_15259,N_13385,N_14953);
xnor U15260 (N_15260,N_13935,N_13391);
nor U15261 (N_15261,N_12640,N_13936);
and U15262 (N_15262,N_12037,N_14903);
xnor U15263 (N_15263,N_12517,N_14308);
or U15264 (N_15264,N_14310,N_14531);
xor U15265 (N_15265,N_14399,N_13737);
nand U15266 (N_15266,N_12599,N_12002);
and U15267 (N_15267,N_13522,N_12119);
and U15268 (N_15268,N_12823,N_13335);
nand U15269 (N_15269,N_13273,N_13513);
xor U15270 (N_15270,N_14030,N_12458);
nand U15271 (N_15271,N_13146,N_13111);
or U15272 (N_15272,N_14196,N_14305);
xnor U15273 (N_15273,N_14895,N_13031);
and U15274 (N_15274,N_14083,N_14930);
or U15275 (N_15275,N_12617,N_13938);
xnor U15276 (N_15276,N_13684,N_13059);
and U15277 (N_15277,N_13357,N_14753);
or U15278 (N_15278,N_14197,N_14176);
nand U15279 (N_15279,N_12951,N_14330);
xnor U15280 (N_15280,N_12413,N_13981);
nand U15281 (N_15281,N_12204,N_14199);
nor U15282 (N_15282,N_14422,N_13885);
nand U15283 (N_15283,N_12745,N_13753);
nand U15284 (N_15284,N_14454,N_14738);
or U15285 (N_15285,N_13459,N_13941);
and U15286 (N_15286,N_14947,N_12177);
nand U15287 (N_15287,N_13420,N_13778);
nor U15288 (N_15288,N_14789,N_13145);
or U15289 (N_15289,N_14465,N_12621);
nor U15290 (N_15290,N_13075,N_14568);
nor U15291 (N_15291,N_13554,N_12958);
xor U15292 (N_15292,N_12329,N_12573);
and U15293 (N_15293,N_13901,N_12287);
xor U15294 (N_15294,N_14955,N_14683);
xnor U15295 (N_15295,N_14427,N_12082);
xor U15296 (N_15296,N_14697,N_12320);
xor U15297 (N_15297,N_14814,N_13280);
xnor U15298 (N_15298,N_14125,N_13399);
or U15299 (N_15299,N_13413,N_14892);
and U15300 (N_15300,N_12220,N_14442);
nor U15301 (N_15301,N_14398,N_14104);
and U15302 (N_15302,N_12954,N_12911);
xor U15303 (N_15303,N_14434,N_14353);
nand U15304 (N_15304,N_13202,N_12130);
or U15305 (N_15305,N_12340,N_12117);
xor U15306 (N_15306,N_13797,N_14306);
or U15307 (N_15307,N_13360,N_12758);
and U15308 (N_15308,N_14222,N_13172);
nand U15309 (N_15309,N_14687,N_12345);
xor U15310 (N_15310,N_13390,N_12947);
nand U15311 (N_15311,N_13854,N_14109);
nor U15312 (N_15312,N_14896,N_12191);
or U15313 (N_15313,N_14051,N_14562);
nor U15314 (N_15314,N_13542,N_14518);
and U15315 (N_15315,N_13682,N_13246);
and U15316 (N_15316,N_14173,N_13494);
xor U15317 (N_15317,N_13576,N_12707);
nor U15318 (N_15318,N_13456,N_14374);
nand U15319 (N_15319,N_14958,N_12875);
nor U15320 (N_15320,N_12371,N_12511);
xnor U15321 (N_15321,N_13552,N_12459);
and U15322 (N_15322,N_13851,N_12516);
or U15323 (N_15323,N_12008,N_14880);
xor U15324 (N_15324,N_13225,N_13787);
nor U15325 (N_15325,N_12856,N_14203);
and U15326 (N_15326,N_14480,N_12376);
xor U15327 (N_15327,N_14086,N_14797);
xnor U15328 (N_15328,N_14956,N_13023);
or U15329 (N_15329,N_13481,N_13001);
xor U15330 (N_15330,N_12125,N_12721);
nor U15331 (N_15331,N_13067,N_14394);
and U15332 (N_15332,N_13675,N_14280);
xnor U15333 (N_15333,N_14406,N_14523);
nand U15334 (N_15334,N_12530,N_14171);
and U15335 (N_15335,N_14255,N_14671);
and U15336 (N_15336,N_13313,N_13019);
nand U15337 (N_15337,N_12398,N_14711);
and U15338 (N_15338,N_12533,N_14676);
and U15339 (N_15339,N_14409,N_13272);
xor U15340 (N_15340,N_12613,N_13696);
xor U15341 (N_15341,N_14297,N_12543);
or U15342 (N_15342,N_12834,N_14499);
xor U15343 (N_15343,N_13593,N_12337);
or U15344 (N_15344,N_12981,N_13134);
xor U15345 (N_15345,N_14233,N_13253);
and U15346 (N_15346,N_14592,N_13630);
and U15347 (N_15347,N_12346,N_14492);
nand U15348 (N_15348,N_12838,N_12249);
nand U15349 (N_15349,N_14587,N_14647);
xnor U15350 (N_15350,N_13082,N_12622);
xnor U15351 (N_15351,N_14134,N_14963);
nor U15352 (N_15352,N_12990,N_14831);
nand U15353 (N_15353,N_13414,N_13887);
nand U15354 (N_15354,N_14858,N_13499);
nor U15355 (N_15355,N_14686,N_12343);
nand U15356 (N_15356,N_13342,N_13311);
and U15357 (N_15357,N_12788,N_14567);
nand U15358 (N_15358,N_12472,N_13009);
nand U15359 (N_15359,N_14009,N_13516);
and U15360 (N_15360,N_14722,N_12556);
nor U15361 (N_15361,N_14245,N_12976);
xnor U15362 (N_15362,N_13384,N_13131);
and U15363 (N_15363,N_14494,N_12677);
xnor U15364 (N_15364,N_12600,N_12294);
or U15365 (N_15365,N_14098,N_12205);
or U15366 (N_15366,N_14391,N_13193);
nor U15367 (N_15367,N_12446,N_12909);
nor U15368 (N_15368,N_12575,N_14759);
or U15369 (N_15369,N_13433,N_12108);
or U15370 (N_15370,N_14451,N_13727);
or U15371 (N_15371,N_14777,N_14396);
nand U15372 (N_15372,N_13331,N_12876);
or U15373 (N_15373,N_13115,N_13828);
nor U15374 (N_15374,N_13578,N_14635);
or U15375 (N_15375,N_14628,N_14706);
or U15376 (N_15376,N_12720,N_12372);
nand U15377 (N_15377,N_13651,N_14526);
or U15378 (N_15378,N_14923,N_13222);
nor U15379 (N_15379,N_14555,N_13519);
xnor U15380 (N_15380,N_14547,N_14013);
nor U15381 (N_15381,N_12549,N_14663);
nor U15382 (N_15382,N_14024,N_13929);
nor U15383 (N_15383,N_13387,N_14574);
nor U15384 (N_15384,N_14390,N_13086);
xnor U15385 (N_15385,N_14785,N_14268);
nand U15386 (N_15386,N_12014,N_12534);
and U15387 (N_15387,N_14850,N_14914);
xnor U15388 (N_15388,N_12546,N_14135);
xor U15389 (N_15389,N_13038,N_12381);
xor U15390 (N_15390,N_13472,N_13905);
nor U15391 (N_15391,N_13673,N_12020);
xor U15392 (N_15392,N_14757,N_14915);
nand U15393 (N_15393,N_13896,N_13892);
or U15394 (N_15394,N_12773,N_14446);
xnor U15395 (N_15395,N_12388,N_14780);
or U15396 (N_15396,N_14804,N_13247);
nand U15397 (N_15397,N_12070,N_12935);
and U15398 (N_15398,N_14040,N_14241);
and U15399 (N_15399,N_14215,N_14826);
nand U15400 (N_15400,N_12251,N_14110);
nand U15401 (N_15401,N_12092,N_13462);
nand U15402 (N_15402,N_13122,N_13807);
nand U15403 (N_15403,N_14190,N_12949);
nor U15404 (N_15404,N_13734,N_12923);
xor U15405 (N_15405,N_12208,N_14283);
nor U15406 (N_15406,N_12004,N_14581);
and U15407 (N_15407,N_13263,N_13441);
nor U15408 (N_15408,N_13351,N_12808);
nand U15409 (N_15409,N_14476,N_14964);
and U15410 (N_15410,N_13983,N_14946);
nand U15411 (N_15411,N_12978,N_13690);
nand U15412 (N_15412,N_13798,N_14762);
xnor U15413 (N_15413,N_13958,N_12995);
nand U15414 (N_15414,N_13048,N_13898);
nand U15415 (N_15415,N_14488,N_14829);
nand U15416 (N_15416,N_12803,N_12310);
nand U15417 (N_15417,N_13438,N_13518);
nor U15418 (N_15418,N_12226,N_12918);
nor U15419 (N_15419,N_12258,N_13490);
nor U15420 (N_15420,N_13742,N_14133);
xnor U15421 (N_15421,N_14705,N_14536);
and U15422 (N_15422,N_12588,N_13479);
xnor U15423 (N_15423,N_12051,N_13703);
or U15424 (N_15424,N_13168,N_13662);
xnor U15425 (N_15425,N_12655,N_12296);
xnor U15426 (N_15426,N_14460,N_14415);
nand U15427 (N_15427,N_13527,N_14935);
xnor U15428 (N_15428,N_13163,N_13874);
xnor U15429 (N_15429,N_13304,N_12068);
and U15430 (N_15430,N_12384,N_13265);
nand U15431 (N_15431,N_13242,N_12852);
xnor U15432 (N_15432,N_12943,N_13735);
xor U15433 (N_15433,N_12986,N_12900);
and U15434 (N_15434,N_14272,N_12919);
or U15435 (N_15435,N_13899,N_12775);
or U15436 (N_15436,N_13824,N_14161);
or U15437 (N_15437,N_14772,N_12688);
nor U15438 (N_15438,N_14265,N_14904);
and U15439 (N_15439,N_12266,N_13792);
or U15440 (N_15440,N_12889,N_13317);
or U15441 (N_15441,N_14801,N_12646);
nand U15442 (N_15442,N_12886,N_13689);
xor U15443 (N_15443,N_12102,N_14202);
nand U15444 (N_15444,N_12138,N_12356);
and U15445 (N_15445,N_14204,N_13804);
nand U15446 (N_15446,N_13150,N_12774);
nand U15447 (N_15447,N_14445,N_13417);
xor U15448 (N_15448,N_12855,N_12722);
nand U15449 (N_15449,N_14668,N_14386);
nor U15450 (N_15450,N_13694,N_12733);
nand U15451 (N_15451,N_14662,N_12568);
or U15452 (N_15452,N_13449,N_12469);
xnor U15453 (N_15453,N_12895,N_14372);
or U15454 (N_15454,N_14382,N_12042);
xnor U15455 (N_15455,N_14017,N_14231);
and U15456 (N_15456,N_14320,N_14029);
nand U15457 (N_15457,N_14002,N_12936);
or U15458 (N_15458,N_12648,N_12328);
nor U15459 (N_15459,N_13326,N_14275);
or U15460 (N_15460,N_13695,N_12521);
or U15461 (N_15461,N_12419,N_14418);
nand U15462 (N_15462,N_12216,N_12765);
xor U15463 (N_15463,N_12259,N_13514);
nor U15464 (N_15464,N_14443,N_14225);
xor U15465 (N_15465,N_13607,N_14240);
and U15466 (N_15466,N_12010,N_12252);
or U15467 (N_15467,N_14730,N_13239);
nand U15468 (N_15468,N_12939,N_12970);
nor U15469 (N_15469,N_14867,N_14585);
and U15470 (N_15470,N_12157,N_13308);
nand U15471 (N_15471,N_12462,N_12429);
and U15472 (N_15472,N_14088,N_14105);
and U15473 (N_15473,N_13367,N_13495);
or U15474 (N_15474,N_12041,N_12242);
nor U15475 (N_15475,N_12547,N_12984);
and U15476 (N_15476,N_14261,N_12716);
xnor U15477 (N_15477,N_12438,N_14608);
nand U15478 (N_15478,N_14812,N_13748);
or U15479 (N_15479,N_14216,N_12760);
nand U15480 (N_15480,N_12047,N_12293);
xor U15481 (N_15481,N_14477,N_14037);
nand U15482 (N_15482,N_13614,N_13999);
nor U15483 (N_15483,N_12318,N_13786);
and U15484 (N_15484,N_13965,N_13592);
and U15485 (N_15485,N_14633,N_13826);
nand U15486 (N_15486,N_12782,N_13819);
or U15487 (N_15487,N_13006,N_12437);
nor U15488 (N_15488,N_14470,N_12914);
and U15489 (N_15489,N_13224,N_14169);
or U15490 (N_15490,N_12930,N_13170);
nand U15491 (N_15491,N_12455,N_13307);
nor U15492 (N_15492,N_12602,N_13624);
nor U15493 (N_15493,N_14198,N_13341);
or U15494 (N_15494,N_13058,N_12668);
nand U15495 (N_15495,N_13035,N_12304);
nor U15496 (N_15496,N_12196,N_12111);
nor U15497 (N_15497,N_12626,N_13231);
xor U15498 (N_15498,N_12906,N_14429);
and U15499 (N_15499,N_12841,N_12589);
or U15500 (N_15500,N_14168,N_12956);
xnor U15501 (N_15501,N_14143,N_13228);
xor U15502 (N_15502,N_13037,N_12312);
and U15503 (N_15503,N_12849,N_12316);
and U15504 (N_15504,N_12240,N_14267);
nand U15505 (N_15505,N_13435,N_12406);
xnor U15506 (N_15506,N_13029,N_13586);
and U15507 (N_15507,N_12938,N_13266);
xor U15508 (N_15508,N_14961,N_13770);
nor U15509 (N_15509,N_12998,N_14891);
xor U15510 (N_15510,N_14342,N_14426);
nor U15511 (N_15511,N_12235,N_13364);
or U15512 (N_15512,N_12375,N_13362);
nor U15513 (N_15513,N_13677,N_13052);
xnor U15514 (N_15514,N_13296,N_13603);
nand U15515 (N_15515,N_14220,N_13072);
nand U15516 (N_15516,N_12831,N_13140);
nor U15517 (N_15517,N_14764,N_12811);
xnor U15518 (N_15518,N_13401,N_14783);
nor U15519 (N_15519,N_12877,N_12291);
nand U15520 (N_15520,N_14995,N_13309);
and U15521 (N_15521,N_13922,N_13760);
nand U15522 (N_15522,N_14596,N_12402);
xor U15523 (N_15523,N_14579,N_14639);
xnor U15524 (N_15524,N_14735,N_14097);
or U15525 (N_15525,N_14741,N_14296);
nand U15526 (N_15526,N_12022,N_14603);
nor U15527 (N_15527,N_14159,N_12456);
or U15528 (N_15528,N_13114,N_14620);
and U15529 (N_15529,N_12922,N_14586);
or U15530 (N_15530,N_13830,N_12422);
nor U15531 (N_15531,N_14069,N_14871);
nor U15532 (N_15532,N_14260,N_13721);
and U15533 (N_15533,N_14611,N_14184);
xor U15534 (N_15534,N_14107,N_13252);
and U15535 (N_15535,N_14441,N_13021);
and U15536 (N_15536,N_12397,N_14922);
nor U15537 (N_15537,N_13227,N_13063);
and U15538 (N_15538,N_14006,N_13966);
nor U15539 (N_15539,N_14577,N_13668);
nand U15540 (N_15540,N_13568,N_13995);
and U15541 (N_15541,N_13541,N_14485);
nand U15542 (N_15542,N_14132,N_13482);
nand U15543 (N_15543,N_13352,N_14055);
and U15544 (N_15544,N_12289,N_14100);
xnor U15545 (N_15545,N_12974,N_13584);
and U15546 (N_15546,N_14535,N_12696);
xor U15547 (N_15547,N_12942,N_13129);
or U15548 (N_15548,N_13230,N_14163);
nor U15549 (N_15549,N_13884,N_13566);
or U15550 (N_15550,N_13392,N_13338);
xnor U15551 (N_15551,N_14721,N_12968);
nor U15552 (N_15552,N_13489,N_12941);
and U15553 (N_15553,N_12987,N_13815);
nor U15554 (N_15554,N_14702,N_12498);
nand U15555 (N_15555,N_12146,N_12279);
nor U15556 (N_15556,N_14279,N_12557);
nand U15557 (N_15557,N_14319,N_13964);
nor U15558 (N_15558,N_12169,N_13327);
and U15559 (N_15559,N_13025,N_12203);
or U15560 (N_15560,N_13460,N_12779);
nor U15561 (N_15561,N_12508,N_14630);
xnor U15562 (N_15562,N_12096,N_13934);
nand U15563 (N_15563,N_14361,N_12912);
xor U15564 (N_15564,N_14347,N_13641);
nor U15565 (N_15565,N_14435,N_14497);
or U15566 (N_15566,N_13219,N_14765);
or U15567 (N_15567,N_12858,N_13191);
nor U15568 (N_15568,N_12925,N_13436);
xor U15569 (N_15569,N_13407,N_14734);
or U15570 (N_15570,N_12843,N_12647);
and U15571 (N_15571,N_12112,N_14836);
nor U15572 (N_15572,N_13084,N_13207);
nor U15573 (N_15573,N_13747,N_14540);
nand U15574 (N_15574,N_12714,N_13171);
nor U15575 (N_15575,N_12276,N_12631);
nand U15576 (N_15576,N_14794,N_12396);
or U15577 (N_15577,N_13985,N_12966);
or U15578 (N_15578,N_14071,N_14607);
nor U15579 (N_15579,N_14076,N_14939);
xnor U15580 (N_15580,N_14369,N_12980);
xor U15581 (N_15581,N_13834,N_14063);
nand U15582 (N_15582,N_14072,N_13032);
nand U15583 (N_15583,N_14000,N_13994);
or U15584 (N_15584,N_13710,N_12139);
and U15585 (N_15585,N_12785,N_12218);
nand U15586 (N_15586,N_12207,N_12673);
or U15587 (N_15587,N_14695,N_13424);
and U15588 (N_15588,N_12350,N_13663);
and U15589 (N_15589,N_12386,N_14569);
or U15590 (N_15590,N_12975,N_12846);
xnor U15591 (N_15591,N_13238,N_13153);
nor U15592 (N_15592,N_13788,N_14436);
nor U15593 (N_15593,N_13169,N_14787);
xnor U15594 (N_15594,N_14819,N_13074);
nor U15595 (N_15595,N_13963,N_13976);
and U15596 (N_15596,N_12269,N_14602);
or U15597 (N_15597,N_14974,N_12408);
nand U15598 (N_15598,N_13921,N_13405);
or U15599 (N_15599,N_12822,N_12537);
or U15600 (N_15600,N_13740,N_12959);
nor U15601 (N_15601,N_12152,N_12040);
and U15602 (N_15602,N_13028,N_12536);
and U15603 (N_15603,N_12993,N_13871);
and U15604 (N_15604,N_12659,N_12161);
nand U15605 (N_15605,N_12799,N_13372);
nand U15606 (N_15606,N_13857,N_14583);
nand U15607 (N_15607,N_12078,N_13164);
nand U15608 (N_15608,N_14929,N_12359);
nor U15609 (N_15609,N_14318,N_13979);
nor U15610 (N_15610,N_14123,N_14572);
nor U15611 (N_15611,N_12364,N_14590);
nand U15612 (N_15612,N_14806,N_12574);
or U15613 (N_15613,N_13337,N_12879);
nor U15614 (N_15614,N_14907,N_12416);
nor U15615 (N_15615,N_12627,N_14578);
nor U15616 (N_15616,N_14551,N_13285);
or U15617 (N_15617,N_14747,N_13325);
nor U15618 (N_15618,N_14967,N_12066);
xnor U15619 (N_15619,N_14793,N_13717);
and U15620 (N_15620,N_12800,N_14731);
nand U15621 (N_15621,N_13756,N_13508);
xnor U15622 (N_15622,N_14285,N_12427);
or U15623 (N_15623,N_14186,N_12878);
and U15624 (N_15624,N_14713,N_12431);
xnor U15625 (N_15625,N_14991,N_14213);
and U15626 (N_15626,N_12527,N_14938);
xor U15627 (N_15627,N_14357,N_12392);
or U15628 (N_15628,N_14228,N_13465);
nand U15629 (N_15629,N_12145,N_12213);
or U15630 (N_15630,N_12212,N_12186);
nor U15631 (N_15631,N_12341,N_13563);
nand U15632 (N_15632,N_13130,N_14872);
nand U15633 (N_15633,N_13089,N_12835);
and U15634 (N_15634,N_14252,N_12718);
xor U15635 (N_15635,N_14193,N_13923);
nor U15636 (N_15636,N_14250,N_14290);
nand U15637 (N_15637,N_13113,N_14440);
xor U15638 (N_15638,N_13497,N_14102);
or U15639 (N_15639,N_13555,N_14542);
or U15640 (N_15640,N_13701,N_12300);
nor U15641 (N_15641,N_14994,N_13123);
xor U15642 (N_15642,N_12767,N_13262);
nand U15643 (N_15643,N_13623,N_14221);
and U15644 (N_15644,N_14035,N_12382);
or U15645 (N_15645,N_13982,N_12285);
and U15646 (N_15646,N_12420,N_12043);
nand U15647 (N_15647,N_13763,N_13974);
nand U15648 (N_15648,N_14281,N_12052);
nand U15649 (N_15649,N_12753,N_13303);
xor U15650 (N_15650,N_14985,N_14230);
nand U15651 (N_15651,N_13264,N_13869);
xnor U15652 (N_15652,N_13155,N_13503);
nand U15653 (N_15653,N_12748,N_13950);
and U15654 (N_15654,N_12369,N_13862);
and U15655 (N_15655,N_14666,N_14148);
nand U15656 (N_15656,N_14218,N_12492);
nand U15657 (N_15657,N_13475,N_13245);
nand U15658 (N_15658,N_14509,N_14329);
nor U15659 (N_15659,N_14768,N_12222);
or U15660 (N_15660,N_13109,N_13258);
and U15661 (N_15661,N_14681,N_13660);
nor U15662 (N_15662,N_13715,N_12089);
nand U15663 (N_15663,N_12781,N_14075);
nand U15664 (N_15664,N_14352,N_12901);
nor U15665 (N_15665,N_13398,N_12031);
nor U15666 (N_15666,N_13017,N_13454);
or U15667 (N_15667,N_12311,N_12848);
nor U15668 (N_15668,N_14380,N_13930);
and U15669 (N_15669,N_12192,N_12643);
and U15670 (N_15670,N_13187,N_12277);
nand U15671 (N_15671,N_13108,N_14684);
xnor U15672 (N_15672,N_14001,N_14559);
nand U15673 (N_15673,N_13538,N_13671);
and U15674 (N_15674,N_14452,N_12675);
or U15675 (N_15675,N_14312,N_13507);
or U15676 (N_15676,N_13277,N_14007);
xnor U15677 (N_15677,N_12581,N_13397);
nand U15678 (N_15678,N_14463,N_12791);
and U15679 (N_15679,N_12188,N_12908);
and U15680 (N_15680,N_14888,N_14194);
nor U15681 (N_15681,N_12077,N_12453);
nand U15682 (N_15682,N_14857,N_14326);
nand U15683 (N_15683,N_13270,N_12736);
nor U15684 (N_15684,N_14882,N_12690);
and U15685 (N_15685,N_13599,N_13033);
nand U15686 (N_15686,N_13906,N_13050);
xor U15687 (N_15687,N_14401,N_13536);
xor U15688 (N_15688,N_12482,N_12278);
nor U15689 (N_15689,N_14875,N_14637);
nor U15690 (N_15690,N_12762,N_13358);
xnor U15691 (N_15691,N_12170,N_13154);
xor U15692 (N_15692,N_14439,N_12910);
nor U15693 (N_15693,N_14038,N_14833);
or U15694 (N_15694,N_12845,N_14437);
nor U15695 (N_15695,N_14890,N_14106);
nor U15696 (N_15696,N_14842,N_14355);
nor U15697 (N_15697,N_13054,N_14457);
and U15698 (N_15698,N_13642,N_13946);
and U15699 (N_15699,N_13181,N_12969);
xor U15700 (N_15700,N_12347,N_13796);
nand U15701 (N_15701,N_14137,N_12151);
xor U15702 (N_15702,N_12193,N_12467);
and U15703 (N_15703,N_14973,N_12697);
and U15704 (N_15704,N_14719,N_12332);
nor U15705 (N_15705,N_14824,N_12502);
nand U15706 (N_15706,N_12824,N_13125);
xor U15707 (N_15707,N_14156,N_13236);
or U15708 (N_15708,N_14433,N_13653);
and U15709 (N_15709,N_13789,N_13579);
nor U15710 (N_15710,N_14189,N_14234);
nand U15711 (N_15711,N_12867,N_12596);
nor U15712 (N_15712,N_14646,N_13772);
xnor U15713 (N_15713,N_13365,N_13348);
nand U15714 (N_15714,N_14763,N_14685);
nor U15715 (N_15715,N_13755,N_14598);
xor U15716 (N_15716,N_13457,N_13925);
nor U15717 (N_15717,N_12425,N_13098);
and U15718 (N_15718,N_14773,N_13165);
and U15719 (N_15719,N_13670,N_13520);
nor U15720 (N_15720,N_13366,N_13821);
nand U15721 (N_15721,N_14410,N_12250);
xor U15722 (N_15722,N_14128,N_13850);
or U15723 (N_15723,N_12507,N_12734);
or U15724 (N_15724,N_14712,N_13403);
or U15725 (N_15725,N_13545,N_13211);
nor U15726 (N_15726,N_13069,N_12825);
nand U15727 (N_15727,N_14248,N_13883);
or U15728 (N_15728,N_12435,N_13531);
nor U15729 (N_15729,N_12731,N_14056);
nor U15730 (N_15730,N_12624,N_14164);
nand U15731 (N_15731,N_12764,N_13158);
or U15732 (N_15732,N_12592,N_13505);
nand U15733 (N_15733,N_14005,N_14115);
and U15734 (N_15734,N_14754,N_13940);
xnor U15735 (N_15735,N_13324,N_13918);
nand U15736 (N_15736,N_12924,N_13562);
nor U15737 (N_15737,N_13139,N_14383);
and U15738 (N_15738,N_13254,N_13766);
or U15739 (N_15739,N_13195,N_14484);
xor U15740 (N_15740,N_14673,N_12977);
nor U15741 (N_15741,N_12691,N_12967);
nor U15742 (N_15742,N_13334,N_14594);
or U15743 (N_15743,N_14751,N_12274);
nor U15744 (N_15744,N_13661,N_13583);
and U15745 (N_15745,N_14111,N_13196);
nand U15746 (N_15746,N_12850,N_12255);
nor U15747 (N_15747,N_13540,N_14337);
or U15748 (N_15748,N_13200,N_13016);
nor U15749 (N_15749,N_12940,N_14987);
xor U15750 (N_15750,N_12433,N_13719);
or U15751 (N_15751,N_14566,N_14354);
or U15752 (N_15752,N_14188,N_13448);
xor U15753 (N_15753,N_14227,N_12450);
nor U15754 (N_15754,N_14121,N_14778);
xor U15755 (N_15755,N_14210,N_12783);
or U15756 (N_15756,N_13419,N_14322);
and U15757 (N_15757,N_14942,N_13529);
and U15758 (N_15758,N_13097,N_13321);
and U15759 (N_15759,N_14886,N_13914);
nand U15760 (N_15760,N_13237,N_14311);
nand U15761 (N_15761,N_13126,N_14981);
xnor U15762 (N_15762,N_13471,N_12933);
nand U15763 (N_15763,N_12224,N_14200);
xor U15764 (N_15764,N_12578,N_13235);
or U15765 (N_15765,N_14664,N_12579);
and U15766 (N_15766,N_13989,N_13622);
nor U15767 (N_15767,N_13561,N_14900);
and U15768 (N_15768,N_13687,N_13615);
and U15769 (N_15769,N_13349,N_12158);
nand U15770 (N_15770,N_14116,N_13891);
nand U15771 (N_15771,N_12254,N_12357);
nor U15772 (N_15772,N_12457,N_14799);
nor U15773 (N_15773,N_12872,N_12728);
nand U15774 (N_15774,N_12587,N_13003);
and U15775 (N_15775,N_12430,N_13151);
and U15776 (N_15776,N_13000,N_13612);
or U15777 (N_15777,N_14514,N_14969);
and U15778 (N_15778,N_14975,N_13825);
nand U15779 (N_15779,N_14208,N_14236);
xor U15780 (N_15780,N_13356,N_14444);
and U15781 (N_15781,N_12754,N_14651);
and U15782 (N_15782,N_14940,N_14077);
nand U15783 (N_15783,N_14548,N_14288);
or U15784 (N_15784,N_14984,N_13034);
or U15785 (N_15785,N_14696,N_12059);
nand U15786 (N_15786,N_12288,N_14307);
nand U15787 (N_15787,N_12039,N_13679);
or U15788 (N_15788,N_12598,N_12827);
nor U15789 (N_15789,N_14385,N_12436);
or U15790 (N_15790,N_13027,N_12862);
and U15791 (N_15791,N_12564,N_12756);
and U15792 (N_15792,N_12842,N_14096);
nand U15793 (N_15793,N_14879,N_14085);
xor U15794 (N_15794,N_12407,N_12155);
nor U15795 (N_15795,N_14959,N_14359);
or U15796 (N_15796,N_12164,N_12383);
and U15797 (N_15797,N_12200,N_13967);
nand U15798 (N_15798,N_12110,N_12410);
or U15799 (N_15799,N_14652,N_14130);
nor U15800 (N_15800,N_14997,N_13802);
nor U15801 (N_15801,N_12931,N_14674);
or U15802 (N_15802,N_14703,N_13469);
or U15803 (N_15803,N_12062,N_13751);
xor U15804 (N_15804,N_12033,N_12732);
nand U15805 (N_15805,N_14087,N_14317);
xnor U15806 (N_15806,N_13175,N_13785);
xnor U15807 (N_15807,N_12695,N_13041);
nand U15808 (N_15808,N_12678,N_14897);
xnor U15809 (N_15809,N_14654,N_13464);
or U15810 (N_15810,N_12083,N_12094);
and U15811 (N_15811,N_12682,N_13010);
or U15812 (N_15812,N_13844,N_13557);
and U15813 (N_15813,N_13190,N_14701);
xnor U15814 (N_15814,N_14976,N_14516);
and U15815 (N_15815,N_13022,N_13406);
nand U15816 (N_15816,N_14209,N_12528);
nor U15817 (N_15817,N_13829,N_12971);
xor U15818 (N_15818,N_14737,N_13492);
and U15819 (N_15819,N_12053,N_13574);
and U15820 (N_15820,N_14643,N_13167);
xnor U15821 (N_15821,N_13571,N_13259);
xor U15822 (N_15822,N_12468,N_12558);
or U15823 (N_15823,N_13902,N_13299);
nor U15824 (N_15824,N_14771,N_12833);
or U15825 (N_15825,N_13724,N_14045);
nand U15826 (N_15826,N_14650,N_14344);
nand U15827 (N_15827,N_14212,N_12393);
xnor U15828 (N_15828,N_13450,N_12238);
or U15829 (N_15829,N_13705,N_14928);
and U15830 (N_15830,N_13488,N_12566);
nand U15831 (N_15831,N_13953,N_14321);
and U15832 (N_15832,N_12494,N_13411);
nand U15833 (N_15833,N_12167,N_14350);
nand U15834 (N_15834,N_13128,N_12195);
or U15835 (N_15835,N_14182,N_12476);
xor U15836 (N_15836,N_14510,N_12560);
nand U15837 (N_15837,N_13007,N_12542);
and U15838 (N_15838,N_14089,N_14496);
nor U15839 (N_15839,N_14172,N_13597);
nor U15840 (N_15840,N_13106,N_13836);
or U15841 (N_15841,N_13431,N_12513);
and U15842 (N_15842,N_12219,N_14856);
nor U15843 (N_15843,N_12689,N_14487);
nor U15844 (N_15844,N_12750,N_14766);
or U15845 (N_15845,N_13442,N_13312);
nand U15846 (N_15846,N_13550,N_12120);
and U15847 (N_15847,N_12960,N_14595);
nand U15848 (N_15848,N_12394,N_14345);
xor U15849 (N_15849,N_13451,N_12650);
nand U15850 (N_15850,N_14413,N_13628);
nor U15851 (N_15851,N_14505,N_13201);
xor U15852 (N_15852,N_13315,N_13178);
or U15853 (N_15853,N_13525,N_13952);
or U15854 (N_15854,N_12743,N_13739);
xnor U15855 (N_15855,N_12122,N_12466);
nor U15856 (N_15856,N_14129,N_14343);
xnor U15857 (N_15857,N_14691,N_14504);
and U15858 (N_15858,N_13286,N_13858);
xnor U15859 (N_15859,N_14564,N_13913);
nand U15860 (N_15860,N_13205,N_12554);
and U15861 (N_15861,N_13990,N_12870);
xnor U15862 (N_15862,N_13517,N_13942);
or U15863 (N_15863,N_14931,N_13570);
and U15864 (N_15864,N_13370,N_13759);
and U15865 (N_15865,N_14150,N_12797);
nand U15866 (N_15866,N_12025,N_13573);
xnor U15867 (N_15867,N_12814,N_13780);
nand U15868 (N_15868,N_12190,N_14447);
or U15869 (N_15869,N_13817,N_13645);
xor U15870 (N_15870,N_13594,N_12761);
nor U15871 (N_15871,N_13714,N_13189);
and U15872 (N_15872,N_13117,N_13208);
nor U15873 (N_15873,N_13135,N_13808);
nand U15874 (N_15874,N_13344,N_14979);
xor U15875 (N_15875,N_12378,N_13192);
xor U15876 (N_15876,N_12806,N_14170);
xor U15877 (N_15877,N_13138,N_14835);
nand U15878 (N_15878,N_13762,N_12173);
nand U15879 (N_15879,N_14822,N_13535);
or U15880 (N_15880,N_13119,N_13600);
nor U15881 (N_15881,N_14599,N_12559);
and U15882 (N_15882,N_14224,N_13402);
nor U15883 (N_15883,N_13014,N_12485);
xnor U15884 (N_15884,N_12086,N_14468);
and U15885 (N_15885,N_14113,N_14371);
nand U15886 (N_15886,N_13992,N_14411);
and U15887 (N_15887,N_14788,N_13301);
or U15888 (N_15888,N_14818,N_13585);
xor U15889 (N_15889,N_13606,N_12715);
xnor U15890 (N_15890,N_14065,N_14333);
or U15891 (N_15891,N_12524,N_14533);
and U15892 (N_15892,N_12156,N_13910);
xor U15893 (N_15893,N_13257,N_14552);
xnor U15894 (N_15894,N_14014,N_12649);
nor U15895 (N_15895,N_12857,N_12163);
and U15896 (N_15896,N_12738,N_12820);
nand U15897 (N_15897,N_14082,N_14908);
or U15898 (N_15898,N_14925,N_13718);
or U15899 (N_15899,N_14378,N_14183);
nand U15900 (N_15900,N_14911,N_13316);
nor U15901 (N_15901,N_14059,N_14813);
and U15902 (N_15902,N_14120,N_13987);
and U15903 (N_15903,N_14809,N_13839);
or U15904 (N_15904,N_14474,N_12223);
and U15905 (N_15905,N_13524,N_13085);
and U15906 (N_15906,N_14160,N_12243);
xor U15907 (N_15907,N_12324,N_12075);
or U15908 (N_15908,N_12662,N_12307);
and U15909 (N_15909,N_14304,N_14917);
or U15910 (N_15910,N_13162,N_12418);
xnor U15911 (N_15911,N_14966,N_14232);
and U15912 (N_15912,N_14889,N_12884);
xnor U15913 (N_15913,N_12264,N_12506);
and U15914 (N_15914,N_12245,N_12651);
and U15915 (N_15915,N_12118,N_13713);
nand U15916 (N_15916,N_13764,N_12321);
and U15917 (N_15917,N_13962,N_13293);
nand U15918 (N_15918,N_12868,N_14397);
and U15919 (N_15919,N_12209,N_12654);
nand U15920 (N_15920,N_14851,N_13647);
xnor U15921 (N_15921,N_12099,N_13300);
nand U15922 (N_15922,N_13640,N_14368);
nand U15923 (N_15923,N_14792,N_13706);
nand U15924 (N_15924,N_13008,N_13716);
nor U15925 (N_15925,N_14576,N_14294);
nor U15926 (N_15926,N_13305,N_12050);
xor U15927 (N_15927,N_12798,N_14490);
nand U15928 (N_15928,N_13875,N_12126);
nand U15929 (N_15929,N_13491,N_13340);
and U15930 (N_15930,N_14254,N_12815);
and U15931 (N_15931,N_14292,N_13039);
nor U15932 (N_15932,N_12247,N_13374);
or U15933 (N_15933,N_13611,N_13267);
or U15934 (N_15934,N_13292,N_12927);
or U15935 (N_15935,N_13882,N_14885);
or U15936 (N_15936,N_14093,N_13425);
nand U15937 (N_15937,N_13806,N_14774);
xnor U15938 (N_15938,N_13079,N_12017);
nand U15939 (N_15939,N_14849,N_13928);
or U15940 (N_15940,N_12221,N_13124);
xnor U15941 (N_15941,N_14012,N_13213);
and U15942 (N_15942,N_12944,N_14180);
xnor U15943 (N_15943,N_12898,N_13567);
nand U15944 (N_15944,N_14032,N_12474);
and U15945 (N_15945,N_12097,N_12159);
and U15946 (N_15946,N_14803,N_13893);
nor U15947 (N_15947,N_12225,N_13005);
or U15948 (N_15948,N_12354,N_13859);
or U15949 (N_15949,N_12994,N_13980);
nor U15950 (N_15950,N_14776,N_14723);
nor U15951 (N_15951,N_13553,N_14811);
and U15952 (N_15952,N_14524,N_12141);
nor U15953 (N_15953,N_13080,N_12656);
nor U15954 (N_15954,N_14223,N_13377);
or U15955 (N_15955,N_12011,N_13386);
xor U15956 (N_15956,N_13894,N_13793);
nand U15957 (N_15957,N_13680,N_13730);
xnor U15958 (N_15958,N_14079,N_13746);
xnor U15959 (N_15959,N_14493,N_12136);
xnor U15960 (N_15960,N_14458,N_12847);
nor U15961 (N_15961,N_14618,N_14756);
nand U15962 (N_15962,N_12081,N_14407);
or U15963 (N_15963,N_13870,N_12358);
xnor U15964 (N_15964,N_13616,N_12074);
nor U15965 (N_15965,N_13149,N_12172);
nand U15966 (N_15966,N_12470,N_14820);
or U15967 (N_15967,N_13791,N_14467);
or U15968 (N_15968,N_12175,N_14264);
nand U15969 (N_15969,N_14373,N_12829);
xnor U15970 (N_15970,N_14278,N_14728);
nor U15971 (N_15971,N_14752,N_13101);
nand U15972 (N_15972,N_14424,N_13876);
and U15973 (N_15973,N_12786,N_13447);
nor U15974 (N_15974,N_13782,N_14898);
nand U15975 (N_15975,N_12630,N_13444);
nand U15976 (N_15976,N_13061,N_14050);
and U15977 (N_15977,N_13376,N_14591);
nor U15978 (N_15978,N_12684,N_13380);
xor U15979 (N_15979,N_13133,N_13790);
or U15980 (N_15980,N_14377,N_12423);
xor U15981 (N_15981,N_14613,N_14779);
xnor U15982 (N_15982,N_14195,N_13276);
and U15983 (N_15983,N_12267,N_12217);
or U15984 (N_15984,N_13443,N_14048);
nand U15985 (N_15985,N_12693,N_13240);
xor U15986 (N_15986,N_13601,N_14657);
and U15987 (N_15987,N_13795,N_14090);
nor U15988 (N_15988,N_14145,N_12509);
nor U15989 (N_15989,N_13564,N_14092);
xnor U15990 (N_15990,N_12176,N_14781);
nor U15991 (N_15991,N_13900,N_14949);
or U15992 (N_15992,N_14151,N_12488);
xnor U15993 (N_15993,N_12272,N_12548);
xor U15994 (N_15994,N_12333,N_13960);
nand U15995 (N_15995,N_12414,N_13665);
nor U15996 (N_15996,N_12555,N_14679);
nand U15997 (N_15997,N_14909,N_13803);
xor U15998 (N_15998,N_13020,N_13833);
or U15999 (N_15999,N_14839,N_14815);
or U16000 (N_16000,N_13743,N_13463);
and U16001 (N_16001,N_12562,N_12283);
and U16002 (N_16002,N_13493,N_12113);
and U16003 (N_16003,N_13256,N_12452);
nor U16004 (N_16004,N_14954,N_13476);
and U16005 (N_16005,N_13379,N_13587);
or U16006 (N_16006,N_12128,N_14868);
or U16007 (N_16007,N_12635,N_12712);
nor U16008 (N_16008,N_14786,N_13278);
or U16009 (N_16009,N_14162,N_12973);
nor U16010 (N_16010,N_14834,N_14767);
or U16011 (N_16011,N_12028,N_12666);
xor U16012 (N_16012,N_13330,N_13846);
and U16013 (N_16013,N_14044,N_12104);
or U16014 (N_16014,N_12826,N_12539);
nand U16015 (N_16015,N_12934,N_13957);
nor U16016 (N_16016,N_12434,N_13881);
nand U16017 (N_16017,N_12603,N_13306);
nor U16018 (N_16018,N_14688,N_12883);
nor U16019 (N_16019,N_14816,N_14901);
nor U16020 (N_16020,N_14565,N_14899);
or U16021 (N_16021,N_14136,N_12349);
or U16022 (N_16022,N_13849,N_12445);
nor U16023 (N_16023,N_14996,N_12735);
nor U16024 (N_16024,N_14832,N_13949);
nor U16025 (N_16025,N_12729,N_13880);
nand U16026 (N_16026,N_13618,N_13255);
or U16027 (N_16027,N_12553,N_14119);
and U16028 (N_16028,N_14206,N_13961);
and U16029 (N_16029,N_13047,N_14309);
and U16030 (N_16030,N_13157,N_12129);
xnor U16031 (N_16031,N_12015,N_13907);
and U16032 (N_16032,N_13920,N_12983);
or U16033 (N_16033,N_12569,N_12605);
xnor U16034 (N_16034,N_12809,N_12595);
nand U16035 (N_16035,N_13396,N_13591);
nand U16036 (N_16036,N_14817,N_12896);
and U16037 (N_16037,N_12339,N_13666);
nor U16038 (N_16038,N_12717,N_12069);
nand U16039 (N_16039,N_13767,N_12495);
xor U16040 (N_16040,N_13404,N_13838);
nand U16041 (N_16041,N_13521,N_14393);
or U16042 (N_16042,N_12263,N_12805);
and U16043 (N_16043,N_13275,N_12591);
xor U16044 (N_16044,N_13991,N_14277);
and U16045 (N_16045,N_13996,N_12582);
nand U16046 (N_16046,N_12854,N_12700);
nor U16047 (N_16047,N_12030,N_14732);
or U16048 (N_16048,N_12478,N_12839);
nand U16049 (N_16049,N_12830,N_12660);
nand U16050 (N_16050,N_12115,N_12080);
nor U16051 (N_16051,N_14381,N_12796);
or U16052 (N_16052,N_14760,N_12618);
nand U16053 (N_16053,N_12331,N_12772);
xnor U16054 (N_16054,N_12493,N_13287);
nand U16055 (N_16055,N_13799,N_14026);
xor U16056 (N_16056,N_12239,N_12246);
and U16057 (N_16057,N_12813,N_12302);
or U16058 (N_16058,N_12541,N_13209);
nor U16059 (N_16059,N_12109,N_13416);
nor U16060 (N_16060,N_12611,N_12400);
and U16061 (N_16061,N_12710,N_13064);
nor U16062 (N_16062,N_12441,N_12510);
nor U16063 (N_16063,N_14830,N_14392);
nor U16064 (N_16064,N_13412,N_13389);
and U16065 (N_16065,N_14349,N_14770);
or U16066 (N_16066,N_14689,N_14095);
and U16067 (N_16067,N_12928,N_14023);
nand U16068 (N_16068,N_13509,N_13269);
and U16069 (N_16069,N_12297,N_14881);
xnor U16070 (N_16070,N_12515,N_12619);
nor U16071 (N_16071,N_13427,N_14729);
xor U16072 (N_16072,N_13588,N_12864);
xor U16073 (N_16073,N_12667,N_14692);
xnor U16074 (N_16074,N_14034,N_14366);
nor U16075 (N_16075,N_14039,N_14539);
nand U16076 (N_16076,N_12295,N_12363);
and U16077 (N_16077,N_14478,N_13664);
nor U16078 (N_16078,N_12103,N_12319);
nor U16079 (N_16079,N_13810,N_14300);
and U16080 (N_16080,N_13775,N_13589);
nor U16081 (N_16081,N_13288,N_14727);
xnor U16082 (N_16082,N_13260,N_12421);
xnor U16083 (N_16083,N_12670,N_13638);
nand U16084 (N_16084,N_13484,N_14049);
xnor U16085 (N_16085,N_13105,N_12088);
nor U16086 (N_16086,N_12518,N_12787);
or U16087 (N_16087,N_13613,N_12680);
and U16088 (N_16088,N_12133,N_12444);
xor U16089 (N_16089,N_12001,N_13083);
nor U16090 (N_16090,N_13350,N_14943);
nand U16091 (N_16091,N_14636,N_14528);
xor U16092 (N_16092,N_14998,N_13725);
or U16093 (N_16093,N_14971,N_12233);
xnor U16094 (N_16094,N_14866,N_13281);
and U16095 (N_16095,N_13841,N_14874);
or U16096 (N_16096,N_12948,N_13853);
nand U16097 (N_16097,N_14070,N_14363);
nand U16098 (N_16098,N_12491,N_14589);
or U16099 (N_16099,N_14179,N_13220);
nor U16100 (N_16100,N_14214,N_13051);
nand U16101 (N_16101,N_12538,N_13102);
xor U16102 (N_16102,N_13077,N_12636);
nand U16103 (N_16103,N_14247,N_13654);
or U16104 (N_16104,N_14844,N_12006);
xnor U16105 (N_16105,N_13076,N_14469);
xnor U16106 (N_16106,N_14739,N_13602);
and U16107 (N_16107,N_12606,N_14968);
nand U16108 (N_16108,N_13864,N_14859);
nand U16109 (N_16109,N_14698,N_14667);
and U16110 (N_16110,N_12957,N_12988);
nand U16111 (N_16111,N_13160,N_13333);
xor U16112 (N_16112,N_13297,N_14187);
nand U16113 (N_16113,N_13648,N_12497);
nor U16114 (N_16114,N_14351,N_14843);
nor U16115 (N_16115,N_13649,N_14498);
nor U16116 (N_16116,N_14205,N_13152);
or U16117 (N_16117,N_12454,N_12661);
nor U16118 (N_16118,N_13809,N_12389);
or U16119 (N_16119,N_14873,N_12526);
or U16120 (N_16120,N_12131,N_14139);
and U16121 (N_16121,N_13575,N_12076);
nor U16122 (N_16122,N_14346,N_13911);
nand U16123 (N_16123,N_13685,N_12937);
nand U16124 (N_16124,N_14621,N_14623);
and U16125 (N_16125,N_13596,N_13997);
and U16126 (N_16126,N_13556,N_13639);
nand U16127 (N_16127,N_13674,N_13381);
xnor U16128 (N_16128,N_12034,N_12882);
xnor U16129 (N_16129,N_12615,N_12178);
xor U16130 (N_16130,N_12706,N_12892);
xor U16131 (N_16131,N_14293,N_14918);
or U16132 (N_16132,N_12447,N_14481);
nor U16133 (N_16133,N_14060,N_14557);
or U16134 (N_16134,N_14489,N_14348);
or U16135 (N_16135,N_13865,N_14855);
or U16136 (N_16136,N_13378,N_14769);
and U16137 (N_16137,N_12147,N_14140);
xor U16138 (N_16138,N_12859,N_14336);
nor U16139 (N_16139,N_12379,N_14274);
and U16140 (N_16140,N_14884,N_12095);
or U16141 (N_16141,N_12585,N_14626);
xnor U16142 (N_16142,N_14471,N_12802);
or U16143 (N_16143,N_12597,N_12953);
xor U16144 (N_16144,N_12746,N_12091);
nand U16145 (N_16145,N_12019,N_12496);
or U16146 (N_16146,N_14053,N_13217);
xnor U16147 (N_16147,N_12885,N_14235);
or U16148 (N_16148,N_13483,N_14775);
nand U16149 (N_16149,N_13878,N_14127);
and U16150 (N_16150,N_12058,N_13863);
nor U16151 (N_16151,N_13210,N_14036);
nand U16152 (N_16152,N_12632,N_14861);
nor U16153 (N_16153,N_14043,N_14644);
and U16154 (N_16154,N_13619,N_14324);
nor U16155 (N_16155,N_14913,N_13672);
or U16156 (N_16156,N_14502,N_12742);
and U16157 (N_16157,N_14617,N_12314);
and U16158 (N_16158,N_12535,N_14331);
xnor U16159 (N_16159,N_12620,N_13777);
and U16160 (N_16160,N_12520,N_12671);
nand U16161 (N_16161,N_12206,N_12776);
and U16162 (N_16162,N_14725,N_14863);
or U16163 (N_16163,N_12107,N_12317);
nand U16164 (N_16164,N_13697,N_12723);
nand U16165 (N_16165,N_14253,N_14530);
nor U16166 (N_16166,N_12227,N_13818);
nand U16167 (N_16167,N_12415,N_13143);
nor U16168 (N_16168,N_14237,N_13708);
nand U16169 (N_16169,N_13428,N_14724);
nor U16170 (N_16170,N_12992,N_13176);
nor U16171 (N_16171,N_12021,N_13233);
or U16172 (N_16172,N_14951,N_13452);
nand U16173 (N_16173,N_12504,N_14400);
xnor U16174 (N_16174,N_14632,N_13018);
and U16175 (N_16175,N_12609,N_14905);
xnor U16176 (N_16176,N_14068,N_13609);
nand U16177 (N_16177,N_14483,N_12483);
xor U16178 (N_16178,N_13432,N_13440);
nand U16179 (N_16179,N_14627,N_14217);
nand U16180 (N_16180,N_14325,N_14736);
and U16181 (N_16181,N_13182,N_12241);
xnor U16182 (N_16182,N_14796,N_14244);
and U16183 (N_16183,N_12063,N_12674);
nand U16184 (N_16184,N_12550,N_12351);
xor U16185 (N_16185,N_14605,N_13368);
nor U16186 (N_16186,N_13656,N_12060);
nand U16187 (N_16187,N_13693,N_13515);
xnor U16188 (N_16188,N_12523,N_13383);
nand U16189 (N_16189,N_13823,N_14948);
nand U16190 (N_16190,N_12724,N_13955);
nand U16191 (N_16191,N_12625,N_14057);
nor U16192 (N_16192,N_12036,N_14360);
or U16193 (N_16193,N_14519,N_12489);
and U16194 (N_16194,N_13127,N_13629);
or U16195 (N_16195,N_14677,N_14273);
and U16196 (N_16196,N_12945,N_12552);
xnor U16197 (N_16197,N_12920,N_12590);
and U16198 (N_16198,N_14341,N_13229);
nor U16199 (N_16199,N_14108,N_12365);
nor U16200 (N_16200,N_14511,N_13873);
nand U16201 (N_16201,N_12007,N_13752);
or U16202 (N_16202,N_12759,N_13726);
or U16203 (N_16203,N_12348,N_13355);
or U16204 (N_16204,N_13132,N_13537);
and U16205 (N_16205,N_14313,N_12769);
nand U16206 (N_16206,N_14303,N_14448);
xor U16207 (N_16207,N_14052,N_13062);
and U16208 (N_16208,N_13972,N_12887);
and U16209 (N_16209,N_12614,N_12869);
and U16210 (N_16210,N_14011,N_14570);
and U16211 (N_16211,N_13361,N_14957);
and U16212 (N_16212,N_12672,N_14656);
xor U16213 (N_16213,N_13944,N_12999);
xnor U16214 (N_16214,N_12789,N_12166);
xnor U16215 (N_16215,N_13468,N_13669);
or U16216 (N_16216,N_14755,N_14745);
nor U16217 (N_16217,N_12116,N_14152);
nand U16218 (N_16218,N_12880,N_13908);
xor U16219 (N_16219,N_13512,N_12149);
nor U16220 (N_16220,N_13769,N_12181);
nor U16221 (N_16221,N_13004,N_13066);
or U16222 (N_16222,N_12305,N_14103);
or U16223 (N_16223,N_12664,N_13142);
nor U16224 (N_16224,N_12282,N_14926);
nand U16225 (N_16225,N_14058,N_13336);
nor U16226 (N_16226,N_13496,N_12888);
nand U16227 (N_16227,N_12583,N_14099);
xor U16228 (N_16228,N_13060,N_14690);
and U16229 (N_16229,N_12490,N_13856);
or U16230 (N_16230,N_12665,N_14122);
or U16231 (N_16231,N_14167,N_13625);
nand U16232 (N_16232,N_12821,N_13861);
or U16233 (N_16233,N_14334,N_12768);
xnor U16234 (N_16234,N_13055,N_14532);
nor U16235 (N_16235,N_14645,N_14131);
nor U16236 (N_16236,N_14181,N_14157);
and U16237 (N_16237,N_14472,N_13889);
and U16238 (N_16238,N_14553,N_12795);
and U16239 (N_16239,N_13765,N_13388);
nor U16240 (N_16240,N_13652,N_13927);
or U16241 (N_16241,N_14927,N_14153);
nand U16242 (N_16242,N_12132,N_13073);
and U16243 (N_16243,N_14507,N_14175);
xor U16244 (N_16244,N_14693,N_13951);
nor U16245 (N_16245,N_13107,N_12681);
nand U16246 (N_16246,N_14517,N_14201);
or U16247 (N_16247,N_13637,N_14887);
and U16248 (N_16248,N_13353,N_14709);
nand U16249 (N_16249,N_14906,N_12018);
and U16250 (N_16250,N_12143,N_13197);
nand U16251 (N_16251,N_12270,N_12607);
nand U16252 (N_16252,N_12065,N_13026);
xor U16253 (N_16253,N_12290,N_14455);
and U16254 (N_16254,N_14138,N_13429);
nor U16255 (N_16255,N_12009,N_12629);
nor U16256 (N_16256,N_13811,N_13551);
and U16257 (N_16257,N_13617,N_13030);
xnor U16258 (N_16258,N_14229,N_14323);
xor U16259 (N_16259,N_12355,N_13729);
or U16260 (N_16260,N_13926,N_12046);
nand U16261 (N_16261,N_13161,N_14074);
or U16262 (N_16262,N_14166,N_14421);
nand U16263 (N_16263,N_13750,N_14456);
and U16264 (N_16264,N_12463,N_12084);
xnor U16265 (N_16265,N_12793,N_12503);
nor U16266 (N_16266,N_14379,N_13103);
or U16267 (N_16267,N_14810,N_13502);
xor U16268 (N_16268,N_14660,N_14021);
or U16269 (N_16269,N_12401,N_13040);
and U16270 (N_16270,N_12679,N_14920);
xor U16271 (N_16271,N_12481,N_12512);
or U16272 (N_16272,N_14912,N_12701);
nor U16273 (N_16273,N_14537,N_13194);
and U16274 (N_16274,N_13738,N_12399);
xor U16275 (N_16275,N_14748,N_13526);
xnor U16276 (N_16276,N_13011,N_12182);
or U16277 (N_16277,N_12551,N_13223);
nand U16278 (N_16278,N_13470,N_14335);
nor U16279 (N_16279,N_14798,N_13423);
nor U16280 (N_16280,N_12153,N_14512);
and U16281 (N_16281,N_14271,N_12639);
nor U16282 (N_16282,N_13375,N_12072);
nand U16283 (N_16283,N_13845,N_12165);
nor U16284 (N_16284,N_13510,N_12368);
nor U16285 (N_16285,N_14018,N_14491);
and U16286 (N_16286,N_14428,N_14289);
or U16287 (N_16287,N_14388,N_13437);
and U16288 (N_16288,N_12964,N_13635);
and U16289 (N_16289,N_12335,N_13234);
and U16290 (N_16290,N_12818,N_14513);
nand U16291 (N_16291,N_13506,N_13650);
nor U16292 (N_16292,N_13466,N_12871);
xnor U16293 (N_16293,N_13015,N_12705);
nor U16294 (N_16294,N_14291,N_14384);
and U16295 (N_16295,N_12061,N_12073);
or U16296 (N_16296,N_14495,N_13919);
or U16297 (N_16297,N_12426,N_13655);
or U16298 (N_16298,N_14126,N_13580);
and U16299 (N_16299,N_14992,N_13909);
nor U16300 (N_16300,N_12024,N_12522);
nor U16301 (N_16301,N_13185,N_13523);
nor U16302 (N_16302,N_12000,N_12713);
and U16303 (N_16303,N_13771,N_12286);
or U16304 (N_16304,N_14506,N_12529);
nor U16305 (N_16305,N_12334,N_14733);
xnor U16306 (N_16306,N_14790,N_14525);
or U16307 (N_16307,N_12873,N_14315);
nor U16308 (N_16308,N_13621,N_13915);
nor U16309 (N_16309,N_13917,N_13057);
and U16310 (N_16310,N_14982,N_13159);
nor U16311 (N_16311,N_12899,N_13805);
xor U16312 (N_16312,N_14862,N_13543);
nand U16313 (N_16313,N_13852,N_14761);
xnor U16314 (N_16314,N_12045,N_13646);
or U16315 (N_16315,N_12770,N_12023);
xnor U16316 (N_16316,N_14362,N_13547);
xor U16317 (N_16317,N_14600,N_12101);
and U16318 (N_16318,N_13112,N_13943);
or U16319 (N_16319,N_12633,N_14978);
and U16320 (N_16320,N_12985,N_14544);
xnor U16321 (N_16321,N_14276,N_12374);
nor U16322 (N_16322,N_13501,N_13329);
and U16323 (N_16323,N_13768,N_14670);
nand U16324 (N_16324,N_14631,N_13042);
nand U16325 (N_16325,N_13395,N_14655);
and U16326 (N_16326,N_13800,N_13659);
nor U16327 (N_16327,N_14062,N_14112);
nor U16328 (N_16328,N_13141,N_14869);
or U16329 (N_16329,N_13528,N_14027);
or U16330 (N_16330,N_13410,N_12424);
nor U16331 (N_16331,N_12248,N_12727);
nand U16332 (N_16332,N_13608,N_13500);
xnor U16333 (N_16333,N_13279,N_12616);
xor U16334 (N_16334,N_12135,N_14980);
nand U16335 (N_16335,N_12484,N_13347);
nor U16336 (N_16336,N_12837,N_13148);
nand U16337 (N_16337,N_13626,N_12501);
xor U16338 (N_16338,N_14054,N_14061);
nand U16339 (N_16339,N_14614,N_14144);
nor U16340 (N_16340,N_12380,N_14101);
nand U16341 (N_16341,N_13973,N_13816);
nand U16342 (N_16342,N_13783,N_14067);
or U16343 (N_16343,N_13298,N_14877);
nand U16344 (N_16344,N_12576,N_13188);
and U16345 (N_16345,N_12048,N_14716);
xor U16346 (N_16346,N_13956,N_14124);
or U16347 (N_16347,N_12594,N_14612);
nand U16348 (N_16348,N_13581,N_12273);
or U16349 (N_16349,N_13866,N_13110);
nor U16350 (N_16350,N_14720,N_14207);
and U16351 (N_16351,N_12790,N_14450);
or U16352 (N_16352,N_14520,N_12105);
or U16353 (N_16353,N_14845,N_14847);
xor U16354 (N_16354,N_12026,N_12703);
xor U16355 (N_16355,N_14921,N_13681);
nor U16356 (N_16356,N_13044,N_13099);
or U16357 (N_16357,N_14678,N_12479);
and U16358 (N_16358,N_12417,N_13758);
nand U16359 (N_16359,N_12475,N_12687);
xor U16360 (N_16360,N_12531,N_13394);
xnor U16361 (N_16361,N_12391,N_12390);
or U16362 (N_16362,N_12567,N_14575);
xnor U16363 (N_16363,N_13434,N_14965);
xor U16364 (N_16364,N_12725,N_12344);
and U16365 (N_16365,N_12292,N_14521);
or U16366 (N_16366,N_12236,N_14178);
or U16367 (N_16367,N_12979,N_13998);
nand U16368 (N_16368,N_12313,N_14932);
nand U16369 (N_16369,N_12807,N_14019);
xnor U16370 (N_16370,N_14840,N_12256);
xor U16371 (N_16371,N_14742,N_13848);
or U16372 (N_16372,N_13533,N_14008);
nor U16373 (N_16373,N_14423,N_12737);
xnor U16374 (N_16374,N_13081,N_14758);
nand U16375 (N_16375,N_14960,N_12866);
xor U16376 (N_16376,N_13091,N_13728);
and U16377 (N_16377,N_13487,N_12134);
xor U16378 (N_16378,N_12352,N_13749);
nor U16379 (N_16379,N_14185,N_12056);
nand U16380 (N_16380,N_12448,N_12299);
and U16381 (N_16381,N_14416,N_14149);
or U16382 (N_16382,N_14158,N_14066);
nor U16383 (N_16383,N_13843,N_12275);
xor U16384 (N_16384,N_12514,N_13984);
or U16385 (N_16385,N_13147,N_14534);
or U16386 (N_16386,N_14597,N_13604);
xor U16387 (N_16387,N_13886,N_14358);
and U16388 (N_16388,N_14438,N_14395);
nor U16389 (N_16389,N_13559,N_13291);
or U16390 (N_16390,N_14003,N_12142);
or U16391 (N_16391,N_13686,N_12265);
nand U16392 (N_16392,N_14582,N_13177);
xnor U16393 (N_16393,N_12532,N_12404);
nand U16394 (N_16394,N_12214,N_14642);
nand U16395 (N_16395,N_12477,N_12366);
or U16396 (N_16396,N_14933,N_14950);
xnor U16397 (N_16397,N_14584,N_13632);
or U16398 (N_16398,N_12719,N_14894);
xor U16399 (N_16399,N_14515,N_14825);
nor U16400 (N_16400,N_13610,N_12405);
xor U16401 (N_16401,N_14262,N_14286);
and U16402 (N_16402,N_13369,N_13212);
nor U16403 (N_16403,N_13888,N_14033);
and U16404 (N_16404,N_12361,N_13382);
and U16405 (N_16405,N_12403,N_13373);
or U16406 (N_16406,N_12708,N_12699);
and U16407 (N_16407,N_14970,N_12338);
or U16408 (N_16408,N_12894,N_13577);
and U16409 (N_16409,N_12057,N_14704);
xnor U16410 (N_16410,N_14258,N_13294);
or U16411 (N_16411,N_12171,N_13937);
or U16412 (N_16412,N_13598,N_12154);
and U16413 (N_16413,N_14146,N_13271);
nor U16414 (N_16414,N_12189,N_14226);
xnor U16415 (N_16415,N_12473,N_12121);
or U16416 (N_16416,N_13733,N_14287);
nand U16417 (N_16417,N_13071,N_14675);
nor U16418 (N_16418,N_12032,N_13947);
nor U16419 (N_16419,N_12253,N_13289);
and U16420 (N_16420,N_14299,N_12281);
and U16421 (N_16421,N_13215,N_14808);
xor U16422 (N_16422,N_13359,N_12451);
or U16423 (N_16423,N_14249,N_14266);
and U16424 (N_16424,N_13731,N_12197);
or U16425 (N_16425,N_12902,N_13302);
nor U16426 (N_16426,N_12777,N_13393);
xnor U16427 (N_16427,N_14449,N_14726);
nand U16428 (N_16428,N_13590,N_12123);
xnor U16429 (N_16429,N_12752,N_13582);
xnor U16430 (N_16430,N_13249,N_13092);
or U16431 (N_16431,N_13904,N_14473);
and U16432 (N_16432,N_13221,N_12373);
and U16433 (N_16433,N_14699,N_14270);
nor U16434 (N_16434,N_12325,N_14147);
xor U16435 (N_16435,N_12229,N_12915);
nand U16436 (N_16436,N_13595,N_12584);
nor U16437 (N_16437,N_13166,N_13631);
or U16438 (N_16438,N_14999,N_12005);
xnor U16439 (N_16439,N_13572,N_13179);
nand U16440 (N_16440,N_14784,N_14629);
xor U16441 (N_16441,N_12336,N_13813);
and U16442 (N_16442,N_14417,N_14387);
nand U16443 (N_16443,N_12342,N_13924);
xnor U16444 (N_16444,N_12926,N_12711);
and U16445 (N_16445,N_13013,N_12840);
nand U16446 (N_16446,N_14414,N_12741);
and U16447 (N_16447,N_12465,N_13732);
or U16448 (N_16448,N_13539,N_12991);
or U16449 (N_16449,N_14046,N_13692);
nand U16450 (N_16450,N_12035,N_13774);
nand U16451 (N_16451,N_14941,N_13400);
xnor U16452 (N_16452,N_13754,N_12362);
xor U16453 (N_16453,N_14883,N_12180);
xor U16454 (N_16454,N_12315,N_13814);
and U16455 (N_16455,N_12601,N_12412);
nor U16456 (N_16456,N_13088,N_12525);
and U16457 (N_16457,N_13903,N_14743);
and U16458 (N_16458,N_14432,N_13658);
and U16459 (N_16459,N_13295,N_14041);
or U16460 (N_16460,N_12755,N_12577);
nor U16461 (N_16461,N_12917,N_13421);
nand U16462 (N_16462,N_12851,N_14114);
xnor U16463 (N_16463,N_14239,N_14503);
nor U16464 (N_16464,N_12370,N_12921);
xnor U16465 (N_16465,N_12561,N_13691);
xnor U16466 (N_16466,N_13700,N_13094);
nand U16467 (N_16467,N_12198,N_12038);
xnor U16468 (N_16468,N_14073,N_12819);
and U16469 (N_16469,N_12874,N_13180);
xor U16470 (N_16470,N_12637,N_12612);
nor U16471 (N_16471,N_12262,N_12604);
nor U16472 (N_16472,N_13636,N_13096);
or U16473 (N_16473,N_13643,N_14876);
or U16474 (N_16474,N_12685,N_14989);
and U16475 (N_16475,N_14538,N_14298);
or U16476 (N_16476,N_12861,N_13477);
or U16477 (N_16477,N_13832,N_12989);
nand U16478 (N_16478,N_12832,N_13644);
and U16479 (N_16479,N_13709,N_13634);
nor U16480 (N_16480,N_14425,N_14694);
xnor U16481 (N_16481,N_13467,N_12676);
nand U16482 (N_16482,N_14561,N_13565);
or U16483 (N_16483,N_13820,N_13430);
xnor U16484 (N_16484,N_14802,N_13065);
nand U16485 (N_16485,N_14367,N_13282);
and U16486 (N_16486,N_12168,N_14902);
or U16487 (N_16487,N_13284,N_12784);
xnor U16488 (N_16488,N_13363,N_12853);
nand U16489 (N_16489,N_12757,N_14549);
nand U16490 (N_16490,N_12704,N_13558);
xnor U16491 (N_16491,N_12740,N_13827);
xnor U16492 (N_16492,N_14028,N_13549);
nand U16493 (N_16493,N_12460,N_14155);
or U16494 (N_16494,N_13045,N_12067);
xnor U16495 (N_16495,N_12652,N_14376);
and U16496 (N_16496,N_13320,N_14606);
nor U16497 (N_16497,N_14619,N_13093);
and U16498 (N_16498,N_13897,N_12865);
nor U16499 (N_16499,N_14142,N_12593);
and U16500 (N_16500,N_12570,N_12092);
xnor U16501 (N_16501,N_14123,N_14135);
or U16502 (N_16502,N_12008,N_14403);
nand U16503 (N_16503,N_13230,N_14558);
nor U16504 (N_16504,N_12682,N_12840);
or U16505 (N_16505,N_13478,N_14286);
nand U16506 (N_16506,N_12116,N_13541);
nor U16507 (N_16507,N_12134,N_14137);
nor U16508 (N_16508,N_12783,N_13921);
or U16509 (N_16509,N_13600,N_13299);
or U16510 (N_16510,N_12234,N_14215);
nor U16511 (N_16511,N_12357,N_13339);
nor U16512 (N_16512,N_12845,N_14334);
nor U16513 (N_16513,N_13156,N_14893);
nor U16514 (N_16514,N_14522,N_14611);
or U16515 (N_16515,N_12025,N_12304);
nor U16516 (N_16516,N_13723,N_14416);
and U16517 (N_16517,N_14948,N_12768);
xor U16518 (N_16518,N_12141,N_12479);
xnor U16519 (N_16519,N_13653,N_14701);
and U16520 (N_16520,N_13529,N_14185);
nor U16521 (N_16521,N_14092,N_13916);
nand U16522 (N_16522,N_14972,N_13886);
and U16523 (N_16523,N_14606,N_12560);
nor U16524 (N_16524,N_13352,N_13016);
and U16525 (N_16525,N_14514,N_13430);
nand U16526 (N_16526,N_12051,N_14164);
xnor U16527 (N_16527,N_14661,N_14602);
and U16528 (N_16528,N_14553,N_14686);
nor U16529 (N_16529,N_13714,N_13437);
nand U16530 (N_16530,N_12062,N_14949);
xor U16531 (N_16531,N_13463,N_13438);
nand U16532 (N_16532,N_12085,N_12572);
xor U16533 (N_16533,N_12277,N_14393);
nor U16534 (N_16534,N_13522,N_12347);
xor U16535 (N_16535,N_14763,N_14396);
nand U16536 (N_16536,N_13730,N_13168);
nand U16537 (N_16537,N_12539,N_13882);
or U16538 (N_16538,N_14780,N_12405);
and U16539 (N_16539,N_12962,N_14339);
and U16540 (N_16540,N_13115,N_14128);
or U16541 (N_16541,N_14018,N_13933);
nand U16542 (N_16542,N_13164,N_14875);
and U16543 (N_16543,N_13810,N_14551);
xnor U16544 (N_16544,N_13899,N_13676);
or U16545 (N_16545,N_12708,N_12288);
nor U16546 (N_16546,N_12885,N_13265);
nand U16547 (N_16547,N_14512,N_14333);
xnor U16548 (N_16548,N_12311,N_12025);
nor U16549 (N_16549,N_14745,N_13007);
xor U16550 (N_16550,N_13231,N_13435);
xor U16551 (N_16551,N_14033,N_14408);
and U16552 (N_16552,N_14733,N_13655);
or U16553 (N_16553,N_14998,N_12076);
nand U16554 (N_16554,N_14662,N_12182);
nor U16555 (N_16555,N_14476,N_14816);
or U16556 (N_16556,N_14057,N_13965);
nand U16557 (N_16557,N_12077,N_13977);
and U16558 (N_16558,N_12090,N_12909);
or U16559 (N_16559,N_13806,N_12185);
nand U16560 (N_16560,N_14423,N_12709);
nor U16561 (N_16561,N_14475,N_13770);
and U16562 (N_16562,N_14111,N_14430);
nand U16563 (N_16563,N_13752,N_14949);
and U16564 (N_16564,N_12250,N_14186);
nand U16565 (N_16565,N_14763,N_13931);
nand U16566 (N_16566,N_13935,N_12099);
nor U16567 (N_16567,N_14982,N_14642);
nand U16568 (N_16568,N_14225,N_14376);
nand U16569 (N_16569,N_14786,N_13936);
nor U16570 (N_16570,N_13158,N_13677);
or U16571 (N_16571,N_14287,N_12002);
nor U16572 (N_16572,N_14423,N_14106);
nor U16573 (N_16573,N_12393,N_14529);
or U16574 (N_16574,N_12914,N_13542);
and U16575 (N_16575,N_12336,N_12374);
nor U16576 (N_16576,N_12951,N_14535);
and U16577 (N_16577,N_12626,N_12223);
nor U16578 (N_16578,N_13032,N_12822);
nor U16579 (N_16579,N_12016,N_13986);
nor U16580 (N_16580,N_12407,N_13261);
and U16581 (N_16581,N_12128,N_12361);
nor U16582 (N_16582,N_12285,N_14862);
xnor U16583 (N_16583,N_13572,N_14143);
and U16584 (N_16584,N_12329,N_12164);
nand U16585 (N_16585,N_12604,N_14716);
nor U16586 (N_16586,N_13596,N_12161);
nor U16587 (N_16587,N_14742,N_12984);
nand U16588 (N_16588,N_12909,N_13150);
xnor U16589 (N_16589,N_14656,N_14721);
nor U16590 (N_16590,N_12299,N_12974);
xnor U16591 (N_16591,N_12396,N_12951);
and U16592 (N_16592,N_13823,N_12124);
or U16593 (N_16593,N_12774,N_12779);
xnor U16594 (N_16594,N_14641,N_13934);
or U16595 (N_16595,N_13994,N_12126);
nand U16596 (N_16596,N_13752,N_12611);
or U16597 (N_16597,N_12380,N_14344);
and U16598 (N_16598,N_12299,N_12104);
and U16599 (N_16599,N_14042,N_14175);
nor U16600 (N_16600,N_13943,N_14520);
nand U16601 (N_16601,N_13236,N_13411);
nand U16602 (N_16602,N_14095,N_13821);
nand U16603 (N_16603,N_13539,N_14415);
nand U16604 (N_16604,N_14131,N_13533);
xnor U16605 (N_16605,N_14511,N_13613);
xor U16606 (N_16606,N_14588,N_14156);
nor U16607 (N_16607,N_12391,N_14161);
and U16608 (N_16608,N_12033,N_14194);
xnor U16609 (N_16609,N_13387,N_13638);
and U16610 (N_16610,N_14578,N_14074);
and U16611 (N_16611,N_13217,N_13813);
nand U16612 (N_16612,N_14079,N_13621);
and U16613 (N_16613,N_14169,N_13016);
or U16614 (N_16614,N_13709,N_12042);
xor U16615 (N_16615,N_14871,N_14498);
nor U16616 (N_16616,N_13084,N_12147);
or U16617 (N_16617,N_13276,N_13842);
or U16618 (N_16618,N_13233,N_13852);
or U16619 (N_16619,N_12550,N_13668);
and U16620 (N_16620,N_12387,N_13274);
or U16621 (N_16621,N_13994,N_13619);
or U16622 (N_16622,N_13078,N_13351);
and U16623 (N_16623,N_13790,N_12283);
xor U16624 (N_16624,N_13476,N_13545);
nand U16625 (N_16625,N_13857,N_13844);
nor U16626 (N_16626,N_13155,N_12485);
and U16627 (N_16627,N_13337,N_12417);
and U16628 (N_16628,N_14218,N_14101);
nand U16629 (N_16629,N_12949,N_14275);
and U16630 (N_16630,N_12598,N_12707);
xor U16631 (N_16631,N_13246,N_12461);
xnor U16632 (N_16632,N_14170,N_13283);
or U16633 (N_16633,N_13925,N_13074);
nor U16634 (N_16634,N_13385,N_13736);
or U16635 (N_16635,N_13909,N_12403);
nor U16636 (N_16636,N_12442,N_14445);
nor U16637 (N_16637,N_12637,N_13533);
and U16638 (N_16638,N_13486,N_14546);
and U16639 (N_16639,N_12569,N_14865);
nand U16640 (N_16640,N_13375,N_13961);
xnor U16641 (N_16641,N_13733,N_13728);
xor U16642 (N_16642,N_14253,N_12150);
or U16643 (N_16643,N_12594,N_12648);
nand U16644 (N_16644,N_14030,N_14773);
and U16645 (N_16645,N_12217,N_12641);
and U16646 (N_16646,N_14528,N_14299);
xor U16647 (N_16647,N_13648,N_14918);
or U16648 (N_16648,N_14968,N_13189);
nor U16649 (N_16649,N_12650,N_13188);
and U16650 (N_16650,N_14658,N_13096);
nand U16651 (N_16651,N_12839,N_13661);
xnor U16652 (N_16652,N_13772,N_14792);
nand U16653 (N_16653,N_13491,N_13589);
or U16654 (N_16654,N_13732,N_14818);
and U16655 (N_16655,N_14518,N_13789);
or U16656 (N_16656,N_14107,N_12281);
or U16657 (N_16657,N_13864,N_13442);
nand U16658 (N_16658,N_14627,N_13431);
and U16659 (N_16659,N_12449,N_14894);
nand U16660 (N_16660,N_12904,N_14756);
xor U16661 (N_16661,N_12742,N_14715);
and U16662 (N_16662,N_12386,N_12011);
or U16663 (N_16663,N_13273,N_13787);
and U16664 (N_16664,N_12888,N_14466);
and U16665 (N_16665,N_13243,N_12658);
xor U16666 (N_16666,N_13516,N_14611);
nand U16667 (N_16667,N_13539,N_14911);
or U16668 (N_16668,N_13982,N_13571);
nand U16669 (N_16669,N_13603,N_12914);
nand U16670 (N_16670,N_12828,N_13220);
nand U16671 (N_16671,N_13908,N_13578);
xnor U16672 (N_16672,N_13891,N_14922);
or U16673 (N_16673,N_14427,N_13681);
xnor U16674 (N_16674,N_14808,N_14508);
nor U16675 (N_16675,N_13133,N_12501);
nor U16676 (N_16676,N_14220,N_13333);
xnor U16677 (N_16677,N_12656,N_14324);
nor U16678 (N_16678,N_12158,N_12193);
and U16679 (N_16679,N_12724,N_13499);
and U16680 (N_16680,N_14694,N_13461);
or U16681 (N_16681,N_14393,N_14302);
nor U16682 (N_16682,N_13941,N_13978);
xnor U16683 (N_16683,N_12314,N_14818);
xor U16684 (N_16684,N_12693,N_12088);
nor U16685 (N_16685,N_13370,N_14716);
or U16686 (N_16686,N_13382,N_12529);
or U16687 (N_16687,N_14405,N_13147);
xor U16688 (N_16688,N_14313,N_14004);
or U16689 (N_16689,N_13911,N_12536);
xnor U16690 (N_16690,N_13995,N_14935);
nor U16691 (N_16691,N_13915,N_14622);
or U16692 (N_16692,N_14351,N_13539);
xnor U16693 (N_16693,N_14861,N_14745);
xnor U16694 (N_16694,N_14315,N_14375);
nor U16695 (N_16695,N_13466,N_14863);
xnor U16696 (N_16696,N_14038,N_12725);
or U16697 (N_16697,N_13859,N_13605);
or U16698 (N_16698,N_12192,N_12563);
or U16699 (N_16699,N_14067,N_13474);
and U16700 (N_16700,N_14287,N_14070);
xnor U16701 (N_16701,N_12041,N_14357);
nand U16702 (N_16702,N_12455,N_12254);
and U16703 (N_16703,N_12567,N_14650);
xnor U16704 (N_16704,N_13792,N_14957);
xnor U16705 (N_16705,N_14289,N_13321);
nand U16706 (N_16706,N_14501,N_14430);
xnor U16707 (N_16707,N_14722,N_12570);
nor U16708 (N_16708,N_12984,N_12125);
or U16709 (N_16709,N_14695,N_13764);
or U16710 (N_16710,N_12070,N_12469);
nand U16711 (N_16711,N_14766,N_12262);
nor U16712 (N_16712,N_14212,N_14875);
nor U16713 (N_16713,N_14573,N_13449);
xor U16714 (N_16714,N_13832,N_12045);
or U16715 (N_16715,N_13880,N_12387);
or U16716 (N_16716,N_12243,N_12693);
nor U16717 (N_16717,N_13265,N_13796);
and U16718 (N_16718,N_12398,N_12092);
xnor U16719 (N_16719,N_14963,N_12952);
and U16720 (N_16720,N_13981,N_14392);
nand U16721 (N_16721,N_14757,N_12600);
and U16722 (N_16722,N_12877,N_14644);
or U16723 (N_16723,N_14003,N_14168);
and U16724 (N_16724,N_13145,N_14701);
and U16725 (N_16725,N_13241,N_13138);
xnor U16726 (N_16726,N_13767,N_14676);
nor U16727 (N_16727,N_13734,N_12374);
xnor U16728 (N_16728,N_14653,N_14369);
xor U16729 (N_16729,N_14562,N_12138);
nor U16730 (N_16730,N_13050,N_14642);
xnor U16731 (N_16731,N_13566,N_13830);
nor U16732 (N_16732,N_12323,N_12377);
nand U16733 (N_16733,N_13235,N_14899);
nor U16734 (N_16734,N_14509,N_12346);
nand U16735 (N_16735,N_14599,N_14099);
and U16736 (N_16736,N_14204,N_14816);
and U16737 (N_16737,N_12000,N_14088);
or U16738 (N_16738,N_12468,N_12644);
and U16739 (N_16739,N_14990,N_14265);
nand U16740 (N_16740,N_14006,N_13754);
nor U16741 (N_16741,N_14763,N_12097);
or U16742 (N_16742,N_12389,N_14057);
and U16743 (N_16743,N_12136,N_13377);
or U16744 (N_16744,N_12799,N_13107);
or U16745 (N_16745,N_13993,N_13617);
or U16746 (N_16746,N_14272,N_12822);
and U16747 (N_16747,N_14621,N_13020);
xnor U16748 (N_16748,N_14328,N_12978);
xnor U16749 (N_16749,N_12043,N_13468);
nand U16750 (N_16750,N_12130,N_12970);
xnor U16751 (N_16751,N_13410,N_13012);
and U16752 (N_16752,N_12668,N_12816);
nor U16753 (N_16753,N_12563,N_12089);
nand U16754 (N_16754,N_12291,N_12033);
nand U16755 (N_16755,N_12143,N_13666);
xor U16756 (N_16756,N_13294,N_12767);
nor U16757 (N_16757,N_13413,N_13407);
nor U16758 (N_16758,N_12859,N_13215);
nor U16759 (N_16759,N_13737,N_12956);
nor U16760 (N_16760,N_13947,N_13226);
and U16761 (N_16761,N_13886,N_14063);
nand U16762 (N_16762,N_12048,N_14052);
and U16763 (N_16763,N_13575,N_14418);
nand U16764 (N_16764,N_13867,N_14856);
nand U16765 (N_16765,N_12810,N_12208);
nand U16766 (N_16766,N_14772,N_13454);
nor U16767 (N_16767,N_14352,N_13667);
or U16768 (N_16768,N_13573,N_14241);
xnor U16769 (N_16769,N_12212,N_12194);
xor U16770 (N_16770,N_12596,N_13198);
nor U16771 (N_16771,N_14590,N_12295);
and U16772 (N_16772,N_13986,N_12336);
nor U16773 (N_16773,N_12230,N_14500);
xnor U16774 (N_16774,N_13705,N_14454);
nor U16775 (N_16775,N_14384,N_14975);
nor U16776 (N_16776,N_12639,N_12774);
nand U16777 (N_16777,N_13740,N_13222);
nand U16778 (N_16778,N_14186,N_13635);
xnor U16779 (N_16779,N_13826,N_12243);
and U16780 (N_16780,N_14365,N_14091);
or U16781 (N_16781,N_12596,N_14271);
nand U16782 (N_16782,N_13993,N_13609);
and U16783 (N_16783,N_13069,N_14797);
nor U16784 (N_16784,N_14824,N_14977);
nand U16785 (N_16785,N_12933,N_14329);
nand U16786 (N_16786,N_12645,N_14987);
and U16787 (N_16787,N_12336,N_13946);
nor U16788 (N_16788,N_14699,N_13119);
nand U16789 (N_16789,N_14309,N_14656);
or U16790 (N_16790,N_12323,N_12132);
or U16791 (N_16791,N_12364,N_14393);
nor U16792 (N_16792,N_13310,N_12036);
nor U16793 (N_16793,N_13268,N_12027);
nor U16794 (N_16794,N_14241,N_13764);
nor U16795 (N_16795,N_12629,N_13117);
nand U16796 (N_16796,N_12257,N_13380);
or U16797 (N_16797,N_12576,N_12616);
nor U16798 (N_16798,N_14887,N_13936);
nand U16799 (N_16799,N_12923,N_14166);
and U16800 (N_16800,N_13040,N_12060);
xnor U16801 (N_16801,N_12170,N_13173);
and U16802 (N_16802,N_14328,N_14766);
nand U16803 (N_16803,N_13960,N_14410);
nand U16804 (N_16804,N_12724,N_13233);
xnor U16805 (N_16805,N_13516,N_14910);
nand U16806 (N_16806,N_14793,N_13105);
xor U16807 (N_16807,N_13629,N_13420);
and U16808 (N_16808,N_12752,N_13715);
nand U16809 (N_16809,N_12137,N_13465);
xnor U16810 (N_16810,N_13004,N_14277);
xor U16811 (N_16811,N_13456,N_14724);
and U16812 (N_16812,N_12118,N_13094);
or U16813 (N_16813,N_12525,N_13077);
and U16814 (N_16814,N_14039,N_12079);
and U16815 (N_16815,N_14718,N_13641);
or U16816 (N_16816,N_13172,N_14823);
and U16817 (N_16817,N_12002,N_14890);
or U16818 (N_16818,N_14638,N_14634);
nor U16819 (N_16819,N_12229,N_13442);
xor U16820 (N_16820,N_13276,N_14130);
nor U16821 (N_16821,N_13347,N_14181);
and U16822 (N_16822,N_12384,N_14989);
or U16823 (N_16823,N_13112,N_14926);
nor U16824 (N_16824,N_14749,N_12264);
xnor U16825 (N_16825,N_13191,N_13203);
xor U16826 (N_16826,N_12720,N_12448);
and U16827 (N_16827,N_12685,N_13964);
nand U16828 (N_16828,N_12106,N_14069);
xor U16829 (N_16829,N_14459,N_14496);
nand U16830 (N_16830,N_13149,N_14196);
and U16831 (N_16831,N_14991,N_14152);
nor U16832 (N_16832,N_12153,N_14938);
nand U16833 (N_16833,N_14327,N_12099);
nand U16834 (N_16834,N_12781,N_12138);
xor U16835 (N_16835,N_14982,N_12129);
nor U16836 (N_16836,N_12628,N_12767);
and U16837 (N_16837,N_13810,N_12384);
nor U16838 (N_16838,N_14028,N_12725);
xnor U16839 (N_16839,N_13068,N_12553);
and U16840 (N_16840,N_12431,N_14751);
xnor U16841 (N_16841,N_14989,N_14719);
or U16842 (N_16842,N_13924,N_13111);
and U16843 (N_16843,N_13498,N_14609);
or U16844 (N_16844,N_14869,N_14521);
and U16845 (N_16845,N_12699,N_14324);
nand U16846 (N_16846,N_12224,N_14361);
nor U16847 (N_16847,N_13681,N_14271);
and U16848 (N_16848,N_13749,N_13985);
nor U16849 (N_16849,N_14255,N_12892);
or U16850 (N_16850,N_12142,N_12602);
nor U16851 (N_16851,N_12478,N_14641);
and U16852 (N_16852,N_13983,N_13710);
nor U16853 (N_16853,N_12007,N_14657);
nand U16854 (N_16854,N_13837,N_12703);
nor U16855 (N_16855,N_13385,N_13114);
or U16856 (N_16856,N_14753,N_14719);
nand U16857 (N_16857,N_14352,N_13097);
nor U16858 (N_16858,N_13481,N_14284);
or U16859 (N_16859,N_12032,N_14051);
and U16860 (N_16860,N_13816,N_12140);
nor U16861 (N_16861,N_14231,N_12586);
xnor U16862 (N_16862,N_14981,N_13829);
or U16863 (N_16863,N_13075,N_13694);
xor U16864 (N_16864,N_13787,N_14286);
xor U16865 (N_16865,N_14362,N_14072);
nand U16866 (N_16866,N_14561,N_14617);
nor U16867 (N_16867,N_13289,N_13329);
nand U16868 (N_16868,N_13389,N_12523);
and U16869 (N_16869,N_12298,N_14477);
nand U16870 (N_16870,N_12998,N_12428);
xor U16871 (N_16871,N_14075,N_12946);
nand U16872 (N_16872,N_12421,N_12872);
nor U16873 (N_16873,N_14356,N_13062);
or U16874 (N_16874,N_12069,N_14558);
xor U16875 (N_16875,N_13318,N_12152);
nor U16876 (N_16876,N_13161,N_12253);
nand U16877 (N_16877,N_14654,N_12054);
and U16878 (N_16878,N_13862,N_14094);
or U16879 (N_16879,N_14391,N_12667);
nand U16880 (N_16880,N_12707,N_13655);
or U16881 (N_16881,N_14318,N_14812);
nand U16882 (N_16882,N_13486,N_14098);
nand U16883 (N_16883,N_14159,N_12440);
xnor U16884 (N_16884,N_14054,N_14475);
xor U16885 (N_16885,N_12104,N_12310);
nand U16886 (N_16886,N_12321,N_12775);
nand U16887 (N_16887,N_14456,N_12784);
xnor U16888 (N_16888,N_13266,N_12834);
nand U16889 (N_16889,N_13972,N_13631);
xnor U16890 (N_16890,N_12878,N_12809);
or U16891 (N_16891,N_14636,N_13588);
nor U16892 (N_16892,N_12814,N_12681);
and U16893 (N_16893,N_12333,N_13244);
xor U16894 (N_16894,N_13665,N_13140);
or U16895 (N_16895,N_12964,N_14734);
or U16896 (N_16896,N_13067,N_14183);
and U16897 (N_16897,N_14850,N_14658);
nor U16898 (N_16898,N_12068,N_14294);
xnor U16899 (N_16899,N_13971,N_12365);
xnor U16900 (N_16900,N_13885,N_12548);
nand U16901 (N_16901,N_14480,N_12789);
nand U16902 (N_16902,N_14911,N_14943);
xnor U16903 (N_16903,N_13614,N_12245);
nand U16904 (N_16904,N_13299,N_12258);
nor U16905 (N_16905,N_12899,N_14039);
nand U16906 (N_16906,N_12633,N_14755);
nand U16907 (N_16907,N_12729,N_14298);
nand U16908 (N_16908,N_12672,N_13180);
and U16909 (N_16909,N_12469,N_14762);
xnor U16910 (N_16910,N_13563,N_13012);
or U16911 (N_16911,N_12513,N_12792);
nor U16912 (N_16912,N_12659,N_13154);
and U16913 (N_16913,N_12770,N_12945);
nor U16914 (N_16914,N_14636,N_12417);
or U16915 (N_16915,N_13144,N_13744);
and U16916 (N_16916,N_12139,N_13202);
xor U16917 (N_16917,N_14087,N_14758);
and U16918 (N_16918,N_12630,N_12097);
or U16919 (N_16919,N_14819,N_12024);
or U16920 (N_16920,N_12214,N_14411);
nand U16921 (N_16921,N_13300,N_13749);
and U16922 (N_16922,N_14663,N_13287);
nor U16923 (N_16923,N_14306,N_14538);
and U16924 (N_16924,N_13622,N_14144);
nand U16925 (N_16925,N_14037,N_14934);
or U16926 (N_16926,N_13494,N_14992);
or U16927 (N_16927,N_12268,N_12746);
or U16928 (N_16928,N_13705,N_13535);
or U16929 (N_16929,N_12404,N_12421);
and U16930 (N_16930,N_12421,N_13390);
nor U16931 (N_16931,N_13683,N_13627);
nand U16932 (N_16932,N_13906,N_13566);
and U16933 (N_16933,N_12104,N_12750);
nor U16934 (N_16934,N_13322,N_14940);
nand U16935 (N_16935,N_12700,N_14726);
xor U16936 (N_16936,N_13213,N_14736);
xor U16937 (N_16937,N_13522,N_13269);
nor U16938 (N_16938,N_13161,N_14747);
and U16939 (N_16939,N_13615,N_12947);
or U16940 (N_16940,N_13515,N_13247);
xor U16941 (N_16941,N_13973,N_14738);
or U16942 (N_16942,N_13086,N_12246);
nand U16943 (N_16943,N_14357,N_13491);
nand U16944 (N_16944,N_14732,N_14191);
nand U16945 (N_16945,N_14147,N_14222);
and U16946 (N_16946,N_12011,N_12005);
nand U16947 (N_16947,N_13270,N_12753);
nand U16948 (N_16948,N_14464,N_14355);
nand U16949 (N_16949,N_12187,N_14127);
nand U16950 (N_16950,N_12734,N_12031);
xor U16951 (N_16951,N_14429,N_13419);
or U16952 (N_16952,N_12264,N_12623);
xor U16953 (N_16953,N_13063,N_12503);
and U16954 (N_16954,N_12127,N_14259);
nand U16955 (N_16955,N_12497,N_13340);
or U16956 (N_16956,N_12838,N_12613);
or U16957 (N_16957,N_14157,N_14821);
xnor U16958 (N_16958,N_12296,N_14536);
or U16959 (N_16959,N_12011,N_12427);
nor U16960 (N_16960,N_12121,N_14380);
nor U16961 (N_16961,N_12932,N_14879);
xor U16962 (N_16962,N_14731,N_12077);
or U16963 (N_16963,N_12705,N_14343);
nor U16964 (N_16964,N_12638,N_12135);
nor U16965 (N_16965,N_12902,N_13498);
nand U16966 (N_16966,N_14194,N_14574);
and U16967 (N_16967,N_14625,N_13343);
and U16968 (N_16968,N_13218,N_14759);
nand U16969 (N_16969,N_12132,N_12668);
nor U16970 (N_16970,N_14410,N_12122);
xnor U16971 (N_16971,N_12443,N_14659);
xnor U16972 (N_16972,N_13171,N_13308);
nor U16973 (N_16973,N_14802,N_12300);
or U16974 (N_16974,N_13697,N_14036);
xnor U16975 (N_16975,N_12125,N_13786);
nor U16976 (N_16976,N_12975,N_13187);
xor U16977 (N_16977,N_14803,N_13464);
or U16978 (N_16978,N_12753,N_12990);
xor U16979 (N_16979,N_14592,N_14327);
nor U16980 (N_16980,N_14364,N_13953);
nand U16981 (N_16981,N_14323,N_13835);
or U16982 (N_16982,N_14002,N_13202);
and U16983 (N_16983,N_14805,N_13317);
nand U16984 (N_16984,N_14024,N_12420);
nor U16985 (N_16985,N_14909,N_12213);
and U16986 (N_16986,N_12938,N_12752);
xor U16987 (N_16987,N_13679,N_13473);
nor U16988 (N_16988,N_14423,N_12117);
and U16989 (N_16989,N_14036,N_14262);
and U16990 (N_16990,N_12569,N_14121);
nor U16991 (N_16991,N_14754,N_14623);
xnor U16992 (N_16992,N_14779,N_14221);
and U16993 (N_16993,N_13560,N_12359);
xnor U16994 (N_16994,N_14418,N_12674);
xor U16995 (N_16995,N_14438,N_12721);
xor U16996 (N_16996,N_14820,N_14595);
or U16997 (N_16997,N_14469,N_14557);
nor U16998 (N_16998,N_14748,N_12811);
nor U16999 (N_16999,N_12559,N_12764);
nand U17000 (N_17000,N_14689,N_13020);
nor U17001 (N_17001,N_12839,N_14547);
or U17002 (N_17002,N_14911,N_13234);
nand U17003 (N_17003,N_14118,N_14223);
or U17004 (N_17004,N_12798,N_14463);
xor U17005 (N_17005,N_13517,N_13599);
or U17006 (N_17006,N_12119,N_13608);
nand U17007 (N_17007,N_14488,N_13685);
or U17008 (N_17008,N_14285,N_12965);
xnor U17009 (N_17009,N_13470,N_12817);
and U17010 (N_17010,N_12247,N_12803);
xor U17011 (N_17011,N_13521,N_14587);
xor U17012 (N_17012,N_14120,N_13953);
or U17013 (N_17013,N_12036,N_14143);
or U17014 (N_17014,N_12982,N_12668);
and U17015 (N_17015,N_14179,N_13110);
xnor U17016 (N_17016,N_14005,N_13678);
xor U17017 (N_17017,N_14313,N_12761);
or U17018 (N_17018,N_12614,N_14661);
or U17019 (N_17019,N_12911,N_14215);
or U17020 (N_17020,N_14537,N_14196);
nor U17021 (N_17021,N_13434,N_12535);
and U17022 (N_17022,N_14628,N_12235);
nand U17023 (N_17023,N_13213,N_14101);
or U17024 (N_17024,N_13757,N_14536);
or U17025 (N_17025,N_12817,N_12358);
nand U17026 (N_17026,N_14006,N_14943);
nand U17027 (N_17027,N_13825,N_13790);
nand U17028 (N_17028,N_12173,N_13037);
and U17029 (N_17029,N_12247,N_13626);
xnor U17030 (N_17030,N_13313,N_13010);
or U17031 (N_17031,N_12017,N_12425);
xnor U17032 (N_17032,N_13948,N_13468);
nor U17033 (N_17033,N_14964,N_13133);
xnor U17034 (N_17034,N_14468,N_12853);
and U17035 (N_17035,N_13209,N_13143);
and U17036 (N_17036,N_13370,N_14035);
xnor U17037 (N_17037,N_13164,N_12798);
or U17038 (N_17038,N_14778,N_13517);
xor U17039 (N_17039,N_13783,N_14893);
and U17040 (N_17040,N_13170,N_12554);
or U17041 (N_17041,N_12431,N_12426);
nand U17042 (N_17042,N_14953,N_12846);
nand U17043 (N_17043,N_13786,N_12960);
and U17044 (N_17044,N_12267,N_13037);
xor U17045 (N_17045,N_12398,N_14739);
nand U17046 (N_17046,N_14374,N_13624);
nor U17047 (N_17047,N_13969,N_13282);
xor U17048 (N_17048,N_12769,N_13019);
nor U17049 (N_17049,N_12440,N_12912);
nand U17050 (N_17050,N_14493,N_12924);
or U17051 (N_17051,N_13910,N_12003);
nand U17052 (N_17052,N_13818,N_13861);
xor U17053 (N_17053,N_13578,N_13139);
xor U17054 (N_17054,N_14911,N_14079);
and U17055 (N_17055,N_12586,N_12384);
xor U17056 (N_17056,N_13925,N_13881);
nor U17057 (N_17057,N_13739,N_14835);
xnor U17058 (N_17058,N_14537,N_14892);
xor U17059 (N_17059,N_14690,N_14553);
or U17060 (N_17060,N_12026,N_14245);
xor U17061 (N_17061,N_12172,N_14996);
nand U17062 (N_17062,N_12991,N_14204);
nor U17063 (N_17063,N_13820,N_12758);
nand U17064 (N_17064,N_14823,N_13477);
nand U17065 (N_17065,N_14145,N_14741);
nand U17066 (N_17066,N_14709,N_14119);
or U17067 (N_17067,N_12905,N_12286);
nand U17068 (N_17068,N_12206,N_14578);
xor U17069 (N_17069,N_13620,N_12614);
and U17070 (N_17070,N_13747,N_14269);
xnor U17071 (N_17071,N_14838,N_14975);
nand U17072 (N_17072,N_14050,N_13067);
or U17073 (N_17073,N_12977,N_12445);
and U17074 (N_17074,N_13254,N_12986);
nand U17075 (N_17075,N_12092,N_12876);
or U17076 (N_17076,N_12925,N_14375);
nand U17077 (N_17077,N_13296,N_14358);
nor U17078 (N_17078,N_12872,N_14643);
nand U17079 (N_17079,N_12325,N_13598);
or U17080 (N_17080,N_14415,N_13535);
and U17081 (N_17081,N_12975,N_14982);
nor U17082 (N_17082,N_12746,N_12387);
xnor U17083 (N_17083,N_12201,N_12551);
and U17084 (N_17084,N_12688,N_14045);
nor U17085 (N_17085,N_12743,N_12632);
nand U17086 (N_17086,N_14030,N_12789);
xor U17087 (N_17087,N_12145,N_14684);
nor U17088 (N_17088,N_12352,N_14946);
xnor U17089 (N_17089,N_13433,N_14477);
xor U17090 (N_17090,N_14208,N_12213);
nand U17091 (N_17091,N_13524,N_12065);
xor U17092 (N_17092,N_14314,N_13075);
nand U17093 (N_17093,N_14058,N_14650);
nor U17094 (N_17094,N_14163,N_12630);
nor U17095 (N_17095,N_14078,N_14431);
nand U17096 (N_17096,N_12789,N_12621);
or U17097 (N_17097,N_14171,N_14929);
and U17098 (N_17098,N_14639,N_13024);
xor U17099 (N_17099,N_13632,N_14785);
nand U17100 (N_17100,N_14686,N_14195);
nand U17101 (N_17101,N_13692,N_12344);
or U17102 (N_17102,N_14912,N_13340);
nand U17103 (N_17103,N_14713,N_14152);
nor U17104 (N_17104,N_12907,N_12248);
xor U17105 (N_17105,N_13012,N_12129);
xnor U17106 (N_17106,N_14980,N_12283);
nor U17107 (N_17107,N_14307,N_12710);
and U17108 (N_17108,N_13581,N_14405);
nand U17109 (N_17109,N_13221,N_13309);
xnor U17110 (N_17110,N_13369,N_13813);
nand U17111 (N_17111,N_12376,N_13485);
or U17112 (N_17112,N_13446,N_12241);
nor U17113 (N_17113,N_12921,N_12309);
or U17114 (N_17114,N_12776,N_14630);
nor U17115 (N_17115,N_13728,N_14488);
xnor U17116 (N_17116,N_14057,N_12770);
nor U17117 (N_17117,N_13866,N_12737);
nand U17118 (N_17118,N_14611,N_13740);
xnor U17119 (N_17119,N_12122,N_13151);
or U17120 (N_17120,N_13908,N_14396);
nor U17121 (N_17121,N_13347,N_14745);
and U17122 (N_17122,N_12954,N_12803);
xnor U17123 (N_17123,N_12804,N_14498);
and U17124 (N_17124,N_12795,N_13452);
nor U17125 (N_17125,N_12481,N_12410);
xnor U17126 (N_17126,N_12535,N_14140);
nand U17127 (N_17127,N_14042,N_13300);
nand U17128 (N_17128,N_12880,N_14288);
nand U17129 (N_17129,N_14434,N_14873);
nand U17130 (N_17130,N_12688,N_14810);
nand U17131 (N_17131,N_13955,N_14388);
and U17132 (N_17132,N_13145,N_12517);
xor U17133 (N_17133,N_14627,N_13312);
xor U17134 (N_17134,N_12997,N_12192);
nand U17135 (N_17135,N_14584,N_14651);
nand U17136 (N_17136,N_12498,N_13196);
and U17137 (N_17137,N_13804,N_14340);
xnor U17138 (N_17138,N_13801,N_13333);
and U17139 (N_17139,N_12038,N_12891);
or U17140 (N_17140,N_14973,N_12094);
nor U17141 (N_17141,N_14690,N_14026);
nor U17142 (N_17142,N_12692,N_14970);
and U17143 (N_17143,N_13424,N_13787);
nand U17144 (N_17144,N_13430,N_12777);
or U17145 (N_17145,N_13682,N_13693);
or U17146 (N_17146,N_14266,N_12230);
nand U17147 (N_17147,N_14042,N_14499);
xnor U17148 (N_17148,N_13374,N_13428);
nand U17149 (N_17149,N_13086,N_12441);
or U17150 (N_17150,N_13316,N_13846);
or U17151 (N_17151,N_12794,N_14735);
nand U17152 (N_17152,N_12692,N_14623);
nor U17153 (N_17153,N_13946,N_13789);
xnor U17154 (N_17154,N_14970,N_12873);
or U17155 (N_17155,N_12621,N_13839);
nor U17156 (N_17156,N_14637,N_14740);
xnor U17157 (N_17157,N_12020,N_13245);
xnor U17158 (N_17158,N_12078,N_13802);
and U17159 (N_17159,N_13568,N_14214);
nor U17160 (N_17160,N_13783,N_14777);
and U17161 (N_17161,N_12194,N_14490);
and U17162 (N_17162,N_13241,N_14729);
nand U17163 (N_17163,N_12079,N_12713);
nor U17164 (N_17164,N_13215,N_14298);
and U17165 (N_17165,N_14646,N_14018);
nor U17166 (N_17166,N_13464,N_12507);
and U17167 (N_17167,N_12464,N_14937);
nand U17168 (N_17168,N_13385,N_14262);
nand U17169 (N_17169,N_12486,N_12803);
nand U17170 (N_17170,N_12826,N_14170);
nand U17171 (N_17171,N_12134,N_12402);
and U17172 (N_17172,N_14922,N_14548);
or U17173 (N_17173,N_13744,N_12885);
xor U17174 (N_17174,N_13391,N_13307);
or U17175 (N_17175,N_14879,N_12825);
nor U17176 (N_17176,N_14588,N_14855);
xor U17177 (N_17177,N_13121,N_12142);
and U17178 (N_17178,N_14436,N_14471);
or U17179 (N_17179,N_14657,N_12797);
nand U17180 (N_17180,N_13176,N_12137);
or U17181 (N_17181,N_14928,N_13841);
xor U17182 (N_17182,N_12026,N_12587);
nor U17183 (N_17183,N_12797,N_12210);
nor U17184 (N_17184,N_12834,N_14500);
nor U17185 (N_17185,N_14795,N_12435);
nor U17186 (N_17186,N_14528,N_14722);
nor U17187 (N_17187,N_13377,N_13782);
nor U17188 (N_17188,N_13203,N_12396);
and U17189 (N_17189,N_14048,N_12563);
nand U17190 (N_17190,N_13825,N_13153);
nor U17191 (N_17191,N_14844,N_12276);
nand U17192 (N_17192,N_13291,N_14800);
or U17193 (N_17193,N_14797,N_12884);
or U17194 (N_17194,N_12287,N_13463);
xnor U17195 (N_17195,N_14298,N_13176);
and U17196 (N_17196,N_13161,N_12320);
nor U17197 (N_17197,N_14347,N_12822);
or U17198 (N_17198,N_12964,N_12886);
nor U17199 (N_17199,N_13580,N_12660);
nor U17200 (N_17200,N_13410,N_13396);
and U17201 (N_17201,N_12854,N_14261);
nand U17202 (N_17202,N_13756,N_14827);
nor U17203 (N_17203,N_13923,N_12400);
and U17204 (N_17204,N_14343,N_13768);
or U17205 (N_17205,N_13801,N_13169);
xnor U17206 (N_17206,N_13955,N_12082);
nand U17207 (N_17207,N_14565,N_12048);
nand U17208 (N_17208,N_12201,N_12225);
nand U17209 (N_17209,N_13709,N_12378);
nand U17210 (N_17210,N_12688,N_12906);
and U17211 (N_17211,N_13582,N_14139);
nor U17212 (N_17212,N_12752,N_12056);
nand U17213 (N_17213,N_14121,N_13228);
nand U17214 (N_17214,N_13507,N_14255);
xnor U17215 (N_17215,N_14347,N_13006);
and U17216 (N_17216,N_14573,N_14470);
nor U17217 (N_17217,N_13361,N_13415);
nand U17218 (N_17218,N_12954,N_12802);
and U17219 (N_17219,N_12683,N_13812);
or U17220 (N_17220,N_12448,N_14257);
and U17221 (N_17221,N_13408,N_14812);
xor U17222 (N_17222,N_13067,N_14990);
or U17223 (N_17223,N_12119,N_12425);
xnor U17224 (N_17224,N_14061,N_14455);
and U17225 (N_17225,N_12076,N_14067);
xor U17226 (N_17226,N_13749,N_12543);
xor U17227 (N_17227,N_14329,N_14460);
and U17228 (N_17228,N_14057,N_14749);
nand U17229 (N_17229,N_12935,N_13148);
xor U17230 (N_17230,N_14741,N_13599);
or U17231 (N_17231,N_14443,N_12556);
xnor U17232 (N_17232,N_14230,N_13275);
nand U17233 (N_17233,N_12511,N_12439);
xnor U17234 (N_17234,N_14625,N_12366);
xor U17235 (N_17235,N_13562,N_13590);
nand U17236 (N_17236,N_13920,N_12762);
and U17237 (N_17237,N_13312,N_12595);
nor U17238 (N_17238,N_14414,N_12612);
or U17239 (N_17239,N_14133,N_13006);
nand U17240 (N_17240,N_14227,N_12154);
and U17241 (N_17241,N_12325,N_14821);
nand U17242 (N_17242,N_13567,N_14094);
nand U17243 (N_17243,N_12486,N_13781);
and U17244 (N_17244,N_12773,N_12116);
nand U17245 (N_17245,N_12945,N_13599);
xor U17246 (N_17246,N_13442,N_14711);
nor U17247 (N_17247,N_13764,N_12813);
nor U17248 (N_17248,N_14986,N_12410);
nand U17249 (N_17249,N_13972,N_13743);
xor U17250 (N_17250,N_12704,N_14263);
xnor U17251 (N_17251,N_12799,N_14960);
and U17252 (N_17252,N_12075,N_13033);
nand U17253 (N_17253,N_14702,N_14786);
xnor U17254 (N_17254,N_14626,N_12104);
nor U17255 (N_17255,N_14059,N_12349);
and U17256 (N_17256,N_12249,N_12987);
xor U17257 (N_17257,N_12467,N_12357);
nand U17258 (N_17258,N_12604,N_12095);
and U17259 (N_17259,N_14923,N_12970);
and U17260 (N_17260,N_12626,N_13367);
nand U17261 (N_17261,N_13241,N_14816);
xor U17262 (N_17262,N_13276,N_14900);
xor U17263 (N_17263,N_14399,N_13860);
nor U17264 (N_17264,N_13686,N_12010);
nor U17265 (N_17265,N_14285,N_13241);
and U17266 (N_17266,N_12554,N_12791);
nand U17267 (N_17267,N_12133,N_13689);
nor U17268 (N_17268,N_14737,N_12692);
nor U17269 (N_17269,N_13842,N_12942);
or U17270 (N_17270,N_12884,N_12281);
or U17271 (N_17271,N_13159,N_14085);
and U17272 (N_17272,N_13929,N_13352);
and U17273 (N_17273,N_12765,N_12437);
nor U17274 (N_17274,N_14070,N_13882);
and U17275 (N_17275,N_12385,N_13013);
and U17276 (N_17276,N_14134,N_12637);
xnor U17277 (N_17277,N_14862,N_14548);
xor U17278 (N_17278,N_13217,N_13538);
and U17279 (N_17279,N_14233,N_12407);
nand U17280 (N_17280,N_13398,N_13703);
nor U17281 (N_17281,N_13877,N_14869);
or U17282 (N_17282,N_13960,N_14207);
and U17283 (N_17283,N_13792,N_13943);
or U17284 (N_17284,N_12455,N_12194);
nor U17285 (N_17285,N_12941,N_13775);
or U17286 (N_17286,N_13708,N_13709);
nand U17287 (N_17287,N_12286,N_12813);
nor U17288 (N_17288,N_13664,N_12360);
nor U17289 (N_17289,N_12229,N_13952);
and U17290 (N_17290,N_12787,N_14364);
nor U17291 (N_17291,N_14365,N_12692);
or U17292 (N_17292,N_13869,N_13936);
and U17293 (N_17293,N_12550,N_12445);
and U17294 (N_17294,N_14610,N_12755);
and U17295 (N_17295,N_14852,N_12963);
or U17296 (N_17296,N_13930,N_13149);
xor U17297 (N_17297,N_12575,N_13886);
and U17298 (N_17298,N_12713,N_12751);
xnor U17299 (N_17299,N_13681,N_14793);
nand U17300 (N_17300,N_13441,N_12460);
nand U17301 (N_17301,N_13639,N_14315);
and U17302 (N_17302,N_13491,N_12815);
nand U17303 (N_17303,N_14913,N_14426);
or U17304 (N_17304,N_12031,N_14055);
xnor U17305 (N_17305,N_13502,N_12695);
xnor U17306 (N_17306,N_14546,N_13662);
nand U17307 (N_17307,N_14020,N_14716);
xor U17308 (N_17308,N_12228,N_14539);
xor U17309 (N_17309,N_14569,N_13061);
nand U17310 (N_17310,N_13091,N_14217);
xnor U17311 (N_17311,N_12308,N_14175);
nand U17312 (N_17312,N_14084,N_14417);
and U17313 (N_17313,N_13311,N_12670);
nor U17314 (N_17314,N_13088,N_12433);
or U17315 (N_17315,N_13376,N_13463);
or U17316 (N_17316,N_14168,N_13389);
or U17317 (N_17317,N_13069,N_12898);
or U17318 (N_17318,N_13535,N_12987);
and U17319 (N_17319,N_12357,N_14399);
and U17320 (N_17320,N_14405,N_14704);
and U17321 (N_17321,N_14254,N_13318);
nand U17322 (N_17322,N_12389,N_12743);
or U17323 (N_17323,N_14257,N_13995);
xnor U17324 (N_17324,N_14769,N_12054);
and U17325 (N_17325,N_14216,N_13347);
or U17326 (N_17326,N_13958,N_14765);
xor U17327 (N_17327,N_12269,N_12649);
xor U17328 (N_17328,N_12995,N_13492);
nand U17329 (N_17329,N_12692,N_14480);
or U17330 (N_17330,N_12972,N_14479);
xnor U17331 (N_17331,N_13016,N_13658);
nand U17332 (N_17332,N_12596,N_13623);
and U17333 (N_17333,N_14816,N_14662);
xor U17334 (N_17334,N_14772,N_14864);
xor U17335 (N_17335,N_14110,N_14919);
and U17336 (N_17336,N_12873,N_13861);
and U17337 (N_17337,N_14348,N_14614);
xor U17338 (N_17338,N_13993,N_14290);
and U17339 (N_17339,N_13294,N_12060);
xnor U17340 (N_17340,N_13125,N_13193);
nand U17341 (N_17341,N_13244,N_13401);
xnor U17342 (N_17342,N_12929,N_14434);
nor U17343 (N_17343,N_14844,N_14026);
nand U17344 (N_17344,N_14456,N_13140);
xor U17345 (N_17345,N_14099,N_14327);
nor U17346 (N_17346,N_13780,N_13969);
nor U17347 (N_17347,N_13680,N_14036);
and U17348 (N_17348,N_12268,N_12686);
nor U17349 (N_17349,N_12941,N_14519);
nand U17350 (N_17350,N_13205,N_14882);
nand U17351 (N_17351,N_13492,N_14773);
xor U17352 (N_17352,N_13559,N_12581);
xnor U17353 (N_17353,N_13091,N_12284);
nor U17354 (N_17354,N_13112,N_12769);
nand U17355 (N_17355,N_14404,N_14640);
and U17356 (N_17356,N_14937,N_12695);
or U17357 (N_17357,N_13115,N_13772);
xor U17358 (N_17358,N_12725,N_14914);
or U17359 (N_17359,N_14410,N_14096);
nand U17360 (N_17360,N_12116,N_14795);
or U17361 (N_17361,N_13822,N_13262);
or U17362 (N_17362,N_13466,N_14469);
xnor U17363 (N_17363,N_14676,N_12499);
xnor U17364 (N_17364,N_14570,N_12307);
nand U17365 (N_17365,N_14031,N_14643);
or U17366 (N_17366,N_12153,N_13326);
and U17367 (N_17367,N_13921,N_14482);
or U17368 (N_17368,N_14249,N_13383);
or U17369 (N_17369,N_14536,N_12812);
nand U17370 (N_17370,N_13681,N_13618);
nand U17371 (N_17371,N_14409,N_12858);
nand U17372 (N_17372,N_12362,N_13771);
nand U17373 (N_17373,N_12962,N_12792);
nand U17374 (N_17374,N_12776,N_13098);
or U17375 (N_17375,N_12642,N_13541);
nand U17376 (N_17376,N_14998,N_12163);
nand U17377 (N_17377,N_13991,N_12864);
nand U17378 (N_17378,N_13317,N_14124);
and U17379 (N_17379,N_12931,N_13543);
nor U17380 (N_17380,N_14161,N_13382);
nand U17381 (N_17381,N_13489,N_13525);
xnor U17382 (N_17382,N_13937,N_13231);
nand U17383 (N_17383,N_13315,N_12465);
xnor U17384 (N_17384,N_13316,N_14207);
or U17385 (N_17385,N_12187,N_12442);
nand U17386 (N_17386,N_13096,N_13056);
and U17387 (N_17387,N_14178,N_14956);
nor U17388 (N_17388,N_14214,N_12017);
and U17389 (N_17389,N_13575,N_14333);
or U17390 (N_17390,N_14127,N_13403);
xnor U17391 (N_17391,N_12304,N_12970);
nor U17392 (N_17392,N_12480,N_12804);
xnor U17393 (N_17393,N_14474,N_13815);
nand U17394 (N_17394,N_14415,N_14200);
and U17395 (N_17395,N_13967,N_14277);
and U17396 (N_17396,N_13371,N_12501);
and U17397 (N_17397,N_12477,N_13811);
nor U17398 (N_17398,N_12888,N_12304);
or U17399 (N_17399,N_13936,N_13046);
and U17400 (N_17400,N_12213,N_12062);
xor U17401 (N_17401,N_14661,N_13692);
and U17402 (N_17402,N_14742,N_13932);
or U17403 (N_17403,N_12531,N_12186);
xnor U17404 (N_17404,N_12119,N_13414);
and U17405 (N_17405,N_13862,N_14000);
and U17406 (N_17406,N_14606,N_13477);
xnor U17407 (N_17407,N_14377,N_12539);
nor U17408 (N_17408,N_14216,N_13092);
nand U17409 (N_17409,N_14890,N_14962);
nor U17410 (N_17410,N_14426,N_13691);
nor U17411 (N_17411,N_14994,N_13163);
or U17412 (N_17412,N_14551,N_12605);
nor U17413 (N_17413,N_13918,N_14555);
nand U17414 (N_17414,N_13682,N_14237);
nor U17415 (N_17415,N_12484,N_12630);
nor U17416 (N_17416,N_14229,N_12369);
and U17417 (N_17417,N_13297,N_12948);
nor U17418 (N_17418,N_14258,N_12585);
nand U17419 (N_17419,N_12523,N_14543);
nand U17420 (N_17420,N_14691,N_13582);
nand U17421 (N_17421,N_12014,N_14632);
xnor U17422 (N_17422,N_13276,N_14868);
nand U17423 (N_17423,N_12224,N_14178);
or U17424 (N_17424,N_14070,N_13656);
or U17425 (N_17425,N_12418,N_12679);
nand U17426 (N_17426,N_14793,N_12725);
and U17427 (N_17427,N_13219,N_12274);
or U17428 (N_17428,N_14318,N_13951);
and U17429 (N_17429,N_14084,N_14530);
nor U17430 (N_17430,N_12221,N_14000);
nand U17431 (N_17431,N_12770,N_12312);
xnor U17432 (N_17432,N_14678,N_12790);
and U17433 (N_17433,N_13920,N_14277);
nor U17434 (N_17434,N_12676,N_12775);
and U17435 (N_17435,N_14289,N_13771);
and U17436 (N_17436,N_14063,N_12963);
nor U17437 (N_17437,N_12370,N_12287);
or U17438 (N_17438,N_14207,N_12631);
xor U17439 (N_17439,N_13669,N_12484);
nand U17440 (N_17440,N_12297,N_14012);
or U17441 (N_17441,N_14968,N_14801);
xnor U17442 (N_17442,N_12417,N_14789);
and U17443 (N_17443,N_13265,N_12358);
and U17444 (N_17444,N_13536,N_12357);
nand U17445 (N_17445,N_12720,N_12806);
or U17446 (N_17446,N_12906,N_12162);
and U17447 (N_17447,N_14371,N_14079);
nor U17448 (N_17448,N_13731,N_14583);
and U17449 (N_17449,N_12634,N_13291);
nand U17450 (N_17450,N_13647,N_13009);
nand U17451 (N_17451,N_13602,N_13204);
nand U17452 (N_17452,N_13417,N_13468);
and U17453 (N_17453,N_12913,N_14486);
nor U17454 (N_17454,N_12207,N_12592);
xnor U17455 (N_17455,N_12051,N_13842);
or U17456 (N_17456,N_14925,N_14087);
nand U17457 (N_17457,N_14706,N_12513);
nand U17458 (N_17458,N_12840,N_12128);
or U17459 (N_17459,N_12853,N_14032);
or U17460 (N_17460,N_14446,N_13710);
nand U17461 (N_17461,N_12173,N_12671);
nand U17462 (N_17462,N_14957,N_12590);
xor U17463 (N_17463,N_12379,N_14624);
or U17464 (N_17464,N_14365,N_14912);
or U17465 (N_17465,N_13173,N_12506);
nor U17466 (N_17466,N_14201,N_13407);
nand U17467 (N_17467,N_12209,N_14287);
or U17468 (N_17468,N_13241,N_13502);
nor U17469 (N_17469,N_14542,N_12956);
nand U17470 (N_17470,N_13067,N_12262);
nor U17471 (N_17471,N_12702,N_14477);
nand U17472 (N_17472,N_14341,N_13331);
and U17473 (N_17473,N_14700,N_13165);
nand U17474 (N_17474,N_12086,N_13903);
xor U17475 (N_17475,N_12890,N_12807);
xor U17476 (N_17476,N_12198,N_13307);
xnor U17477 (N_17477,N_14560,N_14079);
and U17478 (N_17478,N_12778,N_12738);
xnor U17479 (N_17479,N_12792,N_13980);
and U17480 (N_17480,N_13672,N_13994);
nor U17481 (N_17481,N_13362,N_12444);
nor U17482 (N_17482,N_12377,N_13830);
and U17483 (N_17483,N_14663,N_13904);
and U17484 (N_17484,N_14837,N_12124);
nor U17485 (N_17485,N_13604,N_12817);
or U17486 (N_17486,N_12370,N_13308);
or U17487 (N_17487,N_13620,N_14480);
or U17488 (N_17488,N_12901,N_13464);
and U17489 (N_17489,N_14880,N_14695);
and U17490 (N_17490,N_13271,N_13192);
xnor U17491 (N_17491,N_14873,N_12298);
or U17492 (N_17492,N_12073,N_13360);
nand U17493 (N_17493,N_12159,N_12990);
or U17494 (N_17494,N_13319,N_14847);
xor U17495 (N_17495,N_12617,N_14101);
and U17496 (N_17496,N_14478,N_12927);
or U17497 (N_17497,N_14768,N_14561);
xor U17498 (N_17498,N_13258,N_13673);
and U17499 (N_17499,N_13917,N_13429);
and U17500 (N_17500,N_13373,N_14814);
or U17501 (N_17501,N_13778,N_12201);
and U17502 (N_17502,N_12717,N_13417);
xnor U17503 (N_17503,N_12938,N_14267);
xor U17504 (N_17504,N_12251,N_13413);
xor U17505 (N_17505,N_13975,N_12382);
xor U17506 (N_17506,N_14672,N_13882);
or U17507 (N_17507,N_14534,N_13310);
or U17508 (N_17508,N_12165,N_13589);
or U17509 (N_17509,N_13107,N_13767);
nand U17510 (N_17510,N_14447,N_13194);
and U17511 (N_17511,N_14406,N_13626);
and U17512 (N_17512,N_12020,N_12873);
nor U17513 (N_17513,N_12021,N_14999);
xor U17514 (N_17514,N_13582,N_12686);
nor U17515 (N_17515,N_13906,N_13679);
nor U17516 (N_17516,N_14931,N_14040);
nor U17517 (N_17517,N_12119,N_12139);
nand U17518 (N_17518,N_13871,N_12824);
nor U17519 (N_17519,N_13479,N_14827);
or U17520 (N_17520,N_12380,N_14330);
nor U17521 (N_17521,N_14063,N_12010);
xor U17522 (N_17522,N_12996,N_12484);
and U17523 (N_17523,N_12119,N_12123);
or U17524 (N_17524,N_14313,N_13099);
or U17525 (N_17525,N_12034,N_12510);
and U17526 (N_17526,N_14910,N_12984);
or U17527 (N_17527,N_14164,N_13253);
or U17528 (N_17528,N_14307,N_13915);
or U17529 (N_17529,N_14262,N_12718);
nor U17530 (N_17530,N_14365,N_12600);
nand U17531 (N_17531,N_14216,N_14668);
xnor U17532 (N_17532,N_14129,N_12522);
or U17533 (N_17533,N_12067,N_12484);
xor U17534 (N_17534,N_12093,N_13224);
nand U17535 (N_17535,N_13864,N_14754);
or U17536 (N_17536,N_12427,N_13415);
xnor U17537 (N_17537,N_12495,N_13417);
xnor U17538 (N_17538,N_13609,N_12588);
nor U17539 (N_17539,N_12115,N_12068);
nor U17540 (N_17540,N_13599,N_12936);
nand U17541 (N_17541,N_13558,N_14070);
and U17542 (N_17542,N_12320,N_12532);
and U17543 (N_17543,N_14728,N_14665);
xnor U17544 (N_17544,N_13146,N_13451);
or U17545 (N_17545,N_12159,N_14148);
or U17546 (N_17546,N_13044,N_13260);
nand U17547 (N_17547,N_12602,N_12979);
xnor U17548 (N_17548,N_12558,N_12165);
nand U17549 (N_17549,N_14765,N_14053);
and U17550 (N_17550,N_13355,N_13718);
nand U17551 (N_17551,N_12067,N_14977);
and U17552 (N_17552,N_12714,N_12151);
and U17553 (N_17553,N_12850,N_14659);
or U17554 (N_17554,N_14345,N_12647);
xnor U17555 (N_17555,N_14961,N_13409);
nand U17556 (N_17556,N_14771,N_12587);
xnor U17557 (N_17557,N_13253,N_14450);
and U17558 (N_17558,N_13998,N_14836);
nor U17559 (N_17559,N_14771,N_12455);
or U17560 (N_17560,N_12379,N_14331);
nand U17561 (N_17561,N_13530,N_13013);
and U17562 (N_17562,N_13497,N_13213);
xor U17563 (N_17563,N_14671,N_14660);
xnor U17564 (N_17564,N_13259,N_13117);
and U17565 (N_17565,N_13769,N_14354);
nor U17566 (N_17566,N_13475,N_13238);
nor U17567 (N_17567,N_12471,N_13792);
nand U17568 (N_17568,N_12275,N_14120);
and U17569 (N_17569,N_14858,N_13236);
nor U17570 (N_17570,N_12966,N_14942);
nand U17571 (N_17571,N_12494,N_14634);
or U17572 (N_17572,N_14207,N_13822);
nor U17573 (N_17573,N_13303,N_14509);
xor U17574 (N_17574,N_12816,N_14772);
nor U17575 (N_17575,N_14414,N_14246);
and U17576 (N_17576,N_14895,N_13233);
or U17577 (N_17577,N_13105,N_14166);
and U17578 (N_17578,N_14373,N_14945);
or U17579 (N_17579,N_13101,N_14353);
or U17580 (N_17580,N_12389,N_14350);
or U17581 (N_17581,N_14940,N_13720);
and U17582 (N_17582,N_12960,N_12031);
nand U17583 (N_17583,N_14467,N_13892);
nor U17584 (N_17584,N_12527,N_14462);
nor U17585 (N_17585,N_13025,N_13843);
nor U17586 (N_17586,N_14617,N_13862);
xor U17587 (N_17587,N_13288,N_12189);
and U17588 (N_17588,N_14441,N_14049);
xor U17589 (N_17589,N_14015,N_12324);
nor U17590 (N_17590,N_14480,N_14125);
xnor U17591 (N_17591,N_12941,N_13659);
nor U17592 (N_17592,N_14482,N_14840);
and U17593 (N_17593,N_12934,N_12002);
nor U17594 (N_17594,N_14934,N_12409);
or U17595 (N_17595,N_14494,N_14317);
nor U17596 (N_17596,N_13562,N_14395);
or U17597 (N_17597,N_13686,N_12501);
and U17598 (N_17598,N_14884,N_14312);
nand U17599 (N_17599,N_12975,N_12300);
nor U17600 (N_17600,N_13986,N_13876);
and U17601 (N_17601,N_12256,N_14412);
xor U17602 (N_17602,N_14108,N_12211);
nor U17603 (N_17603,N_12277,N_13696);
xor U17604 (N_17604,N_12129,N_14426);
nor U17605 (N_17605,N_13338,N_12487);
xnor U17606 (N_17606,N_12067,N_13753);
or U17607 (N_17607,N_12795,N_12235);
xnor U17608 (N_17608,N_14246,N_13799);
nand U17609 (N_17609,N_13798,N_14574);
nor U17610 (N_17610,N_13306,N_14345);
xor U17611 (N_17611,N_12149,N_13145);
nand U17612 (N_17612,N_12307,N_14188);
nor U17613 (N_17613,N_12734,N_13932);
nand U17614 (N_17614,N_14360,N_14758);
xnor U17615 (N_17615,N_14484,N_14118);
or U17616 (N_17616,N_14972,N_13492);
or U17617 (N_17617,N_12917,N_13510);
and U17618 (N_17618,N_13597,N_13955);
xor U17619 (N_17619,N_14331,N_14370);
and U17620 (N_17620,N_14858,N_14054);
nor U17621 (N_17621,N_13214,N_13275);
nor U17622 (N_17622,N_13404,N_12098);
xnor U17623 (N_17623,N_12016,N_12533);
xor U17624 (N_17624,N_14151,N_12128);
and U17625 (N_17625,N_13069,N_14614);
or U17626 (N_17626,N_13976,N_13098);
nor U17627 (N_17627,N_13592,N_14981);
nor U17628 (N_17628,N_12799,N_12316);
and U17629 (N_17629,N_14081,N_13876);
and U17630 (N_17630,N_14831,N_13592);
nand U17631 (N_17631,N_13530,N_13812);
and U17632 (N_17632,N_13067,N_12467);
and U17633 (N_17633,N_12479,N_12712);
xor U17634 (N_17634,N_12855,N_13502);
nand U17635 (N_17635,N_12468,N_14119);
or U17636 (N_17636,N_14159,N_13939);
nand U17637 (N_17637,N_14013,N_14409);
or U17638 (N_17638,N_13333,N_13267);
nand U17639 (N_17639,N_13598,N_12406);
xnor U17640 (N_17640,N_14356,N_14271);
xnor U17641 (N_17641,N_13433,N_14884);
and U17642 (N_17642,N_13671,N_13961);
or U17643 (N_17643,N_13460,N_12212);
nor U17644 (N_17644,N_12282,N_12713);
xnor U17645 (N_17645,N_14235,N_13843);
or U17646 (N_17646,N_12991,N_14756);
or U17647 (N_17647,N_12949,N_13698);
nor U17648 (N_17648,N_13905,N_13756);
nor U17649 (N_17649,N_13941,N_12161);
xor U17650 (N_17650,N_14817,N_13875);
nor U17651 (N_17651,N_14731,N_12253);
xor U17652 (N_17652,N_13149,N_13756);
nor U17653 (N_17653,N_14980,N_14030);
and U17654 (N_17654,N_13892,N_12299);
nand U17655 (N_17655,N_13494,N_13594);
xor U17656 (N_17656,N_12964,N_13823);
and U17657 (N_17657,N_12309,N_12289);
nand U17658 (N_17658,N_12952,N_12194);
xor U17659 (N_17659,N_13147,N_12751);
nand U17660 (N_17660,N_13340,N_14823);
nor U17661 (N_17661,N_12121,N_13819);
xnor U17662 (N_17662,N_14645,N_13559);
xnor U17663 (N_17663,N_12274,N_14911);
and U17664 (N_17664,N_13679,N_14950);
nand U17665 (N_17665,N_13390,N_13542);
nand U17666 (N_17666,N_13760,N_12191);
and U17667 (N_17667,N_14276,N_14589);
nand U17668 (N_17668,N_13818,N_14294);
nand U17669 (N_17669,N_13978,N_14914);
or U17670 (N_17670,N_13254,N_12209);
or U17671 (N_17671,N_14044,N_13227);
xnor U17672 (N_17672,N_12163,N_13589);
xnor U17673 (N_17673,N_13978,N_12565);
nor U17674 (N_17674,N_13458,N_13739);
and U17675 (N_17675,N_13182,N_13118);
nand U17676 (N_17676,N_14738,N_13134);
and U17677 (N_17677,N_14319,N_12797);
nor U17678 (N_17678,N_13829,N_13451);
nor U17679 (N_17679,N_14207,N_12983);
and U17680 (N_17680,N_14557,N_14452);
xor U17681 (N_17681,N_14887,N_12660);
xnor U17682 (N_17682,N_14226,N_13620);
nor U17683 (N_17683,N_13217,N_12511);
nor U17684 (N_17684,N_12590,N_13558);
and U17685 (N_17685,N_13172,N_13853);
nand U17686 (N_17686,N_13134,N_12007);
nor U17687 (N_17687,N_14265,N_12403);
nor U17688 (N_17688,N_13035,N_14889);
or U17689 (N_17689,N_13926,N_14836);
and U17690 (N_17690,N_14316,N_13770);
nand U17691 (N_17691,N_14715,N_13140);
xor U17692 (N_17692,N_14047,N_14361);
nand U17693 (N_17693,N_13136,N_12614);
nand U17694 (N_17694,N_12937,N_14487);
or U17695 (N_17695,N_13812,N_13228);
nand U17696 (N_17696,N_13615,N_12236);
nand U17697 (N_17697,N_12187,N_14706);
and U17698 (N_17698,N_13203,N_12643);
nor U17699 (N_17699,N_14091,N_14546);
nand U17700 (N_17700,N_14686,N_12581);
or U17701 (N_17701,N_14234,N_14112);
nand U17702 (N_17702,N_14481,N_12747);
nand U17703 (N_17703,N_14792,N_13135);
and U17704 (N_17704,N_13562,N_12311);
nor U17705 (N_17705,N_13991,N_13152);
and U17706 (N_17706,N_13934,N_13212);
nor U17707 (N_17707,N_12009,N_14569);
and U17708 (N_17708,N_13309,N_14888);
xor U17709 (N_17709,N_14112,N_13308);
xor U17710 (N_17710,N_13266,N_13663);
and U17711 (N_17711,N_12271,N_12312);
or U17712 (N_17712,N_12874,N_12494);
and U17713 (N_17713,N_12662,N_12000);
xnor U17714 (N_17714,N_13140,N_12214);
and U17715 (N_17715,N_14862,N_13108);
and U17716 (N_17716,N_14419,N_14544);
or U17717 (N_17717,N_12071,N_12708);
xnor U17718 (N_17718,N_13941,N_13950);
nor U17719 (N_17719,N_12927,N_14633);
xor U17720 (N_17720,N_12299,N_12882);
xor U17721 (N_17721,N_13317,N_14266);
nand U17722 (N_17722,N_12918,N_12504);
nor U17723 (N_17723,N_14601,N_12501);
or U17724 (N_17724,N_13487,N_13179);
nor U17725 (N_17725,N_12312,N_14589);
xor U17726 (N_17726,N_14821,N_14601);
xnor U17727 (N_17727,N_12551,N_14334);
nand U17728 (N_17728,N_14429,N_14764);
nor U17729 (N_17729,N_14410,N_12990);
nor U17730 (N_17730,N_13704,N_14623);
nor U17731 (N_17731,N_14193,N_13894);
and U17732 (N_17732,N_12442,N_12386);
nand U17733 (N_17733,N_12955,N_14085);
xor U17734 (N_17734,N_13261,N_12228);
and U17735 (N_17735,N_14631,N_13358);
and U17736 (N_17736,N_14906,N_13318);
nand U17737 (N_17737,N_13409,N_13859);
nand U17738 (N_17738,N_12461,N_12964);
xnor U17739 (N_17739,N_12969,N_13343);
nor U17740 (N_17740,N_13446,N_14739);
and U17741 (N_17741,N_14052,N_13759);
xnor U17742 (N_17742,N_14323,N_12527);
or U17743 (N_17743,N_12222,N_14957);
xor U17744 (N_17744,N_14403,N_14673);
nor U17745 (N_17745,N_14880,N_13949);
and U17746 (N_17746,N_12262,N_13483);
nor U17747 (N_17747,N_14879,N_12359);
nand U17748 (N_17748,N_14740,N_13832);
and U17749 (N_17749,N_13179,N_13539);
and U17750 (N_17750,N_12963,N_14323);
nand U17751 (N_17751,N_13847,N_12177);
xnor U17752 (N_17752,N_12912,N_13139);
nand U17753 (N_17753,N_13981,N_13067);
or U17754 (N_17754,N_12525,N_13133);
and U17755 (N_17755,N_14040,N_12852);
nor U17756 (N_17756,N_12638,N_14479);
nand U17757 (N_17757,N_13365,N_13389);
nor U17758 (N_17758,N_14521,N_13351);
nor U17759 (N_17759,N_13211,N_13514);
nor U17760 (N_17760,N_14406,N_12795);
and U17761 (N_17761,N_12794,N_14901);
and U17762 (N_17762,N_14630,N_12317);
nor U17763 (N_17763,N_12497,N_12154);
nand U17764 (N_17764,N_12446,N_12185);
and U17765 (N_17765,N_13497,N_13721);
or U17766 (N_17766,N_12895,N_13086);
xnor U17767 (N_17767,N_12363,N_12271);
xnor U17768 (N_17768,N_13305,N_14827);
or U17769 (N_17769,N_13178,N_14220);
nand U17770 (N_17770,N_13610,N_12671);
nand U17771 (N_17771,N_13108,N_13573);
and U17772 (N_17772,N_14896,N_14536);
nand U17773 (N_17773,N_12886,N_14642);
xor U17774 (N_17774,N_14782,N_13343);
and U17775 (N_17775,N_14473,N_12481);
xnor U17776 (N_17776,N_14422,N_14781);
nand U17777 (N_17777,N_12117,N_13361);
nand U17778 (N_17778,N_13856,N_14352);
and U17779 (N_17779,N_13527,N_12920);
or U17780 (N_17780,N_14387,N_12882);
and U17781 (N_17781,N_14723,N_13123);
and U17782 (N_17782,N_13699,N_14783);
or U17783 (N_17783,N_12900,N_13400);
xor U17784 (N_17784,N_12347,N_13273);
or U17785 (N_17785,N_13308,N_12748);
or U17786 (N_17786,N_14471,N_14232);
or U17787 (N_17787,N_12696,N_12865);
nor U17788 (N_17788,N_14319,N_14880);
and U17789 (N_17789,N_13507,N_12388);
or U17790 (N_17790,N_12237,N_12643);
or U17791 (N_17791,N_12222,N_12289);
nand U17792 (N_17792,N_12314,N_14964);
xor U17793 (N_17793,N_13121,N_13917);
and U17794 (N_17794,N_13916,N_13922);
xor U17795 (N_17795,N_14322,N_14740);
nor U17796 (N_17796,N_12805,N_12225);
xnor U17797 (N_17797,N_14259,N_12811);
nand U17798 (N_17798,N_14285,N_13650);
nand U17799 (N_17799,N_14075,N_12704);
or U17800 (N_17800,N_12511,N_12219);
nor U17801 (N_17801,N_13592,N_14520);
nor U17802 (N_17802,N_13008,N_14300);
or U17803 (N_17803,N_14704,N_13857);
nor U17804 (N_17804,N_14311,N_14787);
xor U17805 (N_17805,N_13675,N_14917);
xor U17806 (N_17806,N_14562,N_14508);
xnor U17807 (N_17807,N_12398,N_12692);
or U17808 (N_17808,N_12961,N_13907);
and U17809 (N_17809,N_12544,N_14337);
xnor U17810 (N_17810,N_13301,N_13534);
nor U17811 (N_17811,N_14938,N_13878);
nor U17812 (N_17812,N_12880,N_12825);
or U17813 (N_17813,N_13554,N_13925);
or U17814 (N_17814,N_12832,N_14226);
xor U17815 (N_17815,N_14336,N_13732);
xor U17816 (N_17816,N_14152,N_12871);
xnor U17817 (N_17817,N_13767,N_14778);
and U17818 (N_17818,N_12384,N_14860);
and U17819 (N_17819,N_14881,N_14343);
and U17820 (N_17820,N_14594,N_13757);
or U17821 (N_17821,N_14440,N_12603);
or U17822 (N_17822,N_12713,N_12805);
and U17823 (N_17823,N_13074,N_13139);
nor U17824 (N_17824,N_13747,N_14621);
or U17825 (N_17825,N_14699,N_12316);
or U17826 (N_17826,N_13023,N_12123);
nor U17827 (N_17827,N_14568,N_12935);
nor U17828 (N_17828,N_12864,N_12514);
nand U17829 (N_17829,N_12070,N_14950);
or U17830 (N_17830,N_12329,N_12931);
or U17831 (N_17831,N_14432,N_14661);
nor U17832 (N_17832,N_12266,N_13429);
or U17833 (N_17833,N_13380,N_13805);
nand U17834 (N_17834,N_14308,N_12611);
and U17835 (N_17835,N_13120,N_13204);
xor U17836 (N_17836,N_12752,N_14836);
or U17837 (N_17837,N_13864,N_12946);
xor U17838 (N_17838,N_13880,N_12133);
and U17839 (N_17839,N_14097,N_13606);
and U17840 (N_17840,N_13458,N_14635);
nand U17841 (N_17841,N_14016,N_12313);
nor U17842 (N_17842,N_14631,N_12873);
nand U17843 (N_17843,N_12787,N_13512);
nand U17844 (N_17844,N_13863,N_14324);
nor U17845 (N_17845,N_12479,N_14864);
and U17846 (N_17846,N_12689,N_13054);
xor U17847 (N_17847,N_12888,N_14158);
xor U17848 (N_17848,N_12038,N_12607);
xnor U17849 (N_17849,N_13745,N_14237);
nor U17850 (N_17850,N_12257,N_13499);
nor U17851 (N_17851,N_14752,N_12961);
xor U17852 (N_17852,N_13403,N_13849);
nor U17853 (N_17853,N_14761,N_12707);
and U17854 (N_17854,N_13569,N_14722);
nand U17855 (N_17855,N_13499,N_12917);
xnor U17856 (N_17856,N_13811,N_12148);
xor U17857 (N_17857,N_12969,N_12305);
or U17858 (N_17858,N_14454,N_14576);
nand U17859 (N_17859,N_13236,N_12208);
xnor U17860 (N_17860,N_12867,N_12273);
and U17861 (N_17861,N_14322,N_13957);
xnor U17862 (N_17862,N_14615,N_14885);
nand U17863 (N_17863,N_12288,N_12010);
nand U17864 (N_17864,N_12578,N_14540);
and U17865 (N_17865,N_12637,N_14645);
or U17866 (N_17866,N_13185,N_13490);
xor U17867 (N_17867,N_14930,N_12412);
or U17868 (N_17868,N_12255,N_14893);
xor U17869 (N_17869,N_13373,N_14722);
and U17870 (N_17870,N_12053,N_13631);
or U17871 (N_17871,N_14587,N_14493);
or U17872 (N_17872,N_13380,N_13302);
or U17873 (N_17873,N_14134,N_13201);
nand U17874 (N_17874,N_13947,N_13262);
or U17875 (N_17875,N_12506,N_12738);
nand U17876 (N_17876,N_13122,N_14098);
and U17877 (N_17877,N_14323,N_14431);
nand U17878 (N_17878,N_12883,N_13276);
or U17879 (N_17879,N_13416,N_12084);
nor U17880 (N_17880,N_12876,N_14747);
nand U17881 (N_17881,N_12303,N_12353);
nand U17882 (N_17882,N_13881,N_13134);
or U17883 (N_17883,N_13930,N_13660);
nor U17884 (N_17884,N_14344,N_13469);
xor U17885 (N_17885,N_13483,N_14765);
or U17886 (N_17886,N_12287,N_14719);
and U17887 (N_17887,N_12181,N_13921);
xor U17888 (N_17888,N_14203,N_13588);
nor U17889 (N_17889,N_12440,N_12379);
xnor U17890 (N_17890,N_14455,N_14546);
or U17891 (N_17891,N_14802,N_12370);
xnor U17892 (N_17892,N_12391,N_13846);
nand U17893 (N_17893,N_13418,N_14265);
xor U17894 (N_17894,N_12911,N_14990);
xor U17895 (N_17895,N_14189,N_13948);
or U17896 (N_17896,N_13643,N_12435);
and U17897 (N_17897,N_13957,N_13116);
nand U17898 (N_17898,N_13581,N_14788);
xor U17899 (N_17899,N_14752,N_12721);
and U17900 (N_17900,N_14986,N_12179);
nand U17901 (N_17901,N_12560,N_14485);
nand U17902 (N_17902,N_14808,N_14806);
or U17903 (N_17903,N_14760,N_12403);
and U17904 (N_17904,N_12472,N_13367);
nand U17905 (N_17905,N_14147,N_14687);
or U17906 (N_17906,N_13903,N_12510);
xnor U17907 (N_17907,N_13227,N_13095);
or U17908 (N_17908,N_14685,N_13079);
xor U17909 (N_17909,N_14111,N_12293);
xor U17910 (N_17910,N_12473,N_12775);
xor U17911 (N_17911,N_12743,N_12056);
or U17912 (N_17912,N_12663,N_14823);
and U17913 (N_17913,N_14370,N_14488);
nand U17914 (N_17914,N_13729,N_14103);
nand U17915 (N_17915,N_12331,N_13533);
xnor U17916 (N_17916,N_13461,N_14634);
nor U17917 (N_17917,N_12153,N_14531);
or U17918 (N_17918,N_13720,N_14202);
nand U17919 (N_17919,N_14914,N_13142);
and U17920 (N_17920,N_14893,N_14414);
or U17921 (N_17921,N_13230,N_13113);
nand U17922 (N_17922,N_12124,N_14351);
nand U17923 (N_17923,N_12779,N_12562);
nor U17924 (N_17924,N_13138,N_13173);
or U17925 (N_17925,N_14173,N_14694);
xnor U17926 (N_17926,N_14040,N_13533);
or U17927 (N_17927,N_14829,N_12696);
or U17928 (N_17928,N_14595,N_14956);
and U17929 (N_17929,N_13488,N_12924);
nor U17930 (N_17930,N_13344,N_12901);
or U17931 (N_17931,N_12082,N_14744);
xnor U17932 (N_17932,N_14229,N_13905);
xor U17933 (N_17933,N_14734,N_14872);
nand U17934 (N_17934,N_13787,N_13987);
or U17935 (N_17935,N_12442,N_14003);
or U17936 (N_17936,N_13709,N_14139);
nand U17937 (N_17937,N_12902,N_13108);
nor U17938 (N_17938,N_14209,N_13379);
nor U17939 (N_17939,N_14322,N_13535);
nor U17940 (N_17940,N_13958,N_14978);
xor U17941 (N_17941,N_14564,N_14615);
or U17942 (N_17942,N_13273,N_12388);
xor U17943 (N_17943,N_13271,N_12336);
nor U17944 (N_17944,N_13478,N_14439);
nand U17945 (N_17945,N_13897,N_13066);
xor U17946 (N_17946,N_12302,N_14718);
nor U17947 (N_17947,N_13845,N_12478);
xor U17948 (N_17948,N_13459,N_14587);
nand U17949 (N_17949,N_12954,N_14920);
and U17950 (N_17950,N_13725,N_14031);
nand U17951 (N_17951,N_12287,N_14126);
and U17952 (N_17952,N_13113,N_13894);
nand U17953 (N_17953,N_14482,N_14569);
nor U17954 (N_17954,N_12777,N_14825);
and U17955 (N_17955,N_12340,N_13322);
nor U17956 (N_17956,N_13911,N_14461);
nand U17957 (N_17957,N_14308,N_13161);
nand U17958 (N_17958,N_14009,N_13149);
nand U17959 (N_17959,N_12543,N_14523);
nand U17960 (N_17960,N_14075,N_12509);
or U17961 (N_17961,N_14741,N_14456);
and U17962 (N_17962,N_14329,N_14590);
nand U17963 (N_17963,N_12783,N_12921);
nand U17964 (N_17964,N_14582,N_14042);
or U17965 (N_17965,N_12609,N_13859);
nor U17966 (N_17966,N_14470,N_13353);
xor U17967 (N_17967,N_12540,N_14669);
nand U17968 (N_17968,N_12772,N_13181);
nor U17969 (N_17969,N_14385,N_14252);
xor U17970 (N_17970,N_12255,N_14734);
and U17971 (N_17971,N_13042,N_13200);
or U17972 (N_17972,N_13458,N_14419);
nor U17973 (N_17973,N_14532,N_13730);
or U17974 (N_17974,N_14295,N_13643);
nor U17975 (N_17975,N_13286,N_14649);
or U17976 (N_17976,N_14079,N_12273);
nor U17977 (N_17977,N_14916,N_12583);
nand U17978 (N_17978,N_12539,N_12009);
nor U17979 (N_17979,N_12368,N_12688);
or U17980 (N_17980,N_13271,N_14754);
and U17981 (N_17981,N_12884,N_12970);
nand U17982 (N_17982,N_14066,N_13086);
nand U17983 (N_17983,N_14586,N_14393);
and U17984 (N_17984,N_13370,N_12109);
nand U17985 (N_17985,N_12878,N_14282);
nand U17986 (N_17986,N_12105,N_12456);
nand U17987 (N_17987,N_13937,N_12608);
and U17988 (N_17988,N_14814,N_12909);
xor U17989 (N_17989,N_12008,N_12411);
and U17990 (N_17990,N_14678,N_14635);
and U17991 (N_17991,N_12240,N_13610);
nor U17992 (N_17992,N_13241,N_14253);
or U17993 (N_17993,N_13999,N_12993);
xor U17994 (N_17994,N_14607,N_13786);
nand U17995 (N_17995,N_12562,N_14300);
or U17996 (N_17996,N_13167,N_13573);
nand U17997 (N_17997,N_12386,N_12463);
nand U17998 (N_17998,N_13686,N_12844);
nand U17999 (N_17999,N_14754,N_12203);
and U18000 (N_18000,N_16710,N_17034);
nor U18001 (N_18001,N_15225,N_15548);
nor U18002 (N_18002,N_15204,N_16819);
or U18003 (N_18003,N_17552,N_17210);
xnor U18004 (N_18004,N_15198,N_15592);
xor U18005 (N_18005,N_16107,N_16502);
nand U18006 (N_18006,N_15110,N_17207);
and U18007 (N_18007,N_15701,N_15051);
and U18008 (N_18008,N_16992,N_15777);
xnor U18009 (N_18009,N_17592,N_15449);
or U18010 (N_18010,N_16425,N_17040);
xnor U18011 (N_18011,N_17478,N_17279);
nor U18012 (N_18012,N_16128,N_16082);
xor U18013 (N_18013,N_16779,N_16040);
and U18014 (N_18014,N_17159,N_15055);
xor U18015 (N_18015,N_15597,N_16575);
xnor U18016 (N_18016,N_15221,N_17303);
or U18017 (N_18017,N_15950,N_16858);
nor U18018 (N_18018,N_17182,N_16121);
xor U18019 (N_18019,N_17025,N_17358);
nand U18020 (N_18020,N_17075,N_15457);
and U18021 (N_18021,N_16822,N_15177);
or U18022 (N_18022,N_17692,N_17878);
and U18023 (N_18023,N_17440,N_15947);
or U18024 (N_18024,N_16063,N_15222);
or U18025 (N_18025,N_16785,N_15547);
nand U18026 (N_18026,N_16682,N_16772);
or U18027 (N_18027,N_16247,N_15971);
nor U18028 (N_18028,N_15923,N_16230);
and U18029 (N_18029,N_15212,N_15027);
or U18030 (N_18030,N_17931,N_17448);
nand U18031 (N_18031,N_15305,N_15644);
xor U18032 (N_18032,N_16348,N_17548);
xor U18033 (N_18033,N_15507,N_16621);
xor U18034 (N_18034,N_15797,N_17164);
xnor U18035 (N_18035,N_15303,N_15307);
and U18036 (N_18036,N_17869,N_16595);
nand U18037 (N_18037,N_15493,N_15076);
or U18038 (N_18038,N_15530,N_15418);
xnor U18039 (N_18039,N_15640,N_16359);
and U18040 (N_18040,N_17140,N_16852);
nor U18041 (N_18041,N_16314,N_17752);
nand U18042 (N_18042,N_17174,N_16672);
nand U18043 (N_18043,N_16316,N_16665);
nand U18044 (N_18044,N_15991,N_15869);
nand U18045 (N_18045,N_17915,N_16109);
xor U18046 (N_18046,N_17235,N_15151);
and U18047 (N_18047,N_16973,N_16214);
nand U18048 (N_18048,N_15004,N_17476);
nand U18049 (N_18049,N_15282,N_17428);
or U18050 (N_18050,N_16959,N_17888);
nor U18051 (N_18051,N_17744,N_15613);
and U18052 (N_18052,N_15271,N_15014);
nand U18053 (N_18053,N_16315,N_15785);
nand U18054 (N_18054,N_16988,N_17222);
xor U18055 (N_18055,N_16846,N_15501);
or U18056 (N_18056,N_15178,N_16465);
nand U18057 (N_18057,N_15734,N_15099);
xor U18058 (N_18058,N_16748,N_17788);
xor U18059 (N_18059,N_17800,N_15108);
or U18060 (N_18060,N_15060,N_16380);
or U18061 (N_18061,N_16260,N_15363);
xor U18062 (N_18062,N_16454,N_16923);
and U18063 (N_18063,N_15525,N_15480);
nor U18064 (N_18064,N_16309,N_17731);
xor U18065 (N_18065,N_17155,N_15728);
xnor U18066 (N_18066,N_15917,N_16137);
or U18067 (N_18067,N_16663,N_17350);
and U18068 (N_18068,N_17759,N_17540);
nor U18069 (N_18069,N_16352,N_16675);
xnor U18070 (N_18070,N_15850,N_15649);
xnor U18071 (N_18071,N_16531,N_17755);
xnor U18072 (N_18072,N_15145,N_15870);
nor U18073 (N_18073,N_16911,N_17468);
nand U18074 (N_18074,N_16277,N_15364);
and U18075 (N_18075,N_15703,N_17770);
xor U18076 (N_18076,N_17223,N_16242);
nor U18077 (N_18077,N_16151,N_17785);
xor U18078 (N_18078,N_16090,N_17310);
xor U18079 (N_18079,N_17580,N_16524);
and U18080 (N_18080,N_15065,N_17783);
and U18081 (N_18081,N_16202,N_17495);
nor U18082 (N_18082,N_15074,N_15506);
nor U18083 (N_18083,N_17444,N_17097);
nand U18084 (N_18084,N_17370,N_16792);
nor U18085 (N_18085,N_17005,N_16256);
nand U18086 (N_18086,N_15328,N_16039);
xnor U18087 (N_18087,N_15391,N_16170);
and U18088 (N_18088,N_17126,N_17679);
and U18089 (N_18089,N_15126,N_17359);
or U18090 (N_18090,N_16186,N_17704);
nor U18091 (N_18091,N_15340,N_15512);
nand U18092 (N_18092,N_17176,N_15849);
nand U18093 (N_18093,N_16673,N_17417);
xor U18094 (N_18094,N_15643,N_15717);
and U18095 (N_18095,N_17137,N_15022);
or U18096 (N_18096,N_17001,N_17747);
and U18097 (N_18097,N_17424,N_17911);
xor U18098 (N_18098,N_17095,N_16219);
or U18099 (N_18099,N_15087,N_16335);
nand U18100 (N_18100,N_17934,N_17905);
or U18101 (N_18101,N_17172,N_17718);
nor U18102 (N_18102,N_17339,N_16861);
xor U18103 (N_18103,N_16190,N_15240);
nor U18104 (N_18104,N_17967,N_16643);
xor U18105 (N_18105,N_17925,N_17923);
nand U18106 (N_18106,N_15908,N_15799);
xnor U18107 (N_18107,N_15281,N_16047);
and U18108 (N_18108,N_17062,N_16737);
xnor U18109 (N_18109,N_17618,N_17741);
nor U18110 (N_18110,N_15387,N_17936);
and U18111 (N_18111,N_16842,N_17166);
or U18112 (N_18112,N_17248,N_16525);
and U18113 (N_18113,N_15733,N_15732);
xor U18114 (N_18114,N_15628,N_17456);
or U18115 (N_18115,N_16432,N_17139);
nand U18116 (N_18116,N_16704,N_17870);
and U18117 (N_18117,N_17985,N_17865);
nor U18118 (N_18118,N_15651,N_16383);
and U18119 (N_18119,N_16141,N_17883);
and U18120 (N_18120,N_17876,N_15535);
nand U18121 (N_18121,N_17828,N_17067);
nand U18122 (N_18122,N_17304,N_17290);
nand U18123 (N_18123,N_15740,N_17682);
or U18124 (N_18124,N_17503,N_17617);
nor U18125 (N_18125,N_17494,N_15447);
and U18126 (N_18126,N_15784,N_16452);
nand U18127 (N_18127,N_16903,N_16386);
nor U18128 (N_18128,N_15653,N_16323);
nand U18129 (N_18129,N_15372,N_15593);
or U18130 (N_18130,N_15309,N_15793);
nand U18131 (N_18131,N_15350,N_16101);
nor U18132 (N_18132,N_16617,N_17107);
xnor U18133 (N_18133,N_15301,N_15521);
nor U18134 (N_18134,N_16409,N_17365);
or U18135 (N_18135,N_17406,N_17302);
xnor U18136 (N_18136,N_16909,N_17746);
or U18137 (N_18137,N_15005,N_16000);
xnor U18138 (N_18138,N_15952,N_15009);
nor U18139 (N_18139,N_17257,N_16150);
or U18140 (N_18140,N_15105,N_16180);
or U18141 (N_18141,N_15646,N_15623);
nor U18142 (N_18142,N_16793,N_17945);
nand U18143 (N_18143,N_16120,N_15633);
xor U18144 (N_18144,N_17334,N_15824);
or U18145 (N_18145,N_16577,N_15999);
nand U18146 (N_18146,N_15851,N_17829);
and U18147 (N_18147,N_16205,N_17397);
or U18148 (N_18148,N_15490,N_15515);
nor U18149 (N_18149,N_15378,N_17342);
nand U18150 (N_18150,N_16915,N_17994);
or U18151 (N_18151,N_17316,N_16060);
nor U18152 (N_18152,N_16631,N_16178);
nor U18153 (N_18153,N_17863,N_16510);
and U18154 (N_18154,N_16559,N_16354);
xor U18155 (N_18155,N_17465,N_16399);
nor U18156 (N_18156,N_15499,N_17029);
and U18157 (N_18157,N_17063,N_17946);
or U18158 (N_18158,N_17846,N_16865);
or U18159 (N_18159,N_15580,N_16317);
nor U18160 (N_18160,N_15796,N_16468);
nor U18161 (N_18161,N_16290,N_17845);
xor U18162 (N_18162,N_16055,N_15086);
and U18163 (N_18163,N_17249,N_17916);
and U18164 (N_18164,N_17535,N_17028);
nor U18165 (N_18165,N_15787,N_16805);
nor U18166 (N_18166,N_15285,N_17857);
xnor U18167 (N_18167,N_16523,N_17115);
and U18168 (N_18168,N_15517,N_15617);
nand U18169 (N_18169,N_16308,N_17412);
or U18170 (N_18170,N_17577,N_17670);
or U18171 (N_18171,N_15738,N_17099);
nand U18172 (N_18172,N_15829,N_17357);
nand U18173 (N_18173,N_17823,N_16760);
nand U18174 (N_18174,N_17361,N_15250);
or U18175 (N_18175,N_17367,N_16810);
xnor U18176 (N_18176,N_17726,N_17642);
and U18177 (N_18177,N_15558,N_15470);
xor U18178 (N_18178,N_15163,N_16567);
xnor U18179 (N_18179,N_17343,N_17254);
nand U18180 (N_18180,N_15524,N_16435);
nor U18181 (N_18181,N_17344,N_17707);
or U18182 (N_18182,N_16372,N_16881);
and U18183 (N_18183,N_15583,N_15555);
xor U18184 (N_18184,N_15046,N_16770);
nand U18185 (N_18185,N_16393,N_15531);
and U18186 (N_18186,N_15909,N_16773);
nor U18187 (N_18187,N_16897,N_16823);
and U18188 (N_18188,N_16778,N_16657);
nand U18189 (N_18189,N_16255,N_16882);
or U18190 (N_18190,N_17982,N_15397);
and U18191 (N_18191,N_15533,N_15868);
xor U18192 (N_18192,N_16262,N_15919);
or U18193 (N_18193,N_15456,N_15011);
nand U18194 (N_18194,N_16200,N_17204);
nand U18195 (N_18195,N_16099,N_16946);
nor U18196 (N_18196,N_16596,N_15172);
and U18197 (N_18197,N_17449,N_15509);
and U18198 (N_18198,N_16056,N_16723);
nor U18199 (N_18199,N_17947,N_15473);
nor U18200 (N_18200,N_17308,N_15492);
or U18201 (N_18201,N_17672,N_15805);
nand U18202 (N_18202,N_16431,N_15820);
nor U18203 (N_18203,N_16173,N_17639);
nor U18204 (N_18204,N_17033,N_17162);
nand U18205 (N_18205,N_17724,N_16686);
and U18206 (N_18206,N_17401,N_16470);
xor U18207 (N_18207,N_17206,N_15903);
xor U18208 (N_18208,N_16720,N_15636);
or U18209 (N_18209,N_16949,N_17524);
and U18210 (N_18210,N_15168,N_16730);
nor U18211 (N_18211,N_15959,N_15306);
and U18212 (N_18212,N_16463,N_17558);
xnor U18213 (N_18213,N_15957,N_17708);
or U18214 (N_18214,N_16649,N_16586);
nand U18215 (N_18215,N_17442,N_16397);
nand U18216 (N_18216,N_17133,N_15462);
nor U18217 (N_18217,N_15056,N_15135);
xor U18218 (N_18218,N_15203,N_15812);
and U18219 (N_18219,N_15357,N_15128);
nand U18220 (N_18220,N_16123,N_16118);
nor U18221 (N_18221,N_15990,N_16052);
nand U18222 (N_18222,N_17842,N_16320);
xor U18223 (N_18223,N_17196,N_16257);
and U18224 (N_18224,N_17723,N_16957);
and U18225 (N_18225,N_17362,N_16168);
nand U18226 (N_18226,N_17472,N_16441);
nand U18227 (N_18227,N_15472,N_17898);
or U18228 (N_18228,N_16342,N_15152);
or U18229 (N_18229,N_15043,N_17651);
nand U18230 (N_18230,N_17252,N_16940);
xor U18231 (N_18231,N_16215,N_16513);
and U18232 (N_18232,N_17125,N_16696);
nand U18233 (N_18233,N_16222,N_17854);
or U18234 (N_18234,N_15468,N_15325);
and U18235 (N_18235,N_15070,N_16297);
and U18236 (N_18236,N_17022,N_16722);
nor U18237 (N_18237,N_16824,N_15474);
and U18238 (N_18238,N_17766,N_15230);
xor U18239 (N_18239,N_15657,N_16300);
nor U18240 (N_18240,N_16693,N_17169);
and U18241 (N_18241,N_16856,N_16018);
nand U18242 (N_18242,N_16493,N_16305);
or U18243 (N_18243,N_17259,N_17669);
nor U18244 (N_18244,N_17879,N_16351);
or U18245 (N_18245,N_15833,N_17505);
and U18246 (N_18246,N_16880,N_17268);
xor U18247 (N_18247,N_17804,N_16296);
or U18248 (N_18248,N_15131,N_15708);
and U18249 (N_18249,N_15928,N_15430);
xnor U18250 (N_18250,N_17073,N_17044);
nand U18251 (N_18251,N_17289,N_17461);
nor U18252 (N_18252,N_17602,N_16014);
nand U18253 (N_18253,N_16166,N_17212);
and U18254 (N_18254,N_16991,N_15402);
nand U18255 (N_18255,N_16122,N_15299);
or U18256 (N_18256,N_16248,N_17398);
nor U18257 (N_18257,N_15932,N_16232);
nand U18258 (N_18258,N_16618,N_16484);
nand U18259 (N_18259,N_17112,N_16045);
or U18260 (N_18260,N_15293,N_16240);
and U18261 (N_18261,N_17630,N_16345);
nand U18262 (N_18262,N_16560,N_15366);
xnor U18263 (N_18263,N_17691,N_17856);
or U18264 (N_18264,N_17563,N_17754);
and U18265 (N_18265,N_16945,N_17794);
xnor U18266 (N_18266,N_17861,N_16442);
or U18267 (N_18267,N_17955,N_16002);
and U18268 (N_18268,N_17699,N_15232);
nor U18269 (N_18269,N_16612,N_15542);
and U18270 (N_18270,N_15763,N_15977);
xor U18271 (N_18271,N_15111,N_16189);
nand U18272 (N_18272,N_17502,N_16936);
nor U18273 (N_18273,N_17802,N_16542);
xnor U18274 (N_18274,N_17853,N_15253);
nor U18275 (N_18275,N_15611,N_16456);
or U18276 (N_18276,N_15469,N_16754);
or U18277 (N_18277,N_16830,N_16377);
nand U18278 (N_18278,N_15434,N_17745);
nor U18279 (N_18279,N_17090,N_16854);
xnor U18280 (N_18280,N_16826,N_15933);
and U18281 (N_18281,N_16637,N_16685);
xnor U18282 (N_18282,N_15544,N_17253);
nand U18283 (N_18283,N_17706,N_16263);
xnor U18284 (N_18284,N_16193,N_15992);
nor U18285 (N_18285,N_15026,N_15445);
or U18286 (N_18286,N_17065,N_16648);
nand U18287 (N_18287,N_15599,N_16184);
nand U18288 (N_18288,N_17922,N_17740);
xnor U18289 (N_18289,N_17305,N_17015);
or U18290 (N_18290,N_17141,N_16281);
or U18291 (N_18291,N_17056,N_17607);
or U18292 (N_18292,N_16952,N_16117);
xnor U18293 (N_18293,N_16816,N_17330);
nand U18294 (N_18294,N_16788,N_16552);
nor U18295 (N_18295,N_15416,N_16546);
nor U18296 (N_18296,N_15714,N_17559);
xnor U18297 (N_18297,N_17710,N_16644);
nor U18298 (N_18298,N_16970,N_16774);
xnor U18299 (N_18299,N_16691,N_16750);
and U18300 (N_18300,N_15813,N_17980);
xor U18301 (N_18301,N_17241,N_15088);
nor U18302 (N_18302,N_16238,N_16016);
or U18303 (N_18303,N_17003,N_17652);
or U18304 (N_18304,N_17657,N_16356);
nor U18305 (N_18305,N_15514,N_16346);
or U18306 (N_18306,N_16850,N_16536);
nand U18307 (N_18307,N_17180,N_17732);
nor U18308 (N_18308,N_17292,N_17455);
and U18309 (N_18309,N_17531,N_16600);
nor U18310 (N_18310,N_17262,N_16494);
or U18311 (N_18311,N_16216,N_15421);
xnor U18312 (N_18312,N_17519,N_16258);
xnor U18313 (N_18313,N_15414,N_16243);
nor U18314 (N_18314,N_17250,N_17722);
nand U18315 (N_18315,N_15886,N_15655);
or U18316 (N_18316,N_17434,N_15031);
xnor U18317 (N_18317,N_17625,N_17506);
or U18318 (N_18318,N_17728,N_16831);
or U18319 (N_18319,N_17532,N_16934);
and U18320 (N_18320,N_17909,N_15518);
nor U18321 (N_18321,N_17390,N_16716);
or U18322 (N_18322,N_17020,N_16944);
nand U18323 (N_18323,N_17463,N_16509);
xor U18324 (N_18324,N_15774,N_16384);
or U18325 (N_18325,N_15124,N_15395);
and U18326 (N_18326,N_15975,N_16094);
nand U18327 (N_18327,N_16653,N_16956);
or U18328 (N_18328,N_16592,N_16076);
xnor U18329 (N_18329,N_17427,N_17321);
and U18330 (N_18330,N_15386,N_16872);
or U18331 (N_18331,N_17817,N_16385);
nor U18332 (N_18332,N_16809,N_17232);
nor U18333 (N_18333,N_15685,N_17464);
nand U18334 (N_18334,N_17533,N_15401);
xnor U18335 (N_18335,N_16964,N_17293);
xor U18336 (N_18336,N_15164,N_17366);
nor U18337 (N_18337,N_17084,N_16904);
xnor U18338 (N_18338,N_15446,N_16475);
and U18339 (N_18339,N_16153,N_15193);
and U18340 (N_18340,N_15876,N_15195);
and U18341 (N_18341,N_15931,N_16280);
or U18342 (N_18342,N_15697,N_16514);
and U18343 (N_18343,N_15883,N_17121);
xnor U18344 (N_18344,N_15093,N_15254);
and U18345 (N_18345,N_17144,N_17481);
or U18346 (N_18346,N_17534,N_17437);
xnor U18347 (N_18347,N_17806,N_17076);
nand U18348 (N_18348,N_17010,N_17251);
nor U18349 (N_18349,N_15537,N_16044);
xnor U18350 (N_18350,N_16995,N_16229);
and U18351 (N_18351,N_17753,N_15737);
xor U18352 (N_18352,N_15696,N_15113);
nand U18353 (N_18353,N_16553,N_15940);
nand U18354 (N_18354,N_17064,N_15405);
or U18355 (N_18355,N_17388,N_16389);
nor U18356 (N_18356,N_17407,N_15141);
or U18357 (N_18357,N_17697,N_16129);
or U18358 (N_18358,N_17522,N_17123);
nor U18359 (N_18359,N_16789,N_17263);
nor U18360 (N_18360,N_17938,N_15879);
nand U18361 (N_18361,N_17668,N_15077);
and U18362 (N_18362,N_16448,N_15795);
or U18363 (N_18363,N_15780,N_16848);
nor U18364 (N_18364,N_15138,N_17995);
xor U18365 (N_18365,N_17487,N_16261);
nor U18366 (N_18366,N_17491,N_16570);
nor U18367 (N_18367,N_16837,N_16426);
or U18368 (N_18368,N_16495,N_15602);
nor U18369 (N_18369,N_17106,N_16656);
or U18370 (N_18370,N_17644,N_16558);
xor U18371 (N_18371,N_17709,N_17261);
nor U18372 (N_18372,N_17544,N_15461);
or U18373 (N_18373,N_17269,N_16642);
nand U18374 (N_18374,N_15144,N_16864);
nor U18375 (N_18375,N_17683,N_16607);
or U18376 (N_18376,N_16931,N_16947);
or U18377 (N_18377,N_15609,N_17874);
nor U18378 (N_18378,N_16102,N_17430);
and U18379 (N_18379,N_15190,N_16587);
nand U18380 (N_18380,N_16252,N_15559);
nor U18381 (N_18381,N_16270,N_17647);
or U18382 (N_18382,N_16086,N_16025);
nand U18383 (N_18383,N_17404,N_17812);
nor U18384 (N_18384,N_17658,N_17217);
xor U18385 (N_18385,N_17323,N_16884);
nand U18386 (N_18386,N_16417,N_17892);
xnor U18387 (N_18387,N_17243,N_17153);
and U18388 (N_18388,N_16119,N_15755);
nor U18389 (N_18389,N_17963,N_15771);
nand U18390 (N_18390,N_17114,N_16438);
and U18391 (N_18391,N_15384,N_16590);
or U18392 (N_18392,N_15188,N_17192);
xor U18393 (N_18393,N_15718,N_17059);
xor U18394 (N_18394,N_17187,N_17486);
and U18395 (N_18395,N_16954,N_17315);
xnor U18396 (N_18396,N_16874,N_15625);
and U18397 (N_18397,N_16888,N_17171);
and U18398 (N_18398,N_15690,N_17805);
xnor U18399 (N_18399,N_15598,N_15516);
or U18400 (N_18400,N_15098,N_15921);
or U18401 (N_18401,N_15966,N_16289);
nand U18402 (N_18402,N_16985,N_17046);
xnor U18403 (N_18403,N_16591,N_16133);
or U18404 (N_18404,N_16980,N_16478);
nor U18405 (N_18405,N_16896,N_16440);
nand U18406 (N_18406,N_17193,N_15295);
or U18407 (N_18407,N_15429,N_16906);
and U18408 (N_18408,N_16111,N_16622);
xnor U18409 (N_18409,N_17662,N_15639);
or U18410 (N_18410,N_16530,N_17234);
or U18411 (N_18411,N_16635,N_17637);
nand U18412 (N_18412,N_15143,N_16311);
xnor U18413 (N_18413,N_15853,N_17498);
or U18414 (N_18414,N_15608,N_15897);
and U18415 (N_18415,N_15283,N_15032);
nor U18416 (N_18416,N_16914,N_15692);
nor U18417 (N_18417,N_15782,N_16035);
nor U18418 (N_18418,N_17284,N_17680);
nor U18419 (N_18419,N_16902,N_17395);
or U18420 (N_18420,N_16011,N_15510);
and U18421 (N_18421,N_15223,N_15007);
or U18422 (N_18422,N_16528,N_17958);
nor U18423 (N_18423,N_16955,N_15688);
xor U18424 (N_18424,N_15552,N_16030);
nand U18425 (N_18425,N_15370,N_17979);
nor U18426 (N_18426,N_16376,N_16332);
and U18427 (N_18427,N_16267,N_17283);
and U18428 (N_18428,N_16436,N_15687);
or U18429 (N_18429,N_17055,N_17897);
and U18430 (N_18430,N_16428,N_16654);
nor U18431 (N_18431,N_17542,N_17821);
or U18432 (N_18432,N_16961,N_17500);
and U18433 (N_18433,N_16913,N_15330);
nand U18434 (N_18434,N_16547,N_15067);
xnor U18435 (N_18435,N_15615,N_17240);
nand U18436 (N_18436,N_16767,N_17891);
nor U18437 (N_18437,N_17031,N_17151);
nor U18438 (N_18438,N_15332,N_17932);
nor U18439 (N_18439,N_15383,N_16646);
nor U18440 (N_18440,N_15484,N_17173);
nor U18441 (N_18441,N_17296,N_17274);
or U18442 (N_18442,N_15245,N_17860);
nand U18443 (N_18443,N_15288,N_16501);
or U18444 (N_18444,N_17808,N_15995);
nand U18445 (N_18445,N_17087,N_16917);
nand U18446 (N_18446,N_17036,N_16391);
xnor U18447 (N_18447,N_17526,N_17624);
and U18448 (N_18448,N_17083,N_15816);
and U18449 (N_18449,N_17632,N_17886);
and U18450 (N_18450,N_16678,N_15845);
or U18451 (N_18451,N_17110,N_16937);
or U18452 (N_18452,N_15567,N_16160);
and U18453 (N_18453,N_17893,N_15902);
or U18454 (N_18454,N_16185,N_16163);
nor U18455 (N_18455,N_16085,N_17373);
xor U18456 (N_18456,N_15907,N_15441);
xor U18457 (N_18457,N_15064,N_15508);
xor U18458 (N_18458,N_17676,N_15175);
xor U18459 (N_18459,N_17997,N_16797);
nand U18460 (N_18460,N_15308,N_16042);
nor U18461 (N_18461,N_17285,N_16387);
and U18462 (N_18462,N_17940,N_16043);
nand U18463 (N_18463,N_17978,N_15422);
nand U18464 (N_18464,N_16585,N_17213);
or U18465 (N_18465,N_17445,N_15182);
nand U18466 (N_18466,N_17007,N_16887);
xor U18467 (N_18467,N_15197,N_17807);
nor U18468 (N_18468,N_15626,N_15498);
nand U18469 (N_18469,N_17017,N_16994);
xnor U18470 (N_18470,N_17514,N_17962);
or U18471 (N_18471,N_16814,N_15585);
xor U18472 (N_18472,N_16694,N_15437);
or U18473 (N_18473,N_16464,N_17094);
and U18474 (N_18474,N_17271,N_15008);
nor U18475 (N_18475,N_15930,N_15601);
or U18476 (N_18476,N_15003,N_17457);
and U18477 (N_18477,N_17372,N_15236);
and U18478 (N_18478,N_17411,N_16540);
or U18479 (N_18479,N_15491,N_15169);
nand U18480 (N_18480,N_17971,N_17131);
or U18481 (N_18481,N_15237,N_17555);
xnor U18482 (N_18482,N_16195,N_15258);
and U18483 (N_18483,N_16863,N_15400);
nand U18484 (N_18484,N_17386,N_16924);
or U18485 (N_18485,N_15691,N_15037);
or U18486 (N_18486,N_15286,N_15112);
nand U18487 (N_18487,N_16899,N_17363);
xor U18488 (N_18488,N_16427,N_16535);
nor U18489 (N_18489,N_17267,N_15803);
or U18490 (N_18490,N_15800,N_17170);
nor U18491 (N_18491,N_17499,N_17633);
or U18492 (N_18492,N_15716,N_16796);
or U18493 (N_18493,N_16217,N_16496);
nand U18494 (N_18494,N_15442,N_16048);
nor U18495 (N_18495,N_17554,N_15511);
nand U18496 (N_18496,N_16538,N_17954);
nor U18497 (N_18497,N_16095,N_17135);
nand U18498 (N_18498,N_15749,N_16533);
or U18499 (N_18499,N_15668,N_17684);
nand U18500 (N_18500,N_16413,N_17834);
nand U18501 (N_18501,N_15465,N_16410);
nor U18502 (N_18502,N_17772,N_15888);
or U18503 (N_18503,N_15209,N_17523);
nor U18504 (N_18504,N_15606,N_17439);
nand U18505 (N_18505,N_16294,N_15810);
nand U18506 (N_18506,N_15089,N_17681);
nand U18507 (N_18507,N_17629,N_17881);
nand U18508 (N_18508,N_15454,N_15998);
xor U18509 (N_18509,N_15631,N_17027);
xnor U18510 (N_18510,N_15247,N_17609);
nor U18511 (N_18511,N_15541,N_16777);
nand U18512 (N_18512,N_15068,N_15746);
and U18513 (N_18513,N_16791,N_17214);
xnor U18514 (N_18514,N_16889,N_16813);
xor U18515 (N_18515,N_16006,N_16106);
nor U18516 (N_18516,N_16479,N_17275);
xor U18517 (N_18517,N_15864,N_17917);
or U18518 (N_18518,N_15607,N_17590);
nand U18519 (N_18519,N_17787,N_16999);
nand U18520 (N_18520,N_15565,N_16689);
xor U18521 (N_18521,N_17205,N_15083);
nor U18522 (N_18522,N_15321,N_15277);
or U18523 (N_18523,N_15039,N_17968);
nor U18524 (N_18524,N_15289,N_17689);
nand U18525 (N_18525,N_16581,N_16683);
and U18526 (N_18526,N_16825,N_17900);
nor U18527 (N_18527,N_15276,N_17935);
xnor U18528 (N_18528,N_16091,N_15844);
nand U18529 (N_18529,N_15148,N_17749);
and U18530 (N_18530,N_15153,N_16755);
or U18531 (N_18531,N_15762,N_15486);
and U18532 (N_18532,N_15589,N_17983);
nor U18533 (N_18533,N_17714,N_17122);
and U18534 (N_18534,N_15877,N_15926);
nor U18535 (N_18535,N_17286,N_17830);
xor U18536 (N_18536,N_15048,N_17128);
nor U18537 (N_18537,N_15960,N_17826);
xnor U18538 (N_18538,N_16659,N_16027);
or U18539 (N_18539,N_15489,N_17760);
xnor U18540 (N_18540,N_17574,N_17178);
nor U18541 (N_18541,N_17483,N_16605);
nand U18542 (N_18542,N_15072,N_15215);
xnor U18543 (N_18543,N_15720,N_16782);
xor U18544 (N_18544,N_16148,N_17762);
and U18545 (N_18545,N_17018,N_16976);
and U18546 (N_18546,N_17237,N_17833);
nand U18547 (N_18547,N_17231,N_17646);
or U18548 (N_18548,N_15794,N_16097);
nor U18549 (N_18549,N_17795,N_17438);
or U18550 (N_18550,N_15231,N_17179);
and U18551 (N_18551,N_17039,N_17453);
nand U18552 (N_18552,N_16334,N_16670);
nor U18553 (N_18553,N_16124,N_15412);
and U18554 (N_18554,N_15938,N_17282);
xnor U18555 (N_18555,N_15379,N_16511);
xor U18556 (N_18556,N_16588,N_15951);
and U18557 (N_18557,N_17216,N_16114);
nor U18558 (N_18558,N_16667,N_16818);
nor U18559 (N_18559,N_15673,N_17104);
and U18560 (N_18560,N_17729,N_17661);
and U18561 (N_18561,N_16972,N_15572);
xor U18562 (N_18562,N_17621,N_17675);
nor U18563 (N_18563,N_15553,N_16405);
nor U18564 (N_18564,N_16333,N_16894);
nand U18565 (N_18565,N_17318,N_15171);
xor U18566 (N_18566,N_15858,N_17380);
nor U18567 (N_18567,N_16574,N_15410);
or U18568 (N_18568,N_16028,N_16662);
xnor U18569 (N_18569,N_16004,N_16740);
nor U18570 (N_18570,N_16224,N_15843);
nor U18571 (N_18571,N_17884,N_15176);
nor U18572 (N_18572,N_17026,N_15248);
xor U18573 (N_18573,N_15373,N_16871);
and U18574 (N_18574,N_15246,N_16344);
nand U18575 (N_18575,N_16614,N_17100);
nor U18576 (N_18576,N_16299,N_15439);
and U18577 (N_18577,N_15768,N_16005);
nand U18578 (N_18578,N_15981,N_15546);
xnor U18579 (N_18579,N_16695,N_17069);
xnor U18580 (N_18580,N_17415,N_17197);
nor U18581 (N_18581,N_15823,N_16236);
or U18582 (N_18582,N_17432,N_15773);
and U18583 (N_18583,N_17391,N_17685);
nor U18584 (N_18584,N_15217,N_15841);
and U18585 (N_18585,N_15899,N_15375);
and U18586 (N_18586,N_15494,N_17451);
or U18587 (N_18587,N_17570,N_16507);
and U18588 (N_18588,N_15911,N_15677);
nor U18589 (N_18589,N_17085,N_15826);
xor U18590 (N_18590,N_15913,N_15670);
and U18591 (N_18591,N_15806,N_16794);
xnor U18592 (N_18592,N_17433,N_17188);
nor U18593 (N_18593,N_17466,N_15319);
nand U18594 (N_18594,N_15071,N_15754);
nand U18595 (N_18595,N_16024,N_17793);
nand U18596 (N_18596,N_16447,N_17421);
and U18597 (N_18597,N_15482,N_16420);
or U18598 (N_18598,N_16237,N_17414);
and U18599 (N_18599,N_16396,N_16753);
nand U18600 (N_18600,N_17376,N_15466);
nand U18601 (N_18601,N_17588,N_16563);
nand U18602 (N_18602,N_16449,N_17070);
and U18603 (N_18603,N_16568,N_16149);
or U18604 (N_18604,N_17566,N_16167);
or U18605 (N_18605,N_16572,N_17560);
and U18606 (N_18606,N_16977,N_15616);
xor U18607 (N_18607,N_15294,N_15239);
or U18608 (N_18608,N_17462,N_15028);
and U18609 (N_18609,N_16729,N_16968);
nor U18610 (N_18610,N_17004,N_16034);
xnor U18611 (N_18611,N_15622,N_15570);
nand U18612 (N_18612,N_15963,N_17377);
or U18613 (N_18613,N_15413,N_15582);
or U18614 (N_18614,N_15575,N_17998);
xnor U18615 (N_18615,N_16065,N_16071);
xor U18616 (N_18616,N_16481,N_16877);
nor U18617 (N_18617,N_16213,N_15100);
and U18618 (N_18618,N_15641,N_15619);
or U18619 (N_18619,N_16715,N_16981);
nand U18620 (N_18620,N_15808,N_17043);
nand U18621 (N_18621,N_15574,N_15958);
nor U18622 (N_18622,N_16081,N_17098);
and U18623 (N_18623,N_15130,N_16112);
xnor U18624 (N_18624,N_17727,N_17953);
xor U18625 (N_18625,N_16268,N_15929);
and U18626 (N_18626,N_17335,N_16015);
nand U18627 (N_18627,N_15343,N_16020);
or U18628 (N_18628,N_15573,N_17918);
and U18629 (N_18629,N_15669,N_17165);
xor U18630 (N_18630,N_16209,N_15117);
and U18631 (N_18631,N_16269,N_17903);
xor U18632 (N_18632,N_17300,N_17586);
xnor U18633 (N_18633,N_16226,N_15726);
or U18634 (N_18634,N_16009,N_15270);
or U18635 (N_18635,N_16241,N_15094);
nor U18636 (N_18636,N_16634,N_15035);
nand U18637 (N_18637,N_16851,N_17389);
and U18638 (N_18638,N_16343,N_17572);
or U18639 (N_18639,N_15165,N_17666);
and U18640 (N_18640,N_16327,N_15545);
xnor U18641 (N_18641,N_16049,N_17508);
or U18642 (N_18642,N_17118,N_16304);
nand U18643 (N_18643,N_17024,N_17482);
xnor U18644 (N_18644,N_15526,N_16744);
xnor U18645 (N_18645,N_15600,N_17183);
or U18646 (N_18646,N_15234,N_16893);
nand U18647 (N_18647,N_16278,N_15427);
or U18648 (N_18648,N_16749,N_16225);
or U18649 (N_18649,N_17635,N_17425);
and U18650 (N_18650,N_15791,N_15275);
xor U18651 (N_18651,N_16943,N_17778);
or U18652 (N_18652,N_16026,N_17847);
or U18653 (N_18653,N_17512,N_16768);
nand U18654 (N_18654,N_16404,N_17610);
nand U18655 (N_18655,N_15119,N_15403);
nand U18656 (N_18656,N_15896,N_15082);
or U18657 (N_18657,N_17603,N_15941);
and U18658 (N_18658,N_17902,N_16414);
xnor U18659 (N_18659,N_17981,N_15464);
xnor U18660 (N_18660,N_16482,N_16284);
or U18661 (N_18661,N_15778,N_15001);
and U18662 (N_18662,N_15536,N_16875);
xor U18663 (N_18663,N_16400,N_16669);
nor U18664 (N_18664,N_16998,N_15576);
xnor U18665 (N_18665,N_15310,N_17988);
nand U18666 (N_18666,N_17648,N_16506);
nand U18667 (N_18667,N_16781,N_17147);
nand U18668 (N_18668,N_15811,N_17711);
nor U18669 (N_18669,N_16761,N_15867);
or U18670 (N_18670,N_15139,N_15819);
nor U18671 (N_18671,N_17721,N_17048);
nand U18672 (N_18672,N_17096,N_15311);
and U18673 (N_18673,N_17735,N_16790);
nand U18674 (N_18674,N_15296,N_15300);
xnor U18675 (N_18675,N_15557,N_16029);
and U18676 (N_18676,N_17815,N_16834);
nand U18677 (N_18677,N_15924,N_17047);
or U18678 (N_18678,N_15362,N_17077);
or U18679 (N_18679,N_15292,N_15982);
or U18680 (N_18680,N_17751,N_15371);
nor U18681 (N_18681,N_17926,N_16445);
nand U18682 (N_18682,N_16145,N_17387);
and U18683 (N_18683,N_15114,N_16394);
and U18684 (N_18684,N_16233,N_16734);
and U18685 (N_18685,N_16313,N_15101);
or U18686 (N_18686,N_17734,N_16249);
and U18687 (N_18687,N_15632,N_17663);
nor U18688 (N_18688,N_15775,N_17576);
or U18689 (N_18689,N_17477,N_15360);
nand U18690 (N_18690,N_16161,N_16444);
nor U18691 (N_18691,N_17012,N_16870);
nor U18692 (N_18692,N_15715,N_15624);
and U18693 (N_18693,N_15885,N_17278);
and U18694 (N_18694,N_15842,N_16927);
nor U18695 (N_18695,N_16103,N_16053);
xor U18696 (N_18696,N_16878,N_16803);
and U18697 (N_18697,N_17416,N_16602);
or U18698 (N_18698,N_17490,N_17631);
or U18699 (N_18699,N_17696,N_15132);
nor U18700 (N_18700,N_17227,N_17791);
nand U18701 (N_18701,N_16077,N_17975);
xor U18702 (N_18702,N_15047,N_15409);
or U18703 (N_18703,N_17189,N_15652);
xor U18704 (N_18704,N_16157,N_16179);
and U18705 (N_18705,N_16548,N_17748);
nor U18706 (N_18706,N_15830,N_15873);
nor U18707 (N_18707,N_16584,N_17109);
or U18708 (N_18708,N_15199,N_17294);
or U18709 (N_18709,N_15080,N_16537);
and U18710 (N_18710,N_16922,N_17977);
or U18711 (N_18711,N_15770,N_16828);
xor U18712 (N_18712,N_15173,N_15393);
nand U18713 (N_18713,N_17260,N_16727);
or U18714 (N_18714,N_17939,N_15206);
xnor U18715 (N_18715,N_17774,N_16544);
xnor U18716 (N_18716,N_16197,N_16159);
nand U18717 (N_18717,N_15679,N_16008);
xor U18718 (N_18718,N_17858,N_16366);
nand U18719 (N_18719,N_15273,N_15835);
xnor U18720 (N_18720,N_15807,N_17654);
nand U18721 (N_18721,N_15662,N_17200);
and U18722 (N_18722,N_15459,N_17021);
and U18723 (N_18723,N_15694,N_16182);
xor U18724 (N_18724,N_15967,N_15396);
xor U18725 (N_18725,N_17352,N_15233);
nand U18726 (N_18726,N_17175,N_16876);
nor U18727 (N_18727,N_15380,N_16328);
xnor U18728 (N_18728,N_16728,N_16138);
xor U18729 (N_18729,N_16608,N_15936);
nor U18730 (N_18730,N_17620,N_17313);
nor U18731 (N_18731,N_15949,N_16175);
or U18732 (N_18732,N_16105,N_16485);
nor U18733 (N_18733,N_16879,N_16679);
or U18734 (N_18734,N_17203,N_16554);
nor U18735 (N_18735,N_15798,N_17006);
xnor U18736 (N_18736,N_16555,N_15002);
xnor U18737 (N_18737,N_16374,N_15066);
nor U18738 (N_18738,N_17215,N_17314);
nor U18739 (N_18739,N_17818,N_16703);
xor U18740 (N_18740,N_16520,N_15346);
or U18741 (N_18741,N_16579,N_15658);
nor U18742 (N_18742,N_17612,N_16259);
and U18743 (N_18743,N_16935,N_16726);
and U18744 (N_18744,N_15698,N_16467);
and U18745 (N_18745,N_17765,N_17695);
xnor U18746 (N_18746,N_15505,N_17513);
nor U18747 (N_18747,N_17068,N_15318);
or U18748 (N_18748,N_17536,N_17134);
or U18749 (N_18749,N_15398,N_15417);
or U18750 (N_18750,N_17674,N_16078);
nor U18751 (N_18751,N_15424,N_17509);
xor U18752 (N_18752,N_17547,N_17961);
xor U18753 (N_18753,N_15859,N_16821);
and U18754 (N_18754,N_16713,N_15551);
nor U18755 (N_18755,N_15502,N_16664);
nand U18756 (N_18756,N_16312,N_17181);
xnor U18757 (N_18757,N_17913,N_17019);
nor U18758 (N_18758,N_17720,N_17767);
nand U18759 (N_18759,N_17384,N_16933);
xor U18760 (N_18760,N_17340,N_16330);
or U18761 (N_18761,N_16181,N_15365);
nor U18762 (N_18762,N_17429,N_15865);
nor U18763 (N_18763,N_16827,N_17908);
and U18764 (N_18764,N_15133,N_16136);
nor U18765 (N_18765,N_15179,N_17375);
and U18766 (N_18766,N_16786,N_16812);
xor U18767 (N_18767,N_17790,N_15269);
nand U18768 (N_18768,N_16598,N_17667);
or U18769 (N_18769,N_16164,N_16687);
and U18770 (N_18770,N_15889,N_15905);
nand U18771 (N_18771,N_17264,N_17103);
nand U18772 (N_18772,N_17000,N_16966);
and U18773 (N_18773,N_17964,N_15109);
and U18774 (N_18774,N_17613,N_15970);
xnor U18775 (N_18775,N_17185,N_15590);
nand U18776 (N_18776,N_15290,N_15337);
or U18777 (N_18777,N_15219,N_17705);
and U18778 (N_18778,N_16938,N_16301);
xnor U18779 (N_18779,N_17443,N_15761);
nor U18780 (N_18780,N_16476,N_17156);
and U18781 (N_18781,N_16466,N_17297);
nand U18782 (N_18782,N_17937,N_15711);
nand U18783 (N_18783,N_15767,N_15727);
or U18784 (N_18784,N_16158,N_17545);
nand U18785 (N_18785,N_15106,N_17797);
or U18786 (N_18786,N_15050,N_16050);
xor U18787 (N_18787,N_15621,N_16364);
nor U18788 (N_18788,N_15729,N_17149);
or U18789 (N_18789,N_17822,N_15614);
and U18790 (N_18790,N_15045,N_15756);
nand U18791 (N_18791,N_17895,N_16844);
xor U18792 (N_18792,N_15015,N_16759);
nor U18793 (N_18793,N_15689,N_17864);
or U18794 (N_18794,N_16883,N_17885);
and U18795 (N_18795,N_15249,N_15302);
xnor U18796 (N_18796,N_15906,N_15018);
xnor U18797 (N_18797,N_16671,N_15500);
nand U18798 (N_18798,N_15471,N_16134);
and U18799 (N_18799,N_17198,N_16551);
nand U18800 (N_18800,N_17420,N_15120);
or U18801 (N_18801,N_16174,N_16477);
and U18802 (N_18802,N_15587,N_17773);
or U18803 (N_18803,N_15338,N_16916);
nor U18804 (N_18804,N_16762,N_17009);
nand U18805 (N_18805,N_15023,N_15968);
nand U18806 (N_18806,N_15882,N_15399);
xnor U18807 (N_18807,N_16576,N_15154);
or U18808 (N_18808,N_15475,N_16776);
xor U18809 (N_18809,N_16453,N_17349);
xnor U18810 (N_18810,N_16593,N_17896);
or U18811 (N_18811,N_17591,N_15187);
and U18812 (N_18812,N_15419,N_17105);
or U18813 (N_18813,N_17138,N_15030);
nand U18814 (N_18814,N_16177,N_17920);
or U18815 (N_18815,N_15647,N_17694);
and U18816 (N_18816,N_15664,N_17287);
or U18817 (N_18817,N_15201,N_17032);
xor U18818 (N_18818,N_17291,N_15985);
nor U18819 (N_18819,N_17868,N_16183);
and U18820 (N_18820,N_17168,N_15684);
or U18821 (N_18821,N_16460,N_17364);
and U18822 (N_18822,N_16565,N_16569);
or U18823 (N_18823,N_16104,N_17594);
nor U18824 (N_18824,N_15196,N_17867);
and U18825 (N_18825,N_16331,N_15983);
nand U18826 (N_18826,N_15013,N_16739);
nor U18827 (N_18827,N_15331,N_15192);
nand U18828 (N_18828,N_15451,N_16100);
nand U18829 (N_18829,N_17459,N_16702);
nor U18830 (N_18830,N_15627,N_15185);
xor U18831 (N_18831,N_15722,N_15280);
and U18832 (N_18832,N_17763,N_16698);
and U18833 (N_18833,N_17965,N_15642);
or U18834 (N_18834,N_16057,N_15894);
and U18835 (N_18835,N_15666,N_15448);
nand U18836 (N_18836,N_17071,N_17758);
nor U18837 (N_18837,N_15334,N_16092);
nor U18838 (N_18838,N_16680,N_17347);
or U18839 (N_18839,N_16469,N_15436);
nand U18840 (N_18840,N_17541,N_15091);
nor U18841 (N_18841,N_16582,N_17686);
and U18842 (N_18842,N_17742,N_17927);
or U18843 (N_18843,N_17436,N_17608);
nor U18844 (N_18844,N_16390,N_16010);
or U18845 (N_18845,N_17809,N_16677);
xnor U18846 (N_18846,N_15699,N_17660);
nand U18847 (N_18847,N_15428,N_15554);
and U18848 (N_18848,N_15274,N_16220);
and U18849 (N_18849,N_15359,N_15228);
nand U18850 (N_18850,N_16601,N_16736);
nor U18851 (N_18851,N_17041,N_17281);
nand U18852 (N_18852,N_16369,N_16403);
xnor U18853 (N_18853,N_16604,N_15095);
nand U18854 (N_18854,N_17848,N_15871);
nor U18855 (N_18855,N_16371,N_16204);
nor U18856 (N_18856,N_17108,N_17565);
nor U18857 (N_18857,N_16341,N_16853);
nand U18858 (N_18858,N_16505,N_17527);
nor U18859 (N_18859,N_15790,N_17906);
and U18860 (N_18860,N_17146,N_15158);
xnor U18861 (N_18861,N_17750,N_15863);
or U18862 (N_18862,N_15584,N_16732);
nor U18863 (N_18863,N_17556,N_16974);
xnor U18864 (N_18864,N_15556,N_17640);
and U18865 (N_18865,N_16849,N_17859);
or U18866 (N_18866,N_16627,N_15779);
nand U18867 (N_18867,N_15988,N_17244);
nand U18868 (N_18868,N_15660,N_16135);
xor U18869 (N_18869,N_15674,N_16721);
and U18870 (N_18870,N_17550,N_16873);
xor U18871 (N_18871,N_17014,N_17801);
or U18872 (N_18872,N_17307,N_16388);
nor U18873 (N_18873,N_17331,N_17471);
or U18874 (N_18874,N_16953,N_17907);
nand U18875 (N_18875,N_17228,N_16490);
xor U18876 (N_18876,N_16503,N_17113);
nand U18877 (N_18877,N_15654,N_15610);
nor U18878 (N_18878,N_16543,N_15136);
nor U18879 (N_18879,N_16451,N_16561);
and U18880 (N_18880,N_17956,N_15948);
or U18881 (N_18881,N_17873,N_15831);
nand U18882 (N_18882,N_15385,N_17130);
nor U18883 (N_18883,N_16326,N_17379);
xor U18884 (N_18884,N_16171,N_16156);
or U18885 (N_18885,N_15166,N_16125);
and U18886 (N_18886,N_17419,N_16206);
and U18887 (N_18887,N_16073,N_15220);
nand U18888 (N_18888,N_17351,N_16589);
xor U18889 (N_18889,N_16143,N_17195);
or U18890 (N_18890,N_15915,N_17208);
nor U18891 (N_18891,N_15935,N_15825);
and U18892 (N_18892,N_16571,N_15821);
xnor U18893 (N_18893,N_15953,N_15884);
nand U18894 (N_18894,N_15766,N_16898);
xnor U18895 (N_18895,N_16668,N_17776);
nor U18896 (N_18896,N_17993,N_17813);
xor U18897 (N_18897,N_17687,N_16474);
xor U18898 (N_18898,N_15174,N_15344);
or U18899 (N_18899,N_17469,N_17872);
nand U18900 (N_18900,N_15042,N_15038);
and U18901 (N_18901,N_15327,N_15257);
and U18902 (N_18902,N_16666,N_15369);
or U18903 (N_18903,N_15481,N_16645);
xor U18904 (N_18904,N_16712,N_15638);
xor U18905 (N_18905,N_16526,N_17816);
xor U18906 (N_18906,N_17698,N_16001);
nand U18907 (N_18907,N_15463,N_17819);
and U18908 (N_18908,N_16488,N_17889);
xnor U18909 (N_18909,N_17634,N_16623);
nand U18910 (N_18910,N_16415,N_16228);
nand U18911 (N_18911,N_16731,N_15562);
nand U18912 (N_18912,N_16639,N_15675);
xnor U18913 (N_18913,N_16594,N_16839);
and U18914 (N_18914,N_16890,N_15149);
nand U18915 (N_18915,N_17091,N_15944);
nor U18916 (N_18916,N_15712,N_16246);
or U18917 (N_18917,N_16422,N_17593);
and U18918 (N_18918,N_16472,N_15837);
or U18919 (N_18919,N_17280,N_15062);
nor U18920 (N_18920,N_16211,N_15743);
nor U18921 (N_18921,N_15996,N_17236);
nor U18922 (N_18922,N_16457,N_17242);
nand U18923 (N_18923,N_16382,N_15759);
nand U18924 (N_18924,N_15298,N_15838);
or U18925 (N_18925,N_17219,N_17538);
and U18926 (N_18926,N_16338,N_17987);
xor U18927 (N_18927,N_17288,N_16362);
nor U18928 (N_18928,N_17066,N_16370);
nand U18929 (N_18929,N_17371,N_16273);
and U18930 (N_18930,N_15407,N_16714);
nor U18931 (N_18931,N_15578,N_16699);
xnor U18932 (N_18932,N_15167,N_15374);
and U18933 (N_18933,N_17431,N_17890);
and U18934 (N_18934,N_15540,N_17798);
and U18935 (N_18935,N_17986,N_16245);
or U18936 (N_18936,N_16583,N_16706);
nor U18937 (N_18937,N_16471,N_17957);
or U18938 (N_18938,N_16439,N_17838);
or U18939 (N_18939,N_17899,N_15336);
xor U18940 (N_18940,N_16155,N_15750);
nand U18941 (N_18941,N_15892,N_15984);
xor U18942 (N_18942,N_16901,N_16483);
or U18943 (N_18943,N_15202,N_17974);
or U18944 (N_18944,N_17418,N_17894);
nor U18945 (N_18945,N_16310,N_17843);
xor U18946 (N_18946,N_16804,N_17161);
or U18947 (N_18947,N_16811,N_16820);
and U18948 (N_18948,N_15961,N_17301);
nor U18949 (N_18949,N_17409,N_15700);
and U18950 (N_18950,N_16658,N_17353);
or U18951 (N_18951,N_16418,N_17969);
and U18952 (N_18952,N_16969,N_17882);
nor U18953 (N_18953,N_17410,N_16434);
or U18954 (N_18954,N_16626,N_16318);
nand U18955 (N_18955,N_16629,N_15840);
xor U18956 (N_18956,N_16802,N_17328);
nand U18957 (N_18957,N_17700,N_16461);
nand U18958 (N_18958,N_17537,N_16251);
and U18959 (N_18959,N_16051,N_15549);
nand U18960 (N_18960,N_16930,N_15571);
and U18961 (N_18961,N_15259,N_15081);
and U18962 (N_18962,N_16176,N_16378);
or U18963 (N_18963,N_15010,N_15783);
and U18964 (N_18964,N_15006,N_15263);
or U18965 (N_18965,N_15686,N_15347);
and U18966 (N_18966,N_15213,N_16108);
nand U18967 (N_18967,N_15134,N_15388);
xor U18968 (N_18968,N_15078,N_16407);
or U18969 (N_18969,N_16069,N_17678);
xnor U18970 (N_18970,N_16061,N_17650);
xor U18971 (N_18971,N_17081,N_15781);
xnor U18972 (N_18972,N_16062,N_17990);
nand U18973 (N_18973,N_15776,N_17184);
nor U18974 (N_18974,N_16424,N_17627);
nand U18975 (N_18975,N_15455,N_17220);
and U18976 (N_18976,N_15367,N_17810);
nor U18977 (N_18977,N_16965,N_16188);
nor U18978 (N_18978,N_16578,N_16087);
nand U18979 (N_18979,N_15788,N_16967);
nand U18980 (N_18980,N_15814,N_16630);
nand U18981 (N_18981,N_17653,N_17317);
xor U18982 (N_18982,N_15972,N_16368);
nor U18983 (N_18983,N_17743,N_16292);
and U18984 (N_18984,N_17575,N_16408);
nor U18985 (N_18985,N_15342,N_16433);
nand U18986 (N_18986,N_16652,N_16829);
and U18987 (N_18987,N_17739,N_15887);
xnor U18988 (N_18988,N_16624,N_17582);
nand U18989 (N_18989,N_17378,N_16023);
or U18990 (N_18990,N_15769,N_17042);
or U18991 (N_18991,N_15987,N_15129);
xnor U18992 (N_18992,N_16306,N_15404);
xor U18993 (N_18993,N_16751,N_16272);
nor U18994 (N_18994,N_17295,N_17875);
and U18995 (N_18995,N_16847,N_17597);
nor U18996 (N_18996,N_17341,N_16676);
xor U18997 (N_18997,N_15890,N_16031);
nor U18998 (N_18998,N_17764,N_16054);
nor U18999 (N_18999,N_15426,N_16541);
or U19000 (N_19000,N_15485,N_16841);
xnor U19001 (N_19001,N_15629,N_15279);
or U19002 (N_19002,N_17002,N_16527);
and U19003 (N_19003,N_17480,N_16769);
nand U19004 (N_19004,N_15671,N_15965);
and U19005 (N_19005,N_15893,N_17756);
nor U19006 (N_19006,N_17737,N_15962);
xor U19007 (N_19007,N_16365,N_15118);
and U19008 (N_19008,N_17615,N_17050);
nand U19009 (N_19009,N_16381,N_16636);
or U19010 (N_19010,N_17346,N_17779);
and U19011 (N_19011,N_15156,N_15857);
xnor U19012 (N_19012,N_17072,N_15880);
xnor U19013 (N_19013,N_17426,N_16521);
and U19014 (N_19014,N_17796,N_17408);
nand U19015 (N_19015,N_17454,N_16986);
and U19016 (N_19016,N_17450,N_16611);
and U19017 (N_19017,N_17811,N_16504);
nand U19018 (N_19018,N_15650,N_16038);
and U19019 (N_19019,N_17970,N_15964);
nand U19020 (N_19020,N_15927,N_16950);
xor U19021 (N_19021,N_17525,N_16154);
and U19022 (N_19022,N_16473,N_15939);
xor U19023 (N_19023,N_16347,N_16446);
xnor U19024 (N_19024,N_17605,N_17702);
nand U19025 (N_19025,N_15969,N_15438);
nor U19026 (N_19026,N_15181,N_15241);
and U19027 (N_19027,N_17299,N_16633);
nor U19028 (N_19028,N_15487,N_17664);
nand U19029 (N_19029,N_15235,N_16907);
xor U19030 (N_19030,N_16808,N_15875);
and U19031 (N_19031,N_16866,N_16492);
and U19032 (N_19032,N_15420,N_17470);
and U19033 (N_19033,N_17655,N_16939);
xnor U19034 (N_19034,N_17771,N_17191);
and U19035 (N_19035,N_15976,N_16353);
or U19036 (N_19036,N_15272,N_16512);
nor U19037 (N_19037,N_15260,N_16517);
xor U19038 (N_19038,N_16660,N_16227);
xnor U19039 (N_19039,N_16690,N_15974);
nor U19040 (N_19040,N_16411,N_16764);
and U19041 (N_19041,N_17587,N_17256);
and U19042 (N_19042,N_15242,N_16707);
nand U19043 (N_19043,N_15147,N_15758);
nor U19044 (N_19044,N_16144,N_15150);
and U19045 (N_19045,N_15265,N_15160);
nor U19046 (N_19046,N_15721,N_17265);
and U19047 (N_19047,N_15942,N_15945);
xor U19048 (N_19048,N_17221,N_15329);
or U19049 (N_19049,N_15450,N_17622);
xnor U19050 (N_19050,N_17972,N_15532);
nor U19051 (N_19051,N_17117,N_16375);
or U19052 (N_19052,N_15116,N_17921);
or U19053 (N_19053,N_16187,N_15313);
nor U19054 (N_19054,N_15874,N_15208);
and U19055 (N_19055,N_16363,N_17693);
nor U19056 (N_19056,N_15723,N_16169);
and U19057 (N_19057,N_17599,N_17976);
or U19058 (N_19058,N_17871,N_16392);
xor U19059 (N_19059,N_16080,N_16800);
and U19060 (N_19060,N_17298,N_17948);
nor U19061 (N_19061,N_17484,N_15255);
xnor U19062 (N_19062,N_16840,N_17855);
or U19063 (N_19063,N_17089,N_15483);
nand U19064 (N_19064,N_16855,N_15956);
and U19065 (N_19065,N_15024,N_15063);
and U19066 (N_19066,N_16757,N_15476);
and U19067 (N_19067,N_16172,N_15390);
or U19068 (N_19068,N_17403,N_16264);
nand U19069 (N_19069,N_16859,N_17562);
or U19070 (N_19070,N_16982,N_15846);
and U19071 (N_19071,N_16017,N_16084);
or U19072 (N_19072,N_16549,N_15423);
or U19073 (N_19073,N_15862,N_17229);
xnor U19074 (N_19074,N_16244,N_15266);
or U19075 (N_19075,N_16993,N_17356);
and U19076 (N_19076,N_16845,N_15180);
or U19077 (N_19077,N_17511,N_15184);
xnor U19078 (N_19078,N_17585,N_15458);
or U19079 (N_19079,N_15786,N_17589);
nand U19080 (N_19080,N_16275,N_16336);
or U19081 (N_19081,N_15324,N_17497);
xnor U19082 (N_19082,N_15667,N_16298);
xor U19083 (N_19083,N_15765,N_16450);
and U19084 (N_19084,N_16603,N_17930);
nand U19085 (N_19085,N_15012,N_17571);
nand U19086 (N_19086,N_15218,N_15211);
nand U19087 (N_19087,N_16089,N_17831);
xnor U19088 (N_19088,N_16795,N_16534);
and U19089 (N_19089,N_16886,N_17780);
nand U19090 (N_19090,N_15757,N_15016);
nor U19091 (N_19091,N_16110,N_15705);
nand U19092 (N_19092,N_15827,N_16286);
nor U19093 (N_19093,N_17553,N_17145);
nand U19094 (N_19094,N_16239,N_15477);
nor U19095 (N_19095,N_17769,N_17186);
xnor U19096 (N_19096,N_15425,N_16733);
xor U19097 (N_19097,N_15937,N_15586);
nor U19098 (N_19098,N_17792,N_17035);
nor U19099 (N_19099,N_15683,N_15912);
and U19100 (N_19100,N_17049,N_15581);
nand U19101 (N_19101,N_17485,N_16557);
nand U19102 (N_19102,N_16920,N_17054);
and U19103 (N_19103,N_16738,N_17690);
nand U19104 (N_19104,N_15157,N_16799);
nor U19105 (N_19105,N_16868,N_15801);
or U19106 (N_19106,N_16628,N_17825);
xnor U19107 (N_19107,N_17474,N_17080);
or U19108 (N_19108,N_17567,N_15297);
nor U19109 (N_19109,N_16895,N_17276);
or U19110 (N_19110,N_16037,N_15017);
nand U19111 (N_19111,N_15528,N_16146);
or U19112 (N_19112,N_16743,N_17245);
nor U19113 (N_19113,N_17082,N_15522);
xnor U19114 (N_19114,N_15495,N_16072);
nor U19115 (N_19115,N_17201,N_15744);
and U19116 (N_19116,N_15381,N_16990);
and U19117 (N_19117,N_16032,N_15659);
nand U19118 (N_19118,N_16801,N_17959);
nand U19119 (N_19119,N_15041,N_15822);
and U19120 (N_19120,N_16379,N_16192);
xor U19121 (N_19121,N_15033,N_17270);
or U19122 (N_19122,N_17551,N_16700);
or U19123 (N_19123,N_16684,N_15361);
xnor U19124 (N_19124,N_17614,N_15079);
xor U19125 (N_19125,N_16711,N_16735);
nor U19126 (N_19126,N_16253,N_16194);
or U19127 (N_19127,N_16518,N_15127);
or U19128 (N_19128,N_16064,N_17160);
and U19129 (N_19129,N_17127,N_16395);
nor U19130 (N_19130,N_17057,N_17671);
or U19131 (N_19131,N_17832,N_16287);
or U19132 (N_19132,N_17719,N_16910);
nor U19133 (N_19133,N_17518,N_17101);
or U19134 (N_19134,N_16941,N_16979);
xor U19135 (N_19135,N_15713,N_17277);
and U19136 (N_19136,N_17850,N_17688);
nor U19137 (N_19137,N_15946,N_15637);
or U19138 (N_19138,N_16283,N_17045);
or U19139 (N_19139,N_16191,N_15251);
nand U19140 (N_19140,N_17626,N_15704);
nand U19141 (N_19141,N_16860,N_15317);
or U19142 (N_19142,N_15955,N_16096);
and U19143 (N_19143,N_17422,N_17782);
xnor U19144 (N_19144,N_17327,N_17789);
or U19145 (N_19145,N_17102,N_17202);
nor U19146 (N_19146,N_15978,N_15029);
and U19147 (N_19147,N_15543,N_15406);
or U19148 (N_19148,N_17919,N_16508);
and U19149 (N_19149,N_16775,N_16632);
or U19150 (N_19150,N_15997,N_17583);
or U19151 (N_19151,N_17266,N_15496);
or U19152 (N_19152,N_16013,N_17596);
nor U19153 (N_19153,N_17733,N_17543);
nand U19154 (N_19154,N_15061,N_16912);
or U19155 (N_19155,N_16718,N_16921);
nor U19156 (N_19156,N_16758,N_15092);
and U19157 (N_19157,N_17120,N_16349);
or U19158 (N_19158,N_16807,N_15539);
xor U19159 (N_19159,N_16207,N_15855);
xor U19160 (N_19160,N_17224,N_16650);
xnor U19161 (N_19161,N_17211,N_16116);
nand U19162 (N_19162,N_17246,N_15058);
nand U19163 (N_19163,N_15736,N_16919);
nor U19164 (N_19164,N_15349,N_15834);
xnor U19165 (N_19165,N_15818,N_15594);
nor U19166 (N_19166,N_15161,N_16498);
nand U19167 (N_19167,N_15314,N_16500);
nor U19168 (N_19168,N_15103,N_16115);
xor U19169 (N_19169,N_17306,N_16532);
nand U19170 (N_19170,N_17092,N_16942);
xor U19171 (N_19171,N_16963,N_15563);
and U19172 (N_19172,N_15568,N_16234);
and U19173 (N_19173,N_16430,N_15682);
or U19174 (N_19174,N_17368,N_16319);
or U19175 (N_19175,N_16285,N_16041);
or U19176 (N_19176,N_16763,N_16325);
or U19177 (N_19177,N_15856,N_17643);
and U19178 (N_19178,N_16835,N_17703);
nand U19179 (N_19179,N_17942,N_16951);
nand U19180 (N_19180,N_17914,N_17836);
or U19181 (N_19181,N_17999,N_17382);
xor U19182 (N_19182,N_15261,N_15630);
or U19183 (N_19183,N_15994,N_16223);
nor U19184 (N_19184,N_15934,N_16022);
nand U19185 (N_19185,N_17142,N_16983);
nand U19186 (N_19186,N_15183,N_17348);
or U19187 (N_19187,N_16885,N_17852);
or U19188 (N_19188,N_15588,N_15986);
xor U19189 (N_19189,N_17949,N_15910);
nor U19190 (N_19190,N_15034,N_16556);
nand U19191 (N_19191,N_15860,N_15665);
nor U19192 (N_19192,N_16139,N_15695);
nand U19193 (N_19193,N_15709,N_17226);
or U19194 (N_19194,N_16402,N_16131);
nor U19195 (N_19195,N_16817,N_16978);
nor U19196 (N_19196,N_17573,N_15852);
and U19197 (N_19197,N_15680,N_16708);
or U19198 (N_19198,N_17177,N_17124);
nor U19199 (N_19199,N_15751,N_16059);
or U19200 (N_19200,N_17493,N_17600);
nor U19201 (N_19201,N_17837,N_16516);
and U19202 (N_19202,N_16806,N_17441);
nand U19203 (N_19203,N_15049,N_16337);
xor U19204 (N_19204,N_17736,N_15316);
or U19205 (N_19205,N_16545,N_16398);
or U19206 (N_19206,N_15904,N_15264);
or U19207 (N_19207,N_16210,N_17561);
and U19208 (N_19208,N_17136,N_15764);
and U19209 (N_19209,N_15523,N_15368);
xnor U19210 (N_19210,N_17510,N_15389);
and U19211 (N_19211,N_16709,N_16783);
nor U19212 (N_19212,N_15753,N_15973);
and U19213 (N_19213,N_17673,N_16198);
and U19214 (N_19214,N_16619,N_17844);
xnor U19215 (N_19215,N_16113,N_17966);
nand U19216 (N_19216,N_17827,N_17521);
nand U19217 (N_19217,N_16208,N_16254);
or U19218 (N_19218,N_17799,N_17479);
nand U19219 (N_19219,N_16908,N_17951);
nor U19220 (N_19220,N_15693,N_17052);
nand U19221 (N_19221,N_15125,N_15730);
or U19222 (N_19222,N_17399,N_15194);
and U19223 (N_19223,N_17996,N_16692);
or U19224 (N_19224,N_16725,N_16655);
xnor U19225 (N_19225,N_15284,N_16012);
or U19226 (N_19226,N_16152,N_17929);
nand U19227 (N_19227,N_17952,N_15618);
xor U19228 (N_19228,N_16491,N_15916);
xor U19229 (N_19229,N_17777,N_17111);
nor U19230 (N_19230,N_15612,N_17489);
and U19231 (N_19231,N_17452,N_17037);
nor U19232 (N_19232,N_16613,N_17013);
xnor U19233 (N_19233,N_17628,N_16597);
xor U19234 (N_19234,N_17569,N_16126);
and U19235 (N_19235,N_16869,N_16499);
and U19236 (N_19236,N_15706,N_17803);
nand U19237 (N_19237,N_17880,N_17488);
or U19238 (N_19238,N_17255,N_17086);
nand U19239 (N_19239,N_17761,N_16046);
xor U19240 (N_19240,N_15341,N_15090);
and U19241 (N_19241,N_16098,N_16265);
or U19242 (N_19242,N_17467,N_15210);
nor U19243 (N_19243,N_16519,N_16480);
nand U19244 (N_19244,N_16971,N_16021);
and U19245 (N_19245,N_16661,N_16423);
or U19246 (N_19246,N_17360,N_17336);
nor U19247 (N_19247,N_17738,N_15925);
and U19248 (N_19248,N_17712,N_15861);
nand U19249 (N_19249,N_15443,N_15719);
or U19250 (N_19250,N_17717,N_16235);
nor U19251 (N_19251,N_16487,N_16293);
nor U19252 (N_19252,N_16647,N_17904);
or U19253 (N_19253,N_15216,N_17008);
nand U19254 (N_19254,N_15848,N_17458);
or U19255 (N_19255,N_15993,N_17530);
xor U19256 (N_19256,N_16742,N_16688);
xor U19257 (N_19257,N_15137,N_17383);
nor U19258 (N_19258,N_15044,N_15432);
or U19259 (N_19259,N_17598,N_16962);
nand U19260 (N_19260,N_17849,N_17247);
and U19261 (N_19261,N_17447,N_16437);
and U19262 (N_19262,N_15745,N_16321);
or U19263 (N_19263,N_15200,N_16787);
xnor U19264 (N_19264,N_15377,N_16162);
nand U19265 (N_19265,N_15339,N_15252);
nand U19266 (N_19266,N_15954,N_15503);
nor U19267 (N_19267,N_15052,N_16093);
and U19268 (N_19268,N_16609,N_16350);
nor U19269 (N_19269,N_16302,N_16340);
or U19270 (N_19270,N_16329,N_16891);
nand U19271 (N_19271,N_17841,N_15085);
or U19272 (N_19272,N_15097,N_17557);
nor U19273 (N_19273,N_15186,N_15898);
nand U19274 (N_19274,N_16199,N_15291);
nand U19275 (N_19275,N_17768,N_15352);
and U19276 (N_19276,N_15760,N_16641);
nand U19277 (N_19277,N_17320,N_17369);
nand U19278 (N_19278,N_16066,N_17933);
xor U19279 (N_19279,N_17078,N_15741);
and U19280 (N_19280,N_16564,N_17715);
xnor U19281 (N_19281,N_17578,N_15278);
nor U19282 (N_19282,N_16987,N_16083);
nor U19283 (N_19283,N_17473,N_17725);
xnor U19284 (N_19284,N_17989,N_17038);
or U19285 (N_19285,N_15519,N_15304);
and U19286 (N_19286,N_15809,N_16218);
nor U19287 (N_19287,N_15943,N_15724);
xor U19288 (N_19288,N_17824,N_16832);
and U19289 (N_19289,N_15731,N_15591);
or U19290 (N_19290,N_15891,N_17475);
xnor U19291 (N_19291,N_17595,N_16892);
and U19292 (N_19292,N_16147,N_15839);
and U19293 (N_19293,N_16925,N_17775);
and U19294 (N_19294,N_17152,N_16036);
nand U19295 (N_19295,N_15057,N_16843);
xor U19296 (N_19296,N_17150,N_17496);
or U19297 (N_19297,N_16640,N_16282);
xnor U19298 (N_19298,N_16443,N_15084);
nor U19299 (N_19299,N_17132,N_16140);
xnor U19300 (N_19300,N_15914,N_16355);
nor U19301 (N_19301,N_17154,N_15315);
nor U19302 (N_19302,N_16486,N_16580);
and U19303 (N_19303,N_17515,N_16562);
nor U19304 (N_19304,N_15102,N_15020);
xor U19305 (N_19305,N_16307,N_17568);
and U19306 (N_19306,N_17950,N_17701);
and U19307 (N_19307,N_15189,N_15595);
xnor U19308 (N_19308,N_17209,N_15534);
nor U19309 (N_19309,N_16697,N_15415);
xnor U19310 (N_19310,N_15287,N_15345);
and U19311 (N_19311,N_16948,N_15478);
xnor U19312 (N_19312,N_17088,N_17638);
or U19313 (N_19313,N_16674,N_16271);
and U19314 (N_19314,N_15433,N_15747);
xnor U19315 (N_19315,N_17460,N_17645);
or U19316 (N_19316,N_16719,N_15205);
xor U19317 (N_19317,N_15635,N_17539);
xnor U19318 (N_19318,N_15392,N_16079);
nand U19319 (N_19319,N_16625,N_17385);
xnor U19320 (N_19320,N_15267,N_15802);
and U19321 (N_19321,N_15244,N_15832);
nand U19322 (N_19322,N_15351,N_15817);
or U19323 (N_19323,N_17272,N_15040);
xnor U19324 (N_19324,N_15394,N_15742);
nor U19325 (N_19325,N_17839,N_17030);
nand U19326 (N_19326,N_15579,N_17492);
or U19327 (N_19327,N_16867,N_15672);
nand U19328 (N_19328,N_15268,N_15440);
nor U19329 (N_19329,N_17912,N_17167);
xnor U19330 (N_19330,N_17659,N_15224);
nand U19331 (N_19331,N_16756,N_17381);
nor U19332 (N_19332,N_15497,N_17501);
xor U19333 (N_19333,N_16932,N_16165);
xor U19334 (N_19334,N_15656,N_15354);
xnor U19335 (N_19335,N_17520,N_16068);
and U19336 (N_19336,N_16573,N_16462);
and U19337 (N_19337,N_16765,N_17402);
nor U19338 (N_19338,N_17258,N_15735);
xnor U19339 (N_19339,N_15872,N_15710);
xor U19340 (N_19340,N_15243,N_15980);
nand U19341 (N_19341,N_16324,N_16960);
nor U19342 (N_19342,N_17393,N_16291);
or U19343 (N_19343,N_15634,N_15227);
and U19344 (N_19344,N_17309,N_16745);
nor U19345 (N_19345,N_17337,N_17941);
or U19346 (N_19346,N_15648,N_17326);
nor U19347 (N_19347,N_17345,N_17194);
xor U19348 (N_19348,N_17011,N_16746);
nor U19349 (N_19349,N_15320,N_16497);
xor U19350 (N_19350,N_16958,N_17273);
nor U19351 (N_19351,N_17616,N_15564);
nand U19352 (N_19352,N_17338,N_17190);
nand U19353 (N_19353,N_16455,N_16599);
nand U19354 (N_19354,N_15847,N_16926);
or U19355 (N_19355,N_15256,N_17784);
and U19356 (N_19356,N_17862,N_17311);
or U19357 (N_19357,N_15238,N_15752);
or U19358 (N_19358,N_15408,N_15155);
nand U19359 (N_19359,N_16429,N_15019);
nor U19360 (N_19360,N_15467,N_15162);
nand U19361 (N_19361,N_17233,N_16231);
or U19362 (N_19362,N_15620,N_15529);
nand U19363 (N_19363,N_17392,N_16610);
nand U19364 (N_19364,N_16067,N_15739);
nand U19365 (N_19365,N_15053,N_15356);
nor U19366 (N_19366,N_17312,N_15828);
and U19367 (N_19367,N_17238,N_15661);
or U19368 (N_19368,N_15488,N_16221);
and U19369 (N_19369,N_17074,N_16928);
and U19370 (N_19370,N_15104,N_15836);
nand U19371 (N_19371,N_17374,N_15059);
nor U19372 (N_19372,N_15323,N_16784);
nor U19373 (N_19373,N_16367,N_15025);
nand U19374 (N_19374,N_15142,N_15504);
nor U19375 (N_19375,N_15121,N_15900);
xor U19376 (N_19376,N_16838,N_17835);
nand U19377 (N_19377,N_17910,N_15881);
nand U19378 (N_19378,N_15678,N_15707);
xor U19379 (N_19379,N_17239,N_15123);
nor U19380 (N_19380,N_16997,N_16459);
or U19381 (N_19381,N_16070,N_16373);
nand U19382 (N_19382,N_16201,N_17319);
xnor U19383 (N_19383,N_17116,N_15122);
nand U19384 (N_19384,N_15566,N_17901);
nor U19385 (N_19385,N_16833,N_15226);
or U19386 (N_19386,N_15036,N_17564);
nor U19387 (N_19387,N_16566,N_15605);
xnor U19388 (N_19388,N_17529,N_15140);
xnor U19389 (N_19389,N_17984,N_17016);
or U19390 (N_19390,N_17677,N_15382);
nor U19391 (N_19391,N_16918,N_17400);
and U19392 (N_19392,N_16798,N_15878);
or U19393 (N_19393,N_16412,N_17611);
and U19394 (N_19394,N_15663,N_15096);
nor U19395 (N_19395,N_17757,N_17053);
or U19396 (N_19396,N_16019,N_15170);
or U19397 (N_19397,N_17546,N_17641);
or U19398 (N_19398,N_15979,N_15815);
nand U19399 (N_19399,N_16747,N_15538);
nand U19400 (N_19400,N_17584,N_17324);
or U19401 (N_19401,N_17325,N_17143);
nor U19402 (N_19402,N_16550,N_16620);
nor U19403 (N_19403,N_16058,N_15645);
xor U19404 (N_19404,N_16771,N_15560);
and U19405 (N_19405,N_16288,N_17924);
xnor U19406 (N_19406,N_16529,N_16419);
xor U19407 (N_19407,N_17333,N_15989);
xor U19408 (N_19408,N_16196,N_16606);
nor U19409 (N_19409,N_16515,N_16539);
xor U19410 (N_19410,N_16458,N_16522);
nand U19411 (N_19411,N_16295,N_15312);
nand U19412 (N_19412,N_15207,N_15335);
and U19413 (N_19413,N_17786,N_17649);
nor U19414 (N_19414,N_15772,N_16996);
xnor U19415 (N_19415,N_16421,N_16857);
or U19416 (N_19416,N_16075,N_16989);
and U19417 (N_19417,N_15569,N_16929);
nand U19418 (N_19418,N_15348,N_16088);
and U19419 (N_19419,N_17814,N_16212);
and U19420 (N_19420,N_15411,N_15214);
nand U19421 (N_19421,N_16752,N_15159);
or U19422 (N_19422,N_17129,N_15513);
nor U19423 (N_19423,N_15479,N_16033);
nand U19424 (N_19424,N_17058,N_17960);
nor U19425 (N_19425,N_17716,N_15191);
and U19426 (N_19426,N_15115,N_15676);
and U19427 (N_19427,N_15460,N_16003);
xnor U19428 (N_19428,N_17549,N_16274);
and U19429 (N_19429,N_17199,N_15901);
or U19430 (N_19430,N_17619,N_17332);
and U19431 (N_19431,N_16127,N_15895);
nand U19432 (N_19432,N_17973,N_17504);
nand U19433 (N_19433,N_15333,N_15075);
and U19434 (N_19434,N_17061,N_16766);
nor U19435 (N_19435,N_15725,N_17355);
nand U19436 (N_19436,N_17507,N_16651);
or U19437 (N_19437,N_15520,N_15069);
or U19438 (N_19438,N_16905,N_16130);
or U19439 (N_19439,N_15054,N_16975);
and U19440 (N_19440,N_15146,N_15596);
nand U19441 (N_19441,N_16741,N_16615);
nor U19442 (N_19442,N_16276,N_16900);
nand U19443 (N_19443,N_17665,N_17991);
nor U19444 (N_19444,N_17944,N_15322);
xnor U19445 (N_19445,N_16701,N_17781);
xor U19446 (N_19446,N_17218,N_17623);
xnor U19447 (N_19447,N_15603,N_16724);
nor U19448 (N_19448,N_16616,N_16132);
or U19449 (N_19449,N_16360,N_17601);
and U19450 (N_19450,N_15229,N_17730);
xor U19451 (N_19451,N_17581,N_16984);
nand U19452 (N_19452,N_17435,N_16836);
nor U19453 (N_19453,N_17051,N_17656);
xor U19454 (N_19454,N_15431,N_15326);
or U19455 (N_19455,N_16203,N_17820);
xnor U19456 (N_19456,N_15604,N_16638);
nor U19457 (N_19457,N_17866,N_16322);
xnor U19458 (N_19458,N_15107,N_15073);
and U19459 (N_19459,N_15681,N_15021);
or U19460 (N_19460,N_16357,N_15918);
nand U19461 (N_19461,N_15922,N_15444);
nand U19462 (N_19462,N_17579,N_17517);
or U19463 (N_19463,N_15702,N_17992);
xnor U19464 (N_19464,N_16074,N_16358);
nand U19465 (N_19465,N_15561,N_17158);
xor U19466 (N_19466,N_17023,N_17329);
nand U19467 (N_19467,N_17119,N_15550);
or U19468 (N_19468,N_16681,N_15789);
xor U19469 (N_19469,N_16862,N_17604);
xor U19470 (N_19470,N_17093,N_16279);
xnor U19471 (N_19471,N_15792,N_15262);
nor U19472 (N_19472,N_16705,N_17157);
or U19473 (N_19473,N_15452,N_15355);
nand U19474 (N_19474,N_17148,N_17423);
nor U19475 (N_19475,N_15527,N_15453);
xnor U19476 (N_19476,N_17230,N_15748);
and U19477 (N_19477,N_17636,N_15000);
or U19478 (N_19478,N_16815,N_17713);
nand U19479 (N_19479,N_17405,N_16416);
nor U19480 (N_19480,N_17840,N_15804);
xnor U19481 (N_19481,N_17322,N_16339);
or U19482 (N_19482,N_17877,N_17396);
nand U19483 (N_19483,N_16142,N_15920);
nor U19484 (N_19484,N_15577,N_17060);
or U19485 (N_19485,N_17079,N_15866);
or U19486 (N_19486,N_17528,N_15854);
nor U19487 (N_19487,N_16401,N_17394);
nand U19488 (N_19488,N_17887,N_17516);
and U19489 (N_19489,N_15376,N_16406);
xnor U19490 (N_19490,N_16007,N_17354);
and U19491 (N_19491,N_17928,N_17225);
nor U19492 (N_19492,N_17446,N_16717);
nor U19493 (N_19493,N_17413,N_17943);
xnor U19494 (N_19494,N_16780,N_15358);
xor U19495 (N_19495,N_16266,N_16250);
and U19496 (N_19496,N_16361,N_17163);
xor U19497 (N_19497,N_15435,N_15353);
nand U19498 (N_19498,N_16489,N_17606);
or U19499 (N_19499,N_16303,N_17851);
nand U19500 (N_19500,N_15190,N_17258);
nor U19501 (N_19501,N_17820,N_16206);
xor U19502 (N_19502,N_15609,N_17700);
nand U19503 (N_19503,N_17217,N_17066);
xnor U19504 (N_19504,N_16534,N_15185);
nand U19505 (N_19505,N_17473,N_17259);
nand U19506 (N_19506,N_15277,N_17861);
xor U19507 (N_19507,N_15166,N_17695);
nand U19508 (N_19508,N_17759,N_17891);
nor U19509 (N_19509,N_17667,N_16428);
nand U19510 (N_19510,N_17680,N_17750);
or U19511 (N_19511,N_16184,N_16012);
or U19512 (N_19512,N_15597,N_17796);
nand U19513 (N_19513,N_17918,N_17910);
or U19514 (N_19514,N_15864,N_17357);
nor U19515 (N_19515,N_16395,N_15662);
and U19516 (N_19516,N_16744,N_16196);
nand U19517 (N_19517,N_15220,N_17628);
and U19518 (N_19518,N_15917,N_16855);
nand U19519 (N_19519,N_16048,N_16537);
nor U19520 (N_19520,N_17504,N_16455);
nor U19521 (N_19521,N_16838,N_15760);
and U19522 (N_19522,N_17435,N_16556);
and U19523 (N_19523,N_16410,N_15707);
nand U19524 (N_19524,N_17417,N_17291);
or U19525 (N_19525,N_17595,N_17152);
nand U19526 (N_19526,N_17707,N_15058);
nor U19527 (N_19527,N_15269,N_16668);
or U19528 (N_19528,N_16150,N_16449);
or U19529 (N_19529,N_16381,N_16485);
xor U19530 (N_19530,N_16117,N_17264);
nand U19531 (N_19531,N_17330,N_15932);
xor U19532 (N_19532,N_17736,N_17825);
or U19533 (N_19533,N_15215,N_17185);
and U19534 (N_19534,N_15857,N_16507);
nor U19535 (N_19535,N_16620,N_16659);
xor U19536 (N_19536,N_16578,N_15213);
nand U19537 (N_19537,N_15845,N_16034);
nor U19538 (N_19538,N_17368,N_15367);
nor U19539 (N_19539,N_16890,N_16793);
xor U19540 (N_19540,N_17182,N_15830);
xnor U19541 (N_19541,N_17791,N_16025);
nor U19542 (N_19542,N_17359,N_15545);
and U19543 (N_19543,N_16555,N_17081);
nor U19544 (N_19544,N_16634,N_16258);
xor U19545 (N_19545,N_15806,N_15608);
xor U19546 (N_19546,N_17626,N_16431);
nand U19547 (N_19547,N_17802,N_17423);
and U19548 (N_19548,N_17068,N_17893);
and U19549 (N_19549,N_16130,N_15522);
xor U19550 (N_19550,N_17154,N_17467);
nor U19551 (N_19551,N_17378,N_17282);
xnor U19552 (N_19552,N_15261,N_17400);
nand U19553 (N_19553,N_16373,N_15915);
and U19554 (N_19554,N_17945,N_17972);
nand U19555 (N_19555,N_15941,N_17958);
nor U19556 (N_19556,N_16801,N_15188);
or U19557 (N_19557,N_16147,N_15201);
or U19558 (N_19558,N_16466,N_16564);
nand U19559 (N_19559,N_16257,N_16002);
nand U19560 (N_19560,N_17963,N_16453);
nand U19561 (N_19561,N_15950,N_16408);
or U19562 (N_19562,N_15990,N_16178);
nor U19563 (N_19563,N_16315,N_16287);
and U19564 (N_19564,N_17015,N_15633);
or U19565 (N_19565,N_15012,N_17393);
nand U19566 (N_19566,N_17363,N_17308);
and U19567 (N_19567,N_16796,N_15234);
and U19568 (N_19568,N_16350,N_15058);
nor U19569 (N_19569,N_16292,N_15267);
and U19570 (N_19570,N_16040,N_15740);
xor U19571 (N_19571,N_17050,N_17839);
or U19572 (N_19572,N_15591,N_15340);
nand U19573 (N_19573,N_17645,N_15955);
nor U19574 (N_19574,N_16086,N_15671);
and U19575 (N_19575,N_16247,N_16016);
and U19576 (N_19576,N_16544,N_15780);
or U19577 (N_19577,N_16188,N_17322);
nor U19578 (N_19578,N_16976,N_15880);
or U19579 (N_19579,N_16895,N_16555);
nand U19580 (N_19580,N_17822,N_16288);
and U19581 (N_19581,N_15315,N_16831);
or U19582 (N_19582,N_17222,N_15419);
nor U19583 (N_19583,N_15251,N_17061);
or U19584 (N_19584,N_15292,N_15033);
nor U19585 (N_19585,N_16034,N_16663);
or U19586 (N_19586,N_16163,N_15953);
nand U19587 (N_19587,N_16261,N_15796);
xnor U19588 (N_19588,N_15053,N_16258);
nand U19589 (N_19589,N_16891,N_17305);
nor U19590 (N_19590,N_17802,N_17396);
or U19591 (N_19591,N_17289,N_16822);
nand U19592 (N_19592,N_16693,N_17919);
nor U19593 (N_19593,N_17596,N_17450);
xnor U19594 (N_19594,N_17990,N_15903);
xor U19595 (N_19595,N_17394,N_15431);
nand U19596 (N_19596,N_15447,N_17089);
or U19597 (N_19597,N_16305,N_17409);
and U19598 (N_19598,N_15877,N_17412);
or U19599 (N_19599,N_15210,N_17828);
xnor U19600 (N_19600,N_16554,N_16714);
and U19601 (N_19601,N_15723,N_15340);
nor U19602 (N_19602,N_16454,N_15382);
and U19603 (N_19603,N_15810,N_16475);
xor U19604 (N_19604,N_17762,N_15186);
nand U19605 (N_19605,N_17886,N_17573);
nand U19606 (N_19606,N_16765,N_16020);
or U19607 (N_19607,N_15177,N_16816);
or U19608 (N_19608,N_16911,N_15420);
or U19609 (N_19609,N_17952,N_17140);
and U19610 (N_19610,N_16437,N_16267);
and U19611 (N_19611,N_15677,N_16959);
or U19612 (N_19612,N_16305,N_15767);
xor U19613 (N_19613,N_16044,N_17201);
xor U19614 (N_19614,N_15788,N_17597);
and U19615 (N_19615,N_15176,N_17961);
nor U19616 (N_19616,N_16708,N_15407);
or U19617 (N_19617,N_16292,N_15114);
or U19618 (N_19618,N_17087,N_16279);
nor U19619 (N_19619,N_15824,N_15622);
and U19620 (N_19620,N_17880,N_16734);
nand U19621 (N_19621,N_16699,N_17405);
and U19622 (N_19622,N_17455,N_16882);
nor U19623 (N_19623,N_17747,N_15415);
or U19624 (N_19624,N_15602,N_17429);
xor U19625 (N_19625,N_17520,N_15525);
or U19626 (N_19626,N_15360,N_17360);
xor U19627 (N_19627,N_17779,N_15297);
nor U19628 (N_19628,N_17590,N_15458);
xor U19629 (N_19629,N_16337,N_16270);
and U19630 (N_19630,N_17986,N_15318);
and U19631 (N_19631,N_17270,N_16149);
nand U19632 (N_19632,N_15447,N_16433);
xnor U19633 (N_19633,N_16255,N_17487);
nand U19634 (N_19634,N_17767,N_16654);
xnor U19635 (N_19635,N_16848,N_15374);
nand U19636 (N_19636,N_16731,N_15831);
nand U19637 (N_19637,N_16468,N_15505);
or U19638 (N_19638,N_17875,N_16632);
xor U19639 (N_19639,N_16891,N_16503);
and U19640 (N_19640,N_17158,N_16887);
or U19641 (N_19641,N_17232,N_15091);
and U19642 (N_19642,N_16870,N_15275);
xnor U19643 (N_19643,N_15579,N_17449);
or U19644 (N_19644,N_17120,N_15548);
xnor U19645 (N_19645,N_17243,N_15360);
nand U19646 (N_19646,N_15058,N_16040);
xnor U19647 (N_19647,N_17436,N_17780);
and U19648 (N_19648,N_15535,N_17095);
nor U19649 (N_19649,N_17256,N_15977);
xnor U19650 (N_19650,N_15248,N_16416);
nand U19651 (N_19651,N_17359,N_16244);
and U19652 (N_19652,N_16720,N_17446);
and U19653 (N_19653,N_17251,N_16381);
and U19654 (N_19654,N_17990,N_15827);
xnor U19655 (N_19655,N_17907,N_17993);
and U19656 (N_19656,N_15949,N_17362);
and U19657 (N_19657,N_16218,N_17705);
and U19658 (N_19658,N_15231,N_17470);
or U19659 (N_19659,N_17841,N_15048);
nand U19660 (N_19660,N_16294,N_16642);
xnor U19661 (N_19661,N_16312,N_15881);
and U19662 (N_19662,N_15103,N_17774);
and U19663 (N_19663,N_16753,N_17490);
and U19664 (N_19664,N_17189,N_15199);
or U19665 (N_19665,N_17368,N_15025);
nand U19666 (N_19666,N_15227,N_15493);
and U19667 (N_19667,N_17375,N_16406);
xor U19668 (N_19668,N_16185,N_17772);
or U19669 (N_19669,N_15765,N_17401);
nor U19670 (N_19670,N_16957,N_17868);
nor U19671 (N_19671,N_16761,N_17108);
xnor U19672 (N_19672,N_16805,N_17551);
or U19673 (N_19673,N_15474,N_17369);
or U19674 (N_19674,N_15084,N_16161);
nor U19675 (N_19675,N_17220,N_17713);
xor U19676 (N_19676,N_15318,N_16524);
nand U19677 (N_19677,N_15453,N_15661);
nand U19678 (N_19678,N_15542,N_17406);
nand U19679 (N_19679,N_16074,N_15984);
xnor U19680 (N_19680,N_17528,N_16688);
nand U19681 (N_19681,N_17781,N_15738);
and U19682 (N_19682,N_17984,N_17018);
nand U19683 (N_19683,N_17382,N_16981);
nor U19684 (N_19684,N_16965,N_16072);
and U19685 (N_19685,N_16930,N_17982);
and U19686 (N_19686,N_15509,N_17746);
xor U19687 (N_19687,N_15861,N_16474);
xnor U19688 (N_19688,N_17133,N_15239);
xnor U19689 (N_19689,N_17339,N_17823);
or U19690 (N_19690,N_15765,N_17369);
xnor U19691 (N_19691,N_17676,N_17635);
and U19692 (N_19692,N_16618,N_15290);
and U19693 (N_19693,N_15351,N_17808);
xnor U19694 (N_19694,N_17966,N_17787);
nor U19695 (N_19695,N_15252,N_17388);
xor U19696 (N_19696,N_16121,N_17061);
or U19697 (N_19697,N_16709,N_16154);
and U19698 (N_19698,N_15987,N_15958);
xor U19699 (N_19699,N_15111,N_17467);
and U19700 (N_19700,N_17566,N_15450);
nor U19701 (N_19701,N_15013,N_15295);
and U19702 (N_19702,N_17758,N_16153);
nand U19703 (N_19703,N_17047,N_16955);
xor U19704 (N_19704,N_16682,N_16189);
xnor U19705 (N_19705,N_17057,N_17594);
and U19706 (N_19706,N_15718,N_16205);
xnor U19707 (N_19707,N_15738,N_16813);
nand U19708 (N_19708,N_17099,N_15090);
nor U19709 (N_19709,N_16589,N_17723);
xor U19710 (N_19710,N_16879,N_16089);
nand U19711 (N_19711,N_17791,N_15064);
and U19712 (N_19712,N_17749,N_17971);
xor U19713 (N_19713,N_17983,N_16856);
nor U19714 (N_19714,N_17551,N_15536);
or U19715 (N_19715,N_15964,N_17355);
or U19716 (N_19716,N_17046,N_17936);
xnor U19717 (N_19717,N_16005,N_16100);
or U19718 (N_19718,N_17478,N_16659);
xor U19719 (N_19719,N_17454,N_17076);
and U19720 (N_19720,N_17385,N_16967);
xnor U19721 (N_19721,N_17128,N_15123);
or U19722 (N_19722,N_16783,N_15737);
nor U19723 (N_19723,N_16412,N_16249);
xnor U19724 (N_19724,N_16472,N_17180);
or U19725 (N_19725,N_17376,N_16910);
nor U19726 (N_19726,N_17960,N_17002);
nand U19727 (N_19727,N_16701,N_16915);
xor U19728 (N_19728,N_17273,N_15722);
nand U19729 (N_19729,N_16228,N_17512);
or U19730 (N_19730,N_15109,N_17889);
xor U19731 (N_19731,N_17533,N_15323);
and U19732 (N_19732,N_16198,N_16187);
nor U19733 (N_19733,N_17805,N_15081);
and U19734 (N_19734,N_15035,N_17828);
nor U19735 (N_19735,N_16554,N_15489);
or U19736 (N_19736,N_15951,N_15453);
or U19737 (N_19737,N_16773,N_17297);
nand U19738 (N_19738,N_16845,N_15218);
nor U19739 (N_19739,N_15758,N_17064);
xor U19740 (N_19740,N_17023,N_15087);
xor U19741 (N_19741,N_17260,N_16547);
xor U19742 (N_19742,N_15402,N_16864);
nor U19743 (N_19743,N_17731,N_16955);
nor U19744 (N_19744,N_17154,N_15935);
nand U19745 (N_19745,N_16601,N_16293);
or U19746 (N_19746,N_15722,N_15252);
nor U19747 (N_19747,N_15405,N_16709);
nor U19748 (N_19748,N_17388,N_16848);
or U19749 (N_19749,N_16788,N_17218);
nor U19750 (N_19750,N_15116,N_17536);
nor U19751 (N_19751,N_15105,N_17857);
nor U19752 (N_19752,N_16485,N_15222);
nand U19753 (N_19753,N_15450,N_15506);
and U19754 (N_19754,N_15373,N_17234);
and U19755 (N_19755,N_17498,N_16265);
nand U19756 (N_19756,N_17657,N_16235);
and U19757 (N_19757,N_16394,N_16517);
and U19758 (N_19758,N_16849,N_17375);
and U19759 (N_19759,N_15085,N_16514);
and U19760 (N_19760,N_16678,N_16930);
or U19761 (N_19761,N_16328,N_15317);
xor U19762 (N_19762,N_15345,N_15975);
and U19763 (N_19763,N_15672,N_17895);
xnor U19764 (N_19764,N_16751,N_15569);
or U19765 (N_19765,N_16546,N_16417);
or U19766 (N_19766,N_17783,N_15182);
and U19767 (N_19767,N_16475,N_16133);
or U19768 (N_19768,N_17009,N_16902);
and U19769 (N_19769,N_16932,N_17668);
nand U19770 (N_19770,N_15180,N_17087);
xor U19771 (N_19771,N_16289,N_16370);
and U19772 (N_19772,N_17391,N_15597);
or U19773 (N_19773,N_17545,N_17474);
nand U19774 (N_19774,N_17942,N_16621);
or U19775 (N_19775,N_15823,N_15789);
and U19776 (N_19776,N_17750,N_17250);
and U19777 (N_19777,N_16345,N_15961);
or U19778 (N_19778,N_16528,N_17569);
xnor U19779 (N_19779,N_15506,N_17132);
nor U19780 (N_19780,N_17183,N_16499);
nand U19781 (N_19781,N_16772,N_17066);
nand U19782 (N_19782,N_17427,N_17316);
and U19783 (N_19783,N_16517,N_17611);
and U19784 (N_19784,N_15618,N_16944);
xnor U19785 (N_19785,N_15239,N_15442);
nand U19786 (N_19786,N_17850,N_15202);
or U19787 (N_19787,N_16141,N_17155);
nand U19788 (N_19788,N_16363,N_17481);
and U19789 (N_19789,N_16919,N_15211);
nand U19790 (N_19790,N_16384,N_15070);
nand U19791 (N_19791,N_15617,N_16449);
xor U19792 (N_19792,N_17525,N_16355);
xor U19793 (N_19793,N_17578,N_17260);
nand U19794 (N_19794,N_15390,N_17121);
or U19795 (N_19795,N_16021,N_16181);
nor U19796 (N_19796,N_17282,N_15918);
and U19797 (N_19797,N_15501,N_17940);
nand U19798 (N_19798,N_15840,N_17538);
and U19799 (N_19799,N_17799,N_17900);
nand U19800 (N_19800,N_15610,N_15767);
nand U19801 (N_19801,N_16882,N_16539);
xor U19802 (N_19802,N_15541,N_16510);
nor U19803 (N_19803,N_17675,N_15518);
nand U19804 (N_19804,N_16480,N_15939);
or U19805 (N_19805,N_16017,N_17209);
and U19806 (N_19806,N_16674,N_17698);
and U19807 (N_19807,N_16507,N_16137);
and U19808 (N_19808,N_15219,N_17802);
or U19809 (N_19809,N_16341,N_15786);
or U19810 (N_19810,N_16947,N_16169);
nor U19811 (N_19811,N_17243,N_17219);
and U19812 (N_19812,N_17280,N_16674);
nor U19813 (N_19813,N_16361,N_16447);
and U19814 (N_19814,N_15352,N_15283);
xor U19815 (N_19815,N_15261,N_15112);
nor U19816 (N_19816,N_16565,N_17384);
xor U19817 (N_19817,N_16362,N_16177);
or U19818 (N_19818,N_16184,N_17398);
and U19819 (N_19819,N_16318,N_15518);
and U19820 (N_19820,N_16547,N_17689);
or U19821 (N_19821,N_15499,N_15461);
nand U19822 (N_19822,N_15231,N_15472);
and U19823 (N_19823,N_17857,N_17667);
and U19824 (N_19824,N_15480,N_17039);
nand U19825 (N_19825,N_17130,N_17915);
nand U19826 (N_19826,N_17371,N_15243);
xor U19827 (N_19827,N_15268,N_16994);
nor U19828 (N_19828,N_16750,N_17134);
nor U19829 (N_19829,N_16026,N_17221);
nand U19830 (N_19830,N_17128,N_15628);
or U19831 (N_19831,N_15170,N_16663);
xor U19832 (N_19832,N_16950,N_16041);
xor U19833 (N_19833,N_16084,N_16064);
and U19834 (N_19834,N_15187,N_15066);
nand U19835 (N_19835,N_17621,N_16354);
xnor U19836 (N_19836,N_17795,N_15711);
xnor U19837 (N_19837,N_17015,N_15242);
or U19838 (N_19838,N_16648,N_15554);
and U19839 (N_19839,N_16130,N_15738);
nor U19840 (N_19840,N_17946,N_16192);
and U19841 (N_19841,N_15752,N_16072);
nor U19842 (N_19842,N_16342,N_17196);
or U19843 (N_19843,N_16884,N_17300);
nand U19844 (N_19844,N_16595,N_16975);
xor U19845 (N_19845,N_16169,N_16893);
xor U19846 (N_19846,N_17594,N_16068);
xor U19847 (N_19847,N_16722,N_16503);
xor U19848 (N_19848,N_16991,N_16556);
and U19849 (N_19849,N_17251,N_15283);
xor U19850 (N_19850,N_17223,N_17968);
and U19851 (N_19851,N_16166,N_17823);
or U19852 (N_19852,N_17666,N_16688);
or U19853 (N_19853,N_17812,N_15739);
nor U19854 (N_19854,N_16847,N_16614);
nand U19855 (N_19855,N_16034,N_16312);
nand U19856 (N_19856,N_17565,N_16438);
xnor U19857 (N_19857,N_16699,N_16637);
and U19858 (N_19858,N_15137,N_15200);
or U19859 (N_19859,N_17631,N_17569);
xnor U19860 (N_19860,N_16824,N_16461);
or U19861 (N_19861,N_15210,N_17466);
xor U19862 (N_19862,N_15946,N_15215);
and U19863 (N_19863,N_17057,N_17947);
nor U19864 (N_19864,N_15576,N_17027);
nand U19865 (N_19865,N_16656,N_17628);
and U19866 (N_19866,N_16958,N_15534);
and U19867 (N_19867,N_17049,N_17586);
and U19868 (N_19868,N_16045,N_15225);
nand U19869 (N_19869,N_15373,N_16428);
nor U19870 (N_19870,N_15981,N_17711);
xor U19871 (N_19871,N_17313,N_15986);
nand U19872 (N_19872,N_16513,N_15180);
nor U19873 (N_19873,N_15841,N_16515);
nor U19874 (N_19874,N_17951,N_16550);
and U19875 (N_19875,N_17304,N_17936);
and U19876 (N_19876,N_15647,N_15035);
nand U19877 (N_19877,N_17915,N_15752);
and U19878 (N_19878,N_16045,N_16200);
xnor U19879 (N_19879,N_17380,N_16017);
nand U19880 (N_19880,N_16862,N_15075);
xnor U19881 (N_19881,N_16911,N_17392);
xnor U19882 (N_19882,N_17892,N_17534);
nor U19883 (N_19883,N_16715,N_16746);
nand U19884 (N_19884,N_16668,N_17788);
nand U19885 (N_19885,N_16663,N_16514);
nor U19886 (N_19886,N_15362,N_17171);
or U19887 (N_19887,N_17608,N_15258);
nor U19888 (N_19888,N_15373,N_16204);
nor U19889 (N_19889,N_16695,N_17829);
nor U19890 (N_19890,N_17479,N_15618);
xor U19891 (N_19891,N_17138,N_16092);
xor U19892 (N_19892,N_17264,N_16983);
nand U19893 (N_19893,N_17754,N_16057);
nor U19894 (N_19894,N_17865,N_16925);
nand U19895 (N_19895,N_17039,N_16128);
nor U19896 (N_19896,N_15050,N_16926);
nand U19897 (N_19897,N_16771,N_16346);
xor U19898 (N_19898,N_17371,N_16417);
or U19899 (N_19899,N_17320,N_17476);
xor U19900 (N_19900,N_15999,N_17995);
or U19901 (N_19901,N_15264,N_15480);
xor U19902 (N_19902,N_17044,N_17486);
and U19903 (N_19903,N_16346,N_17744);
and U19904 (N_19904,N_17730,N_16431);
nor U19905 (N_19905,N_16559,N_17394);
and U19906 (N_19906,N_17376,N_17442);
xnor U19907 (N_19907,N_15353,N_15241);
nor U19908 (N_19908,N_16393,N_17345);
nand U19909 (N_19909,N_17878,N_15138);
xnor U19910 (N_19910,N_16920,N_17058);
xor U19911 (N_19911,N_15211,N_16470);
xnor U19912 (N_19912,N_16750,N_17844);
nor U19913 (N_19913,N_17668,N_16297);
nand U19914 (N_19914,N_15112,N_17784);
xor U19915 (N_19915,N_15536,N_16764);
or U19916 (N_19916,N_15780,N_16838);
and U19917 (N_19917,N_16107,N_16916);
nand U19918 (N_19918,N_16433,N_15667);
nand U19919 (N_19919,N_16711,N_15588);
and U19920 (N_19920,N_15675,N_16914);
xor U19921 (N_19921,N_17425,N_16491);
and U19922 (N_19922,N_17647,N_15038);
xnor U19923 (N_19923,N_17481,N_17252);
and U19924 (N_19924,N_16680,N_15489);
nand U19925 (N_19925,N_15426,N_17913);
nor U19926 (N_19926,N_16739,N_17596);
nor U19927 (N_19927,N_17246,N_16426);
and U19928 (N_19928,N_16562,N_16376);
and U19929 (N_19929,N_15059,N_15491);
xnor U19930 (N_19930,N_17745,N_15991);
and U19931 (N_19931,N_15147,N_17152);
nand U19932 (N_19932,N_17376,N_17435);
and U19933 (N_19933,N_15303,N_15587);
xnor U19934 (N_19934,N_15707,N_16169);
nor U19935 (N_19935,N_16568,N_17004);
or U19936 (N_19936,N_16782,N_15472);
xor U19937 (N_19937,N_16092,N_16954);
nor U19938 (N_19938,N_16351,N_16624);
and U19939 (N_19939,N_15282,N_15200);
and U19940 (N_19940,N_17820,N_15566);
xor U19941 (N_19941,N_17790,N_15239);
or U19942 (N_19942,N_16176,N_16521);
nand U19943 (N_19943,N_17074,N_15453);
xnor U19944 (N_19944,N_15944,N_17432);
and U19945 (N_19945,N_15825,N_15925);
xnor U19946 (N_19946,N_15013,N_16205);
or U19947 (N_19947,N_17738,N_15839);
nor U19948 (N_19948,N_17277,N_15373);
xnor U19949 (N_19949,N_16727,N_17306);
and U19950 (N_19950,N_17182,N_16865);
nor U19951 (N_19951,N_15454,N_15041);
nand U19952 (N_19952,N_15998,N_16392);
or U19953 (N_19953,N_15303,N_16140);
nor U19954 (N_19954,N_16762,N_15939);
xnor U19955 (N_19955,N_17576,N_17181);
xor U19956 (N_19956,N_16442,N_15416);
nand U19957 (N_19957,N_16975,N_15582);
or U19958 (N_19958,N_16434,N_17982);
nand U19959 (N_19959,N_17984,N_15421);
xnor U19960 (N_19960,N_16902,N_17435);
or U19961 (N_19961,N_16184,N_16162);
and U19962 (N_19962,N_17426,N_15664);
xor U19963 (N_19963,N_16624,N_15276);
and U19964 (N_19964,N_16496,N_15191);
xnor U19965 (N_19965,N_15465,N_17860);
and U19966 (N_19966,N_16202,N_17198);
nor U19967 (N_19967,N_15396,N_17009);
nand U19968 (N_19968,N_17780,N_17159);
or U19969 (N_19969,N_16844,N_16818);
or U19970 (N_19970,N_17711,N_16708);
xnor U19971 (N_19971,N_16302,N_15850);
and U19972 (N_19972,N_15139,N_16745);
nand U19973 (N_19973,N_16370,N_16647);
and U19974 (N_19974,N_17432,N_15407);
or U19975 (N_19975,N_16826,N_15884);
nor U19976 (N_19976,N_17297,N_15773);
or U19977 (N_19977,N_17353,N_16866);
and U19978 (N_19978,N_16185,N_17740);
and U19979 (N_19979,N_16906,N_15599);
and U19980 (N_19980,N_17253,N_17039);
and U19981 (N_19981,N_17037,N_16985);
nand U19982 (N_19982,N_15667,N_15145);
or U19983 (N_19983,N_17968,N_15103);
nand U19984 (N_19984,N_15017,N_16452);
and U19985 (N_19985,N_16430,N_17661);
or U19986 (N_19986,N_15253,N_15569);
nand U19987 (N_19987,N_15941,N_17455);
nor U19988 (N_19988,N_17242,N_17395);
nand U19989 (N_19989,N_17399,N_15668);
nor U19990 (N_19990,N_15795,N_16634);
or U19991 (N_19991,N_17968,N_15498);
xor U19992 (N_19992,N_15240,N_17539);
or U19993 (N_19993,N_15377,N_16145);
or U19994 (N_19994,N_17741,N_16458);
or U19995 (N_19995,N_17312,N_17711);
nor U19996 (N_19996,N_15226,N_16120);
and U19997 (N_19997,N_16293,N_17616);
or U19998 (N_19998,N_15924,N_15330);
and U19999 (N_19999,N_15677,N_17662);
and U20000 (N_20000,N_17568,N_16145);
and U20001 (N_20001,N_16270,N_15452);
xor U20002 (N_20002,N_15247,N_15409);
nand U20003 (N_20003,N_17960,N_15996);
and U20004 (N_20004,N_15342,N_16339);
nor U20005 (N_20005,N_16404,N_17162);
or U20006 (N_20006,N_15156,N_15984);
nor U20007 (N_20007,N_17689,N_15223);
nand U20008 (N_20008,N_17551,N_15109);
xor U20009 (N_20009,N_15348,N_15813);
xnor U20010 (N_20010,N_15602,N_15649);
or U20011 (N_20011,N_17998,N_15912);
or U20012 (N_20012,N_15344,N_15583);
and U20013 (N_20013,N_15859,N_17201);
nor U20014 (N_20014,N_15351,N_17032);
nor U20015 (N_20015,N_16762,N_17090);
and U20016 (N_20016,N_15367,N_15033);
xor U20017 (N_20017,N_16985,N_15612);
or U20018 (N_20018,N_16963,N_15778);
nor U20019 (N_20019,N_15147,N_17377);
nor U20020 (N_20020,N_17079,N_15913);
nand U20021 (N_20021,N_17049,N_15543);
nand U20022 (N_20022,N_17984,N_16785);
nor U20023 (N_20023,N_17350,N_15685);
nor U20024 (N_20024,N_16262,N_15513);
nor U20025 (N_20025,N_16381,N_16376);
and U20026 (N_20026,N_17577,N_16959);
or U20027 (N_20027,N_17441,N_16173);
and U20028 (N_20028,N_15855,N_16918);
nand U20029 (N_20029,N_15316,N_15285);
or U20030 (N_20030,N_17254,N_16325);
nand U20031 (N_20031,N_15342,N_17383);
and U20032 (N_20032,N_17943,N_16070);
or U20033 (N_20033,N_15884,N_16581);
and U20034 (N_20034,N_16973,N_15682);
nand U20035 (N_20035,N_15817,N_15329);
and U20036 (N_20036,N_15872,N_16192);
and U20037 (N_20037,N_17571,N_16925);
or U20038 (N_20038,N_16184,N_17448);
nand U20039 (N_20039,N_16010,N_16205);
xor U20040 (N_20040,N_16553,N_17992);
or U20041 (N_20041,N_17926,N_16571);
and U20042 (N_20042,N_15939,N_15292);
nand U20043 (N_20043,N_15856,N_16532);
and U20044 (N_20044,N_16210,N_15125);
or U20045 (N_20045,N_16280,N_15171);
nor U20046 (N_20046,N_16745,N_15954);
nor U20047 (N_20047,N_17358,N_17929);
nor U20048 (N_20048,N_17799,N_16773);
nand U20049 (N_20049,N_15175,N_17550);
and U20050 (N_20050,N_15341,N_17798);
or U20051 (N_20051,N_16321,N_15307);
or U20052 (N_20052,N_15819,N_15373);
nand U20053 (N_20053,N_15950,N_15122);
nand U20054 (N_20054,N_16452,N_16453);
or U20055 (N_20055,N_17186,N_17262);
nor U20056 (N_20056,N_17371,N_16656);
nor U20057 (N_20057,N_16643,N_16057);
xor U20058 (N_20058,N_17606,N_17884);
and U20059 (N_20059,N_16331,N_16277);
nand U20060 (N_20060,N_15841,N_16150);
nand U20061 (N_20061,N_15184,N_17700);
and U20062 (N_20062,N_17096,N_16130);
or U20063 (N_20063,N_16553,N_16778);
or U20064 (N_20064,N_17220,N_17958);
nand U20065 (N_20065,N_17871,N_16703);
nor U20066 (N_20066,N_16321,N_17282);
or U20067 (N_20067,N_17665,N_17452);
nor U20068 (N_20068,N_16310,N_16272);
nand U20069 (N_20069,N_15557,N_15140);
or U20070 (N_20070,N_16573,N_16414);
nor U20071 (N_20071,N_15268,N_17471);
xnor U20072 (N_20072,N_15947,N_16357);
and U20073 (N_20073,N_16051,N_16326);
and U20074 (N_20074,N_16090,N_15513);
or U20075 (N_20075,N_16182,N_15711);
or U20076 (N_20076,N_16422,N_15140);
nor U20077 (N_20077,N_16659,N_15622);
nor U20078 (N_20078,N_15662,N_15221);
xor U20079 (N_20079,N_17080,N_16409);
nor U20080 (N_20080,N_15328,N_16676);
nand U20081 (N_20081,N_17297,N_17205);
nor U20082 (N_20082,N_16243,N_15906);
nand U20083 (N_20083,N_15056,N_15992);
nor U20084 (N_20084,N_17621,N_15143);
and U20085 (N_20085,N_16731,N_16172);
or U20086 (N_20086,N_16504,N_15064);
nand U20087 (N_20087,N_17438,N_17181);
nor U20088 (N_20088,N_17715,N_16744);
nand U20089 (N_20089,N_16213,N_15468);
nor U20090 (N_20090,N_17508,N_16088);
nand U20091 (N_20091,N_15201,N_17042);
and U20092 (N_20092,N_17548,N_17901);
nand U20093 (N_20093,N_17209,N_16602);
or U20094 (N_20094,N_16583,N_17601);
nand U20095 (N_20095,N_15914,N_17042);
or U20096 (N_20096,N_15233,N_16337);
nand U20097 (N_20097,N_15456,N_16417);
and U20098 (N_20098,N_17692,N_17201);
nor U20099 (N_20099,N_16732,N_16598);
xor U20100 (N_20100,N_16879,N_16931);
nor U20101 (N_20101,N_16749,N_16043);
nor U20102 (N_20102,N_15530,N_15612);
and U20103 (N_20103,N_16556,N_15202);
nor U20104 (N_20104,N_15833,N_16223);
xor U20105 (N_20105,N_17725,N_17755);
xnor U20106 (N_20106,N_17471,N_17596);
xnor U20107 (N_20107,N_17974,N_15086);
and U20108 (N_20108,N_16564,N_15556);
and U20109 (N_20109,N_17345,N_15366);
or U20110 (N_20110,N_15746,N_15138);
nor U20111 (N_20111,N_15454,N_17807);
and U20112 (N_20112,N_16927,N_15852);
xnor U20113 (N_20113,N_15881,N_16586);
or U20114 (N_20114,N_17939,N_17854);
and U20115 (N_20115,N_15740,N_15545);
nor U20116 (N_20116,N_16218,N_16466);
or U20117 (N_20117,N_16756,N_17966);
and U20118 (N_20118,N_16218,N_17205);
nand U20119 (N_20119,N_17019,N_16081);
xnor U20120 (N_20120,N_16268,N_17571);
xnor U20121 (N_20121,N_16963,N_15140);
nand U20122 (N_20122,N_17135,N_17859);
and U20123 (N_20123,N_15526,N_15512);
and U20124 (N_20124,N_17690,N_16098);
or U20125 (N_20125,N_15237,N_15178);
and U20126 (N_20126,N_16699,N_17776);
nand U20127 (N_20127,N_17433,N_17894);
nand U20128 (N_20128,N_16263,N_16230);
nand U20129 (N_20129,N_17755,N_15129);
nor U20130 (N_20130,N_16781,N_16290);
or U20131 (N_20131,N_17052,N_17645);
nand U20132 (N_20132,N_16369,N_17270);
xnor U20133 (N_20133,N_16217,N_15891);
or U20134 (N_20134,N_16383,N_15143);
xnor U20135 (N_20135,N_17120,N_15361);
nand U20136 (N_20136,N_17513,N_17034);
xnor U20137 (N_20137,N_16660,N_15108);
nor U20138 (N_20138,N_17445,N_16709);
xnor U20139 (N_20139,N_17213,N_16314);
nor U20140 (N_20140,N_15622,N_15280);
nor U20141 (N_20141,N_15130,N_17273);
xnor U20142 (N_20142,N_16656,N_17133);
and U20143 (N_20143,N_17744,N_16409);
nor U20144 (N_20144,N_15684,N_17005);
xnor U20145 (N_20145,N_17864,N_16239);
or U20146 (N_20146,N_17915,N_17467);
xnor U20147 (N_20147,N_16443,N_15789);
nand U20148 (N_20148,N_16334,N_15086);
and U20149 (N_20149,N_17858,N_16530);
and U20150 (N_20150,N_15848,N_15843);
nor U20151 (N_20151,N_16567,N_15499);
nor U20152 (N_20152,N_15683,N_15248);
or U20153 (N_20153,N_16837,N_17557);
or U20154 (N_20154,N_17183,N_17272);
nor U20155 (N_20155,N_16266,N_17512);
or U20156 (N_20156,N_16145,N_16356);
or U20157 (N_20157,N_17268,N_16632);
nand U20158 (N_20158,N_15629,N_15360);
or U20159 (N_20159,N_16227,N_16628);
or U20160 (N_20160,N_16116,N_16692);
and U20161 (N_20161,N_17707,N_17342);
xnor U20162 (N_20162,N_17816,N_15400);
nand U20163 (N_20163,N_17926,N_16980);
nand U20164 (N_20164,N_16164,N_16090);
and U20165 (N_20165,N_16122,N_15670);
or U20166 (N_20166,N_17887,N_15188);
or U20167 (N_20167,N_17325,N_17478);
nor U20168 (N_20168,N_16817,N_17001);
xnor U20169 (N_20169,N_15258,N_17137);
or U20170 (N_20170,N_15184,N_15946);
nor U20171 (N_20171,N_15497,N_15736);
nor U20172 (N_20172,N_15686,N_17659);
or U20173 (N_20173,N_15830,N_16362);
xnor U20174 (N_20174,N_15716,N_17989);
nand U20175 (N_20175,N_15344,N_17358);
xor U20176 (N_20176,N_17358,N_16749);
and U20177 (N_20177,N_16656,N_17012);
and U20178 (N_20178,N_16946,N_15310);
and U20179 (N_20179,N_15576,N_16603);
xor U20180 (N_20180,N_16525,N_15741);
nor U20181 (N_20181,N_15727,N_15922);
nor U20182 (N_20182,N_15204,N_16187);
and U20183 (N_20183,N_17892,N_16499);
nor U20184 (N_20184,N_17403,N_15894);
nor U20185 (N_20185,N_16265,N_17377);
xor U20186 (N_20186,N_16189,N_15941);
and U20187 (N_20187,N_17542,N_16952);
and U20188 (N_20188,N_17831,N_16984);
and U20189 (N_20189,N_17679,N_15067);
or U20190 (N_20190,N_15641,N_17414);
or U20191 (N_20191,N_16091,N_16281);
xor U20192 (N_20192,N_15085,N_17723);
nor U20193 (N_20193,N_15086,N_16811);
or U20194 (N_20194,N_17129,N_15459);
xor U20195 (N_20195,N_15308,N_15416);
and U20196 (N_20196,N_15700,N_15824);
xnor U20197 (N_20197,N_16680,N_17249);
nor U20198 (N_20198,N_15064,N_15781);
or U20199 (N_20199,N_15367,N_17223);
and U20200 (N_20200,N_15763,N_16437);
or U20201 (N_20201,N_16537,N_16103);
or U20202 (N_20202,N_17248,N_15269);
and U20203 (N_20203,N_15963,N_15695);
and U20204 (N_20204,N_16895,N_17398);
and U20205 (N_20205,N_17194,N_15535);
and U20206 (N_20206,N_15986,N_16003);
and U20207 (N_20207,N_16395,N_16849);
xnor U20208 (N_20208,N_17324,N_17053);
xor U20209 (N_20209,N_16665,N_15448);
xnor U20210 (N_20210,N_15197,N_17167);
nand U20211 (N_20211,N_17219,N_16428);
xnor U20212 (N_20212,N_15940,N_15464);
and U20213 (N_20213,N_15125,N_15854);
nand U20214 (N_20214,N_17300,N_16351);
nand U20215 (N_20215,N_17095,N_16165);
xor U20216 (N_20216,N_17437,N_16351);
xor U20217 (N_20217,N_16344,N_17914);
or U20218 (N_20218,N_15002,N_16922);
or U20219 (N_20219,N_16175,N_15233);
xnor U20220 (N_20220,N_17616,N_17078);
nor U20221 (N_20221,N_17117,N_15526);
nand U20222 (N_20222,N_17065,N_17537);
xor U20223 (N_20223,N_16848,N_16452);
xor U20224 (N_20224,N_17906,N_15108);
nor U20225 (N_20225,N_15908,N_16146);
nand U20226 (N_20226,N_17738,N_16951);
nand U20227 (N_20227,N_17842,N_16156);
and U20228 (N_20228,N_16016,N_15079);
and U20229 (N_20229,N_17180,N_15383);
and U20230 (N_20230,N_15159,N_15511);
and U20231 (N_20231,N_15987,N_17629);
nor U20232 (N_20232,N_15694,N_17741);
and U20233 (N_20233,N_17304,N_16692);
nand U20234 (N_20234,N_15958,N_17467);
nor U20235 (N_20235,N_16946,N_16762);
or U20236 (N_20236,N_17430,N_16826);
and U20237 (N_20237,N_15422,N_15518);
nor U20238 (N_20238,N_15519,N_15532);
and U20239 (N_20239,N_15343,N_17166);
and U20240 (N_20240,N_15546,N_15983);
nand U20241 (N_20241,N_16851,N_15874);
xor U20242 (N_20242,N_15254,N_16811);
nor U20243 (N_20243,N_17093,N_17525);
nor U20244 (N_20244,N_17176,N_16713);
nor U20245 (N_20245,N_17233,N_17567);
nand U20246 (N_20246,N_16708,N_16162);
nor U20247 (N_20247,N_15982,N_16360);
or U20248 (N_20248,N_17318,N_16118);
nand U20249 (N_20249,N_16590,N_17128);
xnor U20250 (N_20250,N_16535,N_16648);
xor U20251 (N_20251,N_17644,N_16026);
xnor U20252 (N_20252,N_17228,N_15214);
or U20253 (N_20253,N_16958,N_16221);
and U20254 (N_20254,N_17550,N_15684);
or U20255 (N_20255,N_15923,N_15888);
nor U20256 (N_20256,N_15688,N_17121);
and U20257 (N_20257,N_17708,N_16388);
or U20258 (N_20258,N_16619,N_16147);
or U20259 (N_20259,N_15088,N_15028);
or U20260 (N_20260,N_16711,N_16811);
or U20261 (N_20261,N_17111,N_17740);
nor U20262 (N_20262,N_17516,N_15851);
nand U20263 (N_20263,N_15992,N_16954);
or U20264 (N_20264,N_16090,N_15230);
or U20265 (N_20265,N_16144,N_16829);
nor U20266 (N_20266,N_16873,N_16332);
xnor U20267 (N_20267,N_16645,N_16460);
or U20268 (N_20268,N_17159,N_17325);
or U20269 (N_20269,N_16161,N_15999);
and U20270 (N_20270,N_15288,N_17566);
nand U20271 (N_20271,N_17272,N_16892);
or U20272 (N_20272,N_15688,N_15672);
xor U20273 (N_20273,N_17765,N_15213);
and U20274 (N_20274,N_15013,N_16513);
nor U20275 (N_20275,N_15953,N_15955);
nand U20276 (N_20276,N_15973,N_16015);
and U20277 (N_20277,N_15462,N_17283);
nand U20278 (N_20278,N_15483,N_17172);
nand U20279 (N_20279,N_17859,N_15955);
and U20280 (N_20280,N_17773,N_17523);
or U20281 (N_20281,N_16300,N_17591);
nand U20282 (N_20282,N_15353,N_17104);
or U20283 (N_20283,N_17610,N_17297);
and U20284 (N_20284,N_15192,N_15239);
nor U20285 (N_20285,N_15904,N_16152);
nor U20286 (N_20286,N_17388,N_15340);
xor U20287 (N_20287,N_17270,N_15098);
nand U20288 (N_20288,N_15038,N_15719);
or U20289 (N_20289,N_17052,N_15371);
xnor U20290 (N_20290,N_16835,N_17415);
xor U20291 (N_20291,N_17836,N_15514);
nand U20292 (N_20292,N_15909,N_15175);
xor U20293 (N_20293,N_15102,N_17189);
and U20294 (N_20294,N_15471,N_17364);
and U20295 (N_20295,N_16052,N_17934);
nor U20296 (N_20296,N_16758,N_17379);
and U20297 (N_20297,N_15020,N_15550);
nand U20298 (N_20298,N_17697,N_17301);
or U20299 (N_20299,N_15685,N_16048);
xnor U20300 (N_20300,N_17571,N_16699);
xor U20301 (N_20301,N_17695,N_17847);
or U20302 (N_20302,N_15437,N_17372);
nand U20303 (N_20303,N_17806,N_15260);
nor U20304 (N_20304,N_16994,N_15993);
nand U20305 (N_20305,N_17928,N_15811);
nand U20306 (N_20306,N_16791,N_17801);
xnor U20307 (N_20307,N_17291,N_16223);
and U20308 (N_20308,N_16739,N_15961);
xor U20309 (N_20309,N_15374,N_16533);
nor U20310 (N_20310,N_17752,N_16230);
nand U20311 (N_20311,N_17511,N_15872);
nand U20312 (N_20312,N_17053,N_15158);
nand U20313 (N_20313,N_16409,N_15069);
nor U20314 (N_20314,N_15831,N_17601);
and U20315 (N_20315,N_16614,N_15666);
xnor U20316 (N_20316,N_16156,N_15623);
nand U20317 (N_20317,N_16053,N_17515);
nor U20318 (N_20318,N_15129,N_17222);
nand U20319 (N_20319,N_15952,N_17390);
nand U20320 (N_20320,N_15092,N_16577);
and U20321 (N_20321,N_15230,N_16867);
nand U20322 (N_20322,N_16880,N_17218);
xor U20323 (N_20323,N_16449,N_15072);
nor U20324 (N_20324,N_17198,N_16263);
nor U20325 (N_20325,N_16909,N_15950);
and U20326 (N_20326,N_16178,N_16901);
nor U20327 (N_20327,N_16186,N_15044);
nor U20328 (N_20328,N_16653,N_16821);
and U20329 (N_20329,N_17669,N_17807);
or U20330 (N_20330,N_16518,N_15693);
nor U20331 (N_20331,N_17672,N_15178);
xor U20332 (N_20332,N_15950,N_15593);
or U20333 (N_20333,N_15845,N_16096);
nand U20334 (N_20334,N_17361,N_16963);
nor U20335 (N_20335,N_16093,N_15094);
and U20336 (N_20336,N_16021,N_17324);
nand U20337 (N_20337,N_17140,N_17822);
and U20338 (N_20338,N_16754,N_15240);
or U20339 (N_20339,N_16039,N_17574);
nand U20340 (N_20340,N_15024,N_15642);
and U20341 (N_20341,N_17056,N_15475);
xor U20342 (N_20342,N_17646,N_17525);
xnor U20343 (N_20343,N_15512,N_17373);
xor U20344 (N_20344,N_15707,N_17352);
nand U20345 (N_20345,N_17760,N_17195);
and U20346 (N_20346,N_16370,N_15796);
xnor U20347 (N_20347,N_15922,N_15602);
nor U20348 (N_20348,N_15161,N_15140);
xor U20349 (N_20349,N_15315,N_17233);
or U20350 (N_20350,N_15806,N_17054);
nand U20351 (N_20351,N_17878,N_15358);
or U20352 (N_20352,N_15002,N_16108);
and U20353 (N_20353,N_17788,N_15143);
nor U20354 (N_20354,N_16894,N_17283);
nand U20355 (N_20355,N_15541,N_17292);
nor U20356 (N_20356,N_16592,N_17876);
nand U20357 (N_20357,N_15315,N_15427);
nor U20358 (N_20358,N_15809,N_17082);
or U20359 (N_20359,N_15621,N_17169);
nor U20360 (N_20360,N_17239,N_15695);
nand U20361 (N_20361,N_16886,N_16416);
and U20362 (N_20362,N_16164,N_17681);
nor U20363 (N_20363,N_17095,N_16924);
nand U20364 (N_20364,N_15744,N_15979);
nor U20365 (N_20365,N_17934,N_15439);
nand U20366 (N_20366,N_16969,N_16688);
or U20367 (N_20367,N_16217,N_17128);
xor U20368 (N_20368,N_17087,N_15840);
xor U20369 (N_20369,N_16092,N_15986);
xor U20370 (N_20370,N_16375,N_16238);
and U20371 (N_20371,N_17720,N_16212);
nor U20372 (N_20372,N_17671,N_17406);
or U20373 (N_20373,N_15682,N_16709);
or U20374 (N_20374,N_16777,N_16058);
xnor U20375 (N_20375,N_16342,N_16476);
nor U20376 (N_20376,N_15184,N_16519);
xnor U20377 (N_20377,N_15960,N_15705);
or U20378 (N_20378,N_16723,N_16454);
and U20379 (N_20379,N_17087,N_17891);
or U20380 (N_20380,N_16343,N_17497);
nor U20381 (N_20381,N_17206,N_15475);
nand U20382 (N_20382,N_17348,N_16739);
and U20383 (N_20383,N_17838,N_15445);
or U20384 (N_20384,N_17756,N_15079);
and U20385 (N_20385,N_17377,N_16873);
and U20386 (N_20386,N_17600,N_16572);
nand U20387 (N_20387,N_16456,N_17417);
nor U20388 (N_20388,N_17234,N_16075);
nand U20389 (N_20389,N_16329,N_17952);
nor U20390 (N_20390,N_17207,N_17929);
and U20391 (N_20391,N_15354,N_15512);
or U20392 (N_20392,N_16706,N_17117);
xnor U20393 (N_20393,N_17674,N_15690);
nor U20394 (N_20394,N_17012,N_17205);
or U20395 (N_20395,N_16018,N_16434);
nor U20396 (N_20396,N_16820,N_17372);
nand U20397 (N_20397,N_15064,N_17488);
nor U20398 (N_20398,N_15170,N_16004);
nor U20399 (N_20399,N_15758,N_16475);
or U20400 (N_20400,N_15220,N_16806);
xnor U20401 (N_20401,N_16272,N_16824);
and U20402 (N_20402,N_17890,N_16908);
and U20403 (N_20403,N_17866,N_17816);
xnor U20404 (N_20404,N_16541,N_17747);
or U20405 (N_20405,N_16853,N_17002);
and U20406 (N_20406,N_16689,N_16616);
nor U20407 (N_20407,N_17144,N_15196);
and U20408 (N_20408,N_16278,N_16620);
nor U20409 (N_20409,N_17045,N_17036);
and U20410 (N_20410,N_17207,N_17357);
or U20411 (N_20411,N_15624,N_16585);
and U20412 (N_20412,N_16825,N_16123);
nand U20413 (N_20413,N_16552,N_16068);
nor U20414 (N_20414,N_17233,N_17152);
or U20415 (N_20415,N_17748,N_17196);
or U20416 (N_20416,N_16957,N_16273);
xnor U20417 (N_20417,N_15491,N_15841);
nor U20418 (N_20418,N_15134,N_15846);
and U20419 (N_20419,N_16194,N_16012);
and U20420 (N_20420,N_16256,N_17151);
or U20421 (N_20421,N_16290,N_15913);
xnor U20422 (N_20422,N_15334,N_17696);
nand U20423 (N_20423,N_16057,N_16577);
or U20424 (N_20424,N_17341,N_16776);
nand U20425 (N_20425,N_15458,N_17383);
nor U20426 (N_20426,N_17021,N_17098);
xor U20427 (N_20427,N_16409,N_17983);
and U20428 (N_20428,N_16001,N_17423);
and U20429 (N_20429,N_16942,N_15131);
and U20430 (N_20430,N_17126,N_17148);
nor U20431 (N_20431,N_17406,N_17605);
nor U20432 (N_20432,N_15777,N_17496);
or U20433 (N_20433,N_15083,N_17571);
nand U20434 (N_20434,N_16749,N_15157);
xnor U20435 (N_20435,N_15854,N_15161);
or U20436 (N_20436,N_15659,N_16817);
nor U20437 (N_20437,N_16497,N_15427);
xor U20438 (N_20438,N_15233,N_17771);
and U20439 (N_20439,N_17446,N_16442);
xor U20440 (N_20440,N_16644,N_15762);
nor U20441 (N_20441,N_17574,N_15964);
nor U20442 (N_20442,N_15073,N_16674);
nor U20443 (N_20443,N_15414,N_16425);
or U20444 (N_20444,N_16411,N_15971);
or U20445 (N_20445,N_17688,N_16290);
or U20446 (N_20446,N_17793,N_16339);
nor U20447 (N_20447,N_15577,N_17461);
and U20448 (N_20448,N_15331,N_15642);
or U20449 (N_20449,N_17532,N_16501);
or U20450 (N_20450,N_16063,N_16695);
and U20451 (N_20451,N_17649,N_15920);
nor U20452 (N_20452,N_17569,N_16057);
nand U20453 (N_20453,N_16340,N_16651);
nand U20454 (N_20454,N_17108,N_16243);
or U20455 (N_20455,N_16685,N_16817);
xnor U20456 (N_20456,N_17582,N_16188);
and U20457 (N_20457,N_17155,N_17892);
xnor U20458 (N_20458,N_15838,N_16950);
or U20459 (N_20459,N_15680,N_17353);
nor U20460 (N_20460,N_15050,N_17619);
nor U20461 (N_20461,N_15268,N_16674);
xor U20462 (N_20462,N_16693,N_17083);
and U20463 (N_20463,N_15658,N_15196);
and U20464 (N_20464,N_17030,N_17965);
xnor U20465 (N_20465,N_15607,N_16754);
nor U20466 (N_20466,N_16793,N_16338);
or U20467 (N_20467,N_16695,N_16602);
nor U20468 (N_20468,N_17452,N_15289);
xnor U20469 (N_20469,N_15232,N_17861);
or U20470 (N_20470,N_17664,N_16496);
xnor U20471 (N_20471,N_15112,N_16694);
and U20472 (N_20472,N_16555,N_17028);
nand U20473 (N_20473,N_17610,N_15164);
and U20474 (N_20474,N_17755,N_15928);
and U20475 (N_20475,N_15307,N_17376);
xor U20476 (N_20476,N_16500,N_17846);
and U20477 (N_20477,N_17335,N_17902);
nor U20478 (N_20478,N_15536,N_17194);
or U20479 (N_20479,N_17414,N_16212);
nand U20480 (N_20480,N_16845,N_16659);
and U20481 (N_20481,N_15118,N_16880);
nor U20482 (N_20482,N_16927,N_15951);
nand U20483 (N_20483,N_16922,N_15448);
and U20484 (N_20484,N_17069,N_16764);
or U20485 (N_20485,N_15329,N_17611);
nand U20486 (N_20486,N_17520,N_17228);
nand U20487 (N_20487,N_17418,N_16221);
nand U20488 (N_20488,N_15490,N_17757);
or U20489 (N_20489,N_15389,N_17966);
nor U20490 (N_20490,N_16052,N_15509);
or U20491 (N_20491,N_17865,N_17891);
and U20492 (N_20492,N_17155,N_17427);
or U20493 (N_20493,N_16352,N_15714);
and U20494 (N_20494,N_17851,N_15021);
and U20495 (N_20495,N_15125,N_15460);
xnor U20496 (N_20496,N_16402,N_17077);
nand U20497 (N_20497,N_17506,N_17488);
xor U20498 (N_20498,N_17702,N_16466);
or U20499 (N_20499,N_15060,N_17958);
nor U20500 (N_20500,N_17087,N_15461);
nor U20501 (N_20501,N_16733,N_17308);
nor U20502 (N_20502,N_15426,N_16478);
or U20503 (N_20503,N_17415,N_17326);
xor U20504 (N_20504,N_15487,N_15488);
xnor U20505 (N_20505,N_17318,N_15741);
xor U20506 (N_20506,N_15367,N_17466);
or U20507 (N_20507,N_15699,N_17161);
and U20508 (N_20508,N_16606,N_17309);
nor U20509 (N_20509,N_16651,N_16664);
xor U20510 (N_20510,N_16155,N_17972);
nand U20511 (N_20511,N_15924,N_15686);
xnor U20512 (N_20512,N_16543,N_16248);
and U20513 (N_20513,N_16053,N_16120);
or U20514 (N_20514,N_16139,N_15049);
or U20515 (N_20515,N_15445,N_15915);
and U20516 (N_20516,N_15684,N_15981);
xor U20517 (N_20517,N_16471,N_16983);
and U20518 (N_20518,N_17849,N_16448);
nand U20519 (N_20519,N_16827,N_15035);
nand U20520 (N_20520,N_15364,N_16251);
xnor U20521 (N_20521,N_17378,N_15884);
or U20522 (N_20522,N_16159,N_15046);
and U20523 (N_20523,N_16896,N_15598);
nor U20524 (N_20524,N_16988,N_16368);
nor U20525 (N_20525,N_15949,N_15545);
nand U20526 (N_20526,N_16853,N_15574);
and U20527 (N_20527,N_15290,N_16178);
nor U20528 (N_20528,N_17550,N_17497);
or U20529 (N_20529,N_16771,N_15823);
and U20530 (N_20530,N_15065,N_15121);
or U20531 (N_20531,N_17698,N_16361);
nand U20532 (N_20532,N_15666,N_16355);
xor U20533 (N_20533,N_17734,N_16421);
xnor U20534 (N_20534,N_15425,N_15216);
xor U20535 (N_20535,N_16169,N_15376);
xnor U20536 (N_20536,N_16896,N_15928);
nand U20537 (N_20537,N_15378,N_17344);
nor U20538 (N_20538,N_17415,N_15138);
and U20539 (N_20539,N_16885,N_17334);
xor U20540 (N_20540,N_15501,N_17008);
nand U20541 (N_20541,N_15533,N_15202);
and U20542 (N_20542,N_15213,N_17113);
or U20543 (N_20543,N_17673,N_16770);
xnor U20544 (N_20544,N_17736,N_17877);
and U20545 (N_20545,N_17379,N_16458);
xor U20546 (N_20546,N_16701,N_16619);
nor U20547 (N_20547,N_15797,N_16771);
xor U20548 (N_20548,N_17721,N_16207);
or U20549 (N_20549,N_15423,N_17891);
nand U20550 (N_20550,N_16485,N_17852);
and U20551 (N_20551,N_15409,N_15732);
nor U20552 (N_20552,N_17896,N_17058);
and U20553 (N_20553,N_15397,N_16688);
or U20554 (N_20554,N_16847,N_15713);
nor U20555 (N_20555,N_17274,N_17193);
nor U20556 (N_20556,N_16873,N_17262);
nor U20557 (N_20557,N_15513,N_16592);
xor U20558 (N_20558,N_17617,N_15150);
and U20559 (N_20559,N_15746,N_17406);
or U20560 (N_20560,N_16762,N_16485);
or U20561 (N_20561,N_17103,N_17763);
and U20562 (N_20562,N_17378,N_17100);
xnor U20563 (N_20563,N_15217,N_16595);
or U20564 (N_20564,N_17910,N_17483);
and U20565 (N_20565,N_16004,N_15491);
nor U20566 (N_20566,N_16645,N_17841);
and U20567 (N_20567,N_15732,N_15349);
or U20568 (N_20568,N_15625,N_16747);
nand U20569 (N_20569,N_15867,N_16749);
nand U20570 (N_20570,N_15842,N_17921);
and U20571 (N_20571,N_16043,N_17319);
nor U20572 (N_20572,N_16703,N_17247);
nor U20573 (N_20573,N_16315,N_15179);
or U20574 (N_20574,N_17092,N_15069);
nor U20575 (N_20575,N_16841,N_17521);
nor U20576 (N_20576,N_16201,N_17346);
nor U20577 (N_20577,N_15036,N_16072);
or U20578 (N_20578,N_16511,N_17051);
xor U20579 (N_20579,N_17897,N_15382);
xor U20580 (N_20580,N_15814,N_16328);
and U20581 (N_20581,N_17957,N_16588);
and U20582 (N_20582,N_15559,N_17167);
nor U20583 (N_20583,N_15852,N_17278);
and U20584 (N_20584,N_16623,N_15731);
or U20585 (N_20585,N_16209,N_15456);
nand U20586 (N_20586,N_16477,N_16608);
nand U20587 (N_20587,N_16667,N_15539);
or U20588 (N_20588,N_17684,N_17949);
or U20589 (N_20589,N_15298,N_16239);
and U20590 (N_20590,N_16518,N_16691);
or U20591 (N_20591,N_15406,N_15176);
and U20592 (N_20592,N_16143,N_15267);
nor U20593 (N_20593,N_15192,N_16570);
or U20594 (N_20594,N_17011,N_16177);
and U20595 (N_20595,N_17741,N_17065);
xor U20596 (N_20596,N_15927,N_15964);
nand U20597 (N_20597,N_15422,N_15802);
and U20598 (N_20598,N_15058,N_16178);
nand U20599 (N_20599,N_15686,N_17102);
nor U20600 (N_20600,N_16516,N_15774);
xnor U20601 (N_20601,N_17567,N_17082);
and U20602 (N_20602,N_15292,N_16739);
or U20603 (N_20603,N_16650,N_15147);
nand U20604 (N_20604,N_17443,N_15755);
nand U20605 (N_20605,N_15433,N_17146);
xnor U20606 (N_20606,N_17422,N_15592);
nor U20607 (N_20607,N_16977,N_17549);
and U20608 (N_20608,N_15045,N_15726);
nor U20609 (N_20609,N_16266,N_15618);
nor U20610 (N_20610,N_15085,N_15793);
xor U20611 (N_20611,N_16451,N_17350);
xnor U20612 (N_20612,N_16628,N_17207);
nor U20613 (N_20613,N_17304,N_17381);
and U20614 (N_20614,N_15641,N_15119);
and U20615 (N_20615,N_15551,N_17577);
or U20616 (N_20616,N_17933,N_16284);
nand U20617 (N_20617,N_16474,N_16951);
or U20618 (N_20618,N_17579,N_15646);
nor U20619 (N_20619,N_17110,N_16096);
nor U20620 (N_20620,N_16709,N_17116);
nand U20621 (N_20621,N_17707,N_17928);
nand U20622 (N_20622,N_17094,N_15467);
nor U20623 (N_20623,N_16087,N_15719);
xor U20624 (N_20624,N_16590,N_16462);
nand U20625 (N_20625,N_16457,N_17822);
nor U20626 (N_20626,N_15561,N_16248);
and U20627 (N_20627,N_15017,N_16060);
xor U20628 (N_20628,N_15511,N_16995);
nor U20629 (N_20629,N_16793,N_17488);
xor U20630 (N_20630,N_15733,N_15305);
nor U20631 (N_20631,N_16819,N_15580);
or U20632 (N_20632,N_15245,N_15137);
nor U20633 (N_20633,N_16335,N_17516);
nor U20634 (N_20634,N_17156,N_15944);
nor U20635 (N_20635,N_16623,N_17987);
nand U20636 (N_20636,N_17187,N_17989);
nor U20637 (N_20637,N_16277,N_15625);
or U20638 (N_20638,N_16691,N_15351);
nand U20639 (N_20639,N_15889,N_17040);
xor U20640 (N_20640,N_17302,N_16408);
nor U20641 (N_20641,N_17686,N_15750);
nor U20642 (N_20642,N_17428,N_16330);
nand U20643 (N_20643,N_15573,N_17266);
nand U20644 (N_20644,N_15394,N_16356);
or U20645 (N_20645,N_15249,N_15195);
nor U20646 (N_20646,N_16499,N_15663);
or U20647 (N_20647,N_17824,N_16148);
or U20648 (N_20648,N_15732,N_17399);
nor U20649 (N_20649,N_17709,N_15274);
nor U20650 (N_20650,N_17640,N_17397);
or U20651 (N_20651,N_17302,N_16416);
or U20652 (N_20652,N_17755,N_15927);
or U20653 (N_20653,N_15711,N_16280);
nor U20654 (N_20654,N_16776,N_17398);
or U20655 (N_20655,N_17250,N_15505);
nor U20656 (N_20656,N_15825,N_17017);
nand U20657 (N_20657,N_17703,N_17397);
xor U20658 (N_20658,N_17041,N_15454);
and U20659 (N_20659,N_15284,N_15301);
and U20660 (N_20660,N_16055,N_15903);
and U20661 (N_20661,N_15485,N_17521);
xor U20662 (N_20662,N_16709,N_15661);
and U20663 (N_20663,N_16181,N_15769);
nor U20664 (N_20664,N_16197,N_15702);
or U20665 (N_20665,N_17406,N_17846);
nand U20666 (N_20666,N_17345,N_16706);
xor U20667 (N_20667,N_15093,N_15539);
nor U20668 (N_20668,N_15668,N_17163);
nand U20669 (N_20669,N_17061,N_16130);
and U20670 (N_20670,N_16254,N_17419);
nor U20671 (N_20671,N_17303,N_16438);
nor U20672 (N_20672,N_17270,N_15048);
or U20673 (N_20673,N_16811,N_15810);
xnor U20674 (N_20674,N_17072,N_15129);
or U20675 (N_20675,N_15581,N_15350);
xnor U20676 (N_20676,N_17456,N_15329);
nand U20677 (N_20677,N_16748,N_15942);
nand U20678 (N_20678,N_16086,N_17106);
xor U20679 (N_20679,N_15195,N_15198);
or U20680 (N_20680,N_15581,N_16051);
nor U20681 (N_20681,N_16591,N_15476);
nor U20682 (N_20682,N_16016,N_17166);
or U20683 (N_20683,N_17500,N_16577);
nor U20684 (N_20684,N_17922,N_16686);
or U20685 (N_20685,N_15318,N_15791);
or U20686 (N_20686,N_17417,N_16170);
xor U20687 (N_20687,N_17301,N_15793);
xnor U20688 (N_20688,N_15637,N_16698);
and U20689 (N_20689,N_17386,N_15266);
nor U20690 (N_20690,N_16316,N_16981);
nor U20691 (N_20691,N_17259,N_17825);
nand U20692 (N_20692,N_16810,N_16625);
nand U20693 (N_20693,N_16844,N_17661);
and U20694 (N_20694,N_15798,N_15504);
and U20695 (N_20695,N_17223,N_17510);
nand U20696 (N_20696,N_15637,N_16461);
and U20697 (N_20697,N_15243,N_17376);
and U20698 (N_20698,N_17352,N_16805);
nor U20699 (N_20699,N_16851,N_15910);
nand U20700 (N_20700,N_15229,N_15042);
or U20701 (N_20701,N_17260,N_17085);
nand U20702 (N_20702,N_17077,N_16182);
xnor U20703 (N_20703,N_15498,N_15046);
nand U20704 (N_20704,N_15568,N_16618);
nand U20705 (N_20705,N_15384,N_16628);
and U20706 (N_20706,N_17634,N_16590);
or U20707 (N_20707,N_17391,N_15811);
nor U20708 (N_20708,N_16900,N_16662);
xor U20709 (N_20709,N_16886,N_17286);
nor U20710 (N_20710,N_15250,N_16029);
or U20711 (N_20711,N_17243,N_17291);
and U20712 (N_20712,N_17179,N_15281);
nand U20713 (N_20713,N_15687,N_15959);
and U20714 (N_20714,N_16831,N_16597);
and U20715 (N_20715,N_15437,N_17033);
xnor U20716 (N_20716,N_17518,N_17210);
and U20717 (N_20717,N_17606,N_17716);
xnor U20718 (N_20718,N_17663,N_15628);
nor U20719 (N_20719,N_16956,N_16840);
xnor U20720 (N_20720,N_16885,N_15472);
xnor U20721 (N_20721,N_15863,N_16744);
or U20722 (N_20722,N_15274,N_15917);
nand U20723 (N_20723,N_17157,N_17906);
nor U20724 (N_20724,N_15635,N_15850);
nor U20725 (N_20725,N_17775,N_17633);
nor U20726 (N_20726,N_16962,N_15548);
or U20727 (N_20727,N_15418,N_15976);
nand U20728 (N_20728,N_17075,N_17970);
or U20729 (N_20729,N_16036,N_17246);
xor U20730 (N_20730,N_17710,N_15648);
xnor U20731 (N_20731,N_17957,N_17049);
or U20732 (N_20732,N_15454,N_15609);
nand U20733 (N_20733,N_15182,N_16291);
or U20734 (N_20734,N_16119,N_17291);
xnor U20735 (N_20735,N_17272,N_17640);
and U20736 (N_20736,N_16560,N_16537);
nand U20737 (N_20737,N_16458,N_17615);
or U20738 (N_20738,N_16542,N_16315);
nor U20739 (N_20739,N_17094,N_16593);
or U20740 (N_20740,N_16457,N_17818);
xor U20741 (N_20741,N_17437,N_16834);
and U20742 (N_20742,N_17769,N_17922);
and U20743 (N_20743,N_15059,N_16473);
xor U20744 (N_20744,N_16368,N_16876);
or U20745 (N_20745,N_16525,N_15916);
and U20746 (N_20746,N_15785,N_16941);
nand U20747 (N_20747,N_17645,N_17108);
nand U20748 (N_20748,N_17478,N_17884);
or U20749 (N_20749,N_17115,N_15962);
nand U20750 (N_20750,N_17344,N_15031);
xnor U20751 (N_20751,N_17484,N_15505);
and U20752 (N_20752,N_15437,N_16508);
nand U20753 (N_20753,N_17582,N_15783);
nand U20754 (N_20754,N_16453,N_15445);
and U20755 (N_20755,N_17928,N_16941);
or U20756 (N_20756,N_17840,N_17398);
and U20757 (N_20757,N_15052,N_17889);
or U20758 (N_20758,N_17992,N_15777);
nor U20759 (N_20759,N_15455,N_15920);
and U20760 (N_20760,N_17384,N_15111);
xnor U20761 (N_20761,N_17421,N_15616);
xnor U20762 (N_20762,N_16246,N_17159);
nor U20763 (N_20763,N_17148,N_17852);
nand U20764 (N_20764,N_15322,N_16486);
nand U20765 (N_20765,N_15454,N_16566);
or U20766 (N_20766,N_15298,N_16802);
xor U20767 (N_20767,N_16692,N_16588);
xor U20768 (N_20768,N_16386,N_16148);
and U20769 (N_20769,N_16732,N_16526);
nor U20770 (N_20770,N_16210,N_17596);
nand U20771 (N_20771,N_15782,N_17491);
and U20772 (N_20772,N_15307,N_15050);
xnor U20773 (N_20773,N_17843,N_17784);
xor U20774 (N_20774,N_15478,N_15858);
or U20775 (N_20775,N_16206,N_15377);
nand U20776 (N_20776,N_17107,N_17794);
nor U20777 (N_20777,N_17907,N_15689);
nand U20778 (N_20778,N_16799,N_15759);
and U20779 (N_20779,N_17868,N_16680);
xor U20780 (N_20780,N_17348,N_17377);
nor U20781 (N_20781,N_17340,N_15973);
xnor U20782 (N_20782,N_16089,N_15042);
and U20783 (N_20783,N_16582,N_17509);
or U20784 (N_20784,N_16844,N_16382);
nand U20785 (N_20785,N_17626,N_15509);
and U20786 (N_20786,N_17859,N_15390);
or U20787 (N_20787,N_15233,N_17668);
or U20788 (N_20788,N_15779,N_16809);
nand U20789 (N_20789,N_17307,N_15906);
or U20790 (N_20790,N_16882,N_17409);
xor U20791 (N_20791,N_16329,N_17501);
nand U20792 (N_20792,N_17022,N_15444);
nor U20793 (N_20793,N_16431,N_17559);
or U20794 (N_20794,N_17816,N_15153);
xnor U20795 (N_20795,N_17830,N_15752);
and U20796 (N_20796,N_17285,N_16214);
nor U20797 (N_20797,N_17992,N_17115);
and U20798 (N_20798,N_16563,N_16930);
nor U20799 (N_20799,N_15821,N_16175);
xnor U20800 (N_20800,N_17267,N_15101);
nor U20801 (N_20801,N_15826,N_17907);
xor U20802 (N_20802,N_16150,N_16580);
xor U20803 (N_20803,N_16697,N_17136);
nor U20804 (N_20804,N_17539,N_17978);
nor U20805 (N_20805,N_15894,N_17453);
xor U20806 (N_20806,N_16157,N_15726);
or U20807 (N_20807,N_16711,N_15719);
and U20808 (N_20808,N_15486,N_17649);
xnor U20809 (N_20809,N_16437,N_15400);
nor U20810 (N_20810,N_15606,N_15203);
or U20811 (N_20811,N_16600,N_16268);
nand U20812 (N_20812,N_17417,N_16664);
xor U20813 (N_20813,N_17023,N_16275);
nand U20814 (N_20814,N_16120,N_16243);
nand U20815 (N_20815,N_15241,N_16771);
xnor U20816 (N_20816,N_15278,N_15510);
nand U20817 (N_20817,N_17320,N_17049);
or U20818 (N_20818,N_15587,N_17969);
nand U20819 (N_20819,N_17063,N_16230);
nand U20820 (N_20820,N_16126,N_15737);
xor U20821 (N_20821,N_15463,N_17230);
nor U20822 (N_20822,N_17560,N_17205);
nor U20823 (N_20823,N_15695,N_16049);
nor U20824 (N_20824,N_16900,N_16782);
xor U20825 (N_20825,N_16354,N_17986);
nand U20826 (N_20826,N_16323,N_16090);
nand U20827 (N_20827,N_15177,N_16099);
nor U20828 (N_20828,N_17975,N_17681);
and U20829 (N_20829,N_16395,N_16496);
and U20830 (N_20830,N_17839,N_15485);
nor U20831 (N_20831,N_15325,N_15381);
or U20832 (N_20832,N_16040,N_15258);
nand U20833 (N_20833,N_15158,N_16004);
and U20834 (N_20834,N_17691,N_15574);
and U20835 (N_20835,N_15852,N_16844);
nand U20836 (N_20836,N_16782,N_17368);
nor U20837 (N_20837,N_16589,N_17960);
or U20838 (N_20838,N_15061,N_17781);
nor U20839 (N_20839,N_17828,N_16698);
or U20840 (N_20840,N_17251,N_16228);
xnor U20841 (N_20841,N_15400,N_16152);
or U20842 (N_20842,N_15190,N_16593);
xnor U20843 (N_20843,N_16309,N_15984);
nor U20844 (N_20844,N_16217,N_16536);
nor U20845 (N_20845,N_16117,N_16203);
xor U20846 (N_20846,N_15455,N_17718);
or U20847 (N_20847,N_17476,N_16381);
xor U20848 (N_20848,N_17998,N_17381);
and U20849 (N_20849,N_17010,N_15596);
xor U20850 (N_20850,N_16254,N_15442);
or U20851 (N_20851,N_16382,N_16374);
and U20852 (N_20852,N_17240,N_17790);
and U20853 (N_20853,N_16634,N_15983);
and U20854 (N_20854,N_17172,N_16909);
xnor U20855 (N_20855,N_15155,N_16443);
or U20856 (N_20856,N_16317,N_17231);
nor U20857 (N_20857,N_15836,N_15919);
nand U20858 (N_20858,N_15323,N_15198);
and U20859 (N_20859,N_15289,N_16165);
nor U20860 (N_20860,N_17023,N_15057);
or U20861 (N_20861,N_15166,N_16983);
or U20862 (N_20862,N_15383,N_17234);
and U20863 (N_20863,N_17957,N_16039);
nand U20864 (N_20864,N_17401,N_17627);
or U20865 (N_20865,N_16190,N_16753);
nand U20866 (N_20866,N_16862,N_15380);
or U20867 (N_20867,N_16887,N_15164);
nor U20868 (N_20868,N_17247,N_15658);
or U20869 (N_20869,N_15159,N_16895);
xnor U20870 (N_20870,N_15575,N_15455);
xnor U20871 (N_20871,N_15292,N_15026);
nor U20872 (N_20872,N_17865,N_15600);
or U20873 (N_20873,N_15553,N_17260);
or U20874 (N_20874,N_16355,N_16112);
nand U20875 (N_20875,N_17020,N_15906);
or U20876 (N_20876,N_16381,N_16443);
or U20877 (N_20877,N_15281,N_15821);
nor U20878 (N_20878,N_15200,N_16395);
xnor U20879 (N_20879,N_17697,N_16497);
nor U20880 (N_20880,N_15893,N_17492);
xnor U20881 (N_20881,N_17143,N_16342);
nor U20882 (N_20882,N_17183,N_16460);
and U20883 (N_20883,N_17114,N_16887);
xnor U20884 (N_20884,N_16286,N_17532);
xnor U20885 (N_20885,N_17870,N_17115);
xor U20886 (N_20886,N_16273,N_17688);
or U20887 (N_20887,N_15335,N_15759);
or U20888 (N_20888,N_15363,N_15238);
and U20889 (N_20889,N_15940,N_16417);
nor U20890 (N_20890,N_17057,N_15609);
nor U20891 (N_20891,N_16376,N_16090);
or U20892 (N_20892,N_17746,N_15535);
and U20893 (N_20893,N_15806,N_17014);
xnor U20894 (N_20894,N_15084,N_16758);
and U20895 (N_20895,N_17309,N_17167);
or U20896 (N_20896,N_15917,N_15550);
or U20897 (N_20897,N_16670,N_17359);
and U20898 (N_20898,N_15572,N_17409);
and U20899 (N_20899,N_16469,N_16365);
or U20900 (N_20900,N_16243,N_17801);
or U20901 (N_20901,N_16637,N_16905);
and U20902 (N_20902,N_17948,N_15545);
nor U20903 (N_20903,N_16257,N_17504);
and U20904 (N_20904,N_15869,N_17841);
and U20905 (N_20905,N_16173,N_17124);
xnor U20906 (N_20906,N_17837,N_17160);
nand U20907 (N_20907,N_17922,N_17645);
nor U20908 (N_20908,N_15108,N_16124);
nor U20909 (N_20909,N_16798,N_17406);
xor U20910 (N_20910,N_16997,N_15632);
and U20911 (N_20911,N_15762,N_15864);
and U20912 (N_20912,N_16838,N_17525);
or U20913 (N_20913,N_16558,N_16847);
and U20914 (N_20914,N_17230,N_16957);
nor U20915 (N_20915,N_15258,N_16248);
nand U20916 (N_20916,N_17984,N_15827);
or U20917 (N_20917,N_16779,N_15574);
nand U20918 (N_20918,N_16848,N_15588);
or U20919 (N_20919,N_17320,N_16784);
nor U20920 (N_20920,N_16114,N_15290);
or U20921 (N_20921,N_17599,N_17186);
and U20922 (N_20922,N_15575,N_17922);
and U20923 (N_20923,N_15124,N_17929);
xor U20924 (N_20924,N_15809,N_17524);
or U20925 (N_20925,N_17654,N_15571);
xor U20926 (N_20926,N_16377,N_17162);
nor U20927 (N_20927,N_15574,N_15961);
or U20928 (N_20928,N_17769,N_16767);
nand U20929 (N_20929,N_15201,N_15588);
or U20930 (N_20930,N_17179,N_16778);
nand U20931 (N_20931,N_17813,N_16932);
xor U20932 (N_20932,N_17493,N_16852);
xor U20933 (N_20933,N_16628,N_15070);
nand U20934 (N_20934,N_16978,N_17432);
xnor U20935 (N_20935,N_15186,N_17128);
nor U20936 (N_20936,N_16448,N_16712);
nor U20937 (N_20937,N_16873,N_16644);
nand U20938 (N_20938,N_16321,N_17623);
and U20939 (N_20939,N_15108,N_16089);
nand U20940 (N_20940,N_15369,N_16520);
nand U20941 (N_20941,N_16811,N_17177);
xnor U20942 (N_20942,N_16815,N_16553);
nand U20943 (N_20943,N_15921,N_15409);
or U20944 (N_20944,N_15879,N_16665);
nand U20945 (N_20945,N_17275,N_15397);
xnor U20946 (N_20946,N_16833,N_17990);
or U20947 (N_20947,N_16544,N_16716);
nor U20948 (N_20948,N_16765,N_17650);
nand U20949 (N_20949,N_17153,N_16816);
xnor U20950 (N_20950,N_17460,N_17676);
nor U20951 (N_20951,N_16921,N_16667);
and U20952 (N_20952,N_17536,N_16376);
nand U20953 (N_20953,N_17903,N_16287);
nand U20954 (N_20954,N_17064,N_16552);
or U20955 (N_20955,N_17652,N_15349);
nand U20956 (N_20956,N_17404,N_17240);
nand U20957 (N_20957,N_16298,N_15084);
nor U20958 (N_20958,N_15496,N_17643);
nor U20959 (N_20959,N_15529,N_17771);
nor U20960 (N_20960,N_17380,N_16437);
and U20961 (N_20961,N_16607,N_15917);
nand U20962 (N_20962,N_17377,N_15901);
xor U20963 (N_20963,N_15284,N_17832);
xnor U20964 (N_20964,N_16266,N_17925);
nand U20965 (N_20965,N_15561,N_15633);
nand U20966 (N_20966,N_17008,N_17197);
and U20967 (N_20967,N_16417,N_15674);
or U20968 (N_20968,N_15401,N_16925);
nor U20969 (N_20969,N_16704,N_17021);
nand U20970 (N_20970,N_17555,N_15688);
xnor U20971 (N_20971,N_15733,N_16080);
or U20972 (N_20972,N_15407,N_15675);
and U20973 (N_20973,N_15741,N_15441);
nor U20974 (N_20974,N_17454,N_15287);
xor U20975 (N_20975,N_16165,N_15523);
and U20976 (N_20976,N_16290,N_15635);
nor U20977 (N_20977,N_16318,N_16466);
xor U20978 (N_20978,N_15952,N_16770);
xnor U20979 (N_20979,N_17288,N_15777);
or U20980 (N_20980,N_17955,N_15533);
nand U20981 (N_20981,N_17463,N_16981);
nor U20982 (N_20982,N_17650,N_16639);
or U20983 (N_20983,N_17741,N_15774);
and U20984 (N_20984,N_15928,N_15302);
xor U20985 (N_20985,N_17679,N_17034);
xnor U20986 (N_20986,N_16891,N_16854);
xnor U20987 (N_20987,N_15293,N_16785);
nand U20988 (N_20988,N_17324,N_15926);
and U20989 (N_20989,N_16052,N_17224);
xor U20990 (N_20990,N_17513,N_16011);
and U20991 (N_20991,N_15443,N_15183);
and U20992 (N_20992,N_17056,N_15558);
and U20993 (N_20993,N_17316,N_16520);
and U20994 (N_20994,N_17106,N_15036);
xnor U20995 (N_20995,N_17573,N_16580);
nor U20996 (N_20996,N_15453,N_15796);
or U20997 (N_20997,N_15992,N_17372);
or U20998 (N_20998,N_17965,N_17483);
or U20999 (N_20999,N_17818,N_17098);
and U21000 (N_21000,N_19708,N_18831);
nand U21001 (N_21001,N_20855,N_18123);
and U21002 (N_21002,N_18812,N_19563);
xnor U21003 (N_21003,N_19470,N_20360);
nor U21004 (N_21004,N_18363,N_18510);
nor U21005 (N_21005,N_19627,N_19087);
or U21006 (N_21006,N_19049,N_20807);
or U21007 (N_21007,N_19681,N_20796);
nand U21008 (N_21008,N_18302,N_18272);
nand U21009 (N_21009,N_20948,N_20954);
and U21010 (N_21010,N_19688,N_18059);
xor U21011 (N_21011,N_20291,N_19034);
nand U21012 (N_21012,N_20776,N_20862);
or U21013 (N_21013,N_18435,N_18460);
xnor U21014 (N_21014,N_20817,N_18707);
nor U21015 (N_21015,N_18754,N_20974);
and U21016 (N_21016,N_20980,N_20617);
nor U21017 (N_21017,N_18315,N_19959);
and U21018 (N_21018,N_19951,N_18336);
and U21019 (N_21019,N_19305,N_19985);
nand U21020 (N_21020,N_19668,N_20261);
nand U21021 (N_21021,N_19833,N_19099);
xor U21022 (N_21022,N_18883,N_18020);
or U21023 (N_21023,N_18457,N_20942);
and U21024 (N_21024,N_20663,N_18192);
nand U21025 (N_21025,N_20445,N_18456);
and U21026 (N_21026,N_20408,N_19780);
nand U21027 (N_21027,N_19020,N_20389);
or U21028 (N_21028,N_19726,N_20429);
and U21029 (N_21029,N_18865,N_20146);
nor U21030 (N_21030,N_18650,N_20368);
nand U21031 (N_21031,N_19878,N_19690);
xnor U21032 (N_21032,N_19743,N_18140);
or U21033 (N_21033,N_20475,N_19923);
xor U21034 (N_21034,N_18894,N_19716);
xnor U21035 (N_21035,N_19301,N_20101);
or U21036 (N_21036,N_19546,N_19801);
nand U21037 (N_21037,N_18601,N_20552);
xor U21038 (N_21038,N_19388,N_19033);
nand U21039 (N_21039,N_18830,N_20646);
or U21040 (N_21040,N_20941,N_18241);
xor U21041 (N_21041,N_20861,N_19530);
nor U21042 (N_21042,N_19151,N_19707);
or U21043 (N_21043,N_20875,N_20680);
or U21044 (N_21044,N_20238,N_19216);
nand U21045 (N_21045,N_18430,N_18277);
and U21046 (N_21046,N_18719,N_20791);
xor U21047 (N_21047,N_20359,N_19974);
or U21048 (N_21048,N_20905,N_18909);
nor U21049 (N_21049,N_18670,N_18109);
or U21050 (N_21050,N_19105,N_19129);
or U21051 (N_21051,N_19602,N_18347);
nand U21052 (N_21052,N_20844,N_19564);
or U21053 (N_21053,N_18455,N_19066);
nor U21054 (N_21054,N_19585,N_19746);
nand U21055 (N_21055,N_19313,N_19032);
nor U21056 (N_21056,N_18124,N_18847);
nor U21057 (N_21057,N_20433,N_20818);
and U21058 (N_21058,N_18502,N_20149);
nand U21059 (N_21059,N_19506,N_19336);
nor U21060 (N_21060,N_19767,N_19088);
or U21061 (N_21061,N_19758,N_19779);
xnor U21062 (N_21062,N_19050,N_20537);
nand U21063 (N_21063,N_19936,N_18944);
nand U21064 (N_21064,N_19064,N_20115);
xnor U21065 (N_21065,N_18688,N_18674);
xnor U21066 (N_21066,N_19760,N_20060);
nor U21067 (N_21067,N_19686,N_20309);
nand U21068 (N_21068,N_18032,N_18822);
or U21069 (N_21069,N_18580,N_20148);
nand U21070 (N_21070,N_18984,N_20381);
xnor U21071 (N_21071,N_20068,N_19499);
and U21072 (N_21072,N_20100,N_18704);
nand U21073 (N_21073,N_19244,N_19870);
nand U21074 (N_21074,N_18735,N_18423);
and U21075 (N_21075,N_20059,N_20836);
nor U21076 (N_21076,N_19278,N_19755);
or U21077 (N_21077,N_20850,N_18204);
xnor U21078 (N_21078,N_19132,N_19989);
and U21079 (N_21079,N_20521,N_18304);
xnor U21080 (N_21080,N_20724,N_19634);
and U21081 (N_21081,N_18266,N_18615);
nor U21082 (N_21082,N_20356,N_20332);
nor U21083 (N_21083,N_20456,N_20409);
nor U21084 (N_21084,N_20872,N_18721);
or U21085 (N_21085,N_19248,N_19826);
xnor U21086 (N_21086,N_20786,N_19000);
or U21087 (N_21087,N_19799,N_20026);
nor U21088 (N_21088,N_20588,N_19465);
and U21089 (N_21089,N_18904,N_18646);
nand U21090 (N_21090,N_19840,N_18669);
nor U21091 (N_21091,N_18742,N_19915);
or U21092 (N_21092,N_20928,N_18786);
and U21093 (N_21093,N_18999,N_19004);
and U21094 (N_21094,N_20548,N_18353);
or U21095 (N_21095,N_20930,N_19071);
and U21096 (N_21096,N_18112,N_20587);
or U21097 (N_21097,N_19102,N_18527);
xor U21098 (N_21098,N_19832,N_18949);
nor U21099 (N_21099,N_20853,N_20504);
and U21100 (N_21100,N_19392,N_20883);
and U21101 (N_21101,N_18872,N_19454);
xor U21102 (N_21102,N_18337,N_20625);
nor U21103 (N_21103,N_20438,N_20686);
and U21104 (N_21104,N_20420,N_20366);
and U21105 (N_21105,N_18235,N_18619);
nor U21106 (N_21106,N_19361,N_19992);
or U21107 (N_21107,N_19453,N_19447);
xnor U21108 (N_21108,N_19830,N_18198);
xnor U21109 (N_21109,N_20804,N_20347);
and U21110 (N_21110,N_19572,N_19558);
or U21111 (N_21111,N_19817,N_20185);
or U21112 (N_21112,N_20970,N_20214);
or U21113 (N_21113,N_19055,N_20211);
and U21114 (N_21114,N_20539,N_18273);
nor U21115 (N_21115,N_20119,N_20351);
and U21116 (N_21116,N_19661,N_18194);
or U21117 (N_21117,N_19471,N_19622);
or U21118 (N_21118,N_19256,N_19013);
and U21119 (N_21119,N_18325,N_20694);
xor U21120 (N_21120,N_18620,N_20890);
nor U21121 (N_21121,N_20832,N_18916);
nor U21122 (N_21122,N_19287,N_20803);
or U21123 (N_21123,N_20687,N_19252);
and U21124 (N_21124,N_19270,N_19773);
nand U21125 (N_21125,N_20303,N_19439);
nor U21126 (N_21126,N_19235,N_18495);
nand U21127 (N_21127,N_19551,N_19365);
or U21128 (N_21128,N_20150,N_20976);
nor U21129 (N_21129,N_19526,N_18932);
nor U21130 (N_21130,N_20428,N_18618);
xor U21131 (N_21131,N_18884,N_20708);
nand U21132 (N_21132,N_20337,N_18518);
nor U21133 (N_21133,N_19115,N_20221);
xor U21134 (N_21134,N_20056,N_20673);
xor U21135 (N_21135,N_19092,N_18038);
nand U21136 (N_21136,N_18714,N_18604);
nand U21137 (N_21137,N_18424,N_20006);
and U21138 (N_21138,N_18309,N_18230);
and U21139 (N_21139,N_19068,N_18401);
or U21140 (N_21140,N_19728,N_18534);
or U21141 (N_21141,N_19685,N_20017);
or U21142 (N_21142,N_19589,N_19180);
nor U21143 (N_21143,N_18757,N_18356);
and U21144 (N_21144,N_20851,N_20772);
or U21145 (N_21145,N_20121,N_18470);
xnor U21146 (N_21146,N_19560,N_18605);
nor U21147 (N_21147,N_18199,N_18159);
or U21148 (N_21148,N_20264,N_19474);
nor U21149 (N_21149,N_20493,N_18979);
nand U21150 (N_21150,N_19357,N_20446);
xor U21151 (N_21151,N_19583,N_18851);
or U21152 (N_21152,N_18323,N_18480);
or U21153 (N_21153,N_18092,N_18765);
nand U21154 (N_21154,N_19139,N_19397);
xor U21155 (N_21155,N_20518,N_20285);
xnor U21156 (N_21156,N_20506,N_20752);
nand U21157 (N_21157,N_18229,N_18095);
nand U21158 (N_21158,N_18240,N_20472);
or U21159 (N_21159,N_18049,N_18284);
nor U21160 (N_21160,N_19539,N_20234);
and U21161 (N_21161,N_18779,N_19842);
or U21162 (N_21162,N_19428,N_18511);
or U21163 (N_21163,N_19373,N_18803);
xor U21164 (N_21164,N_18209,N_20141);
xor U21165 (N_21165,N_19909,N_20959);
or U21166 (N_21166,N_20509,N_20384);
nor U21167 (N_21167,N_18611,N_19948);
or U21168 (N_21168,N_18813,N_18130);
or U21169 (N_21169,N_18770,N_18584);
nor U21170 (N_21170,N_18819,N_20527);
and U21171 (N_21171,N_18000,N_18683);
or U21172 (N_21172,N_20681,N_19623);
and U21173 (N_21173,N_20206,N_20714);
or U21174 (N_21174,N_19926,N_19429);
nand U21175 (N_21175,N_18835,N_19663);
nand U21176 (N_21176,N_19885,N_18799);
nand U21177 (N_21177,N_20816,N_18278);
xnor U21178 (N_21178,N_19666,N_19512);
and U21179 (N_21179,N_19215,N_19326);
nand U21180 (N_21180,N_20029,N_20399);
nand U21181 (N_21181,N_18689,N_19884);
nor U21182 (N_21182,N_18778,N_19605);
xor U21183 (N_21183,N_18982,N_20645);
xnor U21184 (N_21184,N_18343,N_18661);
or U21185 (N_21185,N_20375,N_20175);
nor U21186 (N_21186,N_19770,N_19073);
and U21187 (N_21187,N_20186,N_19754);
and U21188 (N_21188,N_19944,N_18355);
nor U21189 (N_21189,N_20835,N_20674);
nor U21190 (N_21190,N_19983,N_19147);
and U21191 (N_21191,N_18562,N_20296);
nand U21192 (N_21192,N_18482,N_18216);
nand U21193 (N_21193,N_19440,N_18785);
or U21194 (N_21194,N_20131,N_18559);
nor U21195 (N_21195,N_20734,N_19442);
nand U21196 (N_21196,N_20626,N_18163);
or U21197 (N_21197,N_20725,N_20333);
or U21198 (N_21198,N_18113,N_20658);
nand U21199 (N_21199,N_18221,N_20897);
nor U21200 (N_21200,N_19054,N_19127);
and U21201 (N_21201,N_19435,N_20720);
and U21202 (N_21202,N_19500,N_20642);
xnor U21203 (N_21203,N_19396,N_19929);
nor U21204 (N_21204,N_20372,N_18964);
nor U21205 (N_21205,N_19402,N_20120);
or U21206 (N_21206,N_18342,N_18839);
or U21207 (N_21207,N_20287,N_20876);
nor U21208 (N_21208,N_19269,N_20641);
and U21209 (N_21209,N_20729,N_20018);
and U21210 (N_21210,N_19881,N_19199);
xor U21211 (N_21211,N_20797,N_19810);
xnor U21212 (N_21212,N_19192,N_19364);
xnor U21213 (N_21213,N_20094,N_20917);
xnor U21214 (N_21214,N_20723,N_20397);
or U21215 (N_21215,N_19721,N_19953);
nor U21216 (N_21216,N_20099,N_18723);
or U21217 (N_21217,N_19279,N_20412);
or U21218 (N_21218,N_20595,N_20022);
xor U21219 (N_21219,N_19818,N_20089);
xor U21220 (N_21220,N_18657,N_18598);
nor U21221 (N_21221,N_20893,N_19375);
and U21222 (N_21222,N_18500,N_18115);
xnor U21223 (N_21223,N_19108,N_18525);
and U21224 (N_21224,N_20700,N_20302);
xnor U21225 (N_21225,N_18409,N_19718);
nor U21226 (N_21226,N_20608,N_19616);
xor U21227 (N_21227,N_19460,N_19785);
and U21228 (N_21228,N_18264,N_18174);
nand U21229 (N_21229,N_20448,N_20699);
nor U21230 (N_21230,N_19290,N_19993);
nand U21231 (N_21231,N_18655,N_18530);
and U21232 (N_21232,N_18026,N_19395);
or U21233 (N_21233,N_20127,N_19224);
and U21234 (N_21234,N_20469,N_18191);
xnor U21235 (N_21235,N_18826,N_20480);
and U21236 (N_21236,N_18673,N_18232);
nor U21237 (N_21237,N_18003,N_20317);
nand U21238 (N_21238,N_18696,N_18665);
and U21239 (N_21239,N_19712,N_19237);
nand U21240 (N_21240,N_20961,N_20039);
and U21241 (N_21241,N_18952,N_19709);
nor U21242 (N_21242,N_18733,N_19384);
nor U21243 (N_21243,N_20001,N_18295);
and U21244 (N_21244,N_18989,N_18705);
nand U21245 (N_21245,N_19965,N_18906);
or U21246 (N_21246,N_20993,N_19537);
xor U21247 (N_21247,N_18781,N_18552);
xor U21248 (N_21248,N_20852,N_19360);
and U21249 (N_21249,N_18042,N_18196);
nor U21250 (N_21250,N_19731,N_20111);
and U21251 (N_21251,N_19677,N_18561);
and U21252 (N_21252,N_20972,N_19413);
and U21253 (N_21253,N_20262,N_18535);
or U21254 (N_21254,N_19484,N_18352);
and U21255 (N_21255,N_20338,N_18545);
nor U21256 (N_21256,N_20889,N_19593);
xor U21257 (N_21257,N_20170,N_19625);
or U21258 (N_21258,N_18971,N_18748);
and U21259 (N_21259,N_18951,N_19696);
or U21260 (N_21260,N_19640,N_19489);
nor U21261 (N_21261,N_19816,N_18182);
or U21262 (N_21262,N_19084,N_19964);
or U21263 (N_21263,N_19424,N_19587);
xor U21264 (N_21264,N_19378,N_20664);
and U21265 (N_21265,N_18311,N_20934);
nand U21266 (N_21266,N_20500,N_18980);
and U21267 (N_21267,N_19538,N_19138);
xnor U21268 (N_21268,N_18672,N_18255);
xnor U21269 (N_21269,N_18052,N_19655);
xnor U21270 (N_21270,N_20147,N_18992);
or U21271 (N_21271,N_20744,N_20757);
and U21272 (N_21272,N_20873,N_18616);
nor U21273 (N_21273,N_18947,N_20478);
or U21274 (N_21274,N_19877,N_18149);
and U21275 (N_21275,N_19880,N_20432);
xor U21276 (N_21276,N_20132,N_19608);
or U21277 (N_21277,N_18606,N_18887);
nor U21278 (N_21278,N_20837,N_20682);
and U21279 (N_21279,N_20055,N_19186);
nor U21280 (N_21280,N_19463,N_19350);
or U21281 (N_21281,N_20114,N_19701);
nor U21282 (N_21282,N_20016,N_18419);
and U21283 (N_21283,N_18730,N_18184);
or U21284 (N_21284,N_18231,N_18823);
nand U21285 (N_21285,N_20668,N_19698);
or U21286 (N_21286,N_18567,N_18633);
and U21287 (N_21287,N_18860,N_20095);
nand U21288 (N_21288,N_18102,N_19981);
or U21289 (N_21289,N_20799,N_20604);
nand U21290 (N_21290,N_20410,N_18166);
nor U21291 (N_21291,N_20679,N_19824);
xnor U21292 (N_21292,N_18108,N_19838);
nor U21293 (N_21293,N_19492,N_20449);
and U21294 (N_21294,N_20161,N_20011);
nand U21295 (N_21295,N_19568,N_19042);
xor U21296 (N_21296,N_20065,N_19807);
nor U21297 (N_21297,N_18399,N_18802);
or U21298 (N_21298,N_20224,N_18051);
nor U21299 (N_21299,N_19120,N_19204);
nor U21300 (N_21300,N_19897,N_19014);
xor U21301 (N_21301,N_19477,N_18837);
and U21302 (N_21302,N_18806,N_20345);
and U21303 (N_21303,N_20907,N_20485);
or U21304 (N_21304,N_20035,N_20415);
nor U21305 (N_21305,N_18950,N_20722);
nor U21306 (N_21306,N_18339,N_20774);
nand U21307 (N_21307,N_18529,N_20675);
and U21308 (N_21308,N_18918,N_19565);
or U21309 (N_21309,N_18481,N_18054);
xnor U21310 (N_21310,N_19994,N_18316);
nor U21311 (N_21311,N_19058,N_18886);
xor U21312 (N_21312,N_18555,N_18469);
xor U21313 (N_21313,N_20042,N_19241);
or U21314 (N_21314,N_18538,N_20981);
xor U21315 (N_21315,N_18465,N_20257);
xor U21316 (N_21316,N_20193,N_18997);
or U21317 (N_21317,N_18248,N_18553);
or U21318 (N_21318,N_19719,N_20632);
and U21319 (N_21319,N_19191,N_18087);
nand U21320 (N_21320,N_18970,N_20582);
or U21321 (N_21321,N_18760,N_18675);
xnor U21322 (N_21322,N_20159,N_18647);
nand U21323 (N_21323,N_20323,N_18953);
nor U21324 (N_21324,N_18321,N_18642);
nand U21325 (N_21325,N_18514,N_18797);
or U21326 (N_21326,N_19511,N_18946);
nand U21327 (N_21327,N_19096,N_19534);
or U21328 (N_21328,N_20209,N_18846);
nor U21329 (N_21329,N_18899,N_20887);
or U21330 (N_21330,N_19910,N_20436);
xor U21331 (N_21331,N_19200,N_20598);
nor U21332 (N_21332,N_19906,N_20523);
xor U21333 (N_21333,N_20484,N_20010);
nand U21334 (N_21334,N_18348,N_18549);
xor U21335 (N_21335,N_20310,N_20488);
nor U21336 (N_21336,N_19418,N_18210);
and U21337 (N_21337,N_18712,N_20922);
nand U21338 (N_21338,N_19660,N_20716);
or U21339 (N_21339,N_19464,N_20874);
xnor U21340 (N_21340,N_19434,N_18445);
xnor U21341 (N_21341,N_19161,N_19829);
or U21342 (N_21342,N_18002,N_20594);
nor U21343 (N_21343,N_19822,N_19706);
and U21344 (N_21344,N_18156,N_19069);
nor U21345 (N_21345,N_20584,N_18239);
xnor U21346 (N_21346,N_19750,N_20986);
nor U21347 (N_21347,N_18041,N_20142);
xnor U21348 (N_21348,N_20076,N_18522);
nand U21349 (N_21349,N_20777,N_18226);
and U21350 (N_21350,N_20104,N_19561);
xnor U21351 (N_21351,N_19043,N_19643);
xnor U21352 (N_21352,N_19740,N_20268);
xnor U21353 (N_21353,N_20203,N_19871);
and U21354 (N_21354,N_19514,N_20705);
or U21355 (N_21355,N_19520,N_18701);
and U21356 (N_21356,N_20913,N_19732);
or U21357 (N_21357,N_20294,N_18082);
xor U21358 (N_21358,N_18681,N_20657);
nand U21359 (N_21359,N_18022,N_19242);
or U21360 (N_21360,N_18013,N_19255);
xnor U21361 (N_21361,N_18211,N_18274);
or U21362 (N_21362,N_18991,N_20929);
xor U21363 (N_21363,N_19575,N_20812);
or U21364 (N_21364,N_20847,N_20854);
nand U21365 (N_21365,N_19697,N_19059);
nand U21366 (N_21366,N_18039,N_19497);
xnor U21367 (N_21367,N_18526,N_19346);
xor U21368 (N_21368,N_18298,N_18033);
and U21369 (N_21369,N_20763,N_19788);
xnor U21370 (N_21370,N_18876,N_18137);
xor U21371 (N_21371,N_18722,N_18296);
and U21372 (N_21372,N_19552,N_18357);
or U21373 (N_21373,N_20540,N_20355);
nand U21374 (N_21374,N_20692,N_19580);
xor U21375 (N_21375,N_20983,N_19104);
or U21376 (N_21376,N_18859,N_19286);
nand U21377 (N_21377,N_19918,N_18475);
xnor U21378 (N_21378,N_19662,N_20053);
xnor U21379 (N_21379,N_20163,N_18116);
nand U21380 (N_21380,N_18310,N_20513);
xor U21381 (N_21381,N_20260,N_18055);
or U21382 (N_21382,N_19293,N_19813);
nand U21383 (N_21383,N_18697,N_18004);
or U21384 (N_21384,N_20609,N_19607);
xnor U21385 (N_21385,N_20858,N_18824);
and U21386 (N_21386,N_18708,N_20492);
nand U21387 (N_21387,N_19430,N_19012);
or U21388 (N_21388,N_20395,N_18270);
or U21389 (N_21389,N_20762,N_18738);
nand U21390 (N_21390,N_19341,N_20487);
or U21391 (N_21391,N_19462,N_19179);
or U21392 (N_21392,N_18663,N_19521);
nor U21393 (N_21393,N_20314,N_20201);
and U21394 (N_21394,N_18061,N_18252);
or U21395 (N_21395,N_20027,N_19815);
nand U21396 (N_21396,N_18888,N_18957);
and U21397 (N_21397,N_20087,N_20256);
nand U21398 (N_21398,N_19030,N_18570);
xnor U21399 (N_21399,N_20025,N_18983);
nand U21400 (N_21400,N_18850,N_18008);
and U21401 (N_21401,N_18063,N_19029);
nand U21402 (N_21402,N_20107,N_18073);
or U21403 (N_21403,N_18364,N_18990);
xnor U21404 (N_21404,N_19163,N_20550);
xnor U21405 (N_21405,N_19933,N_18256);
nor U21406 (N_21406,N_19995,N_19991);
nand U21407 (N_21407,N_19831,N_19942);
xnor U21408 (N_21408,N_19901,N_20184);
nor U21409 (N_21409,N_19232,N_19727);
xnor U21410 (N_21410,N_19808,N_20770);
nand U21411 (N_21411,N_20813,N_19914);
and U21412 (N_21412,N_19040,N_20299);
nor U21413 (N_21413,N_18064,N_20322);
nor U21414 (N_21414,N_20339,N_19382);
and U21415 (N_21415,N_18144,N_19896);
and U21416 (N_21416,N_20290,N_18384);
or U21417 (N_21417,N_19264,N_18703);
xor U21418 (N_21418,N_18926,N_19063);
or U21419 (N_21419,N_19544,N_20557);
xor U21420 (N_21420,N_20721,N_18623);
and U21421 (N_21421,N_18843,N_18154);
or U21422 (N_21422,N_18940,N_19372);
xor U21423 (N_21423,N_19312,N_18820);
nor U21424 (N_21424,N_19028,N_20881);
and U21425 (N_21425,N_19854,N_19422);
nand U21426 (N_21426,N_18282,N_18692);
and U21427 (N_21427,N_19786,N_20283);
nor U21428 (N_21428,N_19271,N_18603);
xnor U21429 (N_21429,N_19090,N_18869);
xnor U21430 (N_21430,N_19285,N_20794);
xnor U21431 (N_21431,N_20482,N_20180);
nand U21432 (N_21432,N_19021,N_20621);
nor U21433 (N_21433,N_18658,N_19672);
nand U21434 (N_21434,N_18898,N_19776);
nand U21435 (N_21435,N_18973,N_18471);
nor U21436 (N_21436,N_19864,N_20849);
xnor U21437 (N_21437,N_20536,N_18297);
and U21438 (N_21438,N_19749,N_19174);
xnor U21439 (N_21439,N_19130,N_20977);
xnor U21440 (N_21440,N_18333,N_18105);
or U21441 (N_21441,N_20319,N_18845);
and U21442 (N_21442,N_19140,N_18128);
nand U21443 (N_21443,N_20885,N_20965);
nor U21444 (N_21444,N_18582,N_20926);
or U21445 (N_21445,N_19579,N_19855);
and U21446 (N_21446,N_18043,N_18120);
and U21447 (N_21447,N_18023,N_18494);
or U21448 (N_21448,N_20181,N_18414);
or U21449 (N_21449,N_20033,N_20864);
or U21450 (N_21450,N_20407,N_19053);
and U21451 (N_21451,N_19142,N_19631);
or U21452 (N_21452,N_20130,N_19062);
or U21453 (N_21453,N_19651,N_20739);
nor U21454 (N_21454,N_20624,N_20247);
nand U21455 (N_21455,N_20566,N_20108);
nand U21456 (N_21456,N_18010,N_18801);
nor U21457 (N_21457,N_20457,N_19190);
and U21458 (N_21458,N_19737,N_19343);
or U21459 (N_21459,N_20671,N_18548);
nand U21460 (N_21460,N_18662,N_19282);
and U21461 (N_21461,N_19937,N_19005);
or U21462 (N_21462,N_18463,N_19766);
or U21463 (N_21463,N_20019,N_19611);
and U21464 (N_21464,N_18451,N_18879);
or U21465 (N_21465,N_19761,N_19052);
or U21466 (N_21466,N_18132,N_20097);
xor U21467 (N_21467,N_18744,N_20191);
nor U21468 (N_21468,N_20473,N_18237);
xor U21469 (N_21469,N_20070,N_20467);
nor U21470 (N_21470,N_18736,N_19695);
xnor U21471 (N_21471,N_19452,N_18461);
and U21472 (N_21472,N_20988,N_20301);
nor U21473 (N_21473,N_19924,N_20622);
or U21474 (N_21474,N_19863,N_20075);
nand U21475 (N_21475,N_18516,N_20088);
xnor U21476 (N_21476,N_19763,N_18448);
nand U21477 (N_21477,N_19480,N_18262);
and U21478 (N_21478,N_20508,N_19874);
or U21479 (N_21479,N_18981,N_18976);
or U21480 (N_21480,N_18224,N_19898);
nand U21481 (N_21481,N_20041,N_20713);
xor U21482 (N_21482,N_19988,N_19851);
xnor U21483 (N_21483,N_20020,N_18581);
nand U21484 (N_21484,N_20547,N_20568);
or U21485 (N_21485,N_19239,N_18094);
nor U21486 (N_21486,N_20569,N_20602);
nand U21487 (N_21487,N_20304,N_20447);
nor U21488 (N_21488,N_19400,N_18126);
or U21489 (N_21489,N_20960,N_19201);
xor U21490 (N_21490,N_18147,N_20249);
and U21491 (N_21491,N_20628,N_20396);
or U21492 (N_21492,N_18720,N_18713);
and U21493 (N_21493,N_18878,N_19665);
or U21494 (N_21494,N_20440,N_18597);
nand U21495 (N_21495,N_20023,N_19610);
nor U21496 (N_21496,N_20280,N_19516);
and U21497 (N_21497,N_20870,N_18157);
nor U21498 (N_21498,N_19504,N_19950);
xor U21499 (N_21499,N_19019,N_20902);
or U21500 (N_21500,N_19711,N_18206);
or U21501 (N_21501,N_19230,N_20217);
nand U21502 (N_21502,N_19876,N_20884);
nand U21503 (N_21503,N_18575,N_20819);
nor U21504 (N_21504,N_19405,N_19868);
xor U21505 (N_21505,N_20049,N_19448);
nor U21506 (N_21506,N_19389,N_18978);
and U21507 (N_21507,N_19074,N_19211);
nand U21508 (N_21508,N_19258,N_18626);
nand U21509 (N_21509,N_19917,N_20455);
nor U21510 (N_21510,N_18833,N_19214);
nor U21511 (N_21511,N_19652,N_19249);
nor U21512 (N_21512,N_19307,N_18577);
nand U21513 (N_21513,N_19381,N_20576);
and U21514 (N_21514,N_18691,N_20524);
nor U21515 (N_21515,N_18135,N_20514);
nor U21516 (N_21516,N_18375,N_20554);
xor U21517 (N_21517,N_20778,N_20559);
and U21518 (N_21518,N_18501,N_18397);
nand U21519 (N_21519,N_20685,N_19753);
and U21520 (N_21520,N_20189,N_19912);
or U21521 (N_21521,N_20753,N_19802);
nand U21522 (N_21522,N_19152,N_20112);
xor U21523 (N_21523,N_20899,N_19450);
and U21524 (N_21524,N_19800,N_19086);
nor U21525 (N_21525,N_20556,N_20510);
nand U21526 (N_21526,N_19212,N_20666);
nor U21527 (N_21527,N_18328,N_20958);
nand U21528 (N_21528,N_19184,N_20834);
nand U21529 (N_21529,N_20240,N_18016);
and U21530 (N_21530,N_20908,N_20005);
xnor U21531 (N_21531,N_18866,N_18070);
xor U21532 (N_21532,N_18287,N_20801);
and U21533 (N_21533,N_20570,N_19535);
or U21534 (N_21534,N_18508,N_19003);
nand U21535 (N_21535,N_18308,N_20940);
nand U21536 (N_21536,N_19476,N_18929);
nand U21537 (N_21537,N_20982,N_18622);
xor U21538 (N_21538,N_18727,N_20935);
or U21539 (N_21539,N_18260,N_18617);
or U21540 (N_21540,N_20665,N_20865);
nand U21541 (N_21541,N_18168,N_20200);
nor U21542 (N_21542,N_18777,N_18400);
nor U21543 (N_21543,N_20627,N_19172);
and U21544 (N_21544,N_19782,N_18560);
and U21545 (N_21545,N_18687,N_19649);
xor U21546 (N_21546,N_19218,N_20305);
and U21547 (N_21547,N_19836,N_18875);
nand U21548 (N_21548,N_20241,N_20458);
nor U21549 (N_21549,N_19016,N_20392);
xnor U21550 (N_21550,N_20468,N_19518);
and U21551 (N_21551,N_20466,N_19189);
xor U21552 (N_21552,N_19233,N_19206);
or U21553 (N_21553,N_18236,N_19469);
nor U21554 (N_21554,N_19496,N_18630);
xor U21555 (N_21555,N_19067,N_19545);
nor U21556 (N_21556,N_18732,N_20670);
nand U21557 (N_21557,N_20346,N_18450);
or U21558 (N_21558,N_18504,N_19328);
and U21559 (N_21559,N_20096,N_19205);
xor U21560 (N_21560,N_19134,N_19911);
nand U21561 (N_21561,N_18499,N_18935);
nor U21562 (N_21562,N_18519,N_20971);
nor U21563 (N_21563,N_19531,N_20698);
and U21564 (N_21564,N_20340,N_20605);
xor U21565 (N_21565,N_20943,N_18773);
and U21566 (N_21566,N_19494,N_19303);
and U21567 (N_21567,N_18425,N_20950);
or U21568 (N_21568,N_18954,N_19723);
or U21569 (N_21569,N_18217,N_19619);
and U21570 (N_21570,N_20078,N_18053);
xnor U21571 (N_21571,N_18195,N_20952);
and U21572 (N_21572,N_19493,N_18709);
nor U21573 (N_21573,N_19198,N_18706);
and U21574 (N_21574,N_19458,N_20773);
nor U21575 (N_21575,N_18180,N_20585);
nor U21576 (N_21576,N_18873,N_20422);
or U21577 (N_21577,N_19292,N_20382);
xor U21578 (N_21578,N_18923,N_19508);
and U21579 (N_21579,N_18269,N_18011);
nand U21580 (N_21580,N_19300,N_20640);
or U21581 (N_21581,N_18173,N_20411);
and U21582 (N_21582,N_19943,N_20168);
nor U21583 (N_21583,N_18171,N_19722);
nand U21584 (N_21584,N_19347,N_20610);
xnor U21585 (N_21585,N_20750,N_18864);
xor U21586 (N_21586,N_18222,N_19883);
nand U21587 (N_21587,N_19812,N_19687);
nand U21588 (N_21588,N_18868,N_19693);
nor U21589 (N_21589,N_18208,N_19986);
xnor U21590 (N_21590,N_18246,N_18200);
or U21591 (N_21591,N_18855,N_18145);
nand U21592 (N_21592,N_18651,N_19907);
and U21593 (N_21593,N_18852,N_18551);
and U21594 (N_21594,N_18391,N_18076);
nand U21595 (N_21595,N_20780,N_18825);
or U21596 (N_21596,N_19441,N_18203);
or U21597 (N_21597,N_20354,N_19963);
nand U21598 (N_21598,N_19247,N_18268);
and U21599 (N_21599,N_18569,N_19008);
nor U21600 (N_21600,N_18573,N_19419);
and U21601 (N_21601,N_20140,N_18117);
or U21602 (N_21602,N_20424,N_19135);
or U21603 (N_21603,N_19805,N_19353);
nand U21604 (N_21604,N_19945,N_20306);
nor U21605 (N_21605,N_20113,N_20737);
nand U21606 (N_21606,N_18065,N_19730);
nand U21607 (N_21607,N_20215,N_18305);
nor U21608 (N_21608,N_18679,N_19315);
nand U21609 (N_21609,N_18690,N_20430);
and U21610 (N_21610,N_18726,N_18739);
nand U21611 (N_21611,N_20233,N_18125);
nor U21612 (N_21612,N_20442,N_18446);
nor U21613 (N_21613,N_19960,N_18856);
or U21614 (N_21614,N_18496,N_20158);
or U21615 (N_21615,N_20174,N_19796);
nand U21616 (N_21616,N_19423,N_18093);
and U21617 (N_21617,N_18406,N_19036);
nor U21618 (N_21618,N_20073,N_20906);
nor U21619 (N_21619,N_19524,N_19488);
and U21620 (N_21620,N_18816,N_18871);
and U21621 (N_21621,N_19949,N_19436);
nor U21622 (N_21622,N_20204,N_19632);
xnor U21623 (N_21623,N_20342,N_19207);
nor U21624 (N_21624,N_20654,N_19768);
xnor U21625 (N_21625,N_19107,N_18452);
and U21626 (N_21626,N_19051,N_19540);
nand U21627 (N_21627,N_20079,N_18808);
and U21628 (N_21628,N_18121,N_18503);
and U21629 (N_21629,N_18741,N_20678);
nand U21630 (N_21630,N_20549,N_20297);
nand U21631 (N_21631,N_19678,N_19111);
nand U21632 (N_21632,N_19717,N_19203);
xor U21633 (N_21633,N_20009,N_18426);
and U21634 (N_21634,N_18885,N_18119);
nor U21635 (N_21635,N_20530,N_20307);
or U21636 (N_21636,N_18827,N_18238);
nor U21637 (N_21637,N_20116,N_19969);
and U21638 (N_21638,N_18286,N_19956);
or U21639 (N_21639,N_20901,N_20028);
nor U21640 (N_21640,N_18212,N_18842);
or U21641 (N_21641,N_19759,N_19363);
nand U21642 (N_21642,N_20197,N_18447);
and U21643 (N_21643,N_19329,N_20134);
and U21644 (N_21644,N_20927,N_19890);
nor U21645 (N_21645,N_20995,N_20754);
xor U21646 (N_21646,N_19574,N_19437);
and U21647 (N_21647,N_20086,N_20519);
or U21648 (N_21648,N_19112,N_18299);
xor U21649 (N_21649,N_19426,N_19866);
or U21650 (N_21650,N_18228,N_18543);
xnor U21651 (N_21651,N_19939,N_19903);
nor U21652 (N_21652,N_18901,N_18832);
nand U21653 (N_21653,N_19962,N_19284);
xor U21654 (N_21654,N_20949,N_18919);
nor U21655 (N_21655,N_20898,N_20643);
nand U21656 (N_21656,N_19570,N_18922);
nor U21657 (N_21657,N_18639,N_18034);
nand U21658 (N_21658,N_18218,N_19653);
xor U21659 (N_21659,N_19354,N_18249);
or U21660 (N_21660,N_19837,N_20071);
nand U21661 (N_21661,N_18533,N_18386);
and U21662 (N_21662,N_20701,N_18454);
nor U21663 (N_21663,N_18939,N_18634);
or U21664 (N_21664,N_20903,N_20840);
nor U21665 (N_21665,N_18595,N_20045);
and U21666 (N_21666,N_20984,N_18882);
xor U21667 (N_21667,N_19443,N_19569);
nand U21668 (N_21668,N_20072,N_18702);
or U21669 (N_21669,N_18060,N_20543);
nor U21670 (N_21670,N_18334,N_19340);
or U21671 (N_21671,N_19057,N_18390);
nand U21672 (N_21672,N_18749,N_20178);
or U21673 (N_21673,N_19259,N_19356);
xor U21674 (N_21674,N_20000,N_20782);
and U21675 (N_21675,N_20656,N_19629);
and U21676 (N_21676,N_20669,N_19861);
nor U21677 (N_21677,N_19362,N_20607);
and U21678 (N_21678,N_18574,N_19277);
or U21679 (N_21679,N_18961,N_19961);
nor U21680 (N_21680,N_20118,N_19416);
xnor U21681 (N_21681,N_20109,N_19345);
and U21682 (N_21682,N_18589,N_19860);
nand U21683 (N_21683,N_18540,N_19635);
xor U21684 (N_21684,N_19809,N_20318);
nand U21685 (N_21685,N_19338,N_20597);
nand U21686 (N_21686,N_19451,N_18912);
or U21687 (N_21687,N_18127,N_18288);
and U21688 (N_21688,N_18213,N_19185);
nand U21689 (N_21689,N_20683,N_19221);
nand U21690 (N_21690,N_19240,N_18664);
or U21691 (N_21691,N_18443,N_18058);
nand U21692 (N_21692,N_19751,N_19618);
or U21693 (N_21693,N_19324,N_18924);
and U21694 (N_21694,N_20464,N_19849);
xnor U21695 (N_21695,N_20593,N_18012);
nor U21696 (N_21696,N_19257,N_20697);
and U21697 (N_21697,N_18332,N_20315);
nand U21698 (N_21698,N_19641,N_20474);
or U21699 (N_21699,N_19156,N_20047);
nor U21700 (N_21700,N_20560,N_20957);
nand U21701 (N_21701,N_20371,N_18969);
or U21702 (N_21702,N_19321,N_19024);
and U21703 (N_21703,N_19957,N_20343);
nor U21704 (N_21704,N_18367,N_19713);
nor U21705 (N_21705,N_20008,N_20894);
or U21706 (N_21706,N_18118,N_20541);
and U21707 (N_21707,N_20270,N_19010);
or U21708 (N_21708,N_18596,N_18388);
nand U21709 (N_21709,N_18484,N_18358);
xnor U21710 (N_21710,N_20459,N_20591);
nor U21711 (N_21711,N_20994,N_20123);
nor U21712 (N_21712,N_18294,N_18258);
nor U21713 (N_21713,N_20208,N_19852);
nor U21714 (N_21714,N_18244,N_18539);
nand U21715 (N_21715,N_20789,N_18190);
nor U21716 (N_21716,N_20373,N_19578);
xor U21717 (N_21717,N_19757,N_20501);
xor U21718 (N_21718,N_20848,N_20098);
or U21719 (N_21719,N_18750,N_19916);
nand U21720 (N_21720,N_18377,N_19922);
xnor U21721 (N_21721,N_20978,N_20745);
xor U21722 (N_21722,N_18069,N_18572);
and U21723 (N_21723,N_19314,N_19376);
nand U21724 (N_21724,N_20759,N_19410);
nor U21725 (N_21725,N_19947,N_20612);
nor U21726 (N_21726,N_20213,N_18766);
nor U21727 (N_21727,N_18737,N_20316);
or U21728 (N_21728,N_20499,N_20615);
or U21729 (N_21729,N_19299,N_19609);
xnor U21730 (N_21730,N_18627,N_19853);
xor U21731 (N_21731,N_18433,N_19900);
xor U21732 (N_21732,N_18769,N_20599);
nand U21733 (N_21733,N_20188,N_20538);
nand U21734 (N_21734,N_19082,N_19586);
nor U21735 (N_21735,N_20361,N_18660);
xnor U21736 (N_21736,N_20122,N_18458);
nor U21737 (N_21737,N_19330,N_18546);
nor U21738 (N_21738,N_18635,N_20202);
xnor U21739 (N_21739,N_20173,N_18700);
and U21740 (N_21740,N_20574,N_19846);
nor U21741 (N_21741,N_19065,N_18488);
nand U21742 (N_21742,N_20516,N_19094);
or U21743 (N_21743,N_19674,N_20243);
xnor U21744 (N_21744,N_20169,N_19035);
and U21745 (N_21745,N_19208,N_18996);
nor U21746 (N_21746,N_19041,N_20512);
or U21747 (N_21747,N_20255,N_20775);
nand U21748 (N_21748,N_19715,N_18587);
or U21749 (N_21749,N_19902,N_18892);
nand U21750 (N_21750,N_19188,N_18437);
nand U21751 (N_21751,N_18275,N_19821);
nor U21752 (N_21752,N_20502,N_19882);
xor U21753 (N_21753,N_20401,N_18745);
nand U21754 (N_21754,N_20369,N_20718);
xnor U21755 (N_21755,N_18403,N_18592);
nand U21756 (N_21756,N_20660,N_18654);
xnor U21757 (N_21757,N_20827,N_19291);
and U21758 (N_21758,N_18276,N_18815);
or U21759 (N_21759,N_20914,N_19283);
nor U21760 (N_21760,N_18136,N_20962);
and U21761 (N_21761,N_19975,N_18207);
or U21762 (N_21762,N_19752,N_20082);
and U21763 (N_21763,N_19173,N_18479);
and U21764 (N_21764,N_18960,N_19348);
and U21765 (N_21765,N_20564,N_20761);
nor U21766 (N_21766,N_20793,N_20945);
xor U21767 (N_21767,N_18591,N_20324);
and U21768 (N_21768,N_18751,N_18734);
xor U21769 (N_21769,N_20644,N_20278);
xnor U21770 (N_21770,N_18994,N_19085);
nor U21771 (N_21771,N_20335,N_20038);
or U21772 (N_21772,N_18853,N_18318);
and U21773 (N_21773,N_19848,N_19979);
or U21774 (N_21774,N_19409,N_18931);
nor U21775 (N_21775,N_20871,N_20768);
or U21776 (N_21776,N_18523,N_20805);
and U21777 (N_21777,N_18775,N_19525);
or U21778 (N_21778,N_18131,N_19980);
nand U21779 (N_21779,N_20491,N_18018);
nand U21780 (N_21780,N_20784,N_18279);
and U21781 (N_21781,N_19160,N_18331);
nand U21782 (N_21782,N_20600,N_19263);
or U21783 (N_21783,N_19072,N_19327);
and U21784 (N_21784,N_19168,N_20707);
nor U21785 (N_21785,N_19867,N_18764);
and U21786 (N_21786,N_19557,N_18027);
nand U21787 (N_21787,N_18600,N_18747);
xnor U21788 (N_21788,N_20563,N_18187);
nand U21789 (N_21789,N_18599,N_19110);
nand U21790 (N_21790,N_19266,N_18429);
and U21791 (N_21791,N_19645,N_19318);
or U21792 (N_21792,N_20963,N_18412);
nand U21793 (N_21793,N_18890,N_18362);
nand U21794 (N_21794,N_18283,N_19093);
nor U21795 (N_21795,N_19143,N_19475);
xnor U21796 (N_21796,N_20376,N_18483);
xnor U21797 (N_21797,N_19342,N_18188);
xor U21798 (N_21798,N_20572,N_18811);
or U21799 (N_21799,N_18303,N_18014);
xnor U21800 (N_21800,N_20228,N_18176);
and U21801 (N_21801,N_20463,N_19650);
or U21802 (N_21802,N_20868,N_19144);
or U21803 (N_21803,N_19647,N_18077);
or U21804 (N_21804,N_20117,N_20405);
nor U21805 (N_21805,N_19691,N_19103);
nor U21806 (N_21806,N_19344,N_18817);
and U21807 (N_21807,N_20483,N_18233);
xnor U21808 (N_21808,N_19527,N_19850);
nand U21809 (N_21809,N_18854,N_20350);
xor U21810 (N_21810,N_19771,N_20614);
and U21811 (N_21811,N_18474,N_19536);
nand U21812 (N_21812,N_18389,N_20542);
nor U21813 (N_21813,N_20427,N_20239);
nor U21814 (N_21814,N_20756,N_18468);
nor U21815 (N_21815,N_19061,N_18699);
and U21816 (N_21816,N_20691,N_18372);
nand U21817 (N_21817,N_19793,N_19566);
nor U21818 (N_21818,N_20242,N_20128);
or U21819 (N_21819,N_20253,N_19735);
xor U21820 (N_21820,N_19457,N_20712);
nand U21821 (N_21821,N_20662,N_20495);
nor U21822 (N_21822,N_20470,N_19486);
nor U21823 (N_21823,N_20385,N_18792);
xor U21824 (N_21824,N_18078,N_18150);
and U21825 (N_21825,N_20061,N_18897);
xnor U21826 (N_21826,N_19756,N_20235);
and U21827 (N_21827,N_19532,N_18590);
nand U21828 (N_21828,N_20653,N_19505);
and U21829 (N_21829,N_19633,N_18291);
nand U21830 (N_21830,N_18219,N_18030);
xor U21831 (N_21831,N_18285,N_18035);
or U21832 (N_21832,N_19276,N_19828);
nor U21833 (N_21833,N_18578,N_20439);
nand U21834 (N_21834,N_19747,N_20650);
or U21835 (N_21835,N_19118,N_19669);
nor U21836 (N_21836,N_18547,N_19080);
or U21837 (N_21837,N_20964,N_19097);
nor U21838 (N_21838,N_19891,N_20553);
or U21839 (N_21839,N_19319,N_20706);
nand U21840 (N_21840,N_19549,N_18382);
nand U21841 (N_21841,N_20271,N_20441);
or U21842 (N_21842,N_19571,N_20138);
and U21843 (N_21843,N_19733,N_20155);
and U21844 (N_21844,N_20531,N_19220);
nor U21845 (N_21845,N_19227,N_20067);
and U21846 (N_21846,N_19705,N_20406);
nand U21847 (N_21847,N_18345,N_18828);
or U21848 (N_21848,N_20190,N_19865);
xor U21849 (N_21849,N_20717,N_18880);
xor U21850 (N_21850,N_19967,N_18716);
and U21851 (N_21851,N_18693,N_19657);
and U21852 (N_21852,N_20137,N_19461);
nor U21853 (N_21853,N_18805,N_18344);
xor U21854 (N_21854,N_18185,N_20171);
and U21855 (N_21855,N_20726,N_20968);
xnor U21856 (N_21856,N_19638,N_18366);
and U21857 (N_21857,N_18902,N_18106);
and U21858 (N_21858,N_20947,N_19325);
nor U21859 (N_21859,N_18346,N_20896);
xnor U21860 (N_21860,N_19150,N_18183);
xor U21861 (N_21861,N_18056,N_19131);
xnor U21862 (N_21862,N_19317,N_18189);
and U21863 (N_21863,N_19406,N_19515);
xnor U21864 (N_21864,N_18312,N_18867);
nand U21865 (N_21865,N_20545,N_18787);
xnor U21866 (N_21866,N_20996,N_18177);
xor U21867 (N_21867,N_18640,N_18564);
or U21868 (N_21868,N_18612,N_18024);
nand U21869 (N_21869,N_19935,N_20649);
nand U21870 (N_21870,N_18968,N_19648);
nand U21871 (N_21871,N_19275,N_20528);
nor U21872 (N_21872,N_19859,N_19126);
nor U21873 (N_21873,N_20618,N_20489);
nand U21874 (N_21874,N_20915,N_19022);
and U21875 (N_21875,N_19136,N_19895);
nand U21876 (N_21876,N_19642,N_19692);
and U21877 (N_21877,N_18711,N_20619);
xnor U21878 (N_21878,N_19598,N_20461);
and U21879 (N_21879,N_18507,N_20814);
nand U21880 (N_21880,N_20069,N_18057);
nand U21881 (N_21881,N_19302,N_20771);
xnor U21882 (N_21882,N_19250,N_20143);
xnor U21883 (N_21883,N_20985,N_18478);
and U21884 (N_21884,N_18834,N_20689);
nand U21885 (N_21885,N_18624,N_18934);
nor U21886 (N_21886,N_18434,N_20606);
and U21887 (N_21887,N_20462,N_19075);
nand U21888 (N_21888,N_19844,N_20866);
xnor U21889 (N_21889,N_20505,N_18571);
nor U21890 (N_21890,N_20573,N_18761);
nand U21891 (N_21891,N_18963,N_18369);
nand U21892 (N_21892,N_18895,N_19646);
nand U21893 (N_21893,N_19272,N_19394);
nor U21894 (N_21894,N_19377,N_19501);
and U21895 (N_21895,N_18541,N_20471);
xnor U21896 (N_21896,N_19742,N_19600);
and U21897 (N_21897,N_20904,N_18520);
and U21898 (N_21898,N_18381,N_18394);
xor U21899 (N_21899,N_20676,N_20806);
nand U21900 (N_21900,N_19311,N_18795);
nand U21901 (N_21901,N_19847,N_18067);
or U21902 (N_21902,N_18648,N_18752);
nor U21903 (N_21903,N_20236,N_19857);
or U21904 (N_21904,N_19445,N_20532);
or U21905 (N_21905,N_20084,N_19543);
xnor U21906 (N_21906,N_20919,N_18261);
and U21907 (N_21907,N_19387,N_20416);
xor U21908 (N_21908,N_19145,N_19814);
nor U21909 (N_21909,N_19165,N_20145);
and U21910 (N_21910,N_18659,N_20525);
xor U21911 (N_21911,N_20077,N_19507);
or U21912 (N_21912,N_18974,N_19385);
or U21913 (N_21913,N_20783,N_20419);
nand U21914 (N_21914,N_20051,N_18780);
and U21915 (N_21915,N_18685,N_19576);
and U21916 (N_21916,N_20633,N_18907);
or U21917 (N_21917,N_19873,N_18684);
nor U21918 (N_21918,N_18420,N_18995);
and U21919 (N_21919,N_20533,N_20702);
nand U21920 (N_21920,N_18903,N_18791);
and U21921 (N_21921,N_18416,N_19254);
nor U21922 (N_21922,N_20511,N_19966);
nand U21923 (N_21923,N_19547,N_20838);
and U21924 (N_21924,N_20719,N_18370);
nor U21925 (N_21925,N_20620,N_20437);
nand U21926 (N_21926,N_19408,N_18427);
and U21927 (N_21927,N_20746,N_19197);
nor U21928 (N_21928,N_19913,N_19790);
and U21929 (N_21929,N_19417,N_18936);
and U21930 (N_21930,N_18784,N_20648);
nor U21931 (N_21931,N_20334,N_20380);
and U21932 (N_21932,N_18905,N_18638);
and U21933 (N_21933,N_18155,N_18472);
nand U21934 (N_21934,N_19060,N_20251);
nor U21935 (N_21935,N_20311,N_19225);
or U21936 (N_21936,N_18643,N_18671);
nor U21937 (N_21937,N_19182,N_18881);
or U21938 (N_21938,N_20199,N_20031);
nor U21939 (N_21939,N_19117,N_20975);
or U21940 (N_21940,N_18084,N_20231);
or U21941 (N_21941,N_20788,N_20279);
nor U21942 (N_21942,N_18365,N_18814);
nor U21943 (N_21943,N_20937,N_20167);
nand U21944 (N_21944,N_19351,N_18031);
xnor U21945 (N_21945,N_18920,N_19238);
xnor U21946 (N_21946,N_19644,N_20050);
nand U21947 (N_21947,N_20275,N_19591);
xnor U21948 (N_21948,N_18943,N_20693);
and U21949 (N_21949,N_18987,N_20423);
nand U21950 (N_21950,N_19412,N_19371);
xor U21951 (N_21951,N_19181,N_18396);
nor U21952 (N_21952,N_20431,N_19509);
xnor U21953 (N_21953,N_18083,N_19932);
xnor U21954 (N_21954,N_20711,N_19825);
nor U21955 (N_21955,N_18807,N_20749);
and U21956 (N_21956,N_18579,N_18915);
or U21957 (N_21957,N_18464,N_20767);
xor U21958 (N_21958,N_19862,N_19899);
xnor U21959 (N_21959,N_20833,N_18161);
or U21960 (N_21960,N_20579,N_18462);
xor U21961 (N_21961,N_20244,N_18172);
and U21962 (N_21962,N_18378,N_18335);
and U21963 (N_21963,N_20450,N_18006);
xor U21964 (N_21964,N_20809,N_20830);
nand U21965 (N_21965,N_19741,N_18609);
nand U21966 (N_21966,N_20800,N_19940);
nor U21967 (N_21967,N_19658,N_19380);
nor U21968 (N_21968,N_20534,N_18374);
or U21969 (N_21969,N_20363,N_19106);
nand U21970 (N_21970,N_19577,N_20034);
or U21971 (N_21971,N_20910,N_18758);
nor U21972 (N_21972,N_18667,N_20292);
xor U21973 (N_21973,N_19834,N_20064);
or U21974 (N_21974,N_18793,N_20237);
xnor U21975 (N_21975,N_20823,N_20272);
nand U21976 (N_21976,N_19748,N_20090);
nand U21977 (N_21977,N_19481,N_20558);
nand U21978 (N_21978,N_20704,N_20846);
nor U21979 (N_21979,N_18411,N_18677);
or U21980 (N_21980,N_20953,N_19195);
nand U21981 (N_21981,N_19628,N_19596);
xnor U21982 (N_21982,N_19274,N_19187);
nand U21983 (N_21983,N_18993,N_20987);
xor U21984 (N_21984,N_18167,N_18361);
nor U21985 (N_21985,N_18234,N_18490);
nor U21986 (N_21986,N_18829,N_19368);
and U21987 (N_21987,N_20867,N_20736);
nand U21988 (N_21988,N_19843,N_19123);
xor U21989 (N_21989,N_20507,N_20912);
nand U21990 (N_21990,N_19670,N_20647);
nand U21991 (N_21991,N_19459,N_20398);
and U21992 (N_21992,N_18306,N_19006);
nor U21993 (N_21993,N_19386,N_19091);
xor U21994 (N_21994,N_20344,N_20944);
nor U21995 (N_21995,N_18453,N_20133);
nor U21996 (N_21996,N_19044,N_18402);
and U21997 (N_21997,N_20859,N_18836);
and U21998 (N_21998,N_19309,N_20151);
nand U21999 (N_21999,N_18972,N_19245);
and U22000 (N_22000,N_19310,N_19100);
or U22001 (N_22001,N_20328,N_18644);
nand U22002 (N_22002,N_20085,N_18821);
nor U22003 (N_22003,N_18028,N_19513);
or U22004 (N_22004,N_20973,N_20798);
and U22005 (N_22005,N_19783,N_18254);
nand U22006 (N_22006,N_20781,N_18729);
xnor U22007 (N_22007,N_19390,N_18439);
or U22008 (N_22008,N_19490,N_20989);
or U22009 (N_22009,N_20263,N_18694);
and U22010 (N_22010,N_20024,N_18848);
nor U22011 (N_22011,N_18089,N_19774);
or U22012 (N_22012,N_19529,N_18327);
nor U22013 (N_22013,N_20490,N_20728);
xnor U22014 (N_22014,N_20580,N_18280);
or U22015 (N_22015,N_19694,N_20358);
xor U22016 (N_22016,N_18068,N_19095);
nor U22017 (N_22017,N_20313,N_18874);
and U22018 (N_22018,N_19791,N_20258);
nor U22019 (N_22019,N_19076,N_18652);
nand U22020 (N_22020,N_18975,N_18844);
xor U22021 (N_22021,N_19261,N_19968);
xor U22022 (N_22022,N_18486,N_18098);
and U22023 (N_22023,N_19888,N_20715);
or U22024 (N_22024,N_18608,N_20387);
nand U22025 (N_22025,N_20057,N_19294);
or U22026 (N_22026,N_20969,N_20325);
nor U22027 (N_22027,N_18162,N_20755);
nor U22028 (N_22028,N_18941,N_20481);
xnor U22029 (N_22029,N_18629,N_18202);
or U22030 (N_22030,N_18440,N_19624);
or U22031 (N_22031,N_20414,N_18066);
nor U22032 (N_22032,N_19972,N_18165);
nor U22033 (N_22033,N_18019,N_18186);
and U22034 (N_22034,N_18506,N_19038);
and U22035 (N_22035,N_20979,N_20709);
nand U22036 (N_22036,N_20266,N_18505);
nand U22037 (N_22037,N_19045,N_18804);
or U22038 (N_22038,N_19456,N_19039);
xor U22039 (N_22039,N_18986,N_19320);
nor U22040 (N_22040,N_20790,N_19700);
xor U22041 (N_22041,N_20222,N_18628);
or U22042 (N_22042,N_19027,N_20856);
nor U22043 (N_22043,N_19482,N_20695);
nor U22044 (N_22044,N_20083,N_20394);
nor U22045 (N_22045,N_20703,N_20931);
nor U22046 (N_22046,N_18725,N_18324);
and U22047 (N_22047,N_20402,N_20967);
xor U22048 (N_22048,N_19401,N_19358);
and U22049 (N_22049,N_19637,N_20154);
xnor U22050 (N_22050,N_19875,N_19789);
nor U22051 (N_22051,N_19455,N_18326);
nand U22052 (N_22052,N_19213,N_19778);
or U22053 (N_22053,N_19777,N_20374);
or U22054 (N_22054,N_20434,N_18554);
and U22055 (N_22055,N_18653,N_18072);
nand U22056 (N_22056,N_18141,N_18442);
xor U22057 (N_22057,N_20738,N_19114);
nor U22058 (N_22058,N_18544,N_19251);
nor U22059 (N_22059,N_20879,N_18017);
xor U22060 (N_22060,N_18515,N_20164);
nand U22061 (N_22061,N_20144,N_20195);
nand U22062 (N_22062,N_19904,N_18175);
or U22063 (N_22063,N_18536,N_19262);
xor U22064 (N_22064,N_18550,N_18253);
nor U22065 (N_22065,N_19804,N_20293);
nand U22066 (N_22066,N_20196,N_20863);
or U22067 (N_22067,N_19243,N_18243);
nand U22068 (N_22068,N_19246,N_18225);
or U22069 (N_22069,N_18517,N_19845);
nand U22070 (N_22070,N_20869,N_18214);
or U22071 (N_22071,N_19764,N_19827);
xor U22072 (N_22072,N_20546,N_20839);
nand U22073 (N_22073,N_20811,N_19169);
or U22074 (N_22074,N_18632,N_20476);
nand U22075 (N_22075,N_19166,N_18849);
nand U22076 (N_22076,N_20289,N_18565);
nor U22077 (N_22077,N_18794,N_20886);
and U22078 (N_22078,N_18563,N_18602);
xor U22079 (N_22079,N_19550,N_19734);
nand U22080 (N_22080,N_19425,N_20179);
and U22081 (N_22081,N_19485,N_20074);
nor U22082 (N_22082,N_20636,N_20769);
and U22083 (N_22083,N_20183,N_19689);
and U22084 (N_22084,N_19582,N_20841);
or U22085 (N_22085,N_18656,N_18405);
and U22086 (N_22086,N_19503,N_18290);
and U22087 (N_22087,N_19997,N_20365);
and U22088 (N_22088,N_18088,N_20452);
nand U22089 (N_22089,N_18313,N_18417);
nor U22090 (N_22090,N_19905,N_19702);
nor U22091 (N_22091,N_19887,N_20177);
and U22092 (N_22092,N_19141,N_18798);
or U22093 (N_22093,N_19001,N_19070);
or U22094 (N_22094,N_19193,N_19025);
xor U22095 (N_22095,N_18800,N_18724);
and U22096 (N_22096,N_18558,N_20066);
nor U22097 (N_22097,N_19542,N_18930);
or U22098 (N_22098,N_20391,N_18289);
and U22099 (N_22099,N_18293,N_19056);
xor U22100 (N_22100,N_20880,N_18928);
nor U22101 (N_22101,N_18317,N_18586);
nand U22102 (N_22102,N_19522,N_19281);
or U22103 (N_22103,N_20367,N_19177);
or U22104 (N_22104,N_20938,N_20312);
nand U22105 (N_22105,N_19113,N_19253);
xnor U22106 (N_22106,N_19077,N_20562);
xnor U22107 (N_22107,N_18438,N_20276);
or U22108 (N_22108,N_20030,N_18513);
and U22109 (N_22109,N_19725,N_20857);
nor U22110 (N_22110,N_19234,N_19744);
nor U22111 (N_22111,N_19603,N_18908);
and U22112 (N_22112,N_19797,N_19331);
and U22113 (N_22113,N_18753,N_19781);
or U22114 (N_22114,N_19122,N_19502);
nand U22115 (N_22115,N_20517,N_19444);
nand U22116 (N_22116,N_20329,N_18134);
xnor U22117 (N_22117,N_19673,N_19175);
nand U22118 (N_22118,N_18080,N_18142);
or U22119 (N_22119,N_18338,N_20826);
and U22120 (N_22120,N_18914,N_18432);
and U22121 (N_22121,N_20048,N_19798);
or U22122 (N_22122,N_18838,N_19308);
or U22123 (N_22123,N_19819,N_19273);
or U22124 (N_22124,N_19162,N_20535);
xor U22125 (N_22125,N_19332,N_19370);
nor U22126 (N_22126,N_20496,N_18649);
or U22127 (N_22127,N_20479,N_18641);
xor U22128 (N_22128,N_20596,N_19297);
nor U22129 (N_22129,N_18090,N_20012);
nand U22130 (N_22130,N_20742,N_20667);
nor U22131 (N_22131,N_19971,N_20250);
xnor U22132 (N_22132,N_18965,N_18418);
or U22133 (N_22133,N_19335,N_19548);
nor U22134 (N_22134,N_19519,N_19858);
or U22135 (N_22135,N_20760,N_20308);
xor U22136 (N_22136,N_20829,N_20730);
nor U22137 (N_22137,N_20497,N_20486);
nand U22138 (N_22138,N_20808,N_20370);
nand U22139 (N_22139,N_19977,N_20498);
nand U22140 (N_22140,N_20103,N_20418);
nand U22141 (N_22141,N_20040,N_19367);
nand U22142 (N_22142,N_20577,N_18921);
nand U22143 (N_22143,N_19938,N_20106);
and U22144 (N_22144,N_20227,N_18408);
nand U22145 (N_22145,N_18259,N_19533);
and U22146 (N_22146,N_18818,N_20223);
nand U22147 (N_22147,N_20684,N_18097);
and U22148 (N_22148,N_18197,N_19399);
and U22149 (N_22149,N_20637,N_20413);
and U22150 (N_22150,N_20021,N_20921);
nor U22151 (N_22151,N_18636,N_19415);
xor U22152 (N_22152,N_20092,N_19002);
and U22153 (N_22153,N_19954,N_18407);
nand U22154 (N_22154,N_20590,N_18193);
xor U22155 (N_22155,N_18307,N_19615);
nand U22156 (N_22156,N_20162,N_19958);
or U22157 (N_22157,N_18160,N_18398);
nor U22158 (N_22158,N_18395,N_19955);
nand U22159 (N_22159,N_18967,N_20327);
nor U22160 (N_22160,N_19023,N_20254);
nand U22161 (N_22161,N_18893,N_18841);
and U22162 (N_22162,N_19337,N_19289);
nand U22163 (N_22163,N_18220,N_20567);
nor U22164 (N_22164,N_20277,N_18422);
xor U22165 (N_22165,N_18731,N_18029);
and U22166 (N_22166,N_18998,N_19098);
and U22167 (N_22167,N_19925,N_18863);
nor U22168 (N_22168,N_20990,N_20321);
and U22169 (N_22169,N_20063,N_18955);
and U22170 (N_22170,N_19167,N_19226);
nand U22171 (N_22171,N_18889,N_19599);
and U22172 (N_22172,N_19498,N_18036);
nand U22173 (N_22173,N_20860,N_19398);
xor U22174 (N_22174,N_19714,N_18759);
nor U22175 (N_22175,N_18062,N_20226);
xor U22176 (N_22176,N_19018,N_18181);
nor U22177 (N_22177,N_19769,N_18383);
xnor U22178 (N_22178,N_18861,N_18466);
nand U22179 (N_22179,N_20421,N_18122);
nand U22180 (N_22180,N_18956,N_19229);
xor U22181 (N_22181,N_18169,N_18351);
nand U22182 (N_22182,N_18349,N_18896);
and U22183 (N_22183,N_20758,N_19664);
nand U22184 (N_22184,N_20451,N_20219);
nand U22185 (N_22185,N_19472,N_20129);
and U22186 (N_22186,N_19604,N_18568);
xnor U22187 (N_22187,N_19738,N_20282);
nor U22188 (N_22188,N_20465,N_18158);
nor U22189 (N_22189,N_19011,N_18393);
xor U22190 (N_22190,N_20561,N_20651);
nand U22191 (N_22191,N_18959,N_19194);
or U22192 (N_22192,N_19978,N_19765);
nand U22193 (N_22193,N_20218,N_19009);
nand U22194 (N_22194,N_20652,N_20135);
and U22195 (N_22195,N_18927,N_18359);
and U22196 (N_22196,N_20966,N_19806);
nand U22197 (N_22197,N_19260,N_19222);
and U22198 (N_22198,N_18314,N_19581);
and U22199 (N_22199,N_20581,N_19288);
nand U22200 (N_22200,N_18099,N_20043);
xnor U22201 (N_22201,N_19015,N_18360);
nand U22202 (N_22202,N_20259,N_19359);
and U22203 (N_22203,N_19823,N_20054);
xnor U22204 (N_22204,N_19710,N_20300);
nor U22205 (N_22205,N_20895,N_19296);
nand U22206 (N_22206,N_18614,N_19614);
nor U22207 (N_22207,N_19210,N_20802);
nor U22208 (N_22208,N_20743,N_18933);
nand U22209 (N_22209,N_18557,N_18810);
or U22210 (N_22210,N_19606,N_18245);
xnor U22211 (N_22211,N_18152,N_20176);
xor U22212 (N_22212,N_20611,N_18436);
nor U22213 (N_22213,N_18891,N_18341);
nand U22214 (N_22214,N_18678,N_20153);
nor U22215 (N_22215,N_19280,N_20882);
xnor U22216 (N_22216,N_20824,N_20845);
or U22217 (N_22217,N_19116,N_19671);
nor U22218 (N_22218,N_18937,N_19920);
nand U22219 (N_22219,N_20997,N_20603);
xor U22220 (N_22220,N_19048,N_18537);
nand U22221 (N_22221,N_18368,N_18491);
or U22222 (N_22222,N_19031,N_19473);
nor U22223 (N_22223,N_19892,N_20843);
and U22224 (N_22224,N_19209,N_18050);
or U22225 (N_22225,N_19007,N_18788);
nor U22226 (N_22226,N_19101,N_19762);
and U22227 (N_22227,N_19554,N_20877);
nand U22228 (N_22228,N_18005,N_19704);
xor U22229 (N_22229,N_20205,N_19133);
and U22230 (N_22230,N_20878,N_20364);
nor U22231 (N_22231,N_19820,N_19433);
nor U22232 (N_22232,N_19155,N_19265);
or U22233 (N_22233,N_19927,N_18917);
nand U22234 (N_22234,N_19584,N_18385);
or U22235 (N_22235,N_18046,N_20265);
xor U22236 (N_22236,N_18444,N_20403);
or U22237 (N_22237,N_19620,N_20349);
xor U22238 (N_22238,N_18413,N_20732);
xnor U22239 (N_22239,N_19612,N_19592);
nand U22240 (N_22240,N_18242,N_19636);
nor U22241 (N_22241,N_19772,N_19170);
xor U22242 (N_22242,N_20655,N_20295);
or U22243 (N_22243,N_19374,N_19339);
nand U22244 (N_22244,N_18910,N_18103);
or U22245 (N_22245,N_18215,N_20157);
xnor U22246 (N_22246,N_20629,N_19236);
nor U22247 (N_22247,N_20044,N_19998);
xor U22248 (N_22248,N_18319,N_18007);
and U22249 (N_22249,N_18380,N_20386);
nand U22250 (N_22250,N_19553,N_18840);
or U22251 (N_22251,N_19149,N_18698);
and U22252 (N_22252,N_19656,N_20352);
xor U22253 (N_22253,N_19231,N_19164);
or U22254 (N_22254,N_20589,N_18945);
xor U22255 (N_22255,N_19999,N_18645);
nand U22256 (N_22256,N_18717,N_18201);
nand U22257 (N_22257,N_19931,N_18768);
or U22258 (N_22258,N_20298,N_20635);
xnor U22259 (N_22259,N_20765,N_18477);
or U22260 (N_22260,N_19352,N_20032);
xor U22261 (N_22261,N_18756,N_20330);
nor U22262 (N_22262,N_18101,N_18459);
xor U22263 (N_22263,N_18710,N_20139);
nand U22264 (N_22264,N_18695,N_19083);
xor U22265 (N_22265,N_18114,N_20544);
nand U22266 (N_22266,N_18911,N_18783);
or U22267 (N_22267,N_20639,N_18583);
xor U22268 (N_22268,N_20933,N_19449);
or U22269 (N_22269,N_18588,N_18776);
and U22270 (N_22270,N_18322,N_19555);
or U22271 (N_22271,N_20172,N_18350);
nand U22272 (N_22272,N_18542,N_20551);
xnor U22273 (N_22273,N_18740,N_18045);
nor U22274 (N_22274,N_20246,N_20828);
xor U22275 (N_22275,N_18133,N_20460);
and U22276 (N_22276,N_19626,N_20453);
nand U22277 (N_22277,N_19523,N_18682);
xnor U22278 (N_22278,N_19393,N_20062);
nand U22279 (N_22279,N_20831,N_19081);
xnor U22280 (N_22280,N_19934,N_20274);
xor U22281 (N_22281,N_18942,N_18044);
nor U22282 (N_22282,N_19125,N_18096);
or U22283 (N_22283,N_19699,N_19414);
or U22284 (N_22284,N_18493,N_18958);
and U22285 (N_22285,N_19046,N_18178);
xor U22286 (N_22286,N_18329,N_18771);
and U22287 (N_22287,N_19047,N_18790);
nor U22288 (N_22288,N_18637,N_18079);
and U22289 (N_22289,N_18387,N_18948);
or U22290 (N_22290,N_20825,N_20810);
or U22291 (N_22291,N_18521,N_19438);
nand U22292 (N_22292,N_20923,N_18938);
nand U22293 (N_22293,N_19894,N_19178);
nor U22294 (N_22294,N_20946,N_18862);
nand U22295 (N_22295,N_19990,N_18715);
xor U22296 (N_22296,N_20110,N_19567);
or U22297 (N_22297,N_19928,N_19987);
and U22298 (N_22298,N_18680,N_20638);
or U22299 (N_22299,N_18081,N_20388);
or U22300 (N_22300,N_20230,N_18728);
nor U22301 (N_22301,N_18129,N_18404);
and U22302 (N_22302,N_20102,N_19158);
nor U22303 (N_22303,N_20526,N_19588);
nand U22304 (N_22304,N_20216,N_20932);
or U22305 (N_22305,N_20555,N_19573);
and U22306 (N_22306,N_19682,N_20052);
xor U22307 (N_22307,N_19304,N_19879);
nand U22308 (N_22308,N_18676,N_20182);
or U22309 (N_22309,N_19921,N_18763);
nand U22310 (N_22310,N_19183,N_18354);
nor U22311 (N_22311,N_20815,N_18143);
nor U22312 (N_22312,N_18048,N_19157);
nor U22313 (N_22313,N_18809,N_19366);
xnor U22314 (N_22314,N_18762,N_20918);
and U22315 (N_22315,N_20393,N_18613);
nor U22316 (N_22316,N_20093,N_19171);
xor U22317 (N_22317,N_20288,N_19930);
nor U22318 (N_22318,N_19079,N_18774);
xor U22319 (N_22319,N_20578,N_20727);
and U22320 (N_22320,N_20336,N_20733);
and U22321 (N_22321,N_19479,N_20522);
and U22322 (N_22322,N_18071,N_20821);
and U22323 (N_22323,N_19196,N_18485);
xnor U22324 (N_22324,N_18593,N_18153);
xor U22325 (N_22325,N_19973,N_18524);
xnor U22326 (N_22326,N_19146,N_19383);
nand U22327 (N_22327,N_19856,N_19369);
xnor U22328 (N_22328,N_20916,N_20571);
nor U22329 (N_22329,N_18492,N_20529);
xor U22330 (N_22330,N_19594,N_18767);
nor U22331 (N_22331,N_19298,N_18755);
xor U22332 (N_22332,N_20630,N_19893);
or U22333 (N_22333,N_19491,N_20037);
or U22334 (N_22334,N_18415,N_20267);
nand U22335 (N_22335,N_19792,N_19736);
xor U22336 (N_22336,N_19617,N_20004);
nand U22337 (N_22337,N_19970,N_20592);
and U22338 (N_22338,N_18925,N_20688);
or U22339 (N_22339,N_19562,N_19803);
nand U22340 (N_22340,N_20165,N_19729);
nand U22341 (N_22341,N_19976,N_18267);
nand U22342 (N_22342,N_19889,N_20124);
or U22343 (N_22343,N_20273,N_20956);
and U22344 (N_22344,N_18467,N_19676);
xor U22345 (N_22345,N_20503,N_19119);
and U22346 (N_22346,N_18497,N_20575);
and U22347 (N_22347,N_20046,N_20091);
or U22348 (N_22348,N_18247,N_18040);
xnor U22349 (N_22349,N_18371,N_20220);
xor U22350 (N_22350,N_19427,N_20696);
or U22351 (N_22351,N_20998,N_18281);
and U22352 (N_22352,N_18498,N_19919);
nor U22353 (N_22353,N_18340,N_20909);
nor U22354 (N_22354,N_20207,N_19223);
nand U22355 (N_22355,N_20081,N_19121);
and U22356 (N_22356,N_18566,N_20787);
or U22357 (N_22357,N_18576,N_20400);
nor U22358 (N_22358,N_19124,N_19109);
xor U22359 (N_22359,N_19217,N_20731);
or U22360 (N_22360,N_18428,N_19323);
and U22361 (N_22361,N_20792,N_19379);
or U22362 (N_22362,N_20892,N_18441);
nor U22363 (N_22363,N_20766,N_20991);
nor U22364 (N_22364,N_18857,N_19478);
and U22365 (N_22365,N_20192,N_18977);
xor U22366 (N_22366,N_20383,N_18047);
and U22367 (N_22367,N_20160,N_18037);
or U22368 (N_22368,N_20586,N_20735);
and U22369 (N_22369,N_18251,N_20152);
xnor U22370 (N_22370,N_19794,N_19026);
xor U22371 (N_22371,N_19355,N_19404);
and U22372 (N_22372,N_19483,N_20425);
nand U22373 (N_22373,N_19784,N_18610);
nand U22374 (N_22374,N_19590,N_20284);
or U22375 (N_22375,N_19835,N_19630);
nor U22376 (N_22376,N_20225,N_20939);
nor U22377 (N_22377,N_19153,N_18301);
nor U22378 (N_22378,N_20002,N_20015);
nor U22379 (N_22379,N_18796,N_20229);
xor U22380 (N_22380,N_19739,N_20747);
nor U22381 (N_22381,N_19306,N_18151);
xor U22382 (N_22382,N_19528,N_18631);
and U22383 (N_22383,N_18205,N_20822);
or U22384 (N_22384,N_20842,N_20248);
xor U22385 (N_22385,N_20390,N_20820);
xor U22386 (N_22386,N_20166,N_20286);
nor U22387 (N_22387,N_20320,N_20377);
or U22388 (N_22388,N_18086,N_19420);
xor U22389 (N_22389,N_20379,N_18320);
and U22390 (N_22390,N_19316,N_19411);
nand U22391 (N_22391,N_18476,N_19601);
nor U22392 (N_22392,N_19703,N_20785);
nand U22393 (N_22393,N_18962,N_19941);
xor U22394 (N_22394,N_19787,N_20661);
or U22395 (N_22395,N_20245,N_19952);
nor U22396 (N_22396,N_18074,N_19795);
xor U22397 (N_22397,N_20992,N_20426);
nor U22398 (N_22398,N_20672,N_20156);
nor U22399 (N_22399,N_18164,N_20888);
nor U22400 (N_22400,N_18373,N_18107);
xor U22401 (N_22401,N_19468,N_18877);
nor U22402 (N_22402,N_19268,N_18625);
xnor U22403 (N_22403,N_19349,N_18170);
nor U22404 (N_22404,N_20136,N_18075);
and U22405 (N_22405,N_18330,N_18743);
or U22406 (N_22406,N_19159,N_20616);
and U22407 (N_22407,N_19684,N_19267);
nand U22408 (N_22408,N_20269,N_19908);
xor U22409 (N_22409,N_20751,N_20404);
or U22410 (N_22410,N_18431,N_20520);
nor U22411 (N_22411,N_20631,N_20634);
xor U22412 (N_22412,N_18025,N_19334);
xnor U22413 (N_22413,N_20362,N_18666);
xnor U22414 (N_22414,N_20740,N_18686);
or U22415 (N_22415,N_19541,N_20955);
nor U22416 (N_22416,N_19467,N_20341);
or U22417 (N_22417,N_20764,N_19724);
and U22418 (N_22418,N_20326,N_19720);
and U22419 (N_22419,N_18512,N_18223);
nand U22420 (N_22420,N_19839,N_19984);
nor U22421 (N_22421,N_18532,N_18966);
or U22422 (N_22422,N_18556,N_19446);
and U22423 (N_22423,N_20565,N_20951);
or U22424 (N_22424,N_18271,N_18100);
xnor U22425 (N_22425,N_19421,N_19886);
and U22426 (N_22426,N_18487,N_19510);
nor U22427 (N_22427,N_18021,N_20494);
nand U22428 (N_22428,N_19811,N_18585);
and U22429 (N_22429,N_18489,N_18913);
nand U22430 (N_22430,N_19745,N_19431);
xor U22431 (N_22431,N_20212,N_20353);
xnor U22432 (N_22432,N_18782,N_18473);
and U22433 (N_22433,N_19679,N_18746);
xnor U22434 (N_22434,N_18668,N_20583);
xor U22435 (N_22435,N_18772,N_18410);
and U22436 (N_22436,N_19996,N_18148);
nand U22437 (N_22437,N_18858,N_18110);
or U22438 (N_22438,N_19654,N_18421);
and U22439 (N_22439,N_19228,N_20677);
nor U22440 (N_22440,N_20779,N_18376);
nand U22441 (N_22441,N_18392,N_19333);
xnor U22442 (N_22442,N_20795,N_18227);
nand U22443 (N_22443,N_18139,N_20378);
nor U22444 (N_22444,N_18607,N_18531);
nor U22445 (N_22445,N_20443,N_19202);
xnor U22446 (N_22446,N_19219,N_19869);
nand U22447 (N_22447,N_20690,N_20623);
nor U22448 (N_22448,N_19597,N_19128);
xnor U22449 (N_22449,N_18988,N_20007);
xor U22450 (N_22450,N_20925,N_19667);
xnor U22451 (N_22451,N_20210,N_20741);
xnor U22452 (N_22452,N_19872,N_20187);
and U22453 (N_22453,N_20080,N_20999);
or U22454 (N_22454,N_19621,N_18001);
nand U22455 (N_22455,N_20613,N_18870);
and U22456 (N_22456,N_20659,N_19613);
nor U22457 (N_22457,N_20710,N_19466);
nand U22458 (N_22458,N_20748,N_19775);
or U22459 (N_22459,N_18009,N_20252);
or U22460 (N_22460,N_19154,N_18263);
nor U22461 (N_22461,N_20924,N_18900);
nand U22462 (N_22462,N_18104,N_19322);
nor U22463 (N_22463,N_20444,N_20125);
nor U22464 (N_22464,N_19432,N_18179);
and U22465 (N_22465,N_19407,N_19391);
or U22466 (N_22466,N_18146,N_18789);
or U22467 (N_22467,N_20417,N_19078);
nor U22468 (N_22468,N_19683,N_19295);
or U22469 (N_22469,N_19137,N_18985);
and U22470 (N_22470,N_20281,N_20936);
xnor U22471 (N_22471,N_19595,N_19559);
and U22472 (N_22472,N_20357,N_20232);
nand U22473 (N_22473,N_18091,N_20126);
xor U22474 (N_22474,N_20014,N_20515);
nor U22475 (N_22475,N_18300,N_19841);
nor U22476 (N_22476,N_19403,N_20348);
nand U22477 (N_22477,N_18379,N_18594);
or U22478 (N_22478,N_18292,N_20900);
and U22479 (N_22479,N_18015,N_20601);
and U22480 (N_22480,N_19675,N_18449);
or U22481 (N_22481,N_18111,N_19556);
nor U22482 (N_22482,N_18250,N_19148);
or U22483 (N_22483,N_18138,N_19017);
nor U22484 (N_22484,N_19495,N_19487);
xnor U22485 (N_22485,N_20331,N_19680);
and U22486 (N_22486,N_19946,N_18085);
or U22487 (N_22487,N_19659,N_19037);
or U22488 (N_22488,N_19176,N_19982);
and U22489 (N_22489,N_19517,N_18509);
and U22490 (N_22490,N_18257,N_18265);
and U22491 (N_22491,N_18621,N_20920);
xnor U22492 (N_22492,N_19639,N_20003);
xor U22493 (N_22493,N_20013,N_18528);
or U22494 (N_22494,N_20911,N_18718);
xor U22495 (N_22495,N_20058,N_20477);
and U22496 (N_22496,N_20454,N_20198);
and U22497 (N_22497,N_20036,N_20435);
and U22498 (N_22498,N_20194,N_20891);
or U22499 (N_22499,N_19089,N_20105);
and U22500 (N_22500,N_19161,N_19062);
or U22501 (N_22501,N_20804,N_18107);
or U22502 (N_22502,N_18624,N_20356);
xnor U22503 (N_22503,N_18520,N_20260);
and U22504 (N_22504,N_19308,N_18421);
nand U22505 (N_22505,N_20827,N_19611);
and U22506 (N_22506,N_20709,N_18871);
and U22507 (N_22507,N_20196,N_20784);
nor U22508 (N_22508,N_19511,N_18473);
nor U22509 (N_22509,N_19611,N_18489);
nand U22510 (N_22510,N_18865,N_20801);
and U22511 (N_22511,N_19317,N_18491);
and U22512 (N_22512,N_19551,N_19508);
or U22513 (N_22513,N_18834,N_18143);
or U22514 (N_22514,N_18361,N_19467);
xnor U22515 (N_22515,N_19207,N_19271);
xor U22516 (N_22516,N_19780,N_18019);
xnor U22517 (N_22517,N_20504,N_18766);
nand U22518 (N_22518,N_19006,N_18743);
xnor U22519 (N_22519,N_19349,N_20619);
xor U22520 (N_22520,N_20729,N_19776);
or U22521 (N_22521,N_20981,N_19814);
nand U22522 (N_22522,N_20730,N_20466);
nor U22523 (N_22523,N_20395,N_18185);
xor U22524 (N_22524,N_20145,N_20284);
xor U22525 (N_22525,N_20820,N_19198);
nand U22526 (N_22526,N_20057,N_19443);
or U22527 (N_22527,N_19708,N_19447);
or U22528 (N_22528,N_20191,N_18299);
nor U22529 (N_22529,N_19871,N_18192);
nand U22530 (N_22530,N_20179,N_20718);
or U22531 (N_22531,N_19171,N_19958);
nor U22532 (N_22532,N_20947,N_20292);
nand U22533 (N_22533,N_20732,N_18654);
xor U22534 (N_22534,N_19843,N_19190);
and U22535 (N_22535,N_20505,N_18193);
xnor U22536 (N_22536,N_20593,N_19689);
nor U22537 (N_22537,N_19976,N_18270);
nor U22538 (N_22538,N_20844,N_20457);
nor U22539 (N_22539,N_19690,N_20157);
nor U22540 (N_22540,N_19069,N_20658);
xnor U22541 (N_22541,N_18428,N_19440);
or U22542 (N_22542,N_20408,N_18390);
xnor U22543 (N_22543,N_19866,N_19561);
or U22544 (N_22544,N_19177,N_19500);
xor U22545 (N_22545,N_18184,N_19762);
nor U22546 (N_22546,N_18113,N_19843);
or U22547 (N_22547,N_18596,N_19686);
or U22548 (N_22548,N_18301,N_18872);
or U22549 (N_22549,N_19395,N_19651);
or U22550 (N_22550,N_19289,N_20217);
nand U22551 (N_22551,N_19993,N_19492);
or U22552 (N_22552,N_18410,N_20345);
and U22553 (N_22553,N_19232,N_18622);
nand U22554 (N_22554,N_19520,N_19645);
nand U22555 (N_22555,N_18798,N_19193);
or U22556 (N_22556,N_20268,N_18988);
xnor U22557 (N_22557,N_20336,N_19222);
and U22558 (N_22558,N_18040,N_20957);
nor U22559 (N_22559,N_18771,N_19785);
nor U22560 (N_22560,N_19462,N_20828);
nor U22561 (N_22561,N_19838,N_18527);
xnor U22562 (N_22562,N_19681,N_18873);
nand U22563 (N_22563,N_19257,N_19354);
or U22564 (N_22564,N_20291,N_18858);
xor U22565 (N_22565,N_20130,N_20789);
xnor U22566 (N_22566,N_20357,N_18148);
or U22567 (N_22567,N_18252,N_20523);
and U22568 (N_22568,N_19110,N_18524);
and U22569 (N_22569,N_20200,N_18467);
and U22570 (N_22570,N_18105,N_19733);
nor U22571 (N_22571,N_19961,N_18481);
and U22572 (N_22572,N_19066,N_20172);
nand U22573 (N_22573,N_18586,N_19104);
and U22574 (N_22574,N_18257,N_18385);
nor U22575 (N_22575,N_19062,N_18374);
xor U22576 (N_22576,N_18646,N_20669);
and U22577 (N_22577,N_20735,N_18273);
xor U22578 (N_22578,N_18906,N_19802);
xnor U22579 (N_22579,N_18548,N_18685);
nor U22580 (N_22580,N_19604,N_18149);
nor U22581 (N_22581,N_18629,N_18381);
or U22582 (N_22582,N_18361,N_19915);
nand U22583 (N_22583,N_20569,N_19402);
nor U22584 (N_22584,N_18545,N_20654);
or U22585 (N_22585,N_18779,N_19738);
xor U22586 (N_22586,N_19658,N_20790);
xor U22587 (N_22587,N_18947,N_20289);
xnor U22588 (N_22588,N_20274,N_19465);
nand U22589 (N_22589,N_20374,N_18268);
or U22590 (N_22590,N_20491,N_20459);
or U22591 (N_22591,N_20808,N_18280);
and U22592 (N_22592,N_18502,N_19003);
or U22593 (N_22593,N_20928,N_19968);
nand U22594 (N_22594,N_19249,N_18270);
xnor U22595 (N_22595,N_20817,N_18266);
nand U22596 (N_22596,N_20744,N_19107);
and U22597 (N_22597,N_18473,N_18947);
xnor U22598 (N_22598,N_19565,N_18526);
or U22599 (N_22599,N_18998,N_18267);
xnor U22600 (N_22600,N_20244,N_19526);
and U22601 (N_22601,N_18646,N_20624);
nand U22602 (N_22602,N_20955,N_20394);
and U22603 (N_22603,N_18146,N_19990);
nor U22604 (N_22604,N_18864,N_20733);
nand U22605 (N_22605,N_18488,N_19751);
and U22606 (N_22606,N_19694,N_18236);
xor U22607 (N_22607,N_18172,N_20401);
or U22608 (N_22608,N_20197,N_20667);
nand U22609 (N_22609,N_20447,N_19336);
xnor U22610 (N_22610,N_20955,N_20485);
or U22611 (N_22611,N_20353,N_18661);
xor U22612 (N_22612,N_20199,N_18756);
nand U22613 (N_22613,N_20731,N_19793);
xor U22614 (N_22614,N_18150,N_20741);
or U22615 (N_22615,N_19977,N_19549);
or U22616 (N_22616,N_19236,N_18749);
xor U22617 (N_22617,N_18448,N_20022);
and U22618 (N_22618,N_19939,N_20311);
nor U22619 (N_22619,N_19158,N_20819);
and U22620 (N_22620,N_18177,N_18373);
and U22621 (N_22621,N_20262,N_18037);
or U22622 (N_22622,N_20786,N_19803);
and U22623 (N_22623,N_19634,N_18618);
nand U22624 (N_22624,N_19382,N_18031);
nor U22625 (N_22625,N_19966,N_20734);
xnor U22626 (N_22626,N_18342,N_20704);
nor U22627 (N_22627,N_18246,N_19688);
nor U22628 (N_22628,N_20002,N_19090);
xor U22629 (N_22629,N_20422,N_19406);
nand U22630 (N_22630,N_18444,N_20184);
nand U22631 (N_22631,N_18970,N_20174);
xor U22632 (N_22632,N_19757,N_18000);
xor U22633 (N_22633,N_20397,N_18758);
and U22634 (N_22634,N_20212,N_18607);
and U22635 (N_22635,N_18048,N_18474);
xnor U22636 (N_22636,N_19086,N_19034);
nor U22637 (N_22637,N_20686,N_19952);
nand U22638 (N_22638,N_20461,N_19530);
or U22639 (N_22639,N_19336,N_19723);
nand U22640 (N_22640,N_18804,N_19219);
xor U22641 (N_22641,N_19456,N_19908);
nand U22642 (N_22642,N_19508,N_20962);
xnor U22643 (N_22643,N_18593,N_20770);
or U22644 (N_22644,N_20409,N_20010);
or U22645 (N_22645,N_19297,N_18306);
xnor U22646 (N_22646,N_20828,N_20108);
nand U22647 (N_22647,N_18044,N_19766);
xnor U22648 (N_22648,N_20176,N_19978);
and U22649 (N_22649,N_18738,N_18946);
nand U22650 (N_22650,N_19323,N_19766);
nor U22651 (N_22651,N_19345,N_20149);
xnor U22652 (N_22652,N_20763,N_18431);
xor U22653 (N_22653,N_19151,N_18231);
xor U22654 (N_22654,N_20503,N_18409);
nand U22655 (N_22655,N_18955,N_20232);
xor U22656 (N_22656,N_19256,N_20517);
and U22657 (N_22657,N_18119,N_18736);
nor U22658 (N_22658,N_19311,N_19331);
nand U22659 (N_22659,N_20172,N_18721);
nand U22660 (N_22660,N_20562,N_18420);
nand U22661 (N_22661,N_18751,N_19650);
xnor U22662 (N_22662,N_20982,N_20074);
and U22663 (N_22663,N_18460,N_20150);
and U22664 (N_22664,N_20397,N_18710);
and U22665 (N_22665,N_20118,N_18322);
and U22666 (N_22666,N_20231,N_18049);
xnor U22667 (N_22667,N_20690,N_20544);
nor U22668 (N_22668,N_18711,N_19270);
xor U22669 (N_22669,N_19631,N_20282);
nand U22670 (N_22670,N_20148,N_19561);
nor U22671 (N_22671,N_20399,N_18641);
nand U22672 (N_22672,N_20581,N_18540);
nand U22673 (N_22673,N_19008,N_18209);
and U22674 (N_22674,N_19016,N_18982);
and U22675 (N_22675,N_20079,N_18518);
nor U22676 (N_22676,N_18659,N_19784);
xor U22677 (N_22677,N_20606,N_20532);
and U22678 (N_22678,N_19813,N_18619);
and U22679 (N_22679,N_18470,N_18590);
nand U22680 (N_22680,N_19401,N_18023);
nand U22681 (N_22681,N_20608,N_19645);
xnor U22682 (N_22682,N_19011,N_18957);
nor U22683 (N_22683,N_18913,N_20964);
nor U22684 (N_22684,N_20989,N_20830);
nand U22685 (N_22685,N_19507,N_18812);
nor U22686 (N_22686,N_20921,N_18117);
nor U22687 (N_22687,N_18479,N_19922);
nor U22688 (N_22688,N_19323,N_20205);
xnor U22689 (N_22689,N_20897,N_18488);
or U22690 (N_22690,N_20884,N_18028);
or U22691 (N_22691,N_20759,N_20262);
nand U22692 (N_22692,N_19421,N_19255);
xor U22693 (N_22693,N_19269,N_20924);
nand U22694 (N_22694,N_18389,N_19533);
nand U22695 (N_22695,N_18403,N_20126);
nor U22696 (N_22696,N_19841,N_18418);
nand U22697 (N_22697,N_20244,N_18505);
or U22698 (N_22698,N_19893,N_20506);
nor U22699 (N_22699,N_20328,N_18632);
and U22700 (N_22700,N_19116,N_20612);
or U22701 (N_22701,N_19447,N_18943);
xnor U22702 (N_22702,N_18762,N_19438);
xor U22703 (N_22703,N_18156,N_19522);
xnor U22704 (N_22704,N_19777,N_20629);
or U22705 (N_22705,N_19795,N_20671);
nor U22706 (N_22706,N_19284,N_19430);
xnor U22707 (N_22707,N_20998,N_19483);
xnor U22708 (N_22708,N_18191,N_20861);
and U22709 (N_22709,N_20339,N_19323);
or U22710 (N_22710,N_19243,N_19444);
nor U22711 (N_22711,N_20857,N_19786);
xnor U22712 (N_22712,N_18106,N_20925);
and U22713 (N_22713,N_18512,N_18876);
nand U22714 (N_22714,N_19343,N_20693);
nor U22715 (N_22715,N_18400,N_19169);
xnor U22716 (N_22716,N_18003,N_19478);
or U22717 (N_22717,N_20624,N_19313);
xnor U22718 (N_22718,N_20025,N_20606);
or U22719 (N_22719,N_20201,N_20129);
and U22720 (N_22720,N_19945,N_19116);
nand U22721 (N_22721,N_18170,N_18933);
nand U22722 (N_22722,N_20761,N_18265);
or U22723 (N_22723,N_20610,N_19867);
or U22724 (N_22724,N_19107,N_19311);
nor U22725 (N_22725,N_20716,N_18615);
xor U22726 (N_22726,N_19475,N_19919);
nor U22727 (N_22727,N_20444,N_19089);
or U22728 (N_22728,N_18153,N_19634);
nor U22729 (N_22729,N_18731,N_18619);
xnor U22730 (N_22730,N_19829,N_19585);
nand U22731 (N_22731,N_20325,N_20039);
and U22732 (N_22732,N_19044,N_18467);
and U22733 (N_22733,N_18559,N_18696);
nor U22734 (N_22734,N_18490,N_18635);
nor U22735 (N_22735,N_19395,N_18461);
nor U22736 (N_22736,N_19694,N_20071);
nor U22737 (N_22737,N_20932,N_20919);
nor U22738 (N_22738,N_19423,N_18133);
and U22739 (N_22739,N_20237,N_18140);
nor U22740 (N_22740,N_18909,N_20197);
xor U22741 (N_22741,N_18907,N_19527);
nand U22742 (N_22742,N_18490,N_18660);
xor U22743 (N_22743,N_18749,N_19411);
and U22744 (N_22744,N_19095,N_18749);
xnor U22745 (N_22745,N_19821,N_20589);
nand U22746 (N_22746,N_19704,N_20081);
or U22747 (N_22747,N_19454,N_18863);
xor U22748 (N_22748,N_19560,N_18861);
nor U22749 (N_22749,N_20870,N_18592);
xnor U22750 (N_22750,N_20670,N_18125);
xor U22751 (N_22751,N_20240,N_19299);
or U22752 (N_22752,N_20050,N_20369);
and U22753 (N_22753,N_19329,N_20728);
xnor U22754 (N_22754,N_18253,N_19186);
or U22755 (N_22755,N_20472,N_18098);
nor U22756 (N_22756,N_19811,N_20143);
or U22757 (N_22757,N_20059,N_18180);
xor U22758 (N_22758,N_20364,N_18937);
nor U22759 (N_22759,N_18354,N_18187);
nand U22760 (N_22760,N_18139,N_19552);
xor U22761 (N_22761,N_18761,N_19653);
nand U22762 (N_22762,N_20644,N_18070);
xor U22763 (N_22763,N_19412,N_18857);
nand U22764 (N_22764,N_20112,N_18892);
or U22765 (N_22765,N_18101,N_19726);
nor U22766 (N_22766,N_20000,N_19922);
and U22767 (N_22767,N_19061,N_19300);
nor U22768 (N_22768,N_20515,N_20617);
xor U22769 (N_22769,N_20530,N_18646);
nor U22770 (N_22770,N_19710,N_20598);
xor U22771 (N_22771,N_20664,N_18544);
nand U22772 (N_22772,N_20105,N_18504);
and U22773 (N_22773,N_19388,N_20198);
nor U22774 (N_22774,N_19798,N_18048);
nor U22775 (N_22775,N_18972,N_20025);
and U22776 (N_22776,N_20762,N_20801);
nand U22777 (N_22777,N_19122,N_19465);
nor U22778 (N_22778,N_20498,N_19907);
or U22779 (N_22779,N_19737,N_19938);
or U22780 (N_22780,N_18185,N_20856);
nand U22781 (N_22781,N_20100,N_19340);
and U22782 (N_22782,N_18981,N_20940);
xor U22783 (N_22783,N_20980,N_20511);
xor U22784 (N_22784,N_18096,N_19631);
and U22785 (N_22785,N_19257,N_20130);
xnor U22786 (N_22786,N_18150,N_20554);
and U22787 (N_22787,N_19043,N_18562);
xor U22788 (N_22788,N_18202,N_19499);
nor U22789 (N_22789,N_20199,N_19257);
and U22790 (N_22790,N_20261,N_20025);
nand U22791 (N_22791,N_20108,N_19300);
or U22792 (N_22792,N_20059,N_20565);
or U22793 (N_22793,N_20242,N_20245);
or U22794 (N_22794,N_18052,N_20279);
nor U22795 (N_22795,N_18892,N_20215);
nand U22796 (N_22796,N_20868,N_20913);
xnor U22797 (N_22797,N_19911,N_18630);
and U22798 (N_22798,N_18161,N_20898);
or U22799 (N_22799,N_18174,N_19179);
and U22800 (N_22800,N_18984,N_19925);
or U22801 (N_22801,N_19853,N_19462);
and U22802 (N_22802,N_19516,N_19919);
nor U22803 (N_22803,N_18060,N_19447);
nand U22804 (N_22804,N_19238,N_18729);
and U22805 (N_22805,N_18381,N_19402);
nor U22806 (N_22806,N_18365,N_18008);
and U22807 (N_22807,N_20502,N_20802);
and U22808 (N_22808,N_18363,N_20438);
or U22809 (N_22809,N_18219,N_19566);
and U22810 (N_22810,N_20642,N_19085);
and U22811 (N_22811,N_18628,N_19273);
nand U22812 (N_22812,N_18703,N_19180);
nor U22813 (N_22813,N_19174,N_20292);
and U22814 (N_22814,N_18475,N_20368);
nand U22815 (N_22815,N_20289,N_18021);
nand U22816 (N_22816,N_20130,N_20024);
nand U22817 (N_22817,N_20914,N_20620);
nor U22818 (N_22818,N_20828,N_18773);
nand U22819 (N_22819,N_18354,N_20732);
and U22820 (N_22820,N_18368,N_18598);
and U22821 (N_22821,N_18818,N_18297);
xnor U22822 (N_22822,N_20460,N_19980);
nand U22823 (N_22823,N_20968,N_20436);
and U22824 (N_22824,N_18499,N_19655);
and U22825 (N_22825,N_20987,N_19653);
and U22826 (N_22826,N_18275,N_20280);
or U22827 (N_22827,N_20155,N_20704);
xor U22828 (N_22828,N_20457,N_20856);
and U22829 (N_22829,N_19075,N_18689);
xnor U22830 (N_22830,N_18583,N_18076);
and U22831 (N_22831,N_19595,N_18588);
nor U22832 (N_22832,N_20195,N_20944);
nor U22833 (N_22833,N_18659,N_20470);
nor U22834 (N_22834,N_20157,N_19506);
nor U22835 (N_22835,N_19060,N_19924);
and U22836 (N_22836,N_19370,N_20178);
xor U22837 (N_22837,N_20678,N_19620);
nor U22838 (N_22838,N_19072,N_18446);
nand U22839 (N_22839,N_20216,N_19174);
nand U22840 (N_22840,N_19086,N_20962);
or U22841 (N_22841,N_18827,N_18313);
or U22842 (N_22842,N_18522,N_18165);
nor U22843 (N_22843,N_19819,N_18192);
and U22844 (N_22844,N_18331,N_20519);
or U22845 (N_22845,N_19631,N_19301);
and U22846 (N_22846,N_20175,N_19276);
and U22847 (N_22847,N_20390,N_19110);
xor U22848 (N_22848,N_20880,N_19108);
and U22849 (N_22849,N_20654,N_18909);
and U22850 (N_22850,N_20202,N_19641);
or U22851 (N_22851,N_19558,N_19904);
and U22852 (N_22852,N_19310,N_18163);
xor U22853 (N_22853,N_18488,N_18904);
nor U22854 (N_22854,N_20910,N_20069);
or U22855 (N_22855,N_18507,N_20205);
or U22856 (N_22856,N_18241,N_18789);
nor U22857 (N_22857,N_19043,N_19970);
and U22858 (N_22858,N_20631,N_20617);
xnor U22859 (N_22859,N_19331,N_19732);
xor U22860 (N_22860,N_20892,N_18016);
xnor U22861 (N_22861,N_20473,N_18091);
and U22862 (N_22862,N_19998,N_18668);
and U22863 (N_22863,N_19759,N_18380);
xor U22864 (N_22864,N_20916,N_18977);
and U22865 (N_22865,N_20260,N_18043);
nor U22866 (N_22866,N_19744,N_20024);
and U22867 (N_22867,N_20145,N_19416);
xor U22868 (N_22868,N_18283,N_19153);
nand U22869 (N_22869,N_20755,N_19758);
or U22870 (N_22870,N_18479,N_20182);
and U22871 (N_22871,N_18670,N_19703);
xnor U22872 (N_22872,N_19739,N_20848);
nor U22873 (N_22873,N_20328,N_20779);
xnor U22874 (N_22874,N_18868,N_19423);
nand U22875 (N_22875,N_20307,N_20586);
xnor U22876 (N_22876,N_20539,N_19414);
and U22877 (N_22877,N_20434,N_20763);
nand U22878 (N_22878,N_19918,N_20005);
and U22879 (N_22879,N_20467,N_18021);
nand U22880 (N_22880,N_19188,N_18991);
nand U22881 (N_22881,N_18951,N_19312);
and U22882 (N_22882,N_20157,N_18980);
xnor U22883 (N_22883,N_18156,N_18757);
or U22884 (N_22884,N_19785,N_19076);
xor U22885 (N_22885,N_18309,N_18636);
and U22886 (N_22886,N_18957,N_20925);
or U22887 (N_22887,N_18021,N_19276);
and U22888 (N_22888,N_19872,N_19256);
nand U22889 (N_22889,N_20039,N_19628);
xor U22890 (N_22890,N_19444,N_18810);
or U22891 (N_22891,N_18777,N_18395);
xor U22892 (N_22892,N_18790,N_18844);
and U22893 (N_22893,N_19285,N_20561);
nor U22894 (N_22894,N_18709,N_19799);
and U22895 (N_22895,N_18584,N_18006);
nor U22896 (N_22896,N_20722,N_20189);
and U22897 (N_22897,N_20419,N_18267);
and U22898 (N_22898,N_20938,N_20698);
nor U22899 (N_22899,N_18336,N_19663);
and U22900 (N_22900,N_18497,N_19015);
xnor U22901 (N_22901,N_18252,N_19428);
xnor U22902 (N_22902,N_18543,N_20930);
nand U22903 (N_22903,N_20273,N_18736);
or U22904 (N_22904,N_19926,N_20357);
nor U22905 (N_22905,N_19789,N_19880);
nand U22906 (N_22906,N_20268,N_18886);
xnor U22907 (N_22907,N_20434,N_20045);
nand U22908 (N_22908,N_19334,N_19920);
nand U22909 (N_22909,N_18599,N_18771);
xnor U22910 (N_22910,N_18982,N_18540);
or U22911 (N_22911,N_19496,N_20165);
and U22912 (N_22912,N_19062,N_19451);
nand U22913 (N_22913,N_20372,N_20422);
xnor U22914 (N_22914,N_18582,N_20259);
and U22915 (N_22915,N_18237,N_20895);
xor U22916 (N_22916,N_20134,N_18511);
and U22917 (N_22917,N_20655,N_20810);
and U22918 (N_22918,N_18361,N_19809);
xnor U22919 (N_22919,N_19449,N_18198);
and U22920 (N_22920,N_19613,N_19796);
nor U22921 (N_22921,N_19380,N_19076);
nand U22922 (N_22922,N_20898,N_19599);
nor U22923 (N_22923,N_19342,N_19985);
and U22924 (N_22924,N_18064,N_18599);
nand U22925 (N_22925,N_20587,N_18079);
and U22926 (N_22926,N_19882,N_20218);
or U22927 (N_22927,N_18649,N_20126);
nor U22928 (N_22928,N_20758,N_18285);
or U22929 (N_22929,N_20881,N_20174);
nor U22930 (N_22930,N_20338,N_20940);
nand U22931 (N_22931,N_20767,N_20879);
nor U22932 (N_22932,N_20279,N_19246);
xnor U22933 (N_22933,N_18702,N_18923);
or U22934 (N_22934,N_18018,N_19007);
nand U22935 (N_22935,N_18696,N_19205);
xor U22936 (N_22936,N_18284,N_19570);
or U22937 (N_22937,N_18023,N_20388);
xor U22938 (N_22938,N_19637,N_19181);
or U22939 (N_22939,N_19402,N_20410);
nor U22940 (N_22940,N_20036,N_19776);
nand U22941 (N_22941,N_18347,N_20474);
nor U22942 (N_22942,N_18551,N_18448);
nand U22943 (N_22943,N_20790,N_19716);
nor U22944 (N_22944,N_19536,N_20544);
nand U22945 (N_22945,N_18997,N_18396);
and U22946 (N_22946,N_20922,N_19260);
nor U22947 (N_22947,N_19720,N_19721);
and U22948 (N_22948,N_19059,N_20396);
nor U22949 (N_22949,N_18229,N_19107);
nand U22950 (N_22950,N_19169,N_20402);
xor U22951 (N_22951,N_18281,N_18009);
and U22952 (N_22952,N_20699,N_20551);
nor U22953 (N_22953,N_20110,N_20298);
nor U22954 (N_22954,N_20372,N_19989);
nand U22955 (N_22955,N_18031,N_20463);
nand U22956 (N_22956,N_20203,N_19219);
and U22957 (N_22957,N_20221,N_18689);
nor U22958 (N_22958,N_19226,N_18035);
and U22959 (N_22959,N_19850,N_19953);
xor U22960 (N_22960,N_18471,N_18347);
or U22961 (N_22961,N_19994,N_20699);
and U22962 (N_22962,N_20527,N_19192);
xor U22963 (N_22963,N_19847,N_20364);
and U22964 (N_22964,N_20816,N_19397);
and U22965 (N_22965,N_19740,N_20193);
nand U22966 (N_22966,N_18709,N_20622);
and U22967 (N_22967,N_20342,N_20222);
nor U22968 (N_22968,N_19286,N_19035);
and U22969 (N_22969,N_20146,N_18159);
nor U22970 (N_22970,N_18058,N_19038);
nor U22971 (N_22971,N_19291,N_18932);
or U22972 (N_22972,N_18440,N_19235);
nor U22973 (N_22973,N_19248,N_20649);
xor U22974 (N_22974,N_20147,N_20278);
xnor U22975 (N_22975,N_20212,N_18413);
nand U22976 (N_22976,N_18116,N_18842);
nand U22977 (N_22977,N_20529,N_19180);
nand U22978 (N_22978,N_19563,N_18813);
xor U22979 (N_22979,N_19381,N_19058);
nor U22980 (N_22980,N_18599,N_19881);
nor U22981 (N_22981,N_20769,N_19549);
nor U22982 (N_22982,N_19676,N_18845);
and U22983 (N_22983,N_18129,N_18373);
nand U22984 (N_22984,N_19352,N_18688);
and U22985 (N_22985,N_18560,N_19496);
and U22986 (N_22986,N_19732,N_18996);
and U22987 (N_22987,N_20776,N_20948);
nand U22988 (N_22988,N_19346,N_20254);
nand U22989 (N_22989,N_20134,N_18351);
nor U22990 (N_22990,N_18459,N_19997);
or U22991 (N_22991,N_19724,N_18559);
nor U22992 (N_22992,N_20902,N_20497);
nand U22993 (N_22993,N_18166,N_19828);
nand U22994 (N_22994,N_20687,N_18688);
nand U22995 (N_22995,N_18190,N_20218);
and U22996 (N_22996,N_18025,N_19495);
nor U22997 (N_22997,N_18580,N_20381);
or U22998 (N_22998,N_20961,N_20518);
nand U22999 (N_22999,N_18107,N_19106);
or U23000 (N_23000,N_19537,N_18077);
nand U23001 (N_23001,N_18112,N_20617);
xor U23002 (N_23002,N_18306,N_20963);
or U23003 (N_23003,N_20971,N_18624);
and U23004 (N_23004,N_18732,N_20994);
or U23005 (N_23005,N_18051,N_20105);
xnor U23006 (N_23006,N_20169,N_19151);
or U23007 (N_23007,N_19929,N_19849);
and U23008 (N_23008,N_19182,N_18939);
and U23009 (N_23009,N_20683,N_18021);
xor U23010 (N_23010,N_18306,N_20396);
xor U23011 (N_23011,N_19452,N_19745);
nand U23012 (N_23012,N_19019,N_19845);
nand U23013 (N_23013,N_19736,N_18116);
nand U23014 (N_23014,N_20344,N_18131);
and U23015 (N_23015,N_18492,N_20325);
and U23016 (N_23016,N_20481,N_20282);
nor U23017 (N_23017,N_18434,N_20127);
xnor U23018 (N_23018,N_18951,N_18214);
xor U23019 (N_23019,N_20462,N_18532);
or U23020 (N_23020,N_19251,N_18289);
xnor U23021 (N_23021,N_18700,N_18116);
or U23022 (N_23022,N_18760,N_20510);
xnor U23023 (N_23023,N_18076,N_20161);
or U23024 (N_23024,N_18061,N_19420);
and U23025 (N_23025,N_18464,N_19009);
nand U23026 (N_23026,N_19072,N_20008);
xnor U23027 (N_23027,N_19399,N_20105);
and U23028 (N_23028,N_20337,N_18946);
or U23029 (N_23029,N_18554,N_20594);
xor U23030 (N_23030,N_19318,N_19498);
xnor U23031 (N_23031,N_18008,N_18589);
nor U23032 (N_23032,N_18609,N_19510);
nor U23033 (N_23033,N_20976,N_19931);
or U23034 (N_23034,N_19827,N_19927);
or U23035 (N_23035,N_19035,N_18191);
or U23036 (N_23036,N_19076,N_20747);
or U23037 (N_23037,N_18485,N_19532);
xnor U23038 (N_23038,N_19611,N_18000);
xor U23039 (N_23039,N_18698,N_20071);
or U23040 (N_23040,N_19947,N_19429);
nand U23041 (N_23041,N_19405,N_18308);
xnor U23042 (N_23042,N_19613,N_19820);
and U23043 (N_23043,N_20130,N_20145);
or U23044 (N_23044,N_19272,N_19980);
or U23045 (N_23045,N_20925,N_20850);
or U23046 (N_23046,N_20180,N_19398);
nor U23047 (N_23047,N_20247,N_19992);
or U23048 (N_23048,N_18899,N_19882);
or U23049 (N_23049,N_18788,N_20682);
nor U23050 (N_23050,N_20353,N_19789);
and U23051 (N_23051,N_18817,N_19841);
and U23052 (N_23052,N_20898,N_19984);
nor U23053 (N_23053,N_19381,N_18574);
and U23054 (N_23054,N_20559,N_20607);
nand U23055 (N_23055,N_19042,N_18569);
or U23056 (N_23056,N_18892,N_19852);
xnor U23057 (N_23057,N_19474,N_20122);
nor U23058 (N_23058,N_18237,N_18968);
xor U23059 (N_23059,N_19637,N_18192);
and U23060 (N_23060,N_18423,N_20000);
nor U23061 (N_23061,N_19614,N_19138);
and U23062 (N_23062,N_18814,N_20880);
xor U23063 (N_23063,N_20835,N_19856);
nor U23064 (N_23064,N_20282,N_18004);
and U23065 (N_23065,N_18301,N_18361);
nor U23066 (N_23066,N_20711,N_20553);
xor U23067 (N_23067,N_19001,N_19807);
xnor U23068 (N_23068,N_18317,N_20300);
nor U23069 (N_23069,N_20005,N_19428);
nand U23070 (N_23070,N_18409,N_18628);
or U23071 (N_23071,N_20805,N_19147);
nor U23072 (N_23072,N_19015,N_20206);
nor U23073 (N_23073,N_19151,N_19882);
nor U23074 (N_23074,N_19462,N_18337);
xnor U23075 (N_23075,N_20842,N_19881);
xor U23076 (N_23076,N_18775,N_20228);
and U23077 (N_23077,N_18901,N_19360);
nor U23078 (N_23078,N_20568,N_18222);
nor U23079 (N_23079,N_18353,N_20785);
nand U23080 (N_23080,N_18287,N_18719);
and U23081 (N_23081,N_20974,N_19850);
xor U23082 (N_23082,N_18922,N_20330);
xnor U23083 (N_23083,N_20905,N_18900);
xnor U23084 (N_23084,N_20209,N_20063);
nor U23085 (N_23085,N_18207,N_18235);
or U23086 (N_23086,N_18778,N_20885);
xor U23087 (N_23087,N_20590,N_18709);
nand U23088 (N_23088,N_18125,N_18801);
nor U23089 (N_23089,N_19429,N_18334);
and U23090 (N_23090,N_18902,N_19673);
and U23091 (N_23091,N_19073,N_18823);
nand U23092 (N_23092,N_20961,N_19463);
nand U23093 (N_23093,N_19399,N_18770);
nand U23094 (N_23094,N_20607,N_20818);
nand U23095 (N_23095,N_19241,N_18523);
and U23096 (N_23096,N_18419,N_19919);
and U23097 (N_23097,N_20414,N_20268);
or U23098 (N_23098,N_20593,N_19633);
and U23099 (N_23099,N_20173,N_20705);
xor U23100 (N_23100,N_19361,N_18226);
nor U23101 (N_23101,N_18282,N_19387);
xor U23102 (N_23102,N_19924,N_19730);
nor U23103 (N_23103,N_20563,N_18622);
or U23104 (N_23104,N_19208,N_18004);
and U23105 (N_23105,N_18465,N_20444);
or U23106 (N_23106,N_19747,N_19538);
nand U23107 (N_23107,N_18861,N_19127);
nand U23108 (N_23108,N_18184,N_18012);
nor U23109 (N_23109,N_18011,N_19354);
nor U23110 (N_23110,N_20358,N_19841);
xnor U23111 (N_23111,N_20572,N_19097);
xnor U23112 (N_23112,N_20522,N_18088);
or U23113 (N_23113,N_19289,N_20584);
xnor U23114 (N_23114,N_20463,N_20288);
nand U23115 (N_23115,N_20416,N_19622);
nor U23116 (N_23116,N_19410,N_19011);
xnor U23117 (N_23117,N_18389,N_18901);
and U23118 (N_23118,N_19483,N_18242);
or U23119 (N_23119,N_19109,N_20825);
or U23120 (N_23120,N_18331,N_19352);
nand U23121 (N_23121,N_19186,N_19482);
and U23122 (N_23122,N_18418,N_18159);
xnor U23123 (N_23123,N_19274,N_18021);
xnor U23124 (N_23124,N_18468,N_18159);
nor U23125 (N_23125,N_18611,N_19068);
nor U23126 (N_23126,N_20372,N_20423);
xor U23127 (N_23127,N_20779,N_18491);
or U23128 (N_23128,N_18572,N_18381);
and U23129 (N_23129,N_19805,N_18844);
nand U23130 (N_23130,N_19849,N_20730);
or U23131 (N_23131,N_18617,N_20309);
nand U23132 (N_23132,N_18327,N_18795);
and U23133 (N_23133,N_20500,N_18572);
nor U23134 (N_23134,N_19412,N_19873);
and U23135 (N_23135,N_20062,N_19137);
nor U23136 (N_23136,N_20077,N_20052);
xor U23137 (N_23137,N_20579,N_18441);
xnor U23138 (N_23138,N_20578,N_20924);
and U23139 (N_23139,N_19311,N_19751);
nand U23140 (N_23140,N_18555,N_20662);
and U23141 (N_23141,N_18223,N_19216);
and U23142 (N_23142,N_19596,N_18378);
nor U23143 (N_23143,N_20323,N_19574);
xor U23144 (N_23144,N_19666,N_18292);
or U23145 (N_23145,N_20975,N_19080);
or U23146 (N_23146,N_20735,N_18862);
nor U23147 (N_23147,N_18737,N_19979);
xnor U23148 (N_23148,N_18665,N_19714);
and U23149 (N_23149,N_18808,N_19662);
nand U23150 (N_23150,N_18593,N_18976);
and U23151 (N_23151,N_18940,N_18542);
nor U23152 (N_23152,N_20387,N_19193);
and U23153 (N_23153,N_19095,N_20555);
xnor U23154 (N_23154,N_19866,N_18503);
nand U23155 (N_23155,N_19021,N_18973);
and U23156 (N_23156,N_18498,N_20322);
and U23157 (N_23157,N_18058,N_18281);
and U23158 (N_23158,N_19113,N_18790);
xnor U23159 (N_23159,N_19771,N_19770);
or U23160 (N_23160,N_20859,N_20083);
xor U23161 (N_23161,N_20353,N_18203);
nand U23162 (N_23162,N_19025,N_18160);
nor U23163 (N_23163,N_19059,N_19545);
nand U23164 (N_23164,N_18354,N_20908);
xnor U23165 (N_23165,N_19420,N_18893);
nor U23166 (N_23166,N_19922,N_19585);
nor U23167 (N_23167,N_20804,N_20718);
nand U23168 (N_23168,N_19856,N_19691);
and U23169 (N_23169,N_19088,N_19044);
nand U23170 (N_23170,N_20265,N_20424);
nor U23171 (N_23171,N_19735,N_19699);
xor U23172 (N_23172,N_20298,N_20368);
xor U23173 (N_23173,N_20854,N_18528);
nor U23174 (N_23174,N_18889,N_20672);
or U23175 (N_23175,N_19809,N_20066);
or U23176 (N_23176,N_20363,N_18345);
nand U23177 (N_23177,N_20903,N_19409);
nand U23178 (N_23178,N_18143,N_19645);
xor U23179 (N_23179,N_20432,N_19889);
or U23180 (N_23180,N_20087,N_18287);
nand U23181 (N_23181,N_20368,N_19913);
nand U23182 (N_23182,N_19073,N_19976);
xnor U23183 (N_23183,N_19221,N_19484);
or U23184 (N_23184,N_19333,N_20273);
nor U23185 (N_23185,N_18783,N_20404);
nor U23186 (N_23186,N_18157,N_19495);
nor U23187 (N_23187,N_18985,N_19807);
and U23188 (N_23188,N_19222,N_20362);
nand U23189 (N_23189,N_19742,N_19709);
nand U23190 (N_23190,N_19227,N_18108);
xor U23191 (N_23191,N_20128,N_19718);
xnor U23192 (N_23192,N_20782,N_19091);
and U23193 (N_23193,N_20455,N_20078);
nor U23194 (N_23194,N_18816,N_19444);
nand U23195 (N_23195,N_18253,N_19809);
xnor U23196 (N_23196,N_18396,N_19658);
or U23197 (N_23197,N_19671,N_20228);
or U23198 (N_23198,N_18928,N_20400);
and U23199 (N_23199,N_20500,N_19077);
nor U23200 (N_23200,N_18927,N_18199);
and U23201 (N_23201,N_19793,N_20774);
nand U23202 (N_23202,N_19344,N_20209);
nor U23203 (N_23203,N_19345,N_20080);
and U23204 (N_23204,N_19270,N_20739);
nand U23205 (N_23205,N_20859,N_18912);
xnor U23206 (N_23206,N_19367,N_19945);
nand U23207 (N_23207,N_20184,N_20707);
and U23208 (N_23208,N_19174,N_18279);
and U23209 (N_23209,N_19033,N_18216);
xnor U23210 (N_23210,N_19721,N_18982);
nand U23211 (N_23211,N_19420,N_20341);
xnor U23212 (N_23212,N_18971,N_18784);
xor U23213 (N_23213,N_20833,N_18270);
nor U23214 (N_23214,N_18350,N_20207);
nand U23215 (N_23215,N_19914,N_18246);
nand U23216 (N_23216,N_19521,N_19594);
nand U23217 (N_23217,N_18443,N_20831);
or U23218 (N_23218,N_20138,N_20091);
or U23219 (N_23219,N_18384,N_19035);
or U23220 (N_23220,N_20284,N_20206);
and U23221 (N_23221,N_19757,N_20818);
nand U23222 (N_23222,N_18697,N_20273);
and U23223 (N_23223,N_20271,N_18006);
nand U23224 (N_23224,N_19643,N_18307);
nor U23225 (N_23225,N_19653,N_19736);
nand U23226 (N_23226,N_19593,N_20594);
xnor U23227 (N_23227,N_19982,N_20340);
or U23228 (N_23228,N_18452,N_18925);
xnor U23229 (N_23229,N_20183,N_20519);
nand U23230 (N_23230,N_19962,N_19356);
nor U23231 (N_23231,N_20261,N_19754);
xnor U23232 (N_23232,N_19793,N_18846);
nor U23233 (N_23233,N_20702,N_19287);
nor U23234 (N_23234,N_19852,N_18382);
xor U23235 (N_23235,N_19587,N_18029);
or U23236 (N_23236,N_20281,N_19590);
nand U23237 (N_23237,N_20217,N_20717);
or U23238 (N_23238,N_20563,N_20644);
and U23239 (N_23239,N_19857,N_20226);
and U23240 (N_23240,N_18908,N_20731);
or U23241 (N_23241,N_18698,N_18427);
and U23242 (N_23242,N_19000,N_19187);
nand U23243 (N_23243,N_19842,N_20824);
nand U23244 (N_23244,N_19893,N_20336);
xnor U23245 (N_23245,N_20438,N_18959);
and U23246 (N_23246,N_19429,N_19377);
and U23247 (N_23247,N_19772,N_20025);
xnor U23248 (N_23248,N_20163,N_19523);
nand U23249 (N_23249,N_18576,N_19541);
nand U23250 (N_23250,N_19142,N_19593);
nor U23251 (N_23251,N_20667,N_19526);
nand U23252 (N_23252,N_19048,N_18411);
nand U23253 (N_23253,N_20158,N_20873);
and U23254 (N_23254,N_20782,N_19157);
xor U23255 (N_23255,N_19408,N_19314);
nor U23256 (N_23256,N_20206,N_19635);
xor U23257 (N_23257,N_19505,N_18291);
xnor U23258 (N_23258,N_18807,N_18477);
or U23259 (N_23259,N_19339,N_20369);
nand U23260 (N_23260,N_20855,N_20946);
or U23261 (N_23261,N_19982,N_18409);
nor U23262 (N_23262,N_19524,N_18037);
nand U23263 (N_23263,N_18568,N_18063);
nor U23264 (N_23264,N_20870,N_19740);
and U23265 (N_23265,N_20254,N_18901);
nand U23266 (N_23266,N_19733,N_19576);
xor U23267 (N_23267,N_18359,N_20416);
nand U23268 (N_23268,N_20736,N_19742);
or U23269 (N_23269,N_18518,N_19799);
nor U23270 (N_23270,N_20141,N_19900);
and U23271 (N_23271,N_18649,N_18548);
and U23272 (N_23272,N_20880,N_18725);
nand U23273 (N_23273,N_18155,N_19648);
nand U23274 (N_23274,N_19601,N_18712);
xor U23275 (N_23275,N_19998,N_18829);
xnor U23276 (N_23276,N_18292,N_18177);
nand U23277 (N_23277,N_18617,N_18812);
or U23278 (N_23278,N_20750,N_18098);
xnor U23279 (N_23279,N_20688,N_18414);
and U23280 (N_23280,N_20645,N_18445);
and U23281 (N_23281,N_20238,N_18230);
and U23282 (N_23282,N_20040,N_18201);
and U23283 (N_23283,N_20278,N_18542);
or U23284 (N_23284,N_18593,N_18094);
or U23285 (N_23285,N_20161,N_19847);
xnor U23286 (N_23286,N_19034,N_18095);
xnor U23287 (N_23287,N_20045,N_18015);
xor U23288 (N_23288,N_20055,N_19122);
xnor U23289 (N_23289,N_20640,N_18252);
nand U23290 (N_23290,N_20596,N_20267);
xor U23291 (N_23291,N_19163,N_20893);
nand U23292 (N_23292,N_20173,N_19107);
xnor U23293 (N_23293,N_18561,N_20068);
or U23294 (N_23294,N_20169,N_20698);
xnor U23295 (N_23295,N_18660,N_18330);
xnor U23296 (N_23296,N_20632,N_19049);
nand U23297 (N_23297,N_18196,N_18052);
nor U23298 (N_23298,N_20738,N_18659);
and U23299 (N_23299,N_20537,N_20182);
and U23300 (N_23300,N_18285,N_18207);
nand U23301 (N_23301,N_19315,N_19780);
nor U23302 (N_23302,N_20680,N_18421);
and U23303 (N_23303,N_18525,N_19520);
or U23304 (N_23304,N_20420,N_19877);
and U23305 (N_23305,N_20815,N_20985);
nor U23306 (N_23306,N_19543,N_20006);
or U23307 (N_23307,N_19967,N_18316);
and U23308 (N_23308,N_20401,N_20372);
nor U23309 (N_23309,N_18738,N_20897);
xor U23310 (N_23310,N_20455,N_19805);
nor U23311 (N_23311,N_20113,N_20731);
xor U23312 (N_23312,N_18529,N_20390);
nor U23313 (N_23313,N_19367,N_20028);
and U23314 (N_23314,N_20693,N_18252);
nor U23315 (N_23315,N_19142,N_20324);
and U23316 (N_23316,N_20700,N_19532);
or U23317 (N_23317,N_19420,N_20561);
nand U23318 (N_23318,N_18861,N_18453);
and U23319 (N_23319,N_18641,N_18807);
nor U23320 (N_23320,N_20110,N_20713);
and U23321 (N_23321,N_19479,N_19960);
or U23322 (N_23322,N_18780,N_18778);
xor U23323 (N_23323,N_20031,N_19277);
nor U23324 (N_23324,N_18334,N_19631);
and U23325 (N_23325,N_18866,N_18606);
or U23326 (N_23326,N_18580,N_18720);
or U23327 (N_23327,N_18881,N_18418);
nand U23328 (N_23328,N_18616,N_20483);
nand U23329 (N_23329,N_20653,N_18822);
and U23330 (N_23330,N_19312,N_18321);
or U23331 (N_23331,N_20857,N_18220);
or U23332 (N_23332,N_19422,N_19960);
nor U23333 (N_23333,N_18364,N_18104);
nor U23334 (N_23334,N_20604,N_18832);
or U23335 (N_23335,N_20684,N_19523);
nand U23336 (N_23336,N_19099,N_18479);
and U23337 (N_23337,N_19557,N_18104);
nand U23338 (N_23338,N_19624,N_18760);
or U23339 (N_23339,N_18322,N_19862);
nor U23340 (N_23340,N_19704,N_20028);
nand U23341 (N_23341,N_19412,N_20296);
nor U23342 (N_23342,N_18835,N_18955);
nor U23343 (N_23343,N_20810,N_20585);
or U23344 (N_23344,N_18385,N_20776);
xnor U23345 (N_23345,N_19146,N_20830);
nand U23346 (N_23346,N_19939,N_19091);
nand U23347 (N_23347,N_19304,N_19973);
xor U23348 (N_23348,N_18472,N_19956);
or U23349 (N_23349,N_20288,N_18379);
nand U23350 (N_23350,N_19484,N_19807);
or U23351 (N_23351,N_20328,N_19785);
nand U23352 (N_23352,N_20498,N_18405);
nor U23353 (N_23353,N_18468,N_18068);
and U23354 (N_23354,N_18705,N_19668);
xnor U23355 (N_23355,N_20735,N_20283);
nor U23356 (N_23356,N_18731,N_20489);
or U23357 (N_23357,N_18459,N_19180);
nor U23358 (N_23358,N_19938,N_18096);
xnor U23359 (N_23359,N_18761,N_18497);
nor U23360 (N_23360,N_20397,N_19419);
or U23361 (N_23361,N_18787,N_20750);
xor U23362 (N_23362,N_18836,N_19500);
nand U23363 (N_23363,N_20451,N_20361);
nor U23364 (N_23364,N_19682,N_18354);
and U23365 (N_23365,N_18611,N_19066);
nor U23366 (N_23366,N_20170,N_20428);
and U23367 (N_23367,N_19523,N_19167);
nor U23368 (N_23368,N_19041,N_19849);
or U23369 (N_23369,N_20599,N_19329);
and U23370 (N_23370,N_19971,N_18242);
nor U23371 (N_23371,N_20758,N_19722);
nor U23372 (N_23372,N_20318,N_19399);
nor U23373 (N_23373,N_18880,N_19804);
xnor U23374 (N_23374,N_20062,N_20519);
xnor U23375 (N_23375,N_20723,N_18684);
xnor U23376 (N_23376,N_19155,N_19884);
and U23377 (N_23377,N_20521,N_18939);
nor U23378 (N_23378,N_19586,N_18077);
nor U23379 (N_23379,N_18769,N_18370);
or U23380 (N_23380,N_20529,N_19515);
or U23381 (N_23381,N_18729,N_19824);
nand U23382 (N_23382,N_18482,N_18461);
or U23383 (N_23383,N_20476,N_20310);
xnor U23384 (N_23384,N_20604,N_20805);
nand U23385 (N_23385,N_18793,N_20224);
nor U23386 (N_23386,N_20592,N_20215);
or U23387 (N_23387,N_19738,N_20342);
xor U23388 (N_23388,N_19668,N_18133);
nand U23389 (N_23389,N_19293,N_18161);
nor U23390 (N_23390,N_19404,N_20763);
and U23391 (N_23391,N_20057,N_19574);
or U23392 (N_23392,N_19672,N_19455);
or U23393 (N_23393,N_20138,N_20045);
or U23394 (N_23394,N_18259,N_20830);
nand U23395 (N_23395,N_20322,N_20812);
xor U23396 (N_23396,N_20419,N_20641);
nor U23397 (N_23397,N_20155,N_18226);
nor U23398 (N_23398,N_18055,N_19160);
or U23399 (N_23399,N_19557,N_19766);
and U23400 (N_23400,N_18027,N_20521);
xor U23401 (N_23401,N_20852,N_19004);
xor U23402 (N_23402,N_19461,N_18088);
and U23403 (N_23403,N_19121,N_18397);
nand U23404 (N_23404,N_18230,N_19586);
or U23405 (N_23405,N_19369,N_20782);
xor U23406 (N_23406,N_20109,N_19272);
nor U23407 (N_23407,N_20333,N_19330);
xor U23408 (N_23408,N_20770,N_19582);
nand U23409 (N_23409,N_20472,N_20063);
and U23410 (N_23410,N_20605,N_19279);
nor U23411 (N_23411,N_19986,N_18061);
or U23412 (N_23412,N_19926,N_18414);
nand U23413 (N_23413,N_20095,N_19078);
nand U23414 (N_23414,N_20147,N_18269);
xor U23415 (N_23415,N_19692,N_18146);
nor U23416 (N_23416,N_19615,N_19522);
or U23417 (N_23417,N_20265,N_20292);
nand U23418 (N_23418,N_19887,N_18150);
nor U23419 (N_23419,N_19602,N_20457);
and U23420 (N_23420,N_20324,N_18144);
nor U23421 (N_23421,N_18959,N_19108);
nor U23422 (N_23422,N_19758,N_20714);
xnor U23423 (N_23423,N_19316,N_20993);
and U23424 (N_23424,N_18919,N_20446);
and U23425 (N_23425,N_18737,N_18312);
nand U23426 (N_23426,N_19687,N_19617);
xnor U23427 (N_23427,N_18683,N_18746);
xor U23428 (N_23428,N_18322,N_18869);
and U23429 (N_23429,N_20731,N_18552);
and U23430 (N_23430,N_18985,N_20877);
nor U23431 (N_23431,N_20154,N_19699);
nor U23432 (N_23432,N_20965,N_18798);
xnor U23433 (N_23433,N_19247,N_20730);
xor U23434 (N_23434,N_18962,N_19399);
xor U23435 (N_23435,N_20981,N_20674);
nor U23436 (N_23436,N_18196,N_20809);
xnor U23437 (N_23437,N_18560,N_20700);
nand U23438 (N_23438,N_18446,N_19861);
nor U23439 (N_23439,N_19176,N_19023);
and U23440 (N_23440,N_20262,N_18072);
nor U23441 (N_23441,N_20388,N_20965);
xor U23442 (N_23442,N_19034,N_20846);
xor U23443 (N_23443,N_19189,N_19679);
xor U23444 (N_23444,N_20302,N_20318);
nor U23445 (N_23445,N_18435,N_19522);
nand U23446 (N_23446,N_19151,N_19245);
nand U23447 (N_23447,N_20926,N_19134);
nand U23448 (N_23448,N_18225,N_20469);
nor U23449 (N_23449,N_19761,N_18027);
xor U23450 (N_23450,N_19760,N_18506);
nand U23451 (N_23451,N_20140,N_20531);
nand U23452 (N_23452,N_20467,N_19536);
nand U23453 (N_23453,N_18275,N_19486);
nor U23454 (N_23454,N_19720,N_20213);
nor U23455 (N_23455,N_18051,N_18776);
nor U23456 (N_23456,N_19162,N_20193);
nor U23457 (N_23457,N_20266,N_18400);
or U23458 (N_23458,N_20325,N_19743);
or U23459 (N_23459,N_19562,N_20085);
nor U23460 (N_23460,N_20098,N_20108);
or U23461 (N_23461,N_18028,N_18246);
and U23462 (N_23462,N_18018,N_18267);
nand U23463 (N_23463,N_18975,N_20997);
nand U23464 (N_23464,N_19746,N_18093);
or U23465 (N_23465,N_18364,N_20197);
or U23466 (N_23466,N_19830,N_19338);
nor U23467 (N_23467,N_19052,N_18495);
nand U23468 (N_23468,N_20245,N_20843);
nand U23469 (N_23469,N_18192,N_18291);
nor U23470 (N_23470,N_18942,N_20890);
and U23471 (N_23471,N_18544,N_18478);
or U23472 (N_23472,N_18860,N_18479);
nand U23473 (N_23473,N_18635,N_20060);
xor U23474 (N_23474,N_19240,N_18405);
nor U23475 (N_23475,N_18487,N_19134);
xor U23476 (N_23476,N_18570,N_20855);
nand U23477 (N_23477,N_18131,N_20433);
or U23478 (N_23478,N_18052,N_19611);
xnor U23479 (N_23479,N_20221,N_20396);
or U23480 (N_23480,N_20811,N_20362);
xnor U23481 (N_23481,N_20383,N_20365);
nand U23482 (N_23482,N_19421,N_20373);
and U23483 (N_23483,N_19116,N_20105);
and U23484 (N_23484,N_20620,N_18467);
nor U23485 (N_23485,N_19001,N_19900);
or U23486 (N_23486,N_18862,N_20278);
or U23487 (N_23487,N_18557,N_20580);
nand U23488 (N_23488,N_19413,N_18430);
nand U23489 (N_23489,N_20282,N_19951);
and U23490 (N_23490,N_20196,N_20459);
and U23491 (N_23491,N_20035,N_18664);
xnor U23492 (N_23492,N_18690,N_19649);
xnor U23493 (N_23493,N_18157,N_19533);
and U23494 (N_23494,N_19543,N_18178);
and U23495 (N_23495,N_19608,N_18913);
nand U23496 (N_23496,N_19740,N_18030);
or U23497 (N_23497,N_18980,N_20813);
nand U23498 (N_23498,N_19831,N_19156);
and U23499 (N_23499,N_18611,N_20600);
xor U23500 (N_23500,N_20791,N_18368);
xnor U23501 (N_23501,N_19497,N_20367);
xor U23502 (N_23502,N_20531,N_20743);
nand U23503 (N_23503,N_19342,N_19260);
nor U23504 (N_23504,N_18829,N_18016);
xnor U23505 (N_23505,N_19648,N_19541);
and U23506 (N_23506,N_20633,N_19029);
or U23507 (N_23507,N_20392,N_19367);
nor U23508 (N_23508,N_19951,N_20052);
nand U23509 (N_23509,N_19943,N_19679);
or U23510 (N_23510,N_19276,N_18334);
nand U23511 (N_23511,N_18973,N_20740);
nand U23512 (N_23512,N_18078,N_20183);
and U23513 (N_23513,N_18159,N_19826);
and U23514 (N_23514,N_18328,N_19810);
xnor U23515 (N_23515,N_20229,N_18614);
xor U23516 (N_23516,N_18539,N_18031);
xor U23517 (N_23517,N_20749,N_18352);
and U23518 (N_23518,N_18696,N_19507);
xnor U23519 (N_23519,N_18322,N_19857);
and U23520 (N_23520,N_20672,N_20978);
or U23521 (N_23521,N_20131,N_18732);
or U23522 (N_23522,N_20503,N_20955);
nand U23523 (N_23523,N_20882,N_18587);
nor U23524 (N_23524,N_20445,N_20543);
xnor U23525 (N_23525,N_20971,N_20535);
nor U23526 (N_23526,N_18154,N_20021);
and U23527 (N_23527,N_18998,N_18910);
and U23528 (N_23528,N_20593,N_18933);
nor U23529 (N_23529,N_19091,N_18968);
xor U23530 (N_23530,N_18735,N_18661);
nor U23531 (N_23531,N_19908,N_18362);
nand U23532 (N_23532,N_18697,N_18135);
and U23533 (N_23533,N_19376,N_19676);
xor U23534 (N_23534,N_19302,N_18371);
or U23535 (N_23535,N_19814,N_19382);
and U23536 (N_23536,N_19916,N_18364);
and U23537 (N_23537,N_20863,N_19130);
and U23538 (N_23538,N_18150,N_19594);
or U23539 (N_23539,N_20087,N_18414);
xnor U23540 (N_23540,N_18457,N_18652);
nor U23541 (N_23541,N_20863,N_18098);
xnor U23542 (N_23542,N_20123,N_19439);
or U23543 (N_23543,N_20423,N_19483);
or U23544 (N_23544,N_18566,N_19535);
nand U23545 (N_23545,N_19366,N_18739);
nor U23546 (N_23546,N_18873,N_19335);
nor U23547 (N_23547,N_18555,N_19411);
nand U23548 (N_23548,N_18115,N_18724);
or U23549 (N_23549,N_19531,N_19169);
nand U23550 (N_23550,N_20135,N_18686);
or U23551 (N_23551,N_20531,N_20396);
nand U23552 (N_23552,N_19793,N_20275);
and U23553 (N_23553,N_20673,N_20054);
xnor U23554 (N_23554,N_20975,N_20705);
nor U23555 (N_23555,N_20499,N_19749);
xor U23556 (N_23556,N_19624,N_20587);
and U23557 (N_23557,N_20245,N_19199);
or U23558 (N_23558,N_19868,N_20420);
and U23559 (N_23559,N_20395,N_19897);
and U23560 (N_23560,N_20845,N_19032);
nor U23561 (N_23561,N_20354,N_18470);
or U23562 (N_23562,N_18488,N_19304);
and U23563 (N_23563,N_19151,N_19776);
nand U23564 (N_23564,N_18465,N_20751);
nor U23565 (N_23565,N_20331,N_20172);
xnor U23566 (N_23566,N_20653,N_20662);
nor U23567 (N_23567,N_20320,N_18206);
or U23568 (N_23568,N_19105,N_19474);
and U23569 (N_23569,N_19365,N_20392);
nor U23570 (N_23570,N_20051,N_20329);
nand U23571 (N_23571,N_18219,N_18828);
nand U23572 (N_23572,N_19996,N_19333);
nor U23573 (N_23573,N_20789,N_18173);
nor U23574 (N_23574,N_18523,N_20386);
and U23575 (N_23575,N_20121,N_20136);
or U23576 (N_23576,N_20304,N_20986);
nand U23577 (N_23577,N_20636,N_20964);
or U23578 (N_23578,N_18843,N_20616);
nor U23579 (N_23579,N_20581,N_18340);
nor U23580 (N_23580,N_20856,N_20789);
xnor U23581 (N_23581,N_19373,N_18103);
and U23582 (N_23582,N_18212,N_18214);
and U23583 (N_23583,N_18863,N_20592);
nor U23584 (N_23584,N_19612,N_20405);
and U23585 (N_23585,N_19117,N_19505);
nor U23586 (N_23586,N_20677,N_19165);
xnor U23587 (N_23587,N_20220,N_19121);
nand U23588 (N_23588,N_20978,N_18212);
nor U23589 (N_23589,N_18585,N_20989);
and U23590 (N_23590,N_20643,N_20830);
xnor U23591 (N_23591,N_19964,N_20473);
and U23592 (N_23592,N_19576,N_19047);
nor U23593 (N_23593,N_19664,N_19111);
xor U23594 (N_23594,N_20121,N_18262);
xnor U23595 (N_23595,N_20832,N_18948);
nor U23596 (N_23596,N_18875,N_18716);
xor U23597 (N_23597,N_19853,N_18839);
nand U23598 (N_23598,N_19458,N_20798);
and U23599 (N_23599,N_19699,N_19468);
nor U23600 (N_23600,N_19172,N_18623);
or U23601 (N_23601,N_20741,N_18637);
and U23602 (N_23602,N_20574,N_19924);
and U23603 (N_23603,N_20420,N_18161);
nand U23604 (N_23604,N_18884,N_19725);
nand U23605 (N_23605,N_18906,N_20082);
nor U23606 (N_23606,N_19543,N_20286);
or U23607 (N_23607,N_18877,N_19567);
nor U23608 (N_23608,N_20860,N_19091);
nand U23609 (N_23609,N_19609,N_18299);
nor U23610 (N_23610,N_19899,N_19551);
xor U23611 (N_23611,N_19984,N_18945);
and U23612 (N_23612,N_18785,N_19500);
nor U23613 (N_23613,N_20121,N_18166);
xor U23614 (N_23614,N_19645,N_19129);
nand U23615 (N_23615,N_18335,N_18851);
xor U23616 (N_23616,N_18246,N_19239);
or U23617 (N_23617,N_20423,N_19288);
nand U23618 (N_23618,N_20655,N_20868);
nor U23619 (N_23619,N_19767,N_20269);
or U23620 (N_23620,N_20140,N_18947);
and U23621 (N_23621,N_18147,N_18118);
nor U23622 (N_23622,N_19410,N_20469);
xnor U23623 (N_23623,N_18897,N_18698);
xor U23624 (N_23624,N_18431,N_19487);
xnor U23625 (N_23625,N_20076,N_20991);
nor U23626 (N_23626,N_18345,N_20340);
nor U23627 (N_23627,N_19102,N_20467);
xnor U23628 (N_23628,N_19057,N_19165);
or U23629 (N_23629,N_20775,N_19655);
nor U23630 (N_23630,N_18274,N_19787);
xor U23631 (N_23631,N_18965,N_20084);
nand U23632 (N_23632,N_19490,N_18813);
nand U23633 (N_23633,N_20691,N_20779);
and U23634 (N_23634,N_18959,N_20514);
nor U23635 (N_23635,N_18967,N_19300);
or U23636 (N_23636,N_19118,N_20274);
nor U23637 (N_23637,N_20145,N_19467);
nand U23638 (N_23638,N_20115,N_20851);
nor U23639 (N_23639,N_19042,N_19897);
nor U23640 (N_23640,N_18986,N_18723);
xor U23641 (N_23641,N_19388,N_20359);
or U23642 (N_23642,N_19123,N_20348);
xnor U23643 (N_23643,N_19376,N_18524);
xor U23644 (N_23644,N_20774,N_20305);
nor U23645 (N_23645,N_20156,N_19456);
xnor U23646 (N_23646,N_19662,N_18288);
nor U23647 (N_23647,N_19745,N_18402);
and U23648 (N_23648,N_20944,N_18911);
or U23649 (N_23649,N_19963,N_19618);
nor U23650 (N_23650,N_19603,N_18303);
nor U23651 (N_23651,N_18820,N_20941);
nand U23652 (N_23652,N_18829,N_20793);
nand U23653 (N_23653,N_20748,N_19827);
or U23654 (N_23654,N_19211,N_20656);
xnor U23655 (N_23655,N_19619,N_18185);
nand U23656 (N_23656,N_18686,N_20515);
or U23657 (N_23657,N_18801,N_19703);
or U23658 (N_23658,N_19083,N_19260);
and U23659 (N_23659,N_20347,N_19354);
xnor U23660 (N_23660,N_19389,N_19954);
and U23661 (N_23661,N_18475,N_19258);
or U23662 (N_23662,N_18237,N_19731);
xor U23663 (N_23663,N_18482,N_18231);
nor U23664 (N_23664,N_20444,N_18836);
xor U23665 (N_23665,N_18960,N_20641);
nand U23666 (N_23666,N_20979,N_19957);
and U23667 (N_23667,N_20745,N_20614);
and U23668 (N_23668,N_18434,N_20858);
xnor U23669 (N_23669,N_20949,N_19103);
and U23670 (N_23670,N_19372,N_20242);
nand U23671 (N_23671,N_19030,N_20894);
nand U23672 (N_23672,N_20316,N_20183);
xnor U23673 (N_23673,N_20119,N_19205);
nand U23674 (N_23674,N_18329,N_19537);
nand U23675 (N_23675,N_19118,N_19143);
xor U23676 (N_23676,N_18756,N_20668);
and U23677 (N_23677,N_18082,N_20617);
nand U23678 (N_23678,N_20757,N_19156);
and U23679 (N_23679,N_19801,N_20445);
nor U23680 (N_23680,N_18855,N_20190);
nand U23681 (N_23681,N_18648,N_18457);
xor U23682 (N_23682,N_18817,N_18858);
xnor U23683 (N_23683,N_19957,N_19489);
or U23684 (N_23684,N_20938,N_20476);
nor U23685 (N_23685,N_20269,N_20518);
and U23686 (N_23686,N_20971,N_19981);
and U23687 (N_23687,N_18118,N_19679);
nand U23688 (N_23688,N_18367,N_19121);
nand U23689 (N_23689,N_20828,N_20019);
xnor U23690 (N_23690,N_19263,N_18539);
and U23691 (N_23691,N_20314,N_18857);
nand U23692 (N_23692,N_19746,N_18434);
nand U23693 (N_23693,N_18143,N_18111);
xnor U23694 (N_23694,N_19496,N_19549);
nor U23695 (N_23695,N_18228,N_20358);
xnor U23696 (N_23696,N_19048,N_18904);
nand U23697 (N_23697,N_20407,N_18519);
nand U23698 (N_23698,N_18463,N_19744);
nor U23699 (N_23699,N_18803,N_19984);
and U23700 (N_23700,N_19917,N_19527);
xor U23701 (N_23701,N_20095,N_20676);
xor U23702 (N_23702,N_18639,N_18805);
nand U23703 (N_23703,N_18741,N_18961);
nand U23704 (N_23704,N_18478,N_19033);
or U23705 (N_23705,N_20089,N_18314);
nor U23706 (N_23706,N_19152,N_18347);
nand U23707 (N_23707,N_20934,N_20427);
nor U23708 (N_23708,N_19322,N_19599);
nor U23709 (N_23709,N_19908,N_20079);
nand U23710 (N_23710,N_18394,N_18872);
nor U23711 (N_23711,N_18540,N_19380);
nand U23712 (N_23712,N_18767,N_18327);
or U23713 (N_23713,N_20632,N_20626);
or U23714 (N_23714,N_19802,N_19882);
and U23715 (N_23715,N_19861,N_20066);
nor U23716 (N_23716,N_19931,N_20546);
or U23717 (N_23717,N_20804,N_18130);
nor U23718 (N_23718,N_19659,N_20253);
xor U23719 (N_23719,N_20578,N_18000);
or U23720 (N_23720,N_20324,N_19834);
or U23721 (N_23721,N_19642,N_20961);
nor U23722 (N_23722,N_19687,N_18370);
and U23723 (N_23723,N_18835,N_19625);
xnor U23724 (N_23724,N_19094,N_20485);
nand U23725 (N_23725,N_18385,N_20310);
and U23726 (N_23726,N_18300,N_20821);
and U23727 (N_23727,N_19937,N_18743);
xnor U23728 (N_23728,N_20262,N_20610);
nor U23729 (N_23729,N_20004,N_18193);
nor U23730 (N_23730,N_19670,N_20706);
nor U23731 (N_23731,N_19179,N_18265);
and U23732 (N_23732,N_19802,N_18837);
and U23733 (N_23733,N_20187,N_19287);
nand U23734 (N_23734,N_18996,N_20584);
nor U23735 (N_23735,N_18095,N_18676);
nor U23736 (N_23736,N_20493,N_18928);
xor U23737 (N_23737,N_20294,N_20395);
or U23738 (N_23738,N_20811,N_18898);
and U23739 (N_23739,N_18849,N_18212);
nor U23740 (N_23740,N_20780,N_20494);
or U23741 (N_23741,N_20906,N_19668);
and U23742 (N_23742,N_18151,N_20827);
xnor U23743 (N_23743,N_18416,N_19021);
xor U23744 (N_23744,N_18882,N_18974);
nor U23745 (N_23745,N_18272,N_19279);
or U23746 (N_23746,N_19200,N_19206);
nand U23747 (N_23747,N_19472,N_20582);
nor U23748 (N_23748,N_18304,N_20462);
and U23749 (N_23749,N_18921,N_19796);
nor U23750 (N_23750,N_20836,N_18661);
or U23751 (N_23751,N_20093,N_20040);
nor U23752 (N_23752,N_20513,N_20792);
nand U23753 (N_23753,N_20341,N_19911);
nor U23754 (N_23754,N_19658,N_18230);
or U23755 (N_23755,N_19384,N_19329);
or U23756 (N_23756,N_18878,N_20955);
nand U23757 (N_23757,N_19750,N_20943);
xnor U23758 (N_23758,N_19176,N_18179);
and U23759 (N_23759,N_18858,N_19407);
nand U23760 (N_23760,N_18970,N_19100);
or U23761 (N_23761,N_20021,N_20993);
or U23762 (N_23762,N_19794,N_19103);
xnor U23763 (N_23763,N_18560,N_18064);
and U23764 (N_23764,N_18687,N_18575);
xor U23765 (N_23765,N_19623,N_18733);
xnor U23766 (N_23766,N_20655,N_19103);
nand U23767 (N_23767,N_19569,N_19088);
xnor U23768 (N_23768,N_20847,N_19538);
nand U23769 (N_23769,N_18989,N_18943);
nand U23770 (N_23770,N_20242,N_20044);
nand U23771 (N_23771,N_19581,N_18177);
nor U23772 (N_23772,N_20313,N_19077);
or U23773 (N_23773,N_19815,N_18138);
nor U23774 (N_23774,N_18114,N_18750);
and U23775 (N_23775,N_18284,N_20992);
nand U23776 (N_23776,N_18378,N_20819);
nand U23777 (N_23777,N_18616,N_19938);
or U23778 (N_23778,N_20060,N_18384);
and U23779 (N_23779,N_20363,N_20623);
or U23780 (N_23780,N_19987,N_20652);
xnor U23781 (N_23781,N_20832,N_18075);
nor U23782 (N_23782,N_19294,N_18555);
and U23783 (N_23783,N_20575,N_18694);
or U23784 (N_23784,N_19605,N_18101);
nand U23785 (N_23785,N_20797,N_19180);
xor U23786 (N_23786,N_18784,N_20979);
xnor U23787 (N_23787,N_20478,N_20158);
nor U23788 (N_23788,N_20647,N_18858);
and U23789 (N_23789,N_20534,N_20754);
nand U23790 (N_23790,N_19873,N_18073);
xnor U23791 (N_23791,N_20751,N_20970);
nand U23792 (N_23792,N_19563,N_20507);
xnor U23793 (N_23793,N_20942,N_19234);
and U23794 (N_23794,N_19570,N_18126);
nand U23795 (N_23795,N_20396,N_18639);
nor U23796 (N_23796,N_19404,N_19931);
nor U23797 (N_23797,N_18847,N_20852);
nand U23798 (N_23798,N_18527,N_18669);
or U23799 (N_23799,N_18147,N_20847);
nand U23800 (N_23800,N_20049,N_18651);
xor U23801 (N_23801,N_19015,N_19771);
nor U23802 (N_23802,N_18240,N_18805);
nand U23803 (N_23803,N_19382,N_20763);
xor U23804 (N_23804,N_19168,N_20994);
nand U23805 (N_23805,N_18556,N_20807);
or U23806 (N_23806,N_20536,N_20841);
nand U23807 (N_23807,N_19062,N_18220);
xor U23808 (N_23808,N_19985,N_19089);
nor U23809 (N_23809,N_18064,N_18102);
nand U23810 (N_23810,N_18266,N_19924);
xor U23811 (N_23811,N_19372,N_20584);
and U23812 (N_23812,N_20930,N_20891);
or U23813 (N_23813,N_20845,N_19620);
nand U23814 (N_23814,N_19938,N_19949);
or U23815 (N_23815,N_19600,N_20837);
or U23816 (N_23816,N_19412,N_18465);
and U23817 (N_23817,N_20051,N_18523);
xnor U23818 (N_23818,N_18566,N_18552);
and U23819 (N_23819,N_18142,N_18433);
nand U23820 (N_23820,N_19200,N_19484);
and U23821 (N_23821,N_18006,N_18189);
and U23822 (N_23822,N_20589,N_19619);
or U23823 (N_23823,N_19345,N_19274);
and U23824 (N_23824,N_19806,N_20680);
xor U23825 (N_23825,N_20950,N_20353);
nand U23826 (N_23826,N_18616,N_19294);
nand U23827 (N_23827,N_19637,N_20938);
nand U23828 (N_23828,N_20079,N_18384);
and U23829 (N_23829,N_19486,N_20557);
nand U23830 (N_23830,N_20277,N_18388);
nand U23831 (N_23831,N_19217,N_20262);
nor U23832 (N_23832,N_19303,N_19317);
nand U23833 (N_23833,N_20547,N_18501);
or U23834 (N_23834,N_20033,N_18844);
nand U23835 (N_23835,N_20355,N_20688);
xnor U23836 (N_23836,N_18482,N_19602);
and U23837 (N_23837,N_18416,N_20588);
or U23838 (N_23838,N_19039,N_18218);
and U23839 (N_23839,N_20103,N_19865);
nor U23840 (N_23840,N_19105,N_19242);
nand U23841 (N_23841,N_20508,N_19223);
nand U23842 (N_23842,N_18793,N_20583);
xnor U23843 (N_23843,N_20697,N_20701);
and U23844 (N_23844,N_19182,N_18227);
xor U23845 (N_23845,N_19050,N_19812);
xnor U23846 (N_23846,N_19697,N_20197);
or U23847 (N_23847,N_19811,N_20546);
nand U23848 (N_23848,N_18645,N_19002);
xor U23849 (N_23849,N_20649,N_18156);
nand U23850 (N_23850,N_19913,N_20226);
xnor U23851 (N_23851,N_18817,N_18310);
and U23852 (N_23852,N_19824,N_19183);
nor U23853 (N_23853,N_18820,N_19748);
nor U23854 (N_23854,N_19410,N_20760);
or U23855 (N_23855,N_20337,N_20011);
and U23856 (N_23856,N_18104,N_18559);
or U23857 (N_23857,N_18532,N_19345);
nand U23858 (N_23858,N_18891,N_18067);
and U23859 (N_23859,N_18244,N_19998);
nor U23860 (N_23860,N_20476,N_20389);
or U23861 (N_23861,N_19508,N_20953);
and U23862 (N_23862,N_20561,N_20599);
xor U23863 (N_23863,N_18654,N_20178);
nand U23864 (N_23864,N_18795,N_19418);
or U23865 (N_23865,N_20559,N_18717);
xnor U23866 (N_23866,N_20248,N_19906);
xor U23867 (N_23867,N_19404,N_19930);
nor U23868 (N_23868,N_20134,N_18661);
nor U23869 (N_23869,N_19856,N_19704);
nand U23870 (N_23870,N_18726,N_20150);
or U23871 (N_23871,N_19242,N_18174);
xnor U23872 (N_23872,N_18660,N_19938);
nand U23873 (N_23873,N_18290,N_20321);
nand U23874 (N_23874,N_20562,N_20721);
or U23875 (N_23875,N_20446,N_18293);
nor U23876 (N_23876,N_20188,N_20420);
and U23877 (N_23877,N_20714,N_19193);
nand U23878 (N_23878,N_20083,N_18641);
or U23879 (N_23879,N_20893,N_20776);
nand U23880 (N_23880,N_18975,N_19884);
or U23881 (N_23881,N_19985,N_18859);
or U23882 (N_23882,N_18731,N_19329);
nand U23883 (N_23883,N_19284,N_20482);
xnor U23884 (N_23884,N_20770,N_18533);
xor U23885 (N_23885,N_19545,N_18302);
or U23886 (N_23886,N_19571,N_18760);
xor U23887 (N_23887,N_20739,N_20702);
or U23888 (N_23888,N_20550,N_18905);
and U23889 (N_23889,N_18668,N_20218);
nand U23890 (N_23890,N_18650,N_20161);
xnor U23891 (N_23891,N_18614,N_19137);
xor U23892 (N_23892,N_20423,N_19145);
and U23893 (N_23893,N_19918,N_19855);
nand U23894 (N_23894,N_20227,N_18302);
and U23895 (N_23895,N_20087,N_18510);
or U23896 (N_23896,N_19383,N_20544);
nand U23897 (N_23897,N_20228,N_19449);
nand U23898 (N_23898,N_20194,N_18987);
xor U23899 (N_23899,N_19914,N_18380);
or U23900 (N_23900,N_20445,N_18599);
nand U23901 (N_23901,N_18133,N_18821);
and U23902 (N_23902,N_19694,N_20533);
nor U23903 (N_23903,N_18440,N_18212);
nor U23904 (N_23904,N_19048,N_19959);
xnor U23905 (N_23905,N_19118,N_19130);
xnor U23906 (N_23906,N_20577,N_20370);
nor U23907 (N_23907,N_18143,N_19336);
nand U23908 (N_23908,N_19217,N_20106);
xor U23909 (N_23909,N_19683,N_20629);
or U23910 (N_23910,N_20544,N_19103);
nand U23911 (N_23911,N_19953,N_18663);
nor U23912 (N_23912,N_20898,N_19197);
xnor U23913 (N_23913,N_20683,N_18602);
or U23914 (N_23914,N_19130,N_20072);
and U23915 (N_23915,N_20906,N_19712);
and U23916 (N_23916,N_20285,N_19306);
and U23917 (N_23917,N_19111,N_18524);
nor U23918 (N_23918,N_19119,N_19715);
or U23919 (N_23919,N_19073,N_18840);
or U23920 (N_23920,N_19181,N_19317);
nor U23921 (N_23921,N_19416,N_18801);
nor U23922 (N_23922,N_19429,N_18412);
nor U23923 (N_23923,N_19413,N_20704);
nor U23924 (N_23924,N_18228,N_19959);
and U23925 (N_23925,N_18823,N_19381);
xor U23926 (N_23926,N_19531,N_20768);
or U23927 (N_23927,N_18637,N_20870);
nand U23928 (N_23928,N_20152,N_18553);
xor U23929 (N_23929,N_18427,N_19144);
xor U23930 (N_23930,N_19639,N_20095);
or U23931 (N_23931,N_20551,N_18896);
and U23932 (N_23932,N_19181,N_18906);
xor U23933 (N_23933,N_20861,N_20628);
or U23934 (N_23934,N_19330,N_19654);
nor U23935 (N_23935,N_19110,N_18314);
or U23936 (N_23936,N_20744,N_18389);
or U23937 (N_23937,N_20224,N_20082);
nand U23938 (N_23938,N_18148,N_20646);
nand U23939 (N_23939,N_20176,N_19421);
nand U23940 (N_23940,N_19354,N_20309);
nor U23941 (N_23941,N_19724,N_20548);
or U23942 (N_23942,N_18359,N_19408);
or U23943 (N_23943,N_20225,N_20793);
nor U23944 (N_23944,N_20505,N_18892);
nand U23945 (N_23945,N_18851,N_18120);
nand U23946 (N_23946,N_19527,N_20204);
nor U23947 (N_23947,N_20118,N_20071);
xor U23948 (N_23948,N_19345,N_18343);
nand U23949 (N_23949,N_19493,N_19117);
nor U23950 (N_23950,N_20249,N_18011);
nor U23951 (N_23951,N_20455,N_20442);
or U23952 (N_23952,N_18499,N_18150);
and U23953 (N_23953,N_20685,N_20559);
nor U23954 (N_23954,N_20457,N_18004);
xor U23955 (N_23955,N_20143,N_19438);
xor U23956 (N_23956,N_20566,N_19776);
or U23957 (N_23957,N_18565,N_20142);
xnor U23958 (N_23958,N_19659,N_19497);
nand U23959 (N_23959,N_18677,N_18534);
xor U23960 (N_23960,N_18797,N_20848);
xnor U23961 (N_23961,N_18215,N_18438);
xor U23962 (N_23962,N_19139,N_20764);
nand U23963 (N_23963,N_18334,N_18756);
nand U23964 (N_23964,N_20402,N_18440);
xor U23965 (N_23965,N_20330,N_19378);
or U23966 (N_23966,N_19324,N_19402);
nand U23967 (N_23967,N_20456,N_19245);
nor U23968 (N_23968,N_19043,N_20923);
nor U23969 (N_23969,N_20988,N_19401);
nor U23970 (N_23970,N_20853,N_20545);
nand U23971 (N_23971,N_19686,N_18518);
or U23972 (N_23972,N_20249,N_19480);
xnor U23973 (N_23973,N_19245,N_20019);
and U23974 (N_23974,N_20239,N_20936);
nand U23975 (N_23975,N_20320,N_19332);
nor U23976 (N_23976,N_19258,N_20718);
xor U23977 (N_23977,N_19417,N_19515);
and U23978 (N_23978,N_20778,N_18063);
nand U23979 (N_23979,N_20612,N_20626);
nand U23980 (N_23980,N_19806,N_20084);
nand U23981 (N_23981,N_18876,N_18194);
xor U23982 (N_23982,N_18870,N_20815);
nand U23983 (N_23983,N_20609,N_20986);
xor U23984 (N_23984,N_20790,N_18861);
or U23985 (N_23985,N_18181,N_20657);
and U23986 (N_23986,N_19565,N_18043);
or U23987 (N_23987,N_20198,N_20180);
nand U23988 (N_23988,N_20231,N_18081);
xnor U23989 (N_23989,N_18415,N_19004);
nand U23990 (N_23990,N_18796,N_19578);
xor U23991 (N_23991,N_19627,N_18968);
nor U23992 (N_23992,N_20438,N_19136);
or U23993 (N_23993,N_18789,N_18912);
or U23994 (N_23994,N_19165,N_19119);
and U23995 (N_23995,N_20125,N_19159);
and U23996 (N_23996,N_18699,N_19919);
nand U23997 (N_23997,N_18253,N_18904);
nor U23998 (N_23998,N_18076,N_19345);
and U23999 (N_23999,N_19772,N_19605);
or U24000 (N_24000,N_21843,N_22585);
and U24001 (N_24001,N_22006,N_21737);
nor U24002 (N_24002,N_21151,N_22948);
xor U24003 (N_24003,N_22038,N_21568);
and U24004 (N_24004,N_23832,N_23483);
nand U24005 (N_24005,N_22844,N_22499);
xnor U24006 (N_24006,N_21941,N_23339);
nor U24007 (N_24007,N_23647,N_22828);
nand U24008 (N_24008,N_21320,N_22895);
or U24009 (N_24009,N_23337,N_21772);
or U24010 (N_24010,N_23012,N_23438);
nand U24011 (N_24011,N_22603,N_22105);
nand U24012 (N_24012,N_21909,N_21088);
xor U24013 (N_24013,N_23713,N_21240);
and U24014 (N_24014,N_23905,N_23096);
nand U24015 (N_24015,N_21628,N_21191);
xor U24016 (N_24016,N_21729,N_23263);
xor U24017 (N_24017,N_22591,N_23535);
or U24018 (N_24018,N_23675,N_21810);
and U24019 (N_24019,N_23506,N_22349);
nor U24020 (N_24020,N_22713,N_21807);
xnor U24021 (N_24021,N_22733,N_23701);
nand U24022 (N_24022,N_23139,N_22057);
or U24023 (N_24023,N_23401,N_22811);
xnor U24024 (N_24024,N_23454,N_21624);
and U24025 (N_24025,N_21434,N_22635);
xnor U24026 (N_24026,N_23459,N_21879);
or U24027 (N_24027,N_22532,N_23710);
nand U24028 (N_24028,N_23502,N_23304);
nor U24029 (N_24029,N_21868,N_23555);
xnor U24030 (N_24030,N_21104,N_23008);
xnor U24031 (N_24031,N_23448,N_23284);
and U24032 (N_24032,N_22595,N_21117);
and U24033 (N_24033,N_21548,N_23296);
nor U24034 (N_24034,N_22695,N_22818);
nor U24035 (N_24035,N_22769,N_22268);
or U24036 (N_24036,N_21108,N_23731);
nor U24037 (N_24037,N_23471,N_21754);
xnor U24038 (N_24038,N_23519,N_21705);
nand U24039 (N_24039,N_22454,N_21346);
xnor U24040 (N_24040,N_21043,N_23033);
nor U24041 (N_24041,N_21045,N_21990);
nor U24042 (N_24042,N_22739,N_21933);
nor U24043 (N_24043,N_21736,N_21822);
and U24044 (N_24044,N_21793,N_21518);
and U24045 (N_24045,N_22484,N_22537);
or U24046 (N_24046,N_23922,N_21247);
nand U24047 (N_24047,N_22605,N_23100);
xor U24048 (N_24048,N_22805,N_21225);
nand U24049 (N_24049,N_23606,N_23679);
xnor U24050 (N_24050,N_22196,N_23940);
nor U24051 (N_24051,N_21918,N_22048);
nand U24052 (N_24052,N_21286,N_22837);
and U24053 (N_24053,N_23219,N_23332);
and U24054 (N_24054,N_22683,N_22181);
nand U24055 (N_24055,N_21188,N_23893);
nor U24056 (N_24056,N_23474,N_21873);
xor U24057 (N_24057,N_21184,N_23997);
nor U24058 (N_24058,N_23255,N_22031);
or U24059 (N_24059,N_23610,N_23685);
or U24060 (N_24060,N_22405,N_22341);
nand U24061 (N_24061,N_21057,N_23035);
and U24062 (N_24062,N_21882,N_23583);
or U24063 (N_24063,N_22479,N_21731);
or U24064 (N_24064,N_21245,N_23865);
nand U24065 (N_24065,N_21641,N_23671);
or U24066 (N_24066,N_21812,N_22620);
and U24067 (N_24067,N_21402,N_23397);
nand U24068 (N_24068,N_21921,N_23258);
nor U24069 (N_24069,N_22997,N_22711);
xnor U24070 (N_24070,N_22018,N_21242);
nor U24071 (N_24071,N_23741,N_21887);
or U24072 (N_24072,N_23120,N_23559);
xnor U24073 (N_24073,N_22988,N_23578);
nor U24074 (N_24074,N_22353,N_22821);
and U24075 (N_24075,N_22530,N_23488);
nor U24076 (N_24076,N_23879,N_22518);
xor U24077 (N_24077,N_22086,N_23913);
nor U24078 (N_24078,N_21886,N_22715);
nor U24079 (N_24079,N_21479,N_23094);
or U24080 (N_24080,N_21620,N_23973);
nand U24081 (N_24081,N_22047,N_21331);
or U24082 (N_24082,N_22602,N_21800);
nand U24083 (N_24083,N_21373,N_22410);
nand U24084 (N_24084,N_21536,N_21858);
and U24085 (N_24085,N_21981,N_23803);
nor U24086 (N_24086,N_21806,N_23440);
nand U24087 (N_24087,N_23492,N_23383);
nor U24088 (N_24088,N_23461,N_22972);
nand U24089 (N_24089,N_22721,N_22355);
xnor U24090 (N_24090,N_21734,N_21257);
and U24091 (N_24091,N_23906,N_21529);
xnor U24092 (N_24092,N_22473,N_23393);
and U24093 (N_24093,N_23058,N_23989);
nor U24094 (N_24094,N_23023,N_21427);
xnor U24095 (N_24095,N_22045,N_23765);
or U24096 (N_24096,N_22426,N_22564);
or U24097 (N_24097,N_23342,N_22124);
nand U24098 (N_24098,N_22166,N_21651);
nand U24099 (N_24099,N_21249,N_22313);
nor U24100 (N_24100,N_22187,N_23453);
or U24101 (N_24101,N_23404,N_23395);
nor U24102 (N_24102,N_22280,N_23788);
nor U24103 (N_24103,N_23573,N_23599);
or U24104 (N_24104,N_21394,N_21369);
or U24105 (N_24105,N_23346,N_22157);
or U24106 (N_24106,N_22016,N_23982);
or U24107 (N_24107,N_21046,N_21011);
xor U24108 (N_24108,N_23861,N_21476);
or U24109 (N_24109,N_22303,N_22394);
or U24110 (N_24110,N_21867,N_21497);
xor U24111 (N_24111,N_23827,N_23752);
nor U24112 (N_24112,N_21673,N_21392);
and U24113 (N_24113,N_23988,N_23247);
nor U24114 (N_24114,N_23612,N_22286);
and U24115 (N_24115,N_23313,N_21998);
and U24116 (N_24116,N_22352,N_22545);
nor U24117 (N_24117,N_23748,N_23884);
and U24118 (N_24118,N_22601,N_22516);
nor U24119 (N_24119,N_21052,N_23436);
or U24120 (N_24120,N_21592,N_21738);
xor U24121 (N_24121,N_22523,N_21743);
nor U24122 (N_24122,N_22368,N_21333);
and U24123 (N_24123,N_21955,N_23807);
nand U24124 (N_24124,N_22522,N_22011);
or U24125 (N_24125,N_21622,N_23031);
or U24126 (N_24126,N_21525,N_21869);
xor U24127 (N_24127,N_23956,N_23880);
nor U24128 (N_24128,N_23895,N_21327);
and U24129 (N_24129,N_23246,N_21038);
nand U24130 (N_24130,N_22279,N_23712);
or U24131 (N_24131,N_22566,N_23787);
xor U24132 (N_24132,N_23717,N_22965);
or U24133 (N_24133,N_22001,N_21398);
and U24134 (N_24134,N_22665,N_23113);
nand U24135 (N_24135,N_23529,N_21894);
nand U24136 (N_24136,N_22727,N_23584);
xor U24137 (N_24137,N_23692,N_22969);
nand U24138 (N_24138,N_23209,N_22232);
xor U24139 (N_24139,N_23472,N_22054);
or U24140 (N_24140,N_21436,N_23550);
xor U24141 (N_24141,N_21376,N_21228);
nand U24142 (N_24142,N_21657,N_22593);
and U24143 (N_24143,N_22346,N_23836);
nor U24144 (N_24144,N_21001,N_23282);
and U24145 (N_24145,N_21156,N_22931);
xnor U24146 (N_24146,N_23540,N_22831);
nand U24147 (N_24147,N_21077,N_22569);
nor U24148 (N_24148,N_23985,N_23727);
nand U24149 (N_24149,N_21189,N_23345);
nand U24150 (N_24150,N_22358,N_22515);
and U24151 (N_24151,N_23766,N_21074);
nor U24152 (N_24152,N_22427,N_21845);
or U24153 (N_24153,N_22804,N_23117);
nand U24154 (N_24154,N_22940,N_23272);
nand U24155 (N_24155,N_22798,N_22779);
nor U24156 (N_24156,N_21898,N_23872);
nor U24157 (N_24157,N_21498,N_22504);
nor U24158 (N_24158,N_22608,N_21647);
nor U24159 (N_24159,N_23622,N_22224);
nand U24160 (N_24160,N_23774,N_21037);
or U24161 (N_24161,N_22924,N_21674);
or U24162 (N_24162,N_23205,N_21839);
and U24163 (N_24163,N_21545,N_22258);
or U24164 (N_24164,N_22501,N_23888);
nand U24165 (N_24165,N_23466,N_23660);
xnor U24166 (N_24166,N_22376,N_21658);
and U24167 (N_24167,N_22478,N_21277);
nand U24168 (N_24168,N_22892,N_23891);
and U24169 (N_24169,N_22551,N_22028);
and U24170 (N_24170,N_23181,N_22203);
and U24171 (N_24171,N_22099,N_21106);
nand U24172 (N_24172,N_21666,N_21337);
or U24173 (N_24173,N_22369,N_22707);
and U24174 (N_24174,N_22442,N_22435);
xor U24175 (N_24175,N_22140,N_22850);
and U24176 (N_24176,N_21913,N_21361);
nand U24177 (N_24177,N_23322,N_23736);
nor U24178 (N_24178,N_22905,N_23743);
and U24179 (N_24179,N_22581,N_23726);
or U24180 (N_24180,N_23870,N_23770);
nand U24181 (N_24181,N_21238,N_21492);
xnor U24182 (N_24182,N_22743,N_21141);
or U24183 (N_24183,N_21127,N_21122);
and U24184 (N_24184,N_21699,N_23078);
nand U24185 (N_24185,N_22982,N_22732);
and U24186 (N_24186,N_23458,N_21484);
nor U24187 (N_24187,N_21103,N_22549);
xnor U24188 (N_24188,N_22383,N_22331);
and U24189 (N_24189,N_22876,N_22158);
nand U24190 (N_24190,N_21595,N_23422);
and U24191 (N_24191,N_22729,N_23953);
nand U24192 (N_24192,N_22451,N_21703);
and U24193 (N_24193,N_21051,N_21632);
nand U24194 (N_24194,N_23202,N_21284);
nand U24195 (N_24195,N_21670,N_22912);
xor U24196 (N_24196,N_22525,N_22423);
and U24197 (N_24197,N_21888,N_23412);
or U24198 (N_24198,N_22781,N_23082);
or U24199 (N_24199,N_22507,N_21421);
nand U24200 (N_24200,N_23235,N_23864);
and U24201 (N_24201,N_21692,N_22030);
or U24202 (N_24202,N_22192,N_22447);
nand U24203 (N_24203,N_23021,N_22907);
xnor U24204 (N_24204,N_22951,N_22643);
nand U24205 (N_24205,N_23268,N_22167);
or U24206 (N_24206,N_22471,N_23541);
nor U24207 (N_24207,N_23848,N_23806);
and U24208 (N_24208,N_23036,N_23330);
and U24209 (N_24209,N_21375,N_21490);
nor U24210 (N_24210,N_23802,N_23556);
xor U24211 (N_24211,N_21943,N_22939);
and U24212 (N_24212,N_22092,N_23961);
or U24213 (N_24213,N_23088,N_23232);
and U24214 (N_24214,N_23248,N_22142);
or U24215 (N_24215,N_21662,N_21062);
or U24216 (N_24216,N_22150,N_21643);
nand U24217 (N_24217,N_22852,N_23210);
nor U24218 (N_24218,N_21811,N_21796);
nor U24219 (N_24219,N_22329,N_22898);
and U24220 (N_24220,N_23747,N_21203);
or U24221 (N_24221,N_23663,N_21708);
or U24222 (N_24222,N_22210,N_21338);
and U24223 (N_24223,N_23965,N_23249);
nand U24224 (N_24224,N_21396,N_23020);
nor U24225 (N_24225,N_21695,N_21672);
or U24226 (N_24226,N_21768,N_22681);
xor U24227 (N_24227,N_21185,N_23421);
or U24228 (N_24228,N_22930,N_21163);
nand U24229 (N_24229,N_22194,N_22734);
nand U24230 (N_24230,N_21216,N_23083);
nand U24231 (N_24231,N_21880,N_23061);
nand U24232 (N_24232,N_21447,N_21220);
and U24233 (N_24233,N_21343,N_22934);
xnor U24234 (N_24234,N_22386,N_22690);
or U24235 (N_24235,N_23237,N_23174);
xnor U24236 (N_24236,N_22847,N_22007);
or U24237 (N_24237,N_23112,N_22223);
or U24238 (N_24238,N_21027,N_22052);
nand U24239 (N_24239,N_22311,N_22785);
nor U24240 (N_24240,N_21610,N_23636);
nand U24241 (N_24241,N_23521,N_22256);
nand U24242 (N_24242,N_23060,N_23121);
xor U24243 (N_24243,N_23341,N_22049);
or U24244 (N_24244,N_22983,N_23030);
xnor U24245 (N_24245,N_21302,N_22385);
xnor U24246 (N_24246,N_23000,N_23990);
or U24247 (N_24247,N_22558,N_23114);
nor U24248 (N_24248,N_21656,N_21168);
and U24249 (N_24249,N_22863,N_22546);
xor U24250 (N_24250,N_22390,N_23552);
xnor U24251 (N_24251,N_21305,N_23010);
or U24252 (N_24252,N_23992,N_22919);
nand U24253 (N_24253,N_21283,N_21136);
xor U24254 (N_24254,N_21391,N_21110);
xor U24255 (N_24255,N_21645,N_22324);
xor U24256 (N_24256,N_22506,N_23075);
xnor U24257 (N_24257,N_23873,N_21453);
xor U24258 (N_24258,N_23126,N_21144);
or U24259 (N_24259,N_22164,N_21970);
nand U24260 (N_24260,N_21988,N_23225);
and U24261 (N_24261,N_21407,N_22925);
xor U24262 (N_24262,N_23143,N_23745);
nor U24263 (N_24263,N_23868,N_23626);
xor U24264 (N_24264,N_21809,N_22335);
xor U24265 (N_24265,N_23242,N_22017);
and U24266 (N_24266,N_21562,N_22922);
or U24267 (N_24267,N_22219,N_22952);
and U24268 (N_24268,N_22340,N_23338);
or U24269 (N_24269,N_21584,N_23199);
or U24270 (N_24270,N_22254,N_22101);
xor U24271 (N_24271,N_22165,N_23821);
xor U24272 (N_24272,N_21769,N_23105);
or U24273 (N_24273,N_23354,N_23382);
xor U24274 (N_24274,N_21615,N_21332);
nand U24275 (N_24275,N_21084,N_21205);
or U24276 (N_24276,N_21488,N_22133);
nor U24277 (N_24277,N_23431,N_21964);
and U24278 (N_24278,N_21432,N_21623);
and U24279 (N_24279,N_22970,N_23028);
xnor U24280 (N_24280,N_23403,N_21905);
nor U24281 (N_24281,N_22191,N_21437);
or U24282 (N_24282,N_23838,N_23238);
xor U24283 (N_24283,N_22422,N_22984);
xnor U24284 (N_24284,N_23823,N_21356);
nand U24285 (N_24285,N_23744,N_22575);
nand U24286 (N_24286,N_23491,N_23718);
and U24287 (N_24287,N_21325,N_22694);
or U24288 (N_24288,N_21388,N_22577);
nand U24289 (N_24289,N_21140,N_23314);
xnor U24290 (N_24290,N_21837,N_21573);
or U24291 (N_24291,N_23193,N_23623);
or U24292 (N_24292,N_21972,N_21158);
or U24293 (N_24293,N_23275,N_22138);
nand U24294 (N_24294,N_23443,N_23359);
or U24295 (N_24295,N_21741,N_21510);
nor U24296 (N_24296,N_23901,N_21834);
nand U24297 (N_24297,N_21187,N_22417);
and U24298 (N_24298,N_21787,N_23358);
or U24299 (N_24299,N_21815,N_21372);
xor U24300 (N_24300,N_22387,N_23596);
and U24301 (N_24301,N_23958,N_23566);
nor U24302 (N_24302,N_23568,N_21702);
and U24303 (N_24303,N_23480,N_22554);
nand U24304 (N_24304,N_22135,N_23994);
xnor U24305 (N_24305,N_23876,N_23650);
nand U24306 (N_24306,N_22307,N_21495);
xor U24307 (N_24307,N_22093,N_21971);
and U24308 (N_24308,N_21274,N_21619);
nand U24309 (N_24309,N_21761,N_21890);
xnor U24310 (N_24310,N_22539,N_21616);
xor U24311 (N_24311,N_22154,N_22883);
nor U24312 (N_24312,N_22758,N_22649);
nor U24313 (N_24313,N_22691,N_23993);
or U24314 (N_24314,N_21637,N_22037);
or U24315 (N_24315,N_21022,N_22866);
and U24316 (N_24316,N_22584,N_22143);
xor U24317 (N_24317,N_21336,N_21359);
or U24318 (N_24318,N_21145,N_21876);
or U24319 (N_24319,N_21340,N_22046);
and U24320 (N_24320,N_21574,N_23089);
xor U24321 (N_24321,N_22638,N_23054);
nor U24322 (N_24322,N_23327,N_21229);
nor U24323 (N_24323,N_22550,N_22686);
nor U24324 (N_24324,N_22418,N_23361);
nand U24325 (N_24325,N_21630,N_21192);
xor U24326 (N_24326,N_23489,N_22594);
xor U24327 (N_24327,N_22889,N_23071);
nor U24328 (N_24328,N_21393,N_22146);
xnor U24329 (N_24329,N_22244,N_22935);
nand U24330 (N_24330,N_23115,N_22231);
or U24331 (N_24331,N_23311,N_23999);
nand U24332 (N_24332,N_23645,N_21980);
or U24333 (N_24333,N_21193,N_22104);
nand U24334 (N_24334,N_23545,N_23977);
xnor U24335 (N_24335,N_23605,N_23980);
or U24336 (N_24336,N_23302,N_22469);
nor U24337 (N_24337,N_23034,N_23525);
nor U24338 (N_24338,N_23380,N_23441);
and U24339 (N_24339,N_22155,N_22110);
or U24340 (N_24340,N_21884,N_23091);
and U24341 (N_24341,N_21554,N_21073);
or U24342 (N_24342,N_21371,N_21795);
nor U24343 (N_24343,N_21138,N_21441);
nor U24344 (N_24344,N_22401,N_21625);
and U24345 (N_24345,N_22238,N_23851);
xor U24346 (N_24346,N_21017,N_22989);
or U24347 (N_24347,N_23926,N_23634);
xnor U24348 (N_24348,N_21048,N_21116);
or U24349 (N_24349,N_23365,N_21297);
nor U24350 (N_24350,N_22810,N_23220);
nor U24351 (N_24351,N_21230,N_22266);
xor U24352 (N_24352,N_23372,N_21999);
xor U24353 (N_24353,N_21491,N_23881);
nor U24354 (N_24354,N_23084,N_21397);
and U24355 (N_24355,N_23804,N_23451);
xnor U24356 (N_24356,N_22100,N_22901);
nor U24357 (N_24357,N_22869,N_23107);
xor U24358 (N_24358,N_21232,N_21314);
nor U24359 (N_24359,N_23577,N_23233);
or U24360 (N_24360,N_23240,N_22115);
xnor U24361 (N_24361,N_21485,N_23355);
nand U24362 (N_24362,N_21728,N_22822);
nand U24363 (N_24363,N_21856,N_23394);
and U24364 (N_24364,N_21865,N_22621);
and U24365 (N_24365,N_22735,N_22958);
nand U24366 (N_24366,N_22626,N_23677);
and U24367 (N_24367,N_22084,N_21758);
nand U24368 (N_24368,N_23859,N_23493);
and U24369 (N_24369,N_23185,N_22689);
nand U24370 (N_24370,N_21661,N_22679);
and U24371 (N_24371,N_23067,N_22589);
nand U24372 (N_24372,N_21493,N_23871);
xnor U24373 (N_24373,N_21313,N_22375);
and U24374 (N_24374,N_22740,N_22816);
or U24375 (N_24375,N_22916,N_21370);
or U24376 (N_24376,N_22528,N_23026);
nor U24377 (N_24377,N_23666,N_22580);
xor U24378 (N_24378,N_22776,N_21358);
nand U24379 (N_24379,N_22913,N_22730);
or U24380 (N_24380,N_22789,N_23822);
nand U24381 (N_24381,N_21442,N_21032);
nand U24382 (N_24382,N_22298,N_23276);
and U24383 (N_24383,N_22672,N_23419);
nand U24384 (N_24384,N_21633,N_21341);
nor U24385 (N_24385,N_23517,N_22206);
nand U24386 (N_24386,N_22867,N_21742);
nor U24387 (N_24387,N_21458,N_21870);
or U24388 (N_24388,N_22719,N_21013);
xnor U24389 (N_24389,N_23102,N_21570);
nand U24390 (N_24390,N_22559,N_22026);
and U24391 (N_24391,N_21475,N_23638);
or U24392 (N_24392,N_23367,N_23188);
and U24393 (N_24393,N_21063,N_22180);
nor U24394 (N_24394,N_23273,N_23122);
xor U24395 (N_24395,N_21601,N_23750);
nand U24396 (N_24396,N_21250,N_22757);
or U24397 (N_24397,N_23749,N_22129);
or U24398 (N_24398,N_22640,N_21408);
and U24399 (N_24399,N_22583,N_21756);
xnor U24400 (N_24400,N_21169,N_21857);
nand U24401 (N_24401,N_23967,N_23810);
and U24402 (N_24402,N_21727,N_23099);
or U24403 (N_24403,N_21794,N_21689);
nand U24404 (N_24404,N_21223,N_23197);
and U24405 (N_24405,N_23644,N_23654);
or U24406 (N_24406,N_21415,N_21569);
nor U24407 (N_24407,N_21326,N_21298);
and U24408 (N_24408,N_23937,N_23189);
and U24409 (N_24409,N_23907,N_22949);
nor U24410 (N_24410,N_21586,N_22887);
nor U24411 (N_24411,N_22490,N_21903);
or U24412 (N_24412,N_23927,N_21801);
and U24413 (N_24413,N_21764,N_23191);
and U24414 (N_24414,N_23963,N_22775);
xnor U24415 (N_24415,N_23446,N_22995);
nand U24416 (N_24416,N_21118,N_23912);
or U24417 (N_24417,N_23811,N_23315);
nor U24418 (N_24418,N_23257,N_22139);
nand U24419 (N_24419,N_23942,N_22910);
xnor U24420 (N_24420,N_21590,N_22412);
or U24421 (N_24421,N_22747,N_21817);
xor U24422 (N_24422,N_23615,N_23594);
or U24423 (N_24423,N_21322,N_23820);
and U24424 (N_24424,N_21792,N_22860);
or U24425 (N_24425,N_21486,N_21607);
nand U24426 (N_24426,N_23839,N_21414);
nand U24427 (N_24427,N_21919,N_21285);
xor U24428 (N_24428,N_22927,N_22010);
xor U24429 (N_24429,N_21838,N_21515);
and U24430 (N_24430,N_23068,N_22202);
or U24431 (N_24431,N_22293,N_22807);
or U24432 (N_24432,N_21818,N_23768);
and U24433 (N_24433,N_22315,N_23914);
and U24434 (N_24434,N_23767,N_21196);
and U24435 (N_24435,N_23348,N_23608);
and U24436 (N_24436,N_21776,N_23487);
or U24437 (N_24437,N_21509,N_21997);
nand U24438 (N_24438,N_21748,N_23563);
xnor U24439 (N_24439,N_23511,N_23156);
nor U24440 (N_24440,N_23005,N_23840);
nor U24441 (N_24441,N_22235,N_22170);
and U24442 (N_24442,N_22568,N_22183);
nor U24443 (N_24443,N_23179,N_21671);
or U24444 (N_24444,N_21197,N_23425);
or U24445 (N_24445,N_22565,N_21199);
and U24446 (N_24446,N_22824,N_22130);
or U24447 (N_24447,N_23037,N_23288);
and U24448 (N_24448,N_21580,N_22343);
nand U24449 (N_24449,N_23389,N_23950);
nor U24450 (N_24450,N_23109,N_22271);
or U24451 (N_24451,N_22669,N_21640);
or U24452 (N_24452,N_23373,N_22270);
xnor U24453 (N_24453,N_22066,N_22119);
xnor U24454 (N_24454,N_21312,N_21502);
xnor U24455 (N_24455,N_21675,N_22731);
xnor U24456 (N_24456,N_21652,N_21556);
xor U24457 (N_24457,N_22704,N_21364);
or U24458 (N_24458,N_22882,N_21377);
nand U24459 (N_24459,N_21280,N_22648);
or U24460 (N_24460,N_21348,N_23386);
xor U24461 (N_24461,N_22718,N_23853);
xor U24462 (N_24462,N_22257,N_22535);
xor U24463 (N_24463,N_23983,N_23539);
nand U24464 (N_24464,N_21900,N_23607);
nor U24465 (N_24465,N_22438,N_21583);
nor U24466 (N_24466,N_23846,N_21953);
xnor U24467 (N_24467,N_21654,N_21066);
xnor U24468 (N_24468,N_21165,N_21938);
or U24469 (N_24469,N_23391,N_21926);
and U24470 (N_24470,N_22406,N_21871);
nor U24471 (N_24471,N_21836,N_22074);
xor U24472 (N_24472,N_21410,N_22696);
nand U24473 (N_24473,N_22710,N_22198);
nor U24474 (N_24474,N_22436,N_21553);
or U24475 (N_24475,N_22547,N_23867);
nand U24476 (N_24476,N_23720,N_23674);
and U24477 (N_24477,N_22096,N_22697);
nand U24478 (N_24478,N_23420,N_22891);
nand U24479 (N_24479,N_23409,N_22020);
and U24480 (N_24480,N_21688,N_23921);
nand U24481 (N_24481,N_23771,N_21342);
or U24482 (N_24482,N_21053,N_23739);
nor U24483 (N_24483,N_22364,N_22023);
nor U24484 (N_24484,N_23271,N_22722);
nor U24485 (N_24485,N_21516,N_22978);
xor U24486 (N_24486,N_23093,N_21157);
nor U24487 (N_24487,N_23408,N_22619);
nor U24488 (N_24488,N_21655,N_23460);
and U24489 (N_24489,N_21904,N_23923);
nor U24490 (N_24490,N_23298,N_23007);
or U24491 (N_24491,N_23123,N_23176);
nor U24492 (N_24492,N_21496,N_22864);
and U24493 (N_24493,N_23402,N_21842);
nand U24494 (N_24494,N_21696,N_22906);
xnor U24495 (N_24495,N_22795,N_21029);
and U24496 (N_24496,N_22639,N_22136);
or U24497 (N_24497,N_22114,N_21296);
or U24498 (N_24498,N_21010,N_23129);
xor U24499 (N_24499,N_23567,N_23548);
nand U24500 (N_24500,N_21086,N_23633);
nor U24501 (N_24501,N_22742,N_23207);
xnor U24502 (N_24502,N_23855,N_21922);
xor U24503 (N_24503,N_23597,N_21786);
nor U24504 (N_24504,N_21541,N_21676);
and U24505 (N_24505,N_22560,N_21306);
nand U24506 (N_24506,N_21942,N_23587);
nand U24507 (N_24507,N_23920,N_21978);
xnor U24508 (N_24508,N_23503,N_21715);
nor U24509 (N_24509,N_23824,N_22217);
nor U24510 (N_24510,N_22652,N_21613);
nor U24511 (N_24511,N_21224,N_22644);
nand U24512 (N_24512,N_21966,N_23135);
nand U24513 (N_24513,N_23643,N_21149);
nor U24514 (N_24514,N_22737,N_23212);
xor U24515 (N_24515,N_23090,N_21956);
nor U24516 (N_24516,N_23433,N_21469);
and U24517 (N_24517,N_21821,N_21512);
nor U24518 (N_24518,N_21299,N_23763);
nand U24519 (N_24519,N_21125,N_22574);
xnor U24520 (N_24520,N_21522,N_22926);
xnor U24521 (N_24521,N_23226,N_22261);
or U24522 (N_24522,N_23581,N_22008);
nor U24523 (N_24523,N_22182,N_23106);
nand U24524 (N_24524,N_21456,N_22102);
and U24525 (N_24525,N_22365,N_23400);
and U24526 (N_24526,N_22236,N_23092);
nand U24527 (N_24527,N_21540,N_23399);
nor U24528 (N_24528,N_21547,N_21252);
or U24529 (N_24529,N_22529,N_23025);
nor U24530 (N_24530,N_23696,N_23551);
nand U24531 (N_24531,N_22842,N_21862);
xor U24532 (N_24532,N_23343,N_23831);
or U24533 (N_24533,N_22189,N_21925);
nor U24534 (N_24534,N_22441,N_22128);
or U24535 (N_24535,N_21099,N_23877);
or U24536 (N_24536,N_23715,N_21602);
nand U24537 (N_24537,N_22637,N_21146);
nand U24538 (N_24538,N_21021,N_22841);
or U24539 (N_24539,N_23772,N_21438);
and U24540 (N_24540,N_23863,N_23168);
xnor U24541 (N_24541,N_22033,N_21629);
xor U24542 (N_24542,N_23267,N_23569);
nor U24543 (N_24543,N_21321,N_21896);
and U24544 (N_24544,N_23457,N_21113);
or U24545 (N_24545,N_23632,N_22803);
nand U24546 (N_24546,N_21425,N_21155);
nor U24547 (N_24547,N_23667,N_21444);
nor U24548 (N_24548,N_23779,N_22370);
or U24549 (N_24549,N_21235,N_23172);
or U24550 (N_24550,N_21000,N_21684);
and U24551 (N_24551,N_23854,N_21974);
nand U24552 (N_24552,N_21080,N_22751);
nor U24553 (N_24553,N_22242,N_23790);
or U24554 (N_24554,N_23924,N_23479);
xor U24555 (N_24555,N_22087,N_23547);
and U24556 (N_24556,N_21362,N_22322);
nand U24557 (N_24557,N_22943,N_23719);
and U24558 (N_24558,N_21773,N_23843);
and U24559 (N_24559,N_21650,N_22024);
and U24560 (N_24560,N_21931,N_21098);
nor U24561 (N_24561,N_22726,N_23494);
xor U24562 (N_24562,N_23277,N_22072);
nor U24563 (N_24563,N_22362,N_23507);
or U24564 (N_24564,N_22896,N_22409);
and U24565 (N_24565,N_23661,N_22708);
nand U24566 (N_24566,N_21450,N_22274);
xnor U24567 (N_24567,N_21937,N_22019);
and U24568 (N_24568,N_23501,N_22306);
nor U24569 (N_24569,N_23513,N_23270);
or U24570 (N_24570,N_22941,N_21068);
nand U24571 (N_24571,N_21791,N_23481);
nor U24572 (N_24572,N_22900,N_23110);
or U24573 (N_24573,N_21952,N_21928);
nand U24574 (N_24574,N_23857,N_21293);
or U24575 (N_24575,N_21244,N_21288);
nor U24576 (N_24576,N_22034,N_22282);
nor U24577 (N_24577,N_23706,N_23320);
or U24578 (N_24578,N_21642,N_23392);
nor U24579 (N_24579,N_21023,N_22163);
and U24580 (N_24580,N_22389,N_22373);
and U24581 (N_24581,N_22381,N_21464);
nor U24582 (N_24582,N_21404,N_21152);
xor U24583 (N_24583,N_21959,N_23885);
xor U24584 (N_24584,N_22339,N_21531);
nor U24585 (N_24585,N_22653,N_21069);
xnor U24586 (N_24586,N_23261,N_22495);
or U24587 (N_24587,N_23149,N_21055);
xnor U24588 (N_24588,N_21639,N_22402);
and U24589 (N_24589,N_22494,N_23616);
or U24590 (N_24590,N_22687,N_23201);
xor U24591 (N_24591,N_23730,N_21065);
or U24592 (N_24592,N_23150,N_22009);
nand U24593 (N_24593,N_21714,N_21911);
nor U24594 (N_24594,N_21363,N_21949);
nor U24595 (N_24595,N_22325,N_22521);
or U24596 (N_24596,N_22336,N_21008);
nor U24597 (N_24597,N_23652,N_23310);
and U24598 (N_24598,N_23844,N_21054);
and U24599 (N_24599,N_22706,N_23930);
xnor U24600 (N_24600,N_21221,N_21423);
and U24601 (N_24601,N_22897,N_23649);
xor U24602 (N_24602,N_21091,N_23522);
and U24603 (N_24603,N_21443,N_23709);
nand U24604 (N_24604,N_21649,N_23592);
nor U24605 (N_24605,N_23673,N_21454);
xnor U24606 (N_24606,N_22050,N_23689);
nor U24607 (N_24607,N_22498,N_23957);
xnor U24608 (N_24608,N_21016,N_21269);
and U24609 (N_24609,N_22668,N_21912);
or U24610 (N_24610,N_21109,N_21452);
nand U24611 (N_24611,N_21004,N_23256);
xnor U24612 (N_24612,N_23669,N_22461);
nand U24613 (N_24613,N_21160,N_21534);
and U24614 (N_24614,N_21691,N_21874);
nor U24615 (N_24615,N_22027,N_21135);
xor U24616 (N_24616,N_21906,N_22979);
nor U24617 (N_24617,N_23076,N_21612);
xor U24618 (N_24618,N_23196,N_21006);
nor U24619 (N_24619,N_22269,N_22411);
or U24620 (N_24620,N_23722,N_22862);
xor U24621 (N_24621,N_23444,N_23141);
nor U24622 (N_24622,N_21164,N_21889);
nand U24623 (N_24623,N_21483,N_21722);
or U24624 (N_24624,N_23154,N_21350);
or U24625 (N_24625,N_21026,N_22162);
xor U24626 (N_24626,N_22357,N_21753);
and U24627 (N_24627,N_21272,N_21174);
nand U24628 (N_24628,N_21982,N_22300);
xnor U24629 (N_24629,N_22861,N_21877);
xnor U24630 (N_24630,N_23948,N_22439);
and U24631 (N_24631,N_21544,N_21031);
xnor U24632 (N_24632,N_23295,N_23307);
or U24633 (N_24633,N_22745,N_23236);
nand U24634 (N_24634,N_21351,N_21543);
or U24635 (N_24635,N_22873,N_23254);
nand U24636 (N_24636,N_22556,N_22042);
or U24637 (N_24637,N_22216,N_21207);
and U24638 (N_24638,N_22004,N_21218);
or U24639 (N_24639,N_21173,N_22415);
xor U24640 (N_24640,N_22197,N_23016);
or U24641 (N_24641,N_22041,N_23160);
xnor U24642 (N_24642,N_23875,N_22082);
nand U24643 (N_24643,N_22538,N_23059);
nand U24644 (N_24644,N_21819,N_22434);
and U24645 (N_24645,N_23782,N_22627);
and U24646 (N_24646,N_21598,N_22520);
and U24647 (N_24647,N_22814,N_21646);
nor U24648 (N_24648,N_21582,N_21147);
or U24649 (N_24649,N_22929,N_22448);
and U24650 (N_24650,N_23833,N_23445);
nand U24651 (N_24651,N_21899,N_22076);
nor U24652 (N_24652,N_22746,N_22043);
nor U24653 (N_24653,N_22334,N_22308);
or U24654 (N_24654,N_23182,N_23362);
nand U24655 (N_24655,N_22172,N_21690);
or U24656 (N_24656,N_22617,N_22126);
nor U24657 (N_24657,N_22994,N_22328);
xnor U24658 (N_24658,N_21506,N_22002);
and U24659 (N_24659,N_21075,N_22380);
xor U24660 (N_24660,N_22089,N_22276);
nand U24661 (N_24661,N_21210,N_22458);
nand U24662 (N_24662,N_21947,N_21575);
xor U24663 (N_24663,N_22625,N_22613);
and U24664 (N_24664,N_23618,N_23009);
xnor U24665 (N_24665,N_22659,N_23686);
nor U24666 (N_24666,N_21571,N_22947);
xnor U24667 (N_24667,N_23159,N_23066);
nand U24668 (N_24668,N_22788,N_22749);
xnor U24669 (N_24669,N_23700,N_23672);
and U24670 (N_24670,N_23514,N_21460);
nand U24671 (N_24671,N_22067,N_23878);
xnor U24672 (N_24672,N_22337,N_21090);
nand U24673 (N_24673,N_23786,N_22845);
xor U24674 (N_24674,N_23648,N_21526);
and U24675 (N_24675,N_22207,N_23439);
nor U24676 (N_24676,N_21115,N_21480);
xnor U24677 (N_24677,N_23909,N_22567);
nor U24678 (N_24678,N_21587,N_23097);
nor U24679 (N_24679,N_21324,N_22933);
nor U24680 (N_24680,N_22314,N_22440);
or U24681 (N_24681,N_22806,N_23406);
nand U24682 (N_24682,N_21246,N_21166);
and U24683 (N_24683,N_21605,N_22060);
or U24684 (N_24684,N_21344,N_23305);
nor U24685 (N_24685,N_23370,N_22616);
or U24686 (N_24686,N_22481,N_23369);
and U24687 (N_24687,N_21328,N_23428);
nand U24688 (N_24688,N_23835,N_22075);
and U24689 (N_24689,N_21585,N_21386);
or U24690 (N_24690,N_23022,N_21994);
nor U24691 (N_24691,N_21832,N_21712);
and U24692 (N_24692,N_21019,N_23152);
and U24693 (N_24693,N_22367,N_23147);
xnor U24694 (N_24694,N_23473,N_21309);
or U24695 (N_24695,N_22836,N_23769);
nor U24696 (N_24696,N_21180,N_23918);
nand U24697 (N_24697,N_22774,N_23326);
or U24698 (N_24698,N_21775,N_21102);
xor U24699 (N_24699,N_23746,N_21783);
xnor U24700 (N_24700,N_22452,N_22241);
or U24701 (N_24701,N_21957,N_21946);
nand U24702 (N_24702,N_21901,N_21170);
and U24703 (N_24703,N_22599,N_21194);
or U24704 (N_24704,N_21271,N_22541);
nand U24705 (N_24705,N_21308,N_23817);
nand U24706 (N_24706,N_23269,N_22973);
or U24707 (N_24707,N_23262,N_22077);
and U24708 (N_24708,N_23469,N_21875);
nand U24709 (N_24709,N_23534,N_21501);
or U24710 (N_24710,N_21852,N_22121);
xor U24711 (N_24711,N_21700,N_21399);
xnor U24712 (N_24712,N_23975,N_22786);
nand U24713 (N_24713,N_23253,N_23155);
xor U24714 (N_24714,N_23659,N_22808);
xnor U24715 (N_24715,N_21007,N_23218);
nor U24716 (N_24716,N_22682,N_22996);
nand U24717 (N_24717,N_21716,N_23974);
or U24718 (N_24718,N_22243,N_22797);
nand U24719 (N_24719,N_21766,N_22486);
and U24720 (N_24720,N_23496,N_23866);
nor U24721 (N_24721,N_23676,N_22051);
nand U24722 (N_24722,N_22483,N_23784);
nand U24723 (N_24723,N_22275,N_21785);
and U24724 (N_24724,N_22199,N_22354);
and U24725 (N_24725,N_22179,N_23664);
nand U24726 (N_24726,N_21467,N_23011);
nor U24727 (N_24727,N_22646,N_21255);
and U24728 (N_24728,N_21089,N_22693);
or U24729 (N_24729,N_21291,N_22145);
and U24730 (N_24730,N_23301,N_22661);
and U24731 (N_24731,N_23228,N_23613);
nand U24732 (N_24732,N_22248,N_22169);
xor U24733 (N_24733,N_21033,N_22312);
xor U24734 (N_24734,N_22466,N_21261);
and U24735 (N_24735,N_23111,N_23477);
xor U24736 (N_24736,N_22633,N_21891);
nor U24737 (N_24737,N_23385,N_22073);
nor U24738 (N_24738,N_21494,N_22628);
xor U24739 (N_24739,N_21621,N_22514);
xor U24740 (N_24740,N_21694,N_22295);
xor U24741 (N_24741,N_23572,N_22908);
nor U24742 (N_24742,N_21975,N_21470);
or U24743 (N_24743,N_22420,N_23278);
or U24744 (N_24744,N_23933,N_21558);
or U24745 (N_24745,N_21720,N_23427);
and U24746 (N_24746,N_22622,N_23001);
nor U24747 (N_24747,N_23486,N_21093);
or U24748 (N_24748,N_22975,N_22480);
xnor U24749 (N_24749,N_22347,N_23274);
nand U24750 (N_24750,N_23542,N_21028);
nand U24751 (N_24751,N_23095,N_23103);
or U24752 (N_24752,N_21798,N_21914);
or U24753 (N_24753,N_22398,N_22954);
or U24754 (N_24754,N_23729,N_23442);
nor U24755 (N_24755,N_22517,N_21428);
and U24756 (N_24756,N_23565,N_22122);
or U24757 (N_24757,N_23124,N_21927);
and U24758 (N_24758,N_23387,N_21183);
nor U24759 (N_24759,N_23418,N_22156);
nor U24760 (N_24760,N_22809,N_23751);
xor U24761 (N_24761,N_21850,N_23721);
nand U24762 (N_24762,N_23708,N_22579);
nand U24763 (N_24763,N_22526,N_23485);
or U24764 (N_24764,N_22701,N_21706);
or U24765 (N_24765,N_22342,N_21014);
nor U24766 (N_24766,N_22429,N_22416);
xor U24767 (N_24767,N_21167,N_21846);
xnor U24768 (N_24768,N_21365,N_23785);
xor U24769 (N_24769,N_21500,N_23497);
and U24770 (N_24770,N_22147,N_23482);
xor U24771 (N_24771,N_21239,N_21555);
xnor U24772 (N_24772,N_21219,N_21808);
nand U24773 (N_24773,N_21087,N_21440);
or U24774 (N_24774,N_21175,N_21413);
xnor U24775 (N_24775,N_22868,N_23898);
and U24776 (N_24776,N_21148,N_22819);
nand U24777 (N_24777,N_22080,N_21233);
xor U24778 (N_24778,N_21781,N_21626);
or U24779 (N_24779,N_21711,N_22851);
or U24780 (N_24780,N_21523,N_21311);
nor U24781 (N_24781,N_22460,N_21532);
or U24782 (N_24782,N_22309,N_22305);
or U24783 (N_24783,N_23316,N_21726);
and U24784 (N_24784,N_22921,N_21668);
xor U24785 (N_24785,N_23964,N_23705);
and U24786 (N_24786,N_22228,N_21917);
nand U24787 (N_24787,N_22467,N_21119);
nand U24788 (N_24788,N_22724,N_23002);
nand U24789 (N_24789,N_21248,N_23306);
and U24790 (N_24790,N_22208,N_23834);
nand U24791 (N_24791,N_22784,N_23175);
nand U24792 (N_24792,N_23946,N_21861);
and U24793 (N_24793,N_23498,N_22610);
nor U24794 (N_24794,N_21360,N_22025);
nand U24795 (N_24795,N_23388,N_22264);
nor U24796 (N_24796,N_22875,N_22185);
nor U24797 (N_24797,N_23962,N_22759);
xnor U24798 (N_24798,N_21455,N_22959);
or U24799 (N_24799,N_23432,N_22766);
xnor U24800 (N_24800,N_22160,N_23783);
nand U24801 (N_24801,N_23919,N_21749);
nor U24802 (N_24802,N_21967,N_23416);
nor U24803 (N_24803,N_23941,N_21566);
and U24804 (N_24804,N_21383,N_22496);
xor U24805 (N_24805,N_21143,N_21064);
nand U24806 (N_24806,N_23104,N_22920);
or U24807 (N_24807,N_22582,N_23300);
and U24808 (N_24808,N_23826,N_21385);
nor U24809 (N_24809,N_23098,N_23371);
nand U24810 (N_24810,N_23725,N_22465);
nor U24811 (N_24811,N_23625,N_23915);
nand U24812 (N_24812,N_22321,N_23575);
nand U24813 (N_24813,N_21256,N_22193);
nand U24814 (N_24814,N_23687,N_22878);
xor U24815 (N_24815,N_23936,N_22720);
or U24816 (N_24816,N_22598,N_23886);
and U24817 (N_24817,N_21685,N_21560);
xnor U24818 (N_24818,N_23003,N_21463);
nand U24819 (N_24819,N_22174,N_22753);
and U24820 (N_24820,N_23733,N_22472);
xnor U24821 (N_24821,N_23704,N_23134);
xor U24822 (N_24822,N_21317,N_22061);
nor U24823 (N_24823,N_21171,N_22717);
and U24824 (N_24824,N_22615,N_21723);
nor U24825 (N_24825,N_23598,N_23976);
and U24826 (N_24826,N_22725,N_22801);
nand U24827 (N_24827,N_21567,N_22378);
nand U24828 (N_24828,N_22990,N_21231);
xor U24829 (N_24829,N_23812,N_23852);
or U24830 (N_24830,N_21020,N_21984);
and U24831 (N_24831,N_22956,N_22297);
or U24832 (N_24832,N_23423,N_22316);
nor U24833 (N_24833,N_21667,N_22200);
xor U24834 (N_24834,N_21847,N_21504);
nand U24835 (N_24835,N_21503,N_21517);
xor U24836 (N_24836,N_22310,N_21648);
and U24837 (N_24837,N_22557,N_21301);
nand U24838 (N_24838,N_22606,N_22457);
or U24839 (N_24839,N_21508,N_22787);
nor U24840 (N_24840,N_23825,N_21680);
nand U24841 (N_24841,N_23533,N_23214);
or U24842 (N_24842,N_22407,N_23850);
xnor U24843 (N_24843,N_22985,N_22301);
nand U24844 (N_24844,N_21131,N_21907);
nand U24845 (N_24845,N_23987,N_22500);
nand U24846 (N_24846,N_23795,N_21934);
xnor U24847 (N_24847,N_23981,N_23579);
or U24848 (N_24848,N_23690,N_23972);
and U24849 (N_24849,N_22083,N_22113);
nor U24850 (N_24850,N_21588,N_21289);
xor U24851 (N_24851,N_22587,N_22449);
nor U24852 (N_24852,N_21549,N_22796);
and U24853 (N_24853,N_21709,N_22437);
or U24854 (N_24854,N_23984,N_23118);
xnor U24855 (N_24855,N_23164,N_23334);
nand U24856 (N_24856,N_22493,N_23178);
nand U24857 (N_24857,N_23619,N_22573);
xnor U24858 (N_24858,N_21268,N_21211);
or U24859 (N_24859,N_21996,N_22453);
nor U24860 (N_24860,N_23221,N_21349);
xor U24861 (N_24861,N_22408,N_22144);
nor U24862 (N_24862,N_22848,N_23781);
or U24863 (N_24863,N_22252,N_23366);
nand U24864 (N_24864,N_23308,N_22664);
and U24865 (N_24865,N_23761,N_22967);
nor U24866 (N_24866,N_21263,N_23849);
xnor U24867 (N_24867,N_22317,N_23350);
nor U24868 (N_24868,N_22230,N_22957);
xor U24869 (N_24869,N_21514,N_21212);
nor U24870 (N_24870,N_21561,N_23490);
and U24871 (N_24871,N_22190,N_23052);
xnor U24872 (N_24872,N_21181,N_22221);
xor U24873 (N_24873,N_21653,N_23291);
or U24874 (N_24874,N_22215,N_21542);
nand U24875 (N_24875,N_22815,N_23171);
and U24876 (N_24876,N_23437,N_22259);
and U24877 (N_24877,N_23133,N_23591);
xnor U24878 (N_24878,N_21330,N_21993);
xnor U24879 (N_24879,N_23153,N_22212);
xnor U24880 (N_24880,N_23882,N_22040);
nand U24881 (N_24881,N_21802,N_21260);
and U24882 (N_24882,N_21422,N_23234);
nor U24883 (N_24883,N_22600,N_21316);
or U24884 (N_24884,N_22107,N_21679);
nor U24885 (N_24885,N_23703,N_23303);
nor U24886 (N_24886,N_22971,N_23792);
nor U24887 (N_24887,N_22044,N_21760);
or U24888 (N_24888,N_21693,N_22890);
xor U24889 (N_24889,N_21384,N_22548);
nor U24890 (N_24890,N_21035,N_22081);
and U24891 (N_24891,N_22656,N_23955);
or U24892 (N_24892,N_23131,N_21669);
nor U24893 (N_24893,N_21600,N_21347);
nor U24894 (N_24894,N_22813,N_21664);
xnor U24895 (N_24895,N_22508,N_23215);
nor U24896 (N_24896,N_21264,N_22263);
nor U24897 (N_24897,N_21446,N_21368);
and U24898 (N_24898,N_22222,N_23691);
and U24899 (N_24899,N_23951,N_23759);
and U24900 (N_24900,N_22287,N_21418);
nand U24901 (N_24901,N_22251,N_23127);
and U24902 (N_24902,N_21426,N_23630);
xor U24903 (N_24903,N_23186,N_21482);
nand U24904 (N_24904,N_22790,N_21161);
or U24905 (N_24905,N_23800,N_23816);
and U24906 (N_24906,N_21039,N_21465);
nand U24907 (N_24907,N_23830,N_21732);
nor U24908 (N_24908,N_22445,N_21050);
xor U24909 (N_24909,N_23101,N_22562);
xnor U24910 (N_24910,N_22932,N_21036);
nand U24911 (N_24911,N_22382,N_21539);
nand U24912 (N_24912,N_22944,N_22768);
xnor U24913 (N_24913,N_21854,N_23137);
nand U24914 (N_24914,N_21100,N_22421);
nor U24915 (N_24915,N_22470,N_22915);
or U24916 (N_24916,N_21058,N_22247);
or U24917 (N_24917,N_23239,N_21594);
nand U24918 (N_24918,N_21757,N_22304);
nor U24919 (N_24919,N_22761,N_21559);
and U24920 (N_24920,N_22563,N_23244);
nor U24921 (N_24921,N_21072,N_22095);
nor U24922 (N_24922,N_22950,N_21527);
or U24923 (N_24923,N_23537,N_22120);
and U24924 (N_24924,N_23006,N_21908);
nor U24925 (N_24925,N_22670,N_23206);
nor U24926 (N_24926,N_21079,N_23694);
nor U24927 (N_24927,N_22741,N_22112);
xor U24928 (N_24928,N_21430,N_21718);
nand U24929 (N_24929,N_21082,N_23841);
and U24930 (N_24930,N_21581,N_22063);
or U24931 (N_24931,N_23695,N_21387);
nor U24932 (N_24932,N_22777,N_23047);
and U24933 (N_24933,N_22502,N_22879);
xor U24934 (N_24934,N_21034,N_23161);
and U24935 (N_24935,N_22756,N_22464);
nor U24936 (N_24936,N_21797,N_22590);
nor U24937 (N_24937,N_23063,N_22642);
and U24938 (N_24938,N_21081,N_23693);
nor U24939 (N_24939,N_23899,N_21634);
nor U24940 (N_24940,N_23187,N_22791);
nor U24941 (N_24941,N_21986,N_22800);
nand U24942 (N_24942,N_21892,N_23162);
and U24943 (N_24943,N_23508,N_21251);
nand U24944 (N_24944,N_23411,N_23357);
nor U24945 (N_24945,N_21855,N_22835);
or U24946 (N_24946,N_21603,N_21751);
nor U24947 (N_24947,N_22062,N_23190);
and U24948 (N_24948,N_22705,N_22655);
and U24949 (N_24949,N_22782,N_23564);
nand U24950 (N_24950,N_23157,N_23390);
xor U24951 (N_24951,N_23655,N_21121);
or U24952 (N_24952,N_21924,N_22854);
nor U24953 (N_24953,N_22384,N_23050);
or U24954 (N_24954,N_22272,N_22292);
nand U24955 (N_24955,N_22176,N_23019);
xnor U24956 (N_24956,N_23292,N_21770);
and U24957 (N_24957,N_21995,N_23527);
nor U24958 (N_24958,N_22645,N_21593);
xor U24959 (N_24959,N_22123,N_21379);
or U24960 (N_24960,N_22685,N_23954);
xnor U24961 (N_24961,N_21267,N_23158);
and U24962 (N_24962,N_21969,N_21774);
nor U24963 (N_24963,N_21958,N_21950);
and U24964 (N_24964,N_21897,N_23978);
xnor U24965 (N_24965,N_22036,N_23132);
or U24966 (N_24966,N_23072,N_23499);
xnor U24967 (N_24967,N_23723,N_23758);
nor U24968 (N_24968,N_21335,N_21697);
xor U24969 (N_24969,N_22468,N_22253);
xnor U24970 (N_24970,N_23080,N_23931);
xor U24971 (N_24971,N_22379,N_23195);
xor U24972 (N_24972,N_21258,N_21154);
and U24973 (N_24973,N_23762,N_21977);
xnor U24974 (N_24974,N_21419,N_23331);
xnor U24975 (N_24975,N_21777,N_23053);
nor U24976 (N_24976,N_23966,N_23018);
xor U24977 (N_24977,N_21707,N_21417);
xnor U24978 (N_24978,N_21150,N_21353);
xor U24979 (N_24979,N_23546,N_23165);
nor U24980 (N_24980,N_21190,N_23532);
nand U24981 (N_24981,N_23216,N_23860);
nor U24982 (N_24982,N_21429,N_23198);
nand U24983 (N_24983,N_21049,N_21803);
nor U24984 (N_24984,N_23789,N_23808);
nor U24985 (N_24985,N_22013,N_21468);
and U24986 (N_24986,N_21281,N_21577);
nand U24987 (N_24987,N_21965,N_23264);
xor U24988 (N_24988,N_23760,N_22474);
nand U24989 (N_24989,N_21784,N_22987);
nor U24990 (N_24990,N_22543,N_22963);
or U24991 (N_24991,N_22961,N_21816);
or U24992 (N_24992,N_21883,N_23398);
and U24993 (N_24993,N_23476,N_21733);
and U24994 (N_24994,N_21389,N_21241);
xor U24995 (N_24995,N_23818,N_22278);
xnor U24996 (N_24996,N_23177,N_21287);
or U24997 (N_24997,N_23504,N_21354);
nor U24998 (N_24998,N_23637,N_22318);
nor U24999 (N_24999,N_23805,N_21962);
nand U25000 (N_25000,N_21449,N_23883);
xor U25001 (N_25001,N_22475,N_22168);
xnor U25002 (N_25002,N_21745,N_23862);
and U25003 (N_25003,N_22624,N_21782);
nand U25004 (N_25004,N_21872,N_21823);
nor U25005 (N_25005,N_22700,N_22870);
and U25006 (N_25006,N_23553,N_22512);
nor U25007 (N_25007,N_23995,N_23842);
and U25008 (N_25008,N_23593,N_23815);
nand U25009 (N_25009,N_21095,N_23478);
or U25010 (N_25010,N_22955,N_21961);
and U25011 (N_25011,N_21114,N_22676);
nor U25012 (N_25012,N_23538,N_23754);
nor U25013 (N_25013,N_22109,N_22899);
nand U25014 (N_25014,N_22032,N_23904);
xor U25015 (N_25015,N_23684,N_23764);
and U25016 (N_25016,N_22663,N_22923);
nor U25017 (N_25017,N_22476,N_21985);
nand U25018 (N_25018,N_22106,N_22127);
and U25019 (N_25019,N_21944,N_21829);
nand U25020 (N_25020,N_22859,N_22834);
or U25021 (N_25021,N_22999,N_23756);
xor U25022 (N_25022,N_23595,N_22237);
nand U25023 (N_25023,N_22489,N_23702);
or U25024 (N_25024,N_21878,N_22607);
and U25025 (N_25025,N_23375,N_23475);
and U25026 (N_25026,N_22576,N_23939);
nand U25027 (N_25027,N_23929,N_21755);
nand U25028 (N_25028,N_21724,N_21932);
nand U25029 (N_25029,N_23151,N_23325);
xnor U25030 (N_25030,N_21094,N_21002);
nand U25031 (N_25031,N_23169,N_23925);
or U25032 (N_25032,N_22444,N_21217);
nor U25033 (N_25033,N_23585,N_21750);
xnor U25034 (N_25034,N_21382,N_22059);
nand U25035 (N_25035,N_22513,N_22209);
nor U25036 (N_25036,N_22511,N_21951);
xor U25037 (N_25037,N_22673,N_21790);
xor U25038 (N_25038,N_23353,N_23140);
nor U25039 (N_25039,N_21111,N_22942);
xor U25040 (N_25040,N_23297,N_21178);
or U25041 (N_25041,N_22881,N_22424);
or U25042 (N_25042,N_21195,N_21923);
nand U25043 (N_25043,N_21830,N_21162);
nor U25044 (N_25044,N_21462,N_21227);
nor U25045 (N_25045,N_21259,N_21983);
nand U25046 (N_25046,N_23424,N_23631);
nor U25047 (N_25047,N_21176,N_23737);
and U25048 (N_25048,N_21935,N_22246);
nor U25049 (N_25049,N_21433,N_22363);
xnor U25050 (N_25050,N_21735,N_23680);
nor U25051 (N_25051,N_22413,N_23108);
nor U25052 (N_25052,N_23653,N_22641);
or U25053 (N_25053,N_21902,N_23735);
and U25054 (N_25054,N_23250,N_23430);
nand U25055 (N_25055,N_23280,N_22799);
or U25056 (N_25056,N_22015,N_23874);
and U25057 (N_25057,N_22712,N_23699);
nand U25058 (N_25058,N_21499,N_23658);
and U25059 (N_25059,N_21609,N_23470);
nand U25060 (N_25060,N_22960,N_23074);
xor U25061 (N_25061,N_21355,N_22736);
and U25062 (N_25062,N_22071,N_23038);
nand U25063 (N_25063,N_23589,N_21519);
nand U25064 (N_25064,N_23586,N_23642);
nand U25065 (N_25065,N_23347,N_23947);
nand U25066 (N_25066,N_22553,N_21448);
or U25067 (N_25067,N_22825,N_22285);
nand U25068 (N_25068,N_23317,N_21295);
or U25069 (N_25069,N_23590,N_23344);
nand U25070 (N_25070,N_22012,N_21893);
and U25071 (N_25071,N_23434,N_22596);
and U25072 (N_25072,N_21665,N_22085);
or U25073 (N_25073,N_21599,N_22068);
or U25074 (N_25074,N_22065,N_22173);
nor U25075 (N_25075,N_23934,N_23065);
xor U25076 (N_25076,N_23714,N_21253);
or U25077 (N_25077,N_21041,N_23697);
nand U25078 (N_25078,N_23449,N_22911);
xor U25079 (N_25079,N_23328,N_23376);
nor U25080 (N_25080,N_21589,N_22524);
xor U25081 (N_25081,N_22289,N_22953);
xnor U25082 (N_25082,N_22372,N_23711);
xor U25083 (N_25083,N_23417,N_22281);
and U25084 (N_25084,N_22262,N_23289);
and U25085 (N_25085,N_23740,N_22151);
xnor U25086 (N_25086,N_22291,N_22839);
or U25087 (N_25087,N_22647,N_22211);
or U25088 (N_25088,N_22534,N_23902);
and U25089 (N_25089,N_22699,N_21576);
nor U25090 (N_25090,N_22091,N_23279);
nor U25091 (N_25091,N_22455,N_23794);
nor U25092 (N_25092,N_21826,N_23049);
or U25093 (N_25093,N_21976,N_21457);
and U25094 (N_25094,N_23911,N_22918);
or U25095 (N_25095,N_22273,N_22716);
nor U25096 (N_25096,N_21973,N_21968);
or U25097 (N_25097,N_21992,N_21222);
xor U25098 (N_25098,N_22205,N_22893);
xor U25099 (N_25099,N_21378,N_22234);
and U25100 (N_25100,N_21744,N_22946);
nand U25101 (N_25101,N_22755,N_22371);
or U25102 (N_25102,N_22488,N_23055);
nor U25103 (N_25103,N_22213,N_22966);
nand U25104 (N_25104,N_21030,N_21730);
nand U25105 (N_25105,N_22332,N_23429);
xnor U25106 (N_25106,N_21481,N_22888);
xnor U25107 (N_25107,N_21713,N_21910);
and U25108 (N_25108,N_23180,N_21564);
nand U25109 (N_25109,N_23224,N_21323);
or U25110 (N_25110,N_23286,N_23351);
xnor U25111 (N_25111,N_23167,N_22450);
or U25112 (N_25112,N_23640,N_23013);
xor U25113 (N_25113,N_22344,N_22977);
xor U25114 (N_25114,N_21009,N_23281);
or U25115 (N_25115,N_22853,N_22116);
and U25116 (N_25116,N_23183,N_21172);
or U25117 (N_25117,N_22849,N_23364);
nand U25118 (N_25118,N_23360,N_23646);
nor U25119 (N_25119,N_22723,N_22108);
xor U25120 (N_25120,N_22403,N_21334);
or U25121 (N_25121,N_21681,N_23682);
nor U25122 (N_25122,N_23043,N_22226);
xor U25123 (N_25123,N_22069,N_22079);
xnor U25124 (N_25124,N_22404,N_22675);
and U25125 (N_25125,N_21505,N_21266);
and U25126 (N_25126,N_22175,N_21991);
xor U25127 (N_25127,N_23753,N_21044);
and U25128 (N_25128,N_22505,N_22348);
or U25129 (N_25129,N_21524,N_21552);
or U25130 (N_25130,N_22531,N_22877);
and U25131 (N_25131,N_23670,N_23484);
nor U25132 (N_25132,N_21206,N_22666);
nor U25133 (N_25133,N_23889,N_22396);
xor U25134 (N_25134,N_22177,N_22857);
xor U25135 (N_25135,N_22542,N_23571);
or U25136 (N_25136,N_21153,N_23378);
or U25137 (N_25137,N_23601,N_22510);
nand U25138 (N_25138,N_22430,N_21071);
and U25139 (N_25139,N_22903,N_22702);
and U25140 (N_25140,N_22764,N_23707);
nor U25141 (N_25141,N_23208,N_22928);
and U25142 (N_25142,N_22366,N_21352);
or U25143 (N_25143,N_22936,N_23778);
nor U25144 (N_25144,N_23081,N_21139);
xnor U25145 (N_25145,N_21677,N_22361);
nand U25146 (N_25146,N_23410,N_21215);
or U25147 (N_25147,N_22561,N_22359);
nor U25148 (N_25148,N_23340,N_21930);
nand U25149 (N_25149,N_21126,N_22233);
or U25150 (N_25150,N_21473,N_21177);
or U25151 (N_25151,N_22431,N_22485);
nand U25152 (N_25152,N_22482,N_21367);
xor U25153 (N_25153,N_22195,N_22070);
and U25154 (N_25154,N_23015,N_23077);
xor U25155 (N_25155,N_23321,N_21329);
nor U25156 (N_25156,N_22885,N_23056);
or U25157 (N_25157,N_21627,N_21042);
and U25158 (N_25158,N_22623,N_21067);
nor U25159 (N_25159,N_23368,N_21771);
xor U25160 (N_25160,N_21403,N_21380);
nand U25161 (N_25161,N_22218,N_23029);
nor U25162 (N_25162,N_22830,N_23512);
xnor U25163 (N_25163,N_22794,N_23455);
and U25164 (N_25164,N_22651,N_21848);
nor U25165 (N_25165,N_22456,N_21345);
and U25166 (N_25166,N_22400,N_23856);
nand U25167 (N_25167,N_21395,N_23617);
and U25168 (N_25168,N_23557,N_22592);
or U25169 (N_25169,N_21614,N_23407);
nand U25170 (N_25170,N_23204,N_23287);
nor U25171 (N_25171,N_22609,N_23543);
xor U25172 (N_25172,N_22159,N_23163);
or U25173 (N_25173,N_23777,N_22604);
and U25174 (N_25174,N_23603,N_21234);
nand U25175 (N_25175,N_23651,N_21835);
nor U25176 (N_25176,N_22356,N_22053);
and U25177 (N_25177,N_21747,N_22414);
nor U25178 (N_25178,N_21236,N_22832);
xnor U25179 (N_25179,N_21591,N_23624);
nand U25180 (N_25180,N_22856,N_21112);
or U25181 (N_25181,N_22654,N_22377);
nand U25182 (N_25182,N_22425,N_21040);
and U25183 (N_25183,N_22688,N_21824);
and U25184 (N_25184,N_23415,N_21435);
xor U25185 (N_25185,N_22812,N_22667);
nor U25186 (N_25186,N_22519,N_21300);
nand U25187 (N_25187,N_22056,N_22843);
and U25188 (N_25188,N_23166,N_22865);
or U25189 (N_25189,N_23798,N_22880);
xor U25190 (N_25190,N_23604,N_22938);
xor U25191 (N_25191,N_21237,N_23217);
or U25192 (N_25192,N_22904,N_21209);
and U25193 (N_25193,N_22714,N_23379);
nand U25194 (N_25194,N_23996,N_22064);
xor U25195 (N_25195,N_22533,N_23148);
nor U25196 (N_25196,N_23223,N_21198);
and U25197 (N_25197,N_21129,N_23986);
and U25198 (N_25198,N_22294,N_22005);
nand U25199 (N_25199,N_21635,N_23377);
nand U25200 (N_25200,N_23194,N_22578);
or U25201 (N_25201,N_21945,N_22178);
nor U25202 (N_25202,N_23336,N_22477);
xnor U25203 (N_25203,N_21710,N_23251);
nor U25204 (N_25204,N_21478,N_21546);
or U25205 (N_25205,N_21133,N_23299);
and U25206 (N_25206,N_22058,N_23041);
nor U25207 (N_25207,N_23447,N_22744);
nor U25208 (N_25208,N_23523,N_23799);
xnor U25209 (N_25209,N_23588,N_22536);
or U25210 (N_25210,N_22858,N_22184);
nand U25211 (N_25211,N_21159,N_22754);
nand U25212 (N_25212,N_23044,N_21799);
nor U25213 (N_25213,N_22255,N_23678);
and U25214 (N_25214,N_23329,N_21849);
nand U25215 (N_25215,N_22981,N_21881);
nor U25216 (N_25216,N_21278,N_23017);
nor U25217 (N_25217,N_21915,N_21132);
nand U25218 (N_25218,N_23969,N_22662);
and U25219 (N_25219,N_21940,N_22509);
or U25220 (N_25220,N_22884,N_23500);
nor U25221 (N_25221,N_22748,N_23014);
xor U25222 (N_25222,N_21813,N_23991);
and U25223 (N_25223,N_21763,N_23949);
nor U25224 (N_25224,N_23414,N_23732);
xor U25225 (N_25225,N_21767,N_21097);
or U25226 (N_25226,N_21445,N_21572);
nor U25227 (N_25227,N_23452,N_22284);
nand U25228 (N_25228,N_22327,N_21788);
nand U25229 (N_25229,N_23662,N_23069);
nor U25230 (N_25230,N_22260,N_23213);
xor U25231 (N_25231,N_23128,N_22657);
or U25232 (N_25232,N_23683,N_23087);
xnor U25233 (N_25233,N_21424,N_21537);
or U25234 (N_25234,N_21636,N_21003);
xnor U25235 (N_25235,N_21078,N_23138);
xnor U25236 (N_25236,N_23318,N_21960);
nor U25237 (N_25237,N_22132,N_22296);
and U25238 (N_25238,N_22611,N_22760);
xor U25239 (N_25239,N_22117,N_22658);
xnor U25240 (N_25240,N_23791,N_21474);
nand U25241 (N_25241,N_23468,N_22632);
nor U25242 (N_25242,N_22631,N_21719);
nor U25243 (N_25243,N_21739,N_23333);
nand U25244 (N_25244,N_23582,N_21105);
nor U25245 (N_25245,N_23524,N_22555);
and U25246 (N_25246,N_23173,N_23192);
and U25247 (N_25247,N_23495,N_23462);
xnor U25248 (N_25248,N_23032,N_22597);
nand U25249 (N_25249,N_22872,N_22540);
xor U25250 (N_25250,N_21682,N_21987);
nor U25251 (N_25251,N_21137,N_22299);
xor U25252 (N_25252,N_22783,N_21107);
nand U25253 (N_25253,N_23227,N_21400);
xnor U25254 (N_25254,N_21717,N_22634);
nand U25255 (N_25255,N_22463,N_21840);
nor U25256 (N_25256,N_22871,N_22945);
and U25257 (N_25257,N_23456,N_21596);
or U25258 (N_25258,N_23970,N_22588);
xnor U25259 (N_25259,N_23558,N_23968);
nand U25260 (N_25260,N_23554,N_22137);
nand U25261 (N_25261,N_23229,N_21814);
and U25262 (N_25262,N_21472,N_23890);
and U25263 (N_25263,N_21273,N_23793);
nand U25264 (N_25264,N_22817,N_21401);
xor U25265 (N_25265,N_21507,N_23515);
xor U25266 (N_25266,N_23116,N_23324);
xnor U25267 (N_25267,N_22886,N_23814);
and U25268 (N_25268,N_21535,N_22630);
and U25269 (N_25269,N_21805,N_23549);
nor U25270 (N_25270,N_23998,N_22771);
or U25271 (N_25271,N_23837,N_23938);
xnor U25272 (N_25272,N_23858,N_21076);
nand U25273 (N_25273,N_21563,N_23773);
xor U25274 (N_25274,N_23467,N_23509);
xor U25275 (N_25275,N_23903,N_21740);
nor U25276 (N_25276,N_22302,N_21725);
xnor U25277 (N_25277,N_22677,N_22874);
and U25278 (N_25278,N_21226,N_22937);
nand U25279 (N_25279,N_23086,N_22614);
or U25280 (N_25280,N_23887,N_23396);
or U25281 (N_25281,N_21471,N_22350);
nand U25282 (N_25282,N_21142,N_23819);
xor U25283 (N_25283,N_23526,N_23231);
nand U25284 (N_25284,N_22998,N_23285);
nand U25285 (N_25285,N_22902,N_21659);
or U25286 (N_25286,N_21310,N_23611);
or U25287 (N_25287,N_22840,N_23809);
nand U25288 (N_25288,N_22111,N_22290);
or U25289 (N_25289,N_21954,N_21130);
nand U25290 (N_25290,N_23374,N_23294);
or U25291 (N_25291,N_21201,N_21208);
nand U25292 (N_25292,N_23062,N_21530);
and U25293 (N_25293,N_23265,N_23829);
or U25294 (N_25294,N_21303,N_21920);
nor U25295 (N_25295,N_21866,N_23510);
or U25296 (N_25296,N_22088,N_23952);
and U25297 (N_25297,N_23657,N_21565);
nand U25298 (N_25298,N_21686,N_22240);
or U25299 (N_25299,N_22827,N_22459);
xor U25300 (N_25300,N_22323,N_21101);
or U25301 (N_25301,N_22770,N_23776);
or U25302 (N_25302,N_21262,N_22570);
nor U25303 (N_25303,N_22250,N_23073);
xnor U25304 (N_25304,N_23211,N_23917);
and U25305 (N_25305,N_22443,N_23520);
nand U25306 (N_25306,N_22650,N_23222);
nand U25307 (N_25307,N_23119,N_21405);
nand U25308 (N_25308,N_22802,N_22909);
and U25309 (N_25309,N_21292,N_22917);
nor U25310 (N_25310,N_22671,N_23323);
and U25311 (N_25311,N_22204,N_22680);
or U25312 (N_25312,N_23079,N_23609);
nor U25313 (N_25313,N_23928,N_21606);
nand U25314 (N_25314,N_23290,N_21214);
and U25315 (N_25315,N_23463,N_23142);
nand U25316 (N_25316,N_21778,N_23698);
nand U25317 (N_25317,N_23046,N_21128);
or U25318 (N_25318,N_23892,N_21660);
nand U25319 (N_25319,N_22249,N_21611);
or U25320 (N_25320,N_21477,N_22330);
xnor U25321 (N_25321,N_23057,N_23627);
nand U25322 (N_25322,N_21319,N_21704);
and U25323 (N_25323,N_21254,N_22772);
or U25324 (N_25324,N_21604,N_22765);
or U25325 (N_25325,N_22674,N_23283);
nor U25326 (N_25326,N_21827,N_21521);
and U25327 (N_25327,N_23959,N_22267);
nor U25328 (N_25328,N_23757,N_21489);
or U25329 (N_25329,N_21746,N_21290);
xor U25330 (N_25330,N_22894,N_21202);
and U25331 (N_25331,N_22035,N_23602);
and U25332 (N_25332,N_21513,N_22678);
or U25333 (N_25333,N_23576,N_23910);
or U25334 (N_25334,N_23979,N_21929);
nor U25335 (N_25335,N_22055,N_23319);
nor U25336 (N_25336,N_23349,N_21617);
nand U25337 (N_25337,N_23570,N_23464);
xor U25338 (N_25338,N_21698,N_22171);
nand U25339 (N_25339,N_21885,N_21825);
and U25340 (N_25340,N_21487,N_21828);
or U25341 (N_25341,N_21687,N_21864);
and U25342 (N_25342,N_22778,N_23813);
or U25343 (N_25343,N_22846,N_22964);
and U25344 (N_25344,N_21124,N_22684);
xor U25345 (N_25345,N_22131,N_21070);
nand U25346 (N_25346,N_21276,N_23574);
and U25347 (N_25347,N_23004,N_22391);
nand U25348 (N_25348,N_22399,N_22544);
xnor U25349 (N_25349,N_21780,N_21762);
and U25350 (N_25350,N_23801,N_22319);
nor U25351 (N_25351,N_22826,N_23531);
nor U25352 (N_25352,N_21275,N_22491);
nand U25353 (N_25353,N_23562,N_23945);
or U25354 (N_25354,N_21597,N_23230);
xnor U25355 (N_25355,N_23144,N_22572);
nand U25356 (N_25356,N_23085,N_22201);
xor U25357 (N_25357,N_23628,N_22692);
or U25358 (N_25358,N_23894,N_23897);
or U25359 (N_25359,N_21318,N_21551);
nand U25360 (N_25360,N_21092,N_21851);
nor U25361 (N_25361,N_21182,N_22552);
nand U25362 (N_25362,N_22838,N_22265);
nand U25363 (N_25363,N_22792,N_22338);
or U25364 (N_25364,N_21025,N_23363);
nand U25365 (N_25365,N_22446,N_23024);
or U25366 (N_25366,N_21683,N_23916);
xor U25367 (N_25367,N_21752,N_22968);
nor U25368 (N_25368,N_21461,N_22188);
nor U25369 (N_25369,N_21578,N_23681);
nor U25370 (N_25370,N_21412,N_23381);
or U25371 (N_25371,N_23200,N_21638);
nor U25372 (N_25372,N_21018,N_22503);
and U25373 (N_25373,N_22245,N_21948);
xor U25374 (N_25374,N_21339,N_22793);
nor U25375 (N_25375,N_22000,N_21060);
and U25376 (N_25376,N_23450,N_22629);
and U25377 (N_25377,N_22636,N_22103);
and U25378 (N_25378,N_23665,N_21859);
nor U25379 (N_25379,N_22039,N_22780);
xnor U25380 (N_25380,N_23530,N_23908);
nor U25381 (N_25381,N_22527,N_22229);
nor U25382 (N_25382,N_21863,N_23309);
xor U25383 (N_25383,N_21120,N_22829);
and U25384 (N_25384,N_23580,N_22351);
nand U25385 (N_25385,N_21789,N_23796);
and U25386 (N_25386,N_23243,N_22462);
and U25387 (N_25387,N_22118,N_23070);
and U25388 (N_25388,N_21381,N_22149);
and U25389 (N_25389,N_22239,N_22571);
xor U25390 (N_25390,N_22992,N_21678);
or U25391 (N_25391,N_21304,N_21186);
nand U25392 (N_25392,N_23869,N_21270);
nand U25393 (N_25393,N_23944,N_21390);
nor U25394 (N_25394,N_23528,N_23828);
xor U25395 (N_25395,N_23560,N_23656);
or U25396 (N_25396,N_21096,N_21989);
xor U25397 (N_25397,N_22098,N_21024);
nor U25398 (N_25398,N_22320,N_22078);
and U25399 (N_25399,N_23688,N_22029);
nand U25400 (N_25400,N_21279,N_21409);
xnor U25401 (N_25401,N_21820,N_22698);
nor U25402 (N_25402,N_22980,N_23045);
nor U25403 (N_25403,N_23435,N_23130);
nand U25404 (N_25404,N_22288,N_21979);
nand U25405 (N_25405,N_21608,N_21451);
nor U25406 (N_25406,N_23335,N_22660);
nand U25407 (N_25407,N_22974,N_21895);
nand U25408 (N_25408,N_22586,N_22762);
or U25409 (N_25409,N_21315,N_21779);
nor U25410 (N_25410,N_23405,N_22014);
nor U25411 (N_25411,N_23544,N_23896);
nor U25412 (N_25412,N_21939,N_21243);
and U25413 (N_25413,N_21631,N_21213);
and U25414 (N_25414,N_23426,N_22374);
nor U25415 (N_25415,N_23252,N_21538);
and U25416 (N_25416,N_21721,N_22214);
or U25417 (N_25417,N_21411,N_23847);
nand U25418 (N_25418,N_21701,N_22432);
nor U25419 (N_25419,N_21528,N_22976);
or U25420 (N_25420,N_23716,N_22914);
or U25421 (N_25421,N_21860,N_23145);
xnor U25422 (N_25422,N_23724,N_23738);
and U25423 (N_25423,N_23039,N_23797);
and U25424 (N_25424,N_22152,N_23259);
or U25425 (N_25425,N_23780,N_23561);
and U25426 (N_25426,N_21759,N_23845);
xnor U25427 (N_25427,N_22419,N_21618);
or U25428 (N_25428,N_21005,N_23600);
nor U25429 (N_25429,N_23040,N_22752);
and U25430 (N_25430,N_22360,N_21533);
or U25431 (N_25431,N_21061,N_23136);
xnor U25432 (N_25432,N_22618,N_22225);
nand U25433 (N_25433,N_22326,N_22823);
or U25434 (N_25434,N_21841,N_23971);
nand U25435 (N_25435,N_22703,N_22833);
nand U25436 (N_25436,N_21265,N_22388);
nor U25437 (N_25437,N_21831,N_22855);
or U25438 (N_25438,N_23027,N_21520);
or U25439 (N_25439,N_22186,N_21366);
nand U25440 (N_25440,N_21059,N_23639);
or U25441 (N_25441,N_21557,N_23742);
xor U25442 (N_25442,N_22393,N_22345);
nor U25443 (N_25443,N_23293,N_21307);
nor U25444 (N_25444,N_22767,N_22283);
nor U25445 (N_25445,N_22097,N_21012);
or U25446 (N_25446,N_21047,N_23170);
or U25447 (N_25447,N_23356,N_22161);
nand U25448 (N_25448,N_21963,N_21579);
or U25449 (N_25449,N_21123,N_23465);
nor U25450 (N_25450,N_23614,N_23668);
or U25451 (N_25451,N_22738,N_23352);
or U25452 (N_25452,N_22820,N_22397);
xor U25453 (N_25453,N_23641,N_22148);
nor U25454 (N_25454,N_22612,N_23125);
xnor U25455 (N_25455,N_23734,N_22277);
xnor U25456 (N_25456,N_21179,N_23184);
and U25457 (N_25457,N_21644,N_22763);
and U25458 (N_25458,N_22433,N_22094);
xor U25459 (N_25459,N_22141,N_23203);
nor U25460 (N_25460,N_21936,N_23312);
nor U25461 (N_25461,N_21804,N_22709);
xnor U25462 (N_25462,N_21550,N_21085);
and U25463 (N_25463,N_22134,N_23960);
nor U25464 (N_25464,N_21134,N_22986);
and U25465 (N_25465,N_21204,N_23266);
and U25466 (N_25466,N_23755,N_21431);
nor U25467 (N_25467,N_23042,N_22003);
xnor U25468 (N_25468,N_22428,N_21511);
and U25469 (N_25469,N_22333,N_21916);
xor U25470 (N_25470,N_23505,N_22392);
and U25471 (N_25471,N_21420,N_23518);
or U25472 (N_25472,N_23935,N_23775);
nor U25473 (N_25473,N_21015,N_22750);
nor U25474 (N_25474,N_23635,N_22773);
xor U25475 (N_25475,N_22153,N_21282);
and U25476 (N_25476,N_22962,N_22021);
and U25477 (N_25477,N_22728,N_22022);
or U25478 (N_25478,N_23413,N_21833);
nand U25479 (N_25479,N_22125,N_21844);
nand U25480 (N_25480,N_21765,N_21663);
and U25481 (N_25481,N_21853,N_23621);
and U25482 (N_25482,N_22991,N_22395);
or U25483 (N_25483,N_23384,N_23932);
nor U25484 (N_25484,N_21083,N_23536);
nor U25485 (N_25485,N_22227,N_23051);
and U25486 (N_25486,N_21357,N_22487);
nand U25487 (N_25487,N_21294,N_22497);
and U25488 (N_25488,N_23629,N_23620);
or U25489 (N_25489,N_22492,N_23048);
or U25490 (N_25490,N_23064,N_21459);
xnor U25491 (N_25491,N_21200,N_22220);
xnor U25492 (N_25492,N_23245,N_21406);
xnor U25493 (N_25493,N_21416,N_21439);
nand U25494 (N_25494,N_21374,N_23728);
xnor U25495 (N_25495,N_21056,N_21466);
or U25496 (N_25496,N_23241,N_23943);
nor U25497 (N_25497,N_22993,N_23900);
and U25498 (N_25498,N_23146,N_23260);
xnor U25499 (N_25499,N_23516,N_22090);
nor U25500 (N_25500,N_23106,N_22914);
and U25501 (N_25501,N_22127,N_22440);
and U25502 (N_25502,N_23335,N_23478);
or U25503 (N_25503,N_21686,N_23956);
or U25504 (N_25504,N_23222,N_21775);
xor U25505 (N_25505,N_22995,N_22454);
nor U25506 (N_25506,N_22328,N_21965);
xor U25507 (N_25507,N_23484,N_23382);
and U25508 (N_25508,N_21455,N_23465);
and U25509 (N_25509,N_21032,N_22676);
or U25510 (N_25510,N_22268,N_21062);
xnor U25511 (N_25511,N_22256,N_23914);
xor U25512 (N_25512,N_23025,N_22468);
nand U25513 (N_25513,N_21173,N_23169);
xor U25514 (N_25514,N_23483,N_22768);
and U25515 (N_25515,N_22580,N_23729);
xor U25516 (N_25516,N_21078,N_23828);
nor U25517 (N_25517,N_22200,N_23310);
nor U25518 (N_25518,N_22239,N_22241);
and U25519 (N_25519,N_22331,N_21789);
xor U25520 (N_25520,N_21166,N_22188);
and U25521 (N_25521,N_21252,N_22605);
nor U25522 (N_25522,N_22135,N_23977);
or U25523 (N_25523,N_22557,N_23875);
or U25524 (N_25524,N_21949,N_21374);
or U25525 (N_25525,N_22020,N_21088);
nand U25526 (N_25526,N_21928,N_23135);
xnor U25527 (N_25527,N_21038,N_23769);
xnor U25528 (N_25528,N_21535,N_21404);
xor U25529 (N_25529,N_22923,N_22164);
xor U25530 (N_25530,N_22747,N_23529);
or U25531 (N_25531,N_23568,N_23878);
or U25532 (N_25532,N_22923,N_23929);
and U25533 (N_25533,N_23444,N_21229);
and U25534 (N_25534,N_22505,N_23842);
xnor U25535 (N_25535,N_22905,N_23358);
xor U25536 (N_25536,N_23582,N_22966);
nor U25537 (N_25537,N_22676,N_21584);
nor U25538 (N_25538,N_23228,N_22680);
or U25539 (N_25539,N_21266,N_22415);
xor U25540 (N_25540,N_22307,N_23683);
nand U25541 (N_25541,N_21410,N_21523);
xor U25542 (N_25542,N_23655,N_21808);
xor U25543 (N_25543,N_21556,N_23055);
nor U25544 (N_25544,N_21922,N_22357);
nor U25545 (N_25545,N_23251,N_22272);
xnor U25546 (N_25546,N_23172,N_21570);
nand U25547 (N_25547,N_23578,N_22509);
xnor U25548 (N_25548,N_22037,N_23742);
xnor U25549 (N_25549,N_21186,N_22512);
or U25550 (N_25550,N_21581,N_23984);
or U25551 (N_25551,N_21338,N_22333);
nand U25552 (N_25552,N_22007,N_21522);
nand U25553 (N_25553,N_21891,N_23208);
nand U25554 (N_25554,N_21447,N_21571);
xnor U25555 (N_25555,N_22256,N_21114);
nor U25556 (N_25556,N_21142,N_23315);
or U25557 (N_25557,N_21046,N_23016);
or U25558 (N_25558,N_21306,N_23384);
nor U25559 (N_25559,N_21923,N_22633);
nor U25560 (N_25560,N_22009,N_23522);
and U25561 (N_25561,N_22400,N_21145);
xor U25562 (N_25562,N_21625,N_23177);
xnor U25563 (N_25563,N_21432,N_21123);
xor U25564 (N_25564,N_23848,N_21586);
and U25565 (N_25565,N_23200,N_22361);
and U25566 (N_25566,N_22604,N_21998);
and U25567 (N_25567,N_23531,N_23693);
nand U25568 (N_25568,N_21527,N_22998);
nor U25569 (N_25569,N_22790,N_23665);
nand U25570 (N_25570,N_21271,N_23419);
and U25571 (N_25571,N_23593,N_22910);
xor U25572 (N_25572,N_22725,N_22206);
nor U25573 (N_25573,N_23316,N_22547);
nand U25574 (N_25574,N_23233,N_21358);
or U25575 (N_25575,N_21846,N_23622);
and U25576 (N_25576,N_22883,N_22404);
and U25577 (N_25577,N_21233,N_22451);
xor U25578 (N_25578,N_22919,N_21790);
xnor U25579 (N_25579,N_21260,N_22357);
nand U25580 (N_25580,N_21750,N_23950);
nor U25581 (N_25581,N_23370,N_23385);
nand U25582 (N_25582,N_21246,N_21238);
and U25583 (N_25583,N_22126,N_21896);
nand U25584 (N_25584,N_22371,N_23819);
nor U25585 (N_25585,N_21307,N_22080);
and U25586 (N_25586,N_21041,N_21511);
and U25587 (N_25587,N_23275,N_21615);
or U25588 (N_25588,N_23674,N_23926);
or U25589 (N_25589,N_21752,N_21821);
nand U25590 (N_25590,N_22415,N_22334);
or U25591 (N_25591,N_21574,N_21599);
xor U25592 (N_25592,N_22776,N_22764);
xnor U25593 (N_25593,N_21233,N_22389);
nor U25594 (N_25594,N_23611,N_21778);
nand U25595 (N_25595,N_21614,N_21456);
xnor U25596 (N_25596,N_21496,N_21300);
and U25597 (N_25597,N_23357,N_21984);
xnor U25598 (N_25598,N_22318,N_23820);
nor U25599 (N_25599,N_23678,N_21797);
and U25600 (N_25600,N_21019,N_23065);
or U25601 (N_25601,N_22769,N_22440);
xor U25602 (N_25602,N_23559,N_23348);
and U25603 (N_25603,N_23575,N_21003);
xor U25604 (N_25604,N_22485,N_23985);
nand U25605 (N_25605,N_22791,N_21689);
or U25606 (N_25606,N_21258,N_22577);
nand U25607 (N_25607,N_21252,N_23301);
nor U25608 (N_25608,N_21571,N_21039);
and U25609 (N_25609,N_22150,N_23216);
xnor U25610 (N_25610,N_23408,N_23988);
nand U25611 (N_25611,N_22705,N_23430);
or U25612 (N_25612,N_23788,N_21567);
or U25613 (N_25613,N_22005,N_21804);
xnor U25614 (N_25614,N_22172,N_21950);
and U25615 (N_25615,N_21729,N_23494);
nand U25616 (N_25616,N_23284,N_21803);
xnor U25617 (N_25617,N_23952,N_22948);
nand U25618 (N_25618,N_21220,N_22726);
nor U25619 (N_25619,N_21570,N_23543);
nand U25620 (N_25620,N_23539,N_22419);
nor U25621 (N_25621,N_21712,N_22573);
nor U25622 (N_25622,N_22016,N_21472);
xor U25623 (N_25623,N_22855,N_23433);
nand U25624 (N_25624,N_23373,N_22790);
xnor U25625 (N_25625,N_21728,N_23869);
nand U25626 (N_25626,N_21331,N_22526);
or U25627 (N_25627,N_23508,N_23339);
and U25628 (N_25628,N_21477,N_21715);
xnor U25629 (N_25629,N_22232,N_21833);
and U25630 (N_25630,N_23199,N_21745);
or U25631 (N_25631,N_22079,N_22900);
and U25632 (N_25632,N_21291,N_23404);
xnor U25633 (N_25633,N_21380,N_21910);
and U25634 (N_25634,N_21328,N_21999);
xor U25635 (N_25635,N_22475,N_23214);
xnor U25636 (N_25636,N_23439,N_23485);
xor U25637 (N_25637,N_21370,N_22965);
or U25638 (N_25638,N_21968,N_23281);
xor U25639 (N_25639,N_22097,N_23153);
xor U25640 (N_25640,N_23185,N_22093);
xor U25641 (N_25641,N_21106,N_21058);
xor U25642 (N_25642,N_22121,N_22668);
nor U25643 (N_25643,N_21714,N_22640);
xnor U25644 (N_25644,N_21538,N_22922);
nand U25645 (N_25645,N_23224,N_22656);
xor U25646 (N_25646,N_22961,N_23649);
nor U25647 (N_25647,N_23980,N_22335);
nand U25648 (N_25648,N_21485,N_23613);
or U25649 (N_25649,N_23318,N_23301);
xor U25650 (N_25650,N_21762,N_23089);
and U25651 (N_25651,N_21115,N_22816);
nand U25652 (N_25652,N_23773,N_22314);
and U25653 (N_25653,N_21912,N_23308);
or U25654 (N_25654,N_21339,N_22697);
xor U25655 (N_25655,N_22644,N_22708);
nor U25656 (N_25656,N_23002,N_22638);
nor U25657 (N_25657,N_21689,N_22044);
nor U25658 (N_25658,N_23672,N_22864);
and U25659 (N_25659,N_23767,N_23827);
nand U25660 (N_25660,N_21726,N_22478);
xor U25661 (N_25661,N_21640,N_22951);
nor U25662 (N_25662,N_21153,N_23645);
nand U25663 (N_25663,N_21026,N_22339);
xnor U25664 (N_25664,N_21529,N_21361);
or U25665 (N_25665,N_21258,N_21781);
or U25666 (N_25666,N_21669,N_23001);
and U25667 (N_25667,N_21877,N_21599);
and U25668 (N_25668,N_21299,N_21086);
or U25669 (N_25669,N_21920,N_23728);
nor U25670 (N_25670,N_21673,N_22549);
and U25671 (N_25671,N_21222,N_22565);
nand U25672 (N_25672,N_21180,N_21021);
xnor U25673 (N_25673,N_22613,N_22519);
xnor U25674 (N_25674,N_22877,N_22079);
and U25675 (N_25675,N_21624,N_22794);
nand U25676 (N_25676,N_21918,N_23257);
xnor U25677 (N_25677,N_23738,N_23685);
and U25678 (N_25678,N_21636,N_22195);
nor U25679 (N_25679,N_23844,N_21984);
or U25680 (N_25680,N_22402,N_21980);
or U25681 (N_25681,N_21242,N_21411);
nand U25682 (N_25682,N_23582,N_21474);
or U25683 (N_25683,N_23064,N_23287);
and U25684 (N_25684,N_23150,N_22228);
xor U25685 (N_25685,N_23820,N_22877);
nand U25686 (N_25686,N_23253,N_23637);
xnor U25687 (N_25687,N_21004,N_22439);
or U25688 (N_25688,N_23637,N_21507);
and U25689 (N_25689,N_22438,N_23350);
or U25690 (N_25690,N_23856,N_23009);
nand U25691 (N_25691,N_21802,N_23174);
or U25692 (N_25692,N_23728,N_23694);
xor U25693 (N_25693,N_23525,N_21798);
or U25694 (N_25694,N_23189,N_21079);
or U25695 (N_25695,N_21231,N_22508);
and U25696 (N_25696,N_22164,N_22254);
nor U25697 (N_25697,N_21266,N_21310);
or U25698 (N_25698,N_21997,N_23523);
or U25699 (N_25699,N_21085,N_22740);
and U25700 (N_25700,N_21482,N_21509);
nand U25701 (N_25701,N_22133,N_21846);
nand U25702 (N_25702,N_22492,N_22909);
and U25703 (N_25703,N_22302,N_21619);
xnor U25704 (N_25704,N_23885,N_23849);
nor U25705 (N_25705,N_23862,N_23464);
nand U25706 (N_25706,N_23409,N_23579);
or U25707 (N_25707,N_21068,N_23563);
nand U25708 (N_25708,N_21527,N_23992);
nand U25709 (N_25709,N_21415,N_23294);
nor U25710 (N_25710,N_21894,N_21231);
nand U25711 (N_25711,N_22862,N_23627);
nor U25712 (N_25712,N_22469,N_21350);
and U25713 (N_25713,N_22398,N_23956);
or U25714 (N_25714,N_23591,N_22028);
and U25715 (N_25715,N_23868,N_22906);
and U25716 (N_25716,N_22480,N_22785);
and U25717 (N_25717,N_21713,N_23068);
xnor U25718 (N_25718,N_21596,N_23131);
and U25719 (N_25719,N_23081,N_23618);
nor U25720 (N_25720,N_22778,N_22531);
xnor U25721 (N_25721,N_23937,N_23905);
or U25722 (N_25722,N_23666,N_21500);
nor U25723 (N_25723,N_21270,N_21059);
or U25724 (N_25724,N_22095,N_22529);
or U25725 (N_25725,N_22201,N_23199);
nor U25726 (N_25726,N_23657,N_23602);
nand U25727 (N_25727,N_23937,N_22929);
nor U25728 (N_25728,N_21411,N_23708);
or U25729 (N_25729,N_21111,N_22006);
nand U25730 (N_25730,N_23882,N_22817);
nor U25731 (N_25731,N_23011,N_23229);
nand U25732 (N_25732,N_21379,N_22838);
and U25733 (N_25733,N_22703,N_21085);
or U25734 (N_25734,N_22552,N_22077);
nor U25735 (N_25735,N_23806,N_22356);
and U25736 (N_25736,N_21059,N_23562);
xor U25737 (N_25737,N_21026,N_21215);
nor U25738 (N_25738,N_21354,N_23091);
nor U25739 (N_25739,N_23467,N_23892);
or U25740 (N_25740,N_23478,N_22384);
or U25741 (N_25741,N_22217,N_22472);
nor U25742 (N_25742,N_22714,N_22141);
nand U25743 (N_25743,N_23569,N_22510);
and U25744 (N_25744,N_21164,N_22544);
and U25745 (N_25745,N_23610,N_23213);
and U25746 (N_25746,N_22829,N_23079);
and U25747 (N_25747,N_23844,N_22497);
nor U25748 (N_25748,N_22052,N_21392);
or U25749 (N_25749,N_22081,N_23985);
or U25750 (N_25750,N_23658,N_22268);
xnor U25751 (N_25751,N_22589,N_22744);
and U25752 (N_25752,N_21053,N_22667);
nand U25753 (N_25753,N_23921,N_23993);
or U25754 (N_25754,N_22902,N_22091);
and U25755 (N_25755,N_23052,N_23481);
nor U25756 (N_25756,N_22623,N_22944);
nand U25757 (N_25757,N_23403,N_21679);
and U25758 (N_25758,N_23246,N_23924);
and U25759 (N_25759,N_22184,N_23059);
nor U25760 (N_25760,N_21777,N_22057);
nor U25761 (N_25761,N_22143,N_21717);
nand U25762 (N_25762,N_22073,N_23722);
nand U25763 (N_25763,N_23490,N_23908);
and U25764 (N_25764,N_23856,N_21913);
xnor U25765 (N_25765,N_21939,N_23059);
nand U25766 (N_25766,N_21207,N_22169);
nor U25767 (N_25767,N_22132,N_21123);
and U25768 (N_25768,N_21595,N_21770);
xnor U25769 (N_25769,N_23377,N_22711);
and U25770 (N_25770,N_22643,N_22229);
nand U25771 (N_25771,N_23226,N_22747);
and U25772 (N_25772,N_21140,N_21025);
nor U25773 (N_25773,N_22168,N_23270);
nor U25774 (N_25774,N_21057,N_23466);
or U25775 (N_25775,N_21663,N_21108);
xor U25776 (N_25776,N_21769,N_22012);
nand U25777 (N_25777,N_21870,N_23072);
or U25778 (N_25778,N_21823,N_22217);
and U25779 (N_25779,N_23388,N_21354);
nand U25780 (N_25780,N_23118,N_22718);
or U25781 (N_25781,N_21137,N_22559);
xor U25782 (N_25782,N_21342,N_22334);
nand U25783 (N_25783,N_21643,N_23426);
nor U25784 (N_25784,N_22410,N_21595);
xnor U25785 (N_25785,N_22774,N_23742);
and U25786 (N_25786,N_23426,N_23127);
or U25787 (N_25787,N_21305,N_22015);
and U25788 (N_25788,N_22208,N_22394);
or U25789 (N_25789,N_22637,N_23114);
xor U25790 (N_25790,N_23246,N_21518);
nand U25791 (N_25791,N_22266,N_22901);
nor U25792 (N_25792,N_21851,N_22573);
nor U25793 (N_25793,N_23185,N_22430);
and U25794 (N_25794,N_21090,N_22352);
and U25795 (N_25795,N_23474,N_22860);
and U25796 (N_25796,N_21429,N_21681);
and U25797 (N_25797,N_21278,N_21641);
nand U25798 (N_25798,N_21672,N_22796);
nor U25799 (N_25799,N_23093,N_22337);
nor U25800 (N_25800,N_21155,N_22392);
nand U25801 (N_25801,N_23805,N_22718);
xnor U25802 (N_25802,N_22331,N_21492);
xnor U25803 (N_25803,N_22001,N_22354);
and U25804 (N_25804,N_21615,N_21090);
xor U25805 (N_25805,N_22214,N_21535);
nor U25806 (N_25806,N_21680,N_23862);
and U25807 (N_25807,N_21874,N_23262);
xnor U25808 (N_25808,N_21636,N_21928);
nand U25809 (N_25809,N_23810,N_21927);
nand U25810 (N_25810,N_23623,N_22011);
xnor U25811 (N_25811,N_22220,N_23642);
xor U25812 (N_25812,N_21061,N_22889);
nand U25813 (N_25813,N_21754,N_22828);
and U25814 (N_25814,N_23083,N_22136);
or U25815 (N_25815,N_21452,N_21436);
nor U25816 (N_25816,N_21835,N_23078);
nand U25817 (N_25817,N_23830,N_23342);
and U25818 (N_25818,N_22724,N_23036);
and U25819 (N_25819,N_23494,N_22842);
and U25820 (N_25820,N_23175,N_23082);
nor U25821 (N_25821,N_21628,N_22904);
nor U25822 (N_25822,N_21489,N_22958);
nand U25823 (N_25823,N_21403,N_21535);
nor U25824 (N_25824,N_21116,N_22602);
or U25825 (N_25825,N_22997,N_22946);
nor U25826 (N_25826,N_23512,N_21048);
nor U25827 (N_25827,N_22740,N_22301);
or U25828 (N_25828,N_23598,N_22259);
and U25829 (N_25829,N_23960,N_23580);
and U25830 (N_25830,N_23242,N_23323);
nor U25831 (N_25831,N_23657,N_23805);
xnor U25832 (N_25832,N_21266,N_22661);
and U25833 (N_25833,N_22177,N_22417);
nand U25834 (N_25834,N_21149,N_22856);
or U25835 (N_25835,N_23452,N_21519);
and U25836 (N_25836,N_23774,N_23693);
or U25837 (N_25837,N_22427,N_23124);
and U25838 (N_25838,N_23873,N_21208);
nor U25839 (N_25839,N_23943,N_22796);
nor U25840 (N_25840,N_22470,N_23417);
nand U25841 (N_25841,N_22431,N_23240);
or U25842 (N_25842,N_23543,N_21406);
xor U25843 (N_25843,N_22403,N_21791);
xnor U25844 (N_25844,N_23001,N_21947);
nor U25845 (N_25845,N_22969,N_23461);
nand U25846 (N_25846,N_23438,N_23774);
or U25847 (N_25847,N_23005,N_22157);
or U25848 (N_25848,N_22533,N_21413);
and U25849 (N_25849,N_23898,N_22040);
nand U25850 (N_25850,N_22583,N_23531);
nand U25851 (N_25851,N_22687,N_23547);
nor U25852 (N_25852,N_23068,N_23602);
or U25853 (N_25853,N_23737,N_23989);
or U25854 (N_25854,N_21437,N_22853);
and U25855 (N_25855,N_22516,N_21665);
and U25856 (N_25856,N_23559,N_23802);
or U25857 (N_25857,N_23432,N_21037);
and U25858 (N_25858,N_21783,N_22060);
or U25859 (N_25859,N_23892,N_21530);
nand U25860 (N_25860,N_22726,N_23330);
and U25861 (N_25861,N_22933,N_23203);
and U25862 (N_25862,N_21386,N_21545);
nor U25863 (N_25863,N_23789,N_22045);
nand U25864 (N_25864,N_21288,N_21021);
and U25865 (N_25865,N_21334,N_22964);
nand U25866 (N_25866,N_21015,N_23516);
nor U25867 (N_25867,N_23890,N_22410);
and U25868 (N_25868,N_21592,N_23433);
and U25869 (N_25869,N_21278,N_22239);
nand U25870 (N_25870,N_23869,N_22925);
nor U25871 (N_25871,N_23074,N_22570);
nand U25872 (N_25872,N_23884,N_23386);
nand U25873 (N_25873,N_23535,N_23628);
and U25874 (N_25874,N_21157,N_21852);
nand U25875 (N_25875,N_23280,N_22380);
nor U25876 (N_25876,N_23703,N_21308);
and U25877 (N_25877,N_21550,N_21680);
xor U25878 (N_25878,N_21487,N_22170);
and U25879 (N_25879,N_22253,N_23359);
xnor U25880 (N_25880,N_23724,N_23974);
and U25881 (N_25881,N_21460,N_23544);
nor U25882 (N_25882,N_23322,N_22152);
or U25883 (N_25883,N_23368,N_23356);
and U25884 (N_25884,N_23857,N_21072);
nor U25885 (N_25885,N_22831,N_21284);
nor U25886 (N_25886,N_22534,N_23817);
xor U25887 (N_25887,N_21634,N_22398);
nor U25888 (N_25888,N_21934,N_21900);
xor U25889 (N_25889,N_21602,N_21235);
and U25890 (N_25890,N_22863,N_22227);
or U25891 (N_25891,N_21352,N_23964);
nand U25892 (N_25892,N_22191,N_23739);
and U25893 (N_25893,N_22170,N_23134);
and U25894 (N_25894,N_22487,N_22253);
nor U25895 (N_25895,N_21735,N_22517);
xnor U25896 (N_25896,N_22366,N_23924);
and U25897 (N_25897,N_23962,N_21419);
nor U25898 (N_25898,N_22793,N_23709);
xor U25899 (N_25899,N_23855,N_21602);
xor U25900 (N_25900,N_22110,N_22634);
nand U25901 (N_25901,N_22081,N_21232);
nor U25902 (N_25902,N_22493,N_21698);
nor U25903 (N_25903,N_21312,N_23522);
or U25904 (N_25904,N_22743,N_21197);
nand U25905 (N_25905,N_23845,N_21244);
and U25906 (N_25906,N_22724,N_23100);
and U25907 (N_25907,N_21213,N_21556);
nand U25908 (N_25908,N_23465,N_23038);
or U25909 (N_25909,N_21736,N_23913);
xnor U25910 (N_25910,N_21500,N_23009);
nor U25911 (N_25911,N_21816,N_23603);
xnor U25912 (N_25912,N_23066,N_21852);
xor U25913 (N_25913,N_22216,N_22951);
nand U25914 (N_25914,N_21072,N_22906);
nand U25915 (N_25915,N_22014,N_21848);
nor U25916 (N_25916,N_21701,N_21824);
xor U25917 (N_25917,N_21969,N_22821);
xnor U25918 (N_25918,N_22623,N_23229);
nor U25919 (N_25919,N_23522,N_21413);
or U25920 (N_25920,N_23538,N_23285);
nor U25921 (N_25921,N_23290,N_21638);
or U25922 (N_25922,N_21867,N_21007);
xor U25923 (N_25923,N_23353,N_21985);
and U25924 (N_25924,N_22040,N_23361);
nor U25925 (N_25925,N_22050,N_23854);
and U25926 (N_25926,N_22505,N_23334);
xnor U25927 (N_25927,N_21945,N_21668);
nand U25928 (N_25928,N_21190,N_23876);
xor U25929 (N_25929,N_22277,N_22996);
or U25930 (N_25930,N_23355,N_21272);
nor U25931 (N_25931,N_23512,N_22274);
and U25932 (N_25932,N_22662,N_21069);
nand U25933 (N_25933,N_22745,N_22253);
xnor U25934 (N_25934,N_22858,N_22222);
and U25935 (N_25935,N_22086,N_22052);
and U25936 (N_25936,N_23141,N_22753);
nor U25937 (N_25937,N_23323,N_21079);
and U25938 (N_25938,N_22876,N_21335);
and U25939 (N_25939,N_23018,N_23077);
and U25940 (N_25940,N_22801,N_22492);
nand U25941 (N_25941,N_22873,N_22075);
and U25942 (N_25942,N_23238,N_22440);
xnor U25943 (N_25943,N_21475,N_22635);
xor U25944 (N_25944,N_22240,N_23369);
xor U25945 (N_25945,N_21935,N_23953);
nand U25946 (N_25946,N_21160,N_21319);
xor U25947 (N_25947,N_21478,N_22636);
or U25948 (N_25948,N_23403,N_22405);
or U25949 (N_25949,N_22408,N_23844);
nor U25950 (N_25950,N_21355,N_23309);
nand U25951 (N_25951,N_23024,N_21117);
xnor U25952 (N_25952,N_23462,N_23237);
nand U25953 (N_25953,N_23700,N_22308);
nand U25954 (N_25954,N_21588,N_21428);
nand U25955 (N_25955,N_23676,N_21339);
nand U25956 (N_25956,N_23692,N_22108);
or U25957 (N_25957,N_23925,N_23901);
nand U25958 (N_25958,N_23966,N_21701);
nor U25959 (N_25959,N_22348,N_21287);
xnor U25960 (N_25960,N_22562,N_23025);
or U25961 (N_25961,N_22274,N_22746);
nand U25962 (N_25962,N_22045,N_22581);
or U25963 (N_25963,N_23827,N_22137);
and U25964 (N_25964,N_21305,N_21666);
nand U25965 (N_25965,N_21368,N_22197);
nand U25966 (N_25966,N_23431,N_21434);
nand U25967 (N_25967,N_21949,N_23147);
nand U25968 (N_25968,N_21765,N_22648);
and U25969 (N_25969,N_23597,N_21338);
nor U25970 (N_25970,N_22417,N_21721);
nor U25971 (N_25971,N_23865,N_21170);
nor U25972 (N_25972,N_22030,N_23297);
xor U25973 (N_25973,N_22181,N_22203);
nor U25974 (N_25974,N_21334,N_21775);
and U25975 (N_25975,N_22706,N_22105);
xnor U25976 (N_25976,N_21921,N_22433);
and U25977 (N_25977,N_22017,N_22866);
nand U25978 (N_25978,N_21304,N_22572);
or U25979 (N_25979,N_23560,N_23404);
and U25980 (N_25980,N_21942,N_23889);
or U25981 (N_25981,N_21753,N_22702);
nand U25982 (N_25982,N_23838,N_22244);
or U25983 (N_25983,N_22967,N_22005);
or U25984 (N_25984,N_23512,N_22204);
xnor U25985 (N_25985,N_21308,N_23922);
and U25986 (N_25986,N_23209,N_22215);
nand U25987 (N_25987,N_21061,N_21888);
nor U25988 (N_25988,N_22629,N_22603);
nor U25989 (N_25989,N_22802,N_23904);
nor U25990 (N_25990,N_21813,N_21148);
xor U25991 (N_25991,N_21585,N_23015);
xor U25992 (N_25992,N_23729,N_23454);
nor U25993 (N_25993,N_22703,N_23126);
or U25994 (N_25994,N_23642,N_22775);
nand U25995 (N_25995,N_21608,N_22711);
xor U25996 (N_25996,N_21993,N_23035);
or U25997 (N_25997,N_23611,N_21927);
or U25998 (N_25998,N_23454,N_22810);
nand U25999 (N_25999,N_21750,N_21621);
and U26000 (N_26000,N_23347,N_22088);
or U26001 (N_26001,N_23840,N_21235);
and U26002 (N_26002,N_22138,N_21362);
and U26003 (N_26003,N_23095,N_21413);
nand U26004 (N_26004,N_23904,N_21314);
xnor U26005 (N_26005,N_21332,N_21682);
nand U26006 (N_26006,N_22401,N_21943);
and U26007 (N_26007,N_22644,N_22914);
nand U26008 (N_26008,N_21754,N_23205);
xnor U26009 (N_26009,N_22449,N_21249);
xor U26010 (N_26010,N_23032,N_21187);
xor U26011 (N_26011,N_22299,N_23831);
nor U26012 (N_26012,N_23133,N_21757);
and U26013 (N_26013,N_21339,N_22124);
or U26014 (N_26014,N_23202,N_21602);
nor U26015 (N_26015,N_23831,N_23762);
nor U26016 (N_26016,N_22714,N_22284);
nand U26017 (N_26017,N_21582,N_21432);
nand U26018 (N_26018,N_21883,N_22482);
or U26019 (N_26019,N_22437,N_21827);
xor U26020 (N_26020,N_23472,N_21320);
and U26021 (N_26021,N_21514,N_23984);
and U26022 (N_26022,N_22112,N_22219);
nand U26023 (N_26023,N_23626,N_23750);
nor U26024 (N_26024,N_22576,N_22101);
nand U26025 (N_26025,N_21382,N_21936);
or U26026 (N_26026,N_23945,N_22507);
xnor U26027 (N_26027,N_23858,N_23348);
xnor U26028 (N_26028,N_22820,N_23113);
xnor U26029 (N_26029,N_22051,N_22820);
nor U26030 (N_26030,N_21038,N_21109);
nand U26031 (N_26031,N_21127,N_23622);
or U26032 (N_26032,N_21108,N_23707);
nor U26033 (N_26033,N_21972,N_21648);
and U26034 (N_26034,N_21633,N_21829);
and U26035 (N_26035,N_23423,N_22924);
and U26036 (N_26036,N_23877,N_23752);
nor U26037 (N_26037,N_22803,N_23394);
nand U26038 (N_26038,N_23131,N_21124);
xor U26039 (N_26039,N_23169,N_22093);
nor U26040 (N_26040,N_21063,N_22002);
or U26041 (N_26041,N_23883,N_21631);
and U26042 (N_26042,N_22399,N_23752);
nor U26043 (N_26043,N_21049,N_22362);
and U26044 (N_26044,N_21360,N_21917);
or U26045 (N_26045,N_23534,N_23081);
xnor U26046 (N_26046,N_22849,N_21845);
or U26047 (N_26047,N_23972,N_21338);
and U26048 (N_26048,N_22629,N_23035);
nand U26049 (N_26049,N_21740,N_22195);
and U26050 (N_26050,N_22438,N_21531);
nor U26051 (N_26051,N_23444,N_21765);
xor U26052 (N_26052,N_23050,N_23081);
and U26053 (N_26053,N_23769,N_22726);
nand U26054 (N_26054,N_22833,N_22301);
xor U26055 (N_26055,N_22615,N_23127);
or U26056 (N_26056,N_22056,N_21602);
or U26057 (N_26057,N_23067,N_23163);
nor U26058 (N_26058,N_21461,N_23249);
xor U26059 (N_26059,N_21550,N_21157);
or U26060 (N_26060,N_23996,N_23060);
and U26061 (N_26061,N_21984,N_23184);
nand U26062 (N_26062,N_21596,N_21048);
nand U26063 (N_26063,N_23921,N_21348);
and U26064 (N_26064,N_23695,N_22175);
nor U26065 (N_26065,N_23522,N_22044);
nor U26066 (N_26066,N_23993,N_23532);
nand U26067 (N_26067,N_23931,N_22588);
nand U26068 (N_26068,N_21347,N_21448);
or U26069 (N_26069,N_22559,N_21532);
xnor U26070 (N_26070,N_23695,N_23733);
or U26071 (N_26071,N_21831,N_23423);
nor U26072 (N_26072,N_23396,N_22103);
or U26073 (N_26073,N_23176,N_22236);
nand U26074 (N_26074,N_23239,N_21553);
nor U26075 (N_26075,N_21792,N_21727);
xnor U26076 (N_26076,N_22427,N_22134);
nand U26077 (N_26077,N_21200,N_23674);
nor U26078 (N_26078,N_23585,N_21250);
and U26079 (N_26079,N_21681,N_21086);
and U26080 (N_26080,N_22809,N_21414);
xnor U26081 (N_26081,N_21339,N_22719);
and U26082 (N_26082,N_21267,N_23044);
nand U26083 (N_26083,N_23286,N_21162);
nor U26084 (N_26084,N_23358,N_21378);
nor U26085 (N_26085,N_23041,N_23196);
xnor U26086 (N_26086,N_23130,N_21425);
xor U26087 (N_26087,N_23038,N_22440);
nand U26088 (N_26088,N_21399,N_21164);
or U26089 (N_26089,N_22082,N_22392);
nor U26090 (N_26090,N_23879,N_21411);
and U26091 (N_26091,N_23241,N_22989);
nor U26092 (N_26092,N_22386,N_22114);
nor U26093 (N_26093,N_23435,N_22694);
xor U26094 (N_26094,N_22641,N_22217);
xor U26095 (N_26095,N_23774,N_22209);
nor U26096 (N_26096,N_21550,N_23099);
or U26097 (N_26097,N_22873,N_23003);
or U26098 (N_26098,N_21654,N_21290);
and U26099 (N_26099,N_22450,N_22535);
and U26100 (N_26100,N_23283,N_21518);
or U26101 (N_26101,N_23091,N_22709);
or U26102 (N_26102,N_22006,N_23677);
nand U26103 (N_26103,N_22446,N_21706);
nand U26104 (N_26104,N_21945,N_21901);
nor U26105 (N_26105,N_22572,N_21478);
or U26106 (N_26106,N_22340,N_22395);
or U26107 (N_26107,N_21363,N_23857);
or U26108 (N_26108,N_21232,N_21480);
xor U26109 (N_26109,N_21638,N_23356);
nand U26110 (N_26110,N_22924,N_23815);
nor U26111 (N_26111,N_21904,N_23912);
and U26112 (N_26112,N_21562,N_23439);
nor U26113 (N_26113,N_23996,N_22081);
nand U26114 (N_26114,N_21946,N_22304);
xor U26115 (N_26115,N_21543,N_21695);
nand U26116 (N_26116,N_22929,N_22095);
xnor U26117 (N_26117,N_23404,N_22937);
or U26118 (N_26118,N_21559,N_22628);
nor U26119 (N_26119,N_22162,N_23105);
xnor U26120 (N_26120,N_21321,N_21088);
nor U26121 (N_26121,N_22955,N_23296);
xor U26122 (N_26122,N_23446,N_21239);
xor U26123 (N_26123,N_21484,N_21313);
nand U26124 (N_26124,N_22257,N_22411);
nand U26125 (N_26125,N_22669,N_21938);
or U26126 (N_26126,N_21601,N_21170);
and U26127 (N_26127,N_21609,N_22093);
nor U26128 (N_26128,N_23742,N_21748);
nand U26129 (N_26129,N_21267,N_22357);
xor U26130 (N_26130,N_23670,N_21089);
xnor U26131 (N_26131,N_22004,N_23316);
xnor U26132 (N_26132,N_22219,N_21517);
xor U26133 (N_26133,N_21369,N_23878);
and U26134 (N_26134,N_22707,N_21288);
nor U26135 (N_26135,N_21241,N_22494);
and U26136 (N_26136,N_21130,N_21812);
or U26137 (N_26137,N_21384,N_22822);
xor U26138 (N_26138,N_21874,N_22298);
xnor U26139 (N_26139,N_22434,N_21963);
nand U26140 (N_26140,N_21009,N_21497);
xnor U26141 (N_26141,N_23808,N_22098);
nor U26142 (N_26142,N_22116,N_23669);
nand U26143 (N_26143,N_23138,N_23222);
and U26144 (N_26144,N_22797,N_21300);
or U26145 (N_26145,N_23155,N_21916);
xor U26146 (N_26146,N_22306,N_22501);
nor U26147 (N_26147,N_23294,N_22807);
xnor U26148 (N_26148,N_22913,N_23216);
and U26149 (N_26149,N_22907,N_22500);
and U26150 (N_26150,N_23759,N_21973);
or U26151 (N_26151,N_23613,N_23164);
or U26152 (N_26152,N_21532,N_23841);
and U26153 (N_26153,N_21626,N_23848);
xor U26154 (N_26154,N_22955,N_23120);
and U26155 (N_26155,N_21710,N_23700);
nor U26156 (N_26156,N_22756,N_22339);
xor U26157 (N_26157,N_21062,N_22521);
and U26158 (N_26158,N_21595,N_23162);
or U26159 (N_26159,N_22099,N_23219);
or U26160 (N_26160,N_23504,N_21572);
and U26161 (N_26161,N_21082,N_23270);
or U26162 (N_26162,N_23094,N_23358);
and U26163 (N_26163,N_21903,N_21175);
nor U26164 (N_26164,N_22822,N_21459);
nor U26165 (N_26165,N_22539,N_23982);
xnor U26166 (N_26166,N_21494,N_23290);
or U26167 (N_26167,N_23346,N_21149);
nand U26168 (N_26168,N_22361,N_22915);
and U26169 (N_26169,N_23560,N_22630);
xor U26170 (N_26170,N_22902,N_21793);
nand U26171 (N_26171,N_23959,N_21116);
nor U26172 (N_26172,N_23287,N_21433);
xnor U26173 (N_26173,N_23369,N_22822);
nor U26174 (N_26174,N_21177,N_21749);
nand U26175 (N_26175,N_23647,N_22060);
nor U26176 (N_26176,N_22388,N_21363);
nand U26177 (N_26177,N_22210,N_21368);
nor U26178 (N_26178,N_22393,N_22466);
or U26179 (N_26179,N_21961,N_23843);
and U26180 (N_26180,N_22921,N_23698);
and U26181 (N_26181,N_22744,N_23762);
nand U26182 (N_26182,N_23212,N_23037);
or U26183 (N_26183,N_23059,N_21718);
nand U26184 (N_26184,N_21671,N_23695);
xnor U26185 (N_26185,N_21361,N_21587);
or U26186 (N_26186,N_23481,N_22787);
or U26187 (N_26187,N_22290,N_23483);
and U26188 (N_26188,N_22109,N_23174);
nand U26189 (N_26189,N_22541,N_21581);
or U26190 (N_26190,N_21680,N_23356);
and U26191 (N_26191,N_23321,N_23376);
nor U26192 (N_26192,N_23126,N_22302);
or U26193 (N_26193,N_21122,N_22436);
nor U26194 (N_26194,N_22298,N_23603);
nand U26195 (N_26195,N_22484,N_23071);
nor U26196 (N_26196,N_21077,N_23953);
or U26197 (N_26197,N_21419,N_22943);
or U26198 (N_26198,N_23574,N_23217);
nand U26199 (N_26199,N_23571,N_22973);
xnor U26200 (N_26200,N_23109,N_21154);
nor U26201 (N_26201,N_23891,N_21471);
and U26202 (N_26202,N_23435,N_22216);
and U26203 (N_26203,N_21067,N_23645);
nor U26204 (N_26204,N_21622,N_22846);
or U26205 (N_26205,N_21872,N_21973);
xnor U26206 (N_26206,N_21490,N_23584);
nand U26207 (N_26207,N_23413,N_21208);
xor U26208 (N_26208,N_23673,N_23478);
xor U26209 (N_26209,N_22569,N_21942);
nand U26210 (N_26210,N_22552,N_22487);
nor U26211 (N_26211,N_21063,N_22047);
nor U26212 (N_26212,N_23909,N_23872);
or U26213 (N_26213,N_23689,N_21299);
xor U26214 (N_26214,N_22871,N_21530);
and U26215 (N_26215,N_22096,N_22605);
nor U26216 (N_26216,N_21390,N_23048);
and U26217 (N_26217,N_22720,N_21718);
nand U26218 (N_26218,N_23588,N_21775);
nand U26219 (N_26219,N_22771,N_21597);
xnor U26220 (N_26220,N_22353,N_22339);
xor U26221 (N_26221,N_23483,N_21834);
xor U26222 (N_26222,N_22735,N_22026);
nand U26223 (N_26223,N_21152,N_21446);
xnor U26224 (N_26224,N_22607,N_22017);
nand U26225 (N_26225,N_23093,N_21160);
and U26226 (N_26226,N_23402,N_22183);
and U26227 (N_26227,N_23516,N_22919);
nand U26228 (N_26228,N_21987,N_23200);
nor U26229 (N_26229,N_23801,N_21178);
xor U26230 (N_26230,N_21455,N_22209);
and U26231 (N_26231,N_22504,N_22816);
or U26232 (N_26232,N_23036,N_23177);
xnor U26233 (N_26233,N_23620,N_21091);
or U26234 (N_26234,N_23166,N_21210);
xnor U26235 (N_26235,N_23130,N_22213);
nor U26236 (N_26236,N_21524,N_21312);
or U26237 (N_26237,N_23008,N_21368);
nor U26238 (N_26238,N_23690,N_22056);
xnor U26239 (N_26239,N_22529,N_23160);
nor U26240 (N_26240,N_21374,N_23369);
nand U26241 (N_26241,N_21913,N_22162);
xnor U26242 (N_26242,N_22734,N_22365);
xnor U26243 (N_26243,N_22039,N_21628);
and U26244 (N_26244,N_21343,N_22900);
or U26245 (N_26245,N_23238,N_22952);
nor U26246 (N_26246,N_23188,N_22773);
and U26247 (N_26247,N_23660,N_23465);
nand U26248 (N_26248,N_22798,N_22906);
and U26249 (N_26249,N_23049,N_23499);
nor U26250 (N_26250,N_22618,N_22176);
and U26251 (N_26251,N_21984,N_22743);
xnor U26252 (N_26252,N_22786,N_21497);
nor U26253 (N_26253,N_23659,N_22074);
nand U26254 (N_26254,N_21096,N_21395);
or U26255 (N_26255,N_22282,N_22199);
and U26256 (N_26256,N_21449,N_22614);
and U26257 (N_26257,N_21730,N_23534);
nand U26258 (N_26258,N_23161,N_22422);
xnor U26259 (N_26259,N_22656,N_21978);
nor U26260 (N_26260,N_23145,N_23766);
nand U26261 (N_26261,N_21199,N_23263);
nor U26262 (N_26262,N_23217,N_22939);
or U26263 (N_26263,N_22404,N_21730);
and U26264 (N_26264,N_22080,N_23658);
or U26265 (N_26265,N_22112,N_23833);
and U26266 (N_26266,N_22644,N_21303);
nor U26267 (N_26267,N_23223,N_22373);
xor U26268 (N_26268,N_22519,N_21302);
nand U26269 (N_26269,N_22410,N_22674);
and U26270 (N_26270,N_22570,N_21279);
nor U26271 (N_26271,N_21036,N_21363);
nand U26272 (N_26272,N_22354,N_22988);
xor U26273 (N_26273,N_23878,N_23372);
nor U26274 (N_26274,N_22791,N_22566);
xor U26275 (N_26275,N_23921,N_21035);
xor U26276 (N_26276,N_21536,N_22955);
nand U26277 (N_26277,N_22630,N_23505);
xnor U26278 (N_26278,N_22935,N_22016);
and U26279 (N_26279,N_21340,N_22775);
nor U26280 (N_26280,N_23570,N_21765);
nand U26281 (N_26281,N_23937,N_23970);
nand U26282 (N_26282,N_23383,N_21540);
or U26283 (N_26283,N_21767,N_21004);
xor U26284 (N_26284,N_21894,N_21530);
nand U26285 (N_26285,N_21227,N_21217);
or U26286 (N_26286,N_21359,N_21578);
xor U26287 (N_26287,N_21031,N_22461);
nor U26288 (N_26288,N_21464,N_21481);
or U26289 (N_26289,N_22810,N_23608);
and U26290 (N_26290,N_22776,N_22901);
nor U26291 (N_26291,N_23984,N_22063);
and U26292 (N_26292,N_23393,N_21453);
xnor U26293 (N_26293,N_21762,N_23562);
or U26294 (N_26294,N_23006,N_23543);
nor U26295 (N_26295,N_21886,N_23159);
nor U26296 (N_26296,N_23573,N_22921);
nor U26297 (N_26297,N_23339,N_22996);
nand U26298 (N_26298,N_21596,N_23052);
nand U26299 (N_26299,N_21073,N_22526);
or U26300 (N_26300,N_23002,N_23893);
xor U26301 (N_26301,N_21597,N_23662);
or U26302 (N_26302,N_22110,N_23216);
nor U26303 (N_26303,N_23020,N_22131);
xor U26304 (N_26304,N_23293,N_21171);
or U26305 (N_26305,N_23591,N_22829);
nand U26306 (N_26306,N_22806,N_21988);
nor U26307 (N_26307,N_23012,N_21966);
xnor U26308 (N_26308,N_21674,N_21889);
or U26309 (N_26309,N_23577,N_22516);
xor U26310 (N_26310,N_21094,N_21496);
nor U26311 (N_26311,N_22041,N_21817);
and U26312 (N_26312,N_23840,N_22486);
or U26313 (N_26313,N_22412,N_21247);
nand U26314 (N_26314,N_22474,N_23985);
or U26315 (N_26315,N_22406,N_22461);
nand U26316 (N_26316,N_21354,N_21485);
nand U26317 (N_26317,N_22791,N_21369);
nand U26318 (N_26318,N_23211,N_22566);
nor U26319 (N_26319,N_21987,N_21450);
nor U26320 (N_26320,N_22933,N_21624);
nand U26321 (N_26321,N_21475,N_21555);
nand U26322 (N_26322,N_22208,N_23877);
xnor U26323 (N_26323,N_21174,N_21060);
nor U26324 (N_26324,N_21458,N_21701);
and U26325 (N_26325,N_23573,N_23506);
nand U26326 (N_26326,N_22027,N_21859);
and U26327 (N_26327,N_22343,N_21031);
xnor U26328 (N_26328,N_21466,N_23852);
nand U26329 (N_26329,N_22612,N_21963);
or U26330 (N_26330,N_21473,N_21575);
nand U26331 (N_26331,N_22589,N_21015);
and U26332 (N_26332,N_23267,N_23304);
nor U26333 (N_26333,N_22822,N_22206);
or U26334 (N_26334,N_21229,N_21943);
and U26335 (N_26335,N_22676,N_21383);
nor U26336 (N_26336,N_23341,N_22109);
nor U26337 (N_26337,N_22834,N_22403);
nand U26338 (N_26338,N_22650,N_23399);
nor U26339 (N_26339,N_21880,N_23519);
or U26340 (N_26340,N_21195,N_23915);
nor U26341 (N_26341,N_23691,N_21872);
nor U26342 (N_26342,N_22087,N_23927);
and U26343 (N_26343,N_23732,N_23656);
and U26344 (N_26344,N_21494,N_21393);
and U26345 (N_26345,N_21874,N_22655);
and U26346 (N_26346,N_22308,N_22371);
nor U26347 (N_26347,N_23469,N_21683);
or U26348 (N_26348,N_21289,N_22797);
nor U26349 (N_26349,N_23444,N_21700);
or U26350 (N_26350,N_22323,N_22847);
nor U26351 (N_26351,N_22426,N_21366);
and U26352 (N_26352,N_21018,N_23736);
and U26353 (N_26353,N_22772,N_21064);
nor U26354 (N_26354,N_23940,N_22598);
nand U26355 (N_26355,N_22094,N_22866);
nand U26356 (N_26356,N_21278,N_21655);
or U26357 (N_26357,N_23231,N_22666);
or U26358 (N_26358,N_21382,N_21723);
nor U26359 (N_26359,N_22339,N_22875);
xnor U26360 (N_26360,N_21816,N_23399);
xor U26361 (N_26361,N_22429,N_21240);
nand U26362 (N_26362,N_23536,N_23192);
nand U26363 (N_26363,N_22071,N_22313);
nand U26364 (N_26364,N_23278,N_23674);
nor U26365 (N_26365,N_21520,N_23611);
nor U26366 (N_26366,N_21142,N_22847);
and U26367 (N_26367,N_21444,N_23068);
nor U26368 (N_26368,N_22383,N_23818);
nand U26369 (N_26369,N_22995,N_23810);
nand U26370 (N_26370,N_21127,N_22761);
or U26371 (N_26371,N_21682,N_23298);
or U26372 (N_26372,N_21395,N_22533);
and U26373 (N_26373,N_21188,N_22567);
xor U26374 (N_26374,N_21964,N_21780);
nand U26375 (N_26375,N_21243,N_22150);
and U26376 (N_26376,N_23131,N_22118);
nand U26377 (N_26377,N_21597,N_21734);
nand U26378 (N_26378,N_23043,N_23564);
xor U26379 (N_26379,N_23819,N_21145);
or U26380 (N_26380,N_21223,N_22730);
nand U26381 (N_26381,N_22703,N_22734);
or U26382 (N_26382,N_21827,N_22751);
nor U26383 (N_26383,N_22536,N_23074);
or U26384 (N_26384,N_21230,N_23905);
nand U26385 (N_26385,N_23739,N_23816);
or U26386 (N_26386,N_23462,N_23126);
xnor U26387 (N_26387,N_21401,N_21578);
xor U26388 (N_26388,N_23373,N_22000);
nand U26389 (N_26389,N_23296,N_23806);
or U26390 (N_26390,N_23492,N_21213);
nand U26391 (N_26391,N_21476,N_23130);
or U26392 (N_26392,N_21211,N_22208);
xnor U26393 (N_26393,N_21355,N_23263);
or U26394 (N_26394,N_23591,N_23619);
nor U26395 (N_26395,N_22760,N_23447);
nand U26396 (N_26396,N_22859,N_23053);
nand U26397 (N_26397,N_22149,N_22502);
xnor U26398 (N_26398,N_23143,N_21749);
nor U26399 (N_26399,N_22731,N_21312);
and U26400 (N_26400,N_22820,N_23040);
xnor U26401 (N_26401,N_23947,N_22849);
or U26402 (N_26402,N_23760,N_22631);
nor U26403 (N_26403,N_22799,N_21730);
and U26404 (N_26404,N_22681,N_22912);
and U26405 (N_26405,N_21899,N_23321);
nor U26406 (N_26406,N_22712,N_23227);
or U26407 (N_26407,N_22080,N_22425);
xor U26408 (N_26408,N_23640,N_23250);
and U26409 (N_26409,N_23619,N_23302);
nor U26410 (N_26410,N_22372,N_21697);
nor U26411 (N_26411,N_22798,N_23129);
nor U26412 (N_26412,N_23778,N_21084);
nand U26413 (N_26413,N_23727,N_22510);
and U26414 (N_26414,N_22390,N_23888);
nor U26415 (N_26415,N_21571,N_23277);
and U26416 (N_26416,N_21931,N_22659);
nand U26417 (N_26417,N_21792,N_21906);
nand U26418 (N_26418,N_21649,N_22310);
nand U26419 (N_26419,N_21706,N_21086);
and U26420 (N_26420,N_21717,N_22667);
nand U26421 (N_26421,N_22422,N_21506);
and U26422 (N_26422,N_23946,N_21348);
xnor U26423 (N_26423,N_22396,N_21139);
nand U26424 (N_26424,N_21064,N_23076);
and U26425 (N_26425,N_21110,N_22919);
and U26426 (N_26426,N_22299,N_23986);
nor U26427 (N_26427,N_23839,N_23235);
nand U26428 (N_26428,N_23767,N_23319);
or U26429 (N_26429,N_23756,N_22573);
or U26430 (N_26430,N_23206,N_23828);
xor U26431 (N_26431,N_22941,N_21998);
nor U26432 (N_26432,N_22753,N_21609);
and U26433 (N_26433,N_21681,N_23286);
nand U26434 (N_26434,N_23456,N_21842);
xor U26435 (N_26435,N_21729,N_23444);
nor U26436 (N_26436,N_23998,N_23465);
nand U26437 (N_26437,N_23991,N_23765);
xor U26438 (N_26438,N_22804,N_22165);
nand U26439 (N_26439,N_21042,N_23038);
xnor U26440 (N_26440,N_21588,N_21500);
and U26441 (N_26441,N_22989,N_22383);
nand U26442 (N_26442,N_21060,N_23376);
and U26443 (N_26443,N_22229,N_21444);
nor U26444 (N_26444,N_22703,N_23980);
nand U26445 (N_26445,N_21082,N_21485);
nand U26446 (N_26446,N_21413,N_23182);
and U26447 (N_26447,N_23287,N_23412);
nor U26448 (N_26448,N_23454,N_21781);
and U26449 (N_26449,N_22926,N_22417);
nor U26450 (N_26450,N_21231,N_22695);
nor U26451 (N_26451,N_23627,N_23999);
or U26452 (N_26452,N_22527,N_22248);
and U26453 (N_26453,N_21796,N_22883);
xor U26454 (N_26454,N_22326,N_22694);
or U26455 (N_26455,N_21690,N_21627);
nor U26456 (N_26456,N_23529,N_23062);
and U26457 (N_26457,N_23792,N_23616);
nand U26458 (N_26458,N_21215,N_23801);
and U26459 (N_26459,N_21381,N_23424);
and U26460 (N_26460,N_21485,N_23435);
or U26461 (N_26461,N_22663,N_22778);
nor U26462 (N_26462,N_23285,N_21971);
or U26463 (N_26463,N_21907,N_23099);
nand U26464 (N_26464,N_22862,N_21507);
and U26465 (N_26465,N_22668,N_21451);
nand U26466 (N_26466,N_23022,N_21559);
nand U26467 (N_26467,N_23424,N_22871);
nand U26468 (N_26468,N_22891,N_21570);
and U26469 (N_26469,N_23098,N_22343);
nor U26470 (N_26470,N_22716,N_21786);
nand U26471 (N_26471,N_22893,N_22631);
nor U26472 (N_26472,N_22615,N_22035);
xnor U26473 (N_26473,N_22750,N_22483);
and U26474 (N_26474,N_23692,N_21228);
xnor U26475 (N_26475,N_21179,N_23254);
or U26476 (N_26476,N_23305,N_22037);
or U26477 (N_26477,N_21797,N_22303);
nor U26478 (N_26478,N_21336,N_22046);
and U26479 (N_26479,N_22179,N_23054);
or U26480 (N_26480,N_22580,N_22197);
xnor U26481 (N_26481,N_22604,N_21486);
nor U26482 (N_26482,N_21495,N_21650);
nor U26483 (N_26483,N_23725,N_21649);
nor U26484 (N_26484,N_21743,N_21040);
and U26485 (N_26485,N_21898,N_21932);
or U26486 (N_26486,N_23287,N_23887);
nand U26487 (N_26487,N_21394,N_22776);
or U26488 (N_26488,N_22401,N_23274);
and U26489 (N_26489,N_21160,N_22016);
xnor U26490 (N_26490,N_23811,N_21180);
nand U26491 (N_26491,N_22179,N_21352);
or U26492 (N_26492,N_21272,N_21070);
nor U26493 (N_26493,N_22788,N_23511);
nand U26494 (N_26494,N_22062,N_21866);
xnor U26495 (N_26495,N_22165,N_23896);
and U26496 (N_26496,N_23222,N_23371);
xnor U26497 (N_26497,N_22901,N_21835);
xnor U26498 (N_26498,N_22009,N_22508);
and U26499 (N_26499,N_21137,N_22816);
nand U26500 (N_26500,N_23568,N_23038);
or U26501 (N_26501,N_22113,N_21684);
xnor U26502 (N_26502,N_21342,N_21059);
xor U26503 (N_26503,N_21772,N_21851);
xnor U26504 (N_26504,N_23244,N_22597);
nand U26505 (N_26505,N_22370,N_22792);
xor U26506 (N_26506,N_23106,N_22069);
or U26507 (N_26507,N_23413,N_21875);
and U26508 (N_26508,N_23189,N_21819);
xnor U26509 (N_26509,N_23816,N_21007);
nor U26510 (N_26510,N_23079,N_21161);
nor U26511 (N_26511,N_23970,N_22846);
and U26512 (N_26512,N_22429,N_22373);
xor U26513 (N_26513,N_22058,N_23779);
and U26514 (N_26514,N_21832,N_22878);
nand U26515 (N_26515,N_22436,N_23131);
or U26516 (N_26516,N_22822,N_21992);
nor U26517 (N_26517,N_23681,N_23118);
nor U26518 (N_26518,N_23375,N_23383);
xor U26519 (N_26519,N_22400,N_23720);
nand U26520 (N_26520,N_21692,N_23365);
nand U26521 (N_26521,N_21980,N_23159);
nand U26522 (N_26522,N_21678,N_23267);
or U26523 (N_26523,N_21679,N_21218);
and U26524 (N_26524,N_21585,N_21773);
nor U26525 (N_26525,N_21403,N_21154);
nand U26526 (N_26526,N_23848,N_23710);
xor U26527 (N_26527,N_23586,N_21790);
nor U26528 (N_26528,N_22855,N_21778);
nor U26529 (N_26529,N_23911,N_23233);
or U26530 (N_26530,N_23605,N_23198);
nor U26531 (N_26531,N_21978,N_21669);
nand U26532 (N_26532,N_23587,N_23784);
xor U26533 (N_26533,N_21601,N_22755);
nand U26534 (N_26534,N_22576,N_21001);
nor U26535 (N_26535,N_22022,N_22857);
xnor U26536 (N_26536,N_22519,N_23959);
and U26537 (N_26537,N_23915,N_21661);
nor U26538 (N_26538,N_22075,N_21886);
or U26539 (N_26539,N_23968,N_21492);
xor U26540 (N_26540,N_21418,N_21636);
nor U26541 (N_26541,N_23950,N_22319);
xor U26542 (N_26542,N_22354,N_21333);
nand U26543 (N_26543,N_22060,N_22579);
or U26544 (N_26544,N_21488,N_22734);
and U26545 (N_26545,N_23840,N_23203);
xnor U26546 (N_26546,N_23810,N_22782);
xnor U26547 (N_26547,N_22493,N_22044);
and U26548 (N_26548,N_22687,N_22999);
xor U26549 (N_26549,N_23104,N_21242);
or U26550 (N_26550,N_23269,N_21793);
nand U26551 (N_26551,N_22522,N_23144);
and U26552 (N_26552,N_23497,N_22006);
nor U26553 (N_26553,N_22199,N_21848);
xor U26554 (N_26554,N_21719,N_22769);
and U26555 (N_26555,N_22605,N_23530);
and U26556 (N_26556,N_22250,N_22638);
and U26557 (N_26557,N_22709,N_21432);
xnor U26558 (N_26558,N_22807,N_21929);
and U26559 (N_26559,N_21570,N_23229);
nor U26560 (N_26560,N_21929,N_22009);
or U26561 (N_26561,N_22278,N_23326);
nand U26562 (N_26562,N_21789,N_23147);
nor U26563 (N_26563,N_22665,N_21541);
xor U26564 (N_26564,N_23943,N_22629);
and U26565 (N_26565,N_23388,N_23139);
xor U26566 (N_26566,N_22694,N_22823);
nor U26567 (N_26567,N_22518,N_21932);
or U26568 (N_26568,N_21363,N_21927);
xor U26569 (N_26569,N_21176,N_22143);
or U26570 (N_26570,N_23694,N_22427);
nor U26571 (N_26571,N_21201,N_23382);
nor U26572 (N_26572,N_22078,N_22870);
and U26573 (N_26573,N_21016,N_23121);
nand U26574 (N_26574,N_22360,N_21600);
xor U26575 (N_26575,N_23154,N_21742);
or U26576 (N_26576,N_22834,N_21282);
xor U26577 (N_26577,N_21628,N_21235);
nor U26578 (N_26578,N_22753,N_21697);
or U26579 (N_26579,N_22789,N_21186);
and U26580 (N_26580,N_23453,N_23048);
nor U26581 (N_26581,N_22708,N_21753);
and U26582 (N_26582,N_21697,N_22574);
xor U26583 (N_26583,N_22124,N_21640);
xnor U26584 (N_26584,N_21415,N_22198);
xor U26585 (N_26585,N_21800,N_21922);
or U26586 (N_26586,N_21453,N_23138);
and U26587 (N_26587,N_21952,N_22569);
xnor U26588 (N_26588,N_22071,N_23100);
and U26589 (N_26589,N_21863,N_21554);
xor U26590 (N_26590,N_22633,N_23542);
nand U26591 (N_26591,N_23694,N_22918);
nand U26592 (N_26592,N_23424,N_22215);
xor U26593 (N_26593,N_22014,N_22894);
nand U26594 (N_26594,N_22862,N_21341);
nand U26595 (N_26595,N_23289,N_23134);
and U26596 (N_26596,N_22483,N_23653);
nor U26597 (N_26597,N_23660,N_23371);
and U26598 (N_26598,N_23005,N_22274);
or U26599 (N_26599,N_21809,N_22578);
nand U26600 (N_26600,N_22879,N_22832);
and U26601 (N_26601,N_22200,N_21737);
nor U26602 (N_26602,N_21109,N_21301);
nor U26603 (N_26603,N_21824,N_22685);
and U26604 (N_26604,N_23717,N_22983);
xor U26605 (N_26605,N_21305,N_22602);
nor U26606 (N_26606,N_22968,N_23528);
nand U26607 (N_26607,N_21973,N_23150);
nand U26608 (N_26608,N_21264,N_21906);
or U26609 (N_26609,N_23575,N_21657);
or U26610 (N_26610,N_21050,N_21591);
and U26611 (N_26611,N_21878,N_21031);
and U26612 (N_26612,N_21646,N_22295);
nor U26613 (N_26613,N_22311,N_23554);
or U26614 (N_26614,N_23583,N_22678);
xor U26615 (N_26615,N_21775,N_21745);
or U26616 (N_26616,N_22027,N_23942);
and U26617 (N_26617,N_21489,N_23285);
xnor U26618 (N_26618,N_23271,N_21384);
nand U26619 (N_26619,N_21255,N_21174);
xnor U26620 (N_26620,N_23219,N_22458);
nor U26621 (N_26621,N_21630,N_22354);
or U26622 (N_26622,N_22511,N_22763);
or U26623 (N_26623,N_22642,N_21319);
nor U26624 (N_26624,N_23329,N_22651);
and U26625 (N_26625,N_22170,N_23040);
xnor U26626 (N_26626,N_23414,N_22101);
or U26627 (N_26627,N_23346,N_23446);
nor U26628 (N_26628,N_22766,N_23788);
nand U26629 (N_26629,N_22567,N_22581);
and U26630 (N_26630,N_23523,N_22851);
nor U26631 (N_26631,N_22262,N_21344);
or U26632 (N_26632,N_22650,N_22623);
nor U26633 (N_26633,N_22560,N_21767);
xor U26634 (N_26634,N_21810,N_23093);
xnor U26635 (N_26635,N_22753,N_22829);
xor U26636 (N_26636,N_21760,N_23162);
nor U26637 (N_26637,N_21880,N_21421);
nand U26638 (N_26638,N_21066,N_21523);
and U26639 (N_26639,N_21966,N_23148);
xnor U26640 (N_26640,N_21814,N_22510);
and U26641 (N_26641,N_22942,N_23771);
nor U26642 (N_26642,N_23249,N_21419);
nand U26643 (N_26643,N_21243,N_21965);
or U26644 (N_26644,N_23688,N_21452);
nor U26645 (N_26645,N_22758,N_23232);
nor U26646 (N_26646,N_23843,N_23227);
and U26647 (N_26647,N_22964,N_21165);
nor U26648 (N_26648,N_23538,N_21815);
xnor U26649 (N_26649,N_21493,N_22832);
nor U26650 (N_26650,N_23691,N_23021);
nand U26651 (N_26651,N_21030,N_21080);
nor U26652 (N_26652,N_22973,N_21889);
and U26653 (N_26653,N_22575,N_21108);
or U26654 (N_26654,N_22349,N_22789);
nor U26655 (N_26655,N_22136,N_22406);
or U26656 (N_26656,N_22420,N_22699);
or U26657 (N_26657,N_21720,N_21254);
nand U26658 (N_26658,N_23590,N_21055);
nor U26659 (N_26659,N_21640,N_22559);
nand U26660 (N_26660,N_21090,N_22378);
nor U26661 (N_26661,N_23697,N_23219);
nand U26662 (N_26662,N_22813,N_23967);
xor U26663 (N_26663,N_21912,N_22161);
nor U26664 (N_26664,N_21226,N_21416);
nand U26665 (N_26665,N_21500,N_23958);
or U26666 (N_26666,N_23798,N_23732);
nand U26667 (N_26667,N_22589,N_23260);
and U26668 (N_26668,N_22572,N_23044);
nand U26669 (N_26669,N_23319,N_22932);
or U26670 (N_26670,N_23729,N_23557);
and U26671 (N_26671,N_22452,N_21660);
nand U26672 (N_26672,N_21834,N_23679);
nor U26673 (N_26673,N_23595,N_21947);
or U26674 (N_26674,N_21512,N_22986);
nor U26675 (N_26675,N_22919,N_21598);
nand U26676 (N_26676,N_23141,N_21650);
or U26677 (N_26677,N_21057,N_22074);
nor U26678 (N_26678,N_22636,N_21601);
xnor U26679 (N_26679,N_23354,N_21233);
and U26680 (N_26680,N_22871,N_21377);
nand U26681 (N_26681,N_21390,N_23367);
xor U26682 (N_26682,N_21115,N_21345);
xor U26683 (N_26683,N_21801,N_22417);
or U26684 (N_26684,N_22415,N_22944);
or U26685 (N_26685,N_23200,N_21426);
nand U26686 (N_26686,N_22205,N_21006);
xor U26687 (N_26687,N_23854,N_23966);
or U26688 (N_26688,N_21167,N_22452);
and U26689 (N_26689,N_23791,N_22150);
nand U26690 (N_26690,N_23298,N_21820);
xnor U26691 (N_26691,N_21165,N_23230);
nor U26692 (N_26692,N_23647,N_21489);
nor U26693 (N_26693,N_21193,N_23455);
nor U26694 (N_26694,N_22299,N_22894);
nand U26695 (N_26695,N_22549,N_22130);
nor U26696 (N_26696,N_22977,N_23193);
and U26697 (N_26697,N_21536,N_21864);
and U26698 (N_26698,N_22042,N_23773);
xor U26699 (N_26699,N_22534,N_21805);
and U26700 (N_26700,N_23982,N_22343);
and U26701 (N_26701,N_23957,N_22454);
or U26702 (N_26702,N_23064,N_23397);
nor U26703 (N_26703,N_21575,N_22638);
xnor U26704 (N_26704,N_21725,N_21478);
nand U26705 (N_26705,N_22029,N_23383);
xor U26706 (N_26706,N_21872,N_21782);
nor U26707 (N_26707,N_22522,N_21639);
xnor U26708 (N_26708,N_23407,N_22128);
xnor U26709 (N_26709,N_23692,N_21589);
or U26710 (N_26710,N_23612,N_22890);
nand U26711 (N_26711,N_22374,N_22986);
and U26712 (N_26712,N_21410,N_23099);
nand U26713 (N_26713,N_23631,N_21556);
nand U26714 (N_26714,N_22301,N_22502);
nand U26715 (N_26715,N_22159,N_21743);
or U26716 (N_26716,N_21114,N_22215);
xnor U26717 (N_26717,N_23684,N_22736);
or U26718 (N_26718,N_23395,N_22661);
and U26719 (N_26719,N_21927,N_22032);
nor U26720 (N_26720,N_22509,N_23036);
and U26721 (N_26721,N_23448,N_21810);
or U26722 (N_26722,N_23215,N_21505);
nor U26723 (N_26723,N_22760,N_21358);
or U26724 (N_26724,N_21900,N_22298);
nor U26725 (N_26725,N_21177,N_21226);
nor U26726 (N_26726,N_23647,N_22131);
xor U26727 (N_26727,N_22169,N_23694);
xnor U26728 (N_26728,N_22874,N_23169);
xor U26729 (N_26729,N_23414,N_21921);
or U26730 (N_26730,N_21625,N_23031);
and U26731 (N_26731,N_22542,N_23403);
nor U26732 (N_26732,N_23985,N_23400);
nor U26733 (N_26733,N_21778,N_23161);
or U26734 (N_26734,N_23786,N_21955);
xor U26735 (N_26735,N_23633,N_22927);
nor U26736 (N_26736,N_21274,N_21194);
xor U26737 (N_26737,N_22917,N_21870);
nand U26738 (N_26738,N_23347,N_21479);
and U26739 (N_26739,N_23077,N_21570);
nor U26740 (N_26740,N_23020,N_21956);
or U26741 (N_26741,N_22550,N_22958);
nor U26742 (N_26742,N_21368,N_21203);
nor U26743 (N_26743,N_23756,N_23565);
or U26744 (N_26744,N_21153,N_22334);
xor U26745 (N_26745,N_21396,N_23968);
and U26746 (N_26746,N_23613,N_23267);
nand U26747 (N_26747,N_23715,N_21719);
nand U26748 (N_26748,N_23943,N_23351);
nor U26749 (N_26749,N_23415,N_21630);
or U26750 (N_26750,N_21042,N_21004);
nor U26751 (N_26751,N_22812,N_21585);
xor U26752 (N_26752,N_21842,N_21339);
and U26753 (N_26753,N_23526,N_21197);
xor U26754 (N_26754,N_23946,N_23016);
nor U26755 (N_26755,N_21776,N_22605);
xor U26756 (N_26756,N_22618,N_21798);
or U26757 (N_26757,N_22199,N_23860);
nand U26758 (N_26758,N_21233,N_22846);
xor U26759 (N_26759,N_23541,N_23339);
or U26760 (N_26760,N_21436,N_22668);
xor U26761 (N_26761,N_22941,N_21802);
nor U26762 (N_26762,N_22158,N_22676);
nor U26763 (N_26763,N_22889,N_22395);
or U26764 (N_26764,N_21831,N_21609);
nand U26765 (N_26765,N_21944,N_22938);
and U26766 (N_26766,N_23277,N_23728);
xor U26767 (N_26767,N_23493,N_23277);
nand U26768 (N_26768,N_21833,N_21525);
xnor U26769 (N_26769,N_21538,N_21291);
xor U26770 (N_26770,N_22001,N_22572);
or U26771 (N_26771,N_21928,N_23109);
or U26772 (N_26772,N_21219,N_21669);
xor U26773 (N_26773,N_23460,N_22945);
nand U26774 (N_26774,N_23012,N_23859);
and U26775 (N_26775,N_21796,N_22898);
nor U26776 (N_26776,N_23784,N_22154);
nor U26777 (N_26777,N_21302,N_23014);
xor U26778 (N_26778,N_23461,N_23230);
or U26779 (N_26779,N_22105,N_21095);
or U26780 (N_26780,N_22887,N_23725);
and U26781 (N_26781,N_23651,N_22807);
and U26782 (N_26782,N_22703,N_22694);
or U26783 (N_26783,N_22893,N_21550);
or U26784 (N_26784,N_21304,N_22906);
xnor U26785 (N_26785,N_21452,N_22290);
or U26786 (N_26786,N_22923,N_23323);
and U26787 (N_26787,N_21885,N_21173);
nand U26788 (N_26788,N_22604,N_21647);
nand U26789 (N_26789,N_23665,N_21401);
nor U26790 (N_26790,N_23199,N_22601);
nor U26791 (N_26791,N_23563,N_23136);
and U26792 (N_26792,N_23172,N_23201);
nor U26793 (N_26793,N_22136,N_22104);
and U26794 (N_26794,N_23541,N_21008);
nand U26795 (N_26795,N_22367,N_23441);
nand U26796 (N_26796,N_21605,N_21783);
and U26797 (N_26797,N_21883,N_22524);
nand U26798 (N_26798,N_21358,N_21322);
nand U26799 (N_26799,N_21494,N_22051);
xnor U26800 (N_26800,N_22913,N_22781);
xor U26801 (N_26801,N_21180,N_22848);
xor U26802 (N_26802,N_21452,N_21298);
and U26803 (N_26803,N_22294,N_22337);
nand U26804 (N_26804,N_23574,N_22292);
or U26805 (N_26805,N_23438,N_22796);
or U26806 (N_26806,N_21429,N_22410);
nor U26807 (N_26807,N_23846,N_21907);
and U26808 (N_26808,N_22189,N_23048);
and U26809 (N_26809,N_21599,N_21947);
or U26810 (N_26810,N_23849,N_23841);
nor U26811 (N_26811,N_22962,N_23304);
xor U26812 (N_26812,N_22027,N_23235);
xor U26813 (N_26813,N_23228,N_21197);
nand U26814 (N_26814,N_23925,N_22225);
xnor U26815 (N_26815,N_21020,N_21229);
and U26816 (N_26816,N_22977,N_21106);
nand U26817 (N_26817,N_23683,N_22306);
nand U26818 (N_26818,N_23860,N_22866);
nor U26819 (N_26819,N_23467,N_21288);
and U26820 (N_26820,N_22425,N_21391);
and U26821 (N_26821,N_23024,N_23364);
xor U26822 (N_26822,N_23426,N_21073);
nor U26823 (N_26823,N_21833,N_23583);
nor U26824 (N_26824,N_23529,N_23264);
nand U26825 (N_26825,N_23087,N_23245);
and U26826 (N_26826,N_21040,N_22269);
xnor U26827 (N_26827,N_21751,N_22527);
xor U26828 (N_26828,N_22989,N_23156);
and U26829 (N_26829,N_22199,N_23771);
xnor U26830 (N_26830,N_23125,N_21578);
and U26831 (N_26831,N_22706,N_23686);
nor U26832 (N_26832,N_21490,N_21699);
or U26833 (N_26833,N_22607,N_21395);
nand U26834 (N_26834,N_23878,N_23519);
nor U26835 (N_26835,N_21208,N_21663);
and U26836 (N_26836,N_22161,N_22594);
nand U26837 (N_26837,N_21251,N_23178);
or U26838 (N_26838,N_21141,N_23097);
or U26839 (N_26839,N_23343,N_23953);
nor U26840 (N_26840,N_23596,N_22492);
or U26841 (N_26841,N_22575,N_21429);
nand U26842 (N_26842,N_22173,N_23675);
or U26843 (N_26843,N_23292,N_21855);
nand U26844 (N_26844,N_23462,N_21463);
xnor U26845 (N_26845,N_22442,N_23514);
nor U26846 (N_26846,N_22080,N_22288);
xor U26847 (N_26847,N_22606,N_23188);
xnor U26848 (N_26848,N_22402,N_23336);
nor U26849 (N_26849,N_22512,N_23122);
and U26850 (N_26850,N_21620,N_23829);
xor U26851 (N_26851,N_22407,N_21966);
and U26852 (N_26852,N_23085,N_21976);
xnor U26853 (N_26853,N_21050,N_22183);
nand U26854 (N_26854,N_23433,N_21484);
xor U26855 (N_26855,N_22656,N_22150);
nor U26856 (N_26856,N_21544,N_22789);
nor U26857 (N_26857,N_23847,N_21028);
and U26858 (N_26858,N_23475,N_23685);
nand U26859 (N_26859,N_23483,N_23277);
nand U26860 (N_26860,N_22032,N_21507);
and U26861 (N_26861,N_22234,N_23640);
and U26862 (N_26862,N_22708,N_22387);
nor U26863 (N_26863,N_23264,N_23818);
nor U26864 (N_26864,N_23505,N_21449);
nand U26865 (N_26865,N_22724,N_23398);
nor U26866 (N_26866,N_22666,N_23532);
xnor U26867 (N_26867,N_23163,N_23248);
or U26868 (N_26868,N_21343,N_21981);
nand U26869 (N_26869,N_22689,N_21044);
xor U26870 (N_26870,N_22467,N_23640);
or U26871 (N_26871,N_23717,N_21038);
or U26872 (N_26872,N_22691,N_22858);
nand U26873 (N_26873,N_23130,N_23113);
xnor U26874 (N_26874,N_21450,N_21582);
xor U26875 (N_26875,N_21381,N_22155);
nor U26876 (N_26876,N_21966,N_22231);
or U26877 (N_26877,N_21661,N_22950);
xnor U26878 (N_26878,N_23853,N_22103);
xnor U26879 (N_26879,N_21869,N_22026);
or U26880 (N_26880,N_23573,N_22799);
nor U26881 (N_26881,N_23976,N_21714);
and U26882 (N_26882,N_21690,N_22063);
nor U26883 (N_26883,N_23199,N_21799);
nor U26884 (N_26884,N_21665,N_21791);
nor U26885 (N_26885,N_22285,N_21685);
and U26886 (N_26886,N_23019,N_21888);
and U26887 (N_26887,N_23529,N_23722);
xor U26888 (N_26888,N_23707,N_23479);
xor U26889 (N_26889,N_22937,N_22769);
nor U26890 (N_26890,N_22664,N_22444);
or U26891 (N_26891,N_23900,N_23738);
and U26892 (N_26892,N_21907,N_22144);
xnor U26893 (N_26893,N_21498,N_23407);
nand U26894 (N_26894,N_23731,N_21091);
nand U26895 (N_26895,N_22915,N_23313);
xnor U26896 (N_26896,N_21624,N_23224);
xor U26897 (N_26897,N_22194,N_22601);
nand U26898 (N_26898,N_23673,N_21069);
and U26899 (N_26899,N_22259,N_23710);
and U26900 (N_26900,N_22118,N_22317);
xor U26901 (N_26901,N_22131,N_22137);
or U26902 (N_26902,N_22200,N_21360);
nor U26903 (N_26903,N_22096,N_23381);
nor U26904 (N_26904,N_23041,N_22919);
nand U26905 (N_26905,N_23986,N_23584);
xnor U26906 (N_26906,N_21313,N_23977);
or U26907 (N_26907,N_22462,N_22232);
xnor U26908 (N_26908,N_23475,N_23997);
and U26909 (N_26909,N_21244,N_23901);
nor U26910 (N_26910,N_23658,N_21926);
xor U26911 (N_26911,N_22001,N_22482);
nor U26912 (N_26912,N_22526,N_22320);
nor U26913 (N_26913,N_21353,N_23119);
nor U26914 (N_26914,N_22129,N_21776);
and U26915 (N_26915,N_23189,N_22422);
xnor U26916 (N_26916,N_21638,N_22025);
xor U26917 (N_26917,N_23040,N_21104);
nand U26918 (N_26918,N_21563,N_23232);
nand U26919 (N_26919,N_22659,N_21636);
xnor U26920 (N_26920,N_22011,N_22779);
nand U26921 (N_26921,N_21304,N_23753);
xnor U26922 (N_26922,N_22389,N_23081);
or U26923 (N_26923,N_21515,N_21930);
or U26924 (N_26924,N_22458,N_23974);
nor U26925 (N_26925,N_23331,N_21598);
nand U26926 (N_26926,N_22572,N_21142);
or U26927 (N_26927,N_23102,N_23859);
nor U26928 (N_26928,N_21070,N_22866);
nand U26929 (N_26929,N_22475,N_23468);
or U26930 (N_26930,N_22130,N_23683);
and U26931 (N_26931,N_22232,N_21071);
xnor U26932 (N_26932,N_22009,N_22755);
nor U26933 (N_26933,N_22540,N_23039);
and U26934 (N_26934,N_23742,N_23734);
xnor U26935 (N_26935,N_21414,N_21380);
xor U26936 (N_26936,N_21844,N_23075);
and U26937 (N_26937,N_23750,N_21296);
nor U26938 (N_26938,N_21544,N_23689);
or U26939 (N_26939,N_21078,N_23745);
nand U26940 (N_26940,N_21812,N_22700);
nor U26941 (N_26941,N_23546,N_23584);
and U26942 (N_26942,N_21710,N_23459);
nor U26943 (N_26943,N_23451,N_21694);
and U26944 (N_26944,N_23545,N_23959);
and U26945 (N_26945,N_22761,N_22709);
and U26946 (N_26946,N_23743,N_21988);
or U26947 (N_26947,N_23040,N_21219);
nand U26948 (N_26948,N_21708,N_23458);
nand U26949 (N_26949,N_23935,N_22369);
nand U26950 (N_26950,N_22084,N_22645);
xnor U26951 (N_26951,N_21663,N_21721);
xor U26952 (N_26952,N_23754,N_22650);
nor U26953 (N_26953,N_21340,N_23391);
xnor U26954 (N_26954,N_23030,N_22554);
and U26955 (N_26955,N_21464,N_22265);
nand U26956 (N_26956,N_23098,N_23627);
and U26957 (N_26957,N_22326,N_23369);
xnor U26958 (N_26958,N_22237,N_22658);
and U26959 (N_26959,N_21724,N_23079);
or U26960 (N_26960,N_22961,N_22764);
nor U26961 (N_26961,N_22770,N_21285);
nand U26962 (N_26962,N_22555,N_21240);
nand U26963 (N_26963,N_21302,N_23970);
and U26964 (N_26964,N_23964,N_21794);
nand U26965 (N_26965,N_21988,N_23891);
and U26966 (N_26966,N_23661,N_21642);
and U26967 (N_26967,N_23340,N_23889);
nor U26968 (N_26968,N_21923,N_21805);
nand U26969 (N_26969,N_21032,N_23886);
xor U26970 (N_26970,N_23217,N_23703);
xor U26971 (N_26971,N_21424,N_21347);
xor U26972 (N_26972,N_21579,N_23835);
or U26973 (N_26973,N_23434,N_23795);
and U26974 (N_26974,N_21768,N_22340);
xnor U26975 (N_26975,N_22224,N_22187);
xnor U26976 (N_26976,N_22001,N_22265);
nand U26977 (N_26977,N_23138,N_22806);
nor U26978 (N_26978,N_22785,N_23209);
xor U26979 (N_26979,N_21734,N_23643);
xor U26980 (N_26980,N_22662,N_22553);
or U26981 (N_26981,N_22167,N_23648);
nand U26982 (N_26982,N_21727,N_22284);
nor U26983 (N_26983,N_22234,N_23623);
or U26984 (N_26984,N_22532,N_21110);
nor U26985 (N_26985,N_22260,N_21313);
xor U26986 (N_26986,N_22369,N_22154);
and U26987 (N_26987,N_21736,N_21166);
or U26988 (N_26988,N_21781,N_22337);
nand U26989 (N_26989,N_23105,N_22828);
nor U26990 (N_26990,N_21368,N_23261);
nor U26991 (N_26991,N_23380,N_22147);
xor U26992 (N_26992,N_21854,N_23811);
or U26993 (N_26993,N_22976,N_22699);
nor U26994 (N_26994,N_21264,N_23065);
xnor U26995 (N_26995,N_23395,N_23329);
and U26996 (N_26996,N_22657,N_23355);
and U26997 (N_26997,N_22486,N_21841);
and U26998 (N_26998,N_22484,N_21935);
nand U26999 (N_26999,N_22184,N_23459);
and U27000 (N_27000,N_26521,N_26182);
nand U27001 (N_27001,N_24025,N_26365);
xnor U27002 (N_27002,N_25318,N_24811);
nor U27003 (N_27003,N_24817,N_25466);
or U27004 (N_27004,N_24709,N_24832);
nand U27005 (N_27005,N_26671,N_24597);
xnor U27006 (N_27006,N_25601,N_25350);
and U27007 (N_27007,N_26172,N_24496);
and U27008 (N_27008,N_26130,N_25239);
nand U27009 (N_27009,N_24898,N_25749);
or U27010 (N_27010,N_24143,N_24109);
or U27011 (N_27011,N_25739,N_24883);
or U27012 (N_27012,N_24248,N_24341);
and U27013 (N_27013,N_24083,N_24315);
or U27014 (N_27014,N_26886,N_26254);
and U27015 (N_27015,N_26696,N_25583);
or U27016 (N_27016,N_24638,N_26714);
and U27017 (N_27017,N_25002,N_25356);
nor U27018 (N_27018,N_26354,N_26613);
nand U27019 (N_27019,N_25142,N_24673);
or U27020 (N_27020,N_24057,N_24161);
nand U27021 (N_27021,N_25054,N_26245);
nor U27022 (N_27022,N_26732,N_26803);
xor U27023 (N_27023,N_24514,N_26063);
nand U27024 (N_27024,N_26384,N_25953);
or U27025 (N_27025,N_24924,N_25578);
and U27026 (N_27026,N_24054,N_25918);
xnor U27027 (N_27027,N_26769,N_25747);
nor U27028 (N_27028,N_25895,N_26662);
and U27029 (N_27029,N_26726,N_25163);
xor U27030 (N_27030,N_26195,N_25340);
and U27031 (N_27031,N_25378,N_26160);
xor U27032 (N_27032,N_25309,N_26954);
and U27033 (N_27033,N_24798,N_24937);
nor U27034 (N_27034,N_24222,N_25555);
nor U27035 (N_27035,N_26953,N_24228);
nor U27036 (N_27036,N_25347,N_24075);
nor U27037 (N_27037,N_24965,N_25782);
nor U27038 (N_27038,N_25098,N_25812);
xor U27039 (N_27039,N_24157,N_26758);
and U27040 (N_27040,N_24086,N_24050);
and U27041 (N_27041,N_25330,N_25846);
or U27042 (N_27042,N_25716,N_25585);
xor U27043 (N_27043,N_26386,N_26302);
xor U27044 (N_27044,N_26874,N_26528);
and U27045 (N_27045,N_26822,N_24280);
or U27046 (N_27046,N_24327,N_25977);
nor U27047 (N_27047,N_25943,N_25037);
or U27048 (N_27048,N_24993,N_25538);
xor U27049 (N_27049,N_26323,N_26699);
nand U27050 (N_27050,N_25916,N_26913);
nand U27051 (N_27051,N_25489,N_25958);
xor U27052 (N_27052,N_26125,N_24699);
and U27053 (N_27053,N_25638,N_25437);
nor U27054 (N_27054,N_25005,N_25871);
xor U27055 (N_27055,N_24711,N_25307);
nand U27056 (N_27056,N_26153,N_26404);
nor U27057 (N_27057,N_25189,N_26083);
xor U27058 (N_27058,N_26552,N_25912);
or U27059 (N_27059,N_24447,N_25623);
nand U27060 (N_27060,N_25514,N_25324);
or U27061 (N_27061,N_24410,N_24518);
xnor U27062 (N_27062,N_26914,N_26307);
or U27063 (N_27063,N_26562,N_26516);
or U27064 (N_27064,N_25593,N_25435);
or U27065 (N_27065,N_25335,N_25869);
and U27066 (N_27066,N_24038,N_25454);
or U27067 (N_27067,N_26244,N_26347);
and U27068 (N_27068,N_25440,N_26659);
and U27069 (N_27069,N_25104,N_25096);
nor U27070 (N_27070,N_25588,N_26427);
nand U27071 (N_27071,N_24239,N_25751);
xor U27072 (N_27072,N_26867,N_25007);
and U27073 (N_27073,N_24960,N_24353);
xnor U27074 (N_27074,N_26325,N_24111);
or U27075 (N_27075,N_25765,N_24879);
or U27076 (N_27076,N_24464,N_26198);
and U27077 (N_27077,N_25050,N_24918);
or U27078 (N_27078,N_24906,N_25224);
nor U27079 (N_27079,N_24970,N_26898);
or U27080 (N_27080,N_24237,N_24389);
and U27081 (N_27081,N_24819,N_26268);
and U27082 (N_27082,N_25411,N_24933);
nand U27083 (N_27083,N_26443,N_24659);
nand U27084 (N_27084,N_26367,N_26775);
or U27085 (N_27085,N_25471,N_26492);
xor U27086 (N_27086,N_25984,N_24085);
or U27087 (N_27087,N_25463,N_26782);
nand U27088 (N_27088,N_24460,N_24417);
xor U27089 (N_27089,N_26697,N_24227);
nor U27090 (N_27090,N_24837,N_25805);
or U27091 (N_27091,N_24218,N_24403);
or U27092 (N_27092,N_24107,N_25693);
and U27093 (N_27093,N_25785,N_26457);
and U27094 (N_27094,N_26584,N_24116);
nand U27095 (N_27095,N_26747,N_24515);
nand U27096 (N_27096,N_24750,N_24439);
and U27097 (N_27097,N_26567,N_26743);
and U27098 (N_27098,N_26509,N_25205);
nor U27099 (N_27099,N_25906,N_25862);
nand U27100 (N_27100,N_25413,N_25980);
or U27101 (N_27101,N_25140,N_25415);
nor U27102 (N_27102,N_24310,N_25071);
nand U27103 (N_27103,N_26155,N_26936);
nor U27104 (N_27104,N_26080,N_25394);
or U27105 (N_27105,N_24436,N_26771);
xnor U27106 (N_27106,N_25566,N_24755);
or U27107 (N_27107,N_24035,N_25697);
or U27108 (N_27108,N_26685,N_25866);
nor U27109 (N_27109,N_25829,N_26077);
or U27110 (N_27110,N_25879,N_26892);
or U27111 (N_27111,N_25665,N_24060);
nand U27112 (N_27112,N_26770,N_26266);
nand U27113 (N_27113,N_24683,N_26231);
or U27114 (N_27114,N_26833,N_26757);
or U27115 (N_27115,N_26361,N_24513);
nor U27116 (N_27116,N_24211,N_24187);
nor U27117 (N_27117,N_25171,N_25159);
nor U27118 (N_27118,N_26150,N_24047);
xnor U27119 (N_27119,N_26180,N_26494);
nand U27120 (N_27120,N_25049,N_25941);
and U27121 (N_27121,N_26420,N_25883);
and U27122 (N_27122,N_26767,N_24339);
and U27123 (N_27123,N_26890,N_25679);
xnor U27124 (N_27124,N_25882,N_24219);
nand U27125 (N_27125,N_26941,N_24763);
nor U27126 (N_27126,N_26736,N_24619);
xor U27127 (N_27127,N_26927,N_25276);
or U27128 (N_27128,N_25092,N_24781);
nand U27129 (N_27129,N_26860,N_26364);
and U27130 (N_27130,N_25836,N_26107);
nor U27131 (N_27131,N_24984,N_25964);
nor U27132 (N_27132,N_24666,N_25384);
and U27133 (N_27133,N_25312,N_25606);
nor U27134 (N_27134,N_24639,N_25063);
xnor U27135 (N_27135,N_26273,N_24446);
and U27136 (N_27136,N_24968,N_25346);
xnor U27137 (N_27137,N_26006,N_26370);
nor U27138 (N_27138,N_24917,N_24089);
and U27139 (N_27139,N_26911,N_24793);
xnor U27140 (N_27140,N_26491,N_25695);
nand U27141 (N_27141,N_24103,N_24361);
nor U27142 (N_27142,N_24100,N_26353);
nand U27143 (N_27143,N_26709,N_25402);
nor U27144 (N_27144,N_26343,N_26374);
xor U27145 (N_27145,N_24283,N_24556);
nand U27146 (N_27146,N_24426,N_24930);
and U27147 (N_27147,N_26463,N_26460);
or U27148 (N_27148,N_24044,N_24810);
nand U27149 (N_27149,N_26289,N_26147);
and U27150 (N_27150,N_26905,N_26294);
nor U27151 (N_27151,N_26435,N_24608);
nor U27152 (N_27152,N_25420,N_26768);
and U27153 (N_27153,N_25921,N_25886);
and U27154 (N_27154,N_26259,N_24382);
and U27155 (N_27155,N_24370,N_25707);
or U27156 (N_27156,N_25210,N_26549);
nor U27157 (N_27157,N_24764,N_26448);
or U27158 (N_27158,N_25845,N_26336);
xnor U27159 (N_27159,N_25186,N_25719);
xnor U27160 (N_27160,N_25061,N_24486);
xor U27161 (N_27161,N_25209,N_26164);
and U27162 (N_27162,N_24355,N_24000);
xor U27163 (N_27163,N_26242,N_25868);
or U27164 (N_27164,N_26538,N_26828);
or U27165 (N_27165,N_24996,N_24106);
nor U27166 (N_27166,N_25681,N_25784);
nand U27167 (N_27167,N_25951,N_24238);
nor U27168 (N_27168,N_24932,N_26131);
nor U27169 (N_27169,N_26542,N_25678);
and U27170 (N_27170,N_26169,N_24650);
or U27171 (N_27171,N_24234,N_24697);
and U27172 (N_27172,N_26398,N_24138);
or U27173 (N_27173,N_26788,N_24869);
nor U27174 (N_27174,N_26534,N_24196);
nand U27175 (N_27175,N_25341,N_25934);
and U27176 (N_27176,N_24794,N_26235);
or U27177 (N_27177,N_26716,N_24973);
nor U27178 (N_27178,N_24105,N_26526);
nand U27179 (N_27179,N_26895,N_24023);
and U27180 (N_27180,N_25443,N_24149);
nand U27181 (N_27181,N_26002,N_24651);
nand U27182 (N_27182,N_25086,N_26566);
nor U27183 (N_27183,N_25064,N_26744);
xor U27184 (N_27184,N_26215,N_24388);
xor U27185 (N_27185,N_25496,N_25787);
or U27186 (N_27186,N_24309,N_26610);
or U27187 (N_27187,N_26348,N_25295);
nand U27188 (N_27188,N_25745,N_25206);
nand U27189 (N_27189,N_24686,N_24504);
and U27190 (N_27190,N_25746,N_25399);
nor U27191 (N_27191,N_26093,N_24474);
nor U27192 (N_27192,N_26328,N_24304);
nand U27193 (N_27193,N_25563,N_26474);
nand U27194 (N_27194,N_24772,N_25653);
or U27195 (N_27195,N_24600,N_26741);
and U27196 (N_27196,N_26092,N_25148);
or U27197 (N_27197,N_26710,N_26517);
nand U27198 (N_27198,N_26570,N_24243);
nand U27199 (N_27199,N_26986,N_26202);
or U27200 (N_27200,N_26412,N_24451);
nand U27201 (N_27201,N_26520,N_26200);
nand U27202 (N_27202,N_25422,N_26407);
xor U27203 (N_27203,N_24262,N_26020);
nand U27204 (N_27204,N_25861,N_26692);
and U27205 (N_27205,N_24146,N_26156);
or U27206 (N_27206,N_24398,N_25053);
nor U27207 (N_27207,N_26881,N_25664);
nand U27208 (N_27208,N_25303,N_26415);
xor U27209 (N_27209,N_24575,N_26087);
nor U27210 (N_27210,N_26012,N_25521);
or U27211 (N_27211,N_25844,N_26621);
nor U27212 (N_27212,N_24080,N_26228);
xnor U27213 (N_27213,N_24946,N_24661);
or U27214 (N_27214,N_25965,N_25870);
nand U27215 (N_27215,N_24622,N_26438);
xor U27216 (N_27216,N_24311,N_26746);
nor U27217 (N_27217,N_25595,N_26476);
and U27218 (N_27218,N_26322,N_24682);
nor U27219 (N_27219,N_26090,N_26406);
nand U27220 (N_27220,N_24043,N_26535);
xnor U27221 (N_27221,N_25997,N_24266);
nand U27222 (N_27222,N_25961,N_25326);
nand U27223 (N_27223,N_24259,N_25960);
or U27224 (N_27224,N_26992,N_26523);
or U27225 (N_27225,N_24757,N_26192);
and U27226 (N_27226,N_24890,N_26925);
xnor U27227 (N_27227,N_26597,N_25925);
nand U27228 (N_27228,N_26751,N_24002);
xor U27229 (N_27229,N_26078,N_25840);
and U27230 (N_27230,N_26928,N_25445);
and U27231 (N_27231,N_26163,N_26875);
nand U27232 (N_27232,N_24381,N_24990);
and U27233 (N_27233,N_26196,N_25758);
xnor U27234 (N_27234,N_25361,N_24537);
or U27235 (N_27235,N_26296,N_25827);
and U27236 (N_27236,N_25947,N_25207);
and U27237 (N_27237,N_25545,N_24319);
nand U27238 (N_27238,N_24742,N_24145);
and U27239 (N_27239,N_25202,N_24155);
nand U27240 (N_27240,N_24194,N_24843);
or U27241 (N_27241,N_24804,N_25754);
or U27242 (N_27242,N_26065,N_25044);
xor U27243 (N_27243,N_24928,N_26220);
and U27244 (N_27244,N_26880,N_24952);
and U27245 (N_27245,N_26319,N_26606);
nor U27246 (N_27246,N_26991,N_24165);
xnor U27247 (N_27247,N_25258,N_24498);
and U27248 (N_27248,N_25552,N_25806);
nand U27249 (N_27249,N_24466,N_26152);
or U27250 (N_27250,N_26411,N_24885);
and U27251 (N_27251,N_25995,N_26265);
and U27252 (N_27252,N_24118,N_24563);
nor U27253 (N_27253,N_25793,N_26226);
xor U27254 (N_27254,N_24826,N_25817);
xnor U27255 (N_27255,N_25970,N_26035);
nand U27256 (N_27256,N_24292,N_26682);
xnor U27257 (N_27257,N_24156,N_25740);
nand U27258 (N_27258,N_24303,N_26037);
nand U27259 (N_27259,N_26349,N_26816);
nand U27260 (N_27260,N_24765,N_25448);
or U27261 (N_27261,N_25633,N_25717);
xnor U27262 (N_27262,N_26416,N_25062);
nand U27263 (N_27263,N_24391,N_25530);
and U27264 (N_27264,N_24576,N_25856);
or U27265 (N_27265,N_26482,N_25100);
nor U27266 (N_27266,N_26633,N_26135);
nand U27267 (N_27267,N_25558,N_24671);
or U27268 (N_27268,N_26159,N_25987);
nor U27269 (N_27269,N_25501,N_25396);
nor U27270 (N_27270,N_24857,N_24756);
xor U27271 (N_27271,N_26686,N_26238);
or U27272 (N_27272,N_24731,N_24191);
or U27273 (N_27273,N_25926,N_25388);
xnor U27274 (N_27274,N_24335,N_24941);
or U27275 (N_27275,N_25511,N_24245);
nand U27276 (N_27276,N_24703,N_25604);
or U27277 (N_27277,N_26396,N_25284);
or U27278 (N_27278,N_25810,N_25523);
or U27279 (N_27279,N_24349,N_25650);
nand U27280 (N_27280,N_24014,N_24119);
xor U27281 (N_27281,N_25085,N_25973);
xor U27282 (N_27282,N_24380,N_24791);
or U27283 (N_27283,N_25070,N_26924);
nor U27284 (N_27284,N_26944,N_24562);
nand U27285 (N_27285,N_24244,N_25006);
xor U27286 (N_27286,N_25557,N_24359);
or U27287 (N_27287,N_25637,N_26910);
xnor U27288 (N_27288,N_26975,N_24048);
and U27289 (N_27289,N_24484,N_24045);
nor U27290 (N_27290,N_26119,N_26950);
nor U27291 (N_27291,N_25605,N_25509);
nor U27292 (N_27292,N_24774,N_24084);
xnor U27293 (N_27293,N_26047,N_25139);
nand U27294 (N_27294,N_24433,N_25612);
xnor U27295 (N_27295,N_26643,N_26326);
nor U27296 (N_27296,N_26513,N_26074);
xor U27297 (N_27297,N_24599,N_24323);
xor U27298 (N_27298,N_25296,N_26329);
or U27299 (N_27299,N_24795,N_26417);
and U27300 (N_27300,N_25029,N_24573);
or U27301 (N_27301,N_26801,N_25872);
nand U27302 (N_27302,N_25649,N_25451);
xnor U27303 (N_27303,N_24831,N_24269);
or U27304 (N_27304,N_26183,N_25180);
or U27305 (N_27305,N_26837,N_25406);
nand U27306 (N_27306,N_24533,N_26848);
nor U27307 (N_27307,N_26515,N_25654);
nand U27308 (N_27308,N_26978,N_26791);
xor U27309 (N_27309,N_25122,N_25711);
nand U27310 (N_27310,N_26050,N_26399);
or U27311 (N_27311,N_25187,N_26904);
or U27312 (N_27312,N_26702,N_26964);
xnor U27313 (N_27313,N_26749,N_26217);
nor U27314 (N_27314,N_25236,N_26870);
and U27315 (N_27315,N_26461,N_26958);
or U27316 (N_27316,N_25743,N_24108);
or U27317 (N_27317,N_26929,N_25069);
nand U27318 (N_27318,N_25587,N_25516);
nor U27319 (N_27319,N_26304,N_25243);
or U27320 (N_27320,N_26593,N_25648);
nor U27321 (N_27321,N_25502,N_24505);
xnor U27322 (N_27322,N_25319,N_25942);
nand U27323 (N_27323,N_26738,N_26965);
and U27324 (N_27324,N_24724,N_24225);
nor U27325 (N_27325,N_25788,N_25680);
or U27326 (N_27326,N_26730,N_24411);
or U27327 (N_27327,N_26234,N_25288);
or U27328 (N_27328,N_26540,N_25354);
nand U27329 (N_27329,N_24531,N_24298);
and U27330 (N_27330,N_24270,N_25662);
and U27331 (N_27331,N_26634,N_25979);
xor U27332 (N_27332,N_26031,N_24718);
xnor U27333 (N_27333,N_26700,N_26672);
or U27334 (N_27334,N_26920,N_26667);
or U27335 (N_27335,N_25955,N_24099);
xor U27336 (N_27336,N_25216,N_24079);
nand U27337 (N_27337,N_24188,N_24372);
xnor U27338 (N_27338,N_26450,N_26103);
nand U27339 (N_27339,N_24321,N_25204);
nand U27340 (N_27340,N_25500,N_25935);
nor U27341 (N_27341,N_25345,N_25497);
nand U27342 (N_27342,N_26674,N_24307);
and U27343 (N_27343,N_26602,N_26665);
nor U27344 (N_27344,N_25673,N_24594);
nand U27345 (N_27345,N_26088,N_24522);
nor U27346 (N_27346,N_25522,N_24988);
xnor U27347 (N_27347,N_26003,N_24416);
nor U27348 (N_27348,N_24643,N_24549);
nand U27349 (N_27349,N_25657,N_26983);
nand U27350 (N_27350,N_25362,N_25878);
nor U27351 (N_27351,N_25214,N_26514);
and U27352 (N_27352,N_26279,N_26277);
nand U27353 (N_27353,N_25438,N_25718);
or U27354 (N_27354,N_24554,N_25232);
nand U27355 (N_27355,N_24470,N_24092);
or U27356 (N_27356,N_26158,N_26641);
nand U27357 (N_27357,N_25147,N_25000);
and U27358 (N_27358,N_26722,N_25488);
nand U27359 (N_27359,N_26754,N_26127);
nor U27360 (N_27360,N_24740,N_24011);
nand U27361 (N_27361,N_24923,N_24631);
nand U27362 (N_27362,N_26909,N_24265);
nor U27363 (N_27363,N_24552,N_24571);
and U27364 (N_27364,N_25730,N_26419);
nand U27365 (N_27365,N_25093,N_26221);
nand U27366 (N_27366,N_25317,N_26883);
nor U27367 (N_27367,N_26072,N_25778);
nand U27368 (N_27368,N_24500,N_24261);
xor U27369 (N_27369,N_25018,N_24129);
nand U27370 (N_27370,N_26369,N_25565);
and U27371 (N_27371,N_24945,N_24687);
nor U27372 (N_27372,N_25769,N_26434);
xor U27373 (N_27373,N_24713,N_25672);
and U27374 (N_27374,N_25277,N_24076);
nor U27375 (N_27375,N_25339,N_24992);
and U27376 (N_27376,N_26720,N_25626);
nor U27377 (N_27377,N_25423,N_25892);
xor U27378 (N_27378,N_26237,N_25416);
nor U27379 (N_27379,N_26792,N_25141);
nand U27380 (N_27380,N_25548,N_26248);
nand U27381 (N_27381,N_26885,N_25418);
nor U27382 (N_27382,N_26590,N_24935);
nor U27383 (N_27383,N_26500,N_25725);
xor U27384 (N_27384,N_26372,N_25636);
nand U27385 (N_27385,N_26388,N_26132);
and U27386 (N_27386,N_25051,N_26145);
xnor U27387 (N_27387,N_24840,N_25446);
and U27388 (N_27388,N_26436,N_25762);
nor U27389 (N_27389,N_24648,N_24396);
nand U27390 (N_27390,N_25761,N_25904);
nand U27391 (N_27391,N_26267,N_26334);
and U27392 (N_27392,N_24822,N_25518);
nor U27393 (N_27393,N_24275,N_24039);
nand U27394 (N_27394,N_26598,N_24122);
or U27395 (N_27395,N_24178,N_26280);
and U27396 (N_27396,N_26505,N_24636);
nand U27397 (N_27397,N_25683,N_25694);
nor U27398 (N_27398,N_26075,N_25094);
xnor U27399 (N_27399,N_25732,N_25692);
xnor U27400 (N_27400,N_24352,N_25708);
or U27401 (N_27401,N_24434,N_26945);
and U27402 (N_27402,N_24538,N_25696);
or U27403 (N_27403,N_24495,N_26422);
nor U27404 (N_27404,N_26115,N_25483);
and U27405 (N_27405,N_26793,N_26537);
and U27406 (N_27406,N_24963,N_24980);
nand U27407 (N_27407,N_24516,N_26918);
xor U27408 (N_27408,N_26112,N_25222);
or U27409 (N_27409,N_25374,N_26810);
xnor U27410 (N_27410,N_26203,N_24018);
or U27411 (N_27411,N_26844,N_25167);
nand U27412 (N_27412,N_26948,N_24981);
and U27413 (N_27413,N_26232,N_26919);
or U27414 (N_27414,N_26007,N_25381);
and U27415 (N_27415,N_25229,N_25246);
nand U27416 (N_27416,N_25027,N_26647);
nand U27417 (N_27417,N_26016,N_25369);
or U27418 (N_27418,N_26185,N_26009);
or U27419 (N_27419,N_26061,N_25897);
nand U27420 (N_27420,N_26878,N_25447);
or U27421 (N_27421,N_25741,N_26831);
and U27422 (N_27422,N_26798,N_25294);
or U27423 (N_27423,N_24957,N_24870);
nor U27424 (N_27424,N_25410,N_25090);
and U27425 (N_27425,N_26642,N_26687);
or U27426 (N_27426,N_24745,N_26212);
xor U27427 (N_27427,N_24364,N_26177);
and U27428 (N_27428,N_26684,N_26915);
nand U27429 (N_27429,N_25183,N_26197);
or U27430 (N_27430,N_25313,N_24512);
nor U27431 (N_27431,N_26262,N_25311);
xnor U27432 (N_27432,N_25068,N_25770);
xnor U27433 (N_27433,N_25956,N_25109);
nor U27434 (N_27434,N_26376,N_25046);
or U27435 (N_27435,N_24397,N_24069);
and U27436 (N_27436,N_26371,N_24616);
nand U27437 (N_27437,N_24235,N_26990);
xor U27438 (N_27438,N_25195,N_24271);
and U27439 (N_27439,N_26313,N_25475);
or U27440 (N_27440,N_24523,N_26068);
nand U27441 (N_27441,N_24720,N_25969);
nand U27442 (N_27442,N_25155,N_26578);
nand U27443 (N_27443,N_24454,N_26311);
and U27444 (N_27444,N_24019,N_26581);
xor U27445 (N_27445,N_25477,N_25536);
and U27446 (N_27446,N_24342,N_25658);
or U27447 (N_27447,N_25178,N_25596);
xnor U27448 (N_27448,N_26923,N_24291);
xor U27449 (N_27449,N_26022,N_26462);
xor U27450 (N_27450,N_26854,N_24526);
nand U27451 (N_27451,N_25724,N_25080);
xnor U27452 (N_27452,N_26518,N_26790);
xnor U27453 (N_27453,N_26045,N_25848);
or U27454 (N_27454,N_26561,N_26639);
and U27455 (N_27455,N_25173,N_24215);
nand U27456 (N_27456,N_24967,N_24180);
and U27457 (N_27457,N_24406,N_24769);
xor U27458 (N_27458,N_25535,N_25727);
xnor U27459 (N_27459,N_26310,N_24179);
nand U27460 (N_27460,N_26717,N_26243);
and U27461 (N_27461,N_24029,N_26387);
nor U27462 (N_27462,N_26451,N_26309);
nand U27463 (N_27463,N_24889,N_26148);
nand U27464 (N_27464,N_26032,N_24198);
and U27465 (N_27465,N_24739,N_24297);
xor U27466 (N_27466,N_26186,N_25607);
nor U27467 (N_27467,N_25244,N_26171);
or U27468 (N_27468,N_25165,N_26223);
nor U27469 (N_27469,N_26703,N_26737);
nor U27470 (N_27470,N_25397,N_24652);
or U27471 (N_27471,N_24583,N_24233);
nor U27472 (N_27472,N_24231,N_26614);
nor U27473 (N_27473,N_25162,N_25704);
nor U27474 (N_27474,N_24205,N_24334);
or U27475 (N_27475,N_24051,N_25040);
xnor U27476 (N_27476,N_24591,N_26947);
xor U27477 (N_27477,N_25748,N_26413);
and U27478 (N_27478,N_26000,N_26934);
nand U27479 (N_27479,N_26432,N_25677);
nor U27480 (N_27480,N_26644,N_24098);
and U27481 (N_27481,N_26168,N_25081);
xor U27482 (N_27482,N_26230,N_24459);
nand U27483 (N_27483,N_26932,N_26629);
or U27484 (N_27484,N_25651,N_25981);
xnor U27485 (N_27485,N_24839,N_24112);
xor U27486 (N_27486,N_26931,N_25261);
and U27487 (N_27487,N_26539,N_26676);
and U27488 (N_27488,N_25505,N_25110);
and U27489 (N_27489,N_25544,N_25099);
nor U27490 (N_27490,N_26960,N_25851);
xnor U27491 (N_27491,N_26858,N_25512);
and U27492 (N_27492,N_25988,N_24477);
and U27493 (N_27493,N_25486,N_26794);
nand U27494 (N_27494,N_25847,N_24305);
or U27495 (N_27495,N_26467,N_25675);
xnor U27496 (N_27496,N_26143,N_26284);
and U27497 (N_27497,N_26301,N_24488);
or U27498 (N_27498,N_25857,N_25011);
nand U27499 (N_27499,N_24733,N_26058);
or U27500 (N_27500,N_24959,N_25111);
nor U27501 (N_27501,N_25764,N_25661);
nor U27502 (N_27502,N_25305,N_25175);
or U27503 (N_27503,N_24012,N_25986);
nor U27504 (N_27504,N_25275,N_24326);
xnor U27505 (N_27505,N_24910,N_26229);
nand U27506 (N_27506,N_24483,N_24097);
and U27507 (N_27507,N_26625,N_26512);
xor U27508 (N_27508,N_24168,N_26530);
and U27509 (N_27509,N_25083,N_26395);
and U27510 (N_27510,N_26021,N_24159);
and U27511 (N_27511,N_24131,N_24135);
nand U27512 (N_27512,N_25641,N_25299);
xor U27513 (N_27513,N_25469,N_24903);
nand U27514 (N_27514,N_26484,N_24747);
xnor U27515 (N_27515,N_25021,N_24842);
or U27516 (N_27516,N_25811,N_26402);
or U27517 (N_27517,N_26969,N_24418);
or U27518 (N_27518,N_25212,N_26906);
nor U27519 (N_27519,N_25398,N_26627);
nand U27520 (N_27520,N_26646,N_24947);
nand U27521 (N_27521,N_24395,N_26356);
xnor U27522 (N_27522,N_26055,N_25273);
nor U27523 (N_27523,N_24881,N_26366);
and U27524 (N_27524,N_26818,N_24543);
nand U27525 (N_27525,N_25985,N_26465);
or U27526 (N_27526,N_25757,N_24553);
nor U27527 (N_27527,N_24782,N_25170);
and U27528 (N_27528,N_24008,N_25426);
nand U27529 (N_27529,N_26466,N_26678);
nor U27530 (N_27530,N_25101,N_25179);
and U27531 (N_27531,N_25372,N_25867);
xor U27532 (N_27532,N_25079,N_24540);
or U27533 (N_27533,N_26225,N_26239);
nand U27534 (N_27534,N_24295,N_26097);
xnor U27535 (N_27535,N_26557,N_24927);
and U27536 (N_27536,N_24841,N_25794);
xnor U27537 (N_27537,N_26690,N_26585);
and U27538 (N_27538,N_25627,N_25035);
and U27539 (N_27539,N_26497,N_24542);
or U27540 (N_27540,N_25594,N_26760);
or U27541 (N_27541,N_26755,N_26121);
nor U27542 (N_27542,N_24785,N_24662);
nand U27543 (N_27543,N_24414,N_24753);
and U27544 (N_27544,N_25144,N_25994);
xnor U27545 (N_27545,N_26401,N_24654);
and U27546 (N_27546,N_24133,N_24758);
nor U27547 (N_27547,N_24059,N_24982);
xor U27548 (N_27548,N_24121,N_25998);
nor U27549 (N_27549,N_25332,N_24469);
nor U27550 (N_27550,N_26554,N_25789);
xor U27551 (N_27551,N_26630,N_25154);
or U27552 (N_27552,N_24443,N_25854);
xor U27553 (N_27553,N_24400,N_24197);
and U27554 (N_27554,N_26378,N_24030);
nor U27555 (N_27555,N_25834,N_26275);
xnor U27556 (N_27556,N_26891,N_25272);
xor U27557 (N_27557,N_25905,N_24172);
and U27558 (N_27558,N_25527,N_24939);
nor U27559 (N_27559,N_25624,N_24675);
nand U27560 (N_27560,N_25026,N_24005);
nand U27561 (N_27561,N_24536,N_24784);
nor U27562 (N_27562,N_26698,N_26752);
nand U27563 (N_27563,N_26655,N_26901);
or U27564 (N_27564,N_25404,N_25546);
or U27565 (N_27565,N_26711,N_26105);
nand U27566 (N_27566,N_24082,N_25108);
nor U27567 (N_27567,N_26162,N_26489);
and U27568 (N_27568,N_24792,N_25285);
or U27569 (N_27569,N_25771,N_24206);
and U27570 (N_27570,N_25103,N_26385);
nor U27571 (N_27571,N_25449,N_24847);
xor U27572 (N_27572,N_26290,N_24624);
nor U27573 (N_27573,N_26976,N_26252);
nor U27574 (N_27574,N_26297,N_24991);
nand U27575 (N_27575,N_24481,N_25252);
nor U27576 (N_27576,N_25959,N_25371);
xor U27577 (N_27577,N_26175,N_24669);
xor U27578 (N_27578,N_26532,N_25009);
or U27579 (N_27579,N_25982,N_25791);
and U27580 (N_27580,N_24318,N_26247);
xnor U27581 (N_27581,N_25297,N_24192);
nand U27582 (N_27582,N_25218,N_24224);
xnor U27583 (N_27583,N_25666,N_25376);
and U27584 (N_27584,N_24173,N_25571);
nand U27585 (N_27585,N_24871,N_26935);
and U27586 (N_27586,N_26137,N_24592);
or U27587 (N_27587,N_25169,N_25220);
nand U27588 (N_27588,N_25132,N_25830);
and U27589 (N_27589,N_25427,N_25820);
or U27590 (N_27590,N_25260,N_25256);
xor U27591 (N_27591,N_25149,N_24647);
or U27592 (N_27592,N_24344,N_26600);
xor U27593 (N_27593,N_24203,N_26997);
xor U27594 (N_27594,N_25574,N_24095);
and U27595 (N_27595,N_25504,N_24407);
xnor U27596 (N_27596,N_24154,N_25116);
nand U27597 (N_27597,N_25549,N_26638);
xnor U27598 (N_27598,N_26216,N_24028);
nand U27599 (N_27599,N_25391,N_25334);
nor U27600 (N_27600,N_26873,N_26888);
or U27601 (N_27601,N_25620,N_25225);
xnor U27602 (N_27602,N_25266,N_26574);
nor U27603 (N_27603,N_24914,N_24415);
or U27604 (N_27604,N_25822,N_26486);
nand U27605 (N_27605,N_25519,N_26673);
nor U27606 (N_27606,N_24022,N_26649);
or U27607 (N_27607,N_25460,N_26030);
nor U27608 (N_27608,N_25056,N_25153);
and U27609 (N_27609,N_24445,N_25643);
nand U27610 (N_27610,N_24978,N_26456);
nor U27611 (N_27611,N_26314,N_26120);
nor U27612 (N_27612,N_24509,N_26010);
or U27613 (N_27613,N_25901,N_26952);
xor U27614 (N_27614,N_24377,N_25419);
nor U27615 (N_27615,N_26312,N_26013);
and U27616 (N_27616,N_24345,N_26306);
or U27617 (N_27617,N_24830,N_24868);
and U27618 (N_27618,N_26588,N_25876);
nor U27619 (N_27619,N_24853,N_25803);
nand U27620 (N_27620,N_24749,N_24294);
xnor U27621 (N_27621,N_25910,N_26100);
and U27622 (N_27622,N_26863,N_25534);
xor U27623 (N_27623,N_24940,N_24567);
nand U27624 (N_27624,N_24820,N_26802);
nor U27625 (N_27625,N_24767,N_24778);
and U27626 (N_27626,N_24667,N_25242);
nand U27627 (N_27627,N_26332,N_26190);
xnor U27628 (N_27628,N_26067,N_25625);
xor U27629 (N_27629,N_25436,N_24166);
and U27630 (N_27630,N_26827,N_24489);
nor U27631 (N_27631,N_25022,N_26846);
xor U27632 (N_27632,N_24394,N_25373);
or U27633 (N_27633,N_26251,N_25274);
or U27634 (N_27634,N_26921,N_24895);
nand U27635 (N_27635,N_25485,N_26219);
xnor U27636 (N_27636,N_25227,N_24759);
nor U27637 (N_27637,N_26477,N_26531);
or U27638 (N_27638,N_26351,N_24017);
nor U27639 (N_27639,N_25185,N_24453);
xor U27640 (N_27640,N_25136,N_25529);
nand U27641 (N_27641,N_25875,N_24706);
or U27642 (N_27642,N_24821,N_24777);
nor U27643 (N_27643,N_25646,N_24586);
xnor U27644 (N_27644,N_26773,N_26556);
or U27645 (N_27645,N_25893,N_26184);
nor U27646 (N_27646,N_25568,N_24063);
and U27647 (N_27647,N_25949,N_25801);
nor U27648 (N_27648,N_24551,N_25617);
nor U27649 (N_27649,N_24209,N_24340);
and U27650 (N_27650,N_25996,N_25199);
nand U27651 (N_27651,N_25125,N_26141);
nor U27652 (N_27652,N_25674,N_25453);
nor U27653 (N_27653,N_26734,N_24741);
nor U27654 (N_27654,N_25797,N_24401);
or U27655 (N_27655,N_24823,N_24950);
or U27656 (N_27656,N_24510,N_26507);
and U27657 (N_27657,N_25966,N_24534);
and U27658 (N_27658,N_26836,N_26609);
nand U27659 (N_27659,N_24716,N_26612);
and U27660 (N_27660,N_25392,N_24185);
and U27661 (N_27661,N_24413,N_26826);
or U27662 (N_27662,N_25525,N_26039);
nor U27663 (N_27663,N_26719,N_24274);
nand U27664 (N_27664,N_25796,N_25458);
xnor U27665 (N_27665,N_26547,N_26449);
xor U27666 (N_27666,N_26967,N_24824);
nor U27667 (N_27667,N_25603,N_25020);
nand U27668 (N_27668,N_26670,N_26178);
nor U27669 (N_27669,N_24799,N_24578);
xnor U27670 (N_27670,N_24263,N_25405);
nor U27671 (N_27671,N_24998,N_26114);
or U27672 (N_27672,N_25452,N_25036);
or U27673 (N_27673,N_25188,N_26688);
nor U27674 (N_27674,N_25632,N_24809);
xor U27675 (N_27675,N_26519,N_24517);
xnor U27676 (N_27676,N_26081,N_25072);
and U27677 (N_27677,N_24293,N_26291);
xor U27678 (N_27678,N_25450,N_25559);
nor U27679 (N_27679,N_25351,N_24728);
nand U27680 (N_27680,N_24053,N_24128);
nor U27681 (N_27681,N_25386,N_25580);
nor U27682 (N_27682,N_25890,N_24528);
xnor U27683 (N_27683,N_25700,N_24986);
nor U27684 (N_27684,N_25635,N_25031);
or U27685 (N_27685,N_25166,N_25779);
nor U27686 (N_27686,N_24717,N_25656);
xor U27687 (N_27687,N_25268,N_24656);
xor U27688 (N_27688,N_25127,N_26753);
nand U27689 (N_27689,N_26445,N_25896);
nor U27690 (N_27690,N_26756,N_25735);
and U27691 (N_27691,N_26479,N_24290);
nor U27692 (N_27692,N_26795,N_26330);
nand U27693 (N_27693,N_25498,N_24365);
or U27694 (N_27694,N_24272,N_24428);
or U27695 (N_27695,N_26987,N_25048);
nor U27696 (N_27696,N_24289,N_26656);
nand U27697 (N_27697,N_24867,N_24874);
xnor U27698 (N_27698,N_25121,N_25045);
nor U27699 (N_27699,N_25691,N_26740);
xor U27700 (N_27700,N_26057,N_24987);
and U27701 (N_27701,N_24324,N_25531);
and U27702 (N_27702,N_24160,N_24001);
or U27703 (N_27703,N_26408,N_24431);
xor U27704 (N_27704,N_24320,N_26663);
nand U27705 (N_27705,N_26604,N_24424);
xnor U27706 (N_27706,N_26592,N_24351);
xnor U27707 (N_27707,N_25807,N_26999);
nor U27708 (N_27708,N_24626,N_26998);
nor U27709 (N_27709,N_24865,N_26480);
or U27710 (N_27710,N_24557,N_25102);
and U27711 (N_27711,N_24139,N_24693);
xnor U27712 (N_27712,N_25034,N_25510);
nor U27713 (N_27713,N_26544,N_24302);
or U27714 (N_27714,N_24676,N_26204);
or U27715 (N_27715,N_25621,N_24649);
and U27716 (N_27716,N_25366,N_24816);
or U27717 (N_27717,N_24771,N_24333);
nor U27718 (N_27718,N_25097,N_24268);
nor U27719 (N_27719,N_25733,N_25839);
xor U27720 (N_27720,N_25957,N_25157);
and U27721 (N_27721,N_24186,N_26260);
or U27722 (N_27722,N_24169,N_24456);
xor U27723 (N_27723,N_25541,N_24630);
nand U27724 (N_27724,N_24475,N_25032);
nor U27725 (N_27725,N_26724,N_24938);
xnor U27726 (N_27726,N_26073,N_26628);
or U27727 (N_27727,N_25884,N_25265);
or U27728 (N_27728,N_24181,N_25721);
nand U27729 (N_27729,N_24800,N_25263);
or U27730 (N_27730,N_24951,N_26959);
or U27731 (N_27731,N_26423,N_25703);
nor U27732 (N_27732,N_25540,N_24409);
and U27733 (N_27733,N_25368,N_25582);
nor U27734 (N_27734,N_26576,N_26444);
and U27735 (N_27735,N_25331,N_25434);
and U27736 (N_27736,N_24891,N_24152);
xnor U27737 (N_27737,N_25240,N_24752);
nand U27738 (N_27738,N_26640,N_26622);
and U27739 (N_27739,N_24070,N_25755);
nor U27740 (N_27740,N_25015,N_26062);
or U27741 (N_27741,N_25135,N_25182);
xnor U27742 (N_27742,N_25945,N_24301);
xor U27743 (N_27743,N_26817,N_25059);
nand U27744 (N_27744,N_24210,N_24392);
and U27745 (N_27745,N_25439,N_26071);
xnor U27746 (N_27746,N_26912,N_26043);
and U27747 (N_27747,N_24286,N_26551);
xnor U27748 (N_27748,N_26008,N_24478);
or U27749 (N_27749,N_24384,N_26529);
and U27750 (N_27750,N_24876,N_26805);
nor U27751 (N_27751,N_25775,N_26024);
nor U27752 (N_27752,N_26963,N_26096);
nor U27753 (N_27753,N_26321,N_24896);
xor U27754 (N_27754,N_26616,N_26218);
or U27755 (N_27755,N_25281,N_25950);
xnor U27756 (N_27756,N_25219,N_26701);
or U27757 (N_27757,N_24521,N_26721);
nor U27758 (N_27758,N_26582,N_26098);
nor U27759 (N_27759,N_25513,N_25468);
nor U27760 (N_27760,N_24645,N_26654);
xnor U27761 (N_27761,N_24071,N_26027);
nor U27762 (N_27762,N_25480,N_25430);
nor U27763 (N_27763,N_26618,N_24695);
nor U27764 (N_27764,N_26468,N_24285);
nand U27765 (N_27765,N_24976,N_25494);
or U27766 (N_27766,N_25859,N_26804);
nor U27767 (N_27767,N_24267,N_25023);
nand U27768 (N_27768,N_25792,N_24690);
nor U27769 (N_27769,N_24480,N_24972);
nand U27770 (N_27770,N_25198,N_25241);
xor U27771 (N_27771,N_26859,N_26765);
xor U27772 (N_27772,N_24603,N_26144);
and U27773 (N_27773,N_24572,N_25611);
nor U27774 (N_27774,N_24790,N_24748);
or U27775 (N_27775,N_25575,N_25479);
or U27776 (N_27776,N_25134,N_26206);
xor U27777 (N_27777,N_26355,N_24449);
or U27778 (N_27778,N_24174,N_24153);
and U27779 (N_27779,N_24812,N_25891);
or U27780 (N_27780,N_25293,N_26763);
or U27781 (N_27781,N_24455,N_24026);
or U27782 (N_27782,N_25255,N_25992);
nor U27783 (N_27783,N_25482,N_26599);
and U27784 (N_27784,N_26651,N_25639);
nor U27785 (N_27785,N_26586,N_25667);
and U27786 (N_27786,N_25481,N_26926);
nand U27787 (N_27787,N_25302,N_24574);
nand U27788 (N_27788,N_24589,N_24712);
or U27789 (N_27789,N_24467,N_26052);
nor U27790 (N_27790,N_24182,N_24796);
nand U27791 (N_27791,N_24241,N_25168);
and U27792 (N_27792,N_25888,N_24884);
or U27793 (N_27793,N_24465,N_25060);
nand U27794 (N_27794,N_24329,N_24052);
xor U27795 (N_27795,N_25766,N_26205);
nor U27796 (N_27796,N_24633,N_24253);
nand U27797 (N_27797,N_24336,N_26681);
xnor U27798 (N_27798,N_25089,N_26522);
or U27799 (N_27799,N_24126,N_25520);
and U27800 (N_27800,N_25087,N_25767);
and U27801 (N_27801,N_24284,N_25599);
nor U27802 (N_27802,N_26051,N_26036);
nand U27803 (N_27803,N_26624,N_24282);
nor U27804 (N_27804,N_25798,N_25467);
or U27805 (N_27805,N_26056,N_26111);
xor U27806 (N_27806,N_24908,N_25914);
xnor U27807 (N_27807,N_24560,N_26615);
and U27808 (N_27808,N_24958,N_25828);
nor U27809 (N_27809,N_25253,N_26383);
nor U27810 (N_27810,N_25714,N_24694);
and U27811 (N_27811,N_25590,N_26799);
nand U27812 (N_27812,N_24362,N_25944);
and U27813 (N_27813,N_24725,N_25615);
or U27814 (N_27814,N_26089,N_24743);
nand U27815 (N_27815,N_25223,N_24861);
xnor U27816 (N_27816,N_26263,N_26102);
nor U27817 (N_27817,N_25908,N_26424);
nor U27818 (N_27818,N_25713,N_26930);
or U27819 (N_27819,N_26781,N_24246);
or U27820 (N_27820,N_25917,N_26236);
and U27821 (N_27821,N_24461,N_25873);
xor U27822 (N_27822,N_26170,N_26847);
and U27823 (N_27823,N_24566,N_26902);
xnor U27824 (N_27824,N_24077,N_25508);
xor U27825 (N_27825,N_25474,N_26368);
xor U27826 (N_27826,N_24040,N_24199);
or U27827 (N_27827,N_26830,N_26645);
nor U27828 (N_27828,N_24183,N_24037);
and U27829 (N_27829,N_26525,N_24678);
nor U27830 (N_27830,N_24387,N_26723);
xnor U27831 (N_27831,N_25983,N_24499);
or U27832 (N_27832,N_24803,N_24325);
or U27833 (N_27833,N_24031,N_25790);
xnor U27834 (N_27834,N_26862,N_24404);
and U27835 (N_27835,N_26426,N_26117);
or U27836 (N_27836,N_25095,N_24508);
xor U27837 (N_27837,N_26617,N_24707);
nor U27838 (N_27838,N_26094,N_26869);
nand U27839 (N_27839,N_24184,N_24250);
xnor U27840 (N_27840,N_25772,N_26658);
nand U27841 (N_27841,N_26715,N_24042);
nand U27842 (N_27842,N_26745,N_26750);
and U27843 (N_27843,N_26018,N_24366);
or U27844 (N_27844,N_26458,N_26110);
nand U27845 (N_27845,N_24278,N_26026);
or U27846 (N_27846,N_24430,N_25387);
nand U27847 (N_27847,N_25628,N_25816);
or U27848 (N_27848,N_24919,N_24604);
or U27849 (N_27849,N_24921,N_25920);
and U27850 (N_27850,N_25024,N_25150);
xnor U27851 (N_27851,N_26393,N_25010);
nor U27852 (N_27852,N_24328,N_24024);
nand U27853 (N_27853,N_24217,N_26317);
or U27854 (N_27854,N_25191,N_26315);
and U27855 (N_27855,N_26394,N_24264);
xor U27856 (N_27856,N_26974,N_24252);
or U27857 (N_27857,N_24899,N_25235);
and U27858 (N_27858,N_24479,N_26774);
or U27859 (N_27859,N_26136,N_25579);
nand U27860 (N_27860,N_26868,N_25948);
nor U27861 (N_27861,N_24858,N_25184);
nor U27862 (N_27862,N_26034,N_25652);
nand U27863 (N_27863,N_24815,N_26142);
nand U27864 (N_27864,N_26852,N_24171);
nand U27865 (N_27865,N_24120,N_26842);
and U27866 (N_27866,N_25197,N_25619);
nand U27867 (N_27867,N_25939,N_24776);
nand U27868 (N_27868,N_24689,N_24789);
xnor U27869 (N_27869,N_24163,N_24249);
nor U27870 (N_27870,N_26949,N_25357);
nand U27871 (N_27871,N_25181,N_26276);
or U27872 (N_27872,N_24034,N_26452);
or U27873 (N_27873,N_24420,N_25414);
xor U27874 (N_27874,N_24848,N_26637);
nand U27875 (N_27875,N_26359,N_26808);
and U27876 (N_27876,N_24316,N_25234);
or U27877 (N_27877,N_25344,N_24127);
xor U27878 (N_27878,N_24371,N_25462);
or U27879 (N_27879,N_25196,N_25990);
nand U27880 (N_27880,N_26693,N_24356);
xor U27881 (N_27881,N_26759,N_26595);
nand U27882 (N_27882,N_25131,N_25931);
nor U27883 (N_27883,N_24497,N_26392);
nor U27884 (N_27884,N_24090,N_26896);
nor U27885 (N_27885,N_25151,N_26053);
nand U27886 (N_27886,N_25752,N_24701);
xnor U27887 (N_27887,N_24130,N_24061);
nor U27888 (N_27888,N_25401,N_26961);
nor U27889 (N_27889,N_25456,N_25200);
nand U27890 (N_27890,N_25254,N_24956);
nand U27891 (N_27891,N_24602,N_25476);
and U27892 (N_27892,N_26194,N_24732);
xor U27893 (N_27893,N_25271,N_26464);
and U27894 (N_27894,N_25077,N_25390);
nor U27895 (N_27895,N_26129,N_25517);
and U27896 (N_27896,N_24313,N_25348);
nor U27897 (N_27897,N_26181,N_25783);
xnor U27898 (N_27898,N_25137,N_24632);
nand U27899 (N_27899,N_24236,N_26933);
or U27900 (N_27900,N_25922,N_24580);
nor U27901 (N_27901,N_24487,N_24873);
nand U27902 (N_27902,N_24067,N_26779);
nor U27903 (N_27903,N_24618,N_24317);
and U27904 (N_27904,N_24003,N_24123);
xor U27905 (N_27905,N_24705,N_25047);
or U27906 (N_27906,N_24845,N_25278);
and U27907 (N_27907,N_25117,N_26421);
nor U27908 (N_27908,N_26250,N_24658);
nand U27909 (N_27909,N_24989,N_24322);
and U27910 (N_27910,N_26980,N_26337);
nor U27911 (N_27911,N_24520,N_24360);
and U27912 (N_27912,N_25201,N_26069);
or U27913 (N_27913,N_25923,N_25874);
nor U27914 (N_27914,N_24825,N_25631);
nor U27915 (N_27915,N_25598,N_25823);
and U27916 (N_27916,N_24435,N_25470);
nor U27917 (N_27917,N_24550,N_26899);
xor U27918 (N_27918,N_26733,N_26558);
or U27919 (N_27919,N_24113,N_26555);
or U27920 (N_27920,N_26653,N_24375);
xor U27921 (N_27921,N_25759,N_26134);
or U27922 (N_27922,N_24072,N_25589);
or U27923 (N_27923,N_26299,N_24544);
and U27924 (N_27924,N_24468,N_24688);
nand U27925 (N_27925,N_26488,N_24829);
xnor U27926 (N_27926,N_26300,N_25472);
nand U27927 (N_27927,N_24969,N_25245);
xnor U27928 (N_27928,N_25915,N_25858);
nor U27929 (N_27929,N_24585,N_26064);
xnor U27930 (N_27930,N_26320,N_24214);
nand U27931 (N_27931,N_24535,N_25432);
or U27932 (N_27932,N_25999,N_25881);
xor U27933 (N_27933,N_24672,N_24254);
nor U27934 (N_27934,N_26876,N_26727);
and U27935 (N_27935,N_25283,N_26340);
and U27936 (N_27936,N_25660,N_26577);
xor U27937 (N_27937,N_25014,N_24866);
and U27938 (N_27938,N_24802,N_24114);
xnor U27939 (N_27939,N_24134,N_26138);
and U27940 (N_27940,N_25441,N_24836);
and U27941 (N_27941,N_24628,N_25701);
nand U27942 (N_27942,N_26838,N_24399);
or U27943 (N_27943,N_24663,N_26165);
nand U27944 (N_27944,N_26762,N_24354);
and U27945 (N_27945,N_24546,N_26840);
xnor U27946 (N_27946,N_25622,N_25802);
nor U27947 (N_27947,N_25042,N_26545);
nand U27948 (N_27948,N_26042,N_26635);
nand U27949 (N_27949,N_24846,N_26346);
nor U27950 (N_27950,N_25676,N_26493);
or U27951 (N_27951,N_24548,N_26327);
or U27952 (N_27952,N_24229,N_24786);
nand U27953 (N_27953,N_25860,N_25008);
nor U27954 (N_27954,N_24200,N_24004);
or U27955 (N_27955,N_26082,N_26704);
xor U27956 (N_27956,N_26857,N_25455);
nand U27957 (N_27957,N_24117,N_26553);
or U27958 (N_27958,N_26033,N_26298);
or U27959 (N_27959,N_24140,N_24162);
nand U27960 (N_27960,N_24852,N_25709);
nand U27961 (N_27961,N_24911,N_26806);
and U27962 (N_27962,N_24611,N_26360);
xnor U27963 (N_27963,N_25073,N_24887);
and U27964 (N_27964,N_24558,N_24606);
or U27965 (N_27965,N_24593,N_25710);
or U27966 (N_27966,N_26305,N_24442);
nand U27967 (N_27967,N_24358,N_24568);
xor U27968 (N_27968,N_26979,N_26109);
and U27969 (N_27969,N_24856,N_25280);
and U27970 (N_27970,N_25831,N_24452);
or U27971 (N_27971,N_24714,N_26350);
nor U27972 (N_27972,N_25819,N_26409);
nor U27973 (N_27973,N_25821,N_24948);
or U27974 (N_27974,N_26748,N_25543);
xor U27975 (N_27975,N_25290,N_24429);
xnor U27976 (N_27976,N_25591,N_26278);
nor U27977 (N_27977,N_24620,N_25238);
and U27978 (N_27978,N_24068,N_25576);
nor U27979 (N_27979,N_24405,N_24049);
xor U27980 (N_27980,N_25459,N_25630);
nor U27981 (N_27981,N_26040,N_24828);
and U27982 (N_27982,N_26066,N_26777);
xor U27983 (N_27983,N_24491,N_24680);
or U27984 (N_27984,N_24448,N_24954);
nor U27985 (N_27985,N_26139,N_25814);
xor U27986 (N_27986,N_24944,N_26938);
nor U27987 (N_27987,N_24746,N_25375);
nor U27988 (N_27988,N_26707,N_24081);
and U27989 (N_27989,N_24373,N_26224);
nand U27990 (N_27990,N_26428,N_26560);
and U27991 (N_27991,N_24668,N_26882);
nor U27992 (N_27992,N_26571,N_25327);
and U27993 (N_27993,N_24376,N_26695);
nand U27994 (N_27994,N_24378,N_25304);
xor U27995 (N_27995,N_26113,N_25343);
or U27996 (N_27996,N_26855,N_26725);
or U27997 (N_27997,N_24719,N_26023);
and U27998 (N_27998,N_24595,N_25539);
and U27999 (N_27999,N_25644,N_26594);
or U28000 (N_28000,N_24598,N_24877);
or U28001 (N_28001,N_24949,N_24385);
and U28002 (N_28002,N_26391,N_25003);
xnor U28003 (N_28003,N_25659,N_26713);
nor U28004 (N_28004,N_24646,N_26675);
nand U28005 (N_28005,N_24281,N_26099);
nand U28006 (N_28006,N_25924,N_24193);
nand U28007 (N_28007,N_25217,N_24425);
nor U28008 (N_28008,N_24343,N_24681);
or U28009 (N_28009,N_24096,N_26814);
nor U28010 (N_28010,N_26742,N_25705);
nand U28011 (N_28011,N_24036,N_25353);
and U28012 (N_28012,N_25940,N_26981);
nor U28013 (N_28013,N_26258,N_26824);
nand U28014 (N_28014,N_24338,N_26256);
and U28015 (N_28015,N_24170,N_24332);
and U28016 (N_28016,N_26787,N_25286);
and U28017 (N_28017,N_24110,N_25128);
or U28018 (N_28018,N_24337,N_25726);
and U28019 (N_28019,N_26405,N_24189);
and U28020 (N_28020,N_26591,N_26809);
or U28021 (N_28021,N_26563,N_26546);
xnor U28022 (N_28022,N_26333,N_25156);
nand U28023 (N_28023,N_24006,N_24679);
nand U28024 (N_28024,N_26669,N_24124);
xor U28025 (N_28025,N_24213,N_25190);
and U28026 (N_28026,N_25408,N_26689);
and U28027 (N_28027,N_24670,N_25259);
xnor U28028 (N_28028,N_26543,N_24872);
or U28029 (N_28029,N_26587,N_25528);
nand U28030 (N_28030,N_25078,N_25597);
xnor U28031 (N_28031,N_25499,N_24230);
nor U28032 (N_28032,N_26498,N_24850);
nand U28033 (N_28033,N_26176,N_24966);
nor U28034 (N_28034,N_24715,N_24257);
and U28035 (N_28035,N_25389,N_25492);
nand U28036 (N_28036,N_25074,N_26060);
or U28037 (N_28037,N_24859,N_25561);
xnor U28038 (N_28038,N_25382,N_25562);
and U28039 (N_28039,N_26122,N_25610);
and U28040 (N_28040,N_25936,N_24532);
nor U28041 (N_28041,N_26601,N_24961);
nor U28042 (N_28042,N_25832,N_24559);
nand U28043 (N_28043,N_25738,N_26454);
xnor U28044 (N_28044,N_25300,N_26338);
nor U28045 (N_28045,N_26866,N_25194);
nor U28046 (N_28046,N_26104,N_25105);
and U28047 (N_28047,N_26856,N_25907);
nand U28048 (N_28048,N_24314,N_26029);
xor U28049 (N_28049,N_25550,N_24471);
nor U28050 (N_28050,N_24584,N_24955);
and U28051 (N_28051,N_24684,N_24104);
xnor U28052 (N_28052,N_26996,N_25786);
nor U28053 (N_28053,N_26149,N_26257);
or U28054 (N_28054,N_25487,N_24907);
xnor U28055 (N_28055,N_25114,N_26161);
or U28056 (N_28056,N_25130,N_24519);
nand U28057 (N_28057,N_24300,N_24472);
xnor U28058 (N_28058,N_24204,N_25320);
and U28059 (N_28059,N_25655,N_25937);
nand U28060 (N_28060,N_26937,N_26843);
and U28061 (N_28061,N_25971,N_26442);
nand U28062 (N_28062,N_24473,N_26274);
and U28063 (N_28063,N_24931,N_26495);
or U28064 (N_28064,N_26589,N_26879);
and U28065 (N_28065,N_25287,N_24240);
and U28066 (N_28066,N_24506,N_26017);
xnor U28067 (N_28067,N_24610,N_25533);
or U28068 (N_28068,N_24660,N_25004);
and U28069 (N_28069,N_24925,N_26569);
nand U28070 (N_28070,N_25228,N_24312);
and U28071 (N_28071,N_24561,N_25247);
xnor U28072 (N_28072,N_25115,N_24220);
nand U28073 (N_28073,N_26815,N_26207);
nor U28074 (N_28074,N_26533,N_24041);
or U28075 (N_28075,N_24905,N_24368);
nand U28076 (N_28076,N_24288,N_25808);
nand U28077 (N_28077,N_24223,N_24893);
xnor U28078 (N_28078,N_24212,N_25019);
and U28079 (N_28079,N_26303,N_24490);
and U28080 (N_28080,N_24150,N_25138);
xnor U28081 (N_28081,N_26596,N_25403);
and U28082 (N_28082,N_24175,N_25336);
nor U28083 (N_28083,N_25058,N_26541);
nor U28084 (N_28084,N_26028,N_26660);
or U28085 (N_28085,N_24437,N_26173);
nor U28086 (N_28086,N_26812,N_24493);
and U28087 (N_28087,N_26502,N_24524);
nor U28088 (N_28088,N_24094,N_26841);
or U28089 (N_28089,N_26048,N_25055);
or U28090 (N_28090,N_26778,N_26632);
or U28091 (N_28091,N_24078,N_24142);
and U28092 (N_28092,N_25395,N_25645);
nor U28093 (N_28093,N_24920,N_26575);
xor U28094 (N_28094,N_26623,N_24137);
or U28095 (N_28095,N_24144,N_24835);
xor U28096 (N_28096,N_25600,N_26188);
or U28097 (N_28097,N_26128,N_24564);
nor U28098 (N_28098,N_26041,N_24369);
xor U28099 (N_28099,N_25978,N_26970);
nor U28100 (N_28100,N_25123,N_25668);
nor U28101 (N_28101,N_26403,N_25815);
nand U28102 (N_28102,N_26636,N_25226);
nor U28103 (N_28103,N_25231,N_26439);
nand U28104 (N_28104,N_26887,N_25781);
nor U28105 (N_28105,N_25903,N_25991);
or U28106 (N_28106,N_24277,N_26729);
xnor U28107 (N_28107,N_26825,N_25013);
or U28108 (N_28108,N_24346,N_25262);
nor U28109 (N_28109,N_24539,N_24677);
nand U28110 (N_28110,N_26650,N_25355);
or U28111 (N_28111,N_24977,N_26907);
nor U28112 (N_28112,N_24808,N_24596);
nor U28113 (N_28113,N_25584,N_25855);
and U28114 (N_28114,N_24974,N_26764);
or U28115 (N_28115,N_25824,N_24347);
or U28116 (N_28116,N_26187,N_24427);
and U28117 (N_28117,N_25715,N_26786);
and U28118 (N_28118,N_26772,N_26889);
or U28119 (N_28119,N_25756,N_24545);
nor U28120 (N_28120,N_26973,N_26473);
xnor U28121 (N_28121,N_25315,N_26124);
xnor U28122 (N_28122,N_25490,N_24601);
nand U28123 (N_28123,N_24909,N_26179);
or U28124 (N_28124,N_24999,N_25647);
xnor U28125 (N_28125,N_25237,N_26865);
nand U28126 (N_28126,N_26989,N_25799);
nand U28127 (N_28127,N_25421,N_26853);
nand U28128 (N_28128,N_24247,N_24735);
nand U28129 (N_28129,N_26735,N_24141);
and U28130 (N_28130,N_25850,N_25192);
nand U28131 (N_28131,N_26210,N_24612);
and U28132 (N_28132,N_24912,N_26167);
and U28133 (N_28133,N_25152,N_24055);
xnor U28134 (N_28134,N_25269,N_25164);
nor U28135 (N_28135,N_26140,N_24507);
nand U28136 (N_28136,N_24727,N_24046);
or U28137 (N_28137,N_25329,N_24942);
and U28138 (N_28138,N_26510,N_25126);
or U28139 (N_28139,N_25429,N_26157);
nand U28140 (N_28140,N_25577,N_24627);
xor U28141 (N_28141,N_24062,N_24971);
or U28142 (N_28142,N_26440,N_24087);
xor U28143 (N_28143,N_25551,N_24273);
nand U28144 (N_28144,N_24177,N_26708);
nand U28145 (N_28145,N_25989,N_25763);
nor U28146 (N_28146,N_25774,N_25613);
nand U28147 (N_28147,N_26249,N_24306);
xnor U28148 (N_28148,N_24216,N_25424);
nand U28149 (N_28149,N_26679,N_25842);
and U28150 (N_28150,N_24058,N_26903);
nand U28151 (N_28151,N_25292,N_24851);
and U28152 (N_28152,N_25325,N_24444);
or U28153 (N_28153,N_26397,N_25039);
nand U28154 (N_28154,N_24674,N_26657);
or U28155 (N_28155,N_26871,N_26849);
xnor U28156 (N_28156,N_26101,N_26607);
and U28157 (N_28157,N_24875,N_24251);
or U28158 (N_28158,N_25760,N_25208);
and U28159 (N_28159,N_25308,N_25417);
xnor U28160 (N_28160,N_24775,N_26680);
nand U28161 (N_28161,N_24692,N_26499);
nand U28162 (N_28162,N_24013,N_24569);
nand U28163 (N_28163,N_26437,N_24331);
xor U28164 (N_28164,N_25712,N_24773);
nor U28165 (N_28165,N_24207,N_26059);
nor U28166 (N_28166,N_24056,N_24195);
or U28167 (N_28167,N_26985,N_25323);
and U28168 (N_28168,N_25052,N_25560);
nor U28169 (N_28169,N_24348,N_24276);
nor U28170 (N_28170,N_25177,N_26968);
nor U28171 (N_28171,N_26375,N_24125);
and U28172 (N_28172,N_24700,N_24357);
nand U28173 (N_28173,N_24015,N_25670);
and U28174 (N_28174,N_25728,N_24737);
and U28175 (N_28175,N_24350,N_24814);
or U28176 (N_28176,N_26085,N_24744);
or U28177 (N_28177,N_26241,N_26481);
xnor U28178 (N_28178,N_26269,N_24983);
xnor U28179 (N_28179,N_26776,N_24299);
nand U28180 (N_28180,N_26648,N_24788);
or U28181 (N_28181,N_24623,N_25524);
or U28182 (N_28182,N_26485,N_24296);
nor U28183 (N_28183,N_25363,N_25176);
or U28184 (N_28184,N_26894,N_26118);
and U28185 (N_28185,N_24279,N_24863);
or U28186 (N_28186,N_24813,N_26605);
xor U28187 (N_28187,N_24363,N_26019);
xnor U28188 (N_28188,N_26834,N_25075);
and U28189 (N_28189,N_24844,N_25929);
xnor U28190 (N_28190,N_26731,N_24021);
and U28191 (N_28191,N_24393,N_26946);
and U28192 (N_28192,N_26381,N_25592);
nor U28193 (N_28193,N_24590,N_24621);
or U28194 (N_28194,N_25493,N_24221);
or U28195 (N_28195,N_24412,N_26829);
nand U28196 (N_28196,N_24704,N_25919);
or U28197 (N_28197,N_25968,N_24308);
or U28198 (N_28198,N_26316,N_26951);
nor U28199 (N_28199,N_25065,N_24202);
or U28200 (N_28200,N_25723,N_25572);
xor U28201 (N_28201,N_24698,N_26293);
nor U28202 (N_28202,N_25737,N_26966);
and U28203 (N_28203,N_26046,N_25001);
and U28204 (N_28204,N_26116,N_24797);
and U28205 (N_28205,N_26766,N_25473);
nor U28206 (N_28206,N_24582,N_26893);
and U28207 (N_28207,N_26335,N_26559);
or U28208 (N_28208,N_25671,N_26797);
and U28209 (N_28209,N_25143,N_26453);
and U28210 (N_28210,N_25129,N_26780);
and U28211 (N_28211,N_26796,N_25569);
xor U28212 (N_28212,N_25547,N_26583);
nand U28213 (N_28213,N_25289,N_25425);
xor U28214 (N_28214,N_26993,N_25902);
and U28215 (N_28215,N_26821,N_24330);
xnor U28216 (N_28216,N_24779,N_25400);
nand U28217 (N_28217,N_24787,N_26015);
or U28218 (N_28218,N_26292,N_25119);
or U28219 (N_28219,N_26151,N_26811);
or U28220 (N_28220,N_24833,N_24482);
nor U28221 (N_28221,N_25457,N_24091);
or U28222 (N_28222,N_25889,N_26342);
nand U28223 (N_28223,N_25484,N_24527);
nand U28224 (N_28224,N_26652,N_26418);
nor U28225 (N_28225,N_25251,N_24570);
xnor U28226 (N_28226,N_26884,N_24501);
and U28227 (N_28227,N_24886,N_25193);
and U28228 (N_28228,N_25385,N_25809);
xnor U28229 (N_28229,N_25952,N_26705);
nor U28230 (N_28230,N_25753,N_24115);
xnor U28231 (N_28231,N_24201,N_25301);
and U28232 (N_28232,N_25172,N_25702);
or U28233 (N_28233,N_26380,N_26739);
or U28234 (N_28234,N_25233,N_24943);
nor U28235 (N_28235,N_24033,N_26784);
and U28236 (N_28236,N_26511,N_25352);
nor U28237 (N_28237,N_25379,N_24132);
nor U28238 (N_28238,N_26783,N_25088);
and U28239 (N_28239,N_26850,N_24419);
xor U28240 (N_28240,N_25322,N_25082);
xnor U28241 (N_28241,N_24888,N_24783);
or U28242 (N_28242,N_24073,N_26459);
nor U28243 (N_28243,N_24642,N_24088);
and U28244 (N_28244,N_26957,N_25461);
nand U28245 (N_28245,N_26166,N_25409);
or U28246 (N_28246,N_25107,N_24581);
xor U28247 (N_28247,N_26564,N_24422);
xor U28248 (N_28248,N_24738,N_24768);
or U28249 (N_28249,N_25669,N_26800);
or U28250 (N_28250,N_26414,N_24151);
xor U28251 (N_28251,N_25298,N_26382);
and U28252 (N_28252,N_24962,N_25124);
or U28253 (N_28253,N_25359,N_24730);
nor U28254 (N_28254,N_24256,N_25976);
or U28255 (N_28255,N_26939,N_25804);
or U28256 (N_28256,N_26281,N_24805);
or U28257 (N_28257,N_24101,N_26095);
nor U28258 (N_28258,N_26014,N_24929);
xor U28259 (N_28259,N_26483,N_25750);
and U28260 (N_28260,N_26271,N_25412);
and U28261 (N_28261,N_24766,N_26084);
or U28262 (N_28262,N_24754,N_24644);
xnor U28263 (N_28263,N_24164,N_25328);
or U28264 (N_28264,N_24605,N_25618);
and U28265 (N_28265,N_26282,N_26339);
xor U28266 (N_28266,N_24440,N_25818);
and U28267 (N_28267,N_24985,N_25564);
or U28268 (N_28268,N_26174,N_25795);
nor U28269 (N_28269,N_25038,N_26318);
nor U28270 (N_28270,N_26988,N_25927);
or U28271 (N_28271,N_24136,N_26146);
xor U28272 (N_28272,N_24147,N_25640);
xnor U28273 (N_28273,N_26661,N_25698);
xor U28274 (N_28274,N_26255,N_25174);
nor U28275 (N_28275,N_24226,N_24995);
nor U28276 (N_28276,N_26611,N_26568);
nor U28277 (N_28277,N_24390,N_26940);
nand U28278 (N_28278,N_25899,N_24864);
and U28279 (N_28279,N_26785,N_25573);
and U28280 (N_28280,N_25043,N_24936);
nand U28281 (N_28281,N_24032,N_24547);
nand U28282 (N_28282,N_26789,N_26133);
and U28283 (N_28283,N_26536,N_24635);
nand U28284 (N_28284,N_24020,N_25067);
nand U28285 (N_28285,N_25554,N_24208);
xor U28286 (N_28286,N_26324,N_24242);
nor U28287 (N_28287,N_26608,N_26331);
nand U28288 (N_28288,N_25913,N_24441);
nand U28289 (N_28289,N_25690,N_25358);
nand U28290 (N_28290,N_26579,N_24934);
and U28291 (N_28291,N_25491,N_25776);
xnor U28292 (N_28292,N_25744,N_25773);
and U28293 (N_28293,N_25158,N_24637);
xnor U28294 (N_28294,N_26864,N_26839);
or U28295 (N_28295,N_25687,N_26209);
or U28296 (N_28296,N_25974,N_26001);
or U28297 (N_28297,N_25465,N_26213);
or U28298 (N_28298,N_26877,N_24463);
and U28299 (N_28299,N_25249,N_26038);
nand U28300 (N_28300,N_26345,N_24074);
nand U28301 (N_28301,N_24402,N_24502);
and U28302 (N_28302,N_26631,N_24458);
or U28303 (N_28303,N_24258,N_24827);
xor U28304 (N_28304,N_24374,N_24421);
xnor U28305 (N_28305,N_26995,N_25431);
and U28306 (N_28306,N_26712,N_24780);
xnor U28307 (N_28307,N_24176,N_25837);
nor U28308 (N_28308,N_26049,N_25076);
and U28309 (N_28309,N_25734,N_24565);
nor U28310 (N_28310,N_26942,N_26668);
nor U28311 (N_28311,N_24462,N_25629);
or U28312 (N_28312,N_26288,N_26718);
nor U28313 (N_28313,N_26005,N_24625);
or U28314 (N_28314,N_24016,N_24190);
nor U28315 (N_28315,N_26189,N_26472);
nor U28316 (N_28316,N_26264,N_25933);
nand U28317 (N_28317,N_25203,N_25975);
nand U28318 (N_28318,N_25865,N_24530);
nand U28319 (N_28319,N_24708,N_25291);
nor U28320 (N_28320,N_24696,N_25777);
or U28321 (N_28321,N_26358,N_24255);
or U28322 (N_28322,N_26283,N_24892);
xor U28323 (N_28323,N_24964,N_26478);
or U28324 (N_28324,N_24629,N_25030);
nand U28325 (N_28325,N_25506,N_24997);
nand U28326 (N_28326,N_26079,N_25911);
xor U28327 (N_28327,N_26728,N_26845);
nor U28328 (N_28328,N_25282,N_25257);
xor U28329 (N_28329,N_24367,N_25113);
xor U28330 (N_28330,N_26246,N_26490);
nand U28331 (N_28331,N_24655,N_24379);
nor U28332 (N_28332,N_24457,N_25849);
and U28333 (N_28333,N_26580,N_26897);
nor U28334 (N_28334,N_26565,N_26972);
nor U28335 (N_28335,N_26285,N_25215);
nand U28336 (N_28336,N_24710,N_25863);
and U28337 (N_28337,N_24862,N_24615);
nand U28338 (N_28338,N_26524,N_24664);
nand U28339 (N_28339,N_25133,N_25887);
xnor U28340 (N_28340,N_26916,N_26011);
xnor U28341 (N_28341,N_25383,N_25800);
xor U28342 (N_28342,N_25091,N_24691);
or U28343 (N_28343,N_26548,N_26508);
nor U28344 (N_28344,N_26379,N_25729);
nor U28345 (N_28345,N_25894,N_25442);
nand U28346 (N_28346,N_25542,N_26691);
xor U28347 (N_28347,N_24726,N_24609);
xnor U28348 (N_28348,N_26253,N_25706);
and U28349 (N_28349,N_25967,N_24723);
xnor U28350 (N_28350,N_24167,N_24102);
nand U28351 (N_28351,N_26835,N_26977);
xor U28352 (N_28352,N_24702,N_24607);
or U28353 (N_28353,N_26761,N_25365);
and U28354 (N_28354,N_26455,N_25360);
nor U28355 (N_28355,N_26429,N_25634);
nor U28356 (N_28356,N_26984,N_24761);
xor U28357 (N_28357,N_25310,N_26341);
xor U28358 (N_28358,N_24975,N_24897);
or U28359 (N_28359,N_26076,N_26086);
or U28360 (N_28360,N_24904,N_25066);
nor U28361 (N_28361,N_25833,N_25364);
nor U28362 (N_28362,N_24855,N_24492);
nand U28363 (N_28363,N_26362,N_25145);
nand U28364 (N_28364,N_25731,N_26308);
or U28365 (N_28365,N_25146,N_25267);
xnor U28366 (N_28366,N_24913,N_24009);
and U28367 (N_28367,N_26287,N_26199);
and U28368 (N_28368,N_26227,N_25663);
and U28369 (N_28369,N_26193,N_24880);
nor U28370 (N_28370,N_25841,N_26475);
nand U28371 (N_28371,N_24736,N_26431);
nor U28372 (N_28372,N_25342,N_24665);
and U28373 (N_28373,N_25780,N_25016);
nand U28374 (N_28374,N_26025,N_25684);
nand U28375 (N_28375,N_25688,N_26861);
xnor U28376 (N_28376,N_25614,N_26389);
or U28377 (N_28377,N_24423,N_25722);
and U28378 (N_28378,N_26447,N_24882);
or U28379 (N_28379,N_24751,N_26823);
or U28380 (N_28380,N_25852,N_25478);
and U28381 (N_28381,N_24408,N_24386);
nand U28382 (N_28382,N_26820,N_26851);
and U28383 (N_28383,N_26487,N_24587);
xnor U28384 (N_28384,N_24525,N_24614);
xnor U28385 (N_28385,N_26214,N_25826);
xnor U28386 (N_28386,N_24232,N_26956);
nor U28387 (N_28387,N_25349,N_26446);
or U28388 (N_28388,N_25699,N_25084);
xor U28389 (N_28389,N_26666,N_25930);
nor U28390 (N_28390,N_25581,N_25321);
xnor U28391 (N_28391,N_24849,N_25537);
nor U28392 (N_28392,N_25507,N_26240);
xnor U28393 (N_28393,N_25853,N_24953);
nor U28394 (N_28394,N_26222,N_24287);
xnor U28395 (N_28395,N_24900,N_26400);
nand U28396 (N_28396,N_26208,N_26373);
nor U28397 (N_28397,N_26982,N_24450);
and U28398 (N_28398,N_24729,N_25993);
nand U28399 (N_28399,N_25428,N_26430);
nand U28400 (N_28400,N_25264,N_25028);
xor U28401 (N_28401,N_24979,N_24577);
or U28402 (N_28402,N_24721,N_25306);
or U28403 (N_28403,N_26664,N_26357);
nor U28404 (N_28404,N_24915,N_25407);
and U28405 (N_28405,N_24657,N_26677);
or U28406 (N_28406,N_24007,N_26819);
or U28407 (N_28407,N_24734,N_24994);
xor U28408 (N_28408,N_26154,N_24383);
or U28409 (N_28409,N_26191,N_25025);
nand U28410 (N_28410,N_26572,N_26619);
xnor U28411 (N_28411,N_24818,N_26433);
nor U28412 (N_28412,N_26471,N_25041);
and U28413 (N_28413,N_26123,N_25954);
or U28414 (N_28414,N_25864,N_25567);
and U28415 (N_28415,N_25686,N_24640);
xor U28416 (N_28416,N_26344,N_24916);
and U28417 (N_28417,N_25057,N_25120);
and U28418 (N_28418,N_26900,N_24838);
nand U28419 (N_28419,N_24093,N_25972);
xnor U28420 (N_28420,N_24066,N_24260);
or U28421 (N_28421,N_26469,N_26054);
nand U28422 (N_28422,N_25877,N_26044);
xnor U28423 (N_28423,N_25248,N_24894);
nand U28424 (N_28424,N_26813,N_24438);
or U28425 (N_28425,N_25314,N_25720);
and U28426 (N_28426,N_26233,N_26363);
nand U28427 (N_28427,N_25843,N_26917);
or U28428 (N_28428,N_25556,N_25825);
xnor U28429 (N_28429,N_24922,N_24613);
or U28430 (N_28430,N_26261,N_26603);
or U28431 (N_28431,N_24065,N_25526);
xor U28432 (N_28432,N_26270,N_25161);
xor U28433 (N_28433,N_26106,N_24806);
xnor U28434 (N_28434,N_26108,N_24926);
nand U28435 (N_28435,N_25367,N_25112);
nand U28436 (N_28436,N_25532,N_26626);
or U28437 (N_28437,N_26441,N_24770);
nand U28438 (N_28438,N_25768,N_26872);
nor U28439 (N_28439,N_26295,N_26352);
nand U28440 (N_28440,N_26377,N_25393);
nor U28441 (N_28441,N_25270,N_26683);
or U28442 (N_28442,N_26908,N_25742);
nor U28443 (N_28443,N_25885,N_24641);
nand U28444 (N_28444,N_24064,N_26832);
xnor U28445 (N_28445,N_25685,N_26390);
nor U28446 (N_28446,N_25900,N_25503);
nor U28447 (N_28447,N_26272,N_25963);
nor U28448 (N_28448,N_24588,N_26527);
nand U28449 (N_28449,N_25946,N_25602);
xnor U28450 (N_28450,N_24555,N_25616);
or U28451 (N_28451,N_24432,N_26004);
nand U28452 (N_28452,N_24541,N_26470);
nor U28453 (N_28453,N_25279,N_25642);
or U28454 (N_28454,N_26994,N_25962);
nand U28455 (N_28455,N_25570,N_26694);
and U28456 (N_28456,N_24878,N_25835);
xnor U28457 (N_28457,N_26550,N_25813);
nor U28458 (N_28458,N_26620,N_26425);
nand U28459 (N_28459,N_25250,N_25689);
and U28460 (N_28460,N_24854,N_25838);
or U28461 (N_28461,N_25433,N_25444);
xor U28462 (N_28462,N_24511,N_26503);
and U28463 (N_28463,N_25736,N_25221);
or U28464 (N_28464,N_24503,N_26955);
nor U28465 (N_28465,N_24807,N_24158);
and U28466 (N_28466,N_26501,N_26943);
nand U28467 (N_28467,N_24653,N_25586);
or U28468 (N_28468,N_25230,N_26506);
xor U28469 (N_28469,N_25106,N_24494);
nand U28470 (N_28470,N_24010,N_26286);
or U28471 (N_28471,N_25012,N_25928);
and U28472 (N_28472,N_26573,N_25938);
nand U28473 (N_28473,N_26971,N_25333);
nor U28474 (N_28474,N_25033,N_25608);
nand U28475 (N_28475,N_26410,N_26504);
or U28476 (N_28476,N_24801,N_25609);
and U28477 (N_28477,N_24901,N_25213);
xor U28478 (N_28478,N_24722,N_25017);
xnor U28479 (N_28479,N_24148,N_25880);
nor U28480 (N_28480,N_25932,N_24762);
and U28481 (N_28481,N_24760,N_26706);
xnor U28482 (N_28482,N_24860,N_24476);
nand U28483 (N_28483,N_25898,N_25909);
and U28484 (N_28484,N_24027,N_24485);
nand U28485 (N_28485,N_25211,N_25515);
nand U28486 (N_28486,N_25370,N_24617);
and U28487 (N_28487,N_25337,N_24634);
nand U28488 (N_28488,N_25380,N_26496);
and U28489 (N_28489,N_26201,N_26962);
and U28490 (N_28490,N_26126,N_24529);
nand U28491 (N_28491,N_25553,N_25377);
nand U28492 (N_28492,N_26922,N_24685);
nor U28493 (N_28493,N_24902,N_26091);
nand U28494 (N_28494,N_24834,N_25316);
or U28495 (N_28495,N_25118,N_25682);
or U28496 (N_28496,N_25338,N_25464);
nand U28497 (N_28497,N_25495,N_26807);
xnor U28498 (N_28498,N_25160,N_24579);
xor U28499 (N_28499,N_26070,N_26211);
or U28500 (N_28500,N_24023,N_26461);
and U28501 (N_28501,N_26773,N_26108);
nor U28502 (N_28502,N_25028,N_25807);
nor U28503 (N_28503,N_25200,N_25730);
nand U28504 (N_28504,N_24656,N_26089);
or U28505 (N_28505,N_24099,N_26671);
nand U28506 (N_28506,N_26420,N_26872);
and U28507 (N_28507,N_25956,N_25718);
or U28508 (N_28508,N_25083,N_25043);
and U28509 (N_28509,N_24602,N_24842);
or U28510 (N_28510,N_25069,N_26055);
nor U28511 (N_28511,N_26028,N_24848);
and U28512 (N_28512,N_25219,N_24425);
xor U28513 (N_28513,N_24047,N_26321);
xnor U28514 (N_28514,N_24414,N_26842);
nand U28515 (N_28515,N_26803,N_24469);
and U28516 (N_28516,N_24311,N_26150);
xnor U28517 (N_28517,N_24292,N_25918);
nand U28518 (N_28518,N_24578,N_26469);
or U28519 (N_28519,N_24449,N_26583);
or U28520 (N_28520,N_24451,N_24987);
or U28521 (N_28521,N_26355,N_25165);
nand U28522 (N_28522,N_26545,N_24006);
or U28523 (N_28523,N_25666,N_25713);
xnor U28524 (N_28524,N_25257,N_24523);
nor U28525 (N_28525,N_25052,N_26951);
xnor U28526 (N_28526,N_24867,N_26174);
nand U28527 (N_28527,N_26415,N_26613);
nand U28528 (N_28528,N_25473,N_26313);
or U28529 (N_28529,N_25521,N_26440);
or U28530 (N_28530,N_26285,N_26749);
and U28531 (N_28531,N_25586,N_24773);
xor U28532 (N_28532,N_24289,N_25964);
xor U28533 (N_28533,N_25682,N_24625);
nand U28534 (N_28534,N_26310,N_24840);
or U28535 (N_28535,N_26220,N_24551);
xnor U28536 (N_28536,N_24230,N_24690);
nor U28537 (N_28537,N_26108,N_26772);
and U28538 (N_28538,N_26841,N_25893);
or U28539 (N_28539,N_26833,N_25716);
nand U28540 (N_28540,N_25747,N_26134);
or U28541 (N_28541,N_25793,N_25736);
xor U28542 (N_28542,N_24724,N_24900);
xor U28543 (N_28543,N_26043,N_24877);
or U28544 (N_28544,N_25930,N_26612);
nand U28545 (N_28545,N_25877,N_24578);
nor U28546 (N_28546,N_26346,N_25290);
or U28547 (N_28547,N_26685,N_25761);
nor U28548 (N_28548,N_26234,N_24367);
nand U28549 (N_28549,N_24081,N_24180);
or U28550 (N_28550,N_26752,N_25733);
nor U28551 (N_28551,N_24848,N_24946);
xnor U28552 (N_28552,N_26560,N_25620);
and U28553 (N_28553,N_24903,N_26810);
and U28554 (N_28554,N_24554,N_24102);
or U28555 (N_28555,N_24646,N_24554);
nand U28556 (N_28556,N_25884,N_25167);
or U28557 (N_28557,N_24686,N_24195);
xor U28558 (N_28558,N_26596,N_26791);
and U28559 (N_28559,N_24426,N_25030);
or U28560 (N_28560,N_24140,N_24604);
nand U28561 (N_28561,N_25394,N_25221);
or U28562 (N_28562,N_25236,N_24274);
nand U28563 (N_28563,N_26169,N_25690);
nor U28564 (N_28564,N_26120,N_24572);
nand U28565 (N_28565,N_26801,N_26557);
nor U28566 (N_28566,N_25198,N_26177);
nand U28567 (N_28567,N_26630,N_26264);
and U28568 (N_28568,N_26779,N_24762);
nand U28569 (N_28569,N_26286,N_26477);
xor U28570 (N_28570,N_24408,N_24699);
xnor U28571 (N_28571,N_24162,N_25720);
xor U28572 (N_28572,N_26693,N_26542);
nand U28573 (N_28573,N_25844,N_26568);
xnor U28574 (N_28574,N_24915,N_26819);
nand U28575 (N_28575,N_24055,N_25552);
and U28576 (N_28576,N_25246,N_24783);
nor U28577 (N_28577,N_25949,N_24097);
nand U28578 (N_28578,N_26025,N_26845);
xnor U28579 (N_28579,N_25067,N_26519);
nor U28580 (N_28580,N_25610,N_26428);
nor U28581 (N_28581,N_25201,N_26333);
nor U28582 (N_28582,N_26874,N_24096);
nand U28583 (N_28583,N_25721,N_26683);
nor U28584 (N_28584,N_26363,N_25646);
nor U28585 (N_28585,N_24580,N_25703);
and U28586 (N_28586,N_24721,N_24876);
and U28587 (N_28587,N_25443,N_25826);
nand U28588 (N_28588,N_26972,N_24294);
nand U28589 (N_28589,N_24560,N_24107);
or U28590 (N_28590,N_26723,N_25133);
nand U28591 (N_28591,N_24791,N_25955);
nand U28592 (N_28592,N_25831,N_25481);
xor U28593 (N_28593,N_24540,N_24468);
or U28594 (N_28594,N_25005,N_26330);
and U28595 (N_28595,N_25885,N_26199);
nor U28596 (N_28596,N_25390,N_24086);
and U28597 (N_28597,N_26530,N_24271);
and U28598 (N_28598,N_26878,N_26058);
nor U28599 (N_28599,N_26816,N_25217);
and U28600 (N_28600,N_24549,N_24025);
and U28601 (N_28601,N_26088,N_26482);
and U28602 (N_28602,N_26960,N_24109);
nor U28603 (N_28603,N_24388,N_24670);
nand U28604 (N_28604,N_26712,N_24239);
nor U28605 (N_28605,N_25762,N_25552);
xor U28606 (N_28606,N_25539,N_24230);
and U28607 (N_28607,N_26527,N_25885);
xor U28608 (N_28608,N_25860,N_25527);
nand U28609 (N_28609,N_26624,N_25838);
xor U28610 (N_28610,N_26284,N_26414);
or U28611 (N_28611,N_25583,N_26957);
xor U28612 (N_28612,N_24530,N_26227);
xor U28613 (N_28613,N_24982,N_26368);
xor U28614 (N_28614,N_25607,N_24705);
or U28615 (N_28615,N_25087,N_24607);
or U28616 (N_28616,N_24379,N_25323);
nor U28617 (N_28617,N_25845,N_24094);
nor U28618 (N_28618,N_24823,N_25860);
xnor U28619 (N_28619,N_26460,N_26679);
nand U28620 (N_28620,N_25597,N_26705);
and U28621 (N_28621,N_26229,N_24506);
xnor U28622 (N_28622,N_26971,N_25472);
nor U28623 (N_28623,N_25007,N_24187);
or U28624 (N_28624,N_24979,N_25945);
or U28625 (N_28625,N_26413,N_25041);
or U28626 (N_28626,N_25874,N_25005);
xor U28627 (N_28627,N_25813,N_24948);
nor U28628 (N_28628,N_24347,N_26588);
nor U28629 (N_28629,N_24103,N_24018);
and U28630 (N_28630,N_25547,N_25912);
xnor U28631 (N_28631,N_26096,N_24521);
or U28632 (N_28632,N_24928,N_26217);
nand U28633 (N_28633,N_25259,N_24037);
and U28634 (N_28634,N_25695,N_24239);
or U28635 (N_28635,N_26695,N_24312);
or U28636 (N_28636,N_25350,N_24956);
xor U28637 (N_28637,N_26220,N_24729);
nand U28638 (N_28638,N_24989,N_25952);
or U28639 (N_28639,N_26423,N_26999);
or U28640 (N_28640,N_24423,N_24180);
xnor U28641 (N_28641,N_24042,N_26464);
or U28642 (N_28642,N_25659,N_24902);
or U28643 (N_28643,N_26043,N_24783);
nand U28644 (N_28644,N_26463,N_25358);
or U28645 (N_28645,N_26487,N_25780);
xnor U28646 (N_28646,N_25202,N_25937);
and U28647 (N_28647,N_26834,N_24240);
and U28648 (N_28648,N_25668,N_25210);
and U28649 (N_28649,N_25195,N_25064);
xor U28650 (N_28650,N_26954,N_26117);
nor U28651 (N_28651,N_25818,N_25220);
and U28652 (N_28652,N_24502,N_26116);
or U28653 (N_28653,N_26278,N_26208);
xor U28654 (N_28654,N_26121,N_24863);
and U28655 (N_28655,N_26595,N_25476);
and U28656 (N_28656,N_24619,N_24345);
nor U28657 (N_28657,N_26525,N_25994);
nor U28658 (N_28658,N_24151,N_25245);
and U28659 (N_28659,N_24314,N_25537);
nand U28660 (N_28660,N_24563,N_25159);
nand U28661 (N_28661,N_24436,N_25218);
and U28662 (N_28662,N_24145,N_25555);
nand U28663 (N_28663,N_24216,N_26628);
nor U28664 (N_28664,N_25708,N_24859);
and U28665 (N_28665,N_26896,N_24441);
or U28666 (N_28666,N_26103,N_26278);
or U28667 (N_28667,N_26039,N_26206);
or U28668 (N_28668,N_25929,N_24342);
xnor U28669 (N_28669,N_25630,N_24736);
and U28670 (N_28670,N_26032,N_25540);
or U28671 (N_28671,N_25192,N_25469);
or U28672 (N_28672,N_24087,N_26376);
nor U28673 (N_28673,N_25565,N_26851);
or U28674 (N_28674,N_26446,N_25834);
or U28675 (N_28675,N_24194,N_26358);
nand U28676 (N_28676,N_26515,N_24124);
nand U28677 (N_28677,N_26873,N_26656);
or U28678 (N_28678,N_26521,N_26033);
nor U28679 (N_28679,N_25123,N_25688);
or U28680 (N_28680,N_24672,N_25587);
xor U28681 (N_28681,N_24638,N_26559);
and U28682 (N_28682,N_25969,N_26941);
xor U28683 (N_28683,N_25798,N_26094);
and U28684 (N_28684,N_26983,N_24970);
xnor U28685 (N_28685,N_26880,N_24922);
or U28686 (N_28686,N_24573,N_25880);
or U28687 (N_28687,N_24648,N_24694);
nand U28688 (N_28688,N_24770,N_26836);
nand U28689 (N_28689,N_24170,N_26835);
nand U28690 (N_28690,N_24070,N_25890);
and U28691 (N_28691,N_26394,N_24419);
xnor U28692 (N_28692,N_26066,N_25050);
and U28693 (N_28693,N_24188,N_26457);
nand U28694 (N_28694,N_26928,N_24499);
nor U28695 (N_28695,N_25335,N_25016);
nor U28696 (N_28696,N_25152,N_26395);
xor U28697 (N_28697,N_24301,N_24318);
nand U28698 (N_28698,N_26451,N_25350);
and U28699 (N_28699,N_24553,N_26288);
nor U28700 (N_28700,N_25439,N_25504);
and U28701 (N_28701,N_24214,N_25382);
nand U28702 (N_28702,N_25389,N_26815);
nor U28703 (N_28703,N_25331,N_24218);
nor U28704 (N_28704,N_26514,N_26701);
xnor U28705 (N_28705,N_24234,N_26634);
nand U28706 (N_28706,N_24014,N_24013);
or U28707 (N_28707,N_24197,N_26491);
nor U28708 (N_28708,N_26489,N_24477);
nor U28709 (N_28709,N_24582,N_26786);
xor U28710 (N_28710,N_26305,N_24511);
or U28711 (N_28711,N_24488,N_24272);
xnor U28712 (N_28712,N_24275,N_25911);
nand U28713 (N_28713,N_26235,N_25635);
xor U28714 (N_28714,N_24895,N_24717);
xnor U28715 (N_28715,N_25888,N_26285);
nor U28716 (N_28716,N_25687,N_25152);
nor U28717 (N_28717,N_25657,N_25317);
nand U28718 (N_28718,N_25947,N_25143);
or U28719 (N_28719,N_24578,N_26676);
nand U28720 (N_28720,N_26401,N_25259);
and U28721 (N_28721,N_26107,N_26356);
nor U28722 (N_28722,N_25715,N_24758);
and U28723 (N_28723,N_26869,N_25568);
and U28724 (N_28724,N_24792,N_24016);
xnor U28725 (N_28725,N_24124,N_26645);
nand U28726 (N_28726,N_25279,N_25096);
nand U28727 (N_28727,N_25030,N_26015);
nor U28728 (N_28728,N_25433,N_26995);
nor U28729 (N_28729,N_26412,N_25136);
or U28730 (N_28730,N_26762,N_24914);
or U28731 (N_28731,N_24471,N_26310);
or U28732 (N_28732,N_24756,N_24053);
nand U28733 (N_28733,N_24263,N_26488);
nand U28734 (N_28734,N_25875,N_25303);
nand U28735 (N_28735,N_26768,N_25451);
xnor U28736 (N_28736,N_25510,N_24861);
nand U28737 (N_28737,N_24245,N_25087);
xor U28738 (N_28738,N_25920,N_26807);
nand U28739 (N_28739,N_26617,N_26306);
xor U28740 (N_28740,N_24679,N_24060);
nand U28741 (N_28741,N_25838,N_25695);
and U28742 (N_28742,N_26982,N_24714);
and U28743 (N_28743,N_25457,N_25882);
and U28744 (N_28744,N_26462,N_26999);
nor U28745 (N_28745,N_25138,N_24425);
or U28746 (N_28746,N_24927,N_26637);
nand U28747 (N_28747,N_26438,N_26401);
nor U28748 (N_28748,N_26647,N_25273);
or U28749 (N_28749,N_25433,N_25560);
or U28750 (N_28750,N_24516,N_25032);
xnor U28751 (N_28751,N_24360,N_24510);
nor U28752 (N_28752,N_24561,N_25686);
and U28753 (N_28753,N_26596,N_24781);
and U28754 (N_28754,N_24563,N_24211);
nand U28755 (N_28755,N_26809,N_25677);
xnor U28756 (N_28756,N_24763,N_26735);
and U28757 (N_28757,N_25118,N_25317);
or U28758 (N_28758,N_25044,N_25242);
xnor U28759 (N_28759,N_25205,N_25779);
and U28760 (N_28760,N_24688,N_26139);
or U28761 (N_28761,N_25518,N_26210);
or U28762 (N_28762,N_26394,N_24162);
xnor U28763 (N_28763,N_24813,N_24609);
or U28764 (N_28764,N_26786,N_26103);
nor U28765 (N_28765,N_25078,N_24737);
and U28766 (N_28766,N_25364,N_24996);
nor U28767 (N_28767,N_26387,N_24074);
or U28768 (N_28768,N_26590,N_24755);
and U28769 (N_28769,N_25070,N_25830);
nor U28770 (N_28770,N_25738,N_24368);
and U28771 (N_28771,N_26148,N_26593);
nor U28772 (N_28772,N_26485,N_26235);
or U28773 (N_28773,N_24600,N_25091);
nor U28774 (N_28774,N_26310,N_25905);
nand U28775 (N_28775,N_26800,N_24146);
nand U28776 (N_28776,N_24325,N_26181);
and U28777 (N_28777,N_25956,N_25325);
nand U28778 (N_28778,N_26011,N_26180);
xnor U28779 (N_28779,N_25262,N_26942);
and U28780 (N_28780,N_25547,N_26373);
nor U28781 (N_28781,N_24728,N_24847);
nor U28782 (N_28782,N_24211,N_25434);
nand U28783 (N_28783,N_26840,N_26620);
and U28784 (N_28784,N_24606,N_25042);
or U28785 (N_28785,N_24476,N_24919);
xnor U28786 (N_28786,N_25896,N_24357);
or U28787 (N_28787,N_26895,N_24094);
xor U28788 (N_28788,N_26985,N_26147);
and U28789 (N_28789,N_26601,N_26506);
and U28790 (N_28790,N_24777,N_26525);
nand U28791 (N_28791,N_25649,N_24661);
or U28792 (N_28792,N_24298,N_26789);
nor U28793 (N_28793,N_25309,N_25225);
nand U28794 (N_28794,N_25819,N_26397);
nor U28795 (N_28795,N_26471,N_26280);
nor U28796 (N_28796,N_25254,N_25354);
nand U28797 (N_28797,N_24497,N_24234);
nor U28798 (N_28798,N_24077,N_26459);
and U28799 (N_28799,N_24551,N_25232);
nand U28800 (N_28800,N_25918,N_26558);
or U28801 (N_28801,N_24375,N_26072);
nor U28802 (N_28802,N_26298,N_25844);
nand U28803 (N_28803,N_25223,N_25956);
or U28804 (N_28804,N_26449,N_24683);
or U28805 (N_28805,N_24156,N_24257);
or U28806 (N_28806,N_24446,N_24732);
nand U28807 (N_28807,N_25476,N_24963);
xnor U28808 (N_28808,N_25277,N_26840);
or U28809 (N_28809,N_26735,N_26528);
nor U28810 (N_28810,N_26724,N_25860);
or U28811 (N_28811,N_26446,N_26507);
xor U28812 (N_28812,N_25351,N_24774);
and U28813 (N_28813,N_24334,N_26231);
nand U28814 (N_28814,N_25658,N_25006);
nor U28815 (N_28815,N_24707,N_25716);
nand U28816 (N_28816,N_26047,N_24805);
nand U28817 (N_28817,N_24875,N_26587);
nand U28818 (N_28818,N_26942,N_25122);
xnor U28819 (N_28819,N_26134,N_25689);
nor U28820 (N_28820,N_24032,N_25914);
or U28821 (N_28821,N_24797,N_24189);
or U28822 (N_28822,N_25888,N_26615);
or U28823 (N_28823,N_25764,N_24430);
nor U28824 (N_28824,N_26205,N_24593);
and U28825 (N_28825,N_24295,N_24331);
nand U28826 (N_28826,N_24854,N_25921);
and U28827 (N_28827,N_25567,N_24133);
or U28828 (N_28828,N_25862,N_25842);
xnor U28829 (N_28829,N_24837,N_26514);
nand U28830 (N_28830,N_25837,N_24755);
or U28831 (N_28831,N_26330,N_25006);
and U28832 (N_28832,N_26894,N_25399);
xnor U28833 (N_28833,N_25088,N_24426);
and U28834 (N_28834,N_25577,N_26075);
and U28835 (N_28835,N_25895,N_24504);
nor U28836 (N_28836,N_25620,N_26140);
xor U28837 (N_28837,N_24125,N_24413);
xor U28838 (N_28838,N_26802,N_25517);
or U28839 (N_28839,N_24052,N_25520);
nor U28840 (N_28840,N_26910,N_24243);
nor U28841 (N_28841,N_24178,N_24336);
nand U28842 (N_28842,N_26255,N_24187);
xor U28843 (N_28843,N_25763,N_26541);
xor U28844 (N_28844,N_25570,N_26933);
or U28845 (N_28845,N_24240,N_25896);
or U28846 (N_28846,N_25719,N_26192);
or U28847 (N_28847,N_26035,N_26663);
and U28848 (N_28848,N_25023,N_24885);
nand U28849 (N_28849,N_26134,N_24953);
or U28850 (N_28850,N_24297,N_24632);
nor U28851 (N_28851,N_25542,N_24341);
nand U28852 (N_28852,N_26213,N_24548);
nor U28853 (N_28853,N_24776,N_25399);
or U28854 (N_28854,N_24575,N_26614);
nor U28855 (N_28855,N_26389,N_26740);
nor U28856 (N_28856,N_26220,N_24192);
nand U28857 (N_28857,N_25464,N_25682);
nor U28858 (N_28858,N_26199,N_25198);
and U28859 (N_28859,N_25483,N_24221);
or U28860 (N_28860,N_25791,N_24261);
nor U28861 (N_28861,N_26043,N_26934);
or U28862 (N_28862,N_26472,N_26609);
nand U28863 (N_28863,N_24789,N_25972);
and U28864 (N_28864,N_25564,N_25979);
xnor U28865 (N_28865,N_25155,N_24519);
nand U28866 (N_28866,N_26311,N_25873);
or U28867 (N_28867,N_26416,N_25449);
nor U28868 (N_28868,N_26874,N_24941);
nand U28869 (N_28869,N_26169,N_24056);
nor U28870 (N_28870,N_25488,N_26386);
nand U28871 (N_28871,N_24911,N_25878);
nand U28872 (N_28872,N_26848,N_24479);
or U28873 (N_28873,N_26713,N_25775);
nor U28874 (N_28874,N_25525,N_25693);
or U28875 (N_28875,N_25084,N_25592);
or U28876 (N_28876,N_25338,N_24098);
nand U28877 (N_28877,N_24704,N_25323);
nor U28878 (N_28878,N_24160,N_25665);
nand U28879 (N_28879,N_25074,N_24590);
or U28880 (N_28880,N_25464,N_25375);
or U28881 (N_28881,N_26333,N_25213);
xor U28882 (N_28882,N_25183,N_26511);
nor U28883 (N_28883,N_26698,N_26253);
nor U28884 (N_28884,N_25929,N_24641);
and U28885 (N_28885,N_26168,N_26399);
xor U28886 (N_28886,N_26112,N_26893);
and U28887 (N_28887,N_26006,N_25654);
xnor U28888 (N_28888,N_26142,N_25623);
and U28889 (N_28889,N_25146,N_24848);
xor U28890 (N_28890,N_25394,N_24864);
and U28891 (N_28891,N_25471,N_24775);
nor U28892 (N_28892,N_26582,N_25898);
or U28893 (N_28893,N_26349,N_26924);
xor U28894 (N_28894,N_25621,N_24613);
and U28895 (N_28895,N_26778,N_26347);
nand U28896 (N_28896,N_25273,N_26394);
nand U28897 (N_28897,N_24695,N_26563);
and U28898 (N_28898,N_25868,N_25880);
or U28899 (N_28899,N_26546,N_26241);
nand U28900 (N_28900,N_26309,N_24116);
xor U28901 (N_28901,N_25707,N_24925);
nand U28902 (N_28902,N_24468,N_25390);
or U28903 (N_28903,N_25621,N_25257);
nor U28904 (N_28904,N_25957,N_24126);
and U28905 (N_28905,N_24424,N_25303);
nand U28906 (N_28906,N_26994,N_24297);
xor U28907 (N_28907,N_25045,N_26376);
xnor U28908 (N_28908,N_25247,N_24641);
and U28909 (N_28909,N_24702,N_26709);
xor U28910 (N_28910,N_24286,N_26701);
nor U28911 (N_28911,N_25189,N_26702);
and U28912 (N_28912,N_25494,N_24990);
and U28913 (N_28913,N_26091,N_24279);
or U28914 (N_28914,N_26732,N_25258);
and U28915 (N_28915,N_25631,N_25118);
xnor U28916 (N_28916,N_24019,N_24841);
xnor U28917 (N_28917,N_25609,N_25801);
nor U28918 (N_28918,N_24453,N_25436);
and U28919 (N_28919,N_24149,N_25463);
and U28920 (N_28920,N_25191,N_26309);
nand U28921 (N_28921,N_26788,N_24887);
and U28922 (N_28922,N_26269,N_26984);
and U28923 (N_28923,N_25837,N_26143);
nand U28924 (N_28924,N_25098,N_26767);
nand U28925 (N_28925,N_26916,N_24204);
xnor U28926 (N_28926,N_24704,N_25158);
xnor U28927 (N_28927,N_26805,N_26074);
and U28928 (N_28928,N_24725,N_25408);
and U28929 (N_28929,N_24775,N_25378);
or U28930 (N_28930,N_25722,N_26992);
nand U28931 (N_28931,N_25055,N_26882);
and U28932 (N_28932,N_26954,N_24829);
and U28933 (N_28933,N_24023,N_25297);
or U28934 (N_28934,N_24082,N_26925);
xor U28935 (N_28935,N_26852,N_25379);
nor U28936 (N_28936,N_26364,N_24012);
or U28937 (N_28937,N_26678,N_25436);
nor U28938 (N_28938,N_26737,N_24444);
nand U28939 (N_28939,N_24765,N_24155);
xor U28940 (N_28940,N_24814,N_25028);
or U28941 (N_28941,N_26069,N_26291);
nor U28942 (N_28942,N_24354,N_25963);
and U28943 (N_28943,N_26545,N_26085);
nor U28944 (N_28944,N_26472,N_24673);
or U28945 (N_28945,N_25571,N_26197);
and U28946 (N_28946,N_25246,N_25528);
and U28947 (N_28947,N_25459,N_24991);
xor U28948 (N_28948,N_24802,N_24939);
nor U28949 (N_28949,N_26525,N_24353);
xor U28950 (N_28950,N_25326,N_24470);
or U28951 (N_28951,N_25055,N_24945);
or U28952 (N_28952,N_25792,N_26290);
nand U28953 (N_28953,N_26637,N_24372);
xor U28954 (N_28954,N_24344,N_26244);
and U28955 (N_28955,N_24515,N_25709);
xnor U28956 (N_28956,N_24370,N_24325);
nand U28957 (N_28957,N_25548,N_26655);
nor U28958 (N_28958,N_26320,N_26728);
xnor U28959 (N_28959,N_24513,N_25153);
or U28960 (N_28960,N_26879,N_25323);
nor U28961 (N_28961,N_26686,N_25861);
nor U28962 (N_28962,N_24810,N_25810);
and U28963 (N_28963,N_25942,N_24009);
nand U28964 (N_28964,N_26439,N_24608);
nand U28965 (N_28965,N_24634,N_25551);
or U28966 (N_28966,N_24806,N_26936);
or U28967 (N_28967,N_24824,N_25050);
nor U28968 (N_28968,N_24814,N_24100);
xor U28969 (N_28969,N_25381,N_24131);
nor U28970 (N_28970,N_26844,N_26333);
xor U28971 (N_28971,N_25645,N_24325);
or U28972 (N_28972,N_26768,N_25075);
xor U28973 (N_28973,N_26342,N_26825);
xor U28974 (N_28974,N_25394,N_26261);
xor U28975 (N_28975,N_24649,N_24048);
nand U28976 (N_28976,N_25186,N_25660);
or U28977 (N_28977,N_25918,N_24562);
and U28978 (N_28978,N_26676,N_24719);
or U28979 (N_28979,N_26051,N_24815);
nor U28980 (N_28980,N_25310,N_24621);
nand U28981 (N_28981,N_26375,N_26817);
nand U28982 (N_28982,N_24932,N_25945);
and U28983 (N_28983,N_24024,N_26006);
nor U28984 (N_28984,N_25133,N_25079);
xnor U28985 (N_28985,N_26645,N_26051);
or U28986 (N_28986,N_24873,N_25755);
and U28987 (N_28987,N_24285,N_25070);
and U28988 (N_28988,N_26316,N_25895);
xor U28989 (N_28989,N_26656,N_25203);
xnor U28990 (N_28990,N_24920,N_25355);
xnor U28991 (N_28991,N_24827,N_26059);
xnor U28992 (N_28992,N_26511,N_25825);
nor U28993 (N_28993,N_25567,N_25056);
nor U28994 (N_28994,N_25495,N_25170);
xnor U28995 (N_28995,N_25385,N_26431);
or U28996 (N_28996,N_24997,N_25197);
xnor U28997 (N_28997,N_25529,N_26904);
nor U28998 (N_28998,N_25161,N_24243);
or U28999 (N_28999,N_26424,N_24474);
and U29000 (N_29000,N_25205,N_26117);
nand U29001 (N_29001,N_24758,N_25619);
nor U29002 (N_29002,N_26110,N_24833);
or U29003 (N_29003,N_26485,N_25059);
or U29004 (N_29004,N_25989,N_26761);
and U29005 (N_29005,N_24588,N_24155);
nor U29006 (N_29006,N_25466,N_26312);
nor U29007 (N_29007,N_24289,N_26184);
nand U29008 (N_29008,N_24611,N_26675);
xnor U29009 (N_29009,N_24052,N_26342);
or U29010 (N_29010,N_26630,N_26861);
or U29011 (N_29011,N_25773,N_24204);
nand U29012 (N_29012,N_26292,N_24249);
xnor U29013 (N_29013,N_26058,N_25110);
nor U29014 (N_29014,N_26981,N_25070);
and U29015 (N_29015,N_25376,N_24104);
and U29016 (N_29016,N_24535,N_26893);
xor U29017 (N_29017,N_26946,N_25924);
xor U29018 (N_29018,N_24803,N_24626);
and U29019 (N_29019,N_26402,N_24499);
nand U29020 (N_29020,N_24362,N_26377);
nor U29021 (N_29021,N_25762,N_24357);
nor U29022 (N_29022,N_25800,N_25948);
or U29023 (N_29023,N_25169,N_24265);
and U29024 (N_29024,N_25886,N_24582);
nand U29025 (N_29025,N_24092,N_26963);
nor U29026 (N_29026,N_25389,N_24776);
xnor U29027 (N_29027,N_24358,N_26544);
or U29028 (N_29028,N_26842,N_26267);
and U29029 (N_29029,N_24232,N_26555);
xor U29030 (N_29030,N_25092,N_25762);
xnor U29031 (N_29031,N_26010,N_26709);
and U29032 (N_29032,N_25649,N_26638);
or U29033 (N_29033,N_26017,N_26551);
and U29034 (N_29034,N_25930,N_25751);
or U29035 (N_29035,N_25927,N_25970);
and U29036 (N_29036,N_25193,N_26225);
nand U29037 (N_29037,N_26558,N_24807);
or U29038 (N_29038,N_24697,N_25709);
nand U29039 (N_29039,N_25782,N_24527);
and U29040 (N_29040,N_26852,N_24501);
nor U29041 (N_29041,N_26097,N_24452);
nand U29042 (N_29042,N_26375,N_24923);
and U29043 (N_29043,N_24104,N_26528);
and U29044 (N_29044,N_24327,N_25882);
and U29045 (N_29045,N_24031,N_24549);
nor U29046 (N_29046,N_25951,N_25280);
and U29047 (N_29047,N_24001,N_26004);
and U29048 (N_29048,N_24366,N_26283);
nor U29049 (N_29049,N_25555,N_25023);
or U29050 (N_29050,N_24163,N_24877);
xnor U29051 (N_29051,N_25259,N_24335);
nand U29052 (N_29052,N_26250,N_25711);
nor U29053 (N_29053,N_25109,N_25012);
or U29054 (N_29054,N_24362,N_26778);
nand U29055 (N_29055,N_24821,N_25515);
nand U29056 (N_29056,N_26753,N_26321);
and U29057 (N_29057,N_25222,N_24305);
and U29058 (N_29058,N_24434,N_25028);
and U29059 (N_29059,N_26497,N_26611);
nand U29060 (N_29060,N_24082,N_24749);
xor U29061 (N_29061,N_26412,N_26922);
nor U29062 (N_29062,N_26568,N_25346);
xnor U29063 (N_29063,N_25147,N_26808);
or U29064 (N_29064,N_24504,N_25759);
nand U29065 (N_29065,N_26977,N_25467);
and U29066 (N_29066,N_25450,N_24904);
or U29067 (N_29067,N_24250,N_25290);
or U29068 (N_29068,N_24233,N_24985);
xor U29069 (N_29069,N_24065,N_25280);
nand U29070 (N_29070,N_25055,N_25655);
or U29071 (N_29071,N_26984,N_26998);
and U29072 (N_29072,N_25274,N_25245);
and U29073 (N_29073,N_26536,N_24499);
and U29074 (N_29074,N_25206,N_25476);
or U29075 (N_29075,N_24884,N_24161);
nor U29076 (N_29076,N_26579,N_26084);
nand U29077 (N_29077,N_24414,N_24020);
xor U29078 (N_29078,N_25675,N_24074);
or U29079 (N_29079,N_25716,N_25759);
nand U29080 (N_29080,N_24847,N_25777);
nor U29081 (N_29081,N_26357,N_24627);
xnor U29082 (N_29082,N_26655,N_24330);
nor U29083 (N_29083,N_24520,N_24603);
nand U29084 (N_29084,N_26894,N_25557);
nor U29085 (N_29085,N_24491,N_26067);
nand U29086 (N_29086,N_26539,N_26494);
nand U29087 (N_29087,N_24318,N_26250);
and U29088 (N_29088,N_26603,N_26942);
nand U29089 (N_29089,N_25039,N_26097);
nand U29090 (N_29090,N_25817,N_25357);
xnor U29091 (N_29091,N_24170,N_25310);
and U29092 (N_29092,N_26815,N_25325);
nand U29093 (N_29093,N_24640,N_24070);
nand U29094 (N_29094,N_26296,N_24144);
and U29095 (N_29095,N_24591,N_25276);
xnor U29096 (N_29096,N_26147,N_26990);
nor U29097 (N_29097,N_25514,N_24866);
or U29098 (N_29098,N_25025,N_25775);
and U29099 (N_29099,N_26751,N_25990);
or U29100 (N_29100,N_25798,N_24982);
nand U29101 (N_29101,N_24653,N_26889);
nand U29102 (N_29102,N_25260,N_24150);
and U29103 (N_29103,N_25836,N_24689);
xnor U29104 (N_29104,N_26044,N_25089);
and U29105 (N_29105,N_25711,N_24396);
and U29106 (N_29106,N_25052,N_24905);
and U29107 (N_29107,N_25254,N_26084);
xnor U29108 (N_29108,N_26458,N_24076);
nand U29109 (N_29109,N_26007,N_24719);
and U29110 (N_29110,N_24690,N_24953);
and U29111 (N_29111,N_24207,N_25707);
nor U29112 (N_29112,N_24043,N_24790);
or U29113 (N_29113,N_26364,N_25859);
and U29114 (N_29114,N_25336,N_26754);
or U29115 (N_29115,N_26056,N_24769);
xnor U29116 (N_29116,N_25324,N_26720);
and U29117 (N_29117,N_25840,N_26632);
nor U29118 (N_29118,N_26848,N_26851);
nand U29119 (N_29119,N_24562,N_26105);
nor U29120 (N_29120,N_25228,N_26303);
and U29121 (N_29121,N_24982,N_24290);
xor U29122 (N_29122,N_26505,N_25890);
xor U29123 (N_29123,N_24356,N_24998);
or U29124 (N_29124,N_26699,N_26081);
xnor U29125 (N_29125,N_24634,N_26097);
or U29126 (N_29126,N_24133,N_25197);
or U29127 (N_29127,N_26264,N_24414);
and U29128 (N_29128,N_25029,N_26284);
xnor U29129 (N_29129,N_25177,N_26086);
or U29130 (N_29130,N_25705,N_25273);
or U29131 (N_29131,N_26831,N_24048);
nor U29132 (N_29132,N_26223,N_24482);
nand U29133 (N_29133,N_25158,N_26551);
nand U29134 (N_29134,N_26581,N_24350);
or U29135 (N_29135,N_25828,N_25891);
and U29136 (N_29136,N_24020,N_26407);
xor U29137 (N_29137,N_24481,N_25497);
nor U29138 (N_29138,N_25606,N_26537);
xnor U29139 (N_29139,N_26360,N_26006);
and U29140 (N_29140,N_24736,N_25089);
nor U29141 (N_29141,N_24332,N_25451);
and U29142 (N_29142,N_25060,N_25488);
nor U29143 (N_29143,N_24305,N_24582);
and U29144 (N_29144,N_26381,N_26618);
nor U29145 (N_29145,N_25202,N_24924);
and U29146 (N_29146,N_25313,N_25495);
nand U29147 (N_29147,N_25927,N_24476);
nand U29148 (N_29148,N_24415,N_24445);
or U29149 (N_29149,N_24872,N_26907);
xor U29150 (N_29150,N_24530,N_24831);
nand U29151 (N_29151,N_26996,N_26320);
nand U29152 (N_29152,N_24940,N_24838);
nand U29153 (N_29153,N_26206,N_25576);
and U29154 (N_29154,N_26970,N_26436);
nor U29155 (N_29155,N_26927,N_24679);
xnor U29156 (N_29156,N_24954,N_25883);
nand U29157 (N_29157,N_25605,N_24087);
nor U29158 (N_29158,N_26079,N_25818);
and U29159 (N_29159,N_25852,N_24538);
xnor U29160 (N_29160,N_26689,N_26139);
or U29161 (N_29161,N_26199,N_24214);
xor U29162 (N_29162,N_26380,N_24291);
xor U29163 (N_29163,N_25424,N_25980);
nor U29164 (N_29164,N_26012,N_25355);
and U29165 (N_29165,N_24292,N_25927);
and U29166 (N_29166,N_24248,N_25328);
and U29167 (N_29167,N_24569,N_25125);
nor U29168 (N_29168,N_24385,N_26653);
nor U29169 (N_29169,N_26541,N_26313);
or U29170 (N_29170,N_25036,N_26487);
or U29171 (N_29171,N_26205,N_26247);
or U29172 (N_29172,N_24439,N_25040);
xnor U29173 (N_29173,N_25565,N_24232);
nand U29174 (N_29174,N_24460,N_24764);
nand U29175 (N_29175,N_24910,N_26675);
xnor U29176 (N_29176,N_25226,N_26334);
nor U29177 (N_29177,N_25605,N_26868);
nor U29178 (N_29178,N_24403,N_26987);
xor U29179 (N_29179,N_26635,N_26890);
nor U29180 (N_29180,N_26496,N_24601);
and U29181 (N_29181,N_25057,N_26091);
nand U29182 (N_29182,N_25567,N_25127);
xnor U29183 (N_29183,N_26375,N_25047);
nor U29184 (N_29184,N_24891,N_26235);
and U29185 (N_29185,N_26812,N_25562);
and U29186 (N_29186,N_25451,N_24730);
or U29187 (N_29187,N_26477,N_26437);
and U29188 (N_29188,N_26910,N_25441);
nand U29189 (N_29189,N_25214,N_26450);
or U29190 (N_29190,N_26198,N_26437);
xnor U29191 (N_29191,N_26353,N_26042);
nand U29192 (N_29192,N_24148,N_24405);
nand U29193 (N_29193,N_25529,N_26841);
or U29194 (N_29194,N_24824,N_24715);
xor U29195 (N_29195,N_24276,N_26371);
nor U29196 (N_29196,N_25087,N_25280);
and U29197 (N_29197,N_24442,N_25008);
nor U29198 (N_29198,N_25930,N_26519);
nor U29199 (N_29199,N_24076,N_25609);
nor U29200 (N_29200,N_24239,N_24215);
nor U29201 (N_29201,N_25753,N_26536);
nor U29202 (N_29202,N_24873,N_25525);
or U29203 (N_29203,N_24787,N_26771);
and U29204 (N_29204,N_25891,N_26485);
nor U29205 (N_29205,N_26153,N_25641);
nand U29206 (N_29206,N_24028,N_24989);
nor U29207 (N_29207,N_24705,N_24838);
xor U29208 (N_29208,N_26395,N_24920);
or U29209 (N_29209,N_24679,N_25095);
nor U29210 (N_29210,N_24377,N_24174);
nand U29211 (N_29211,N_26054,N_24257);
xor U29212 (N_29212,N_26811,N_25522);
nand U29213 (N_29213,N_24306,N_26170);
or U29214 (N_29214,N_26444,N_26483);
and U29215 (N_29215,N_24990,N_25421);
nand U29216 (N_29216,N_25019,N_26248);
and U29217 (N_29217,N_25422,N_25324);
and U29218 (N_29218,N_26360,N_24936);
and U29219 (N_29219,N_24762,N_26369);
and U29220 (N_29220,N_25312,N_26834);
xnor U29221 (N_29221,N_25925,N_24076);
xnor U29222 (N_29222,N_26970,N_24465);
and U29223 (N_29223,N_25252,N_24395);
nand U29224 (N_29224,N_26924,N_25522);
nor U29225 (N_29225,N_24716,N_25195);
xor U29226 (N_29226,N_26064,N_24622);
nor U29227 (N_29227,N_25084,N_26542);
or U29228 (N_29228,N_26251,N_26915);
nand U29229 (N_29229,N_24508,N_24220);
or U29230 (N_29230,N_26708,N_25642);
nand U29231 (N_29231,N_24651,N_24450);
and U29232 (N_29232,N_25705,N_24245);
xor U29233 (N_29233,N_26722,N_25207);
nor U29234 (N_29234,N_24498,N_26646);
nand U29235 (N_29235,N_25927,N_26217);
nor U29236 (N_29236,N_26595,N_25718);
xnor U29237 (N_29237,N_25911,N_24092);
nor U29238 (N_29238,N_25200,N_24200);
nand U29239 (N_29239,N_26903,N_24514);
and U29240 (N_29240,N_26958,N_24472);
and U29241 (N_29241,N_26411,N_26166);
nand U29242 (N_29242,N_25424,N_26988);
xnor U29243 (N_29243,N_25019,N_24561);
nor U29244 (N_29244,N_24300,N_24897);
or U29245 (N_29245,N_25277,N_24199);
nand U29246 (N_29246,N_24384,N_26461);
or U29247 (N_29247,N_26904,N_25608);
xor U29248 (N_29248,N_24399,N_25541);
nor U29249 (N_29249,N_25113,N_26236);
and U29250 (N_29250,N_26159,N_25291);
xor U29251 (N_29251,N_24095,N_24505);
nor U29252 (N_29252,N_25040,N_25619);
nor U29253 (N_29253,N_25463,N_25531);
xnor U29254 (N_29254,N_26790,N_26494);
nand U29255 (N_29255,N_24247,N_24156);
nand U29256 (N_29256,N_24500,N_24390);
and U29257 (N_29257,N_25250,N_26187);
xor U29258 (N_29258,N_24834,N_24347);
xor U29259 (N_29259,N_25862,N_25502);
or U29260 (N_29260,N_25650,N_24112);
and U29261 (N_29261,N_24424,N_24138);
and U29262 (N_29262,N_25460,N_25660);
xnor U29263 (N_29263,N_24663,N_25116);
xnor U29264 (N_29264,N_25511,N_25284);
or U29265 (N_29265,N_26197,N_25436);
nand U29266 (N_29266,N_26804,N_25150);
and U29267 (N_29267,N_25492,N_25986);
nor U29268 (N_29268,N_24091,N_26794);
xnor U29269 (N_29269,N_25436,N_24133);
and U29270 (N_29270,N_25226,N_26992);
xnor U29271 (N_29271,N_26755,N_26994);
xor U29272 (N_29272,N_24217,N_26389);
xor U29273 (N_29273,N_26214,N_25953);
or U29274 (N_29274,N_24835,N_25349);
nand U29275 (N_29275,N_24775,N_24678);
or U29276 (N_29276,N_25988,N_25952);
nor U29277 (N_29277,N_26388,N_24234);
nor U29278 (N_29278,N_25764,N_24297);
or U29279 (N_29279,N_24763,N_26671);
and U29280 (N_29280,N_26286,N_25798);
nand U29281 (N_29281,N_24546,N_24081);
or U29282 (N_29282,N_25442,N_24885);
nand U29283 (N_29283,N_25186,N_26256);
nor U29284 (N_29284,N_25766,N_24402);
or U29285 (N_29285,N_25100,N_26475);
or U29286 (N_29286,N_24455,N_26263);
or U29287 (N_29287,N_25865,N_24087);
xor U29288 (N_29288,N_24356,N_26954);
and U29289 (N_29289,N_26428,N_25910);
xor U29290 (N_29290,N_26349,N_26146);
nor U29291 (N_29291,N_25144,N_25515);
and U29292 (N_29292,N_24886,N_24982);
nand U29293 (N_29293,N_26539,N_24568);
nand U29294 (N_29294,N_26225,N_24010);
or U29295 (N_29295,N_25688,N_24590);
or U29296 (N_29296,N_24459,N_25889);
nand U29297 (N_29297,N_26436,N_25771);
xor U29298 (N_29298,N_26395,N_26054);
nand U29299 (N_29299,N_24735,N_24080);
nand U29300 (N_29300,N_24546,N_26384);
xnor U29301 (N_29301,N_24434,N_26617);
xor U29302 (N_29302,N_25841,N_24320);
nor U29303 (N_29303,N_26885,N_26695);
nor U29304 (N_29304,N_25581,N_26249);
or U29305 (N_29305,N_25972,N_26607);
nor U29306 (N_29306,N_25102,N_26203);
and U29307 (N_29307,N_25956,N_26560);
xnor U29308 (N_29308,N_26876,N_26035);
nor U29309 (N_29309,N_25221,N_24882);
and U29310 (N_29310,N_24593,N_25330);
or U29311 (N_29311,N_25126,N_25065);
xor U29312 (N_29312,N_25624,N_24485);
nor U29313 (N_29313,N_25306,N_24718);
and U29314 (N_29314,N_24416,N_25846);
nor U29315 (N_29315,N_26145,N_24958);
nand U29316 (N_29316,N_26233,N_25532);
nand U29317 (N_29317,N_26572,N_26675);
and U29318 (N_29318,N_24927,N_26365);
nor U29319 (N_29319,N_25712,N_25015);
nor U29320 (N_29320,N_24453,N_25549);
nor U29321 (N_29321,N_26347,N_26375);
or U29322 (N_29322,N_26568,N_25679);
and U29323 (N_29323,N_26143,N_25819);
nor U29324 (N_29324,N_26349,N_26490);
xnor U29325 (N_29325,N_25257,N_26042);
and U29326 (N_29326,N_24105,N_24360);
nand U29327 (N_29327,N_25666,N_26695);
nor U29328 (N_29328,N_25199,N_26363);
or U29329 (N_29329,N_24325,N_26000);
and U29330 (N_29330,N_24730,N_24745);
nor U29331 (N_29331,N_24558,N_24872);
nand U29332 (N_29332,N_24139,N_26107);
and U29333 (N_29333,N_24405,N_24127);
nand U29334 (N_29334,N_26620,N_24665);
and U29335 (N_29335,N_25394,N_25477);
and U29336 (N_29336,N_24378,N_24345);
nand U29337 (N_29337,N_26353,N_26932);
or U29338 (N_29338,N_25881,N_24893);
nand U29339 (N_29339,N_25370,N_26441);
xor U29340 (N_29340,N_26888,N_26610);
or U29341 (N_29341,N_24014,N_26875);
or U29342 (N_29342,N_26040,N_26119);
xnor U29343 (N_29343,N_26650,N_26810);
and U29344 (N_29344,N_24965,N_26605);
or U29345 (N_29345,N_26847,N_25774);
or U29346 (N_29346,N_25413,N_24300);
and U29347 (N_29347,N_25206,N_26029);
nand U29348 (N_29348,N_25275,N_24376);
nand U29349 (N_29349,N_24103,N_25385);
xnor U29350 (N_29350,N_24851,N_25561);
nand U29351 (N_29351,N_26935,N_25773);
and U29352 (N_29352,N_24396,N_26558);
or U29353 (N_29353,N_25583,N_25247);
nor U29354 (N_29354,N_24693,N_26915);
xor U29355 (N_29355,N_24437,N_24223);
nor U29356 (N_29356,N_25407,N_25437);
nand U29357 (N_29357,N_26727,N_25878);
and U29358 (N_29358,N_26858,N_26525);
nand U29359 (N_29359,N_24591,N_26731);
or U29360 (N_29360,N_25515,N_25146);
xor U29361 (N_29361,N_24403,N_26609);
nor U29362 (N_29362,N_25064,N_26706);
nand U29363 (N_29363,N_25526,N_26542);
or U29364 (N_29364,N_24702,N_25027);
nand U29365 (N_29365,N_26809,N_26325);
xor U29366 (N_29366,N_26825,N_26513);
nand U29367 (N_29367,N_26875,N_26332);
xnor U29368 (N_29368,N_24945,N_24753);
nand U29369 (N_29369,N_24925,N_24491);
nor U29370 (N_29370,N_26789,N_25001);
and U29371 (N_29371,N_25368,N_26014);
or U29372 (N_29372,N_25521,N_24781);
nand U29373 (N_29373,N_25471,N_25804);
xor U29374 (N_29374,N_24795,N_25717);
xnor U29375 (N_29375,N_24552,N_26821);
and U29376 (N_29376,N_25776,N_24582);
or U29377 (N_29377,N_24521,N_24240);
nor U29378 (N_29378,N_25373,N_25436);
nand U29379 (N_29379,N_26307,N_26410);
xor U29380 (N_29380,N_25792,N_26309);
nor U29381 (N_29381,N_25228,N_25345);
and U29382 (N_29382,N_24716,N_25346);
nand U29383 (N_29383,N_25356,N_25545);
xor U29384 (N_29384,N_24869,N_25648);
xor U29385 (N_29385,N_25591,N_26236);
nand U29386 (N_29386,N_25650,N_24810);
nand U29387 (N_29387,N_25116,N_24974);
and U29388 (N_29388,N_25537,N_26362);
and U29389 (N_29389,N_26240,N_24384);
or U29390 (N_29390,N_25334,N_24240);
xnor U29391 (N_29391,N_26308,N_24050);
or U29392 (N_29392,N_26493,N_24012);
xor U29393 (N_29393,N_26227,N_25964);
nand U29394 (N_29394,N_26787,N_25652);
and U29395 (N_29395,N_24246,N_25794);
xor U29396 (N_29396,N_25955,N_24413);
and U29397 (N_29397,N_25250,N_24114);
or U29398 (N_29398,N_25761,N_24098);
and U29399 (N_29399,N_26761,N_25913);
nand U29400 (N_29400,N_26571,N_26077);
xor U29401 (N_29401,N_25419,N_24973);
nand U29402 (N_29402,N_24882,N_25184);
xnor U29403 (N_29403,N_24430,N_26994);
nor U29404 (N_29404,N_24616,N_26693);
xnor U29405 (N_29405,N_24177,N_26981);
nor U29406 (N_29406,N_26594,N_25195);
or U29407 (N_29407,N_25733,N_25103);
nand U29408 (N_29408,N_24510,N_24507);
and U29409 (N_29409,N_24986,N_24099);
xor U29410 (N_29410,N_24940,N_24436);
nand U29411 (N_29411,N_26780,N_24518);
nand U29412 (N_29412,N_24303,N_26825);
and U29413 (N_29413,N_26922,N_24519);
xor U29414 (N_29414,N_26089,N_25666);
nor U29415 (N_29415,N_25939,N_26682);
and U29416 (N_29416,N_26846,N_25208);
nand U29417 (N_29417,N_24511,N_25291);
or U29418 (N_29418,N_25500,N_26075);
nand U29419 (N_29419,N_24613,N_24154);
nand U29420 (N_29420,N_25982,N_24921);
nand U29421 (N_29421,N_26134,N_24747);
nor U29422 (N_29422,N_25771,N_25220);
nand U29423 (N_29423,N_26182,N_26981);
xnor U29424 (N_29424,N_25810,N_25299);
and U29425 (N_29425,N_24297,N_26370);
xnor U29426 (N_29426,N_25887,N_24433);
or U29427 (N_29427,N_25656,N_24465);
and U29428 (N_29428,N_26334,N_25602);
nand U29429 (N_29429,N_24149,N_25466);
or U29430 (N_29430,N_24475,N_26696);
nor U29431 (N_29431,N_26359,N_26000);
and U29432 (N_29432,N_25752,N_26921);
xor U29433 (N_29433,N_25354,N_25224);
and U29434 (N_29434,N_26129,N_25943);
nor U29435 (N_29435,N_25270,N_26814);
or U29436 (N_29436,N_26565,N_25315);
xnor U29437 (N_29437,N_26437,N_24238);
and U29438 (N_29438,N_25853,N_25011);
and U29439 (N_29439,N_25597,N_24166);
xnor U29440 (N_29440,N_24039,N_26193);
nand U29441 (N_29441,N_24548,N_24128);
and U29442 (N_29442,N_26723,N_24184);
or U29443 (N_29443,N_25195,N_24762);
and U29444 (N_29444,N_24571,N_24986);
xnor U29445 (N_29445,N_26145,N_24129);
or U29446 (N_29446,N_26112,N_25139);
nor U29447 (N_29447,N_24635,N_26507);
nor U29448 (N_29448,N_24241,N_26355);
nor U29449 (N_29449,N_25999,N_24912);
and U29450 (N_29450,N_26030,N_26165);
nor U29451 (N_29451,N_26789,N_26268);
and U29452 (N_29452,N_24823,N_24306);
nand U29453 (N_29453,N_26836,N_26428);
nor U29454 (N_29454,N_24110,N_24124);
and U29455 (N_29455,N_26917,N_25465);
and U29456 (N_29456,N_26384,N_26773);
xor U29457 (N_29457,N_26621,N_26975);
or U29458 (N_29458,N_26232,N_24147);
xnor U29459 (N_29459,N_25745,N_24422);
nand U29460 (N_29460,N_25472,N_24062);
and U29461 (N_29461,N_26300,N_26886);
and U29462 (N_29462,N_25880,N_25145);
xnor U29463 (N_29463,N_24253,N_24661);
nand U29464 (N_29464,N_26599,N_26010);
nand U29465 (N_29465,N_24809,N_25435);
and U29466 (N_29466,N_26807,N_26556);
xor U29467 (N_29467,N_26868,N_24442);
nand U29468 (N_29468,N_24182,N_24566);
nor U29469 (N_29469,N_26933,N_25498);
or U29470 (N_29470,N_24316,N_25941);
nor U29471 (N_29471,N_24571,N_24736);
nor U29472 (N_29472,N_24444,N_25201);
and U29473 (N_29473,N_25998,N_26486);
or U29474 (N_29474,N_24947,N_25228);
nand U29475 (N_29475,N_25307,N_25982);
xnor U29476 (N_29476,N_26119,N_26519);
or U29477 (N_29477,N_24294,N_26650);
nand U29478 (N_29478,N_26894,N_25037);
or U29479 (N_29479,N_24724,N_26152);
and U29480 (N_29480,N_26301,N_24178);
xnor U29481 (N_29481,N_26587,N_25003);
nor U29482 (N_29482,N_24030,N_26151);
nor U29483 (N_29483,N_26028,N_24811);
nand U29484 (N_29484,N_26273,N_25549);
xnor U29485 (N_29485,N_24588,N_25438);
or U29486 (N_29486,N_24280,N_26410);
nand U29487 (N_29487,N_25887,N_24811);
nand U29488 (N_29488,N_26469,N_24177);
xor U29489 (N_29489,N_25360,N_25632);
xor U29490 (N_29490,N_24457,N_26094);
and U29491 (N_29491,N_24244,N_24337);
nand U29492 (N_29492,N_25373,N_24553);
nor U29493 (N_29493,N_25275,N_24080);
and U29494 (N_29494,N_24499,N_26610);
nand U29495 (N_29495,N_24843,N_25672);
or U29496 (N_29496,N_26627,N_26950);
nor U29497 (N_29497,N_25143,N_26660);
nand U29498 (N_29498,N_26701,N_25406);
nor U29499 (N_29499,N_26881,N_25264);
nand U29500 (N_29500,N_25731,N_24800);
or U29501 (N_29501,N_26272,N_24252);
or U29502 (N_29502,N_26263,N_26896);
nand U29503 (N_29503,N_26045,N_24029);
or U29504 (N_29504,N_24202,N_25503);
nor U29505 (N_29505,N_26514,N_24812);
nor U29506 (N_29506,N_25895,N_26743);
xor U29507 (N_29507,N_26034,N_25637);
and U29508 (N_29508,N_26347,N_24397);
xnor U29509 (N_29509,N_24715,N_26763);
nor U29510 (N_29510,N_24563,N_26019);
or U29511 (N_29511,N_26367,N_26490);
xnor U29512 (N_29512,N_25402,N_25013);
or U29513 (N_29513,N_26688,N_24237);
xnor U29514 (N_29514,N_25204,N_24552);
and U29515 (N_29515,N_25215,N_26558);
and U29516 (N_29516,N_26501,N_24458);
or U29517 (N_29517,N_26672,N_25813);
nor U29518 (N_29518,N_26211,N_25380);
nand U29519 (N_29519,N_26519,N_26940);
and U29520 (N_29520,N_26970,N_26743);
and U29521 (N_29521,N_24215,N_26662);
or U29522 (N_29522,N_24219,N_25563);
nor U29523 (N_29523,N_25672,N_24853);
xor U29524 (N_29524,N_26684,N_25601);
and U29525 (N_29525,N_24643,N_26884);
or U29526 (N_29526,N_25426,N_25199);
nand U29527 (N_29527,N_26350,N_24157);
nand U29528 (N_29528,N_25277,N_26561);
or U29529 (N_29529,N_24536,N_25032);
nor U29530 (N_29530,N_25998,N_24675);
or U29531 (N_29531,N_25498,N_26928);
nor U29532 (N_29532,N_25976,N_25718);
or U29533 (N_29533,N_24178,N_25832);
xor U29534 (N_29534,N_25949,N_24640);
nor U29535 (N_29535,N_25776,N_26696);
xor U29536 (N_29536,N_25241,N_26439);
or U29537 (N_29537,N_26622,N_24834);
xnor U29538 (N_29538,N_24667,N_25487);
xor U29539 (N_29539,N_25804,N_25795);
and U29540 (N_29540,N_24160,N_25564);
xor U29541 (N_29541,N_26032,N_24628);
or U29542 (N_29542,N_24566,N_24089);
or U29543 (N_29543,N_25015,N_26305);
and U29544 (N_29544,N_26721,N_26902);
or U29545 (N_29545,N_25230,N_25585);
xnor U29546 (N_29546,N_25634,N_25254);
or U29547 (N_29547,N_24913,N_25570);
or U29548 (N_29548,N_26820,N_25471);
nand U29549 (N_29549,N_26569,N_25497);
and U29550 (N_29550,N_24543,N_26177);
nor U29551 (N_29551,N_25079,N_26346);
nor U29552 (N_29552,N_25991,N_26929);
nor U29553 (N_29553,N_24610,N_25506);
and U29554 (N_29554,N_24115,N_25150);
and U29555 (N_29555,N_24176,N_24809);
or U29556 (N_29556,N_25685,N_24628);
nand U29557 (N_29557,N_26771,N_24868);
and U29558 (N_29558,N_25476,N_26847);
and U29559 (N_29559,N_26078,N_25404);
nor U29560 (N_29560,N_24480,N_24901);
and U29561 (N_29561,N_26214,N_25586);
and U29562 (N_29562,N_25247,N_25057);
xor U29563 (N_29563,N_24519,N_24193);
nand U29564 (N_29564,N_25959,N_25168);
nand U29565 (N_29565,N_26900,N_24341);
nor U29566 (N_29566,N_25264,N_24518);
nor U29567 (N_29567,N_24322,N_26584);
or U29568 (N_29568,N_24948,N_26188);
nor U29569 (N_29569,N_26060,N_24760);
or U29570 (N_29570,N_24257,N_26829);
and U29571 (N_29571,N_25877,N_26853);
nor U29572 (N_29572,N_25560,N_24911);
or U29573 (N_29573,N_25662,N_24740);
nand U29574 (N_29574,N_25550,N_26847);
nor U29575 (N_29575,N_24703,N_25339);
nor U29576 (N_29576,N_25078,N_24957);
nor U29577 (N_29577,N_25281,N_26637);
and U29578 (N_29578,N_26348,N_25477);
nand U29579 (N_29579,N_25643,N_24579);
and U29580 (N_29580,N_26743,N_25427);
nand U29581 (N_29581,N_25203,N_26828);
and U29582 (N_29582,N_25038,N_24930);
nand U29583 (N_29583,N_26043,N_26628);
or U29584 (N_29584,N_26369,N_25206);
nand U29585 (N_29585,N_26041,N_24481);
or U29586 (N_29586,N_26407,N_24951);
or U29587 (N_29587,N_25118,N_25457);
nor U29588 (N_29588,N_24140,N_26349);
nand U29589 (N_29589,N_25688,N_26287);
or U29590 (N_29590,N_25628,N_24132);
and U29591 (N_29591,N_24350,N_24593);
or U29592 (N_29592,N_25876,N_26534);
or U29593 (N_29593,N_25054,N_25558);
nand U29594 (N_29594,N_26724,N_26676);
nor U29595 (N_29595,N_26890,N_26709);
xnor U29596 (N_29596,N_25157,N_25099);
xor U29597 (N_29597,N_25185,N_24602);
and U29598 (N_29598,N_25332,N_24482);
nand U29599 (N_29599,N_25919,N_26299);
and U29600 (N_29600,N_25783,N_25716);
or U29601 (N_29601,N_24590,N_25048);
and U29602 (N_29602,N_26523,N_26092);
nand U29603 (N_29603,N_26453,N_26195);
nand U29604 (N_29604,N_24442,N_25653);
nor U29605 (N_29605,N_25386,N_24654);
xnor U29606 (N_29606,N_24095,N_24412);
xnor U29607 (N_29607,N_25673,N_25410);
nand U29608 (N_29608,N_26842,N_25982);
nor U29609 (N_29609,N_26681,N_26080);
nor U29610 (N_29610,N_26256,N_24700);
xnor U29611 (N_29611,N_26645,N_26046);
nor U29612 (N_29612,N_26174,N_25261);
xnor U29613 (N_29613,N_25909,N_25927);
xor U29614 (N_29614,N_25820,N_26264);
and U29615 (N_29615,N_26002,N_24984);
nor U29616 (N_29616,N_25944,N_25975);
nand U29617 (N_29617,N_24386,N_24976);
xor U29618 (N_29618,N_25212,N_26516);
xor U29619 (N_29619,N_25229,N_24636);
and U29620 (N_29620,N_24255,N_26301);
and U29621 (N_29621,N_24695,N_24930);
and U29622 (N_29622,N_24875,N_24212);
xnor U29623 (N_29623,N_25750,N_26572);
and U29624 (N_29624,N_25285,N_24217);
nand U29625 (N_29625,N_26473,N_24692);
and U29626 (N_29626,N_24931,N_24489);
or U29627 (N_29627,N_25570,N_25177);
nor U29628 (N_29628,N_25828,N_25371);
and U29629 (N_29629,N_24100,N_26097);
xnor U29630 (N_29630,N_24361,N_25988);
nor U29631 (N_29631,N_26465,N_25480);
or U29632 (N_29632,N_26730,N_25453);
or U29633 (N_29633,N_26688,N_26858);
nor U29634 (N_29634,N_26703,N_24465);
nor U29635 (N_29635,N_26455,N_26588);
or U29636 (N_29636,N_24380,N_24060);
or U29637 (N_29637,N_25246,N_25376);
nor U29638 (N_29638,N_24071,N_26347);
nand U29639 (N_29639,N_25079,N_24218);
or U29640 (N_29640,N_24121,N_24587);
or U29641 (N_29641,N_25139,N_24513);
and U29642 (N_29642,N_24569,N_25538);
xor U29643 (N_29643,N_26861,N_26360);
nand U29644 (N_29644,N_26818,N_25220);
nand U29645 (N_29645,N_25137,N_26515);
nor U29646 (N_29646,N_25673,N_25795);
xor U29647 (N_29647,N_25808,N_26786);
and U29648 (N_29648,N_24300,N_26472);
nand U29649 (N_29649,N_26173,N_25695);
or U29650 (N_29650,N_24678,N_24497);
xnor U29651 (N_29651,N_25114,N_25627);
or U29652 (N_29652,N_26017,N_24052);
xor U29653 (N_29653,N_26225,N_25877);
and U29654 (N_29654,N_24576,N_26992);
and U29655 (N_29655,N_26995,N_24566);
nor U29656 (N_29656,N_25277,N_26176);
xor U29657 (N_29657,N_24584,N_26198);
xor U29658 (N_29658,N_24438,N_24913);
nor U29659 (N_29659,N_25884,N_25964);
or U29660 (N_29660,N_25596,N_25512);
nor U29661 (N_29661,N_24552,N_25964);
nor U29662 (N_29662,N_24017,N_25936);
nor U29663 (N_29663,N_26833,N_26850);
or U29664 (N_29664,N_26466,N_24270);
nor U29665 (N_29665,N_26396,N_25763);
and U29666 (N_29666,N_25665,N_24249);
nand U29667 (N_29667,N_24145,N_26963);
xor U29668 (N_29668,N_24205,N_25828);
and U29669 (N_29669,N_26160,N_25950);
nand U29670 (N_29670,N_25487,N_24029);
nand U29671 (N_29671,N_25312,N_25978);
or U29672 (N_29672,N_25919,N_25201);
and U29673 (N_29673,N_25670,N_24874);
xor U29674 (N_29674,N_26342,N_25548);
or U29675 (N_29675,N_26525,N_25559);
xor U29676 (N_29676,N_24528,N_25861);
nand U29677 (N_29677,N_24975,N_26825);
nand U29678 (N_29678,N_25885,N_24351);
nand U29679 (N_29679,N_25157,N_26018);
nand U29680 (N_29680,N_25462,N_26244);
nand U29681 (N_29681,N_24991,N_25813);
nand U29682 (N_29682,N_25180,N_24280);
and U29683 (N_29683,N_25695,N_24124);
nand U29684 (N_29684,N_25144,N_26251);
xor U29685 (N_29685,N_26658,N_25065);
nor U29686 (N_29686,N_24785,N_26729);
or U29687 (N_29687,N_25906,N_24752);
or U29688 (N_29688,N_24731,N_25250);
or U29689 (N_29689,N_26838,N_26878);
or U29690 (N_29690,N_24224,N_24572);
or U29691 (N_29691,N_25083,N_24013);
nor U29692 (N_29692,N_26986,N_25982);
nand U29693 (N_29693,N_24354,N_26259);
nor U29694 (N_29694,N_25772,N_24874);
nor U29695 (N_29695,N_26265,N_26191);
and U29696 (N_29696,N_25372,N_24424);
xor U29697 (N_29697,N_25699,N_24095);
and U29698 (N_29698,N_24015,N_26441);
nand U29699 (N_29699,N_26433,N_24466);
nor U29700 (N_29700,N_26836,N_25167);
and U29701 (N_29701,N_24238,N_26102);
xor U29702 (N_29702,N_26368,N_26965);
nor U29703 (N_29703,N_25315,N_24121);
nand U29704 (N_29704,N_25014,N_24189);
and U29705 (N_29705,N_26534,N_26050);
nand U29706 (N_29706,N_24129,N_24525);
xor U29707 (N_29707,N_26952,N_26990);
or U29708 (N_29708,N_25681,N_24282);
or U29709 (N_29709,N_26208,N_24507);
and U29710 (N_29710,N_24429,N_25234);
or U29711 (N_29711,N_26322,N_24247);
xnor U29712 (N_29712,N_25622,N_24089);
or U29713 (N_29713,N_26955,N_26885);
nand U29714 (N_29714,N_25890,N_24285);
and U29715 (N_29715,N_24786,N_26023);
xor U29716 (N_29716,N_24356,N_24983);
and U29717 (N_29717,N_26450,N_25712);
or U29718 (N_29718,N_25765,N_26547);
xnor U29719 (N_29719,N_25491,N_26722);
and U29720 (N_29720,N_26260,N_25962);
nor U29721 (N_29721,N_24392,N_24578);
nor U29722 (N_29722,N_26818,N_24593);
nand U29723 (N_29723,N_25385,N_26952);
nor U29724 (N_29724,N_26836,N_24201);
or U29725 (N_29725,N_26639,N_26782);
or U29726 (N_29726,N_24462,N_26629);
xnor U29727 (N_29727,N_25458,N_25929);
and U29728 (N_29728,N_24431,N_25606);
or U29729 (N_29729,N_26729,N_24056);
nor U29730 (N_29730,N_25429,N_26747);
xor U29731 (N_29731,N_25771,N_25151);
and U29732 (N_29732,N_24947,N_26580);
nor U29733 (N_29733,N_24899,N_25571);
xor U29734 (N_29734,N_26756,N_24210);
xor U29735 (N_29735,N_24054,N_25029);
nand U29736 (N_29736,N_26905,N_26747);
nor U29737 (N_29737,N_24853,N_26266);
nand U29738 (N_29738,N_24200,N_24847);
or U29739 (N_29739,N_25242,N_24654);
nand U29740 (N_29740,N_26089,N_24516);
xnor U29741 (N_29741,N_26212,N_25656);
nor U29742 (N_29742,N_24761,N_26324);
nor U29743 (N_29743,N_25064,N_25004);
nand U29744 (N_29744,N_25588,N_26592);
xor U29745 (N_29745,N_25239,N_25905);
or U29746 (N_29746,N_24096,N_24181);
and U29747 (N_29747,N_26028,N_24931);
or U29748 (N_29748,N_24263,N_24249);
nor U29749 (N_29749,N_26897,N_24922);
or U29750 (N_29750,N_25928,N_24061);
or U29751 (N_29751,N_25023,N_26162);
nand U29752 (N_29752,N_25669,N_26567);
or U29753 (N_29753,N_24553,N_25195);
and U29754 (N_29754,N_24441,N_26847);
nor U29755 (N_29755,N_25361,N_24615);
or U29756 (N_29756,N_26753,N_25860);
and U29757 (N_29757,N_26126,N_24616);
nand U29758 (N_29758,N_26359,N_25465);
and U29759 (N_29759,N_24378,N_24677);
nor U29760 (N_29760,N_26092,N_24160);
nand U29761 (N_29761,N_26115,N_25971);
or U29762 (N_29762,N_24014,N_24037);
xnor U29763 (N_29763,N_25257,N_24299);
and U29764 (N_29764,N_26438,N_26974);
nand U29765 (N_29765,N_24454,N_25216);
or U29766 (N_29766,N_26697,N_26784);
or U29767 (N_29767,N_26468,N_26103);
or U29768 (N_29768,N_26107,N_25747);
nand U29769 (N_29769,N_25640,N_26591);
nand U29770 (N_29770,N_25508,N_25834);
nand U29771 (N_29771,N_24099,N_25854);
or U29772 (N_29772,N_24855,N_24923);
nor U29773 (N_29773,N_25126,N_24467);
nand U29774 (N_29774,N_24114,N_25259);
nand U29775 (N_29775,N_24352,N_25313);
and U29776 (N_29776,N_26662,N_24933);
or U29777 (N_29777,N_26429,N_26846);
xor U29778 (N_29778,N_26194,N_25650);
nand U29779 (N_29779,N_24648,N_26534);
xor U29780 (N_29780,N_24854,N_26860);
or U29781 (N_29781,N_26080,N_25747);
or U29782 (N_29782,N_25150,N_25514);
nor U29783 (N_29783,N_26336,N_25394);
or U29784 (N_29784,N_25652,N_26708);
xnor U29785 (N_29785,N_26595,N_24810);
xnor U29786 (N_29786,N_26271,N_24044);
nor U29787 (N_29787,N_24712,N_25891);
and U29788 (N_29788,N_26139,N_24151);
and U29789 (N_29789,N_24301,N_26924);
xor U29790 (N_29790,N_25058,N_25413);
nand U29791 (N_29791,N_24666,N_25872);
nor U29792 (N_29792,N_26000,N_24420);
or U29793 (N_29793,N_26726,N_24014);
nand U29794 (N_29794,N_25213,N_24905);
or U29795 (N_29795,N_26673,N_26356);
nor U29796 (N_29796,N_26604,N_26439);
nand U29797 (N_29797,N_25093,N_25872);
and U29798 (N_29798,N_26151,N_24011);
or U29799 (N_29799,N_26259,N_24649);
nor U29800 (N_29800,N_25603,N_26635);
or U29801 (N_29801,N_25288,N_25313);
nor U29802 (N_29802,N_25118,N_24242);
or U29803 (N_29803,N_24210,N_26837);
nand U29804 (N_29804,N_25029,N_26477);
nand U29805 (N_29805,N_25861,N_24830);
or U29806 (N_29806,N_25594,N_26352);
and U29807 (N_29807,N_26996,N_26531);
or U29808 (N_29808,N_24681,N_26254);
nor U29809 (N_29809,N_26619,N_26309);
nor U29810 (N_29810,N_24259,N_25421);
or U29811 (N_29811,N_25638,N_26910);
nand U29812 (N_29812,N_24804,N_24698);
or U29813 (N_29813,N_26973,N_24410);
nor U29814 (N_29814,N_25937,N_24154);
nor U29815 (N_29815,N_24657,N_24036);
xnor U29816 (N_29816,N_26911,N_24729);
or U29817 (N_29817,N_24929,N_24240);
or U29818 (N_29818,N_26151,N_24772);
nand U29819 (N_29819,N_25278,N_24155);
nand U29820 (N_29820,N_24595,N_24198);
xor U29821 (N_29821,N_25641,N_25020);
xnor U29822 (N_29822,N_24870,N_25044);
nand U29823 (N_29823,N_25617,N_26181);
nand U29824 (N_29824,N_26862,N_25258);
or U29825 (N_29825,N_26924,N_26199);
nand U29826 (N_29826,N_25370,N_25304);
nand U29827 (N_29827,N_25356,N_26471);
or U29828 (N_29828,N_25800,N_24448);
xnor U29829 (N_29829,N_25216,N_25503);
or U29830 (N_29830,N_24980,N_24384);
and U29831 (N_29831,N_26747,N_26912);
and U29832 (N_29832,N_26216,N_24790);
xor U29833 (N_29833,N_25687,N_24427);
nor U29834 (N_29834,N_25010,N_26661);
xnor U29835 (N_29835,N_24473,N_26955);
xnor U29836 (N_29836,N_24589,N_25860);
nand U29837 (N_29837,N_26963,N_24134);
or U29838 (N_29838,N_24522,N_26251);
or U29839 (N_29839,N_25911,N_26790);
or U29840 (N_29840,N_25330,N_25401);
and U29841 (N_29841,N_24132,N_24520);
nand U29842 (N_29842,N_24716,N_25538);
xor U29843 (N_29843,N_25030,N_25278);
nor U29844 (N_29844,N_24019,N_24971);
and U29845 (N_29845,N_26474,N_26730);
xor U29846 (N_29846,N_24540,N_26971);
nand U29847 (N_29847,N_26680,N_24217);
or U29848 (N_29848,N_25820,N_24825);
or U29849 (N_29849,N_26758,N_24314);
nand U29850 (N_29850,N_24461,N_26828);
and U29851 (N_29851,N_25278,N_24830);
nor U29852 (N_29852,N_26006,N_25512);
nand U29853 (N_29853,N_25309,N_25051);
nand U29854 (N_29854,N_26776,N_25618);
or U29855 (N_29855,N_25950,N_25935);
nand U29856 (N_29856,N_24981,N_26321);
and U29857 (N_29857,N_24844,N_26396);
xnor U29858 (N_29858,N_24825,N_24393);
xnor U29859 (N_29859,N_24232,N_24338);
nor U29860 (N_29860,N_24160,N_25551);
and U29861 (N_29861,N_26311,N_26780);
nor U29862 (N_29862,N_26301,N_24919);
xor U29863 (N_29863,N_24325,N_24134);
and U29864 (N_29864,N_26208,N_26250);
or U29865 (N_29865,N_25632,N_24540);
xor U29866 (N_29866,N_24070,N_26414);
xor U29867 (N_29867,N_25700,N_25941);
nor U29868 (N_29868,N_24476,N_26561);
xnor U29869 (N_29869,N_24994,N_25198);
xor U29870 (N_29870,N_24730,N_26449);
or U29871 (N_29871,N_24145,N_24058);
or U29872 (N_29872,N_26396,N_24614);
xor U29873 (N_29873,N_25104,N_25394);
xnor U29874 (N_29874,N_26740,N_26936);
xor U29875 (N_29875,N_26772,N_26358);
xor U29876 (N_29876,N_24280,N_25761);
nand U29877 (N_29877,N_24928,N_25471);
nand U29878 (N_29878,N_25816,N_25787);
nand U29879 (N_29879,N_25719,N_26485);
nor U29880 (N_29880,N_24662,N_25058);
nand U29881 (N_29881,N_26156,N_25820);
xor U29882 (N_29882,N_24013,N_26979);
nand U29883 (N_29883,N_24066,N_25115);
xnor U29884 (N_29884,N_24729,N_25357);
or U29885 (N_29885,N_26392,N_26180);
nand U29886 (N_29886,N_24310,N_25941);
and U29887 (N_29887,N_25402,N_25508);
nand U29888 (N_29888,N_25888,N_26989);
xor U29889 (N_29889,N_24045,N_26028);
or U29890 (N_29890,N_25891,N_25617);
or U29891 (N_29891,N_26692,N_24386);
and U29892 (N_29892,N_26347,N_25706);
nor U29893 (N_29893,N_26730,N_25515);
or U29894 (N_29894,N_25713,N_24232);
nand U29895 (N_29895,N_25761,N_24652);
nand U29896 (N_29896,N_26811,N_26332);
and U29897 (N_29897,N_24232,N_24712);
xnor U29898 (N_29898,N_26519,N_26604);
and U29899 (N_29899,N_25445,N_25257);
nand U29900 (N_29900,N_26032,N_25501);
nand U29901 (N_29901,N_24281,N_25622);
nor U29902 (N_29902,N_24793,N_25873);
and U29903 (N_29903,N_26338,N_24493);
or U29904 (N_29904,N_24474,N_25906);
and U29905 (N_29905,N_26384,N_24831);
xnor U29906 (N_29906,N_24664,N_26167);
xor U29907 (N_29907,N_26259,N_24430);
nand U29908 (N_29908,N_24029,N_24958);
xor U29909 (N_29909,N_25649,N_25745);
nor U29910 (N_29910,N_26226,N_24217);
nand U29911 (N_29911,N_25622,N_24915);
or U29912 (N_29912,N_26339,N_24030);
or U29913 (N_29913,N_26896,N_24643);
xor U29914 (N_29914,N_24105,N_26509);
xnor U29915 (N_29915,N_26714,N_24518);
and U29916 (N_29916,N_25366,N_24667);
xnor U29917 (N_29917,N_26773,N_24311);
or U29918 (N_29918,N_24477,N_25931);
or U29919 (N_29919,N_26710,N_24445);
nand U29920 (N_29920,N_25304,N_25897);
and U29921 (N_29921,N_25244,N_25904);
nor U29922 (N_29922,N_24154,N_24260);
xnor U29923 (N_29923,N_26138,N_26803);
or U29924 (N_29924,N_26223,N_25225);
nor U29925 (N_29925,N_24674,N_26013);
or U29926 (N_29926,N_25803,N_25733);
nor U29927 (N_29927,N_24289,N_24731);
nor U29928 (N_29928,N_26995,N_26275);
or U29929 (N_29929,N_24388,N_26303);
nand U29930 (N_29930,N_24496,N_26027);
or U29931 (N_29931,N_25591,N_25814);
xnor U29932 (N_29932,N_24522,N_25225);
nor U29933 (N_29933,N_26296,N_24662);
or U29934 (N_29934,N_26895,N_26352);
xnor U29935 (N_29935,N_26622,N_25444);
nor U29936 (N_29936,N_26727,N_25253);
nand U29937 (N_29937,N_26777,N_25705);
nor U29938 (N_29938,N_25669,N_24427);
nor U29939 (N_29939,N_25753,N_24624);
nand U29940 (N_29940,N_26263,N_25344);
or U29941 (N_29941,N_24666,N_24306);
nand U29942 (N_29942,N_24161,N_25218);
or U29943 (N_29943,N_26221,N_26411);
xor U29944 (N_29944,N_24541,N_24141);
and U29945 (N_29945,N_26921,N_24534);
nand U29946 (N_29946,N_24748,N_24956);
xnor U29947 (N_29947,N_25870,N_24440);
nor U29948 (N_29948,N_24343,N_26041);
or U29949 (N_29949,N_26061,N_24761);
or U29950 (N_29950,N_25019,N_24281);
or U29951 (N_29951,N_24887,N_25181);
xnor U29952 (N_29952,N_24074,N_25116);
and U29953 (N_29953,N_24854,N_25874);
nand U29954 (N_29954,N_25347,N_25978);
or U29955 (N_29955,N_26294,N_24757);
or U29956 (N_29956,N_25952,N_25614);
nand U29957 (N_29957,N_25052,N_24893);
nand U29958 (N_29958,N_24311,N_26951);
nor U29959 (N_29959,N_25936,N_26216);
xnor U29960 (N_29960,N_24404,N_24090);
xnor U29961 (N_29961,N_25339,N_24824);
or U29962 (N_29962,N_25756,N_24840);
and U29963 (N_29963,N_24907,N_26282);
or U29964 (N_29964,N_26489,N_26089);
or U29965 (N_29965,N_24693,N_26026);
nor U29966 (N_29966,N_24881,N_26400);
and U29967 (N_29967,N_24248,N_26242);
nor U29968 (N_29968,N_25800,N_25762);
nand U29969 (N_29969,N_24826,N_24958);
nand U29970 (N_29970,N_25601,N_25872);
xnor U29971 (N_29971,N_25019,N_25412);
and U29972 (N_29972,N_26216,N_26694);
or U29973 (N_29973,N_25176,N_26621);
nand U29974 (N_29974,N_26232,N_26003);
or U29975 (N_29975,N_26685,N_24414);
and U29976 (N_29976,N_24544,N_25431);
nand U29977 (N_29977,N_25610,N_24504);
nand U29978 (N_29978,N_25519,N_25632);
and U29979 (N_29979,N_24924,N_24197);
nand U29980 (N_29980,N_25156,N_25453);
nand U29981 (N_29981,N_26146,N_25967);
or U29982 (N_29982,N_24566,N_25798);
xor U29983 (N_29983,N_26803,N_26429);
nand U29984 (N_29984,N_25839,N_26309);
or U29985 (N_29985,N_24759,N_25334);
xnor U29986 (N_29986,N_24521,N_25041);
nand U29987 (N_29987,N_26624,N_25050);
or U29988 (N_29988,N_25116,N_26567);
nor U29989 (N_29989,N_24940,N_24068);
and U29990 (N_29990,N_24226,N_25616);
xnor U29991 (N_29991,N_26122,N_26763);
xor U29992 (N_29992,N_26426,N_25745);
nand U29993 (N_29993,N_26453,N_25413);
nand U29994 (N_29994,N_24985,N_25226);
xnor U29995 (N_29995,N_26272,N_24154);
and U29996 (N_29996,N_26713,N_25562);
or U29997 (N_29997,N_24712,N_25334);
nand U29998 (N_29998,N_24940,N_25503);
and U29999 (N_29999,N_25438,N_26745);
or UO_0 (O_0,N_29691,N_29213);
or UO_1 (O_1,N_27587,N_27524);
or UO_2 (O_2,N_29124,N_27371);
or UO_3 (O_3,N_27714,N_28264);
nor UO_4 (O_4,N_29052,N_29315);
xor UO_5 (O_5,N_28297,N_28279);
and UO_6 (O_6,N_28833,N_28242);
nand UO_7 (O_7,N_28337,N_27677);
xor UO_8 (O_8,N_27661,N_29741);
or UO_9 (O_9,N_28584,N_28054);
and UO_10 (O_10,N_27427,N_28785);
and UO_11 (O_11,N_27270,N_29833);
nor UO_12 (O_12,N_27618,N_27455);
and UO_13 (O_13,N_27144,N_28621);
or UO_14 (O_14,N_28257,N_27383);
nor UO_15 (O_15,N_29994,N_28805);
and UO_16 (O_16,N_27728,N_27035);
nand UO_17 (O_17,N_28952,N_29875);
xor UO_18 (O_18,N_27890,N_29851);
nor UO_19 (O_19,N_27279,N_28047);
nor UO_20 (O_20,N_29260,N_27411);
or UO_21 (O_21,N_27118,N_29822);
xnor UO_22 (O_22,N_28266,N_28495);
and UO_23 (O_23,N_29419,N_28650);
and UO_24 (O_24,N_28673,N_28608);
nand UO_25 (O_25,N_28413,N_28903);
nor UO_26 (O_26,N_27582,N_29918);
nand UO_27 (O_27,N_29548,N_28084);
or UO_28 (O_28,N_29420,N_28843);
and UO_29 (O_29,N_29271,N_28988);
nor UO_30 (O_30,N_29111,N_28512);
and UO_31 (O_31,N_28652,N_28271);
or UO_32 (O_32,N_28183,N_28565);
and UO_33 (O_33,N_27904,N_29495);
or UO_34 (O_34,N_27598,N_29214);
or UO_35 (O_35,N_28597,N_27401);
nor UO_36 (O_36,N_29900,N_27722);
xor UO_37 (O_37,N_27561,N_29434);
or UO_38 (O_38,N_27006,N_27562);
nand UO_39 (O_39,N_29142,N_29653);
nand UO_40 (O_40,N_29223,N_28760);
nor UO_41 (O_41,N_29464,N_29141);
nand UO_42 (O_42,N_27820,N_27123);
xor UO_43 (O_43,N_29863,N_28824);
nor UO_44 (O_44,N_28677,N_28301);
nor UO_45 (O_45,N_27177,N_27305);
nor UO_46 (O_46,N_27301,N_27647);
nor UO_47 (O_47,N_27718,N_27944);
xnor UO_48 (O_48,N_27130,N_28787);
xnor UO_49 (O_49,N_27005,N_28813);
nor UO_50 (O_50,N_29031,N_29683);
or UO_51 (O_51,N_28466,N_28114);
nand UO_52 (O_52,N_29428,N_27851);
nand UO_53 (O_53,N_27576,N_29184);
nand UO_54 (O_54,N_29583,N_29266);
nor UO_55 (O_55,N_27386,N_27135);
nor UO_56 (O_56,N_27726,N_28284);
or UO_57 (O_57,N_28001,N_28395);
and UO_58 (O_58,N_27671,N_28393);
and UO_59 (O_59,N_29856,N_28486);
or UO_60 (O_60,N_28851,N_29929);
and UO_61 (O_61,N_28801,N_29390);
or UO_62 (O_62,N_27655,N_27484);
nand UO_63 (O_63,N_29757,N_27020);
nor UO_64 (O_64,N_27772,N_27959);
xor UO_65 (O_65,N_27313,N_27507);
xor UO_66 (O_66,N_28921,N_28309);
and UO_67 (O_67,N_29640,N_27907);
or UO_68 (O_68,N_29762,N_29408);
and UO_69 (O_69,N_27656,N_28042);
xor UO_70 (O_70,N_27237,N_28141);
nand UO_71 (O_71,N_28070,N_29125);
nor UO_72 (O_72,N_27815,N_27175);
or UO_73 (O_73,N_27999,N_28751);
nor UO_74 (O_74,N_28000,N_29823);
nand UO_75 (O_75,N_27956,N_28446);
and UO_76 (O_76,N_28109,N_28954);
xor UO_77 (O_77,N_28991,N_29499);
nand UO_78 (O_78,N_28184,N_29054);
or UO_79 (O_79,N_29703,N_27824);
nor UO_80 (O_80,N_28553,N_29338);
nor UO_81 (O_81,N_27004,N_27509);
nand UO_82 (O_82,N_29983,N_29636);
nand UO_83 (O_83,N_29964,N_27056);
xnor UO_84 (O_84,N_27653,N_29944);
xnor UO_85 (O_85,N_29621,N_27148);
xor UO_86 (O_86,N_28769,N_27102);
nand UO_87 (O_87,N_27060,N_29884);
or UO_88 (O_88,N_28224,N_28657);
and UO_89 (O_89,N_29244,N_27865);
or UO_90 (O_90,N_29514,N_29759);
and UO_91 (O_91,N_29307,N_29505);
nand UO_92 (O_92,N_27300,N_28152);
and UO_93 (O_93,N_27188,N_29721);
xor UO_94 (O_94,N_28982,N_28962);
xor UO_95 (O_95,N_27402,N_28926);
nand UO_96 (O_96,N_29865,N_29614);
xnor UO_97 (O_97,N_27555,N_29180);
nor UO_98 (O_98,N_27965,N_29580);
nor UO_99 (O_99,N_29027,N_27725);
or UO_100 (O_100,N_28857,N_28905);
and UO_101 (O_101,N_27014,N_27558);
nor UO_102 (O_102,N_29398,N_29379);
or UO_103 (O_103,N_29360,N_28002);
nor UO_104 (O_104,N_29129,N_29200);
and UO_105 (O_105,N_27183,N_27713);
nand UO_106 (O_106,N_28401,N_27138);
nand UO_107 (O_107,N_27801,N_27500);
nand UO_108 (O_108,N_27443,N_28481);
nor UO_109 (O_109,N_29526,N_27040);
and UO_110 (O_110,N_28111,N_29253);
nand UO_111 (O_111,N_27275,N_29976);
or UO_112 (O_112,N_27365,N_28473);
nand UO_113 (O_113,N_27278,N_28093);
nor UO_114 (O_114,N_28747,N_29704);
xor UO_115 (O_115,N_27462,N_27117);
xnor UO_116 (O_116,N_27614,N_27053);
nor UO_117 (O_117,N_28499,N_27600);
nand UO_118 (O_118,N_29376,N_29527);
and UO_119 (O_119,N_28088,N_29662);
or UO_120 (O_120,N_28579,N_27033);
or UO_121 (O_121,N_29556,N_27591);
and UO_122 (O_122,N_28382,N_28804);
nand UO_123 (O_123,N_28668,N_28492);
nand UO_124 (O_124,N_29261,N_27634);
and UO_125 (O_125,N_28244,N_28333);
nor UO_126 (O_126,N_29279,N_27925);
xnor UO_127 (O_127,N_27882,N_28305);
or UO_128 (O_128,N_28339,N_27250);
nor UO_129 (O_129,N_29712,N_28549);
and UO_130 (O_130,N_28765,N_28731);
nand UO_131 (O_131,N_28231,N_27178);
or UO_132 (O_132,N_29224,N_29073);
nand UO_133 (O_133,N_27242,N_27556);
nor UO_134 (O_134,N_27215,N_29452);
and UO_135 (O_135,N_29101,N_29898);
nor UO_136 (O_136,N_28429,N_28159);
and UO_137 (O_137,N_29915,N_28104);
nand UO_138 (O_138,N_27276,N_29424);
and UO_139 (O_139,N_28326,N_29956);
nand UO_140 (O_140,N_29945,N_28927);
nor UO_141 (O_141,N_28161,N_29592);
xnor UO_142 (O_142,N_29008,N_27757);
nor UO_143 (O_143,N_27601,N_28080);
xor UO_144 (O_144,N_28236,N_27922);
nor UO_145 (O_145,N_29018,N_29620);
or UO_146 (O_146,N_28276,N_29332);
nand UO_147 (O_147,N_27560,N_28825);
or UO_148 (O_148,N_29845,N_27038);
xnor UO_149 (O_149,N_27982,N_29449);
and UO_150 (O_150,N_29631,N_28928);
nand UO_151 (O_151,N_28687,N_27977);
nand UO_152 (O_152,N_27011,N_28729);
and UO_153 (O_153,N_29385,N_27567);
nor UO_154 (O_154,N_29503,N_27075);
or UO_155 (O_155,N_27711,N_27165);
nand UO_156 (O_156,N_28533,N_29017);
xor UO_157 (O_157,N_28531,N_28253);
xnor UO_158 (O_158,N_27776,N_27180);
xor UO_159 (O_159,N_29046,N_29806);
nor UO_160 (O_160,N_28222,N_27819);
or UO_161 (O_161,N_28788,N_28459);
or UO_162 (O_162,N_29349,N_28237);
nand UO_163 (O_163,N_27830,N_29061);
nand UO_164 (O_164,N_29615,N_29730);
or UO_165 (O_165,N_27724,N_27638);
or UO_166 (O_166,N_28210,N_27346);
nand UO_167 (O_167,N_29597,N_27219);
nor UO_168 (O_168,N_27116,N_29751);
nand UO_169 (O_169,N_28756,N_28035);
nand UO_170 (O_170,N_29882,N_28853);
xor UO_171 (O_171,N_28269,N_28006);
nor UO_172 (O_172,N_28947,N_28427);
and UO_173 (O_173,N_27871,N_29827);
and UO_174 (O_174,N_29270,N_28873);
and UO_175 (O_175,N_28876,N_28270);
xor UO_176 (O_176,N_28475,N_28868);
nand UO_177 (O_177,N_29634,N_29909);
xor UO_178 (O_178,N_28559,N_27050);
nor UO_179 (O_179,N_28839,N_27248);
nand UO_180 (O_180,N_28248,N_29013);
xor UO_181 (O_181,N_27212,N_29747);
nand UO_182 (O_182,N_28955,N_28026);
or UO_183 (O_183,N_28700,N_29251);
xor UO_184 (O_184,N_27669,N_27062);
or UO_185 (O_185,N_29324,N_29230);
nor UO_186 (O_186,N_27626,N_29748);
and UO_187 (O_187,N_29248,N_29395);
nand UO_188 (O_188,N_29766,N_27810);
nor UO_189 (O_189,N_28912,N_29354);
nor UO_190 (O_190,N_27928,N_28987);
xnor UO_191 (O_191,N_27895,N_29645);
nor UO_192 (O_192,N_29880,N_27234);
or UO_193 (O_193,N_29439,N_27169);
or UO_194 (O_194,N_29919,N_29318);
nor UO_195 (O_195,N_28258,N_27423);
nor UO_196 (O_196,N_27641,N_28158);
xnor UO_197 (O_197,N_29300,N_27404);
nor UO_198 (O_198,N_27227,N_28591);
or UO_199 (O_199,N_28234,N_28706);
or UO_200 (O_200,N_28166,N_27852);
nor UO_201 (O_201,N_29557,N_28530);
xnor UO_202 (O_202,N_27208,N_29984);
nand UO_203 (O_203,N_28827,N_29082);
xor UO_204 (O_204,N_27262,N_27639);
xor UO_205 (O_205,N_28678,N_29688);
and UO_206 (O_206,N_28125,N_27095);
or UO_207 (O_207,N_28958,N_29134);
nor UO_208 (O_208,N_29859,N_29857);
nand UO_209 (O_209,N_29133,N_28064);
or UO_210 (O_210,N_27249,N_27196);
xnor UO_211 (O_211,N_27839,N_29701);
or UO_212 (O_212,N_29317,N_29559);
or UO_213 (O_213,N_27151,N_28315);
or UO_214 (O_214,N_29902,N_28145);
nand UO_215 (O_215,N_28594,N_27995);
and UO_216 (O_216,N_28208,N_27419);
nor UO_217 (O_217,N_29675,N_29576);
or UO_218 (O_218,N_28795,N_29835);
or UO_219 (O_219,N_28432,N_27485);
nor UO_220 (O_220,N_27741,N_27277);
xnor UO_221 (O_221,N_28993,N_28911);
xnor UO_222 (O_222,N_29654,N_28890);
nor UO_223 (O_223,N_28031,N_28770);
and UO_224 (O_224,N_29241,N_28017);
or UO_225 (O_225,N_29697,N_27777);
or UO_226 (O_226,N_29590,N_29016);
nor UO_227 (O_227,N_28773,N_27460);
and UO_228 (O_228,N_27894,N_27619);
xnor UO_229 (O_229,N_28891,N_27707);
xor UO_230 (O_230,N_27778,N_29734);
and UO_231 (O_231,N_29958,N_27044);
nor UO_232 (O_232,N_29686,N_27515);
xor UO_233 (O_233,N_28972,N_28346);
and UO_234 (O_234,N_28470,N_29276);
and UO_235 (O_235,N_27306,N_27043);
or UO_236 (O_236,N_28612,N_27461);
nor UO_237 (O_237,N_29713,N_27362);
xor UO_238 (O_238,N_27825,N_28592);
and UO_239 (O_239,N_29461,N_29905);
and UO_240 (O_240,N_27575,N_27803);
nand UO_241 (O_241,N_27831,N_27849);
and UO_242 (O_242,N_29245,N_27797);
xnor UO_243 (O_243,N_28938,N_29516);
and UO_244 (O_244,N_29342,N_28195);
nand UO_245 (O_245,N_29507,N_28904);
nor UO_246 (O_246,N_28013,N_28477);
xnor UO_247 (O_247,N_27288,N_28672);
nand UO_248 (O_248,N_27333,N_27037);
nor UO_249 (O_249,N_28915,N_27574);
nor UO_250 (O_250,N_28930,N_28771);
xnor UO_251 (O_251,N_27140,N_28377);
nor UO_252 (O_252,N_29015,N_29961);
and UO_253 (O_253,N_28860,N_27001);
and UO_254 (O_254,N_27263,N_29950);
or UO_255 (O_255,N_29034,N_28397);
nor UO_256 (O_256,N_27632,N_27246);
or UO_257 (O_257,N_28138,N_28659);
or UO_258 (O_258,N_29032,N_27773);
nor UO_259 (O_259,N_29109,N_27845);
nand UO_260 (O_260,N_29044,N_27498);
nand UO_261 (O_261,N_29108,N_27847);
nor UO_262 (O_262,N_27002,N_28670);
or UO_263 (O_263,N_29972,N_27459);
and UO_264 (O_264,N_29731,N_27602);
and UO_265 (O_265,N_28123,N_28286);
xnor UO_266 (O_266,N_27953,N_28307);
xor UO_267 (O_267,N_27727,N_27488);
nor UO_268 (O_268,N_28488,N_28216);
and UO_269 (O_269,N_29295,N_27069);
xor UO_270 (O_270,N_27914,N_28008);
xnor UO_271 (O_271,N_27723,N_28819);
nand UO_272 (O_272,N_27812,N_28455);
nor UO_273 (O_273,N_29409,N_28199);
or UO_274 (O_274,N_27566,N_28029);
or UO_275 (O_275,N_27088,N_28577);
nand UO_276 (O_276,N_27494,N_27265);
xor UO_277 (O_277,N_29227,N_29680);
or UO_278 (O_278,N_27829,N_29282);
nor UO_279 (O_279,N_29820,N_27047);
xnor UO_280 (O_280,N_29067,N_28228);
nand UO_281 (O_281,N_27370,N_28964);
xor UO_282 (O_282,N_29723,N_27395);
or UO_283 (O_283,N_27241,N_29425);
nand UO_284 (O_284,N_28960,N_27802);
nand UO_285 (O_285,N_29773,N_28130);
or UO_286 (O_286,N_28792,N_29739);
or UO_287 (O_287,N_29138,N_29676);
nor UO_288 (O_288,N_29630,N_28797);
and UO_289 (O_289,N_27125,N_29163);
xnor UO_290 (O_290,N_29301,N_27409);
xnor UO_291 (O_291,N_29089,N_27579);
or UO_292 (O_292,N_29176,N_27063);
nor UO_293 (O_293,N_29209,N_27407);
and UO_294 (O_294,N_28806,N_28015);
or UO_295 (O_295,N_29440,N_27673);
nand UO_296 (O_296,N_29429,N_27142);
xor UO_297 (O_297,N_27846,N_28067);
or UO_298 (O_298,N_29211,N_27164);
and UO_299 (O_299,N_29932,N_27372);
xnor UO_300 (O_300,N_29637,N_29491);
nand UO_301 (O_301,N_28388,N_28137);
or UO_302 (O_302,N_27924,N_28663);
or UO_303 (O_303,N_29040,N_28294);
nand UO_304 (O_304,N_27179,N_28011);
nor UO_305 (O_305,N_27912,N_27425);
nand UO_306 (O_306,N_29960,N_29164);
nor UO_307 (O_307,N_29831,N_27770);
or UO_308 (O_308,N_28415,N_29077);
nor UO_309 (O_309,N_28744,N_29647);
nor UO_310 (O_310,N_28906,N_28165);
nand UO_311 (O_311,N_27101,N_29033);
nand UO_312 (O_312,N_27692,N_28046);
or UO_313 (O_313,N_28572,N_27762);
nand UO_314 (O_314,N_29869,N_27059);
and UO_315 (O_315,N_28436,N_28734);
or UO_316 (O_316,N_28334,N_28518);
nand UO_317 (O_317,N_28803,N_28252);
and UO_318 (O_318,N_29152,N_29292);
nand UO_319 (O_319,N_27525,N_29225);
xnor UO_320 (O_320,N_29249,N_29707);
and UO_321 (O_321,N_29840,N_28779);
xor UO_322 (O_322,N_28398,N_27610);
nand UO_323 (O_323,N_28627,N_28025);
nand UO_324 (O_324,N_28027,N_29836);
nor UO_325 (O_325,N_27527,N_28528);
or UO_326 (O_326,N_28351,N_28999);
xor UO_327 (O_327,N_28335,N_28768);
or UO_328 (O_328,N_27704,N_27716);
nor UO_329 (O_329,N_28984,N_29838);
or UO_330 (O_330,N_27475,N_28738);
xor UO_331 (O_331,N_29584,N_27302);
nand UO_332 (O_332,N_29803,N_28794);
nor UO_333 (O_333,N_27049,N_29547);
and UO_334 (O_334,N_29727,N_27154);
nand UO_335 (O_335,N_29239,N_28665);
or UO_336 (O_336,N_29202,N_29981);
and UO_337 (O_337,N_28653,N_29980);
nand UO_338 (O_338,N_27683,N_29951);
or UO_339 (O_339,N_29462,N_28791);
nand UO_340 (O_340,N_28098,N_29215);
xor UO_341 (O_341,N_27256,N_28967);
nor UO_342 (O_342,N_28044,N_28696);
or UO_343 (O_343,N_29510,N_28190);
and UO_344 (O_344,N_28556,N_29387);
nor UO_345 (O_345,N_29603,N_29834);
nor UO_346 (O_346,N_27315,N_28702);
or UO_347 (O_347,N_28444,N_29885);
xnor UO_348 (O_348,N_28884,N_29776);
nor UO_349 (O_349,N_28327,N_29316);
xor UO_350 (O_350,N_28290,N_28676);
nor UO_351 (O_351,N_27392,N_28133);
nand UO_352 (O_352,N_27768,N_29029);
nor UO_353 (O_353,N_29007,N_28213);
and UO_354 (O_354,N_27406,N_27875);
xnor UO_355 (O_355,N_29830,N_28866);
nand UO_356 (O_356,N_28010,N_27205);
nand UO_357 (O_357,N_29183,N_27563);
nor UO_358 (O_358,N_28423,N_27921);
xor UO_359 (O_359,N_28420,N_28838);
xor UO_360 (O_360,N_27644,N_29002);
or UO_361 (O_361,N_29302,N_27862);
or UO_362 (O_362,N_27472,N_28725);
and UO_363 (O_363,N_27139,N_27285);
xnor UO_364 (O_364,N_29805,N_27152);
and UO_365 (O_365,N_29372,N_27899);
nor UO_366 (O_366,N_27480,N_28522);
nor UO_367 (O_367,N_29575,N_28187);
nand UO_368 (O_368,N_27085,N_27200);
nor UO_369 (O_369,N_29255,N_27431);
nor UO_370 (O_370,N_29888,N_29622);
xor UO_371 (O_371,N_27997,N_28447);
and UO_372 (O_372,N_27676,N_29383);
nand UO_373 (O_373,N_28818,N_27583);
nor UO_374 (O_374,N_27304,N_27568);
nor UO_375 (O_375,N_27450,N_27963);
or UO_376 (O_376,N_28360,N_28753);
nor UO_377 (O_377,N_28356,N_29336);
and UO_378 (O_378,N_28135,N_27821);
or UO_379 (O_379,N_29524,N_28886);
xor UO_380 (O_380,N_29188,N_28578);
nor UO_381 (O_381,N_27606,N_27690);
and UO_382 (O_382,N_29598,N_27366);
nand UO_383 (O_383,N_29199,N_29296);
xnor UO_384 (O_384,N_28235,N_29472);
xor UO_385 (O_385,N_28471,N_29485);
or UO_386 (O_386,N_29737,N_27887);
or UO_387 (O_387,N_28521,N_27487);
nor UO_388 (O_388,N_28453,N_29346);
or UO_389 (O_389,N_29482,N_29581);
xor UO_390 (O_390,N_27897,N_29504);
or UO_391 (O_391,N_29413,N_28358);
nand UO_392 (O_392,N_28885,N_27906);
xor UO_393 (O_393,N_29517,N_29114);
nor UO_394 (O_394,N_27238,N_28586);
or UO_395 (O_395,N_27900,N_29502);
or UO_396 (O_396,N_29924,N_28004);
xnor UO_397 (O_397,N_27627,N_28003);
nand UO_398 (O_398,N_28889,N_29521);
or UO_399 (O_399,N_28124,N_29605);
and UO_400 (O_400,N_28349,N_29070);
and UO_401 (O_401,N_28451,N_27788);
and UO_402 (O_402,N_28116,N_29969);
nor UO_403 (O_403,N_28864,N_27573);
nor UO_404 (O_404,N_29309,N_29750);
and UO_405 (O_405,N_29810,N_28063);
nor UO_406 (O_406,N_27390,N_27964);
xor UO_407 (O_407,N_28859,N_28538);
xnor UO_408 (O_408,N_28980,N_28511);
xor UO_409 (O_409,N_28754,N_27808);
nor UO_410 (O_410,N_28778,N_28879);
and UO_411 (O_411,N_29147,N_28632);
nor UO_412 (O_412,N_29374,N_29140);
nand UO_413 (O_413,N_29732,N_28932);
xor UO_414 (O_414,N_27732,N_29438);
and UO_415 (O_415,N_29846,N_27469);
and UO_416 (O_416,N_27268,N_28185);
xnor UO_417 (O_417,N_27132,N_27544);
nand UO_418 (O_418,N_27156,N_27994);
and UO_419 (O_419,N_27605,N_27811);
nand UO_420 (O_420,N_28445,N_27709);
and UO_421 (O_421,N_27961,N_29198);
or UO_422 (O_422,N_28310,N_27584);
nand UO_423 (O_423,N_29635,N_27519);
and UO_424 (O_424,N_28498,N_27415);
nor UO_425 (O_425,N_27933,N_29555);
nand UO_426 (O_426,N_29916,N_27223);
nand UO_427 (O_427,N_28350,N_27160);
nor UO_428 (O_428,N_28361,N_27341);
xor UO_429 (O_429,N_29794,N_29967);
xor UO_430 (O_430,N_27616,N_29871);
and UO_431 (O_431,N_27720,N_29541);
nor UO_432 (O_432,N_28265,N_29802);
xor UO_433 (O_433,N_27211,N_29025);
xnor UO_434 (O_434,N_27010,N_27785);
or UO_435 (O_435,N_28332,N_27297);
nand UO_436 (O_436,N_27027,N_28534);
nand UO_437 (O_437,N_28649,N_27592);
xor UO_438 (O_438,N_27335,N_27946);
nand UO_439 (O_439,N_27076,N_28331);
nand UO_440 (O_440,N_28941,N_28923);
nand UO_441 (O_441,N_28723,N_27079);
nor UO_442 (O_442,N_27859,N_29287);
and UO_443 (O_443,N_27712,N_28571);
and UO_444 (O_444,N_27945,N_28776);
xnor UO_445 (O_445,N_28681,N_29048);
nand UO_446 (O_446,N_28251,N_27310);
nor UO_447 (O_447,N_29157,N_28272);
nand UO_448 (O_448,N_27684,N_27284);
nor UO_449 (O_449,N_27837,N_28014);
and UO_450 (O_450,N_27503,N_27700);
xnor UO_451 (O_451,N_29811,N_29378);
nor UO_452 (O_452,N_29761,N_29446);
nor UO_453 (O_453,N_28516,N_27464);
or UO_454 (O_454,N_29797,N_29359);
nor UO_455 (O_455,N_27572,N_28274);
nor UO_456 (O_456,N_28296,N_28041);
nand UO_457 (O_457,N_28142,N_29971);
and UO_458 (O_458,N_29953,N_29549);
and UO_459 (O_459,N_27195,N_28507);
nand UO_460 (O_460,N_29185,N_27112);
or UO_461 (O_461,N_28916,N_28981);
nor UO_462 (O_462,N_27129,N_29130);
nor UO_463 (O_463,N_27753,N_27446);
nand UO_464 (O_464,N_27696,N_28686);
and UO_465 (O_465,N_27954,N_27721);
nor UO_466 (O_466,N_27388,N_28600);
or UO_467 (O_467,N_28467,N_29341);
nand UO_468 (O_468,N_28345,N_29088);
xnor UO_469 (O_469,N_29277,N_27240);
or UO_470 (O_470,N_29232,N_29456);
and UO_471 (O_471,N_27209,N_28176);
xnor UO_472 (O_472,N_27141,N_28073);
nor UO_473 (O_473,N_27182,N_27643);
xnor UO_474 (O_474,N_29186,N_29267);
nor UO_475 (O_475,N_28633,N_28448);
and UO_476 (O_476,N_27717,N_29386);
and UO_477 (O_477,N_28287,N_28811);
xor UO_478 (O_478,N_28363,N_27795);
nand UO_479 (O_479,N_29441,N_27437);
xnor UO_480 (O_480,N_29263,N_27735);
nand UO_481 (O_481,N_28077,N_29347);
or UO_482 (O_482,N_27084,N_29219);
nor UO_483 (O_483,N_29451,N_29756);
and UO_484 (O_484,N_28799,N_29254);
nor UO_485 (O_485,N_29700,N_29753);
and UO_486 (O_486,N_28157,N_27630);
or UO_487 (O_487,N_29722,N_27400);
or UO_488 (O_488,N_28148,N_28091);
xor UO_489 (O_489,N_29045,N_28683);
xnor UO_490 (O_490,N_28246,N_29786);
xor UO_491 (O_491,N_27942,N_29936);
nor UO_492 (O_492,N_29407,N_27320);
or UO_493 (O_493,N_29377,N_29238);
nor UO_494 (O_494,N_27100,N_29926);
nor UO_495 (O_495,N_27216,N_28666);
or UO_496 (O_496,N_27686,N_28996);
and UO_497 (O_497,N_27586,N_29619);
nand UO_498 (O_498,N_28581,N_28871);
and UO_499 (O_499,N_28709,N_27911);
nor UO_500 (O_500,N_29659,N_29974);
nand UO_501 (O_501,N_27330,N_28800);
or UO_502 (O_502,N_27949,N_29864);
and UO_503 (O_503,N_27477,N_29458);
nor UO_504 (O_504,N_27444,N_27071);
nor UO_505 (O_505,N_27546,N_28865);
and UO_506 (O_506,N_29729,N_27985);
xnor UO_507 (O_507,N_29911,N_27660);
or UO_508 (O_508,N_27976,N_27291);
or UO_509 (O_509,N_29079,N_28715);
and UO_510 (O_510,N_27134,N_29459);
and UO_511 (O_511,N_27491,N_28841);
or UO_512 (O_512,N_27375,N_29004);
and UO_513 (O_513,N_28587,N_29197);
or UO_514 (O_514,N_28400,N_29841);
nor UO_515 (O_515,N_29305,N_29038);
nor UO_516 (O_516,N_28520,N_28362);
nand UO_517 (O_517,N_27067,N_28658);
nor UO_518 (O_518,N_27870,N_29664);
or UO_519 (O_519,N_29115,N_27892);
xnor UO_520 (O_520,N_27805,N_27046);
nand UO_521 (O_521,N_27841,N_27951);
nor UO_522 (O_522,N_29787,N_27162);
nor UO_523 (O_523,N_27744,N_28551);
nor UO_524 (O_524,N_29370,N_29627);
and UO_525 (O_525,N_28948,N_27645);
nor UO_526 (O_526,N_27421,N_28379);
or UO_527 (O_527,N_28376,N_29481);
xnor UO_528 (O_528,N_29062,N_29629);
xor UO_529 (O_529,N_27939,N_28394);
xor UO_530 (O_530,N_27974,N_28082);
xnor UO_531 (O_531,N_29511,N_29611);
xnor UO_532 (O_532,N_28880,N_29616);
xor UO_533 (O_533,N_27203,N_27971);
and UO_534 (O_534,N_27570,N_28758);
nor UO_535 (O_535,N_29358,N_28226);
nor UO_536 (O_536,N_29993,N_28783);
nand UO_537 (O_537,N_28278,N_28324);
xor UO_538 (O_538,N_27025,N_29177);
or UO_539 (O_539,N_28695,N_27633);
nand UO_540 (O_540,N_28690,N_27023);
xor UO_541 (O_541,N_27853,N_29804);
and UO_542 (O_542,N_29283,N_29384);
xor UO_543 (O_543,N_28497,N_29626);
and UO_544 (O_544,N_29718,N_28878);
or UO_545 (O_545,N_27512,N_27978);
nand UO_546 (O_546,N_29633,N_29512);
and UO_547 (O_547,N_29135,N_29962);
xnor UO_548 (O_548,N_29807,N_29763);
or UO_549 (O_549,N_28603,N_27590);
nand UO_550 (O_550,N_29433,N_29705);
nor UO_551 (O_551,N_29923,N_27185);
xor UO_552 (O_552,N_29415,N_27345);
xnor UO_553 (O_553,N_28966,N_28131);
nor UO_554 (O_554,N_29954,N_29174);
xnor UO_555 (O_555,N_29706,N_27064);
or UO_556 (O_556,N_28348,N_27622);
nand UO_557 (O_557,N_27765,N_28986);
nor UO_558 (O_558,N_29131,N_28150);
nor UO_559 (O_559,N_29881,N_28173);
xor UO_560 (O_560,N_28625,N_29946);
xnor UO_561 (O_561,N_28206,N_28007);
xor UO_562 (O_562,N_28721,N_27247);
xnor UO_563 (O_563,N_29353,N_28068);
nand UO_564 (O_564,N_28468,N_29784);
xor UO_565 (O_565,N_27319,N_28403);
or UO_566 (O_566,N_27779,N_29677);
and UO_567 (O_567,N_29818,N_29998);
or UO_568 (O_568,N_28842,N_27880);
xor UO_569 (O_569,N_28204,N_27932);
nand UO_570 (O_570,N_27207,N_29042);
nor UO_571 (O_571,N_27662,N_28946);
nand UO_572 (O_572,N_28043,N_28221);
xnor UO_573 (O_573,N_28117,N_28040);
and UO_574 (O_574,N_29159,N_29985);
nor UO_575 (O_575,N_28215,N_29323);
and UO_576 (O_576,N_29085,N_27257);
xnor UO_577 (O_577,N_28896,N_27642);
nand UO_578 (O_578,N_28645,N_29883);
or UO_579 (O_579,N_27896,N_28934);
or UO_580 (O_580,N_29093,N_27414);
and UO_581 (O_581,N_27432,N_27885);
or UO_582 (O_582,N_27474,N_29474);
or UO_583 (O_583,N_29136,N_28611);
and UO_584 (O_584,N_27452,N_29742);
xnor UO_585 (O_585,N_27528,N_29933);
or UO_586 (O_586,N_27595,N_28939);
nand UO_587 (O_587,N_27454,N_28422);
xor UO_588 (O_588,N_27730,N_27624);
xor UO_589 (O_589,N_28302,N_28583);
nand UO_590 (O_590,N_29858,N_28273);
and UO_591 (O_591,N_27199,N_27547);
or UO_592 (O_592,N_27344,N_27508);
and UO_593 (O_593,N_27133,N_27781);
xnor UO_594 (O_594,N_29080,N_29417);
xnor UO_595 (O_595,N_28519,N_29448);
or UO_596 (O_596,N_27394,N_28629);
nand UO_597 (O_597,N_28132,N_28523);
and UO_598 (O_598,N_27695,N_28097);
or UO_599 (O_599,N_27137,N_28990);
nand UO_600 (O_600,N_28740,N_27008);
xor UO_601 (O_601,N_28711,N_28389);
xnor UO_602 (O_602,N_28536,N_29442);
xnor UO_603 (O_603,N_27338,N_29935);
or UO_604 (O_604,N_28328,N_29165);
and UO_605 (O_605,N_29201,N_28160);
nand UO_606 (O_606,N_29890,N_29308);
or UO_607 (O_607,N_28317,N_29127);
and UO_608 (O_608,N_27863,N_29816);
and UO_609 (O_609,N_27523,N_28410);
xnor UO_610 (O_610,N_27998,N_27814);
and UO_611 (O_611,N_29561,N_28940);
or UO_612 (O_612,N_29047,N_28951);
xnor UO_613 (O_613,N_27149,N_27749);
and UO_614 (O_614,N_27081,N_27530);
nand UO_615 (O_615,N_29119,N_27280);
nor UO_616 (O_616,N_27264,N_29815);
xnor UO_617 (O_617,N_27289,N_27941);
xor UO_618 (O_618,N_28589,N_29542);
and UO_619 (O_619,N_29679,N_28685);
and UO_620 (O_620,N_27981,N_27792);
and UO_621 (O_621,N_29934,N_27550);
xnor UO_622 (O_622,N_27731,N_29060);
xnor UO_623 (O_623,N_27364,N_28012);
or UO_624 (O_624,N_29872,N_27516);
nand UO_625 (O_625,N_29084,N_27860);
nor UO_626 (O_626,N_27658,N_29011);
nand UO_627 (O_627,N_29043,N_27988);
and UO_628 (O_628,N_28207,N_29656);
and UO_629 (O_629,N_27571,N_27518);
or UO_630 (O_630,N_28083,N_28956);
xor UO_631 (O_631,N_29367,N_29735);
and UO_632 (O_632,N_29774,N_29265);
or UO_633 (O_633,N_28169,N_28655);
nand UO_634 (O_634,N_28718,N_28807);
nand UO_635 (O_635,N_28739,N_27434);
nor UO_636 (O_636,N_29252,N_28823);
xnor UO_637 (O_637,N_29887,N_27197);
xnor UO_638 (O_638,N_29798,N_27352);
xor UO_639 (O_639,N_28622,N_28781);
or UO_640 (O_640,N_27670,N_28917);
xnor UO_641 (O_641,N_29105,N_28682);
nor UO_642 (O_642,N_27103,N_27126);
and UO_643 (O_643,N_27314,N_28599);
and UO_644 (O_644,N_29515,N_27226);
or UO_645 (O_645,N_28836,N_27858);
and UO_646 (O_646,N_27426,N_27379);
and UO_647 (O_647,N_28874,N_28129);
xor UO_648 (O_648,N_27840,N_29365);
and UO_649 (O_649,N_28974,N_29059);
or UO_650 (O_650,N_28809,N_28193);
xnor UO_651 (O_651,N_29427,N_27332);
nor UO_652 (O_652,N_27201,N_28852);
nor UO_653 (O_653,N_27466,N_28689);
nor UO_654 (O_654,N_29997,N_28513);
xor UO_655 (O_655,N_29824,N_29613);
nor UO_656 (O_656,N_27283,N_29169);
xor UO_657 (O_657,N_28254,N_28961);
and UO_658 (O_658,N_28719,N_27834);
or UO_659 (O_659,N_28626,N_27329);
nand UO_660 (O_660,N_28557,N_28604);
nor UO_661 (O_661,N_27748,N_28717);
xor UO_662 (O_662,N_29001,N_29591);
or UO_663 (O_663,N_27649,N_28094);
xnor UO_664 (O_664,N_28056,N_29450);
xor UO_665 (O_665,N_27024,N_27521);
nor UO_666 (O_666,N_27496,N_28240);
nand UO_667 (O_667,N_27456,N_29913);
xor UO_668 (O_668,N_29544,N_28661);
and UO_669 (O_669,N_28694,N_27473);
and UO_670 (O_670,N_27052,N_29123);
and UO_671 (O_671,N_27155,N_27159);
nor UO_672 (O_672,N_28679,N_28793);
nor UO_673 (O_673,N_28298,N_28209);
nor UO_674 (O_674,N_28935,N_28933);
nor UO_675 (O_675,N_29530,N_27886);
nor UO_676 (O_676,N_28197,N_27096);
nand UO_677 (O_677,N_28798,N_27955);
nor UO_678 (O_678,N_29853,N_27232);
and UO_679 (O_679,N_28121,N_29930);
or UO_680 (O_680,N_29196,N_29486);
nor UO_681 (O_681,N_28487,N_29178);
or UO_682 (O_682,N_29494,N_29335);
xor UO_683 (O_683,N_27340,N_28113);
nor UO_684 (O_684,N_29465,N_27317);
and UO_685 (O_685,N_27397,N_28406);
nor UO_686 (O_686,N_28179,N_27510);
nor UO_687 (O_687,N_27844,N_28493);
nor UO_688 (O_688,N_28802,N_29212);
and UO_689 (O_689,N_27124,N_27176);
nor UO_690 (O_690,N_27490,N_28110);
xnor UO_691 (O_691,N_28708,N_27073);
and UO_692 (O_692,N_27481,N_27121);
nand UO_693 (O_693,N_27698,N_29468);
xor UO_694 (O_694,N_28218,N_27294);
and UO_695 (O_695,N_28052,N_29010);
xnor UO_696 (O_696,N_27356,N_28503);
nand UO_697 (O_697,N_29912,N_28075);
nand UO_698 (O_698,N_27299,N_28628);
xnor UO_699 (O_699,N_28742,N_27664);
and UO_700 (O_700,N_28136,N_29259);
and UO_701 (O_701,N_28038,N_27536);
nor UO_702 (O_702,N_28407,N_29435);
or UO_703 (O_703,N_28992,N_29155);
xor UO_704 (O_704,N_27222,N_29992);
or UO_705 (O_705,N_29286,N_29350);
and UO_706 (O_706,N_27710,N_28598);
xor UO_707 (O_707,N_29848,N_28680);
or UO_708 (O_708,N_27514,N_29800);
and UO_709 (O_709,N_29120,N_27127);
or UO_710 (O_710,N_27220,N_28402);
nand UO_711 (O_711,N_27057,N_27763);
nand UO_712 (O_712,N_27621,N_28045);
nor UO_713 (O_713,N_28454,N_29696);
and UO_714 (O_714,N_28812,N_29366);
nand UO_715 (O_715,N_27361,N_28555);
nand UO_716 (O_716,N_27565,N_27357);
xnor UO_717 (O_717,N_29709,N_28736);
nand UO_718 (O_718,N_29596,N_28637);
and UO_719 (O_719,N_28460,N_27486);
nand UO_720 (O_720,N_28537,N_29782);
nor UO_721 (O_721,N_27187,N_29273);
and UO_722 (O_722,N_27325,N_29719);
xnor UO_723 (O_723,N_29564,N_28909);
nor UO_724 (O_724,N_29860,N_28737);
or UO_725 (O_725,N_27766,N_28535);
nand UO_726 (O_726,N_27041,N_27729);
and UO_727 (O_727,N_29380,N_28200);
and UO_728 (O_728,N_27992,N_29455);
and UO_729 (O_729,N_29097,N_27842);
or UO_730 (O_730,N_28018,N_28399);
nand UO_731 (O_731,N_29179,N_29650);
or UO_732 (O_732,N_29828,N_28312);
and UO_733 (O_733,N_28569,N_27952);
or UO_734 (O_734,N_29910,N_29496);
and UO_735 (O_735,N_29339,N_28699);
xor UO_736 (O_736,N_27967,N_29081);
or UO_737 (O_737,N_28634,N_27635);
xnor UO_738 (O_738,N_29103,N_27708);
or UO_739 (O_739,N_28178,N_28280);
or UO_740 (O_740,N_29019,N_28201);
or UO_741 (O_741,N_28338,N_27734);
and UO_742 (O_742,N_29588,N_28684);
or UO_743 (O_743,N_28139,N_28034);
nor UO_744 (O_744,N_29189,N_29938);
or UO_745 (O_745,N_28203,N_27739);
and UO_746 (O_746,N_28566,N_28442);
nand UO_747 (O_747,N_27109,N_29226);
or UO_748 (O_748,N_29728,N_28354);
xnor UO_749 (O_749,N_29897,N_27009);
nand UO_750 (O_750,N_28750,N_29531);
xnor UO_751 (O_751,N_29778,N_28863);
nand UO_752 (O_752,N_28283,N_27360);
nand UO_753 (O_753,N_29149,N_29190);
xor UO_754 (O_754,N_28192,N_27687);
or UO_755 (O_755,N_27968,N_28112);
or UO_756 (O_756,N_29285,N_28066);
xor UO_757 (O_757,N_28844,N_27433);
xor UO_758 (O_758,N_27483,N_28289);
or UO_759 (O_759,N_29063,N_27191);
or UO_760 (O_760,N_27261,N_27094);
nor UO_761 (O_761,N_28970,N_27077);
nor UO_762 (O_762,N_27213,N_28100);
or UO_763 (O_763,N_29567,N_29978);
xor UO_764 (O_764,N_27086,N_27902);
xnor UO_765 (O_765,N_27682,N_28546);
nand UO_766 (O_766,N_27915,N_27378);
xor UO_767 (O_767,N_28463,N_29382);
xnor UO_768 (O_768,N_27607,N_28456);
nor UO_769 (O_769,N_29608,N_29546);
nor UO_770 (O_770,N_29973,N_27585);
xnor UO_771 (O_771,N_29306,N_29536);
or UO_772 (O_772,N_29970,N_27048);
or UO_773 (O_773,N_27937,N_27893);
nor UO_774 (O_774,N_28259,N_29218);
nand UO_775 (O_775,N_27428,N_27657);
or UO_776 (O_776,N_27150,N_27935);
and UO_777 (O_777,N_27693,N_29543);
nand UO_778 (O_778,N_27580,N_29995);
and UO_779 (O_779,N_28156,N_29112);
and UO_780 (O_780,N_28945,N_29553);
or UO_781 (O_781,N_28989,N_28120);
nand UO_782 (O_782,N_29290,N_28189);
and UO_783 (O_783,N_29565,N_29699);
nor UO_784 (O_784,N_27445,N_27628);
nor UO_785 (O_785,N_28250,N_29725);
or UO_786 (O_786,N_28963,N_28570);
nand UO_787 (O_787,N_29612,N_28233);
xnor UO_788 (O_788,N_28509,N_27608);
and UO_789 (O_789,N_28378,N_29217);
nor UO_790 (O_790,N_29411,N_28767);
or UO_791 (O_791,N_27504,N_28457);
or UO_792 (O_792,N_29667,N_27553);
nor UO_793 (O_793,N_29394,N_27526);
and UO_794 (O_794,N_29023,N_29602);
nand UO_795 (O_795,N_27243,N_29221);
nand UO_796 (O_796,N_28277,N_28205);
and UO_797 (O_797,N_28144,N_28845);
and UO_798 (O_798,N_28443,N_29825);
nand UO_799 (O_799,N_27679,N_28167);
nor UO_800 (O_800,N_28472,N_29403);
or UO_801 (O_801,N_27835,N_27136);
nand UO_802 (O_802,N_27685,N_29371);
nor UO_803 (O_803,N_27791,N_27522);
nor UO_804 (O_804,N_28032,N_29893);
xnor UO_805 (O_805,N_28730,N_28716);
nor UO_806 (O_806,N_28898,N_28211);
or UO_807 (O_807,N_27429,N_27339);
xor UO_808 (O_808,N_28848,N_29508);
nand UO_809 (O_809,N_27564,N_28452);
nor UO_810 (O_810,N_29098,N_28675);
and UO_811 (O_811,N_28162,N_29470);
nand UO_812 (O_812,N_28057,N_27258);
and UO_813 (O_813,N_28059,N_29162);
nor UO_814 (O_814,N_27623,N_29673);
nand UO_815 (O_815,N_28899,N_27438);
and UO_816 (O_816,N_29191,N_29388);
and UO_817 (O_817,N_29589,N_29710);
or UO_818 (O_818,N_28560,N_28311);
nor UO_819 (O_819,N_29765,N_28942);
xor UO_820 (O_820,N_28636,N_29375);
and UO_821 (O_821,N_27244,N_27453);
nor UO_822 (O_822,N_29839,N_29095);
nand UO_823 (O_823,N_27021,N_27822);
xor UO_824 (O_824,N_29401,N_27989);
nor UO_825 (O_825,N_29574,N_28548);
or UO_826 (O_826,N_29143,N_29116);
nor UO_827 (O_827,N_29132,N_28796);
nand UO_828 (O_828,N_27252,N_27737);
nand UO_829 (O_829,N_29595,N_27236);
and UO_830 (O_830,N_27435,N_28275);
xnor UO_831 (O_831,N_29003,N_27688);
nor UO_832 (O_832,N_27702,N_27774);
nand UO_833 (O_833,N_28504,N_28180);
xnor UO_834 (O_834,N_27163,N_28194);
xnor UO_835 (O_835,N_29792,N_28784);
nand UO_836 (O_836,N_27254,N_29418);
or UO_837 (O_837,N_27599,N_28417);
or UO_838 (O_838,N_28922,N_29651);
and UO_839 (O_839,N_29861,N_29453);
xor UO_840 (O_840,N_28671,N_29518);
nand UO_841 (O_841,N_27224,N_27548);
nand UO_842 (O_842,N_27157,N_28883);
or UO_843 (O_843,N_29256,N_29257);
nor UO_844 (O_844,N_29154,N_27348);
nor UO_845 (O_845,N_28016,N_27396);
nand UO_846 (O_846,N_27030,N_27680);
nor UO_847 (O_847,N_27016,N_29866);
and UO_848 (O_848,N_28295,N_28808);
xnor UO_849 (O_849,N_29966,N_28418);
or UO_850 (O_850,N_28810,N_28892);
and UO_851 (O_851,N_29092,N_27767);
xnor UO_852 (O_852,N_29684,N_29783);
nand UO_853 (O_853,N_29641,N_27996);
xor UO_854 (O_854,N_29069,N_29573);
nand UO_855 (O_855,N_28691,N_28667);
and UO_856 (O_856,N_27328,N_27420);
or UO_857 (O_857,N_27093,N_28118);
nand UO_858 (O_858,N_27761,N_29229);
nand UO_859 (O_859,N_27045,N_29126);
xor UO_860 (O_860,N_27266,N_29362);
nor UO_861 (O_861,N_27309,N_28367);
and UO_862 (O_862,N_29208,N_28728);
nand UO_863 (O_863,N_29724,N_27648);
xnor UO_864 (O_864,N_27520,N_27376);
nor UO_865 (O_865,N_29566,N_29799);
or UO_866 (O_866,N_29182,N_29012);
and UO_867 (O_867,N_29203,N_29422);
nor UO_868 (O_868,N_27983,N_29161);
and UO_869 (O_869,N_27323,N_28186);
nand UO_870 (O_870,N_27569,N_29304);
xor UO_871 (O_871,N_29554,N_29801);
or UO_872 (O_872,N_28355,N_27296);
and UO_873 (O_873,N_29432,N_29231);
nand UO_874 (O_874,N_27119,N_28820);
nand UO_875 (O_875,N_27771,N_27541);
nor UO_876 (O_876,N_29666,N_29600);
nor UO_877 (O_877,N_28450,N_29170);
nand UO_878 (O_878,N_27879,N_27281);
nor UO_879 (O_879,N_29144,N_28641);
and UO_880 (O_880,N_27543,N_29572);
and UO_881 (O_881,N_28527,N_29687);
nand UO_882 (O_882,N_29228,N_27013);
nor UO_883 (O_883,N_27715,N_28726);
nand UO_884 (O_884,N_27405,N_28202);
nor UO_885 (O_885,N_29035,N_29074);
xnor UO_886 (O_886,N_28030,N_29195);
nand UO_887 (O_887,N_27874,N_29873);
and UO_888 (O_888,N_29483,N_27823);
nand UO_889 (O_889,N_27173,N_29443);
and UO_890 (O_890,N_27758,N_27318);
or UO_891 (O_891,N_27854,N_29205);
xnor UO_892 (O_892,N_28483,N_28968);
nand UO_893 (O_893,N_28081,N_28255);
or UO_894 (O_894,N_28256,N_27864);
or UO_895 (O_895,N_27221,N_29829);
nor UO_896 (O_896,N_27307,N_29955);
and UO_897 (O_897,N_28720,N_27936);
or UO_898 (O_898,N_27681,N_27993);
nand UO_899 (O_899,N_27827,N_28605);
or UO_900 (O_900,N_29087,N_29624);
nand UO_901 (O_901,N_27233,N_27979);
or UO_902 (O_902,N_29570,N_27350);
nor UO_903 (O_903,N_28815,N_29837);
xor UO_904 (O_904,N_29310,N_27637);
nor UO_905 (O_905,N_27106,N_27678);
nand UO_906 (O_906,N_27636,N_27986);
nor UO_907 (O_907,N_29181,N_29039);
xor UO_908 (O_908,N_27269,N_29854);
xnor UO_909 (O_909,N_27168,N_27058);
nand UO_910 (O_910,N_28541,N_27917);
nand UO_911 (O_911,N_27082,N_27447);
and UO_912 (O_912,N_28745,N_28821);
xnor UO_913 (O_913,N_27012,N_27408);
xnor UO_914 (O_914,N_29236,N_28370);
or UO_915 (O_915,N_29331,N_27374);
xnor UO_916 (O_916,N_27113,N_27966);
and UO_917 (O_917,N_27051,N_28421);
xor UO_918 (O_918,N_28434,N_29870);
or UO_919 (O_919,N_29582,N_29764);
nor UO_920 (O_920,N_27947,N_28635);
nor UO_921 (O_921,N_28957,N_28971);
nand UO_922 (O_922,N_28426,N_27128);
xnor UO_923 (O_923,N_28319,N_27003);
nor UO_924 (O_924,N_28618,N_28174);
or UO_925 (O_925,N_29490,N_27337);
and UO_926 (O_926,N_28877,N_27322);
nand UO_927 (O_927,N_29426,N_28642);
xnor UO_928 (O_928,N_28977,N_29326);
nand UO_929 (O_929,N_29021,N_29817);
or UO_930 (O_930,N_28664,N_29604);
or UO_931 (O_931,N_27110,N_28931);
and UO_932 (O_932,N_29717,N_27884);
and UO_933 (O_933,N_29558,N_28249);
and UO_934 (O_934,N_27596,N_27813);
nor UO_935 (O_935,N_27919,N_27171);
or UO_936 (O_936,N_28595,N_28372);
nand UO_937 (O_937,N_29246,N_28656);
xor UO_938 (O_938,N_27505,N_29479);
nand UO_939 (O_939,N_27022,N_28614);
xnor UO_940 (O_940,N_27888,N_27511);
and UO_941 (O_941,N_29649,N_27181);
or UO_942 (O_942,N_27399,N_27793);
nor UO_943 (O_943,N_29563,N_27230);
xor UO_944 (O_944,N_28910,N_29532);
or UO_945 (O_945,N_28755,N_29538);
nand UO_946 (O_946,N_29478,N_27535);
nand UO_947 (O_947,N_29537,N_29813);
and UO_948 (O_948,N_29355,N_28847);
nor UO_949 (O_949,N_28959,N_28660);
nand UO_950 (O_950,N_27501,N_27017);
xnor UO_951 (O_951,N_28285,N_28875);
nor UO_952 (O_952,N_29430,N_27551);
nand UO_953 (O_953,N_27104,N_28352);
nor UO_954 (O_954,N_27424,N_28924);
nor UO_955 (O_955,N_28381,N_27206);
xnor UO_956 (O_956,N_27948,N_28529);
or UO_957 (O_957,N_29344,N_28071);
and UO_958 (O_958,N_27479,N_29091);
and UO_959 (O_959,N_29064,N_29569);
nand UO_960 (O_960,N_27733,N_27898);
nor UO_961 (O_961,N_28502,N_27742);
and UO_962 (O_962,N_28703,N_28480);
nor UO_963 (O_963,N_29693,N_28568);
and UO_964 (O_964,N_27782,N_29665);
nand UO_965 (O_965,N_28688,N_28895);
nor UO_966 (O_966,N_29466,N_28238);
nand UO_967 (O_967,N_29711,N_29104);
and UO_968 (O_968,N_27973,N_28188);
and UO_969 (O_969,N_28411,N_29454);
and UO_970 (O_970,N_29118,N_29669);
or UO_971 (O_971,N_27463,N_27807);
nor UO_972 (O_972,N_27218,N_28061);
nand UO_973 (O_973,N_29708,N_28979);
or UO_974 (O_974,N_27691,N_28607);
nor UO_975 (O_975,N_27172,N_27111);
or UO_976 (O_976,N_28322,N_27204);
or UO_977 (O_977,N_29393,N_27231);
and UO_978 (O_978,N_29107,N_29233);
and UO_979 (O_979,N_27629,N_28908);
nand UO_980 (O_980,N_28733,N_29743);
xnor UO_981 (O_981,N_27282,N_29949);
nor UO_982 (O_982,N_28539,N_27705);
nand UO_983 (O_983,N_28357,N_29988);
or UO_984 (O_984,N_29117,N_28710);
xnor UO_985 (O_985,N_28155,N_27927);
nor UO_986 (O_986,N_29243,N_29678);
nand UO_987 (O_987,N_29791,N_29957);
nand UO_988 (O_988,N_28108,N_28867);
nor UO_989 (O_989,N_27186,N_27652);
nand UO_990 (O_990,N_29351,N_27202);
xor UO_991 (O_991,N_29769,N_27384);
and UO_992 (O_992,N_27975,N_27747);
nand UO_993 (O_993,N_28526,N_27061);
xor UO_994 (O_994,N_29437,N_29877);
nand UO_995 (O_995,N_28830,N_29312);
xor UO_996 (O_996,N_29609,N_29814);
and UO_997 (O_997,N_27292,N_29498);
nor UO_998 (O_998,N_27589,N_27931);
nor UO_999 (O_999,N_28085,N_29648);
and UO_1000 (O_1000,N_29628,N_29947);
nand UO_1001 (O_1001,N_29173,N_29071);
and UO_1002 (O_1002,N_27326,N_28175);
nand UO_1003 (O_1003,N_29281,N_28440);
nor UO_1004 (O_1004,N_29030,N_29535);
or UO_1005 (O_1005,N_29768,N_28293);
and UO_1006 (O_1006,N_28882,N_28774);
nand UO_1007 (O_1007,N_28300,N_29368);
and UO_1008 (O_1008,N_29171,N_28692);
nor UO_1009 (O_1009,N_29373,N_27298);
xor UO_1010 (O_1010,N_28419,N_28325);
nand UO_1011 (O_1011,N_28164,N_29821);
or UO_1012 (O_1012,N_28119,N_27410);
or UO_1013 (O_1013,N_28752,N_28263);
xnor UO_1014 (O_1014,N_27442,N_29606);
and UO_1015 (O_1015,N_27877,N_27752);
and UO_1016 (O_1016,N_29364,N_27549);
and UO_1017 (O_1017,N_29009,N_27611);
or UO_1018 (O_1018,N_29577,N_27072);
xor UO_1019 (O_1019,N_28872,N_27499);
and UO_1020 (O_1020,N_28404,N_29193);
or UO_1021 (O_1021,N_27192,N_28384);
nor UO_1022 (O_1022,N_27640,N_28510);
nand UO_1023 (O_1023,N_28585,N_27809);
xnor UO_1024 (O_1024,N_27506,N_28837);
xor UO_1025 (O_1025,N_28973,N_27751);
nor UO_1026 (O_1026,N_28127,N_27166);
xnor UO_1027 (O_1027,N_29585,N_27189);
or UO_1028 (O_1028,N_28099,N_27759);
xor UO_1029 (O_1029,N_28651,N_28020);
or UO_1030 (O_1030,N_29940,N_27706);
or UO_1031 (O_1031,N_28735,N_27531);
xnor UO_1032 (O_1032,N_27923,N_27358);
and UO_1033 (O_1033,N_27832,N_28177);
xnor UO_1034 (O_1034,N_29337,N_27039);
or UO_1035 (O_1035,N_27303,N_29361);
xor UO_1036 (O_1036,N_29832,N_27091);
xnor UO_1037 (O_1037,N_29506,N_29777);
nor UO_1038 (O_1038,N_29210,N_29986);
and UO_1039 (O_1039,N_27389,N_27554);
or UO_1040 (O_1040,N_28033,N_27665);
nor UO_1041 (O_1041,N_28965,N_28514);
and UO_1042 (O_1042,N_28925,N_27625);
nor UO_1043 (O_1043,N_27368,N_29652);
or UO_1044 (O_1044,N_28375,N_28814);
nand UO_1045 (O_1045,N_28478,N_28831);
xnor UO_1046 (O_1046,N_27833,N_28102);
or UO_1047 (O_1047,N_27775,N_27529);
nor UO_1048 (O_1048,N_28323,N_29771);
and UO_1049 (O_1049,N_29431,N_28881);
and UO_1050 (O_1050,N_29026,N_28062);
nor UO_1051 (O_1051,N_29037,N_28674);
and UO_1052 (O_1052,N_29770,N_28212);
xnor UO_1053 (O_1053,N_27934,N_29139);
nand UO_1054 (O_1054,N_27089,N_29948);
nand UO_1055 (O_1055,N_29927,N_27416);
xnor UO_1056 (O_1056,N_27066,N_28573);
and UO_1057 (O_1057,N_28078,N_28858);
nor UO_1058 (O_1058,N_28431,N_28074);
and UO_1059 (O_1059,N_29522,N_27334);
and UO_1060 (O_1060,N_28134,N_28096);
xor UO_1061 (O_1061,N_28870,N_27161);
or UO_1062 (O_1062,N_28722,N_27108);
nand UO_1063 (O_1063,N_29056,N_28777);
nor UO_1064 (O_1064,N_29655,N_29436);
xor UO_1065 (O_1065,N_27032,N_29540);
and UO_1066 (O_1066,N_27436,N_28897);
and UO_1067 (O_1067,N_27239,N_28022);
or UO_1068 (O_1068,N_28832,N_27251);
and UO_1069 (O_1069,N_29990,N_27866);
and UO_1070 (O_1070,N_27331,N_27806);
xnor UO_1071 (O_1071,N_28749,N_28368);
and UO_1072 (O_1072,N_27697,N_28408);
or UO_1073 (O_1073,N_29738,N_29113);
or UO_1074 (O_1074,N_29313,N_27311);
and UO_1075 (O_1075,N_27701,N_27457);
nor UO_1076 (O_1076,N_29151,N_29005);
nor UO_1077 (O_1077,N_27259,N_27382);
or UO_1078 (O_1078,N_29937,N_28943);
xnor UO_1079 (O_1079,N_29410,N_28576);
xnor UO_1080 (O_1080,N_28095,N_27167);
nor UO_1081 (O_1081,N_29493,N_28950);
xnor UO_1082 (O_1082,N_29400,N_28232);
xor UO_1083 (O_1083,N_27158,N_29192);
xor UO_1084 (O_1084,N_27970,N_28090);
or UO_1085 (O_1085,N_29471,N_29534);
xnor UO_1086 (O_1086,N_28588,N_29055);
nand UO_1087 (O_1087,N_29876,N_29333);
or UO_1088 (O_1088,N_29601,N_27413);
xnor UO_1089 (O_1089,N_27597,N_28318);
nor UO_1090 (O_1090,N_28476,N_28314);
nor UO_1091 (O_1091,N_27087,N_29187);
or UO_1092 (O_1092,N_27029,N_29519);
nand UO_1093 (O_1093,N_29745,N_28412);
nor UO_1094 (O_1094,N_28617,N_29586);
nand UO_1095 (O_1095,N_28829,N_27467);
and UO_1096 (O_1096,N_29406,N_27107);
nand UO_1097 (O_1097,N_29793,N_28944);
nand UO_1098 (O_1098,N_27146,N_28501);
nor UO_1099 (O_1099,N_27962,N_29746);
nor UO_1100 (O_1100,N_29785,N_27578);
and UO_1101 (O_1101,N_27552,N_27542);
and UO_1102 (O_1102,N_27210,N_29607);
nor UO_1103 (O_1103,N_29975,N_29991);
xor UO_1104 (O_1104,N_27594,N_29749);
and UO_1105 (O_1105,N_28291,N_29444);
and UO_1106 (O_1106,N_28714,N_27534);
nand UO_1107 (O_1107,N_29469,N_29899);
xor UO_1108 (O_1108,N_29952,N_29891);
nor UO_1109 (O_1109,N_27969,N_27889);
xnor UO_1110 (O_1110,N_29996,N_28439);
or UO_1111 (O_1111,N_29689,N_28901);
or UO_1112 (O_1112,N_28590,N_28544);
or UO_1113 (O_1113,N_29812,N_28146);
and UO_1114 (O_1114,N_28024,N_27666);
xor UO_1115 (O_1115,N_29660,N_29275);
xnor UO_1116 (O_1116,N_28856,N_27861);
nor UO_1117 (O_1117,N_27745,N_28036);
nand UO_1118 (O_1118,N_29345,N_29780);
or UO_1119 (O_1119,N_29847,N_28782);
nand UO_1120 (O_1120,N_27675,N_28140);
nand UO_1121 (O_1121,N_28554,N_27613);
or UO_1122 (O_1122,N_29327,N_28374);
and UO_1123 (O_1123,N_29694,N_28458);
or UO_1124 (O_1124,N_28391,N_28914);
nand UO_1125 (O_1125,N_27533,N_27984);
and UO_1126 (O_1126,N_28643,N_28998);
nor UO_1127 (O_1127,N_29755,N_28545);
and UO_1128 (O_1128,N_28306,N_28713);
and UO_1129 (O_1129,N_27398,N_28396);
and UO_1130 (O_1130,N_29369,N_28540);
or UO_1131 (O_1131,N_27316,N_29523);
nand UO_1132 (O_1132,N_28465,N_29322);
and UO_1133 (O_1133,N_27476,N_29020);
nand UO_1134 (O_1134,N_29278,N_29571);
xor UO_1135 (O_1135,N_28775,N_28894);
xor UO_1136 (O_1136,N_27007,N_28648);
nor UO_1137 (O_1137,N_28741,N_28712);
and UO_1138 (O_1138,N_28126,N_27115);
nand UO_1139 (O_1139,N_28619,N_27369);
nand UO_1140 (O_1140,N_28304,N_29610);
xor UO_1141 (O_1141,N_28341,N_29879);
xnor UO_1142 (O_1142,N_28623,N_29356);
or UO_1143 (O_1143,N_29999,N_29357);
or UO_1144 (O_1144,N_27513,N_28366);
nand UO_1145 (O_1145,N_29644,N_29392);
nor UO_1146 (O_1146,N_28606,N_27603);
or UO_1147 (O_1147,N_29674,N_27960);
nand UO_1148 (O_1148,N_28247,N_27190);
xnor UO_1149 (O_1149,N_28547,N_29051);
and UO_1150 (O_1150,N_28092,N_28854);
nand UO_1151 (O_1151,N_27147,N_29593);
xnor UO_1152 (O_1152,N_29525,N_28762);
or UO_1153 (O_1153,N_27799,N_29638);
or UO_1154 (O_1154,N_28631,N_28353);
or UO_1155 (O_1155,N_29447,N_29796);
nor UO_1156 (O_1156,N_27105,N_28494);
or UO_1157 (O_1157,N_28050,N_28474);
nor UO_1158 (O_1158,N_27492,N_29237);
xor UO_1159 (O_1159,N_27867,N_29167);
xnor UO_1160 (O_1160,N_29560,N_29943);
xnor UO_1161 (O_1161,N_28260,N_29642);
or UO_1162 (O_1162,N_27891,N_29968);
nor UO_1163 (O_1163,N_28855,N_27920);
xor UO_1164 (O_1164,N_29288,N_28154);
nand UO_1165 (O_1165,N_29965,N_29475);
or UO_1166 (O_1166,N_28039,N_29334);
and UO_1167 (O_1167,N_27078,N_29065);
nand UO_1168 (O_1168,N_28496,N_27439);
and UO_1169 (O_1169,N_27143,N_28861);
nor UO_1170 (O_1170,N_27267,N_29698);
or UO_1171 (O_1171,N_29204,N_27750);
nand UO_1172 (O_1172,N_27826,N_28826);
nand UO_1173 (O_1173,N_28638,N_29216);
and UO_1174 (O_1174,N_29274,N_29808);
and UO_1175 (O_1175,N_28616,N_27856);
xnor UO_1176 (O_1176,N_28757,N_29121);
or UO_1177 (O_1177,N_27913,N_27351);
xnor UO_1178 (O_1178,N_27031,N_28405);
and UO_1179 (O_1179,N_29050,N_27545);
nand UO_1180 (O_1180,N_28582,N_29551);
nor UO_1181 (O_1181,N_29982,N_28764);
and UO_1182 (O_1182,N_28229,N_27943);
and UO_1183 (O_1183,N_29852,N_28230);
nand UO_1184 (O_1184,N_27869,N_28392);
xor UO_1185 (O_1185,N_29240,N_28816);
nand UO_1186 (O_1186,N_27786,N_28435);
and UO_1187 (O_1187,N_29234,N_28086);
or UO_1188 (O_1188,N_29423,N_27070);
xnor UO_1189 (O_1189,N_29078,N_27174);
or UO_1190 (O_1190,N_28701,N_27028);
xnor UO_1191 (O_1191,N_27153,N_28170);
nor UO_1192 (O_1192,N_29094,N_27272);
nor UO_1193 (O_1193,N_29299,N_28181);
or UO_1194 (O_1194,N_27214,N_29562);
nor UO_1195 (O_1195,N_27417,N_28994);
and UO_1196 (O_1196,N_28817,N_28416);
or UO_1197 (O_1197,N_27804,N_28508);
xnor UO_1198 (O_1198,N_28262,N_27843);
nand UO_1199 (O_1199,N_29790,N_29194);
or UO_1200 (O_1200,N_29625,N_28515);
xnor UO_1201 (O_1201,N_28048,N_28282);
xnor UO_1202 (O_1202,N_28524,N_28365);
nand UO_1203 (O_1203,N_29959,N_28009);
nand UO_1204 (O_1204,N_29896,N_29587);
and UO_1205 (O_1205,N_29533,N_27418);
nand UO_1206 (O_1206,N_29083,N_27145);
nand UO_1207 (O_1207,N_27253,N_27738);
or UO_1208 (O_1208,N_29467,N_29396);
nor UO_1209 (O_1209,N_29989,N_27926);
nor UO_1210 (O_1210,N_28321,N_27054);
xnor UO_1211 (O_1211,N_27286,N_27646);
nor UO_1212 (O_1212,N_27816,N_28601);
and UO_1213 (O_1213,N_29402,N_29623);
and UO_1214 (O_1214,N_27577,N_29914);
nor UO_1215 (O_1215,N_27929,N_29744);
nor UO_1216 (O_1216,N_28639,N_27980);
nand UO_1217 (O_1217,N_28542,N_29513);
xor UO_1218 (O_1218,N_27631,N_28101);
and UO_1219 (O_1219,N_27055,N_29404);
or UO_1220 (O_1220,N_29445,N_28489);
xor UO_1221 (O_1221,N_28936,N_28149);
or UO_1222 (O_1222,N_27957,N_29568);
and UO_1223 (O_1223,N_29389,N_28163);
and UO_1224 (O_1224,N_29886,N_29692);
and UO_1225 (O_1225,N_29867,N_28902);
nand UO_1226 (O_1226,N_27260,N_27780);
or UO_1227 (O_1227,N_28369,N_27790);
xnor UO_1228 (O_1228,N_29862,N_28316);
nand UO_1229 (O_1229,N_29058,N_28997);
nand UO_1230 (O_1230,N_27740,N_29156);
or UO_1231 (O_1231,N_29284,N_28624);
nor UO_1232 (O_1232,N_27604,N_28438);
or UO_1233 (O_1233,N_29760,N_27451);
or UO_1234 (O_1234,N_29303,N_27380);
nor UO_1235 (O_1235,N_29463,N_29668);
nand UO_1236 (O_1236,N_28983,N_27034);
and UO_1237 (O_1237,N_27581,N_27502);
xnor UO_1238 (O_1238,N_28464,N_28225);
or UO_1239 (O_1239,N_27818,N_29175);
nand UO_1240 (O_1240,N_28724,N_29489);
nand UO_1241 (O_1241,N_27217,N_29148);
and UO_1242 (O_1242,N_27324,N_29110);
nor UO_1243 (O_1243,N_29166,N_27000);
and UO_1244 (O_1244,N_29340,N_27381);
xnor UO_1245 (O_1245,N_29014,N_28103);
and UO_1246 (O_1246,N_28654,N_28850);
nand UO_1247 (O_1247,N_28602,N_28786);
nand UO_1248 (O_1248,N_27517,N_28449);
and UO_1249 (O_1249,N_29480,N_27321);
and UO_1250 (O_1250,N_28055,N_27120);
and UO_1251 (O_1251,N_27950,N_27651);
or UO_1252 (O_1252,N_27497,N_28261);
or UO_1253 (O_1253,N_28051,N_27674);
nand UO_1254 (O_1254,N_28342,N_27938);
nand UO_1255 (O_1255,N_29578,N_28640);
xor UO_1256 (O_1256,N_29736,N_28023);
nand UO_1257 (O_1257,N_28887,N_28491);
or UO_1258 (O_1258,N_29476,N_28340);
xnor UO_1259 (O_1259,N_28975,N_28430);
nor UO_1260 (O_1260,N_28834,N_29268);
or UO_1261 (O_1261,N_29235,N_29767);
or UO_1262 (O_1262,N_27065,N_29484);
or UO_1263 (O_1263,N_28558,N_27537);
and UO_1264 (O_1264,N_28243,N_28596);
nor UO_1265 (O_1265,N_28500,N_29492);
or UO_1266 (O_1266,N_27796,N_29528);
nand UO_1267 (O_1267,N_28128,N_29049);
xnor UO_1268 (O_1268,N_27559,N_27308);
nor UO_1269 (O_1269,N_29720,N_29343);
nor UO_1270 (O_1270,N_29298,N_28373);
nand UO_1271 (O_1271,N_27430,N_27532);
xnor UO_1272 (O_1272,N_29895,N_27668);
xnor UO_1273 (O_1273,N_28364,N_29908);
nand UO_1274 (O_1274,N_27336,N_28613);
or UO_1275 (O_1275,N_27099,N_29850);
xor UO_1276 (O_1276,N_29072,N_29363);
xor UO_1277 (O_1277,N_28409,N_27440);
or UO_1278 (O_1278,N_29137,N_27850);
nor UO_1279 (O_1279,N_28707,N_28575);
nand UO_1280 (O_1280,N_29381,N_29289);
or UO_1281 (O_1281,N_27872,N_27327);
or UO_1282 (O_1282,N_27193,N_29963);
nor UO_1283 (O_1283,N_28433,N_27393);
nor UO_1284 (O_1284,N_29086,N_29297);
nand UO_1285 (O_1285,N_28484,N_29250);
nor UO_1286 (O_1286,N_29671,N_29779);
xnor UO_1287 (O_1287,N_28313,N_27663);
or UO_1288 (O_1288,N_28918,N_29843);
nor UO_1289 (O_1289,N_27857,N_27342);
nor UO_1290 (O_1290,N_27367,N_29501);
and UO_1291 (O_1291,N_29617,N_29291);
xnor UO_1292 (O_1292,N_28669,N_29643);
nor UO_1293 (O_1293,N_29076,N_28191);
or UO_1294 (O_1294,N_28428,N_27255);
nand UO_1295 (O_1295,N_29903,N_28343);
nand UO_1296 (O_1296,N_27881,N_28267);
and UO_1297 (O_1297,N_27672,N_28846);
nor UO_1298 (O_1298,N_29321,N_27290);
nor UO_1299 (O_1299,N_29145,N_29325);
xor UO_1300 (O_1300,N_28076,N_29917);
or UO_1301 (O_1301,N_29892,N_28219);
xnor UO_1302 (O_1302,N_28562,N_28308);
xnor UO_1303 (O_1303,N_28949,N_27609);
or UO_1304 (O_1304,N_28759,N_28552);
nor UO_1305 (O_1305,N_28893,N_28976);
xor UO_1306 (O_1306,N_28888,N_27667);
nand UO_1307 (O_1307,N_27868,N_27828);
nand UO_1308 (O_1308,N_27593,N_27170);
and UO_1309 (O_1309,N_29272,N_29639);
or UO_1310 (O_1310,N_29421,N_28214);
and UO_1311 (O_1311,N_29206,N_27991);
nand UO_1312 (O_1312,N_28561,N_27784);
and UO_1313 (O_1313,N_29280,N_28288);
or UO_1314 (O_1314,N_28615,N_28424);
and UO_1315 (O_1315,N_29646,N_28732);
nand UO_1316 (O_1316,N_27800,N_28705);
xnor UO_1317 (O_1317,N_28079,N_27225);
or UO_1318 (O_1318,N_29868,N_29906);
nand UO_1319 (O_1319,N_27901,N_28069);
and UO_1320 (O_1320,N_29658,N_29920);
nor UO_1321 (O_1321,N_29979,N_27359);
or UO_1322 (O_1322,N_29690,N_27235);
and UO_1323 (O_1323,N_29681,N_28371);
nand UO_1324 (O_1324,N_27916,N_27540);
nand UO_1325 (O_1325,N_29715,N_27271);
nand UO_1326 (O_1326,N_29405,N_29457);
nor UO_1327 (O_1327,N_29901,N_27620);
nor UO_1328 (O_1328,N_28580,N_27184);
nand UO_1329 (O_1329,N_27987,N_29242);
nor UO_1330 (O_1330,N_29500,N_27557);
nand UO_1331 (O_1331,N_27403,N_29594);
and UO_1332 (O_1332,N_29075,N_28172);
nor UO_1333 (O_1333,N_29552,N_29068);
or UO_1334 (O_1334,N_27783,N_29128);
nor UO_1335 (O_1335,N_28303,N_29695);
nand UO_1336 (O_1336,N_29294,N_29090);
xnor UO_1337 (O_1337,N_28385,N_27743);
or UO_1338 (O_1338,N_28609,N_28115);
or UO_1339 (O_1339,N_29795,N_28644);
nand UO_1340 (O_1340,N_29320,N_28336);
nand UO_1341 (O_1341,N_27228,N_29330);
nor UO_1342 (O_1342,N_27930,N_29412);
nor UO_1343 (O_1343,N_27098,N_28490);
nand UO_1344 (O_1344,N_28840,N_29657);
nor UO_1345 (O_1345,N_28168,N_27468);
and UO_1346 (O_1346,N_29348,N_28019);
xor UO_1347 (O_1347,N_27448,N_27689);
or UO_1348 (O_1348,N_27958,N_29100);
nand UO_1349 (O_1349,N_28196,N_27903);
nor UO_1350 (O_1350,N_28789,N_28567);
nor UO_1351 (O_1351,N_27909,N_29172);
and UO_1352 (O_1352,N_28630,N_27097);
nand UO_1353 (O_1353,N_28743,N_29096);
or UO_1354 (O_1354,N_28245,N_28227);
nor UO_1355 (O_1355,N_27794,N_27131);
xnor UO_1356 (O_1356,N_27754,N_28564);
xor UO_1357 (O_1357,N_27387,N_27026);
nand UO_1358 (O_1358,N_27817,N_27617);
nand UO_1359 (O_1359,N_29849,N_28482);
or UO_1360 (O_1360,N_27083,N_28550);
nand UO_1361 (O_1361,N_27449,N_27068);
nor UO_1362 (O_1362,N_27755,N_28593);
nor UO_1363 (O_1363,N_28028,N_27194);
or UO_1364 (O_1364,N_27905,N_28763);
xor UO_1365 (O_1365,N_28479,N_29826);
or UO_1366 (O_1366,N_28383,N_28347);
xor UO_1367 (O_1367,N_29939,N_29150);
nand UO_1368 (O_1368,N_29106,N_27910);
and UO_1369 (O_1369,N_28106,N_27441);
or UO_1370 (O_1370,N_28441,N_29904);
or UO_1371 (O_1371,N_29509,N_29539);
or UO_1372 (O_1372,N_29053,N_27465);
and UO_1373 (O_1373,N_29006,N_28849);
nand UO_1374 (O_1374,N_29497,N_27347);
nand UO_1375 (O_1375,N_28223,N_27471);
nand UO_1376 (O_1376,N_27539,N_29894);
xnor UO_1377 (O_1377,N_29752,N_29942);
and UO_1378 (O_1378,N_27354,N_27312);
and UO_1379 (O_1379,N_29874,N_27873);
xor UO_1380 (O_1380,N_29099,N_28907);
or UO_1381 (O_1381,N_27764,N_27018);
and UO_1382 (O_1382,N_28241,N_28647);
and UO_1383 (O_1383,N_29520,N_28727);
nor UO_1384 (O_1384,N_27883,N_27391);
or UO_1385 (O_1385,N_29740,N_29545);
or UO_1386 (O_1386,N_27470,N_29941);
xnor UO_1387 (O_1387,N_27876,N_29775);
nand UO_1388 (O_1388,N_28171,N_28937);
nor UO_1389 (O_1389,N_29928,N_27245);
xor UO_1390 (O_1390,N_28953,N_28919);
or UO_1391 (O_1391,N_29477,N_29672);
and UO_1392 (O_1392,N_29269,N_28049);
xnor UO_1393 (O_1393,N_28532,N_29314);
xor UO_1394 (O_1394,N_28563,N_28005);
nor UO_1395 (O_1395,N_27972,N_29220);
nor UO_1396 (O_1396,N_29488,N_29319);
nand UO_1397 (O_1397,N_29921,N_29122);
or UO_1398 (O_1398,N_28517,N_27036);
xnor UO_1399 (O_1399,N_29618,N_27789);
and UO_1400 (O_1400,N_28746,N_29414);
nor UO_1401 (O_1401,N_29842,N_28900);
nor UO_1402 (O_1402,N_28437,N_29397);
and UO_1403 (O_1403,N_29028,N_29057);
or UO_1404 (O_1404,N_29352,N_28153);
or UO_1405 (O_1405,N_28662,N_29102);
xnor UO_1406 (O_1406,N_29925,N_27377);
and UO_1407 (O_1407,N_29460,N_28268);
nand UO_1408 (O_1408,N_27412,N_28704);
or UO_1409 (O_1409,N_29066,N_27908);
or UO_1410 (O_1410,N_27855,N_28053);
or UO_1411 (O_1411,N_28330,N_29754);
xor UO_1412 (O_1412,N_27836,N_28610);
and UO_1413 (O_1413,N_29855,N_29987);
or UO_1414 (O_1414,N_27363,N_29247);
xnor UO_1415 (O_1415,N_28414,N_29772);
or UO_1416 (O_1416,N_28761,N_29024);
xnor UO_1417 (O_1417,N_27122,N_27293);
and UO_1418 (O_1418,N_28299,N_28217);
xnor UO_1419 (O_1419,N_27493,N_27838);
nand UO_1420 (O_1420,N_29733,N_27114);
and UO_1421 (O_1421,N_27489,N_29661);
or UO_1422 (O_1422,N_27756,N_29716);
xor UO_1423 (O_1423,N_27990,N_29632);
or UO_1424 (O_1424,N_28105,N_28646);
or UO_1425 (O_1425,N_27699,N_29781);
xnor UO_1426 (O_1426,N_27612,N_28693);
or UO_1427 (O_1427,N_28462,N_27287);
xor UO_1428 (O_1428,N_28543,N_28913);
nand UO_1429 (O_1429,N_29579,N_29809);
nor UO_1430 (O_1430,N_29670,N_27355);
and UO_1431 (O_1431,N_29328,N_28198);
nand UO_1432 (O_1432,N_28485,N_27760);
nor UO_1433 (O_1433,N_29977,N_27736);
and UO_1434 (O_1434,N_27198,N_29264);
nand UO_1435 (O_1435,N_28969,N_28822);
nor UO_1436 (O_1436,N_29878,N_27422);
nor UO_1437 (O_1437,N_29399,N_29311);
nor UO_1438 (O_1438,N_29529,N_28748);
or UO_1439 (O_1439,N_27042,N_28697);
and UO_1440 (O_1440,N_27273,N_28790);
and UO_1441 (O_1441,N_28772,N_29041);
or UO_1442 (O_1442,N_28390,N_29819);
nor UO_1443 (O_1443,N_27659,N_27495);
or UO_1444 (O_1444,N_27848,N_27385);
nand UO_1445 (O_1445,N_29262,N_28239);
nand UO_1446 (O_1446,N_29153,N_28060);
nand UO_1447 (O_1447,N_27769,N_29160);
nor UO_1448 (O_1448,N_29550,N_29022);
or UO_1449 (O_1449,N_28359,N_28320);
or UO_1450 (O_1450,N_28380,N_27019);
nor UO_1451 (O_1451,N_28995,N_29663);
nand UO_1452 (O_1452,N_28386,N_29922);
or UO_1453 (O_1453,N_29258,N_28281);
and UO_1454 (O_1454,N_27878,N_28292);
or UO_1455 (O_1455,N_28869,N_27274);
or UO_1456 (O_1456,N_29416,N_29146);
and UO_1457 (O_1457,N_28461,N_28344);
nor UO_1458 (O_1458,N_29487,N_28828);
nor UO_1459 (O_1459,N_29329,N_27650);
nor UO_1460 (O_1460,N_27703,N_29222);
nand UO_1461 (O_1461,N_27074,N_28037);
nor UO_1462 (O_1462,N_29168,N_28147);
and UO_1463 (O_1463,N_29844,N_28780);
xnor UO_1464 (O_1464,N_28087,N_29931);
nand UO_1465 (O_1465,N_29293,N_29889);
or UO_1466 (O_1466,N_29000,N_27719);
nand UO_1467 (O_1467,N_28920,N_29758);
or UO_1468 (O_1468,N_28065,N_28058);
nand UO_1469 (O_1469,N_29682,N_28862);
nor UO_1470 (O_1470,N_29685,N_28021);
or UO_1471 (O_1471,N_27694,N_27940);
xnor UO_1472 (O_1472,N_27918,N_29391);
or UO_1473 (O_1473,N_28506,N_29788);
or UO_1474 (O_1474,N_27353,N_28766);
nand UO_1475 (O_1475,N_28835,N_28122);
or UO_1476 (O_1476,N_28525,N_28698);
and UO_1477 (O_1477,N_27092,N_28151);
nand UO_1478 (O_1478,N_29207,N_28182);
and UO_1479 (O_1479,N_28387,N_29714);
nand UO_1480 (O_1480,N_29158,N_27349);
and UO_1481 (O_1481,N_27654,N_28220);
nor UO_1482 (O_1482,N_28620,N_27798);
and UO_1483 (O_1483,N_27588,N_27538);
nand UO_1484 (O_1484,N_29599,N_27746);
nand UO_1485 (O_1485,N_28978,N_27482);
or UO_1486 (O_1486,N_27080,N_29726);
and UO_1487 (O_1487,N_28574,N_28505);
or UO_1488 (O_1488,N_27295,N_27615);
xnor UO_1489 (O_1489,N_29036,N_28089);
nand UO_1490 (O_1490,N_27229,N_28985);
nand UO_1491 (O_1491,N_28469,N_28143);
and UO_1492 (O_1492,N_29907,N_28329);
xor UO_1493 (O_1493,N_28929,N_29702);
xnor UO_1494 (O_1494,N_28107,N_27787);
xnor UO_1495 (O_1495,N_27458,N_27343);
nand UO_1496 (O_1496,N_27015,N_28425);
or UO_1497 (O_1497,N_29789,N_27373);
nor UO_1498 (O_1498,N_29473,N_28072);
or UO_1499 (O_1499,N_27478,N_27090);
and UO_1500 (O_1500,N_28099,N_28072);
or UO_1501 (O_1501,N_28699,N_28479);
and UO_1502 (O_1502,N_27429,N_27000);
nand UO_1503 (O_1503,N_28083,N_29360);
xnor UO_1504 (O_1504,N_29521,N_27535);
and UO_1505 (O_1505,N_27710,N_29590);
nand UO_1506 (O_1506,N_29097,N_29727);
nand UO_1507 (O_1507,N_27388,N_28011);
xor UO_1508 (O_1508,N_28255,N_27898);
nor UO_1509 (O_1509,N_28342,N_27105);
or UO_1510 (O_1510,N_29294,N_28931);
and UO_1511 (O_1511,N_28254,N_27625);
nand UO_1512 (O_1512,N_29601,N_28357);
nand UO_1513 (O_1513,N_27906,N_29820);
nand UO_1514 (O_1514,N_28237,N_27055);
nand UO_1515 (O_1515,N_27468,N_28300);
and UO_1516 (O_1516,N_29172,N_27099);
xnor UO_1517 (O_1517,N_27617,N_27111);
nand UO_1518 (O_1518,N_29719,N_28270);
xor UO_1519 (O_1519,N_29423,N_28418);
xnor UO_1520 (O_1520,N_28485,N_29380);
xnor UO_1521 (O_1521,N_27130,N_27091);
or UO_1522 (O_1522,N_28360,N_28605);
nand UO_1523 (O_1523,N_28727,N_29103);
and UO_1524 (O_1524,N_28763,N_28649);
xnor UO_1525 (O_1525,N_28673,N_29734);
and UO_1526 (O_1526,N_28448,N_28007);
or UO_1527 (O_1527,N_28449,N_27857);
nand UO_1528 (O_1528,N_29392,N_27455);
xor UO_1529 (O_1529,N_29387,N_29782);
xnor UO_1530 (O_1530,N_27387,N_28343);
xnor UO_1531 (O_1531,N_27926,N_28589);
nand UO_1532 (O_1532,N_28713,N_28829);
or UO_1533 (O_1533,N_29215,N_29157);
nand UO_1534 (O_1534,N_29884,N_28187);
or UO_1535 (O_1535,N_29595,N_27070);
or UO_1536 (O_1536,N_29597,N_27579);
and UO_1537 (O_1537,N_29196,N_29002);
or UO_1538 (O_1538,N_28973,N_29498);
nor UO_1539 (O_1539,N_27516,N_28361);
or UO_1540 (O_1540,N_29356,N_28338);
xor UO_1541 (O_1541,N_29447,N_28021);
or UO_1542 (O_1542,N_28238,N_28229);
nor UO_1543 (O_1543,N_27204,N_27234);
xnor UO_1544 (O_1544,N_29268,N_28583);
nand UO_1545 (O_1545,N_27458,N_28591);
and UO_1546 (O_1546,N_27708,N_27232);
xor UO_1547 (O_1547,N_28708,N_28920);
and UO_1548 (O_1548,N_28295,N_29886);
or UO_1549 (O_1549,N_27310,N_27626);
xor UO_1550 (O_1550,N_29588,N_28371);
xnor UO_1551 (O_1551,N_28766,N_29242);
or UO_1552 (O_1552,N_27975,N_27649);
xor UO_1553 (O_1553,N_27784,N_29632);
xnor UO_1554 (O_1554,N_29581,N_27566);
nor UO_1555 (O_1555,N_28319,N_28323);
or UO_1556 (O_1556,N_27836,N_28776);
or UO_1557 (O_1557,N_27547,N_28733);
xor UO_1558 (O_1558,N_27116,N_28970);
nor UO_1559 (O_1559,N_29695,N_28985);
nor UO_1560 (O_1560,N_28008,N_29156);
xor UO_1561 (O_1561,N_28052,N_27176);
nand UO_1562 (O_1562,N_28118,N_28382);
xnor UO_1563 (O_1563,N_29767,N_28100);
xnor UO_1564 (O_1564,N_28179,N_28137);
nor UO_1565 (O_1565,N_29915,N_28498);
and UO_1566 (O_1566,N_29367,N_29990);
nor UO_1567 (O_1567,N_28570,N_27908);
and UO_1568 (O_1568,N_27228,N_29852);
xor UO_1569 (O_1569,N_28919,N_29994);
xnor UO_1570 (O_1570,N_29329,N_27440);
nor UO_1571 (O_1571,N_28515,N_29237);
or UO_1572 (O_1572,N_29070,N_27071);
or UO_1573 (O_1573,N_27496,N_29487);
or UO_1574 (O_1574,N_28655,N_27740);
xor UO_1575 (O_1575,N_28210,N_28506);
nor UO_1576 (O_1576,N_28331,N_29215);
xnor UO_1577 (O_1577,N_29844,N_27858);
xnor UO_1578 (O_1578,N_28078,N_29737);
xor UO_1579 (O_1579,N_28531,N_27853);
and UO_1580 (O_1580,N_27328,N_28613);
xor UO_1581 (O_1581,N_28249,N_27736);
and UO_1582 (O_1582,N_29404,N_28159);
nor UO_1583 (O_1583,N_29809,N_29816);
or UO_1584 (O_1584,N_29277,N_27508);
and UO_1585 (O_1585,N_29133,N_27599);
xor UO_1586 (O_1586,N_29013,N_27325);
or UO_1587 (O_1587,N_27469,N_27520);
xnor UO_1588 (O_1588,N_28524,N_28783);
or UO_1589 (O_1589,N_27601,N_29458);
nor UO_1590 (O_1590,N_29202,N_28796);
or UO_1591 (O_1591,N_27294,N_27378);
xnor UO_1592 (O_1592,N_27767,N_27428);
or UO_1593 (O_1593,N_29839,N_29092);
xnor UO_1594 (O_1594,N_28995,N_29736);
or UO_1595 (O_1595,N_29880,N_28618);
or UO_1596 (O_1596,N_29441,N_29985);
and UO_1597 (O_1597,N_27544,N_28236);
xor UO_1598 (O_1598,N_28737,N_28416);
nand UO_1599 (O_1599,N_27012,N_27465);
and UO_1600 (O_1600,N_27473,N_27717);
nor UO_1601 (O_1601,N_28380,N_27384);
and UO_1602 (O_1602,N_28632,N_28280);
xor UO_1603 (O_1603,N_28008,N_28803);
or UO_1604 (O_1604,N_29183,N_29423);
xnor UO_1605 (O_1605,N_29424,N_28939);
or UO_1606 (O_1606,N_27850,N_29686);
or UO_1607 (O_1607,N_27831,N_29156);
xnor UO_1608 (O_1608,N_27689,N_28682);
nor UO_1609 (O_1609,N_27194,N_29618);
nand UO_1610 (O_1610,N_28308,N_27595);
and UO_1611 (O_1611,N_29179,N_29613);
nor UO_1612 (O_1612,N_28805,N_29754);
nor UO_1613 (O_1613,N_29269,N_27654);
nor UO_1614 (O_1614,N_29849,N_29268);
nand UO_1615 (O_1615,N_27710,N_28907);
nand UO_1616 (O_1616,N_27826,N_27341);
xor UO_1617 (O_1617,N_28857,N_27334);
and UO_1618 (O_1618,N_27003,N_29869);
nor UO_1619 (O_1619,N_28690,N_27897);
nand UO_1620 (O_1620,N_27614,N_28079);
nand UO_1621 (O_1621,N_29360,N_28938);
nand UO_1622 (O_1622,N_27805,N_28576);
xnor UO_1623 (O_1623,N_29211,N_28060);
xnor UO_1624 (O_1624,N_28583,N_28255);
nand UO_1625 (O_1625,N_29214,N_27212);
nand UO_1626 (O_1626,N_29181,N_29641);
nor UO_1627 (O_1627,N_28415,N_28991);
or UO_1628 (O_1628,N_27712,N_27154);
nor UO_1629 (O_1629,N_27839,N_28995);
nand UO_1630 (O_1630,N_28529,N_29436);
nor UO_1631 (O_1631,N_28649,N_28616);
nand UO_1632 (O_1632,N_28919,N_28273);
nor UO_1633 (O_1633,N_29741,N_27447);
nor UO_1634 (O_1634,N_28512,N_28600);
or UO_1635 (O_1635,N_27533,N_28107);
nor UO_1636 (O_1636,N_29851,N_28622);
xor UO_1637 (O_1637,N_29433,N_29121);
nand UO_1638 (O_1638,N_27351,N_27181);
nor UO_1639 (O_1639,N_29569,N_27372);
nor UO_1640 (O_1640,N_27192,N_28277);
nor UO_1641 (O_1641,N_29347,N_28867);
xor UO_1642 (O_1642,N_27609,N_27745);
or UO_1643 (O_1643,N_28890,N_27115);
or UO_1644 (O_1644,N_28361,N_27297);
nand UO_1645 (O_1645,N_27582,N_27406);
or UO_1646 (O_1646,N_29476,N_28866);
or UO_1647 (O_1647,N_27622,N_27205);
nor UO_1648 (O_1648,N_27998,N_29002);
nor UO_1649 (O_1649,N_28427,N_29947);
and UO_1650 (O_1650,N_28885,N_27806);
nor UO_1651 (O_1651,N_27861,N_27179);
xnor UO_1652 (O_1652,N_29968,N_28232);
or UO_1653 (O_1653,N_29552,N_29417);
and UO_1654 (O_1654,N_27483,N_28415);
xnor UO_1655 (O_1655,N_29612,N_29470);
or UO_1656 (O_1656,N_28122,N_27868);
xor UO_1657 (O_1657,N_29228,N_29481);
xnor UO_1658 (O_1658,N_27051,N_28389);
or UO_1659 (O_1659,N_28692,N_27170);
and UO_1660 (O_1660,N_28796,N_28616);
or UO_1661 (O_1661,N_28689,N_28451);
nand UO_1662 (O_1662,N_28296,N_29151);
nand UO_1663 (O_1663,N_28289,N_27457);
or UO_1664 (O_1664,N_29551,N_28986);
and UO_1665 (O_1665,N_29614,N_28183);
or UO_1666 (O_1666,N_27813,N_28655);
nor UO_1667 (O_1667,N_27936,N_28855);
nand UO_1668 (O_1668,N_27998,N_29907);
xor UO_1669 (O_1669,N_29913,N_27723);
nor UO_1670 (O_1670,N_28829,N_27096);
or UO_1671 (O_1671,N_29796,N_28928);
xnor UO_1672 (O_1672,N_29264,N_28404);
and UO_1673 (O_1673,N_27617,N_29577);
nand UO_1674 (O_1674,N_29820,N_28687);
nor UO_1675 (O_1675,N_27472,N_28521);
nor UO_1676 (O_1676,N_29394,N_28883);
and UO_1677 (O_1677,N_29371,N_28481);
or UO_1678 (O_1678,N_29261,N_27992);
xor UO_1679 (O_1679,N_27218,N_28564);
or UO_1680 (O_1680,N_29979,N_27040);
xor UO_1681 (O_1681,N_29800,N_27381);
xor UO_1682 (O_1682,N_27566,N_29230);
and UO_1683 (O_1683,N_28444,N_28431);
and UO_1684 (O_1684,N_28122,N_29031);
nor UO_1685 (O_1685,N_29748,N_28961);
or UO_1686 (O_1686,N_28075,N_29518);
nand UO_1687 (O_1687,N_28085,N_28451);
and UO_1688 (O_1688,N_27021,N_29484);
and UO_1689 (O_1689,N_29037,N_27677);
or UO_1690 (O_1690,N_27843,N_27470);
nor UO_1691 (O_1691,N_29144,N_28053);
nor UO_1692 (O_1692,N_29091,N_29662);
and UO_1693 (O_1693,N_28015,N_28363);
or UO_1694 (O_1694,N_28117,N_29151);
nor UO_1695 (O_1695,N_28064,N_28553);
nor UO_1696 (O_1696,N_27504,N_29086);
nand UO_1697 (O_1697,N_27528,N_29213);
and UO_1698 (O_1698,N_29274,N_28623);
and UO_1699 (O_1699,N_28516,N_28435);
nand UO_1700 (O_1700,N_27453,N_28626);
or UO_1701 (O_1701,N_29030,N_29488);
xnor UO_1702 (O_1702,N_28852,N_27563);
nor UO_1703 (O_1703,N_29193,N_27084);
nor UO_1704 (O_1704,N_28900,N_27196);
nor UO_1705 (O_1705,N_27709,N_28779);
xnor UO_1706 (O_1706,N_29976,N_27912);
or UO_1707 (O_1707,N_27753,N_29860);
and UO_1708 (O_1708,N_27087,N_29069);
nor UO_1709 (O_1709,N_28078,N_29579);
nand UO_1710 (O_1710,N_29991,N_28732);
nand UO_1711 (O_1711,N_28213,N_29673);
nand UO_1712 (O_1712,N_29334,N_27845);
or UO_1713 (O_1713,N_27800,N_28336);
xor UO_1714 (O_1714,N_28273,N_28461);
nand UO_1715 (O_1715,N_29609,N_27601);
nand UO_1716 (O_1716,N_27778,N_27789);
or UO_1717 (O_1717,N_29017,N_27303);
and UO_1718 (O_1718,N_28337,N_29666);
xor UO_1719 (O_1719,N_29627,N_28370);
xor UO_1720 (O_1720,N_27348,N_27448);
nor UO_1721 (O_1721,N_28251,N_29072);
or UO_1722 (O_1722,N_28798,N_27977);
nand UO_1723 (O_1723,N_27187,N_27043);
xor UO_1724 (O_1724,N_28523,N_27716);
nor UO_1725 (O_1725,N_28471,N_29344);
xor UO_1726 (O_1726,N_27023,N_29914);
or UO_1727 (O_1727,N_27446,N_29593);
or UO_1728 (O_1728,N_28680,N_29350);
nand UO_1729 (O_1729,N_28227,N_29154);
and UO_1730 (O_1730,N_29598,N_27828);
nand UO_1731 (O_1731,N_29762,N_27275);
or UO_1732 (O_1732,N_27144,N_28321);
xnor UO_1733 (O_1733,N_27845,N_27690);
xnor UO_1734 (O_1734,N_29861,N_28326);
nand UO_1735 (O_1735,N_29942,N_28789);
nand UO_1736 (O_1736,N_28909,N_28071);
or UO_1737 (O_1737,N_27252,N_27541);
nand UO_1738 (O_1738,N_28531,N_27751);
or UO_1739 (O_1739,N_29065,N_29633);
nor UO_1740 (O_1740,N_28618,N_29474);
xnor UO_1741 (O_1741,N_27843,N_27769);
nor UO_1742 (O_1742,N_28903,N_27139);
and UO_1743 (O_1743,N_27296,N_29799);
nor UO_1744 (O_1744,N_29757,N_27451);
or UO_1745 (O_1745,N_29537,N_29449);
and UO_1746 (O_1746,N_29220,N_28901);
and UO_1747 (O_1747,N_28720,N_27207);
xnor UO_1748 (O_1748,N_27866,N_29708);
nor UO_1749 (O_1749,N_29952,N_28346);
nand UO_1750 (O_1750,N_29596,N_29898);
nor UO_1751 (O_1751,N_28716,N_27004);
or UO_1752 (O_1752,N_27603,N_27833);
xor UO_1753 (O_1753,N_29343,N_27001);
and UO_1754 (O_1754,N_27192,N_28527);
and UO_1755 (O_1755,N_29026,N_29393);
nand UO_1756 (O_1756,N_28067,N_27369);
xor UO_1757 (O_1757,N_29473,N_27538);
or UO_1758 (O_1758,N_27569,N_29159);
and UO_1759 (O_1759,N_27941,N_29400);
xor UO_1760 (O_1760,N_29074,N_29877);
and UO_1761 (O_1761,N_28462,N_29336);
nand UO_1762 (O_1762,N_29454,N_28198);
and UO_1763 (O_1763,N_27214,N_27444);
and UO_1764 (O_1764,N_29152,N_29976);
or UO_1765 (O_1765,N_27868,N_28407);
or UO_1766 (O_1766,N_29595,N_28078);
and UO_1767 (O_1767,N_28009,N_29129);
xor UO_1768 (O_1768,N_28053,N_27247);
or UO_1769 (O_1769,N_28604,N_29423);
and UO_1770 (O_1770,N_29531,N_28671);
nand UO_1771 (O_1771,N_28869,N_28694);
or UO_1772 (O_1772,N_27871,N_28601);
nor UO_1773 (O_1773,N_29849,N_27764);
or UO_1774 (O_1774,N_28419,N_29897);
nor UO_1775 (O_1775,N_29502,N_27427);
or UO_1776 (O_1776,N_29337,N_28183);
and UO_1777 (O_1777,N_29798,N_27341);
nor UO_1778 (O_1778,N_29998,N_29835);
nand UO_1779 (O_1779,N_29862,N_28758);
and UO_1780 (O_1780,N_27470,N_29811);
nand UO_1781 (O_1781,N_28857,N_29352);
xnor UO_1782 (O_1782,N_27649,N_28189);
or UO_1783 (O_1783,N_29214,N_28761);
nor UO_1784 (O_1784,N_29908,N_29716);
nand UO_1785 (O_1785,N_27626,N_29459);
nand UO_1786 (O_1786,N_27483,N_29514);
and UO_1787 (O_1787,N_28922,N_27093);
or UO_1788 (O_1788,N_28993,N_29696);
and UO_1789 (O_1789,N_28689,N_28782);
or UO_1790 (O_1790,N_27751,N_27816);
or UO_1791 (O_1791,N_27593,N_27630);
or UO_1792 (O_1792,N_29578,N_27520);
xnor UO_1793 (O_1793,N_27679,N_29691);
nor UO_1794 (O_1794,N_29809,N_29594);
and UO_1795 (O_1795,N_28805,N_28816);
nor UO_1796 (O_1796,N_28231,N_28189);
or UO_1797 (O_1797,N_29418,N_27049);
nand UO_1798 (O_1798,N_28981,N_28422);
nand UO_1799 (O_1799,N_29133,N_27659);
or UO_1800 (O_1800,N_27694,N_28993);
xnor UO_1801 (O_1801,N_29820,N_29747);
and UO_1802 (O_1802,N_27938,N_28768);
nor UO_1803 (O_1803,N_27172,N_29929);
and UO_1804 (O_1804,N_27081,N_28074);
or UO_1805 (O_1805,N_28903,N_28772);
nand UO_1806 (O_1806,N_28735,N_28613);
nand UO_1807 (O_1807,N_28191,N_28093);
nor UO_1808 (O_1808,N_28814,N_29640);
nand UO_1809 (O_1809,N_29309,N_29839);
or UO_1810 (O_1810,N_29077,N_28981);
or UO_1811 (O_1811,N_28714,N_27741);
nand UO_1812 (O_1812,N_28075,N_28540);
xor UO_1813 (O_1813,N_27271,N_27839);
nand UO_1814 (O_1814,N_27108,N_28844);
nor UO_1815 (O_1815,N_29131,N_29859);
or UO_1816 (O_1816,N_28478,N_29455);
and UO_1817 (O_1817,N_27774,N_27201);
xor UO_1818 (O_1818,N_28402,N_29961);
nor UO_1819 (O_1819,N_29162,N_29666);
nand UO_1820 (O_1820,N_27026,N_29533);
or UO_1821 (O_1821,N_29690,N_28756);
or UO_1822 (O_1822,N_27442,N_28216);
and UO_1823 (O_1823,N_29120,N_29261);
nand UO_1824 (O_1824,N_29180,N_28446);
nor UO_1825 (O_1825,N_29965,N_27163);
xnor UO_1826 (O_1826,N_29621,N_28501);
nand UO_1827 (O_1827,N_27678,N_28949);
nor UO_1828 (O_1828,N_29249,N_28880);
xor UO_1829 (O_1829,N_28083,N_27599);
and UO_1830 (O_1830,N_28614,N_29545);
nand UO_1831 (O_1831,N_27844,N_28117);
nor UO_1832 (O_1832,N_28929,N_27070);
xnor UO_1833 (O_1833,N_28357,N_28637);
or UO_1834 (O_1834,N_29512,N_28475);
and UO_1835 (O_1835,N_28207,N_29221);
and UO_1836 (O_1836,N_27146,N_27794);
xor UO_1837 (O_1837,N_28357,N_28743);
and UO_1838 (O_1838,N_27125,N_27050);
nor UO_1839 (O_1839,N_28430,N_29818);
and UO_1840 (O_1840,N_29004,N_28801);
nand UO_1841 (O_1841,N_29571,N_29750);
nand UO_1842 (O_1842,N_29843,N_29079);
xnor UO_1843 (O_1843,N_29603,N_27129);
and UO_1844 (O_1844,N_27166,N_29936);
nand UO_1845 (O_1845,N_29701,N_27438);
nor UO_1846 (O_1846,N_28831,N_27453);
xor UO_1847 (O_1847,N_29995,N_27117);
nand UO_1848 (O_1848,N_27172,N_29166);
nor UO_1849 (O_1849,N_29148,N_29534);
xor UO_1850 (O_1850,N_29764,N_28846);
xor UO_1851 (O_1851,N_29357,N_28619);
and UO_1852 (O_1852,N_28995,N_29592);
and UO_1853 (O_1853,N_27737,N_29081);
xor UO_1854 (O_1854,N_27593,N_28515);
or UO_1855 (O_1855,N_29970,N_28302);
or UO_1856 (O_1856,N_28202,N_27978);
or UO_1857 (O_1857,N_28573,N_29938);
nand UO_1858 (O_1858,N_27063,N_27914);
and UO_1859 (O_1859,N_27403,N_28655);
or UO_1860 (O_1860,N_29763,N_27648);
nand UO_1861 (O_1861,N_28275,N_27551);
nor UO_1862 (O_1862,N_28671,N_29168);
xor UO_1863 (O_1863,N_27441,N_28655);
xnor UO_1864 (O_1864,N_29823,N_27549);
xor UO_1865 (O_1865,N_28726,N_27338);
nand UO_1866 (O_1866,N_29877,N_27503);
nand UO_1867 (O_1867,N_28171,N_29204);
and UO_1868 (O_1868,N_29231,N_27266);
nor UO_1869 (O_1869,N_27519,N_27204);
xnor UO_1870 (O_1870,N_29721,N_28147);
nand UO_1871 (O_1871,N_27398,N_28096);
xnor UO_1872 (O_1872,N_28553,N_27950);
and UO_1873 (O_1873,N_29960,N_27008);
xnor UO_1874 (O_1874,N_27815,N_28022);
nor UO_1875 (O_1875,N_27225,N_28153);
xor UO_1876 (O_1876,N_28278,N_28060);
or UO_1877 (O_1877,N_27694,N_28220);
and UO_1878 (O_1878,N_28832,N_28509);
xnor UO_1879 (O_1879,N_27509,N_29157);
nand UO_1880 (O_1880,N_27006,N_27044);
and UO_1881 (O_1881,N_27622,N_28703);
nand UO_1882 (O_1882,N_28190,N_28992);
nand UO_1883 (O_1883,N_29545,N_27123);
xor UO_1884 (O_1884,N_29441,N_27749);
and UO_1885 (O_1885,N_27072,N_28880);
or UO_1886 (O_1886,N_29235,N_27259);
and UO_1887 (O_1887,N_29001,N_27927);
or UO_1888 (O_1888,N_29640,N_29970);
and UO_1889 (O_1889,N_29189,N_29119);
xor UO_1890 (O_1890,N_28713,N_29787);
nor UO_1891 (O_1891,N_28848,N_28087);
and UO_1892 (O_1892,N_28215,N_29240);
and UO_1893 (O_1893,N_29352,N_29219);
or UO_1894 (O_1894,N_29026,N_27135);
nand UO_1895 (O_1895,N_29401,N_28886);
nor UO_1896 (O_1896,N_28042,N_27146);
and UO_1897 (O_1897,N_27162,N_28985);
nor UO_1898 (O_1898,N_28923,N_29357);
nor UO_1899 (O_1899,N_28338,N_29906);
or UO_1900 (O_1900,N_27762,N_29918);
nor UO_1901 (O_1901,N_28391,N_29522);
nor UO_1902 (O_1902,N_28987,N_27896);
or UO_1903 (O_1903,N_27446,N_27145);
or UO_1904 (O_1904,N_29656,N_29897);
or UO_1905 (O_1905,N_27240,N_29045);
or UO_1906 (O_1906,N_27394,N_27638);
nor UO_1907 (O_1907,N_28962,N_29140);
and UO_1908 (O_1908,N_27405,N_27442);
nand UO_1909 (O_1909,N_28617,N_29314);
xnor UO_1910 (O_1910,N_27267,N_29607);
nor UO_1911 (O_1911,N_28117,N_28101);
and UO_1912 (O_1912,N_28244,N_28512);
nor UO_1913 (O_1913,N_29724,N_27675);
and UO_1914 (O_1914,N_29823,N_29581);
xor UO_1915 (O_1915,N_27464,N_27835);
and UO_1916 (O_1916,N_28148,N_29080);
xor UO_1917 (O_1917,N_29111,N_29552);
or UO_1918 (O_1918,N_27522,N_27768);
nand UO_1919 (O_1919,N_28361,N_27536);
nand UO_1920 (O_1920,N_28935,N_27451);
xnor UO_1921 (O_1921,N_28523,N_27607);
xor UO_1922 (O_1922,N_29426,N_29775);
xnor UO_1923 (O_1923,N_28677,N_27719);
xor UO_1924 (O_1924,N_27055,N_28192);
or UO_1925 (O_1925,N_27105,N_28703);
xor UO_1926 (O_1926,N_27591,N_28391);
or UO_1927 (O_1927,N_27168,N_28186);
nand UO_1928 (O_1928,N_27570,N_27326);
nand UO_1929 (O_1929,N_29849,N_28866);
nor UO_1930 (O_1930,N_28449,N_29784);
nor UO_1931 (O_1931,N_29259,N_29985);
nor UO_1932 (O_1932,N_28727,N_27890);
xnor UO_1933 (O_1933,N_27079,N_27006);
xnor UO_1934 (O_1934,N_27649,N_27272);
nand UO_1935 (O_1935,N_29502,N_28666);
nor UO_1936 (O_1936,N_28227,N_27972);
nand UO_1937 (O_1937,N_29832,N_27785);
xnor UO_1938 (O_1938,N_27974,N_28513);
nor UO_1939 (O_1939,N_27738,N_28055);
and UO_1940 (O_1940,N_27699,N_28004);
xor UO_1941 (O_1941,N_27178,N_27902);
nand UO_1942 (O_1942,N_27910,N_27873);
xnor UO_1943 (O_1943,N_28763,N_29112);
and UO_1944 (O_1944,N_27533,N_27931);
xnor UO_1945 (O_1945,N_29963,N_29356);
or UO_1946 (O_1946,N_29638,N_27980);
nand UO_1947 (O_1947,N_27743,N_28829);
and UO_1948 (O_1948,N_28309,N_29551);
or UO_1949 (O_1949,N_28030,N_27658);
nand UO_1950 (O_1950,N_27031,N_27975);
or UO_1951 (O_1951,N_28696,N_29082);
xnor UO_1952 (O_1952,N_29899,N_27919);
or UO_1953 (O_1953,N_28380,N_28826);
nor UO_1954 (O_1954,N_28000,N_28123);
or UO_1955 (O_1955,N_28695,N_27315);
or UO_1956 (O_1956,N_29698,N_27469);
and UO_1957 (O_1957,N_28660,N_28452);
nand UO_1958 (O_1958,N_27465,N_29584);
nor UO_1959 (O_1959,N_29374,N_28835);
or UO_1960 (O_1960,N_27726,N_29404);
nor UO_1961 (O_1961,N_29105,N_28792);
nor UO_1962 (O_1962,N_27038,N_28880);
nor UO_1963 (O_1963,N_29641,N_29943);
or UO_1964 (O_1964,N_29271,N_27974);
or UO_1965 (O_1965,N_27185,N_29229);
xor UO_1966 (O_1966,N_29230,N_27691);
or UO_1967 (O_1967,N_29316,N_29458);
xnor UO_1968 (O_1968,N_28432,N_28906);
nor UO_1969 (O_1969,N_28764,N_29637);
nand UO_1970 (O_1970,N_29606,N_27962);
xnor UO_1971 (O_1971,N_28195,N_27467);
and UO_1972 (O_1972,N_29122,N_27439);
and UO_1973 (O_1973,N_29817,N_28486);
and UO_1974 (O_1974,N_27850,N_28329);
or UO_1975 (O_1975,N_28315,N_27464);
and UO_1976 (O_1976,N_28396,N_29479);
or UO_1977 (O_1977,N_28469,N_28189);
xnor UO_1978 (O_1978,N_29647,N_29088);
xor UO_1979 (O_1979,N_29929,N_28090);
nand UO_1980 (O_1980,N_27682,N_28695);
xnor UO_1981 (O_1981,N_28204,N_29294);
xnor UO_1982 (O_1982,N_28395,N_29503);
and UO_1983 (O_1983,N_29219,N_27778);
and UO_1984 (O_1984,N_27237,N_29579);
nand UO_1985 (O_1985,N_28946,N_28869);
xor UO_1986 (O_1986,N_29626,N_29172);
or UO_1987 (O_1987,N_29061,N_28101);
nor UO_1988 (O_1988,N_29798,N_27907);
and UO_1989 (O_1989,N_29889,N_28031);
xor UO_1990 (O_1990,N_27153,N_28627);
nand UO_1991 (O_1991,N_27348,N_28388);
or UO_1992 (O_1992,N_28627,N_27386);
nor UO_1993 (O_1993,N_28345,N_29335);
and UO_1994 (O_1994,N_29568,N_27656);
xnor UO_1995 (O_1995,N_27155,N_28509);
xor UO_1996 (O_1996,N_27775,N_27219);
nor UO_1997 (O_1997,N_29187,N_28931);
xor UO_1998 (O_1998,N_29119,N_28199);
xnor UO_1999 (O_1999,N_27050,N_29407);
xor UO_2000 (O_2000,N_28046,N_27433);
nor UO_2001 (O_2001,N_29448,N_28065);
nor UO_2002 (O_2002,N_29412,N_27172);
nor UO_2003 (O_2003,N_28004,N_29890);
or UO_2004 (O_2004,N_28570,N_28962);
nor UO_2005 (O_2005,N_28258,N_29007);
nor UO_2006 (O_2006,N_28364,N_27465);
or UO_2007 (O_2007,N_28697,N_29589);
nor UO_2008 (O_2008,N_29443,N_27749);
nand UO_2009 (O_2009,N_29204,N_27686);
nor UO_2010 (O_2010,N_29387,N_28210);
nand UO_2011 (O_2011,N_27259,N_28162);
nand UO_2012 (O_2012,N_27025,N_29641);
xnor UO_2013 (O_2013,N_29514,N_27666);
nand UO_2014 (O_2014,N_27623,N_28036);
nor UO_2015 (O_2015,N_29104,N_28282);
or UO_2016 (O_2016,N_29256,N_27174);
and UO_2017 (O_2017,N_27988,N_27213);
or UO_2018 (O_2018,N_29735,N_29232);
nand UO_2019 (O_2019,N_28022,N_28613);
nand UO_2020 (O_2020,N_29494,N_27330);
and UO_2021 (O_2021,N_28061,N_27055);
and UO_2022 (O_2022,N_27071,N_29668);
nand UO_2023 (O_2023,N_29950,N_28841);
nand UO_2024 (O_2024,N_28428,N_27095);
or UO_2025 (O_2025,N_27992,N_29429);
xor UO_2026 (O_2026,N_29993,N_27744);
nand UO_2027 (O_2027,N_28028,N_28302);
nand UO_2028 (O_2028,N_27017,N_29701);
nand UO_2029 (O_2029,N_27033,N_27468);
nor UO_2030 (O_2030,N_29001,N_27992);
xnor UO_2031 (O_2031,N_29761,N_27844);
nand UO_2032 (O_2032,N_27485,N_27652);
nor UO_2033 (O_2033,N_27751,N_29208);
and UO_2034 (O_2034,N_29095,N_29328);
nor UO_2035 (O_2035,N_28455,N_28164);
or UO_2036 (O_2036,N_29495,N_29550);
xor UO_2037 (O_2037,N_29967,N_29003);
or UO_2038 (O_2038,N_28619,N_27668);
and UO_2039 (O_2039,N_29860,N_27026);
and UO_2040 (O_2040,N_29931,N_27952);
or UO_2041 (O_2041,N_27541,N_28574);
or UO_2042 (O_2042,N_28265,N_28635);
or UO_2043 (O_2043,N_27636,N_29511);
nand UO_2044 (O_2044,N_27008,N_27180);
xor UO_2045 (O_2045,N_27788,N_29748);
nor UO_2046 (O_2046,N_28196,N_28838);
nand UO_2047 (O_2047,N_27432,N_28903);
or UO_2048 (O_2048,N_29711,N_29645);
nand UO_2049 (O_2049,N_29178,N_28486);
nor UO_2050 (O_2050,N_27677,N_29870);
and UO_2051 (O_2051,N_29315,N_28605);
or UO_2052 (O_2052,N_29099,N_29352);
nand UO_2053 (O_2053,N_28556,N_28704);
or UO_2054 (O_2054,N_29835,N_27915);
or UO_2055 (O_2055,N_29711,N_28001);
xnor UO_2056 (O_2056,N_27325,N_29799);
xnor UO_2057 (O_2057,N_29802,N_27559);
and UO_2058 (O_2058,N_27813,N_29432);
nor UO_2059 (O_2059,N_27132,N_29689);
nor UO_2060 (O_2060,N_27799,N_29500);
or UO_2061 (O_2061,N_29235,N_27668);
nor UO_2062 (O_2062,N_28725,N_27812);
or UO_2063 (O_2063,N_27954,N_27107);
xor UO_2064 (O_2064,N_29286,N_28944);
and UO_2065 (O_2065,N_27894,N_29021);
and UO_2066 (O_2066,N_29852,N_28764);
xnor UO_2067 (O_2067,N_29050,N_27657);
or UO_2068 (O_2068,N_27702,N_27809);
nor UO_2069 (O_2069,N_27460,N_29712);
xnor UO_2070 (O_2070,N_27308,N_27063);
or UO_2071 (O_2071,N_27711,N_28718);
xor UO_2072 (O_2072,N_28597,N_28557);
and UO_2073 (O_2073,N_27201,N_29909);
and UO_2074 (O_2074,N_29362,N_29329);
nand UO_2075 (O_2075,N_28804,N_27496);
nand UO_2076 (O_2076,N_27032,N_28509);
or UO_2077 (O_2077,N_27814,N_27369);
or UO_2078 (O_2078,N_27867,N_28424);
or UO_2079 (O_2079,N_28435,N_27757);
or UO_2080 (O_2080,N_27298,N_28610);
nand UO_2081 (O_2081,N_28433,N_28984);
nor UO_2082 (O_2082,N_27226,N_28520);
nor UO_2083 (O_2083,N_28896,N_28129);
and UO_2084 (O_2084,N_28115,N_28771);
nor UO_2085 (O_2085,N_28228,N_29689);
and UO_2086 (O_2086,N_28234,N_27079);
or UO_2087 (O_2087,N_29015,N_27528);
nand UO_2088 (O_2088,N_28617,N_29063);
xnor UO_2089 (O_2089,N_28003,N_28500);
xnor UO_2090 (O_2090,N_27265,N_27553);
xnor UO_2091 (O_2091,N_28724,N_29874);
and UO_2092 (O_2092,N_29663,N_29523);
or UO_2093 (O_2093,N_29907,N_29830);
nor UO_2094 (O_2094,N_27672,N_27366);
or UO_2095 (O_2095,N_27090,N_28557);
nand UO_2096 (O_2096,N_27362,N_29287);
nand UO_2097 (O_2097,N_29931,N_29513);
nand UO_2098 (O_2098,N_28108,N_28608);
or UO_2099 (O_2099,N_27645,N_29429);
nor UO_2100 (O_2100,N_28483,N_28097);
xor UO_2101 (O_2101,N_28509,N_28784);
xor UO_2102 (O_2102,N_29959,N_27546);
nor UO_2103 (O_2103,N_28265,N_29091);
and UO_2104 (O_2104,N_27141,N_29214);
nor UO_2105 (O_2105,N_28574,N_28210);
nand UO_2106 (O_2106,N_27662,N_28362);
xnor UO_2107 (O_2107,N_29156,N_27432);
nand UO_2108 (O_2108,N_29067,N_29721);
or UO_2109 (O_2109,N_28147,N_27491);
nand UO_2110 (O_2110,N_29213,N_27958);
nand UO_2111 (O_2111,N_27158,N_29606);
xor UO_2112 (O_2112,N_29722,N_28100);
and UO_2113 (O_2113,N_28276,N_27568);
or UO_2114 (O_2114,N_28606,N_29706);
and UO_2115 (O_2115,N_28070,N_27942);
nand UO_2116 (O_2116,N_27813,N_29275);
xor UO_2117 (O_2117,N_29648,N_27849);
nor UO_2118 (O_2118,N_27257,N_27984);
nor UO_2119 (O_2119,N_28157,N_29872);
nor UO_2120 (O_2120,N_27940,N_29532);
nor UO_2121 (O_2121,N_28217,N_27348);
and UO_2122 (O_2122,N_28758,N_28646);
nor UO_2123 (O_2123,N_27954,N_28857);
nor UO_2124 (O_2124,N_29803,N_27312);
and UO_2125 (O_2125,N_27536,N_28936);
and UO_2126 (O_2126,N_28145,N_29823);
nand UO_2127 (O_2127,N_28136,N_29493);
nand UO_2128 (O_2128,N_29230,N_27795);
xnor UO_2129 (O_2129,N_27861,N_29697);
nor UO_2130 (O_2130,N_29209,N_27188);
and UO_2131 (O_2131,N_27231,N_29805);
nor UO_2132 (O_2132,N_27128,N_28509);
nand UO_2133 (O_2133,N_29160,N_28574);
and UO_2134 (O_2134,N_29972,N_28754);
xnor UO_2135 (O_2135,N_29976,N_29258);
nand UO_2136 (O_2136,N_27487,N_29663);
xor UO_2137 (O_2137,N_27492,N_29238);
or UO_2138 (O_2138,N_27811,N_28405);
nor UO_2139 (O_2139,N_27269,N_29031);
nand UO_2140 (O_2140,N_29206,N_28060);
or UO_2141 (O_2141,N_27288,N_28860);
and UO_2142 (O_2142,N_28425,N_27436);
xnor UO_2143 (O_2143,N_29616,N_28775);
or UO_2144 (O_2144,N_28091,N_28802);
or UO_2145 (O_2145,N_27646,N_28146);
nand UO_2146 (O_2146,N_29668,N_28638);
nor UO_2147 (O_2147,N_27863,N_27602);
xnor UO_2148 (O_2148,N_28191,N_28227);
nor UO_2149 (O_2149,N_27170,N_29806);
or UO_2150 (O_2150,N_28806,N_27021);
nand UO_2151 (O_2151,N_28433,N_29831);
nand UO_2152 (O_2152,N_27095,N_29972);
nand UO_2153 (O_2153,N_29851,N_29305);
nand UO_2154 (O_2154,N_28632,N_27422);
nand UO_2155 (O_2155,N_29357,N_28927);
or UO_2156 (O_2156,N_27460,N_29776);
nand UO_2157 (O_2157,N_28530,N_28165);
or UO_2158 (O_2158,N_27524,N_28041);
or UO_2159 (O_2159,N_28491,N_28095);
nor UO_2160 (O_2160,N_28991,N_29992);
or UO_2161 (O_2161,N_29584,N_29135);
or UO_2162 (O_2162,N_27491,N_27080);
nand UO_2163 (O_2163,N_29689,N_27534);
nor UO_2164 (O_2164,N_28080,N_27826);
nor UO_2165 (O_2165,N_29229,N_27128);
xnor UO_2166 (O_2166,N_29206,N_27687);
xnor UO_2167 (O_2167,N_28910,N_27884);
and UO_2168 (O_2168,N_29672,N_29693);
nand UO_2169 (O_2169,N_29950,N_27727);
or UO_2170 (O_2170,N_29848,N_27803);
xor UO_2171 (O_2171,N_28129,N_28142);
and UO_2172 (O_2172,N_28662,N_29735);
or UO_2173 (O_2173,N_28939,N_29997);
nor UO_2174 (O_2174,N_28620,N_27653);
nand UO_2175 (O_2175,N_29355,N_27624);
nand UO_2176 (O_2176,N_27352,N_28514);
nor UO_2177 (O_2177,N_27020,N_29481);
and UO_2178 (O_2178,N_29444,N_29782);
and UO_2179 (O_2179,N_27609,N_28202);
nand UO_2180 (O_2180,N_28114,N_27184);
and UO_2181 (O_2181,N_29455,N_29742);
and UO_2182 (O_2182,N_27998,N_29026);
and UO_2183 (O_2183,N_27850,N_28925);
and UO_2184 (O_2184,N_27758,N_29207);
nand UO_2185 (O_2185,N_29006,N_28636);
or UO_2186 (O_2186,N_29087,N_29676);
xor UO_2187 (O_2187,N_28783,N_29445);
nor UO_2188 (O_2188,N_29955,N_28443);
xnor UO_2189 (O_2189,N_27031,N_29644);
and UO_2190 (O_2190,N_27895,N_29613);
nand UO_2191 (O_2191,N_29709,N_28993);
and UO_2192 (O_2192,N_28352,N_28201);
nand UO_2193 (O_2193,N_29803,N_27076);
or UO_2194 (O_2194,N_27591,N_27734);
and UO_2195 (O_2195,N_28614,N_28878);
and UO_2196 (O_2196,N_28412,N_28850);
xnor UO_2197 (O_2197,N_28507,N_27910);
xnor UO_2198 (O_2198,N_29441,N_27280);
nor UO_2199 (O_2199,N_29679,N_27641);
nand UO_2200 (O_2200,N_27784,N_28291);
nor UO_2201 (O_2201,N_28555,N_28071);
nand UO_2202 (O_2202,N_28999,N_27081);
nand UO_2203 (O_2203,N_28994,N_29187);
nand UO_2204 (O_2204,N_27405,N_29108);
nand UO_2205 (O_2205,N_28004,N_29555);
xor UO_2206 (O_2206,N_27481,N_28361);
nand UO_2207 (O_2207,N_27860,N_29121);
or UO_2208 (O_2208,N_29638,N_29609);
or UO_2209 (O_2209,N_28330,N_29832);
and UO_2210 (O_2210,N_27990,N_27754);
nor UO_2211 (O_2211,N_28592,N_29434);
and UO_2212 (O_2212,N_28571,N_29704);
xor UO_2213 (O_2213,N_29391,N_29565);
xnor UO_2214 (O_2214,N_29788,N_28169);
nor UO_2215 (O_2215,N_29689,N_29811);
and UO_2216 (O_2216,N_28237,N_27733);
nand UO_2217 (O_2217,N_27880,N_27483);
or UO_2218 (O_2218,N_29341,N_27097);
or UO_2219 (O_2219,N_27827,N_29973);
or UO_2220 (O_2220,N_27923,N_27502);
and UO_2221 (O_2221,N_29979,N_29740);
nand UO_2222 (O_2222,N_28295,N_27337);
or UO_2223 (O_2223,N_29825,N_28245);
and UO_2224 (O_2224,N_29654,N_29367);
xnor UO_2225 (O_2225,N_29971,N_27325);
or UO_2226 (O_2226,N_29857,N_28141);
xor UO_2227 (O_2227,N_27971,N_27814);
xor UO_2228 (O_2228,N_27122,N_28403);
nor UO_2229 (O_2229,N_29410,N_27306);
nand UO_2230 (O_2230,N_28083,N_28219);
or UO_2231 (O_2231,N_27151,N_28453);
nand UO_2232 (O_2232,N_29247,N_27795);
nand UO_2233 (O_2233,N_29027,N_28404);
or UO_2234 (O_2234,N_29618,N_27268);
xnor UO_2235 (O_2235,N_27245,N_28246);
and UO_2236 (O_2236,N_28385,N_28912);
xnor UO_2237 (O_2237,N_29290,N_27039);
nor UO_2238 (O_2238,N_28529,N_27519);
xor UO_2239 (O_2239,N_28727,N_27734);
or UO_2240 (O_2240,N_28146,N_27976);
xor UO_2241 (O_2241,N_29027,N_29464);
nand UO_2242 (O_2242,N_27456,N_29018);
nand UO_2243 (O_2243,N_28521,N_27636);
nand UO_2244 (O_2244,N_27330,N_27495);
or UO_2245 (O_2245,N_27674,N_29235);
nor UO_2246 (O_2246,N_28968,N_27595);
nand UO_2247 (O_2247,N_27799,N_28015);
nor UO_2248 (O_2248,N_28226,N_28813);
nand UO_2249 (O_2249,N_29262,N_29587);
nor UO_2250 (O_2250,N_29930,N_29621);
or UO_2251 (O_2251,N_27244,N_28514);
or UO_2252 (O_2252,N_27040,N_28111);
nor UO_2253 (O_2253,N_28583,N_27773);
and UO_2254 (O_2254,N_28889,N_28819);
nor UO_2255 (O_2255,N_27561,N_28672);
and UO_2256 (O_2256,N_27472,N_29580);
xor UO_2257 (O_2257,N_29711,N_27426);
nand UO_2258 (O_2258,N_29805,N_29783);
nand UO_2259 (O_2259,N_27701,N_27250);
xnor UO_2260 (O_2260,N_29836,N_29735);
xor UO_2261 (O_2261,N_28471,N_28604);
nand UO_2262 (O_2262,N_27677,N_27102);
and UO_2263 (O_2263,N_29430,N_27589);
nand UO_2264 (O_2264,N_27694,N_28084);
xor UO_2265 (O_2265,N_28457,N_27273);
nand UO_2266 (O_2266,N_28584,N_27144);
nand UO_2267 (O_2267,N_27916,N_28547);
and UO_2268 (O_2268,N_28483,N_28508);
nor UO_2269 (O_2269,N_29612,N_27960);
nor UO_2270 (O_2270,N_27902,N_28522);
or UO_2271 (O_2271,N_27647,N_27261);
and UO_2272 (O_2272,N_27379,N_29359);
and UO_2273 (O_2273,N_27908,N_27239);
xnor UO_2274 (O_2274,N_27752,N_28695);
nor UO_2275 (O_2275,N_27237,N_29510);
nand UO_2276 (O_2276,N_27276,N_29166);
or UO_2277 (O_2277,N_28835,N_29990);
nand UO_2278 (O_2278,N_28584,N_28724);
nor UO_2279 (O_2279,N_28463,N_28960);
and UO_2280 (O_2280,N_28646,N_27000);
and UO_2281 (O_2281,N_29182,N_29693);
or UO_2282 (O_2282,N_27533,N_27927);
and UO_2283 (O_2283,N_29282,N_28723);
and UO_2284 (O_2284,N_29050,N_28388);
nor UO_2285 (O_2285,N_28143,N_27628);
xor UO_2286 (O_2286,N_28449,N_27275);
or UO_2287 (O_2287,N_27451,N_27637);
xor UO_2288 (O_2288,N_29856,N_27574);
and UO_2289 (O_2289,N_28062,N_28566);
nand UO_2290 (O_2290,N_29889,N_29010);
nand UO_2291 (O_2291,N_28656,N_28884);
xnor UO_2292 (O_2292,N_27041,N_29407);
nand UO_2293 (O_2293,N_28592,N_29245);
nand UO_2294 (O_2294,N_27151,N_28012);
or UO_2295 (O_2295,N_28040,N_29356);
nor UO_2296 (O_2296,N_27667,N_28458);
and UO_2297 (O_2297,N_27944,N_27750);
and UO_2298 (O_2298,N_28115,N_29389);
and UO_2299 (O_2299,N_29394,N_27284);
nand UO_2300 (O_2300,N_27508,N_27012);
or UO_2301 (O_2301,N_28356,N_28201);
nor UO_2302 (O_2302,N_29695,N_28382);
nor UO_2303 (O_2303,N_29171,N_28609);
or UO_2304 (O_2304,N_28605,N_27172);
xor UO_2305 (O_2305,N_27461,N_29880);
nand UO_2306 (O_2306,N_27389,N_27102);
nand UO_2307 (O_2307,N_27895,N_29305);
nor UO_2308 (O_2308,N_28300,N_28907);
or UO_2309 (O_2309,N_28324,N_27722);
or UO_2310 (O_2310,N_29336,N_27312);
xnor UO_2311 (O_2311,N_29990,N_27400);
xor UO_2312 (O_2312,N_28333,N_28997);
or UO_2313 (O_2313,N_27448,N_28851);
and UO_2314 (O_2314,N_29489,N_28266);
nor UO_2315 (O_2315,N_29958,N_29230);
xnor UO_2316 (O_2316,N_28731,N_28108);
and UO_2317 (O_2317,N_28913,N_27358);
xor UO_2318 (O_2318,N_28118,N_29373);
and UO_2319 (O_2319,N_27716,N_28149);
and UO_2320 (O_2320,N_28011,N_27902);
nor UO_2321 (O_2321,N_29011,N_28141);
and UO_2322 (O_2322,N_28114,N_28521);
or UO_2323 (O_2323,N_27905,N_29915);
xor UO_2324 (O_2324,N_27364,N_29782);
or UO_2325 (O_2325,N_28196,N_28011);
nor UO_2326 (O_2326,N_29758,N_28189);
nor UO_2327 (O_2327,N_27532,N_29525);
and UO_2328 (O_2328,N_29294,N_29110);
xor UO_2329 (O_2329,N_29124,N_28306);
xor UO_2330 (O_2330,N_29947,N_29467);
nand UO_2331 (O_2331,N_27500,N_29778);
or UO_2332 (O_2332,N_29130,N_27687);
nand UO_2333 (O_2333,N_29034,N_28691);
nand UO_2334 (O_2334,N_29025,N_28889);
or UO_2335 (O_2335,N_28755,N_27976);
or UO_2336 (O_2336,N_29312,N_29376);
nor UO_2337 (O_2337,N_27863,N_28639);
or UO_2338 (O_2338,N_28843,N_27144);
xor UO_2339 (O_2339,N_29539,N_27895);
nor UO_2340 (O_2340,N_29744,N_29044);
nor UO_2341 (O_2341,N_28891,N_27136);
and UO_2342 (O_2342,N_27852,N_28880);
or UO_2343 (O_2343,N_27075,N_29715);
xnor UO_2344 (O_2344,N_28320,N_29103);
or UO_2345 (O_2345,N_28784,N_29571);
nor UO_2346 (O_2346,N_29026,N_27811);
xor UO_2347 (O_2347,N_27528,N_29834);
or UO_2348 (O_2348,N_29115,N_27707);
xor UO_2349 (O_2349,N_28687,N_29683);
nor UO_2350 (O_2350,N_28035,N_28073);
nor UO_2351 (O_2351,N_28856,N_28920);
or UO_2352 (O_2352,N_27338,N_27100);
or UO_2353 (O_2353,N_29969,N_29766);
xor UO_2354 (O_2354,N_29680,N_27338);
or UO_2355 (O_2355,N_27869,N_27504);
nand UO_2356 (O_2356,N_28317,N_27768);
or UO_2357 (O_2357,N_29575,N_27712);
and UO_2358 (O_2358,N_28540,N_28112);
and UO_2359 (O_2359,N_27736,N_27387);
nand UO_2360 (O_2360,N_29998,N_27931);
nand UO_2361 (O_2361,N_29811,N_29326);
xnor UO_2362 (O_2362,N_28202,N_28191);
nor UO_2363 (O_2363,N_29905,N_27072);
and UO_2364 (O_2364,N_29557,N_27726);
or UO_2365 (O_2365,N_28468,N_27479);
or UO_2366 (O_2366,N_28470,N_29754);
and UO_2367 (O_2367,N_28626,N_28726);
xnor UO_2368 (O_2368,N_27292,N_28402);
nor UO_2369 (O_2369,N_28276,N_29737);
xor UO_2370 (O_2370,N_28024,N_28217);
and UO_2371 (O_2371,N_28349,N_27002);
nor UO_2372 (O_2372,N_27092,N_27307);
nor UO_2373 (O_2373,N_27148,N_29831);
xor UO_2374 (O_2374,N_28500,N_29035);
and UO_2375 (O_2375,N_28846,N_29171);
or UO_2376 (O_2376,N_29594,N_29734);
and UO_2377 (O_2377,N_28396,N_27608);
and UO_2378 (O_2378,N_28163,N_29975);
nand UO_2379 (O_2379,N_29260,N_27633);
and UO_2380 (O_2380,N_27690,N_27015);
or UO_2381 (O_2381,N_27250,N_29486);
nor UO_2382 (O_2382,N_28313,N_29773);
xnor UO_2383 (O_2383,N_27204,N_29622);
xor UO_2384 (O_2384,N_27216,N_28477);
nand UO_2385 (O_2385,N_29557,N_29519);
xnor UO_2386 (O_2386,N_29201,N_29393);
xor UO_2387 (O_2387,N_29212,N_29820);
nor UO_2388 (O_2388,N_29528,N_28070);
xnor UO_2389 (O_2389,N_29407,N_28257);
nor UO_2390 (O_2390,N_27968,N_29620);
and UO_2391 (O_2391,N_27621,N_27746);
nand UO_2392 (O_2392,N_29884,N_27570);
xnor UO_2393 (O_2393,N_28805,N_28333);
nor UO_2394 (O_2394,N_29059,N_27347);
or UO_2395 (O_2395,N_29123,N_28965);
and UO_2396 (O_2396,N_28453,N_29690);
and UO_2397 (O_2397,N_28347,N_27975);
nand UO_2398 (O_2398,N_27417,N_28879);
nor UO_2399 (O_2399,N_29027,N_27516);
and UO_2400 (O_2400,N_28515,N_29333);
and UO_2401 (O_2401,N_27756,N_28194);
and UO_2402 (O_2402,N_28857,N_28505);
nor UO_2403 (O_2403,N_29024,N_29227);
nand UO_2404 (O_2404,N_29590,N_28921);
or UO_2405 (O_2405,N_27957,N_28937);
and UO_2406 (O_2406,N_28494,N_27501);
nor UO_2407 (O_2407,N_29419,N_28986);
xnor UO_2408 (O_2408,N_29384,N_28710);
nand UO_2409 (O_2409,N_28359,N_28750);
and UO_2410 (O_2410,N_28101,N_28177);
xnor UO_2411 (O_2411,N_29628,N_29497);
or UO_2412 (O_2412,N_28253,N_28624);
and UO_2413 (O_2413,N_29647,N_27123);
nand UO_2414 (O_2414,N_29499,N_27149);
nor UO_2415 (O_2415,N_28516,N_29411);
nor UO_2416 (O_2416,N_28874,N_27830);
xnor UO_2417 (O_2417,N_27616,N_27928);
xor UO_2418 (O_2418,N_29975,N_29734);
or UO_2419 (O_2419,N_27805,N_29731);
nor UO_2420 (O_2420,N_29150,N_28782);
nand UO_2421 (O_2421,N_27778,N_27251);
or UO_2422 (O_2422,N_27237,N_29168);
or UO_2423 (O_2423,N_27464,N_28265);
xor UO_2424 (O_2424,N_29926,N_29912);
xnor UO_2425 (O_2425,N_28187,N_28711);
xor UO_2426 (O_2426,N_28470,N_28356);
or UO_2427 (O_2427,N_27437,N_29384);
nand UO_2428 (O_2428,N_28982,N_27689);
xor UO_2429 (O_2429,N_28618,N_29560);
or UO_2430 (O_2430,N_28524,N_27260);
xor UO_2431 (O_2431,N_29854,N_29671);
nor UO_2432 (O_2432,N_29910,N_28439);
nor UO_2433 (O_2433,N_27965,N_29832);
and UO_2434 (O_2434,N_27580,N_28418);
nand UO_2435 (O_2435,N_29927,N_27684);
and UO_2436 (O_2436,N_28624,N_27760);
xor UO_2437 (O_2437,N_27887,N_29660);
nor UO_2438 (O_2438,N_29828,N_27042);
or UO_2439 (O_2439,N_27007,N_28625);
nand UO_2440 (O_2440,N_28401,N_28340);
nor UO_2441 (O_2441,N_29717,N_27802);
and UO_2442 (O_2442,N_29348,N_29725);
nand UO_2443 (O_2443,N_29616,N_29304);
or UO_2444 (O_2444,N_28458,N_27845);
and UO_2445 (O_2445,N_29168,N_28136);
or UO_2446 (O_2446,N_29216,N_28782);
or UO_2447 (O_2447,N_27338,N_28246);
nor UO_2448 (O_2448,N_28684,N_28161);
nor UO_2449 (O_2449,N_29693,N_29098);
nand UO_2450 (O_2450,N_29580,N_27313);
xnor UO_2451 (O_2451,N_29207,N_29179);
or UO_2452 (O_2452,N_29704,N_27602);
nor UO_2453 (O_2453,N_29764,N_28694);
and UO_2454 (O_2454,N_29626,N_29347);
or UO_2455 (O_2455,N_28327,N_28431);
nor UO_2456 (O_2456,N_29232,N_28448);
nor UO_2457 (O_2457,N_29026,N_27132);
nand UO_2458 (O_2458,N_27360,N_28603);
and UO_2459 (O_2459,N_28266,N_29328);
nand UO_2460 (O_2460,N_29240,N_27902);
nor UO_2461 (O_2461,N_27573,N_27618);
and UO_2462 (O_2462,N_27177,N_29383);
or UO_2463 (O_2463,N_27934,N_27894);
nor UO_2464 (O_2464,N_27604,N_27124);
nand UO_2465 (O_2465,N_29292,N_27197);
xor UO_2466 (O_2466,N_27956,N_28322);
nand UO_2467 (O_2467,N_28235,N_27542);
or UO_2468 (O_2468,N_28787,N_27097);
and UO_2469 (O_2469,N_27916,N_27535);
xnor UO_2470 (O_2470,N_29007,N_28498);
or UO_2471 (O_2471,N_28574,N_29564);
xor UO_2472 (O_2472,N_29312,N_29650);
xnor UO_2473 (O_2473,N_27381,N_29996);
or UO_2474 (O_2474,N_28167,N_27595);
or UO_2475 (O_2475,N_29891,N_27861);
nor UO_2476 (O_2476,N_29953,N_28115);
or UO_2477 (O_2477,N_27976,N_29706);
or UO_2478 (O_2478,N_27082,N_29614);
and UO_2479 (O_2479,N_27372,N_28412);
and UO_2480 (O_2480,N_27933,N_27392);
xor UO_2481 (O_2481,N_27966,N_28331);
nor UO_2482 (O_2482,N_28727,N_27749);
nand UO_2483 (O_2483,N_29308,N_29726);
xnor UO_2484 (O_2484,N_29024,N_29364);
nor UO_2485 (O_2485,N_28007,N_28021);
or UO_2486 (O_2486,N_29066,N_27706);
nor UO_2487 (O_2487,N_28910,N_28681);
nor UO_2488 (O_2488,N_27911,N_29306);
xnor UO_2489 (O_2489,N_27695,N_28683);
nand UO_2490 (O_2490,N_29291,N_28939);
and UO_2491 (O_2491,N_27078,N_29021);
xnor UO_2492 (O_2492,N_29101,N_27189);
or UO_2493 (O_2493,N_27068,N_28999);
and UO_2494 (O_2494,N_29461,N_28303);
or UO_2495 (O_2495,N_29913,N_27492);
or UO_2496 (O_2496,N_27726,N_28638);
xnor UO_2497 (O_2497,N_28059,N_28323);
nand UO_2498 (O_2498,N_28355,N_29134);
nor UO_2499 (O_2499,N_28803,N_29416);
nand UO_2500 (O_2500,N_27144,N_29940);
and UO_2501 (O_2501,N_27257,N_28168);
or UO_2502 (O_2502,N_29226,N_27158);
xnor UO_2503 (O_2503,N_28317,N_29753);
xor UO_2504 (O_2504,N_29764,N_28914);
or UO_2505 (O_2505,N_28495,N_27183);
nand UO_2506 (O_2506,N_29450,N_28847);
nand UO_2507 (O_2507,N_27443,N_28700);
nand UO_2508 (O_2508,N_27704,N_29619);
or UO_2509 (O_2509,N_27561,N_27408);
and UO_2510 (O_2510,N_28328,N_28717);
and UO_2511 (O_2511,N_29952,N_29041);
nor UO_2512 (O_2512,N_29842,N_29853);
nor UO_2513 (O_2513,N_28746,N_28134);
and UO_2514 (O_2514,N_27942,N_27306);
and UO_2515 (O_2515,N_27213,N_28411);
or UO_2516 (O_2516,N_27946,N_27762);
nand UO_2517 (O_2517,N_29245,N_27915);
or UO_2518 (O_2518,N_29179,N_29780);
nand UO_2519 (O_2519,N_27879,N_27201);
or UO_2520 (O_2520,N_28866,N_29044);
and UO_2521 (O_2521,N_28868,N_28557);
xnor UO_2522 (O_2522,N_29974,N_27853);
nand UO_2523 (O_2523,N_28788,N_27730);
and UO_2524 (O_2524,N_28741,N_28048);
nor UO_2525 (O_2525,N_28489,N_29918);
xnor UO_2526 (O_2526,N_28827,N_29387);
nand UO_2527 (O_2527,N_27969,N_28905);
nor UO_2528 (O_2528,N_28996,N_28826);
or UO_2529 (O_2529,N_28913,N_29791);
xor UO_2530 (O_2530,N_29314,N_29901);
nand UO_2531 (O_2531,N_28549,N_27872);
xor UO_2532 (O_2532,N_28731,N_28199);
or UO_2533 (O_2533,N_29070,N_29161);
or UO_2534 (O_2534,N_29672,N_27742);
nor UO_2535 (O_2535,N_27493,N_27860);
xor UO_2536 (O_2536,N_27582,N_29047);
xnor UO_2537 (O_2537,N_28352,N_27483);
nor UO_2538 (O_2538,N_29965,N_29725);
and UO_2539 (O_2539,N_27937,N_29853);
nand UO_2540 (O_2540,N_27577,N_29648);
or UO_2541 (O_2541,N_27261,N_27000);
or UO_2542 (O_2542,N_28667,N_29505);
or UO_2543 (O_2543,N_28012,N_27259);
xor UO_2544 (O_2544,N_27555,N_29542);
xnor UO_2545 (O_2545,N_27894,N_27761);
nor UO_2546 (O_2546,N_27217,N_27422);
nand UO_2547 (O_2547,N_27219,N_27478);
nor UO_2548 (O_2548,N_28909,N_29945);
xnor UO_2549 (O_2549,N_29129,N_28975);
or UO_2550 (O_2550,N_28518,N_28900);
nor UO_2551 (O_2551,N_29012,N_28740);
and UO_2552 (O_2552,N_29908,N_28639);
or UO_2553 (O_2553,N_27671,N_27590);
or UO_2554 (O_2554,N_28541,N_28634);
xnor UO_2555 (O_2555,N_27559,N_29808);
nand UO_2556 (O_2556,N_27687,N_27880);
and UO_2557 (O_2557,N_29491,N_29433);
and UO_2558 (O_2558,N_28450,N_29376);
nand UO_2559 (O_2559,N_28245,N_29065);
or UO_2560 (O_2560,N_28389,N_28693);
or UO_2561 (O_2561,N_29528,N_27762);
xnor UO_2562 (O_2562,N_27343,N_28908);
nand UO_2563 (O_2563,N_29739,N_29900);
and UO_2564 (O_2564,N_27663,N_28068);
or UO_2565 (O_2565,N_28427,N_27504);
nand UO_2566 (O_2566,N_28051,N_27966);
nand UO_2567 (O_2567,N_29615,N_27000);
xor UO_2568 (O_2568,N_28606,N_28012);
nand UO_2569 (O_2569,N_27752,N_28634);
xnor UO_2570 (O_2570,N_28844,N_28847);
nand UO_2571 (O_2571,N_29524,N_29725);
xor UO_2572 (O_2572,N_27285,N_29192);
or UO_2573 (O_2573,N_27783,N_28432);
nor UO_2574 (O_2574,N_29579,N_27310);
nor UO_2575 (O_2575,N_29090,N_29188);
or UO_2576 (O_2576,N_28182,N_29805);
and UO_2577 (O_2577,N_28160,N_28420);
nand UO_2578 (O_2578,N_27571,N_27666);
and UO_2579 (O_2579,N_27429,N_28545);
or UO_2580 (O_2580,N_28009,N_27845);
and UO_2581 (O_2581,N_27421,N_27389);
xnor UO_2582 (O_2582,N_28664,N_27452);
or UO_2583 (O_2583,N_29124,N_28262);
nor UO_2584 (O_2584,N_29248,N_27774);
and UO_2585 (O_2585,N_28967,N_28583);
nand UO_2586 (O_2586,N_29722,N_27883);
and UO_2587 (O_2587,N_29519,N_27919);
nor UO_2588 (O_2588,N_28900,N_27950);
nor UO_2589 (O_2589,N_27598,N_28797);
xor UO_2590 (O_2590,N_29940,N_27784);
nor UO_2591 (O_2591,N_27009,N_29698);
nand UO_2592 (O_2592,N_27274,N_29922);
xor UO_2593 (O_2593,N_27458,N_29157);
nand UO_2594 (O_2594,N_27731,N_28659);
nor UO_2595 (O_2595,N_28651,N_28320);
xor UO_2596 (O_2596,N_27499,N_27897);
xor UO_2597 (O_2597,N_27209,N_28668);
nor UO_2598 (O_2598,N_29292,N_29174);
nand UO_2599 (O_2599,N_27708,N_29839);
nor UO_2600 (O_2600,N_29898,N_28466);
nor UO_2601 (O_2601,N_29652,N_28411);
nand UO_2602 (O_2602,N_28274,N_28952);
and UO_2603 (O_2603,N_29836,N_27053);
and UO_2604 (O_2604,N_28020,N_29197);
nand UO_2605 (O_2605,N_29131,N_28499);
xnor UO_2606 (O_2606,N_29673,N_27608);
and UO_2607 (O_2607,N_28651,N_28178);
xnor UO_2608 (O_2608,N_27970,N_29131);
or UO_2609 (O_2609,N_28176,N_29689);
or UO_2610 (O_2610,N_27914,N_28404);
or UO_2611 (O_2611,N_28586,N_28387);
nand UO_2612 (O_2612,N_27042,N_28381);
nor UO_2613 (O_2613,N_28616,N_29243);
xnor UO_2614 (O_2614,N_28021,N_28206);
nor UO_2615 (O_2615,N_27427,N_27596);
xor UO_2616 (O_2616,N_29355,N_28416);
xor UO_2617 (O_2617,N_29436,N_28131);
xor UO_2618 (O_2618,N_29534,N_28905);
nand UO_2619 (O_2619,N_27886,N_29018);
or UO_2620 (O_2620,N_27274,N_27590);
nor UO_2621 (O_2621,N_27929,N_27293);
nand UO_2622 (O_2622,N_29977,N_27365);
nor UO_2623 (O_2623,N_27308,N_28427);
and UO_2624 (O_2624,N_28533,N_29917);
or UO_2625 (O_2625,N_28468,N_27781);
xnor UO_2626 (O_2626,N_29608,N_29640);
and UO_2627 (O_2627,N_29111,N_28546);
nand UO_2628 (O_2628,N_29780,N_27237);
or UO_2629 (O_2629,N_29975,N_28311);
or UO_2630 (O_2630,N_27387,N_27019);
and UO_2631 (O_2631,N_27657,N_27108);
nand UO_2632 (O_2632,N_27777,N_29194);
nand UO_2633 (O_2633,N_27012,N_29905);
nor UO_2634 (O_2634,N_28872,N_28590);
nand UO_2635 (O_2635,N_27057,N_27811);
or UO_2636 (O_2636,N_29767,N_28304);
xor UO_2637 (O_2637,N_27198,N_27361);
or UO_2638 (O_2638,N_28346,N_27565);
and UO_2639 (O_2639,N_29132,N_28885);
nand UO_2640 (O_2640,N_29472,N_28867);
or UO_2641 (O_2641,N_28587,N_28214);
nor UO_2642 (O_2642,N_28265,N_29444);
or UO_2643 (O_2643,N_28954,N_28599);
or UO_2644 (O_2644,N_28495,N_28769);
nor UO_2645 (O_2645,N_28380,N_28321);
and UO_2646 (O_2646,N_29593,N_28992);
nor UO_2647 (O_2647,N_28446,N_27736);
and UO_2648 (O_2648,N_28484,N_29586);
or UO_2649 (O_2649,N_27942,N_27067);
nor UO_2650 (O_2650,N_27589,N_29605);
or UO_2651 (O_2651,N_28530,N_28894);
or UO_2652 (O_2652,N_28905,N_29276);
xnor UO_2653 (O_2653,N_28443,N_28350);
or UO_2654 (O_2654,N_28504,N_27293);
xnor UO_2655 (O_2655,N_29914,N_29529);
nand UO_2656 (O_2656,N_29575,N_29364);
nand UO_2657 (O_2657,N_28550,N_29784);
or UO_2658 (O_2658,N_27663,N_27429);
xor UO_2659 (O_2659,N_27068,N_29690);
or UO_2660 (O_2660,N_29950,N_27580);
xor UO_2661 (O_2661,N_28700,N_29378);
xor UO_2662 (O_2662,N_29336,N_28806);
nand UO_2663 (O_2663,N_29626,N_29402);
nor UO_2664 (O_2664,N_29364,N_28081);
nor UO_2665 (O_2665,N_29533,N_29023);
xor UO_2666 (O_2666,N_28486,N_29748);
and UO_2667 (O_2667,N_28222,N_28782);
nor UO_2668 (O_2668,N_27060,N_29986);
nor UO_2669 (O_2669,N_27361,N_29808);
xor UO_2670 (O_2670,N_28825,N_28282);
and UO_2671 (O_2671,N_27961,N_29270);
nor UO_2672 (O_2672,N_28815,N_27759);
and UO_2673 (O_2673,N_27732,N_27079);
nand UO_2674 (O_2674,N_27497,N_29480);
xor UO_2675 (O_2675,N_29496,N_28165);
xnor UO_2676 (O_2676,N_27024,N_27547);
nor UO_2677 (O_2677,N_28742,N_28918);
nand UO_2678 (O_2678,N_27262,N_29255);
nand UO_2679 (O_2679,N_27988,N_29712);
nor UO_2680 (O_2680,N_29601,N_28200);
or UO_2681 (O_2681,N_28024,N_28092);
or UO_2682 (O_2682,N_27357,N_27023);
and UO_2683 (O_2683,N_29740,N_28444);
nand UO_2684 (O_2684,N_28503,N_27228);
nand UO_2685 (O_2685,N_28020,N_27185);
xor UO_2686 (O_2686,N_27676,N_28005);
nor UO_2687 (O_2687,N_28160,N_28706);
xor UO_2688 (O_2688,N_29851,N_29160);
and UO_2689 (O_2689,N_29705,N_27027);
xnor UO_2690 (O_2690,N_29870,N_28309);
nand UO_2691 (O_2691,N_29115,N_29084);
xnor UO_2692 (O_2692,N_27710,N_28075);
nor UO_2693 (O_2693,N_29526,N_28478);
nor UO_2694 (O_2694,N_28620,N_27327);
nand UO_2695 (O_2695,N_29891,N_29587);
and UO_2696 (O_2696,N_29287,N_28966);
xnor UO_2697 (O_2697,N_27364,N_28935);
xor UO_2698 (O_2698,N_27728,N_29479);
nand UO_2699 (O_2699,N_27803,N_27204);
xor UO_2700 (O_2700,N_29904,N_29819);
or UO_2701 (O_2701,N_29451,N_29870);
nor UO_2702 (O_2702,N_29860,N_29575);
nor UO_2703 (O_2703,N_29138,N_28386);
or UO_2704 (O_2704,N_27654,N_28986);
or UO_2705 (O_2705,N_28046,N_29520);
and UO_2706 (O_2706,N_28783,N_27732);
and UO_2707 (O_2707,N_27700,N_28123);
and UO_2708 (O_2708,N_27546,N_29564);
nand UO_2709 (O_2709,N_27627,N_28881);
or UO_2710 (O_2710,N_27948,N_29489);
and UO_2711 (O_2711,N_27284,N_29421);
and UO_2712 (O_2712,N_28094,N_27134);
xor UO_2713 (O_2713,N_27717,N_29415);
nand UO_2714 (O_2714,N_29049,N_28359);
and UO_2715 (O_2715,N_27880,N_27272);
or UO_2716 (O_2716,N_29940,N_29163);
or UO_2717 (O_2717,N_28604,N_28425);
nor UO_2718 (O_2718,N_27742,N_27763);
xor UO_2719 (O_2719,N_29941,N_27282);
nand UO_2720 (O_2720,N_27262,N_27843);
or UO_2721 (O_2721,N_29799,N_27311);
nor UO_2722 (O_2722,N_29754,N_29788);
nand UO_2723 (O_2723,N_27183,N_27972);
xnor UO_2724 (O_2724,N_28857,N_27849);
nand UO_2725 (O_2725,N_27061,N_29819);
nand UO_2726 (O_2726,N_28479,N_28525);
xnor UO_2727 (O_2727,N_29169,N_27704);
nor UO_2728 (O_2728,N_28875,N_27627);
or UO_2729 (O_2729,N_27332,N_29998);
nand UO_2730 (O_2730,N_29792,N_28666);
nor UO_2731 (O_2731,N_27580,N_29646);
nor UO_2732 (O_2732,N_28405,N_28764);
nor UO_2733 (O_2733,N_29387,N_28609);
nand UO_2734 (O_2734,N_27768,N_29056);
or UO_2735 (O_2735,N_28265,N_29532);
or UO_2736 (O_2736,N_28976,N_28887);
xnor UO_2737 (O_2737,N_29325,N_29257);
nor UO_2738 (O_2738,N_27390,N_27261);
or UO_2739 (O_2739,N_27091,N_29981);
xor UO_2740 (O_2740,N_29147,N_29539);
and UO_2741 (O_2741,N_29738,N_29002);
and UO_2742 (O_2742,N_28164,N_29159);
nor UO_2743 (O_2743,N_29808,N_28623);
xor UO_2744 (O_2744,N_28004,N_27789);
and UO_2745 (O_2745,N_29451,N_27173);
and UO_2746 (O_2746,N_27019,N_28095);
nand UO_2747 (O_2747,N_27565,N_29267);
nand UO_2748 (O_2748,N_27557,N_28241);
nand UO_2749 (O_2749,N_28547,N_27847);
and UO_2750 (O_2750,N_29089,N_28946);
and UO_2751 (O_2751,N_29503,N_29695);
and UO_2752 (O_2752,N_27920,N_28068);
nand UO_2753 (O_2753,N_29832,N_29376);
or UO_2754 (O_2754,N_28306,N_27206);
xor UO_2755 (O_2755,N_29002,N_29015);
nor UO_2756 (O_2756,N_28516,N_28371);
or UO_2757 (O_2757,N_27268,N_28048);
and UO_2758 (O_2758,N_27141,N_28106);
and UO_2759 (O_2759,N_29971,N_27798);
or UO_2760 (O_2760,N_29040,N_28723);
xnor UO_2761 (O_2761,N_28788,N_27558);
or UO_2762 (O_2762,N_27535,N_28836);
or UO_2763 (O_2763,N_27744,N_27096);
and UO_2764 (O_2764,N_27911,N_27466);
xnor UO_2765 (O_2765,N_27213,N_29864);
and UO_2766 (O_2766,N_27156,N_27404);
xnor UO_2767 (O_2767,N_28313,N_29581);
and UO_2768 (O_2768,N_28216,N_28896);
and UO_2769 (O_2769,N_27540,N_28127);
nor UO_2770 (O_2770,N_28854,N_29823);
nor UO_2771 (O_2771,N_29098,N_29131);
or UO_2772 (O_2772,N_29091,N_28482);
nor UO_2773 (O_2773,N_27315,N_27361);
nor UO_2774 (O_2774,N_27194,N_27442);
nor UO_2775 (O_2775,N_29011,N_28120);
xnor UO_2776 (O_2776,N_28082,N_28734);
xnor UO_2777 (O_2777,N_29633,N_27470);
xor UO_2778 (O_2778,N_28875,N_27849);
or UO_2779 (O_2779,N_27979,N_29399);
or UO_2780 (O_2780,N_28564,N_27955);
nor UO_2781 (O_2781,N_29884,N_27063);
nand UO_2782 (O_2782,N_27852,N_27607);
xor UO_2783 (O_2783,N_27671,N_29852);
or UO_2784 (O_2784,N_27325,N_27921);
nand UO_2785 (O_2785,N_27554,N_29474);
nor UO_2786 (O_2786,N_29682,N_29788);
xor UO_2787 (O_2787,N_29812,N_27200);
nor UO_2788 (O_2788,N_29025,N_29132);
and UO_2789 (O_2789,N_27160,N_29234);
xnor UO_2790 (O_2790,N_29927,N_27954);
nor UO_2791 (O_2791,N_29906,N_28274);
xor UO_2792 (O_2792,N_27646,N_29535);
and UO_2793 (O_2793,N_27956,N_29069);
or UO_2794 (O_2794,N_27738,N_29851);
xor UO_2795 (O_2795,N_29203,N_29319);
and UO_2796 (O_2796,N_28448,N_29688);
or UO_2797 (O_2797,N_27500,N_28034);
or UO_2798 (O_2798,N_27132,N_27772);
or UO_2799 (O_2799,N_27054,N_28877);
or UO_2800 (O_2800,N_27078,N_28136);
nand UO_2801 (O_2801,N_29666,N_27558);
nand UO_2802 (O_2802,N_28434,N_29946);
and UO_2803 (O_2803,N_28520,N_28263);
nor UO_2804 (O_2804,N_27344,N_28828);
or UO_2805 (O_2805,N_29779,N_29930);
xor UO_2806 (O_2806,N_28560,N_27149);
nand UO_2807 (O_2807,N_28379,N_27221);
and UO_2808 (O_2808,N_27232,N_28034);
xor UO_2809 (O_2809,N_28278,N_28753);
nor UO_2810 (O_2810,N_27261,N_29205);
nand UO_2811 (O_2811,N_29525,N_28239);
or UO_2812 (O_2812,N_27609,N_27125);
xor UO_2813 (O_2813,N_29017,N_28323);
and UO_2814 (O_2814,N_28346,N_29372);
or UO_2815 (O_2815,N_27814,N_27520);
or UO_2816 (O_2816,N_29041,N_28661);
nor UO_2817 (O_2817,N_27228,N_28671);
or UO_2818 (O_2818,N_27432,N_29217);
nor UO_2819 (O_2819,N_29786,N_29244);
xnor UO_2820 (O_2820,N_27207,N_27955);
or UO_2821 (O_2821,N_27048,N_29696);
nor UO_2822 (O_2822,N_28751,N_29731);
and UO_2823 (O_2823,N_29826,N_28534);
xnor UO_2824 (O_2824,N_28402,N_29057);
xnor UO_2825 (O_2825,N_27417,N_27813);
or UO_2826 (O_2826,N_28069,N_28525);
xnor UO_2827 (O_2827,N_27576,N_29432);
nand UO_2828 (O_2828,N_29731,N_28447);
nand UO_2829 (O_2829,N_29182,N_29044);
xor UO_2830 (O_2830,N_28522,N_28400);
xor UO_2831 (O_2831,N_28099,N_29528);
nor UO_2832 (O_2832,N_29637,N_29347);
xnor UO_2833 (O_2833,N_27782,N_29239);
or UO_2834 (O_2834,N_28431,N_29407);
and UO_2835 (O_2835,N_28968,N_27504);
or UO_2836 (O_2836,N_27967,N_29299);
or UO_2837 (O_2837,N_29858,N_28580);
nand UO_2838 (O_2838,N_27741,N_28516);
nor UO_2839 (O_2839,N_28831,N_27907);
or UO_2840 (O_2840,N_27003,N_29592);
nand UO_2841 (O_2841,N_28344,N_27879);
nand UO_2842 (O_2842,N_28026,N_29120);
nor UO_2843 (O_2843,N_28308,N_29009);
nor UO_2844 (O_2844,N_28182,N_28021);
xor UO_2845 (O_2845,N_28502,N_27372);
nor UO_2846 (O_2846,N_29905,N_29398);
nand UO_2847 (O_2847,N_28538,N_28914);
xnor UO_2848 (O_2848,N_29470,N_28430);
and UO_2849 (O_2849,N_28277,N_29565);
nor UO_2850 (O_2850,N_29914,N_29067);
xnor UO_2851 (O_2851,N_28615,N_27277);
xor UO_2852 (O_2852,N_29768,N_29249);
nor UO_2853 (O_2853,N_27338,N_27493);
and UO_2854 (O_2854,N_29348,N_27268);
or UO_2855 (O_2855,N_28002,N_27483);
nand UO_2856 (O_2856,N_29327,N_29125);
or UO_2857 (O_2857,N_27957,N_27038);
and UO_2858 (O_2858,N_28388,N_27771);
nand UO_2859 (O_2859,N_28781,N_27220);
or UO_2860 (O_2860,N_28549,N_27714);
or UO_2861 (O_2861,N_28704,N_29989);
nand UO_2862 (O_2862,N_28915,N_28270);
nor UO_2863 (O_2863,N_29914,N_29251);
and UO_2864 (O_2864,N_28265,N_29924);
nor UO_2865 (O_2865,N_29433,N_27049);
nor UO_2866 (O_2866,N_27803,N_27243);
nand UO_2867 (O_2867,N_29809,N_28752);
and UO_2868 (O_2868,N_27380,N_29123);
nor UO_2869 (O_2869,N_29983,N_27682);
and UO_2870 (O_2870,N_27460,N_27658);
and UO_2871 (O_2871,N_29896,N_28751);
nor UO_2872 (O_2872,N_27596,N_29631);
xor UO_2873 (O_2873,N_28090,N_29623);
nand UO_2874 (O_2874,N_28012,N_29764);
and UO_2875 (O_2875,N_28859,N_28885);
nor UO_2876 (O_2876,N_28906,N_29294);
nor UO_2877 (O_2877,N_29575,N_29139);
nand UO_2878 (O_2878,N_28733,N_27359);
nor UO_2879 (O_2879,N_29868,N_29324);
or UO_2880 (O_2880,N_28654,N_29892);
and UO_2881 (O_2881,N_27610,N_28159);
nand UO_2882 (O_2882,N_29082,N_29369);
xor UO_2883 (O_2883,N_27013,N_29678);
or UO_2884 (O_2884,N_27662,N_29436);
nand UO_2885 (O_2885,N_29710,N_29309);
nand UO_2886 (O_2886,N_27462,N_28178);
nand UO_2887 (O_2887,N_28568,N_29400);
and UO_2888 (O_2888,N_29426,N_28945);
nor UO_2889 (O_2889,N_28124,N_28601);
and UO_2890 (O_2890,N_27306,N_28699);
or UO_2891 (O_2891,N_28174,N_27708);
xor UO_2892 (O_2892,N_27072,N_27224);
nand UO_2893 (O_2893,N_29138,N_28509);
or UO_2894 (O_2894,N_28810,N_27499);
and UO_2895 (O_2895,N_28627,N_29946);
nor UO_2896 (O_2896,N_27852,N_28897);
xor UO_2897 (O_2897,N_28799,N_29606);
nand UO_2898 (O_2898,N_27001,N_27782);
and UO_2899 (O_2899,N_27494,N_27937);
nand UO_2900 (O_2900,N_27586,N_28757);
or UO_2901 (O_2901,N_28222,N_28828);
nand UO_2902 (O_2902,N_27935,N_28338);
nand UO_2903 (O_2903,N_29967,N_29750);
nand UO_2904 (O_2904,N_28198,N_27536);
nand UO_2905 (O_2905,N_28856,N_29261);
nor UO_2906 (O_2906,N_27875,N_28986);
xor UO_2907 (O_2907,N_29535,N_29717);
nor UO_2908 (O_2908,N_27015,N_27256);
and UO_2909 (O_2909,N_27682,N_28593);
and UO_2910 (O_2910,N_28812,N_29326);
or UO_2911 (O_2911,N_29574,N_27831);
xor UO_2912 (O_2912,N_27972,N_29280);
and UO_2913 (O_2913,N_27225,N_28090);
and UO_2914 (O_2914,N_27597,N_28439);
nand UO_2915 (O_2915,N_27519,N_29673);
or UO_2916 (O_2916,N_28580,N_29848);
and UO_2917 (O_2917,N_27218,N_27285);
and UO_2918 (O_2918,N_27805,N_28578);
or UO_2919 (O_2919,N_28251,N_27596);
or UO_2920 (O_2920,N_27279,N_29201);
or UO_2921 (O_2921,N_29392,N_28350);
and UO_2922 (O_2922,N_27334,N_27497);
or UO_2923 (O_2923,N_29592,N_27142);
nand UO_2924 (O_2924,N_29026,N_29387);
and UO_2925 (O_2925,N_28650,N_28081);
xor UO_2926 (O_2926,N_29598,N_27734);
and UO_2927 (O_2927,N_28589,N_28498);
nor UO_2928 (O_2928,N_27270,N_27720);
xor UO_2929 (O_2929,N_28294,N_28766);
and UO_2930 (O_2930,N_28135,N_29518);
nand UO_2931 (O_2931,N_27878,N_29522);
and UO_2932 (O_2932,N_27137,N_29500);
xor UO_2933 (O_2933,N_27495,N_27605);
xnor UO_2934 (O_2934,N_27156,N_29981);
nand UO_2935 (O_2935,N_28777,N_27574);
nor UO_2936 (O_2936,N_28742,N_27125);
and UO_2937 (O_2937,N_28840,N_29859);
and UO_2938 (O_2938,N_28664,N_29048);
or UO_2939 (O_2939,N_29578,N_29684);
and UO_2940 (O_2940,N_29027,N_28290);
or UO_2941 (O_2941,N_29359,N_27119);
or UO_2942 (O_2942,N_27560,N_28684);
or UO_2943 (O_2943,N_27376,N_29036);
xor UO_2944 (O_2944,N_27712,N_29653);
nor UO_2945 (O_2945,N_27350,N_28505);
nand UO_2946 (O_2946,N_27706,N_28871);
nand UO_2947 (O_2947,N_27947,N_29197);
or UO_2948 (O_2948,N_29329,N_28851);
nor UO_2949 (O_2949,N_27317,N_27895);
xor UO_2950 (O_2950,N_28419,N_28822);
nand UO_2951 (O_2951,N_27131,N_29869);
nand UO_2952 (O_2952,N_28144,N_27736);
nand UO_2953 (O_2953,N_29439,N_29272);
xnor UO_2954 (O_2954,N_27260,N_29707);
or UO_2955 (O_2955,N_29971,N_29370);
and UO_2956 (O_2956,N_28941,N_28173);
nor UO_2957 (O_2957,N_28792,N_28986);
and UO_2958 (O_2958,N_29759,N_28659);
or UO_2959 (O_2959,N_29479,N_29748);
nand UO_2960 (O_2960,N_29210,N_27023);
nand UO_2961 (O_2961,N_29284,N_29254);
and UO_2962 (O_2962,N_28647,N_29732);
or UO_2963 (O_2963,N_29277,N_28734);
nor UO_2964 (O_2964,N_27817,N_28784);
xnor UO_2965 (O_2965,N_27239,N_27232);
nand UO_2966 (O_2966,N_27835,N_29775);
or UO_2967 (O_2967,N_29707,N_27538);
nand UO_2968 (O_2968,N_29865,N_29739);
nand UO_2969 (O_2969,N_27446,N_27003);
or UO_2970 (O_2970,N_27115,N_29417);
xor UO_2971 (O_2971,N_28704,N_28012);
xor UO_2972 (O_2972,N_27247,N_29407);
or UO_2973 (O_2973,N_28924,N_29651);
and UO_2974 (O_2974,N_29178,N_28078);
nand UO_2975 (O_2975,N_28011,N_27938);
nor UO_2976 (O_2976,N_29078,N_29164);
xor UO_2977 (O_2977,N_28337,N_29692);
xor UO_2978 (O_2978,N_27169,N_29256);
or UO_2979 (O_2979,N_29629,N_28734);
or UO_2980 (O_2980,N_29469,N_28876);
xor UO_2981 (O_2981,N_27165,N_27852);
nor UO_2982 (O_2982,N_27573,N_29602);
nand UO_2983 (O_2983,N_28803,N_29608);
xnor UO_2984 (O_2984,N_29998,N_28837);
or UO_2985 (O_2985,N_29901,N_27255);
or UO_2986 (O_2986,N_29879,N_27421);
nor UO_2987 (O_2987,N_29904,N_29871);
xnor UO_2988 (O_2988,N_29418,N_29121);
xor UO_2989 (O_2989,N_27696,N_29077);
nor UO_2990 (O_2990,N_27285,N_28710);
or UO_2991 (O_2991,N_27004,N_27423);
nor UO_2992 (O_2992,N_28984,N_27165);
or UO_2993 (O_2993,N_28688,N_28838);
and UO_2994 (O_2994,N_27219,N_29664);
xor UO_2995 (O_2995,N_27189,N_29372);
and UO_2996 (O_2996,N_27502,N_28032);
or UO_2997 (O_2997,N_29778,N_29982);
and UO_2998 (O_2998,N_28285,N_28539);
and UO_2999 (O_2999,N_28289,N_28374);
or UO_3000 (O_3000,N_28610,N_28192);
nor UO_3001 (O_3001,N_27332,N_29194);
or UO_3002 (O_3002,N_29897,N_28569);
nor UO_3003 (O_3003,N_29895,N_28530);
xnor UO_3004 (O_3004,N_29613,N_27288);
or UO_3005 (O_3005,N_28614,N_27852);
nor UO_3006 (O_3006,N_28099,N_29190);
and UO_3007 (O_3007,N_29966,N_28555);
or UO_3008 (O_3008,N_27695,N_29502);
nor UO_3009 (O_3009,N_29430,N_29588);
and UO_3010 (O_3010,N_28853,N_28751);
and UO_3011 (O_3011,N_27228,N_28970);
xor UO_3012 (O_3012,N_28160,N_27684);
or UO_3013 (O_3013,N_29543,N_28759);
xnor UO_3014 (O_3014,N_28815,N_27765);
or UO_3015 (O_3015,N_29591,N_28015);
and UO_3016 (O_3016,N_27088,N_27593);
nor UO_3017 (O_3017,N_28710,N_29555);
or UO_3018 (O_3018,N_28418,N_27478);
nor UO_3019 (O_3019,N_29159,N_28284);
nand UO_3020 (O_3020,N_28302,N_28843);
or UO_3021 (O_3021,N_28899,N_28947);
nand UO_3022 (O_3022,N_27477,N_29374);
nor UO_3023 (O_3023,N_29097,N_27854);
xnor UO_3024 (O_3024,N_29818,N_27608);
xnor UO_3025 (O_3025,N_28999,N_27896);
or UO_3026 (O_3026,N_27096,N_28151);
nand UO_3027 (O_3027,N_27921,N_29077);
nor UO_3028 (O_3028,N_27060,N_29977);
nor UO_3029 (O_3029,N_29601,N_27027);
or UO_3030 (O_3030,N_29542,N_28164);
xnor UO_3031 (O_3031,N_27800,N_28768);
or UO_3032 (O_3032,N_28318,N_27458);
and UO_3033 (O_3033,N_27341,N_28342);
or UO_3034 (O_3034,N_27166,N_27291);
nand UO_3035 (O_3035,N_28019,N_29808);
xor UO_3036 (O_3036,N_29610,N_29617);
xor UO_3037 (O_3037,N_28801,N_29607);
or UO_3038 (O_3038,N_28399,N_28103);
xor UO_3039 (O_3039,N_28053,N_28916);
and UO_3040 (O_3040,N_29690,N_27398);
nor UO_3041 (O_3041,N_28887,N_29532);
xor UO_3042 (O_3042,N_28224,N_29064);
xnor UO_3043 (O_3043,N_27639,N_27064);
xor UO_3044 (O_3044,N_29282,N_29379);
nor UO_3045 (O_3045,N_27935,N_27868);
xor UO_3046 (O_3046,N_28609,N_27823);
and UO_3047 (O_3047,N_28534,N_27631);
or UO_3048 (O_3048,N_29353,N_27321);
nor UO_3049 (O_3049,N_27949,N_29606);
and UO_3050 (O_3050,N_29745,N_29667);
xor UO_3051 (O_3051,N_29566,N_28205);
or UO_3052 (O_3052,N_27068,N_29219);
nor UO_3053 (O_3053,N_27248,N_28759);
nor UO_3054 (O_3054,N_29116,N_29281);
nand UO_3055 (O_3055,N_29041,N_29548);
nand UO_3056 (O_3056,N_28686,N_27452);
nor UO_3057 (O_3057,N_28666,N_28939);
nand UO_3058 (O_3058,N_27527,N_29639);
xor UO_3059 (O_3059,N_27251,N_27924);
and UO_3060 (O_3060,N_28254,N_28468);
or UO_3061 (O_3061,N_28907,N_29338);
and UO_3062 (O_3062,N_28854,N_28959);
nand UO_3063 (O_3063,N_29369,N_28543);
or UO_3064 (O_3064,N_27542,N_28420);
xor UO_3065 (O_3065,N_28536,N_29281);
xnor UO_3066 (O_3066,N_27416,N_28087);
and UO_3067 (O_3067,N_27407,N_29582);
nor UO_3068 (O_3068,N_29843,N_27843);
xor UO_3069 (O_3069,N_29477,N_27822);
nor UO_3070 (O_3070,N_29868,N_27733);
xor UO_3071 (O_3071,N_28688,N_28152);
nor UO_3072 (O_3072,N_28696,N_28994);
or UO_3073 (O_3073,N_27058,N_28699);
and UO_3074 (O_3074,N_28951,N_28668);
or UO_3075 (O_3075,N_27469,N_29020);
and UO_3076 (O_3076,N_28219,N_29372);
xnor UO_3077 (O_3077,N_28352,N_28852);
or UO_3078 (O_3078,N_28005,N_27179);
nor UO_3079 (O_3079,N_27920,N_29379);
xor UO_3080 (O_3080,N_28236,N_27343);
nand UO_3081 (O_3081,N_27239,N_28718);
nor UO_3082 (O_3082,N_28208,N_29893);
nand UO_3083 (O_3083,N_27235,N_29935);
nor UO_3084 (O_3084,N_29682,N_27237);
nand UO_3085 (O_3085,N_29717,N_27357);
nand UO_3086 (O_3086,N_28808,N_27471);
and UO_3087 (O_3087,N_29368,N_28770);
nand UO_3088 (O_3088,N_29211,N_29341);
xor UO_3089 (O_3089,N_29383,N_29685);
and UO_3090 (O_3090,N_27807,N_29721);
or UO_3091 (O_3091,N_29441,N_29435);
and UO_3092 (O_3092,N_27553,N_28157);
nand UO_3093 (O_3093,N_28746,N_28706);
or UO_3094 (O_3094,N_29008,N_29995);
or UO_3095 (O_3095,N_29896,N_28210);
and UO_3096 (O_3096,N_28186,N_29225);
and UO_3097 (O_3097,N_27351,N_29991);
xnor UO_3098 (O_3098,N_29618,N_29622);
or UO_3099 (O_3099,N_27419,N_27797);
and UO_3100 (O_3100,N_27494,N_29329);
xnor UO_3101 (O_3101,N_28376,N_27103);
xor UO_3102 (O_3102,N_28499,N_28745);
or UO_3103 (O_3103,N_28713,N_29852);
nor UO_3104 (O_3104,N_28170,N_28565);
nor UO_3105 (O_3105,N_27410,N_28632);
xor UO_3106 (O_3106,N_28456,N_29199);
nand UO_3107 (O_3107,N_27000,N_29085);
or UO_3108 (O_3108,N_29165,N_28815);
nor UO_3109 (O_3109,N_28834,N_29204);
nand UO_3110 (O_3110,N_27212,N_29965);
xor UO_3111 (O_3111,N_29986,N_29703);
nand UO_3112 (O_3112,N_27965,N_27036);
or UO_3113 (O_3113,N_28688,N_28013);
or UO_3114 (O_3114,N_27793,N_29689);
xnor UO_3115 (O_3115,N_29116,N_28410);
and UO_3116 (O_3116,N_28407,N_29319);
and UO_3117 (O_3117,N_27513,N_27441);
nor UO_3118 (O_3118,N_28992,N_29971);
nor UO_3119 (O_3119,N_28468,N_27809);
and UO_3120 (O_3120,N_28773,N_28599);
or UO_3121 (O_3121,N_27911,N_28733);
nand UO_3122 (O_3122,N_29054,N_27587);
nor UO_3123 (O_3123,N_27445,N_29084);
or UO_3124 (O_3124,N_29989,N_27067);
nor UO_3125 (O_3125,N_27786,N_27814);
or UO_3126 (O_3126,N_28730,N_29835);
nand UO_3127 (O_3127,N_29726,N_28708);
nor UO_3128 (O_3128,N_29608,N_27734);
nor UO_3129 (O_3129,N_28256,N_28055);
nand UO_3130 (O_3130,N_29670,N_28079);
or UO_3131 (O_3131,N_28317,N_28822);
nand UO_3132 (O_3132,N_28309,N_28987);
and UO_3133 (O_3133,N_29364,N_28565);
xor UO_3134 (O_3134,N_28739,N_28032);
or UO_3135 (O_3135,N_29302,N_29065);
or UO_3136 (O_3136,N_29950,N_29332);
and UO_3137 (O_3137,N_28927,N_27159);
xor UO_3138 (O_3138,N_28073,N_29009);
xor UO_3139 (O_3139,N_29065,N_28419);
or UO_3140 (O_3140,N_29676,N_29070);
xor UO_3141 (O_3141,N_27728,N_27912);
and UO_3142 (O_3142,N_29066,N_29626);
or UO_3143 (O_3143,N_28695,N_28623);
xnor UO_3144 (O_3144,N_27835,N_29230);
nand UO_3145 (O_3145,N_27344,N_27678);
or UO_3146 (O_3146,N_27225,N_28639);
and UO_3147 (O_3147,N_27745,N_29024);
nand UO_3148 (O_3148,N_28664,N_28803);
nor UO_3149 (O_3149,N_28330,N_28283);
or UO_3150 (O_3150,N_28846,N_27064);
or UO_3151 (O_3151,N_27350,N_27453);
or UO_3152 (O_3152,N_27498,N_28013);
or UO_3153 (O_3153,N_28074,N_29497);
or UO_3154 (O_3154,N_27212,N_29028);
xor UO_3155 (O_3155,N_28183,N_27738);
xnor UO_3156 (O_3156,N_27953,N_28191);
or UO_3157 (O_3157,N_29067,N_28688);
nor UO_3158 (O_3158,N_27378,N_29819);
or UO_3159 (O_3159,N_29182,N_27489);
or UO_3160 (O_3160,N_27411,N_28454);
and UO_3161 (O_3161,N_28046,N_28985);
and UO_3162 (O_3162,N_29294,N_29177);
and UO_3163 (O_3163,N_29226,N_27638);
xor UO_3164 (O_3164,N_28652,N_27681);
or UO_3165 (O_3165,N_27301,N_29619);
or UO_3166 (O_3166,N_27498,N_29086);
xor UO_3167 (O_3167,N_27696,N_29463);
xnor UO_3168 (O_3168,N_27310,N_28141);
and UO_3169 (O_3169,N_27452,N_27206);
nor UO_3170 (O_3170,N_27242,N_27446);
nand UO_3171 (O_3171,N_29118,N_28686);
or UO_3172 (O_3172,N_28290,N_29404);
xor UO_3173 (O_3173,N_29927,N_28879);
and UO_3174 (O_3174,N_27252,N_28781);
or UO_3175 (O_3175,N_29517,N_29241);
nand UO_3176 (O_3176,N_27060,N_27421);
and UO_3177 (O_3177,N_27677,N_28562);
xnor UO_3178 (O_3178,N_28583,N_27856);
or UO_3179 (O_3179,N_27171,N_27452);
and UO_3180 (O_3180,N_27507,N_27138);
nand UO_3181 (O_3181,N_28634,N_27229);
nor UO_3182 (O_3182,N_28938,N_27725);
nand UO_3183 (O_3183,N_29038,N_27222);
nand UO_3184 (O_3184,N_29689,N_27374);
nor UO_3185 (O_3185,N_27446,N_28132);
nand UO_3186 (O_3186,N_29529,N_29139);
nor UO_3187 (O_3187,N_29197,N_29190);
nor UO_3188 (O_3188,N_28093,N_29455);
nand UO_3189 (O_3189,N_27852,N_29717);
nor UO_3190 (O_3190,N_28226,N_27824);
and UO_3191 (O_3191,N_27847,N_27690);
and UO_3192 (O_3192,N_27351,N_27730);
and UO_3193 (O_3193,N_28818,N_28998);
and UO_3194 (O_3194,N_28835,N_27084);
nor UO_3195 (O_3195,N_28048,N_27063);
or UO_3196 (O_3196,N_29444,N_27584);
and UO_3197 (O_3197,N_28893,N_29777);
and UO_3198 (O_3198,N_27030,N_28191);
nor UO_3199 (O_3199,N_29563,N_28730);
or UO_3200 (O_3200,N_27497,N_29667);
nor UO_3201 (O_3201,N_29430,N_27378);
nor UO_3202 (O_3202,N_29890,N_29845);
and UO_3203 (O_3203,N_28095,N_29167);
or UO_3204 (O_3204,N_27761,N_27075);
xnor UO_3205 (O_3205,N_28557,N_28077);
xnor UO_3206 (O_3206,N_28661,N_29800);
and UO_3207 (O_3207,N_27801,N_27638);
nand UO_3208 (O_3208,N_27443,N_29708);
nand UO_3209 (O_3209,N_27224,N_29809);
and UO_3210 (O_3210,N_28441,N_27437);
and UO_3211 (O_3211,N_28958,N_27625);
or UO_3212 (O_3212,N_29744,N_28068);
and UO_3213 (O_3213,N_27119,N_27818);
or UO_3214 (O_3214,N_28916,N_27009);
xor UO_3215 (O_3215,N_28447,N_28689);
nor UO_3216 (O_3216,N_27187,N_29828);
nand UO_3217 (O_3217,N_28427,N_29107);
nor UO_3218 (O_3218,N_27035,N_29903);
and UO_3219 (O_3219,N_29021,N_28809);
nand UO_3220 (O_3220,N_27395,N_28430);
xor UO_3221 (O_3221,N_29074,N_27508);
xor UO_3222 (O_3222,N_29003,N_27845);
xnor UO_3223 (O_3223,N_28733,N_28576);
or UO_3224 (O_3224,N_29040,N_29127);
and UO_3225 (O_3225,N_27422,N_29550);
nand UO_3226 (O_3226,N_27744,N_28714);
nand UO_3227 (O_3227,N_27713,N_29053);
xnor UO_3228 (O_3228,N_28225,N_29476);
nor UO_3229 (O_3229,N_28046,N_29912);
xnor UO_3230 (O_3230,N_28561,N_27122);
or UO_3231 (O_3231,N_29215,N_27890);
and UO_3232 (O_3232,N_28120,N_28303);
nor UO_3233 (O_3233,N_29943,N_29348);
nand UO_3234 (O_3234,N_29017,N_28981);
xor UO_3235 (O_3235,N_29305,N_27430);
or UO_3236 (O_3236,N_27878,N_27702);
nand UO_3237 (O_3237,N_27276,N_29983);
nor UO_3238 (O_3238,N_27273,N_28475);
and UO_3239 (O_3239,N_27649,N_29057);
and UO_3240 (O_3240,N_29081,N_28740);
or UO_3241 (O_3241,N_27587,N_29620);
and UO_3242 (O_3242,N_27513,N_27538);
or UO_3243 (O_3243,N_28933,N_29374);
xnor UO_3244 (O_3244,N_29976,N_29535);
nor UO_3245 (O_3245,N_28215,N_28828);
nand UO_3246 (O_3246,N_28829,N_27917);
xor UO_3247 (O_3247,N_27955,N_28387);
nor UO_3248 (O_3248,N_29733,N_27968);
or UO_3249 (O_3249,N_29968,N_27975);
nor UO_3250 (O_3250,N_28832,N_28410);
nor UO_3251 (O_3251,N_29531,N_29367);
and UO_3252 (O_3252,N_29454,N_27023);
or UO_3253 (O_3253,N_29770,N_29875);
nor UO_3254 (O_3254,N_27963,N_27325);
and UO_3255 (O_3255,N_27165,N_27970);
nor UO_3256 (O_3256,N_28590,N_27986);
xor UO_3257 (O_3257,N_28557,N_29650);
nor UO_3258 (O_3258,N_29761,N_29246);
and UO_3259 (O_3259,N_29202,N_28603);
nand UO_3260 (O_3260,N_27581,N_27280);
nand UO_3261 (O_3261,N_27127,N_29372);
or UO_3262 (O_3262,N_29387,N_28396);
xnor UO_3263 (O_3263,N_29027,N_28810);
xnor UO_3264 (O_3264,N_28184,N_29237);
nand UO_3265 (O_3265,N_29421,N_28979);
or UO_3266 (O_3266,N_28620,N_28660);
nor UO_3267 (O_3267,N_27826,N_28316);
or UO_3268 (O_3268,N_28946,N_27124);
nor UO_3269 (O_3269,N_27751,N_27337);
nor UO_3270 (O_3270,N_27245,N_28074);
nand UO_3271 (O_3271,N_29527,N_29438);
nor UO_3272 (O_3272,N_28389,N_28547);
and UO_3273 (O_3273,N_27186,N_29011);
nand UO_3274 (O_3274,N_28086,N_28595);
and UO_3275 (O_3275,N_28594,N_28985);
and UO_3276 (O_3276,N_27268,N_27256);
or UO_3277 (O_3277,N_28109,N_28383);
xnor UO_3278 (O_3278,N_28282,N_29321);
or UO_3279 (O_3279,N_28281,N_29251);
nor UO_3280 (O_3280,N_28020,N_27352);
nand UO_3281 (O_3281,N_29694,N_28042);
nor UO_3282 (O_3282,N_27456,N_28575);
and UO_3283 (O_3283,N_29511,N_27927);
and UO_3284 (O_3284,N_29633,N_29095);
xor UO_3285 (O_3285,N_27337,N_27818);
and UO_3286 (O_3286,N_29207,N_29852);
and UO_3287 (O_3287,N_29559,N_28417);
nor UO_3288 (O_3288,N_29434,N_29945);
nand UO_3289 (O_3289,N_29642,N_29263);
and UO_3290 (O_3290,N_27510,N_29294);
or UO_3291 (O_3291,N_27137,N_28429);
or UO_3292 (O_3292,N_29265,N_28010);
and UO_3293 (O_3293,N_27826,N_27384);
nor UO_3294 (O_3294,N_27956,N_29193);
nand UO_3295 (O_3295,N_27895,N_28826);
and UO_3296 (O_3296,N_29081,N_27441);
and UO_3297 (O_3297,N_27319,N_29578);
nand UO_3298 (O_3298,N_28517,N_27187);
xnor UO_3299 (O_3299,N_27226,N_29017);
nor UO_3300 (O_3300,N_29763,N_27106);
nor UO_3301 (O_3301,N_27881,N_29447);
xnor UO_3302 (O_3302,N_29652,N_27833);
xor UO_3303 (O_3303,N_29117,N_29624);
xor UO_3304 (O_3304,N_28738,N_27196);
xor UO_3305 (O_3305,N_29440,N_28856);
nor UO_3306 (O_3306,N_29947,N_29044);
and UO_3307 (O_3307,N_29031,N_28230);
xor UO_3308 (O_3308,N_27461,N_28803);
xnor UO_3309 (O_3309,N_29480,N_29007);
nor UO_3310 (O_3310,N_28975,N_29956);
nand UO_3311 (O_3311,N_27236,N_29773);
or UO_3312 (O_3312,N_27767,N_27231);
and UO_3313 (O_3313,N_27293,N_28545);
or UO_3314 (O_3314,N_28148,N_27268);
nand UO_3315 (O_3315,N_29808,N_27197);
or UO_3316 (O_3316,N_28751,N_29054);
or UO_3317 (O_3317,N_28942,N_28481);
xnor UO_3318 (O_3318,N_29578,N_29444);
nor UO_3319 (O_3319,N_28844,N_28624);
xnor UO_3320 (O_3320,N_29654,N_27162);
nand UO_3321 (O_3321,N_29835,N_29053);
nand UO_3322 (O_3322,N_27726,N_28551);
nor UO_3323 (O_3323,N_29646,N_27887);
or UO_3324 (O_3324,N_29195,N_27764);
and UO_3325 (O_3325,N_29385,N_29768);
xnor UO_3326 (O_3326,N_28150,N_28569);
nor UO_3327 (O_3327,N_28901,N_29616);
nor UO_3328 (O_3328,N_28202,N_29744);
and UO_3329 (O_3329,N_29618,N_28495);
nor UO_3330 (O_3330,N_29291,N_27503);
or UO_3331 (O_3331,N_27017,N_29792);
xnor UO_3332 (O_3332,N_28367,N_28549);
nand UO_3333 (O_3333,N_27095,N_28478);
xnor UO_3334 (O_3334,N_28099,N_29985);
or UO_3335 (O_3335,N_28977,N_28630);
xor UO_3336 (O_3336,N_29449,N_27538);
or UO_3337 (O_3337,N_28473,N_27761);
nor UO_3338 (O_3338,N_27434,N_28471);
or UO_3339 (O_3339,N_28750,N_27036);
and UO_3340 (O_3340,N_28200,N_28849);
or UO_3341 (O_3341,N_28767,N_27468);
xnor UO_3342 (O_3342,N_28300,N_29889);
or UO_3343 (O_3343,N_28546,N_29044);
nand UO_3344 (O_3344,N_29012,N_29235);
nor UO_3345 (O_3345,N_29407,N_28544);
and UO_3346 (O_3346,N_27079,N_29019);
or UO_3347 (O_3347,N_27442,N_28855);
nand UO_3348 (O_3348,N_28338,N_28401);
and UO_3349 (O_3349,N_29644,N_29647);
xor UO_3350 (O_3350,N_27852,N_27581);
or UO_3351 (O_3351,N_28896,N_28346);
or UO_3352 (O_3352,N_29996,N_28477);
xnor UO_3353 (O_3353,N_27518,N_27173);
nor UO_3354 (O_3354,N_29717,N_29027);
nor UO_3355 (O_3355,N_28062,N_28185);
nor UO_3356 (O_3356,N_29925,N_28914);
xnor UO_3357 (O_3357,N_27186,N_29841);
and UO_3358 (O_3358,N_29570,N_28953);
nor UO_3359 (O_3359,N_29750,N_29009);
nor UO_3360 (O_3360,N_29157,N_29933);
nand UO_3361 (O_3361,N_27695,N_27495);
or UO_3362 (O_3362,N_27149,N_28538);
nor UO_3363 (O_3363,N_29856,N_27969);
xor UO_3364 (O_3364,N_28158,N_28859);
xor UO_3365 (O_3365,N_27662,N_28612);
nand UO_3366 (O_3366,N_29728,N_27761);
nor UO_3367 (O_3367,N_27988,N_27758);
or UO_3368 (O_3368,N_28656,N_29438);
or UO_3369 (O_3369,N_27308,N_27753);
and UO_3370 (O_3370,N_29871,N_29257);
nand UO_3371 (O_3371,N_27819,N_29936);
or UO_3372 (O_3372,N_27905,N_27241);
and UO_3373 (O_3373,N_28078,N_29802);
nand UO_3374 (O_3374,N_29449,N_28754);
nor UO_3375 (O_3375,N_28336,N_28103);
nor UO_3376 (O_3376,N_28094,N_27100);
xnor UO_3377 (O_3377,N_28347,N_29003);
and UO_3378 (O_3378,N_28583,N_29432);
nor UO_3379 (O_3379,N_29922,N_28495);
or UO_3380 (O_3380,N_27333,N_28201);
xor UO_3381 (O_3381,N_29340,N_29318);
or UO_3382 (O_3382,N_28467,N_28715);
nor UO_3383 (O_3383,N_27061,N_27480);
xnor UO_3384 (O_3384,N_27282,N_28061);
nor UO_3385 (O_3385,N_28725,N_27451);
nand UO_3386 (O_3386,N_27400,N_28261);
nor UO_3387 (O_3387,N_27249,N_29463);
nor UO_3388 (O_3388,N_29967,N_29880);
nand UO_3389 (O_3389,N_29636,N_29744);
nand UO_3390 (O_3390,N_27559,N_29530);
xor UO_3391 (O_3391,N_28650,N_28541);
or UO_3392 (O_3392,N_27594,N_27679);
xor UO_3393 (O_3393,N_28735,N_28762);
xnor UO_3394 (O_3394,N_29570,N_28110);
nand UO_3395 (O_3395,N_28276,N_27718);
xnor UO_3396 (O_3396,N_28771,N_28548);
nand UO_3397 (O_3397,N_29313,N_27951);
nor UO_3398 (O_3398,N_28408,N_28339);
nand UO_3399 (O_3399,N_29332,N_27959);
or UO_3400 (O_3400,N_29630,N_28179);
and UO_3401 (O_3401,N_27635,N_27163);
xnor UO_3402 (O_3402,N_28006,N_27809);
xnor UO_3403 (O_3403,N_28137,N_27711);
or UO_3404 (O_3404,N_29318,N_28899);
nor UO_3405 (O_3405,N_27182,N_29797);
xor UO_3406 (O_3406,N_28042,N_27988);
xor UO_3407 (O_3407,N_29181,N_29865);
or UO_3408 (O_3408,N_29025,N_29252);
nor UO_3409 (O_3409,N_27414,N_29447);
xnor UO_3410 (O_3410,N_29537,N_28115);
and UO_3411 (O_3411,N_27753,N_29469);
xor UO_3412 (O_3412,N_28027,N_28879);
nand UO_3413 (O_3413,N_28323,N_27205);
or UO_3414 (O_3414,N_29462,N_27785);
xor UO_3415 (O_3415,N_27376,N_28676);
or UO_3416 (O_3416,N_29934,N_28652);
nand UO_3417 (O_3417,N_27042,N_27376);
nor UO_3418 (O_3418,N_28078,N_27102);
nand UO_3419 (O_3419,N_27963,N_29707);
and UO_3420 (O_3420,N_29370,N_29143);
nand UO_3421 (O_3421,N_29286,N_28097);
xnor UO_3422 (O_3422,N_27450,N_27446);
nor UO_3423 (O_3423,N_28847,N_29993);
or UO_3424 (O_3424,N_28544,N_27577);
and UO_3425 (O_3425,N_28177,N_29575);
nand UO_3426 (O_3426,N_29764,N_28222);
xor UO_3427 (O_3427,N_28735,N_27792);
and UO_3428 (O_3428,N_29917,N_27384);
or UO_3429 (O_3429,N_29771,N_27472);
and UO_3430 (O_3430,N_27129,N_28166);
xnor UO_3431 (O_3431,N_29045,N_27909);
or UO_3432 (O_3432,N_28909,N_28228);
and UO_3433 (O_3433,N_29294,N_27370);
nand UO_3434 (O_3434,N_27815,N_29510);
nand UO_3435 (O_3435,N_29102,N_28720);
nand UO_3436 (O_3436,N_29038,N_29191);
xnor UO_3437 (O_3437,N_29833,N_28492);
nor UO_3438 (O_3438,N_29208,N_29777);
and UO_3439 (O_3439,N_28354,N_28707);
nor UO_3440 (O_3440,N_29661,N_28429);
nor UO_3441 (O_3441,N_28169,N_28350);
xor UO_3442 (O_3442,N_29658,N_28191);
nand UO_3443 (O_3443,N_29305,N_28418);
or UO_3444 (O_3444,N_29190,N_27843);
and UO_3445 (O_3445,N_29991,N_29291);
and UO_3446 (O_3446,N_29430,N_28514);
or UO_3447 (O_3447,N_28646,N_27687);
and UO_3448 (O_3448,N_29034,N_27636);
or UO_3449 (O_3449,N_29314,N_29590);
nand UO_3450 (O_3450,N_28246,N_28059);
or UO_3451 (O_3451,N_28386,N_29722);
nor UO_3452 (O_3452,N_28323,N_29678);
nor UO_3453 (O_3453,N_28252,N_27810);
and UO_3454 (O_3454,N_29886,N_28444);
xnor UO_3455 (O_3455,N_29121,N_29840);
xnor UO_3456 (O_3456,N_28393,N_27133);
nand UO_3457 (O_3457,N_28723,N_27877);
nor UO_3458 (O_3458,N_29524,N_29370);
and UO_3459 (O_3459,N_29803,N_29385);
or UO_3460 (O_3460,N_28117,N_28917);
and UO_3461 (O_3461,N_28273,N_27243);
xor UO_3462 (O_3462,N_28652,N_27492);
and UO_3463 (O_3463,N_29154,N_29386);
nand UO_3464 (O_3464,N_29556,N_29709);
or UO_3465 (O_3465,N_29558,N_28155);
nor UO_3466 (O_3466,N_28741,N_29026);
nor UO_3467 (O_3467,N_29634,N_28539);
or UO_3468 (O_3468,N_28740,N_29236);
nor UO_3469 (O_3469,N_28420,N_27047);
or UO_3470 (O_3470,N_29606,N_29384);
nand UO_3471 (O_3471,N_29465,N_29851);
or UO_3472 (O_3472,N_29961,N_28974);
nand UO_3473 (O_3473,N_28949,N_29373);
nand UO_3474 (O_3474,N_29587,N_29322);
xor UO_3475 (O_3475,N_29643,N_28262);
or UO_3476 (O_3476,N_27398,N_29663);
and UO_3477 (O_3477,N_29095,N_28388);
and UO_3478 (O_3478,N_29569,N_29333);
and UO_3479 (O_3479,N_29422,N_27276);
and UO_3480 (O_3480,N_28894,N_29773);
xnor UO_3481 (O_3481,N_29862,N_28803);
nand UO_3482 (O_3482,N_29756,N_28628);
or UO_3483 (O_3483,N_28144,N_29382);
and UO_3484 (O_3484,N_27334,N_29674);
or UO_3485 (O_3485,N_28800,N_28025);
nand UO_3486 (O_3486,N_27867,N_28175);
xor UO_3487 (O_3487,N_29532,N_28545);
and UO_3488 (O_3488,N_27332,N_28166);
nand UO_3489 (O_3489,N_27573,N_29305);
or UO_3490 (O_3490,N_29719,N_29311);
nand UO_3491 (O_3491,N_28858,N_27980);
and UO_3492 (O_3492,N_27941,N_29658);
nand UO_3493 (O_3493,N_28852,N_27809);
nand UO_3494 (O_3494,N_28092,N_29519);
nand UO_3495 (O_3495,N_29019,N_28572);
nand UO_3496 (O_3496,N_28025,N_28901);
xnor UO_3497 (O_3497,N_29872,N_27964);
and UO_3498 (O_3498,N_29033,N_27781);
or UO_3499 (O_3499,N_29673,N_27946);
endmodule