module basic_750_5000_1000_10_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_361,In_610);
nand U1 (N_1,In_379,In_50);
nor U2 (N_2,In_400,In_736);
or U3 (N_3,In_67,In_539);
nand U4 (N_4,In_307,In_121);
or U5 (N_5,In_576,In_578);
nand U6 (N_6,In_306,In_150);
and U7 (N_7,In_603,In_586);
nand U8 (N_8,In_556,In_739);
or U9 (N_9,In_631,In_674);
xnor U10 (N_10,In_165,In_697);
nand U11 (N_11,In_221,In_503);
nand U12 (N_12,In_429,In_547);
nor U13 (N_13,In_508,In_483);
or U14 (N_14,In_482,In_83);
and U15 (N_15,In_567,In_319);
nor U16 (N_16,In_220,In_284);
nor U17 (N_17,In_575,In_635);
and U18 (N_18,In_722,In_551);
nor U19 (N_19,In_640,In_623);
nand U20 (N_20,In_649,In_634);
nor U21 (N_21,In_600,In_721);
nor U22 (N_22,In_471,In_500);
or U23 (N_23,In_713,In_66);
nor U24 (N_24,In_177,In_317);
nand U25 (N_25,In_84,In_313);
nor U26 (N_26,In_678,In_373);
or U27 (N_27,In_422,In_468);
nand U28 (N_28,In_132,In_691);
xnor U29 (N_29,In_144,In_704);
nor U30 (N_30,In_253,In_134);
or U31 (N_31,In_733,In_271);
and U32 (N_32,In_597,In_224);
and U33 (N_33,In_385,In_671);
and U34 (N_34,In_367,In_16);
or U35 (N_35,In_316,In_241);
and U36 (N_36,In_4,In_44);
nand U37 (N_37,In_608,In_176);
nand U38 (N_38,In_676,In_708);
nor U39 (N_39,In_356,In_267);
or U40 (N_40,In_215,In_131);
nor U41 (N_41,In_302,In_737);
xor U42 (N_42,In_238,In_626);
and U43 (N_43,In_726,In_265);
nand U44 (N_44,In_375,In_596);
and U45 (N_45,In_485,In_652);
nor U46 (N_46,In_469,In_701);
or U47 (N_47,In_178,In_130);
and U48 (N_48,In_390,In_218);
or U49 (N_49,In_728,In_607);
nand U50 (N_50,In_531,In_74);
nor U51 (N_51,In_527,In_6);
and U52 (N_52,In_703,In_278);
or U53 (N_53,In_425,In_181);
nor U54 (N_54,In_263,In_655);
or U55 (N_55,In_28,In_374);
nand U56 (N_56,In_112,In_211);
and U57 (N_57,In_170,In_333);
or U58 (N_58,In_89,In_258);
and U59 (N_59,In_413,In_219);
and U60 (N_60,In_583,In_23);
nand U61 (N_61,In_202,In_561);
or U62 (N_62,In_227,In_738);
or U63 (N_63,In_366,In_504);
or U64 (N_64,In_168,In_473);
nand U65 (N_65,In_376,In_746);
nor U66 (N_66,In_614,In_183);
and U67 (N_67,In_300,In_298);
nand U68 (N_68,In_90,In_53);
nor U69 (N_69,In_257,In_731);
nor U70 (N_70,In_457,In_548);
nand U71 (N_71,In_214,In_229);
or U72 (N_72,In_477,In_45);
nand U73 (N_73,In_236,In_580);
nand U74 (N_74,In_166,In_314);
or U75 (N_75,In_564,In_507);
and U76 (N_76,In_543,In_346);
or U77 (N_77,In_452,In_495);
and U78 (N_78,In_46,In_673);
nand U79 (N_79,In_677,In_106);
or U80 (N_80,In_282,In_71);
nand U81 (N_81,In_514,In_117);
and U82 (N_82,In_136,In_435);
nand U83 (N_83,In_291,In_418);
and U84 (N_84,In_541,In_643);
nor U85 (N_85,In_518,In_647);
nor U86 (N_86,In_570,In_480);
and U87 (N_87,In_235,In_466);
nand U88 (N_88,In_217,In_743);
and U89 (N_89,In_563,In_365);
nor U90 (N_90,In_138,In_421);
or U91 (N_91,In_506,In_711);
and U92 (N_92,In_154,In_99);
nand U93 (N_93,In_330,In_740);
nand U94 (N_94,In_472,In_720);
or U95 (N_95,In_207,In_644);
nand U96 (N_96,In_85,In_206);
nand U97 (N_97,In_140,In_172);
nor U98 (N_98,In_328,In_591);
or U99 (N_99,In_351,In_593);
nor U100 (N_100,In_275,In_515);
or U101 (N_101,In_695,In_279);
or U102 (N_102,In_599,In_137);
nor U103 (N_103,In_656,In_540);
nand U104 (N_104,In_357,In_742);
nor U105 (N_105,In_456,In_297);
and U106 (N_106,In_645,In_148);
or U107 (N_107,In_288,In_700);
or U108 (N_108,In_398,In_173);
or U109 (N_109,In_588,In_244);
nor U110 (N_110,In_404,In_308);
nand U111 (N_111,In_353,In_286);
or U112 (N_112,In_110,In_533);
nor U113 (N_113,In_433,In_345);
nand U114 (N_114,In_526,In_702);
nor U115 (N_115,In_149,In_577);
or U116 (N_116,In_231,In_684);
nor U117 (N_117,In_143,In_546);
nor U118 (N_118,In_553,In_57);
or U119 (N_119,In_301,In_524);
nand U120 (N_120,In_403,In_430);
nand U121 (N_121,In_416,In_560);
or U122 (N_122,In_159,In_399);
or U123 (N_123,In_100,In_324);
and U124 (N_124,In_9,In_748);
and U125 (N_125,In_281,In_64);
and U126 (N_126,In_14,In_654);
and U127 (N_127,In_549,In_715);
or U128 (N_128,In_488,In_40);
nand U129 (N_129,In_190,In_228);
nor U130 (N_130,In_26,In_212);
nor U131 (N_131,In_20,In_545);
nor U132 (N_132,In_182,In_675);
nor U133 (N_133,In_186,In_126);
nand U134 (N_134,In_692,In_283);
nor U135 (N_135,In_29,In_646);
nor U136 (N_136,In_24,In_419);
nand U137 (N_137,In_34,In_261);
or U138 (N_138,In_156,In_426);
nor U139 (N_139,In_123,In_157);
nor U140 (N_140,In_188,In_368);
or U141 (N_141,In_396,In_120);
or U142 (N_142,In_58,In_359);
nand U143 (N_143,In_683,In_25);
or U144 (N_144,In_641,In_438);
or U145 (N_145,In_402,In_441);
nor U146 (N_146,In_522,In_461);
nor U147 (N_147,In_557,In_254);
nor U148 (N_148,In_354,In_584);
or U149 (N_149,In_442,In_609);
or U150 (N_150,In_509,In_242);
or U151 (N_151,In_377,In_363);
or U152 (N_152,In_344,In_450);
nand U153 (N_153,In_295,In_334);
and U154 (N_154,In_668,In_5);
nor U155 (N_155,In_108,In_434);
or U156 (N_156,In_222,In_554);
and U157 (N_157,In_699,In_658);
nor U158 (N_158,In_75,In_371);
nand U159 (N_159,In_667,In_88);
nand U160 (N_160,In_664,In_70);
or U161 (N_161,In_341,In_252);
nand U162 (N_162,In_325,In_338);
nor U163 (N_163,In_0,In_378);
and U164 (N_164,In_417,In_660);
nor U165 (N_165,In_620,In_209);
and U166 (N_166,In_230,In_535);
nor U167 (N_167,In_447,In_428);
and U168 (N_168,In_439,In_36);
and U169 (N_169,In_93,In_725);
nor U170 (N_170,In_550,In_519);
nor U171 (N_171,In_414,In_744);
nand U172 (N_172,In_76,In_536);
and U173 (N_173,In_653,In_666);
and U174 (N_174,In_719,In_613);
and U175 (N_175,In_95,In_362);
or U176 (N_176,In_216,In_462);
nand U177 (N_177,In_54,In_332);
or U178 (N_178,In_256,In_160);
nand U179 (N_179,In_255,In_39);
nor U180 (N_180,In_129,In_384);
nor U181 (N_181,In_494,In_262);
or U182 (N_182,In_496,In_331);
or U183 (N_183,In_512,In_77);
or U184 (N_184,In_349,In_705);
nand U185 (N_185,In_124,In_397);
and U186 (N_186,In_627,In_718);
nand U187 (N_187,In_21,In_393);
or U188 (N_188,In_625,In_147);
or U189 (N_189,In_27,In_478);
nand U190 (N_190,In_350,In_501);
nand U191 (N_191,In_3,In_490);
nor U192 (N_192,In_35,In_723);
and U193 (N_193,In_10,In_246);
or U194 (N_194,In_248,In_56);
nor U195 (N_195,In_343,In_17);
or U196 (N_196,In_693,In_611);
and U197 (N_197,In_115,In_169);
nor U198 (N_198,In_141,In_22);
nand U199 (N_199,In_250,In_61);
nand U200 (N_200,In_432,In_714);
nor U201 (N_201,In_203,In_293);
nor U202 (N_202,In_266,In_259);
nand U203 (N_203,In_101,In_197);
and U204 (N_204,In_49,In_572);
and U205 (N_205,In_237,In_318);
or U206 (N_206,In_559,In_630);
nor U207 (N_207,In_582,In_194);
nor U208 (N_208,In_642,In_240);
nand U209 (N_209,In_735,In_410);
and U210 (N_210,In_423,In_37);
nand U211 (N_211,In_493,In_19);
nor U212 (N_212,In_612,In_663);
nand U213 (N_213,In_679,In_405);
and U214 (N_214,In_680,In_712);
or U215 (N_215,In_304,In_72);
and U216 (N_216,In_339,In_2);
nor U217 (N_217,In_201,In_386);
nor U218 (N_218,In_690,In_96);
or U219 (N_219,In_624,In_322);
nor U220 (N_220,In_463,In_638);
nand U221 (N_221,In_47,In_369);
and U222 (N_222,In_285,In_498);
or U223 (N_223,In_622,In_619);
nand U224 (N_224,In_392,In_401);
or U225 (N_225,In_688,In_65);
or U226 (N_226,In_724,In_534);
nand U227 (N_227,In_274,In_30);
nor U228 (N_228,In_568,In_710);
and U229 (N_229,In_81,In_370);
nor U230 (N_230,In_280,In_233);
nand U231 (N_231,In_628,In_445);
and U232 (N_232,In_552,In_62);
nand U233 (N_233,In_200,In_618);
or U234 (N_234,In_602,In_208);
and U235 (N_235,In_133,In_198);
nand U236 (N_236,In_292,In_538);
or U237 (N_237,In_505,In_270);
nand U238 (N_238,In_303,In_287);
nor U239 (N_239,In_449,In_145);
or U240 (N_240,In_155,In_581);
or U241 (N_241,In_364,In_745);
and U242 (N_242,In_69,In_55);
nand U243 (N_243,In_199,In_78);
nand U244 (N_244,In_311,In_520);
and U245 (N_245,In_565,In_48);
and U246 (N_246,In_380,In_305);
nand U247 (N_247,In_162,In_113);
and U248 (N_248,In_558,In_193);
or U249 (N_249,In_440,In_273);
nor U250 (N_250,In_91,In_342);
nor U251 (N_251,In_87,In_479);
nand U252 (N_252,In_569,In_590);
and U253 (N_253,In_243,In_670);
or U254 (N_254,In_521,In_355);
and U255 (N_255,In_406,In_427);
nor U256 (N_256,In_80,In_436);
nor U257 (N_257,In_294,In_92);
and U258 (N_258,In_180,In_164);
and U259 (N_259,In_73,In_689);
nand U260 (N_260,In_458,In_51);
and U261 (N_261,In_326,In_621);
and U262 (N_262,In_467,In_204);
nand U263 (N_263,In_484,In_446);
nand U264 (N_264,In_142,In_276);
or U265 (N_265,In_451,In_650);
nor U266 (N_266,In_223,In_530);
nor U267 (N_267,In_38,In_727);
or U268 (N_268,In_104,In_8);
and U269 (N_269,In_226,In_329);
and U270 (N_270,In_443,In_573);
and U271 (N_271,In_210,In_272);
nor U272 (N_272,In_470,In_102);
and U273 (N_273,In_682,In_158);
and U274 (N_274,In_383,In_174);
nor U275 (N_275,In_225,In_487);
or U276 (N_276,In_408,In_18);
and U277 (N_277,In_167,In_592);
nor U278 (N_278,In_135,In_388);
nand U279 (N_279,In_98,In_732);
and U280 (N_280,In_323,In_213);
nor U281 (N_281,In_391,In_335);
nand U282 (N_282,In_289,In_605);
or U283 (N_283,In_179,In_601);
and U284 (N_284,In_681,In_617);
and U285 (N_285,In_662,In_659);
nand U286 (N_286,In_33,In_239);
or U287 (N_287,In_606,In_492);
and U288 (N_288,In_1,In_562);
nand U289 (N_289,In_517,In_694);
nand U290 (N_290,In_555,In_516);
or U291 (N_291,In_125,In_513);
and U292 (N_292,In_730,In_296);
and U293 (N_293,In_109,In_107);
and U294 (N_294,In_615,In_598);
and U295 (N_295,In_310,In_94);
and U296 (N_296,In_249,In_637);
nor U297 (N_297,In_389,In_629);
or U298 (N_298,In_12,In_502);
nor U299 (N_299,In_707,In_340);
nor U300 (N_300,In_86,In_232);
or U301 (N_301,In_41,In_116);
or U302 (N_302,In_585,In_415);
or U303 (N_303,In_525,In_636);
and U304 (N_304,In_32,In_337);
and U305 (N_305,In_717,In_63);
nand U306 (N_306,In_7,In_234);
and U307 (N_307,In_651,In_151);
nor U308 (N_308,In_595,In_729);
nand U309 (N_309,In_734,In_184);
nor U310 (N_310,In_542,In_163);
xnor U311 (N_311,In_459,In_139);
nand U312 (N_312,In_544,In_128);
or U313 (N_313,In_444,In_747);
and U314 (N_314,In_594,In_52);
xor U315 (N_315,In_103,In_79);
or U316 (N_316,In_269,In_476);
nor U317 (N_317,In_336,In_187);
nor U318 (N_318,In_464,In_195);
or U319 (N_319,In_465,In_453);
or U320 (N_320,In_60,In_486);
nand U321 (N_321,In_382,In_616);
and U322 (N_322,In_604,In_437);
or U323 (N_323,In_706,In_327);
or U324 (N_324,In_528,In_481);
nand U325 (N_325,In_523,In_15);
nand U326 (N_326,In_491,In_245);
nor U327 (N_327,In_11,In_455);
nor U328 (N_328,In_264,In_431);
or U329 (N_329,In_589,In_566);
nor U330 (N_330,In_474,In_320);
nor U331 (N_331,In_686,In_122);
or U332 (N_332,In_161,In_97);
and U333 (N_333,In_68,In_510);
nor U334 (N_334,In_309,In_146);
nand U335 (N_335,In_687,In_315);
nand U336 (N_336,In_290,In_268);
and U337 (N_337,In_13,In_412);
nor U338 (N_338,In_716,In_387);
and U339 (N_339,In_685,In_118);
nand U340 (N_340,In_537,In_669);
and U341 (N_341,In_372,In_111);
or U342 (N_342,In_454,In_277);
or U343 (N_343,In_119,In_511);
and U344 (N_344,In_657,In_352);
nand U345 (N_345,In_185,In_191);
nor U346 (N_346,In_394,In_82);
and U347 (N_347,In_312,In_105);
and U348 (N_348,In_571,In_696);
nor U349 (N_349,In_672,In_152);
or U350 (N_350,In_632,In_665);
or U351 (N_351,In_59,In_205);
nand U352 (N_352,In_499,In_648);
or U353 (N_353,In_407,In_42);
and U354 (N_354,In_395,In_171);
or U355 (N_355,In_411,In_358);
and U356 (N_356,In_360,In_574);
nor U357 (N_357,In_192,In_639);
or U358 (N_358,In_497,In_175);
nor U359 (N_359,In_424,In_196);
and U360 (N_360,In_460,In_381);
and U361 (N_361,In_127,In_348);
nand U362 (N_362,In_749,In_189);
nor U363 (N_363,In_31,In_448);
and U364 (N_364,In_532,In_587);
and U365 (N_365,In_633,In_409);
nor U366 (N_366,In_489,In_709);
and U367 (N_367,In_698,In_153);
and U368 (N_368,In_43,In_114);
nand U369 (N_369,In_475,In_741);
nand U370 (N_370,In_661,In_420);
or U371 (N_371,In_347,In_251);
nor U372 (N_372,In_260,In_247);
nand U373 (N_373,In_299,In_321);
nor U374 (N_374,In_579,In_529);
nand U375 (N_375,In_468,In_391);
and U376 (N_376,In_574,In_536);
nor U377 (N_377,In_576,In_748);
nor U378 (N_378,In_731,In_207);
nand U379 (N_379,In_73,In_127);
nand U380 (N_380,In_111,In_254);
and U381 (N_381,In_390,In_432);
nor U382 (N_382,In_449,In_730);
nor U383 (N_383,In_550,In_208);
nor U384 (N_384,In_371,In_334);
nor U385 (N_385,In_94,In_704);
and U386 (N_386,In_393,In_53);
or U387 (N_387,In_576,In_176);
nor U388 (N_388,In_592,In_622);
nor U389 (N_389,In_405,In_65);
xor U390 (N_390,In_311,In_273);
or U391 (N_391,In_517,In_194);
or U392 (N_392,In_7,In_553);
or U393 (N_393,In_464,In_140);
or U394 (N_394,In_350,In_579);
nand U395 (N_395,In_610,In_285);
nand U396 (N_396,In_17,In_279);
nand U397 (N_397,In_645,In_483);
nor U398 (N_398,In_533,In_176);
and U399 (N_399,In_44,In_572);
nand U400 (N_400,In_372,In_327);
nor U401 (N_401,In_442,In_538);
nand U402 (N_402,In_416,In_332);
nand U403 (N_403,In_364,In_225);
or U404 (N_404,In_731,In_728);
and U405 (N_405,In_500,In_381);
nor U406 (N_406,In_220,In_447);
and U407 (N_407,In_550,In_359);
and U408 (N_408,In_29,In_117);
nand U409 (N_409,In_41,In_322);
or U410 (N_410,In_587,In_739);
nor U411 (N_411,In_238,In_460);
nor U412 (N_412,In_222,In_304);
and U413 (N_413,In_328,In_442);
and U414 (N_414,In_62,In_45);
or U415 (N_415,In_425,In_449);
nand U416 (N_416,In_330,In_607);
or U417 (N_417,In_640,In_70);
and U418 (N_418,In_182,In_410);
and U419 (N_419,In_519,In_736);
nor U420 (N_420,In_622,In_236);
and U421 (N_421,In_431,In_546);
nand U422 (N_422,In_137,In_248);
nand U423 (N_423,In_736,In_417);
or U424 (N_424,In_746,In_679);
nand U425 (N_425,In_233,In_688);
and U426 (N_426,In_595,In_714);
or U427 (N_427,In_598,In_353);
nand U428 (N_428,In_697,In_375);
or U429 (N_429,In_121,In_478);
and U430 (N_430,In_165,In_535);
or U431 (N_431,In_652,In_217);
and U432 (N_432,In_186,In_541);
nand U433 (N_433,In_7,In_730);
or U434 (N_434,In_289,In_338);
and U435 (N_435,In_323,In_285);
and U436 (N_436,In_431,In_223);
xor U437 (N_437,In_499,In_449);
or U438 (N_438,In_150,In_477);
nand U439 (N_439,In_223,In_597);
or U440 (N_440,In_504,In_632);
or U441 (N_441,In_99,In_740);
nor U442 (N_442,In_134,In_562);
nand U443 (N_443,In_496,In_59);
nand U444 (N_444,In_184,In_395);
or U445 (N_445,In_727,In_55);
nor U446 (N_446,In_295,In_78);
nor U447 (N_447,In_222,In_458);
and U448 (N_448,In_287,In_657);
and U449 (N_449,In_610,In_86);
and U450 (N_450,In_614,In_702);
nor U451 (N_451,In_728,In_50);
nor U452 (N_452,In_122,In_411);
and U453 (N_453,In_276,In_698);
and U454 (N_454,In_748,In_345);
nand U455 (N_455,In_537,In_720);
or U456 (N_456,In_407,In_121);
nor U457 (N_457,In_344,In_297);
or U458 (N_458,In_618,In_412);
and U459 (N_459,In_84,In_631);
and U460 (N_460,In_189,In_512);
nor U461 (N_461,In_567,In_260);
and U462 (N_462,In_698,In_668);
nand U463 (N_463,In_299,In_439);
nor U464 (N_464,In_548,In_130);
and U465 (N_465,In_745,In_730);
nor U466 (N_466,In_350,In_609);
and U467 (N_467,In_179,In_131);
and U468 (N_468,In_674,In_642);
and U469 (N_469,In_255,In_61);
nand U470 (N_470,In_715,In_358);
nor U471 (N_471,In_635,In_489);
nand U472 (N_472,In_590,In_190);
nand U473 (N_473,In_66,In_315);
nand U474 (N_474,In_173,In_77);
and U475 (N_475,In_597,In_723);
nor U476 (N_476,In_578,In_31);
and U477 (N_477,In_170,In_23);
or U478 (N_478,In_209,In_172);
nand U479 (N_479,In_22,In_284);
or U480 (N_480,In_729,In_379);
nor U481 (N_481,In_255,In_710);
nand U482 (N_482,In_163,In_0);
or U483 (N_483,In_431,In_608);
and U484 (N_484,In_255,In_321);
nand U485 (N_485,In_547,In_202);
or U486 (N_486,In_35,In_336);
and U487 (N_487,In_479,In_311);
and U488 (N_488,In_612,In_734);
nor U489 (N_489,In_559,In_93);
and U490 (N_490,In_742,In_220);
nor U491 (N_491,In_140,In_688);
nand U492 (N_492,In_49,In_174);
xnor U493 (N_493,In_49,In_460);
or U494 (N_494,In_632,In_75);
nand U495 (N_495,In_335,In_413);
or U496 (N_496,In_63,In_88);
and U497 (N_497,In_94,In_358);
or U498 (N_498,In_505,In_705);
nor U499 (N_499,In_672,In_196);
and U500 (N_500,N_250,N_488);
nand U501 (N_501,N_152,N_138);
or U502 (N_502,N_66,N_102);
nand U503 (N_503,N_233,N_348);
or U504 (N_504,N_90,N_175);
nor U505 (N_505,N_195,N_338);
nor U506 (N_506,N_265,N_232);
nand U507 (N_507,N_38,N_472);
nand U508 (N_508,N_154,N_81);
and U509 (N_509,N_398,N_179);
and U510 (N_510,N_103,N_475);
nand U511 (N_511,N_401,N_225);
nor U512 (N_512,N_322,N_26);
nor U513 (N_513,N_471,N_67);
or U514 (N_514,N_463,N_56);
nand U515 (N_515,N_220,N_5);
nand U516 (N_516,N_367,N_288);
and U517 (N_517,N_424,N_198);
nor U518 (N_518,N_385,N_492);
nor U519 (N_519,N_221,N_335);
nor U520 (N_520,N_235,N_380);
or U521 (N_521,N_376,N_130);
nand U522 (N_522,N_342,N_439);
nor U523 (N_523,N_469,N_302);
nand U524 (N_524,N_321,N_363);
nor U525 (N_525,N_153,N_479);
nor U526 (N_526,N_337,N_381);
nor U527 (N_527,N_149,N_453);
and U528 (N_528,N_304,N_169);
nor U529 (N_529,N_7,N_356);
nand U530 (N_530,N_25,N_310);
nor U531 (N_531,N_364,N_467);
and U532 (N_532,N_125,N_78);
nand U533 (N_533,N_285,N_20);
nor U534 (N_534,N_243,N_206);
or U535 (N_535,N_89,N_464);
nor U536 (N_536,N_332,N_327);
xnor U537 (N_537,N_57,N_480);
nand U538 (N_538,N_408,N_256);
and U539 (N_539,N_186,N_438);
and U540 (N_540,N_201,N_156);
and U541 (N_541,N_474,N_294);
or U542 (N_542,N_457,N_24);
nand U543 (N_543,N_121,N_300);
nor U544 (N_544,N_183,N_390);
nand U545 (N_545,N_62,N_460);
nand U546 (N_546,N_443,N_495);
nand U547 (N_547,N_194,N_426);
nor U548 (N_548,N_404,N_270);
and U549 (N_549,N_173,N_362);
nand U550 (N_550,N_284,N_448);
or U551 (N_551,N_258,N_54);
nand U552 (N_552,N_461,N_218);
nand U553 (N_553,N_478,N_98);
or U554 (N_554,N_122,N_187);
nand U555 (N_555,N_455,N_127);
and U556 (N_556,N_303,N_217);
or U557 (N_557,N_423,N_454);
and U558 (N_558,N_1,N_373);
nand U559 (N_559,N_85,N_83);
nor U560 (N_560,N_482,N_42);
nand U561 (N_561,N_437,N_386);
and U562 (N_562,N_309,N_55);
or U563 (N_563,N_339,N_357);
nand U564 (N_564,N_485,N_352);
and U565 (N_565,N_99,N_417);
or U566 (N_566,N_176,N_29);
or U567 (N_567,N_476,N_170);
nand U568 (N_568,N_188,N_43);
or U569 (N_569,N_136,N_290);
or U570 (N_570,N_389,N_456);
nor U571 (N_571,N_378,N_383);
and U572 (N_572,N_49,N_76);
and U573 (N_573,N_94,N_244);
and U574 (N_574,N_189,N_286);
nor U575 (N_575,N_126,N_14);
and U576 (N_576,N_402,N_248);
nor U577 (N_577,N_222,N_172);
or U578 (N_578,N_349,N_145);
or U579 (N_579,N_280,N_28);
and U580 (N_580,N_208,N_272);
nand U581 (N_581,N_277,N_110);
and U582 (N_582,N_370,N_45);
or U583 (N_583,N_462,N_161);
and U584 (N_584,N_41,N_4);
or U585 (N_585,N_268,N_331);
and U586 (N_586,N_224,N_27);
nand U587 (N_587,N_433,N_157);
nand U588 (N_588,N_400,N_92);
nor U589 (N_589,N_190,N_366);
or U590 (N_590,N_163,N_255);
and U591 (N_591,N_200,N_320);
or U592 (N_592,N_343,N_46);
nand U593 (N_593,N_174,N_204);
nand U594 (N_594,N_128,N_344);
or U595 (N_595,N_360,N_414);
or U596 (N_596,N_409,N_80);
and U597 (N_597,N_82,N_63);
nor U598 (N_598,N_18,N_296);
or U599 (N_599,N_253,N_61);
and U600 (N_600,N_249,N_245);
or U601 (N_601,N_184,N_91);
nor U602 (N_602,N_452,N_51);
nor U603 (N_603,N_237,N_15);
nor U604 (N_604,N_240,N_498);
nor U605 (N_605,N_295,N_421);
or U606 (N_606,N_199,N_297);
nor U607 (N_607,N_271,N_40);
nor U608 (N_608,N_52,N_114);
and U609 (N_609,N_289,N_35);
or U610 (N_610,N_75,N_151);
nand U611 (N_611,N_22,N_434);
or U612 (N_612,N_496,N_59);
or U613 (N_613,N_316,N_493);
nand U614 (N_614,N_266,N_345);
or U615 (N_615,N_65,N_403);
nand U616 (N_616,N_451,N_226);
or U617 (N_617,N_330,N_312);
nand U618 (N_618,N_158,N_311);
nor U619 (N_619,N_430,N_168);
nor U620 (N_620,N_251,N_229);
or U621 (N_621,N_359,N_139);
or U622 (N_622,N_325,N_422);
nor U623 (N_623,N_10,N_328);
nand U624 (N_624,N_64,N_77);
nand U625 (N_625,N_193,N_132);
or U626 (N_626,N_387,N_148);
and U627 (N_627,N_301,N_72);
nor U628 (N_628,N_0,N_178);
or U629 (N_629,N_375,N_3);
or U630 (N_630,N_101,N_410);
nand U631 (N_631,N_407,N_420);
nand U632 (N_632,N_6,N_274);
and U633 (N_633,N_137,N_267);
nor U634 (N_634,N_13,N_155);
nand U635 (N_635,N_413,N_384);
or U636 (N_636,N_71,N_371);
and U637 (N_637,N_2,N_405);
nand U638 (N_638,N_459,N_432);
nor U639 (N_639,N_435,N_227);
or U640 (N_640,N_326,N_143);
nand U641 (N_641,N_37,N_254);
nor U642 (N_642,N_395,N_213);
nor U643 (N_643,N_68,N_269);
and U644 (N_644,N_305,N_202);
nor U645 (N_645,N_53,N_263);
or U646 (N_646,N_281,N_334);
nand U647 (N_647,N_483,N_234);
and U648 (N_648,N_48,N_203);
and U649 (N_649,N_23,N_87);
or U650 (N_650,N_315,N_9);
nand U651 (N_651,N_215,N_358);
nand U652 (N_652,N_298,N_147);
or U653 (N_653,N_212,N_411);
and U654 (N_654,N_445,N_353);
and U655 (N_655,N_441,N_428);
nor U656 (N_656,N_129,N_144);
or U657 (N_657,N_210,N_30);
nor U658 (N_658,N_238,N_11);
or U659 (N_659,N_34,N_484);
nand U660 (N_660,N_107,N_416);
or U661 (N_661,N_242,N_278);
nand U662 (N_662,N_12,N_499);
nand U663 (N_663,N_39,N_473);
nor U664 (N_664,N_50,N_429);
nand U665 (N_665,N_140,N_350);
nor U666 (N_666,N_230,N_207);
or U667 (N_667,N_167,N_96);
nand U668 (N_668,N_180,N_355);
nor U669 (N_669,N_197,N_425);
nor U670 (N_670,N_69,N_160);
or U671 (N_671,N_369,N_368);
nand U672 (N_672,N_260,N_372);
and U673 (N_673,N_282,N_489);
or U674 (N_674,N_406,N_181);
and U675 (N_675,N_351,N_391);
and U676 (N_676,N_177,N_146);
nor U677 (N_677,N_216,N_123);
nand U678 (N_678,N_182,N_468);
and U679 (N_679,N_135,N_314);
and U680 (N_680,N_159,N_196);
nand U681 (N_681,N_340,N_134);
or U682 (N_682,N_436,N_276);
or U683 (N_683,N_259,N_447);
nor U684 (N_684,N_214,N_185);
and U685 (N_685,N_336,N_393);
and U686 (N_686,N_112,N_150);
or U687 (N_687,N_47,N_33);
nor U688 (N_688,N_487,N_211);
nor U689 (N_689,N_490,N_32);
nor U690 (N_690,N_279,N_88);
or U691 (N_691,N_494,N_74);
or U692 (N_692,N_466,N_19);
nand U693 (N_693,N_418,N_419);
or U694 (N_694,N_109,N_394);
and U695 (N_695,N_446,N_392);
and U696 (N_696,N_219,N_449);
or U697 (N_697,N_317,N_162);
nand U698 (N_698,N_283,N_70);
nand U699 (N_699,N_442,N_396);
nand U700 (N_700,N_105,N_341);
nor U701 (N_701,N_165,N_131);
and U702 (N_702,N_313,N_236);
nand U703 (N_703,N_307,N_486);
and U704 (N_704,N_329,N_497);
xor U705 (N_705,N_113,N_458);
or U706 (N_706,N_79,N_95);
and U707 (N_707,N_333,N_354);
and U708 (N_708,N_246,N_318);
or U709 (N_709,N_21,N_142);
or U710 (N_710,N_308,N_36);
nor U711 (N_711,N_306,N_261);
or U712 (N_712,N_465,N_324);
nand U713 (N_713,N_481,N_231);
and U714 (N_714,N_264,N_120);
nor U715 (N_715,N_293,N_273);
or U716 (N_716,N_397,N_477);
nand U717 (N_717,N_319,N_205);
or U718 (N_718,N_262,N_427);
and U719 (N_719,N_415,N_450);
and U720 (N_720,N_239,N_124);
and U721 (N_721,N_111,N_44);
nor U722 (N_722,N_60,N_379);
nor U723 (N_723,N_440,N_93);
nor U724 (N_724,N_491,N_133);
nand U725 (N_725,N_118,N_431);
or U726 (N_726,N_257,N_164);
nor U727 (N_727,N_104,N_58);
or U728 (N_728,N_377,N_16);
and U729 (N_729,N_106,N_275);
or U730 (N_730,N_287,N_86);
and U731 (N_731,N_73,N_100);
and U732 (N_732,N_8,N_141);
nand U733 (N_733,N_346,N_374);
or U734 (N_734,N_171,N_119);
nor U735 (N_735,N_192,N_191);
or U736 (N_736,N_323,N_228);
and U737 (N_737,N_241,N_247);
or U738 (N_738,N_108,N_299);
and U739 (N_739,N_291,N_382);
and U740 (N_740,N_412,N_31);
and U741 (N_741,N_17,N_166);
and U742 (N_742,N_223,N_116);
or U743 (N_743,N_209,N_444);
nor U744 (N_744,N_117,N_347);
nor U745 (N_745,N_399,N_97);
nor U746 (N_746,N_292,N_115);
and U747 (N_747,N_470,N_365);
nor U748 (N_748,N_84,N_388);
nand U749 (N_749,N_252,N_361);
xor U750 (N_750,N_189,N_14);
nand U751 (N_751,N_1,N_174);
and U752 (N_752,N_265,N_321);
nand U753 (N_753,N_487,N_152);
and U754 (N_754,N_449,N_479);
or U755 (N_755,N_38,N_239);
or U756 (N_756,N_299,N_305);
or U757 (N_757,N_32,N_161);
or U758 (N_758,N_91,N_295);
nand U759 (N_759,N_452,N_50);
nand U760 (N_760,N_321,N_94);
nand U761 (N_761,N_9,N_17);
nor U762 (N_762,N_361,N_327);
nor U763 (N_763,N_242,N_452);
or U764 (N_764,N_362,N_415);
xor U765 (N_765,N_155,N_352);
and U766 (N_766,N_226,N_462);
and U767 (N_767,N_112,N_443);
nand U768 (N_768,N_290,N_424);
or U769 (N_769,N_129,N_375);
nand U770 (N_770,N_430,N_458);
nor U771 (N_771,N_337,N_328);
nor U772 (N_772,N_443,N_130);
or U773 (N_773,N_153,N_299);
nand U774 (N_774,N_162,N_208);
or U775 (N_775,N_304,N_356);
nand U776 (N_776,N_82,N_289);
nand U777 (N_777,N_376,N_475);
or U778 (N_778,N_241,N_176);
nand U779 (N_779,N_482,N_6);
nor U780 (N_780,N_472,N_112);
nand U781 (N_781,N_101,N_49);
nor U782 (N_782,N_421,N_481);
nor U783 (N_783,N_126,N_428);
nand U784 (N_784,N_222,N_270);
and U785 (N_785,N_157,N_337);
nor U786 (N_786,N_445,N_105);
or U787 (N_787,N_433,N_234);
nand U788 (N_788,N_294,N_103);
nor U789 (N_789,N_125,N_395);
nor U790 (N_790,N_475,N_28);
nand U791 (N_791,N_160,N_344);
nor U792 (N_792,N_263,N_397);
and U793 (N_793,N_493,N_442);
nor U794 (N_794,N_278,N_268);
and U795 (N_795,N_438,N_485);
or U796 (N_796,N_312,N_299);
nand U797 (N_797,N_19,N_34);
or U798 (N_798,N_264,N_66);
nand U799 (N_799,N_17,N_398);
nand U800 (N_800,N_239,N_322);
or U801 (N_801,N_319,N_0);
nand U802 (N_802,N_114,N_26);
or U803 (N_803,N_417,N_64);
nand U804 (N_804,N_285,N_119);
nor U805 (N_805,N_229,N_427);
nand U806 (N_806,N_341,N_339);
nor U807 (N_807,N_352,N_268);
nor U808 (N_808,N_250,N_433);
nor U809 (N_809,N_111,N_272);
and U810 (N_810,N_89,N_47);
and U811 (N_811,N_240,N_435);
nand U812 (N_812,N_499,N_236);
or U813 (N_813,N_260,N_312);
or U814 (N_814,N_204,N_439);
nand U815 (N_815,N_353,N_115);
and U816 (N_816,N_176,N_193);
and U817 (N_817,N_465,N_442);
nand U818 (N_818,N_213,N_437);
nand U819 (N_819,N_411,N_117);
nor U820 (N_820,N_372,N_116);
nand U821 (N_821,N_250,N_287);
and U822 (N_822,N_368,N_304);
nand U823 (N_823,N_410,N_353);
nand U824 (N_824,N_326,N_51);
nor U825 (N_825,N_16,N_52);
nand U826 (N_826,N_31,N_483);
and U827 (N_827,N_278,N_414);
nor U828 (N_828,N_142,N_34);
nand U829 (N_829,N_339,N_253);
nor U830 (N_830,N_232,N_371);
nand U831 (N_831,N_200,N_326);
nor U832 (N_832,N_383,N_53);
and U833 (N_833,N_332,N_350);
and U834 (N_834,N_328,N_5);
or U835 (N_835,N_401,N_206);
nor U836 (N_836,N_380,N_286);
nor U837 (N_837,N_19,N_496);
and U838 (N_838,N_326,N_323);
nor U839 (N_839,N_148,N_59);
nor U840 (N_840,N_10,N_257);
nor U841 (N_841,N_360,N_387);
nand U842 (N_842,N_439,N_49);
nor U843 (N_843,N_29,N_4);
or U844 (N_844,N_356,N_41);
nand U845 (N_845,N_204,N_447);
nor U846 (N_846,N_439,N_15);
and U847 (N_847,N_47,N_309);
or U848 (N_848,N_219,N_205);
nand U849 (N_849,N_289,N_212);
and U850 (N_850,N_356,N_50);
nor U851 (N_851,N_439,N_4);
nor U852 (N_852,N_60,N_383);
or U853 (N_853,N_41,N_137);
nand U854 (N_854,N_419,N_265);
nor U855 (N_855,N_111,N_135);
nor U856 (N_856,N_289,N_498);
or U857 (N_857,N_35,N_453);
or U858 (N_858,N_72,N_102);
nor U859 (N_859,N_262,N_98);
nand U860 (N_860,N_126,N_223);
nor U861 (N_861,N_22,N_349);
xnor U862 (N_862,N_315,N_480);
xor U863 (N_863,N_466,N_164);
nand U864 (N_864,N_159,N_412);
and U865 (N_865,N_122,N_376);
nor U866 (N_866,N_363,N_100);
nand U867 (N_867,N_75,N_84);
nor U868 (N_868,N_250,N_370);
and U869 (N_869,N_232,N_225);
nor U870 (N_870,N_158,N_128);
or U871 (N_871,N_87,N_7);
nor U872 (N_872,N_187,N_283);
nor U873 (N_873,N_460,N_255);
and U874 (N_874,N_202,N_323);
and U875 (N_875,N_254,N_364);
or U876 (N_876,N_481,N_1);
nand U877 (N_877,N_135,N_11);
and U878 (N_878,N_237,N_455);
or U879 (N_879,N_423,N_280);
and U880 (N_880,N_136,N_377);
or U881 (N_881,N_363,N_410);
nand U882 (N_882,N_372,N_143);
and U883 (N_883,N_127,N_404);
or U884 (N_884,N_127,N_120);
nor U885 (N_885,N_243,N_27);
and U886 (N_886,N_490,N_497);
nand U887 (N_887,N_25,N_294);
and U888 (N_888,N_438,N_102);
nand U889 (N_889,N_12,N_172);
nand U890 (N_890,N_83,N_188);
or U891 (N_891,N_447,N_439);
and U892 (N_892,N_245,N_258);
and U893 (N_893,N_338,N_2);
nand U894 (N_894,N_209,N_68);
nand U895 (N_895,N_102,N_478);
nor U896 (N_896,N_23,N_415);
and U897 (N_897,N_457,N_90);
or U898 (N_898,N_132,N_149);
nand U899 (N_899,N_183,N_298);
or U900 (N_900,N_356,N_275);
or U901 (N_901,N_213,N_58);
nand U902 (N_902,N_59,N_168);
nand U903 (N_903,N_478,N_75);
or U904 (N_904,N_77,N_294);
nor U905 (N_905,N_181,N_239);
nand U906 (N_906,N_214,N_405);
or U907 (N_907,N_365,N_261);
or U908 (N_908,N_261,N_81);
or U909 (N_909,N_374,N_194);
nor U910 (N_910,N_48,N_174);
xnor U911 (N_911,N_260,N_102);
nand U912 (N_912,N_36,N_149);
and U913 (N_913,N_389,N_194);
nor U914 (N_914,N_95,N_88);
or U915 (N_915,N_288,N_49);
or U916 (N_916,N_403,N_24);
or U917 (N_917,N_283,N_106);
or U918 (N_918,N_90,N_41);
nor U919 (N_919,N_208,N_276);
nand U920 (N_920,N_272,N_61);
nand U921 (N_921,N_7,N_252);
nor U922 (N_922,N_62,N_338);
nor U923 (N_923,N_368,N_410);
nand U924 (N_924,N_361,N_277);
nand U925 (N_925,N_367,N_145);
and U926 (N_926,N_348,N_428);
nand U927 (N_927,N_311,N_22);
and U928 (N_928,N_199,N_259);
nand U929 (N_929,N_290,N_226);
and U930 (N_930,N_196,N_19);
or U931 (N_931,N_297,N_46);
nand U932 (N_932,N_68,N_390);
nand U933 (N_933,N_199,N_497);
nor U934 (N_934,N_196,N_482);
nor U935 (N_935,N_444,N_89);
nor U936 (N_936,N_248,N_477);
nor U937 (N_937,N_379,N_249);
or U938 (N_938,N_397,N_200);
nand U939 (N_939,N_88,N_47);
or U940 (N_940,N_490,N_123);
nand U941 (N_941,N_408,N_217);
and U942 (N_942,N_190,N_394);
nor U943 (N_943,N_416,N_451);
nand U944 (N_944,N_472,N_81);
nor U945 (N_945,N_22,N_296);
and U946 (N_946,N_61,N_312);
or U947 (N_947,N_79,N_104);
and U948 (N_948,N_429,N_283);
and U949 (N_949,N_19,N_239);
nor U950 (N_950,N_414,N_250);
or U951 (N_951,N_193,N_116);
or U952 (N_952,N_248,N_410);
nor U953 (N_953,N_421,N_291);
or U954 (N_954,N_487,N_300);
nand U955 (N_955,N_396,N_364);
xor U956 (N_956,N_117,N_406);
or U957 (N_957,N_259,N_462);
nor U958 (N_958,N_212,N_342);
and U959 (N_959,N_261,N_349);
nor U960 (N_960,N_72,N_65);
and U961 (N_961,N_324,N_314);
or U962 (N_962,N_326,N_337);
nor U963 (N_963,N_311,N_379);
xor U964 (N_964,N_414,N_77);
nor U965 (N_965,N_486,N_60);
and U966 (N_966,N_412,N_279);
or U967 (N_967,N_216,N_116);
and U968 (N_968,N_285,N_203);
and U969 (N_969,N_204,N_496);
and U970 (N_970,N_231,N_64);
nand U971 (N_971,N_149,N_376);
and U972 (N_972,N_183,N_120);
or U973 (N_973,N_325,N_262);
and U974 (N_974,N_221,N_187);
or U975 (N_975,N_477,N_309);
or U976 (N_976,N_440,N_424);
nor U977 (N_977,N_207,N_183);
nor U978 (N_978,N_369,N_62);
nand U979 (N_979,N_116,N_442);
nand U980 (N_980,N_85,N_169);
and U981 (N_981,N_340,N_16);
nor U982 (N_982,N_406,N_258);
nand U983 (N_983,N_485,N_177);
nor U984 (N_984,N_338,N_19);
or U985 (N_985,N_211,N_370);
nand U986 (N_986,N_403,N_480);
nand U987 (N_987,N_497,N_292);
nand U988 (N_988,N_344,N_423);
nor U989 (N_989,N_202,N_250);
or U990 (N_990,N_480,N_355);
and U991 (N_991,N_365,N_325);
nor U992 (N_992,N_286,N_32);
or U993 (N_993,N_329,N_297);
and U994 (N_994,N_19,N_420);
or U995 (N_995,N_384,N_235);
nor U996 (N_996,N_217,N_293);
nor U997 (N_997,N_351,N_224);
or U998 (N_998,N_351,N_229);
nor U999 (N_999,N_357,N_16);
and U1000 (N_1000,N_968,N_749);
and U1001 (N_1001,N_708,N_798);
nand U1002 (N_1002,N_836,N_504);
nand U1003 (N_1003,N_817,N_540);
nor U1004 (N_1004,N_699,N_575);
nor U1005 (N_1005,N_818,N_519);
or U1006 (N_1006,N_594,N_885);
nand U1007 (N_1007,N_988,N_975);
and U1008 (N_1008,N_650,N_891);
nor U1009 (N_1009,N_837,N_720);
nand U1010 (N_1010,N_697,N_691);
or U1011 (N_1011,N_698,N_779);
nand U1012 (N_1012,N_671,N_913);
or U1013 (N_1013,N_998,N_538);
and U1014 (N_1014,N_741,N_992);
nand U1015 (N_1015,N_672,N_900);
and U1016 (N_1016,N_724,N_666);
or U1017 (N_1017,N_587,N_955);
nand U1018 (N_1018,N_703,N_535);
or U1019 (N_1019,N_870,N_729);
nor U1020 (N_1020,N_599,N_688);
xnor U1021 (N_1021,N_922,N_761);
or U1022 (N_1022,N_682,N_990);
or U1023 (N_1023,N_626,N_754);
and U1024 (N_1024,N_665,N_833);
and U1025 (N_1025,N_564,N_809);
and U1026 (N_1026,N_553,N_940);
xor U1027 (N_1027,N_502,N_571);
and U1028 (N_1028,N_570,N_591);
nor U1029 (N_1029,N_684,N_742);
nand U1030 (N_1030,N_911,N_795);
or U1031 (N_1031,N_869,N_927);
or U1032 (N_1032,N_547,N_947);
and U1033 (N_1033,N_614,N_893);
nand U1034 (N_1034,N_924,N_549);
or U1035 (N_1035,N_797,N_744);
or U1036 (N_1036,N_550,N_606);
or U1037 (N_1037,N_616,N_917);
and U1038 (N_1038,N_978,N_677);
and U1039 (N_1039,N_603,N_751);
and U1040 (N_1040,N_518,N_979);
nor U1041 (N_1041,N_581,N_812);
nand U1042 (N_1042,N_952,N_993);
or U1043 (N_1043,N_938,N_541);
nor U1044 (N_1044,N_679,N_989);
nand U1045 (N_1045,N_777,N_711);
nand U1046 (N_1046,N_643,N_826);
and U1047 (N_1047,N_892,N_901);
and U1048 (N_1048,N_690,N_658);
and U1049 (N_1049,N_558,N_838);
nand U1050 (N_1050,N_923,N_889);
and U1051 (N_1051,N_780,N_910);
and U1052 (N_1052,N_685,N_758);
and U1053 (N_1053,N_907,N_618);
nor U1054 (N_1054,N_858,N_775);
nor U1055 (N_1055,N_508,N_530);
and U1056 (N_1056,N_632,N_501);
xor U1057 (N_1057,N_568,N_661);
nand U1058 (N_1058,N_505,N_769);
and U1059 (N_1059,N_802,N_972);
and U1060 (N_1060,N_631,N_974);
nor U1061 (N_1061,N_772,N_759);
nor U1062 (N_1062,N_636,N_694);
and U1063 (N_1063,N_867,N_655);
nand U1064 (N_1064,N_531,N_546);
and U1065 (N_1065,N_552,N_732);
and U1066 (N_1066,N_670,N_987);
and U1067 (N_1067,N_880,N_719);
nor U1068 (N_1068,N_791,N_577);
and U1069 (N_1069,N_919,N_660);
nor U1070 (N_1070,N_945,N_920);
nand U1071 (N_1071,N_962,N_634);
xor U1072 (N_1072,N_561,N_799);
nor U1073 (N_1073,N_608,N_640);
nand U1074 (N_1074,N_601,N_840);
and U1075 (N_1075,N_536,N_537);
nor U1076 (N_1076,N_787,N_877);
nand U1077 (N_1077,N_942,N_909);
nand U1078 (N_1078,N_965,N_544);
or U1079 (N_1079,N_683,N_609);
nor U1080 (N_1080,N_980,N_808);
nor U1081 (N_1081,N_871,N_746);
nand U1082 (N_1082,N_706,N_957);
nand U1083 (N_1083,N_539,N_623);
and U1084 (N_1084,N_647,N_534);
nor U1085 (N_1085,N_997,N_839);
nor U1086 (N_1086,N_764,N_637);
nand U1087 (N_1087,N_981,N_805);
and U1088 (N_1088,N_948,N_600);
and U1089 (N_1089,N_586,N_578);
nand U1090 (N_1090,N_747,N_843);
or U1091 (N_1091,N_573,N_686);
or U1092 (N_1092,N_653,N_783);
nand U1093 (N_1093,N_876,N_710);
nand U1094 (N_1094,N_970,N_941);
and U1095 (N_1095,N_845,N_598);
and U1096 (N_1096,N_716,N_645);
xnor U1097 (N_1097,N_971,N_790);
and U1098 (N_1098,N_543,N_855);
nor U1099 (N_1099,N_832,N_718);
nor U1100 (N_1100,N_921,N_888);
nor U1101 (N_1101,N_695,N_673);
and U1102 (N_1102,N_523,N_905);
nand U1103 (N_1103,N_554,N_781);
or U1104 (N_1104,N_903,N_629);
nand U1105 (N_1105,N_659,N_734);
or U1106 (N_1106,N_983,N_596);
nor U1107 (N_1107,N_850,N_722);
or U1108 (N_1108,N_664,N_784);
nand U1109 (N_1109,N_932,N_675);
nor U1110 (N_1110,N_693,N_517);
and U1111 (N_1111,N_605,N_865);
nor U1112 (N_1112,N_887,N_961);
and U1113 (N_1113,N_574,N_681);
nor U1114 (N_1114,N_960,N_612);
or U1115 (N_1115,N_566,N_882);
nor U1116 (N_1116,N_740,N_620);
and U1117 (N_1117,N_611,N_651);
and U1118 (N_1118,N_762,N_813);
or U1119 (N_1119,N_739,N_883);
and U1120 (N_1120,N_792,N_933);
nand U1121 (N_1121,N_963,N_580);
and U1122 (N_1122,N_627,N_859);
nor U1123 (N_1123,N_757,N_819);
nand U1124 (N_1124,N_778,N_994);
nor U1125 (N_1125,N_615,N_667);
nand U1126 (N_1126,N_806,N_801);
nand U1127 (N_1127,N_966,N_565);
or U1128 (N_1128,N_656,N_854);
and U1129 (N_1129,N_735,N_515);
nor U1130 (N_1130,N_652,N_786);
and U1131 (N_1131,N_743,N_873);
or U1132 (N_1132,N_676,N_841);
nor U1133 (N_1133,N_943,N_804);
or U1134 (N_1134,N_999,N_521);
nor U1135 (N_1135,N_622,N_641);
or U1136 (N_1136,N_953,N_628);
and U1137 (N_1137,N_563,N_604);
nand U1138 (N_1138,N_902,N_834);
or U1139 (N_1139,N_793,N_814);
and U1140 (N_1140,N_856,N_825);
nand U1141 (N_1141,N_527,N_884);
xor U1142 (N_1142,N_593,N_642);
or U1143 (N_1143,N_824,N_890);
and U1144 (N_1144,N_898,N_712);
nand U1145 (N_1145,N_816,N_748);
nor U1146 (N_1146,N_525,N_984);
nand U1147 (N_1147,N_516,N_894);
and U1148 (N_1148,N_648,N_503);
nand U1149 (N_1149,N_860,N_847);
or U1150 (N_1150,N_916,N_576);
and U1151 (N_1151,N_602,N_526);
nor U1152 (N_1152,N_936,N_904);
nand U1153 (N_1153,N_853,N_709);
or U1154 (N_1154,N_560,N_912);
nand U1155 (N_1155,N_875,N_753);
and U1156 (N_1156,N_895,N_934);
and U1157 (N_1157,N_959,N_669);
or U1158 (N_1158,N_644,N_727);
nand U1159 (N_1159,N_830,N_862);
or U1160 (N_1160,N_954,N_794);
or U1161 (N_1161,N_507,N_678);
or U1162 (N_1162,N_680,N_589);
nor U1163 (N_1163,N_528,N_674);
nor U1164 (N_1164,N_638,N_949);
or U1165 (N_1165,N_996,N_595);
or U1166 (N_1166,N_937,N_701);
and U1167 (N_1167,N_931,N_689);
nor U1168 (N_1168,N_733,N_879);
nor U1169 (N_1169,N_506,N_548);
or U1170 (N_1170,N_976,N_821);
and U1171 (N_1171,N_950,N_908);
nand U1172 (N_1172,N_831,N_569);
or U1173 (N_1173,N_500,N_796);
nand U1174 (N_1174,N_995,N_533);
and U1175 (N_1175,N_621,N_991);
nor U1176 (N_1176,N_607,N_585);
nor U1177 (N_1177,N_977,N_767);
and U1178 (N_1178,N_785,N_878);
and U1179 (N_1179,N_861,N_800);
and U1180 (N_1180,N_633,N_696);
nor U1181 (N_1181,N_692,N_717);
nor U1182 (N_1182,N_823,N_588);
nor U1183 (N_1183,N_567,N_773);
or U1184 (N_1184,N_967,N_829);
nor U1185 (N_1185,N_738,N_545);
nand U1186 (N_1186,N_776,N_713);
nand U1187 (N_1187,N_617,N_662);
or U1188 (N_1188,N_509,N_635);
and U1189 (N_1189,N_848,N_771);
and U1190 (N_1190,N_866,N_597);
and U1191 (N_1191,N_846,N_925);
nor U1192 (N_1192,N_584,N_723);
nand U1193 (N_1193,N_745,N_789);
and U1194 (N_1194,N_619,N_572);
nand U1195 (N_1195,N_827,N_881);
nand U1196 (N_1196,N_964,N_520);
nor U1197 (N_1197,N_630,N_982);
and U1198 (N_1198,N_842,N_946);
and U1199 (N_1199,N_654,N_750);
and U1200 (N_1200,N_513,N_768);
and U1201 (N_1201,N_512,N_930);
nand U1202 (N_1202,N_700,N_728);
or U1203 (N_1203,N_852,N_803);
or U1204 (N_1204,N_529,N_774);
and U1205 (N_1205,N_951,N_649);
and U1206 (N_1206,N_583,N_973);
or U1207 (N_1207,N_510,N_551);
nor U1208 (N_1208,N_939,N_863);
nand U1209 (N_1209,N_755,N_857);
and U1210 (N_1210,N_872,N_592);
xnor U1211 (N_1211,N_582,N_726);
or U1212 (N_1212,N_807,N_969);
or U1213 (N_1213,N_899,N_944);
or U1214 (N_1214,N_828,N_935);
and U1215 (N_1215,N_704,N_730);
or U1216 (N_1216,N_765,N_897);
or U1217 (N_1217,N_926,N_815);
and U1218 (N_1218,N_524,N_864);
or U1219 (N_1219,N_736,N_752);
or U1220 (N_1220,N_956,N_687);
and U1221 (N_1221,N_820,N_522);
or U1222 (N_1222,N_760,N_707);
or U1223 (N_1223,N_914,N_851);
nand U1224 (N_1224,N_532,N_986);
or U1225 (N_1225,N_958,N_721);
nand U1226 (N_1226,N_613,N_929);
nand U1227 (N_1227,N_639,N_985);
nor U1228 (N_1228,N_657,N_702);
nand U1229 (N_1229,N_590,N_835);
nand U1230 (N_1230,N_663,N_788);
and U1231 (N_1231,N_725,N_844);
or U1232 (N_1232,N_668,N_542);
xor U1233 (N_1233,N_559,N_906);
and U1234 (N_1234,N_555,N_915);
nand U1235 (N_1235,N_514,N_886);
or U1236 (N_1236,N_928,N_849);
nand U1237 (N_1237,N_624,N_556);
nor U1238 (N_1238,N_610,N_646);
or U1239 (N_1239,N_810,N_782);
and U1240 (N_1240,N_705,N_511);
and U1241 (N_1241,N_714,N_822);
nor U1242 (N_1242,N_715,N_918);
or U1243 (N_1243,N_766,N_874);
and U1244 (N_1244,N_625,N_868);
and U1245 (N_1245,N_731,N_737);
or U1246 (N_1246,N_557,N_562);
or U1247 (N_1247,N_770,N_756);
nand U1248 (N_1248,N_579,N_763);
nand U1249 (N_1249,N_896,N_811);
nor U1250 (N_1250,N_730,N_785);
nand U1251 (N_1251,N_525,N_722);
or U1252 (N_1252,N_918,N_614);
nand U1253 (N_1253,N_975,N_594);
and U1254 (N_1254,N_503,N_812);
nor U1255 (N_1255,N_685,N_640);
nand U1256 (N_1256,N_990,N_918);
nor U1257 (N_1257,N_885,N_987);
nand U1258 (N_1258,N_967,N_869);
or U1259 (N_1259,N_952,N_698);
nand U1260 (N_1260,N_576,N_562);
xnor U1261 (N_1261,N_800,N_698);
or U1262 (N_1262,N_539,N_760);
nor U1263 (N_1263,N_987,N_932);
and U1264 (N_1264,N_852,N_886);
and U1265 (N_1265,N_862,N_624);
or U1266 (N_1266,N_846,N_546);
nor U1267 (N_1267,N_720,N_593);
and U1268 (N_1268,N_876,N_827);
nor U1269 (N_1269,N_855,N_739);
and U1270 (N_1270,N_917,N_560);
or U1271 (N_1271,N_838,N_871);
nand U1272 (N_1272,N_548,N_783);
nor U1273 (N_1273,N_844,N_956);
nand U1274 (N_1274,N_610,N_633);
nor U1275 (N_1275,N_655,N_579);
and U1276 (N_1276,N_919,N_784);
and U1277 (N_1277,N_576,N_591);
or U1278 (N_1278,N_948,N_677);
nor U1279 (N_1279,N_894,N_781);
nand U1280 (N_1280,N_967,N_763);
or U1281 (N_1281,N_922,N_938);
nor U1282 (N_1282,N_963,N_734);
or U1283 (N_1283,N_747,N_696);
and U1284 (N_1284,N_786,N_926);
nand U1285 (N_1285,N_730,N_988);
and U1286 (N_1286,N_546,N_737);
nor U1287 (N_1287,N_545,N_594);
or U1288 (N_1288,N_507,N_897);
nor U1289 (N_1289,N_901,N_686);
nand U1290 (N_1290,N_748,N_789);
and U1291 (N_1291,N_648,N_718);
or U1292 (N_1292,N_831,N_801);
nand U1293 (N_1293,N_866,N_848);
nand U1294 (N_1294,N_890,N_849);
or U1295 (N_1295,N_899,N_715);
nand U1296 (N_1296,N_911,N_950);
or U1297 (N_1297,N_584,N_658);
or U1298 (N_1298,N_759,N_663);
nand U1299 (N_1299,N_920,N_803);
nor U1300 (N_1300,N_516,N_661);
and U1301 (N_1301,N_947,N_932);
nand U1302 (N_1302,N_878,N_883);
and U1303 (N_1303,N_738,N_535);
nor U1304 (N_1304,N_662,N_923);
and U1305 (N_1305,N_583,N_938);
nand U1306 (N_1306,N_673,N_591);
or U1307 (N_1307,N_933,N_808);
nor U1308 (N_1308,N_821,N_914);
and U1309 (N_1309,N_788,N_873);
nor U1310 (N_1310,N_754,N_776);
nor U1311 (N_1311,N_715,N_882);
nor U1312 (N_1312,N_816,N_850);
nor U1313 (N_1313,N_977,N_583);
nor U1314 (N_1314,N_682,N_517);
or U1315 (N_1315,N_667,N_883);
nor U1316 (N_1316,N_654,N_551);
nand U1317 (N_1317,N_780,N_582);
nor U1318 (N_1318,N_975,N_836);
or U1319 (N_1319,N_816,N_654);
nand U1320 (N_1320,N_686,N_836);
and U1321 (N_1321,N_539,N_690);
nor U1322 (N_1322,N_960,N_739);
nand U1323 (N_1323,N_578,N_699);
nor U1324 (N_1324,N_631,N_546);
or U1325 (N_1325,N_599,N_952);
or U1326 (N_1326,N_910,N_757);
and U1327 (N_1327,N_631,N_724);
or U1328 (N_1328,N_856,N_797);
or U1329 (N_1329,N_997,N_552);
nor U1330 (N_1330,N_529,N_911);
or U1331 (N_1331,N_860,N_859);
nor U1332 (N_1332,N_559,N_793);
and U1333 (N_1333,N_925,N_960);
nand U1334 (N_1334,N_961,N_776);
and U1335 (N_1335,N_872,N_809);
or U1336 (N_1336,N_549,N_582);
nand U1337 (N_1337,N_749,N_922);
or U1338 (N_1338,N_899,N_967);
nand U1339 (N_1339,N_736,N_907);
and U1340 (N_1340,N_956,N_834);
and U1341 (N_1341,N_579,N_718);
and U1342 (N_1342,N_555,N_984);
and U1343 (N_1343,N_733,N_526);
nor U1344 (N_1344,N_562,N_551);
and U1345 (N_1345,N_856,N_520);
nand U1346 (N_1346,N_604,N_627);
nand U1347 (N_1347,N_731,N_817);
or U1348 (N_1348,N_578,N_603);
or U1349 (N_1349,N_804,N_620);
and U1350 (N_1350,N_542,N_715);
or U1351 (N_1351,N_960,N_973);
nand U1352 (N_1352,N_510,N_549);
and U1353 (N_1353,N_674,N_775);
nand U1354 (N_1354,N_759,N_501);
nor U1355 (N_1355,N_668,N_588);
nor U1356 (N_1356,N_619,N_782);
or U1357 (N_1357,N_897,N_643);
or U1358 (N_1358,N_592,N_739);
and U1359 (N_1359,N_758,N_669);
nand U1360 (N_1360,N_766,N_793);
nor U1361 (N_1361,N_776,N_968);
and U1362 (N_1362,N_831,N_889);
or U1363 (N_1363,N_752,N_734);
and U1364 (N_1364,N_785,N_721);
or U1365 (N_1365,N_544,N_844);
and U1366 (N_1366,N_613,N_524);
nand U1367 (N_1367,N_596,N_885);
and U1368 (N_1368,N_536,N_883);
or U1369 (N_1369,N_791,N_806);
nand U1370 (N_1370,N_599,N_610);
nor U1371 (N_1371,N_770,N_980);
nand U1372 (N_1372,N_662,N_886);
or U1373 (N_1373,N_559,N_692);
and U1374 (N_1374,N_795,N_981);
and U1375 (N_1375,N_509,N_719);
and U1376 (N_1376,N_523,N_662);
nor U1377 (N_1377,N_834,N_661);
and U1378 (N_1378,N_826,N_814);
nor U1379 (N_1379,N_723,N_857);
nand U1380 (N_1380,N_617,N_666);
or U1381 (N_1381,N_746,N_998);
or U1382 (N_1382,N_622,N_776);
nand U1383 (N_1383,N_697,N_905);
nand U1384 (N_1384,N_997,N_876);
or U1385 (N_1385,N_723,N_825);
and U1386 (N_1386,N_999,N_763);
nand U1387 (N_1387,N_673,N_669);
nand U1388 (N_1388,N_731,N_568);
or U1389 (N_1389,N_978,N_865);
and U1390 (N_1390,N_807,N_817);
nand U1391 (N_1391,N_807,N_689);
nor U1392 (N_1392,N_913,N_786);
nor U1393 (N_1393,N_837,N_871);
and U1394 (N_1394,N_743,N_795);
nor U1395 (N_1395,N_723,N_551);
nand U1396 (N_1396,N_683,N_682);
and U1397 (N_1397,N_634,N_513);
xor U1398 (N_1398,N_801,N_917);
xor U1399 (N_1399,N_635,N_885);
nand U1400 (N_1400,N_813,N_781);
nor U1401 (N_1401,N_685,N_975);
and U1402 (N_1402,N_971,N_764);
nor U1403 (N_1403,N_536,N_789);
or U1404 (N_1404,N_914,N_502);
and U1405 (N_1405,N_913,N_761);
or U1406 (N_1406,N_763,N_709);
or U1407 (N_1407,N_803,N_577);
or U1408 (N_1408,N_509,N_503);
nor U1409 (N_1409,N_658,N_797);
or U1410 (N_1410,N_887,N_621);
or U1411 (N_1411,N_808,N_626);
nor U1412 (N_1412,N_710,N_645);
nor U1413 (N_1413,N_822,N_750);
nor U1414 (N_1414,N_790,N_562);
or U1415 (N_1415,N_941,N_990);
nor U1416 (N_1416,N_890,N_915);
and U1417 (N_1417,N_961,N_506);
nand U1418 (N_1418,N_996,N_579);
nor U1419 (N_1419,N_865,N_901);
nor U1420 (N_1420,N_866,N_820);
nor U1421 (N_1421,N_588,N_657);
nor U1422 (N_1422,N_842,N_933);
or U1423 (N_1423,N_900,N_883);
nand U1424 (N_1424,N_765,N_870);
nor U1425 (N_1425,N_781,N_740);
nand U1426 (N_1426,N_897,N_767);
nand U1427 (N_1427,N_789,N_854);
nand U1428 (N_1428,N_829,N_699);
nor U1429 (N_1429,N_572,N_816);
and U1430 (N_1430,N_953,N_663);
or U1431 (N_1431,N_617,N_865);
or U1432 (N_1432,N_695,N_524);
and U1433 (N_1433,N_929,N_915);
nor U1434 (N_1434,N_967,N_837);
nor U1435 (N_1435,N_929,N_808);
and U1436 (N_1436,N_746,N_848);
or U1437 (N_1437,N_575,N_847);
and U1438 (N_1438,N_694,N_549);
and U1439 (N_1439,N_929,N_962);
nand U1440 (N_1440,N_784,N_698);
nor U1441 (N_1441,N_815,N_662);
nand U1442 (N_1442,N_721,N_793);
nand U1443 (N_1443,N_991,N_890);
or U1444 (N_1444,N_742,N_654);
and U1445 (N_1445,N_980,N_891);
and U1446 (N_1446,N_531,N_731);
nor U1447 (N_1447,N_878,N_918);
or U1448 (N_1448,N_929,N_836);
or U1449 (N_1449,N_667,N_821);
nand U1450 (N_1450,N_648,N_989);
nor U1451 (N_1451,N_676,N_717);
or U1452 (N_1452,N_888,N_692);
nand U1453 (N_1453,N_931,N_712);
and U1454 (N_1454,N_598,N_927);
and U1455 (N_1455,N_694,N_655);
nand U1456 (N_1456,N_938,N_880);
nand U1457 (N_1457,N_650,N_870);
nand U1458 (N_1458,N_640,N_821);
nand U1459 (N_1459,N_809,N_634);
nor U1460 (N_1460,N_531,N_902);
nor U1461 (N_1461,N_850,N_758);
or U1462 (N_1462,N_965,N_740);
nor U1463 (N_1463,N_558,N_837);
and U1464 (N_1464,N_521,N_817);
and U1465 (N_1465,N_589,N_578);
nand U1466 (N_1466,N_809,N_861);
and U1467 (N_1467,N_569,N_685);
or U1468 (N_1468,N_966,N_984);
nand U1469 (N_1469,N_830,N_916);
nor U1470 (N_1470,N_767,N_946);
nor U1471 (N_1471,N_752,N_751);
xor U1472 (N_1472,N_927,N_676);
nor U1473 (N_1473,N_557,N_685);
and U1474 (N_1474,N_873,N_948);
and U1475 (N_1475,N_752,N_844);
and U1476 (N_1476,N_691,N_941);
and U1477 (N_1477,N_564,N_861);
nor U1478 (N_1478,N_879,N_828);
or U1479 (N_1479,N_876,N_903);
nand U1480 (N_1480,N_515,N_722);
and U1481 (N_1481,N_528,N_582);
nor U1482 (N_1482,N_752,N_910);
or U1483 (N_1483,N_617,N_503);
nor U1484 (N_1484,N_950,N_861);
or U1485 (N_1485,N_946,N_753);
nand U1486 (N_1486,N_617,N_540);
and U1487 (N_1487,N_955,N_584);
or U1488 (N_1488,N_986,N_981);
nand U1489 (N_1489,N_871,N_934);
and U1490 (N_1490,N_888,N_880);
or U1491 (N_1491,N_577,N_758);
or U1492 (N_1492,N_714,N_698);
or U1493 (N_1493,N_666,N_615);
nand U1494 (N_1494,N_943,N_668);
nand U1495 (N_1495,N_918,N_521);
or U1496 (N_1496,N_811,N_721);
and U1497 (N_1497,N_624,N_673);
or U1498 (N_1498,N_518,N_559);
or U1499 (N_1499,N_782,N_696);
nor U1500 (N_1500,N_1232,N_1423);
or U1501 (N_1501,N_1397,N_1078);
nor U1502 (N_1502,N_1049,N_1058);
and U1503 (N_1503,N_1344,N_1082);
nand U1504 (N_1504,N_1240,N_1434);
and U1505 (N_1505,N_1160,N_1107);
nor U1506 (N_1506,N_1334,N_1044);
or U1507 (N_1507,N_1452,N_1282);
nor U1508 (N_1508,N_1348,N_1306);
nand U1509 (N_1509,N_1438,N_1229);
or U1510 (N_1510,N_1002,N_1319);
and U1511 (N_1511,N_1329,N_1014);
nor U1512 (N_1512,N_1093,N_1497);
or U1513 (N_1513,N_1451,N_1026);
and U1514 (N_1514,N_1361,N_1198);
or U1515 (N_1515,N_1390,N_1439);
nor U1516 (N_1516,N_1013,N_1033);
nand U1517 (N_1517,N_1285,N_1369);
or U1518 (N_1518,N_1293,N_1405);
or U1519 (N_1519,N_1021,N_1071);
and U1520 (N_1520,N_1478,N_1092);
nor U1521 (N_1521,N_1322,N_1458);
or U1522 (N_1522,N_1430,N_1387);
or U1523 (N_1523,N_1327,N_1420);
nor U1524 (N_1524,N_1455,N_1350);
and U1525 (N_1525,N_1004,N_1426);
nand U1526 (N_1526,N_1403,N_1254);
nand U1527 (N_1527,N_1165,N_1170);
nor U1528 (N_1528,N_1011,N_1089);
or U1529 (N_1529,N_1087,N_1370);
or U1530 (N_1530,N_1340,N_1034);
nand U1531 (N_1531,N_1362,N_1494);
nor U1532 (N_1532,N_1163,N_1166);
or U1533 (N_1533,N_1302,N_1228);
nor U1534 (N_1534,N_1111,N_1437);
and U1535 (N_1535,N_1338,N_1133);
and U1536 (N_1536,N_1268,N_1417);
and U1537 (N_1537,N_1446,N_1355);
xor U1538 (N_1538,N_1227,N_1091);
nand U1539 (N_1539,N_1490,N_1029);
nand U1540 (N_1540,N_1248,N_1485);
nand U1541 (N_1541,N_1180,N_1395);
or U1542 (N_1542,N_1114,N_1492);
or U1543 (N_1543,N_1171,N_1183);
and U1544 (N_1544,N_1202,N_1073);
and U1545 (N_1545,N_1207,N_1023);
or U1546 (N_1546,N_1496,N_1276);
and U1547 (N_1547,N_1298,N_1193);
nor U1548 (N_1548,N_1121,N_1190);
or U1549 (N_1549,N_1252,N_1373);
and U1550 (N_1550,N_1330,N_1470);
or U1551 (N_1551,N_1129,N_1131);
nand U1552 (N_1552,N_1135,N_1048);
nor U1553 (N_1553,N_1483,N_1043);
and U1554 (N_1554,N_1055,N_1052);
or U1555 (N_1555,N_1309,N_1411);
nor U1556 (N_1556,N_1214,N_1375);
or U1557 (N_1557,N_1220,N_1132);
nand U1558 (N_1558,N_1216,N_1262);
nand U1559 (N_1559,N_1466,N_1408);
nand U1560 (N_1560,N_1341,N_1155);
nand U1561 (N_1561,N_1108,N_1196);
or U1562 (N_1562,N_1006,N_1213);
or U1563 (N_1563,N_1365,N_1461);
or U1564 (N_1564,N_1393,N_1404);
or U1565 (N_1565,N_1443,N_1098);
or U1566 (N_1566,N_1360,N_1331);
nor U1567 (N_1567,N_1316,N_1305);
or U1568 (N_1568,N_1187,N_1012);
and U1569 (N_1569,N_1041,N_1459);
nand U1570 (N_1570,N_1473,N_1112);
nor U1571 (N_1571,N_1357,N_1474);
and U1572 (N_1572,N_1223,N_1476);
nand U1573 (N_1573,N_1182,N_1152);
nand U1574 (N_1574,N_1057,N_1323);
and U1575 (N_1575,N_1457,N_1005);
xnor U1576 (N_1576,N_1480,N_1045);
nor U1577 (N_1577,N_1241,N_1454);
or U1578 (N_1578,N_1136,N_1283);
nand U1579 (N_1579,N_1346,N_1139);
nor U1580 (N_1580,N_1032,N_1286);
or U1581 (N_1581,N_1462,N_1016);
and U1582 (N_1582,N_1488,N_1389);
or U1583 (N_1583,N_1491,N_1156);
nor U1584 (N_1584,N_1096,N_1063);
nor U1585 (N_1585,N_1095,N_1471);
or U1586 (N_1586,N_1027,N_1315);
nor U1587 (N_1587,N_1211,N_1413);
and U1588 (N_1588,N_1412,N_1000);
and U1589 (N_1589,N_1303,N_1304);
and U1590 (N_1590,N_1402,N_1209);
and U1591 (N_1591,N_1435,N_1074);
and U1592 (N_1592,N_1090,N_1313);
or U1593 (N_1593,N_1410,N_1288);
or U1594 (N_1594,N_1146,N_1053);
nand U1595 (N_1595,N_1290,N_1167);
and U1596 (N_1596,N_1022,N_1249);
nand U1597 (N_1597,N_1294,N_1308);
and U1598 (N_1598,N_1253,N_1359);
and U1599 (N_1599,N_1115,N_1158);
and U1600 (N_1600,N_1374,N_1448);
and U1601 (N_1601,N_1210,N_1008);
and U1602 (N_1602,N_1105,N_1311);
and U1603 (N_1603,N_1363,N_1173);
or U1604 (N_1604,N_1077,N_1427);
and U1605 (N_1605,N_1257,N_1320);
and U1606 (N_1606,N_1218,N_1384);
nor U1607 (N_1607,N_1259,N_1328);
and U1608 (N_1608,N_1177,N_1342);
nor U1609 (N_1609,N_1356,N_1056);
and U1610 (N_1610,N_1201,N_1270);
and U1611 (N_1611,N_1498,N_1036);
nand U1612 (N_1612,N_1347,N_1398);
nor U1613 (N_1613,N_1019,N_1150);
and U1614 (N_1614,N_1159,N_1025);
nand U1615 (N_1615,N_1366,N_1123);
nand U1616 (N_1616,N_1097,N_1113);
nand U1617 (N_1617,N_1261,N_1083);
nand U1618 (N_1618,N_1181,N_1212);
nor U1619 (N_1619,N_1142,N_1120);
or U1620 (N_1620,N_1274,N_1318);
or U1621 (N_1621,N_1392,N_1310);
nand U1622 (N_1622,N_1186,N_1239);
xor U1623 (N_1623,N_1194,N_1100);
nor U1624 (N_1624,N_1039,N_1128);
nand U1625 (N_1625,N_1487,N_1242);
and U1626 (N_1626,N_1381,N_1453);
or U1627 (N_1627,N_1238,N_1493);
and U1628 (N_1628,N_1028,N_1038);
nand U1629 (N_1629,N_1419,N_1151);
nor U1630 (N_1630,N_1157,N_1208);
and U1631 (N_1631,N_1064,N_1335);
and U1632 (N_1632,N_1371,N_1275);
or U1633 (N_1633,N_1024,N_1380);
nor U1634 (N_1634,N_1247,N_1400);
nand U1635 (N_1635,N_1042,N_1317);
or U1636 (N_1636,N_1143,N_1010);
nand U1637 (N_1637,N_1189,N_1267);
or U1638 (N_1638,N_1060,N_1364);
or U1639 (N_1639,N_1376,N_1351);
and U1640 (N_1640,N_1422,N_1300);
nor U1641 (N_1641,N_1424,N_1367);
nor U1642 (N_1642,N_1484,N_1046);
and U1643 (N_1643,N_1106,N_1069);
nand U1644 (N_1644,N_1429,N_1301);
nor U1645 (N_1645,N_1250,N_1388);
nor U1646 (N_1646,N_1409,N_1345);
nand U1647 (N_1647,N_1126,N_1450);
and U1648 (N_1648,N_1179,N_1172);
nor U1649 (N_1649,N_1110,N_1117);
nor U1650 (N_1650,N_1061,N_1103);
nor U1651 (N_1651,N_1407,N_1076);
or U1652 (N_1652,N_1349,N_1226);
nand U1653 (N_1653,N_1333,N_1176);
and U1654 (N_1654,N_1003,N_1030);
or U1655 (N_1655,N_1234,N_1066);
nand U1656 (N_1656,N_1486,N_1079);
and U1657 (N_1657,N_1145,N_1251);
or U1658 (N_1658,N_1237,N_1125);
nand U1659 (N_1659,N_1007,N_1312);
and U1660 (N_1660,N_1225,N_1062);
nor U1661 (N_1661,N_1447,N_1065);
and U1662 (N_1662,N_1445,N_1192);
nor U1663 (N_1663,N_1258,N_1051);
nand U1664 (N_1664,N_1382,N_1017);
and U1665 (N_1665,N_1084,N_1224);
and U1666 (N_1666,N_1432,N_1260);
and U1667 (N_1667,N_1280,N_1266);
nand U1668 (N_1668,N_1343,N_1094);
nor U1669 (N_1669,N_1001,N_1378);
or U1670 (N_1670,N_1436,N_1020);
or U1671 (N_1671,N_1215,N_1130);
nand U1672 (N_1672,N_1292,N_1205);
nand U1673 (N_1673,N_1144,N_1119);
and U1674 (N_1674,N_1379,N_1314);
and U1675 (N_1675,N_1200,N_1099);
or U1676 (N_1676,N_1399,N_1161);
nor U1677 (N_1677,N_1421,N_1281);
nand U1678 (N_1678,N_1230,N_1164);
nand U1679 (N_1679,N_1217,N_1219);
nand U1680 (N_1680,N_1264,N_1456);
nand U1681 (N_1681,N_1174,N_1354);
and U1682 (N_1682,N_1243,N_1465);
and U1683 (N_1683,N_1386,N_1441);
nor U1684 (N_1684,N_1047,N_1277);
nand U1685 (N_1685,N_1206,N_1153);
and U1686 (N_1686,N_1289,N_1352);
nor U1687 (N_1687,N_1269,N_1050);
or U1688 (N_1688,N_1406,N_1287);
and U1689 (N_1689,N_1460,N_1279);
or U1690 (N_1690,N_1178,N_1244);
nand U1691 (N_1691,N_1358,N_1231);
nor U1692 (N_1692,N_1321,N_1442);
nor U1693 (N_1693,N_1222,N_1086);
nand U1694 (N_1694,N_1265,N_1278);
nand U1695 (N_1695,N_1168,N_1468);
nand U1696 (N_1696,N_1203,N_1297);
or U1697 (N_1697,N_1175,N_1383);
or U1698 (N_1698,N_1273,N_1263);
nand U1699 (N_1699,N_1477,N_1464);
or U1700 (N_1700,N_1147,N_1499);
nor U1701 (N_1701,N_1059,N_1284);
nand U1702 (N_1702,N_1116,N_1122);
nand U1703 (N_1703,N_1101,N_1118);
and U1704 (N_1704,N_1124,N_1080);
and U1705 (N_1705,N_1009,N_1337);
or U1706 (N_1706,N_1489,N_1326);
and U1707 (N_1707,N_1188,N_1031);
nor U1708 (N_1708,N_1271,N_1256);
or U1709 (N_1709,N_1054,N_1204);
and U1710 (N_1710,N_1197,N_1035);
and U1711 (N_1711,N_1481,N_1472);
or U1712 (N_1712,N_1127,N_1444);
or U1713 (N_1713,N_1394,N_1440);
and U1714 (N_1714,N_1233,N_1141);
and U1715 (N_1715,N_1291,N_1495);
nand U1716 (N_1716,N_1085,N_1162);
and U1717 (N_1717,N_1140,N_1236);
nand U1718 (N_1718,N_1414,N_1037);
or U1719 (N_1719,N_1148,N_1015);
or U1720 (N_1720,N_1353,N_1385);
and U1721 (N_1721,N_1324,N_1449);
nand U1722 (N_1722,N_1235,N_1425);
and U1723 (N_1723,N_1255,N_1199);
nor U1724 (N_1724,N_1245,N_1109);
and U1725 (N_1725,N_1040,N_1272);
nor U1726 (N_1726,N_1088,N_1296);
nor U1727 (N_1727,N_1068,N_1169);
nand U1728 (N_1728,N_1184,N_1154);
and U1729 (N_1729,N_1339,N_1081);
nand U1730 (N_1730,N_1102,N_1368);
nand U1731 (N_1731,N_1325,N_1018);
nand U1732 (N_1732,N_1469,N_1482);
or U1733 (N_1733,N_1070,N_1332);
and U1734 (N_1734,N_1137,N_1391);
nand U1735 (N_1735,N_1415,N_1134);
nor U1736 (N_1736,N_1416,N_1377);
xor U1737 (N_1737,N_1295,N_1191);
and U1738 (N_1738,N_1401,N_1463);
and U1739 (N_1739,N_1433,N_1299);
and U1740 (N_1740,N_1138,N_1221);
nand U1741 (N_1741,N_1149,N_1307);
nand U1742 (N_1742,N_1475,N_1195);
or U1743 (N_1743,N_1418,N_1104);
nand U1744 (N_1744,N_1372,N_1246);
or U1745 (N_1745,N_1428,N_1467);
and U1746 (N_1746,N_1336,N_1479);
nand U1747 (N_1747,N_1072,N_1185);
nand U1748 (N_1748,N_1396,N_1075);
nand U1749 (N_1749,N_1431,N_1067);
nand U1750 (N_1750,N_1108,N_1401);
and U1751 (N_1751,N_1418,N_1188);
or U1752 (N_1752,N_1225,N_1124);
nor U1753 (N_1753,N_1001,N_1389);
nor U1754 (N_1754,N_1085,N_1107);
nand U1755 (N_1755,N_1033,N_1329);
nor U1756 (N_1756,N_1006,N_1037);
nand U1757 (N_1757,N_1259,N_1402);
or U1758 (N_1758,N_1340,N_1140);
or U1759 (N_1759,N_1309,N_1005);
nor U1760 (N_1760,N_1157,N_1469);
nor U1761 (N_1761,N_1067,N_1217);
nand U1762 (N_1762,N_1448,N_1421);
nor U1763 (N_1763,N_1056,N_1152);
or U1764 (N_1764,N_1205,N_1427);
and U1765 (N_1765,N_1217,N_1475);
and U1766 (N_1766,N_1321,N_1368);
and U1767 (N_1767,N_1154,N_1055);
nand U1768 (N_1768,N_1095,N_1377);
and U1769 (N_1769,N_1330,N_1061);
and U1770 (N_1770,N_1483,N_1131);
nor U1771 (N_1771,N_1117,N_1371);
nor U1772 (N_1772,N_1257,N_1326);
nor U1773 (N_1773,N_1068,N_1482);
and U1774 (N_1774,N_1039,N_1471);
or U1775 (N_1775,N_1208,N_1054);
or U1776 (N_1776,N_1339,N_1292);
and U1777 (N_1777,N_1231,N_1451);
and U1778 (N_1778,N_1142,N_1246);
or U1779 (N_1779,N_1122,N_1400);
nor U1780 (N_1780,N_1092,N_1257);
and U1781 (N_1781,N_1118,N_1059);
or U1782 (N_1782,N_1400,N_1453);
and U1783 (N_1783,N_1262,N_1437);
and U1784 (N_1784,N_1205,N_1431);
nand U1785 (N_1785,N_1275,N_1062);
nand U1786 (N_1786,N_1357,N_1495);
and U1787 (N_1787,N_1415,N_1480);
or U1788 (N_1788,N_1332,N_1236);
or U1789 (N_1789,N_1056,N_1405);
and U1790 (N_1790,N_1484,N_1377);
or U1791 (N_1791,N_1176,N_1138);
or U1792 (N_1792,N_1220,N_1320);
or U1793 (N_1793,N_1067,N_1475);
and U1794 (N_1794,N_1308,N_1132);
and U1795 (N_1795,N_1188,N_1427);
nor U1796 (N_1796,N_1306,N_1074);
and U1797 (N_1797,N_1418,N_1386);
and U1798 (N_1798,N_1128,N_1216);
nor U1799 (N_1799,N_1450,N_1363);
nand U1800 (N_1800,N_1345,N_1455);
or U1801 (N_1801,N_1190,N_1473);
nand U1802 (N_1802,N_1218,N_1494);
or U1803 (N_1803,N_1079,N_1260);
and U1804 (N_1804,N_1159,N_1007);
nand U1805 (N_1805,N_1410,N_1185);
or U1806 (N_1806,N_1105,N_1049);
and U1807 (N_1807,N_1036,N_1391);
nor U1808 (N_1808,N_1052,N_1410);
or U1809 (N_1809,N_1355,N_1171);
nand U1810 (N_1810,N_1454,N_1178);
and U1811 (N_1811,N_1141,N_1303);
or U1812 (N_1812,N_1244,N_1149);
nor U1813 (N_1813,N_1332,N_1179);
nor U1814 (N_1814,N_1225,N_1215);
or U1815 (N_1815,N_1287,N_1175);
and U1816 (N_1816,N_1017,N_1340);
and U1817 (N_1817,N_1047,N_1413);
or U1818 (N_1818,N_1016,N_1158);
and U1819 (N_1819,N_1390,N_1496);
and U1820 (N_1820,N_1079,N_1308);
nand U1821 (N_1821,N_1038,N_1469);
nand U1822 (N_1822,N_1189,N_1235);
nand U1823 (N_1823,N_1204,N_1459);
and U1824 (N_1824,N_1408,N_1054);
and U1825 (N_1825,N_1426,N_1042);
nor U1826 (N_1826,N_1155,N_1490);
nor U1827 (N_1827,N_1455,N_1002);
and U1828 (N_1828,N_1313,N_1050);
nand U1829 (N_1829,N_1384,N_1072);
nor U1830 (N_1830,N_1270,N_1317);
and U1831 (N_1831,N_1142,N_1191);
and U1832 (N_1832,N_1201,N_1180);
or U1833 (N_1833,N_1288,N_1419);
nand U1834 (N_1834,N_1233,N_1304);
or U1835 (N_1835,N_1493,N_1187);
nand U1836 (N_1836,N_1256,N_1411);
and U1837 (N_1837,N_1160,N_1157);
or U1838 (N_1838,N_1366,N_1382);
or U1839 (N_1839,N_1401,N_1304);
nor U1840 (N_1840,N_1071,N_1184);
nand U1841 (N_1841,N_1161,N_1082);
and U1842 (N_1842,N_1128,N_1025);
nor U1843 (N_1843,N_1228,N_1495);
nand U1844 (N_1844,N_1360,N_1385);
nor U1845 (N_1845,N_1007,N_1054);
or U1846 (N_1846,N_1235,N_1245);
nand U1847 (N_1847,N_1209,N_1371);
and U1848 (N_1848,N_1301,N_1373);
and U1849 (N_1849,N_1350,N_1299);
or U1850 (N_1850,N_1406,N_1092);
and U1851 (N_1851,N_1036,N_1090);
or U1852 (N_1852,N_1399,N_1170);
nor U1853 (N_1853,N_1203,N_1429);
and U1854 (N_1854,N_1221,N_1427);
and U1855 (N_1855,N_1448,N_1219);
or U1856 (N_1856,N_1026,N_1155);
nand U1857 (N_1857,N_1431,N_1369);
nand U1858 (N_1858,N_1006,N_1057);
nor U1859 (N_1859,N_1449,N_1340);
nor U1860 (N_1860,N_1203,N_1210);
nor U1861 (N_1861,N_1257,N_1082);
nor U1862 (N_1862,N_1233,N_1053);
nand U1863 (N_1863,N_1275,N_1395);
and U1864 (N_1864,N_1478,N_1473);
nor U1865 (N_1865,N_1296,N_1369);
or U1866 (N_1866,N_1347,N_1061);
or U1867 (N_1867,N_1176,N_1103);
nor U1868 (N_1868,N_1236,N_1399);
nand U1869 (N_1869,N_1121,N_1438);
and U1870 (N_1870,N_1053,N_1252);
nor U1871 (N_1871,N_1324,N_1450);
and U1872 (N_1872,N_1168,N_1496);
and U1873 (N_1873,N_1109,N_1252);
nand U1874 (N_1874,N_1020,N_1430);
nor U1875 (N_1875,N_1063,N_1301);
and U1876 (N_1876,N_1172,N_1223);
and U1877 (N_1877,N_1441,N_1253);
nor U1878 (N_1878,N_1180,N_1126);
nand U1879 (N_1879,N_1001,N_1076);
nor U1880 (N_1880,N_1018,N_1410);
nor U1881 (N_1881,N_1291,N_1209);
and U1882 (N_1882,N_1321,N_1406);
or U1883 (N_1883,N_1399,N_1182);
nor U1884 (N_1884,N_1467,N_1431);
and U1885 (N_1885,N_1430,N_1116);
and U1886 (N_1886,N_1231,N_1105);
or U1887 (N_1887,N_1238,N_1496);
nor U1888 (N_1888,N_1129,N_1217);
nor U1889 (N_1889,N_1085,N_1417);
and U1890 (N_1890,N_1256,N_1313);
or U1891 (N_1891,N_1247,N_1358);
nor U1892 (N_1892,N_1294,N_1459);
nand U1893 (N_1893,N_1076,N_1430);
nand U1894 (N_1894,N_1366,N_1318);
and U1895 (N_1895,N_1484,N_1417);
or U1896 (N_1896,N_1491,N_1454);
nand U1897 (N_1897,N_1141,N_1319);
and U1898 (N_1898,N_1497,N_1437);
and U1899 (N_1899,N_1298,N_1203);
and U1900 (N_1900,N_1467,N_1140);
or U1901 (N_1901,N_1139,N_1029);
and U1902 (N_1902,N_1313,N_1151);
or U1903 (N_1903,N_1244,N_1074);
and U1904 (N_1904,N_1233,N_1187);
nand U1905 (N_1905,N_1348,N_1059);
or U1906 (N_1906,N_1297,N_1166);
xnor U1907 (N_1907,N_1350,N_1132);
and U1908 (N_1908,N_1343,N_1048);
nand U1909 (N_1909,N_1384,N_1076);
nand U1910 (N_1910,N_1289,N_1031);
or U1911 (N_1911,N_1130,N_1347);
or U1912 (N_1912,N_1062,N_1029);
or U1913 (N_1913,N_1250,N_1268);
or U1914 (N_1914,N_1009,N_1046);
nand U1915 (N_1915,N_1195,N_1179);
nand U1916 (N_1916,N_1305,N_1336);
nor U1917 (N_1917,N_1359,N_1135);
and U1918 (N_1918,N_1165,N_1068);
or U1919 (N_1919,N_1288,N_1382);
and U1920 (N_1920,N_1340,N_1387);
nand U1921 (N_1921,N_1053,N_1066);
or U1922 (N_1922,N_1364,N_1404);
nand U1923 (N_1923,N_1269,N_1147);
or U1924 (N_1924,N_1241,N_1105);
nor U1925 (N_1925,N_1401,N_1039);
nor U1926 (N_1926,N_1200,N_1233);
nor U1927 (N_1927,N_1375,N_1442);
nor U1928 (N_1928,N_1417,N_1263);
nor U1929 (N_1929,N_1413,N_1124);
nand U1930 (N_1930,N_1240,N_1153);
nor U1931 (N_1931,N_1288,N_1461);
nand U1932 (N_1932,N_1207,N_1145);
nor U1933 (N_1933,N_1333,N_1241);
or U1934 (N_1934,N_1453,N_1474);
nor U1935 (N_1935,N_1055,N_1113);
nand U1936 (N_1936,N_1169,N_1108);
nor U1937 (N_1937,N_1402,N_1229);
and U1938 (N_1938,N_1306,N_1277);
or U1939 (N_1939,N_1052,N_1084);
or U1940 (N_1940,N_1159,N_1249);
nor U1941 (N_1941,N_1465,N_1149);
nor U1942 (N_1942,N_1465,N_1486);
nor U1943 (N_1943,N_1448,N_1127);
or U1944 (N_1944,N_1349,N_1494);
nor U1945 (N_1945,N_1425,N_1460);
nor U1946 (N_1946,N_1134,N_1165);
and U1947 (N_1947,N_1340,N_1067);
or U1948 (N_1948,N_1213,N_1112);
nand U1949 (N_1949,N_1096,N_1204);
or U1950 (N_1950,N_1038,N_1248);
nor U1951 (N_1951,N_1309,N_1202);
or U1952 (N_1952,N_1317,N_1481);
and U1953 (N_1953,N_1129,N_1135);
nor U1954 (N_1954,N_1270,N_1082);
and U1955 (N_1955,N_1001,N_1144);
xnor U1956 (N_1956,N_1063,N_1348);
and U1957 (N_1957,N_1027,N_1299);
and U1958 (N_1958,N_1351,N_1273);
or U1959 (N_1959,N_1192,N_1229);
nand U1960 (N_1960,N_1085,N_1284);
and U1961 (N_1961,N_1118,N_1239);
nand U1962 (N_1962,N_1472,N_1051);
and U1963 (N_1963,N_1285,N_1436);
and U1964 (N_1964,N_1475,N_1038);
nand U1965 (N_1965,N_1335,N_1059);
or U1966 (N_1966,N_1385,N_1069);
nor U1967 (N_1967,N_1432,N_1084);
or U1968 (N_1968,N_1220,N_1159);
nor U1969 (N_1969,N_1040,N_1257);
and U1970 (N_1970,N_1079,N_1369);
or U1971 (N_1971,N_1279,N_1016);
and U1972 (N_1972,N_1456,N_1278);
or U1973 (N_1973,N_1448,N_1262);
nand U1974 (N_1974,N_1357,N_1454);
nor U1975 (N_1975,N_1094,N_1442);
or U1976 (N_1976,N_1285,N_1161);
and U1977 (N_1977,N_1097,N_1061);
nand U1978 (N_1978,N_1106,N_1202);
and U1979 (N_1979,N_1227,N_1012);
nor U1980 (N_1980,N_1033,N_1421);
nor U1981 (N_1981,N_1235,N_1056);
nor U1982 (N_1982,N_1413,N_1471);
nand U1983 (N_1983,N_1294,N_1407);
nand U1984 (N_1984,N_1263,N_1367);
nor U1985 (N_1985,N_1256,N_1427);
nor U1986 (N_1986,N_1270,N_1180);
and U1987 (N_1987,N_1366,N_1404);
nand U1988 (N_1988,N_1269,N_1185);
and U1989 (N_1989,N_1338,N_1466);
nand U1990 (N_1990,N_1125,N_1337);
nor U1991 (N_1991,N_1418,N_1224);
nor U1992 (N_1992,N_1298,N_1416);
and U1993 (N_1993,N_1059,N_1146);
and U1994 (N_1994,N_1301,N_1361);
or U1995 (N_1995,N_1212,N_1003);
or U1996 (N_1996,N_1128,N_1368);
nand U1997 (N_1997,N_1181,N_1027);
or U1998 (N_1998,N_1021,N_1328);
nand U1999 (N_1999,N_1284,N_1413);
nand U2000 (N_2000,N_1678,N_1972);
nor U2001 (N_2001,N_1664,N_1910);
nand U2002 (N_2002,N_1590,N_1601);
and U2003 (N_2003,N_1801,N_1650);
nand U2004 (N_2004,N_1848,N_1988);
nor U2005 (N_2005,N_1660,N_1874);
or U2006 (N_2006,N_1662,N_1798);
or U2007 (N_2007,N_1782,N_1805);
nor U2008 (N_2008,N_1938,N_1973);
or U2009 (N_2009,N_1605,N_1920);
or U2010 (N_2010,N_1923,N_1517);
and U2011 (N_2011,N_1976,N_1783);
and U2012 (N_2012,N_1636,N_1842);
or U2013 (N_2013,N_1975,N_1510);
nand U2014 (N_2014,N_1970,N_1692);
or U2015 (N_2015,N_1600,N_1685);
nor U2016 (N_2016,N_1868,N_1697);
nor U2017 (N_2017,N_1931,N_1950);
nand U2018 (N_2018,N_1911,N_1827);
nor U2019 (N_2019,N_1968,N_1707);
and U2020 (N_2020,N_1696,N_1775);
nor U2021 (N_2021,N_1732,N_1574);
xor U2022 (N_2022,N_1759,N_1500);
or U2023 (N_2023,N_1723,N_1623);
and U2024 (N_2024,N_1965,N_1901);
and U2025 (N_2025,N_1992,N_1736);
and U2026 (N_2026,N_1584,N_1611);
nand U2027 (N_2027,N_1888,N_1958);
nand U2028 (N_2028,N_1734,N_1733);
or U2029 (N_2029,N_1808,N_1825);
nand U2030 (N_2030,N_1716,N_1849);
nand U2031 (N_2031,N_1959,N_1755);
and U2032 (N_2032,N_1655,N_1595);
nand U2033 (N_2033,N_1690,N_1737);
or U2034 (N_2034,N_1724,N_1719);
and U2035 (N_2035,N_1699,N_1828);
or U2036 (N_2036,N_1781,N_1772);
or U2037 (N_2037,N_1961,N_1875);
nand U2038 (N_2038,N_1843,N_1916);
and U2039 (N_2039,N_1822,N_1837);
and U2040 (N_2040,N_1657,N_1903);
and U2041 (N_2041,N_1613,N_1794);
nand U2042 (N_2042,N_1960,N_1521);
and U2043 (N_2043,N_1899,N_1908);
or U2044 (N_2044,N_1966,N_1514);
nand U2045 (N_2045,N_1628,N_1952);
or U2046 (N_2046,N_1990,N_1974);
and U2047 (N_2047,N_1639,N_1895);
nor U2048 (N_2048,N_1766,N_1602);
and U2049 (N_2049,N_1744,N_1516);
or U2050 (N_2050,N_1693,N_1620);
nand U2051 (N_2051,N_1980,N_1909);
nor U2052 (N_2052,N_1534,N_1860);
or U2053 (N_2053,N_1728,N_1541);
or U2054 (N_2054,N_1940,N_1807);
or U2055 (N_2055,N_1756,N_1934);
and U2056 (N_2056,N_1897,N_1760);
or U2057 (N_2057,N_1654,N_1629);
nor U2058 (N_2058,N_1730,N_1845);
nand U2059 (N_2059,N_1924,N_1904);
nor U2060 (N_2060,N_1597,N_1945);
and U2061 (N_2061,N_1815,N_1859);
nor U2062 (N_2062,N_1640,N_1870);
or U2063 (N_2063,N_1604,N_1544);
nor U2064 (N_2064,N_1993,N_1906);
and U2065 (N_2065,N_1869,N_1864);
nor U2066 (N_2066,N_1679,N_1813);
and U2067 (N_2067,N_1610,N_1577);
and U2068 (N_2068,N_1700,N_1761);
or U2069 (N_2069,N_1506,N_1619);
xor U2070 (N_2070,N_1853,N_1771);
nand U2071 (N_2071,N_1711,N_1880);
nand U2072 (N_2072,N_1762,N_1505);
nor U2073 (N_2073,N_1790,N_1740);
and U2074 (N_2074,N_1545,N_1648);
nor U2075 (N_2075,N_1515,N_1520);
nor U2076 (N_2076,N_1578,N_1582);
or U2077 (N_2077,N_1836,N_1932);
nor U2078 (N_2078,N_1527,N_1511);
nor U2079 (N_2079,N_1686,N_1663);
nor U2080 (N_2080,N_1995,N_1658);
and U2081 (N_2081,N_1676,N_1502);
and U2082 (N_2082,N_1778,N_1508);
nor U2083 (N_2083,N_1525,N_1913);
and U2084 (N_2084,N_1552,N_1675);
or U2085 (N_2085,N_1557,N_1575);
and U2086 (N_2086,N_1503,N_1963);
or U2087 (N_2087,N_1780,N_1666);
xor U2088 (N_2088,N_1512,N_1930);
nor U2089 (N_2089,N_1643,N_1674);
or U2090 (N_2090,N_1991,N_1537);
and U2091 (N_2091,N_1936,N_1572);
nand U2092 (N_2092,N_1935,N_1592);
and U2093 (N_2093,N_1768,N_1814);
nor U2094 (N_2094,N_1765,N_1809);
nor U2095 (N_2095,N_1524,N_1543);
and U2096 (N_2096,N_1540,N_1562);
and U2097 (N_2097,N_1598,N_1915);
or U2098 (N_2098,N_1641,N_1832);
nor U2099 (N_2099,N_1615,N_1871);
nand U2100 (N_2100,N_1767,N_1890);
and U2101 (N_2101,N_1585,N_1501);
and U2102 (N_2102,N_1627,N_1637);
nor U2103 (N_2103,N_1855,N_1946);
or U2104 (N_2104,N_1670,N_1955);
nand U2105 (N_2105,N_1591,N_1746);
and U2106 (N_2106,N_1919,N_1564);
and U2107 (N_2107,N_1504,N_1831);
and U2108 (N_2108,N_1914,N_1884);
nand U2109 (N_2109,N_1622,N_1854);
nor U2110 (N_2110,N_1683,N_1594);
nand U2111 (N_2111,N_1519,N_1727);
nor U2112 (N_2112,N_1548,N_1721);
xnor U2113 (N_2113,N_1526,N_1824);
nor U2114 (N_2114,N_1509,N_1816);
and U2115 (N_2115,N_1586,N_1918);
nand U2116 (N_2116,N_1635,N_1891);
nand U2117 (N_2117,N_1986,N_1748);
or U2118 (N_2118,N_1747,N_1607);
and U2119 (N_2119,N_1982,N_1704);
nor U2120 (N_2120,N_1896,N_1705);
or U2121 (N_2121,N_1659,N_1580);
nand U2122 (N_2122,N_1917,N_1750);
nand U2123 (N_2123,N_1513,N_1997);
nor U2124 (N_2124,N_1887,N_1538);
or U2125 (N_2125,N_1944,N_1647);
nor U2126 (N_2126,N_1735,N_1787);
nand U2127 (N_2127,N_1715,N_1954);
and U2128 (N_2128,N_1835,N_1587);
nand U2129 (N_2129,N_1630,N_1539);
or U2130 (N_2130,N_1701,N_1989);
nand U2131 (N_2131,N_1645,N_1752);
or U2132 (N_2132,N_1712,N_1588);
or U2133 (N_2133,N_1878,N_1892);
or U2134 (N_2134,N_1925,N_1549);
nor U2135 (N_2135,N_1806,N_1729);
nor U2136 (N_2136,N_1687,N_1788);
nand U2137 (N_2137,N_1883,N_1902);
and U2138 (N_2138,N_1739,N_1862);
and U2139 (N_2139,N_1625,N_1905);
nand U2140 (N_2140,N_1844,N_1943);
and U2141 (N_2141,N_1547,N_1941);
nor U2142 (N_2142,N_1531,N_1987);
or U2143 (N_2143,N_1556,N_1947);
or U2144 (N_2144,N_1651,N_1951);
nor U2145 (N_2145,N_1634,N_1535);
nand U2146 (N_2146,N_1710,N_1872);
or U2147 (N_2147,N_1603,N_1691);
or U2148 (N_2148,N_1969,N_1881);
nor U2149 (N_2149,N_1624,N_1608);
nand U2150 (N_2150,N_1741,N_1826);
nor U2151 (N_2151,N_1698,N_1984);
nand U2152 (N_2152,N_1937,N_1742);
or U2153 (N_2153,N_1898,N_1560);
and U2154 (N_2154,N_1799,N_1665);
or U2155 (N_2155,N_1830,N_1743);
nand U2156 (N_2156,N_1720,N_1738);
nand U2157 (N_2157,N_1817,N_1565);
nand U2158 (N_2158,N_1850,N_1793);
and U2159 (N_2159,N_1764,N_1758);
nor U2160 (N_2160,N_1684,N_1847);
nor U2161 (N_2161,N_1551,N_1770);
nor U2162 (N_2162,N_1800,N_1810);
nor U2163 (N_2163,N_1818,N_1773);
nor U2164 (N_2164,N_1889,N_1861);
nor U2165 (N_2165,N_1823,N_1949);
or U2166 (N_2166,N_1718,N_1829);
or U2167 (N_2167,N_1978,N_1795);
or U2168 (N_2168,N_1867,N_1576);
or U2169 (N_2169,N_1811,N_1558);
nand U2170 (N_2170,N_1948,N_1751);
nand U2171 (N_2171,N_1614,N_1661);
and U2172 (N_2172,N_1863,N_1928);
and U2173 (N_2173,N_1929,N_1550);
and U2174 (N_2174,N_1536,N_1672);
or U2175 (N_2175,N_1618,N_1530);
and U2176 (N_2176,N_1927,N_1820);
and U2177 (N_2177,N_1695,N_1668);
and U2178 (N_2178,N_1529,N_1554);
or U2179 (N_2179,N_1553,N_1985);
nand U2180 (N_2180,N_1796,N_1523);
nor U2181 (N_2181,N_1612,N_1702);
nor U2182 (N_2182,N_1942,N_1745);
nor U2183 (N_2183,N_1865,N_1776);
xnor U2184 (N_2184,N_1900,N_1882);
or U2185 (N_2185,N_1642,N_1819);
and U2186 (N_2186,N_1769,N_1839);
and U2187 (N_2187,N_1567,N_1589);
nor U2188 (N_2188,N_1649,N_1708);
nor U2189 (N_2189,N_1840,N_1979);
nor U2190 (N_2190,N_1821,N_1703);
nand U2191 (N_2191,N_1667,N_1680);
nor U2192 (N_2192,N_1964,N_1653);
or U2193 (N_2193,N_1632,N_1555);
nand U2194 (N_2194,N_1876,N_1717);
nand U2195 (N_2195,N_1856,N_1579);
and U2196 (N_2196,N_1646,N_1573);
and U2197 (N_2197,N_1833,N_1777);
nor U2198 (N_2198,N_1857,N_1616);
nand U2199 (N_2199,N_1893,N_1784);
nor U2200 (N_2200,N_1563,N_1638);
nand U2201 (N_2201,N_1804,N_1994);
and U2202 (N_2202,N_1596,N_1812);
nor U2203 (N_2203,N_1757,N_1656);
or U2204 (N_2204,N_1977,N_1677);
nand U2205 (N_2205,N_1566,N_1689);
nand U2206 (N_2206,N_1606,N_1542);
nor U2207 (N_2207,N_1569,N_1652);
nor U2208 (N_2208,N_1709,N_1522);
and U2209 (N_2209,N_1971,N_1581);
or U2210 (N_2210,N_1852,N_1673);
and U2211 (N_2211,N_1706,N_1983);
and U2212 (N_2212,N_1731,N_1671);
nor U2213 (N_2213,N_1688,N_1921);
and U2214 (N_2214,N_1841,N_1763);
nand U2215 (N_2215,N_1803,N_1907);
nand U2216 (N_2216,N_1507,N_1912);
nand U2217 (N_2217,N_1786,N_1791);
or U2218 (N_2218,N_1571,N_1834);
nor U2219 (N_2219,N_1599,N_1533);
or U2220 (N_2220,N_1885,N_1528);
nor U2221 (N_2221,N_1518,N_1568);
nor U2222 (N_2222,N_1583,N_1996);
nor U2223 (N_2223,N_1694,N_1998);
nor U2224 (N_2224,N_1939,N_1785);
or U2225 (N_2225,N_1894,N_1779);
nor U2226 (N_2226,N_1999,N_1749);
and U2227 (N_2227,N_1532,N_1546);
or U2228 (N_2228,N_1922,N_1802);
or U2229 (N_2229,N_1570,N_1617);
and U2230 (N_2230,N_1866,N_1725);
nor U2231 (N_2231,N_1609,N_1682);
nor U2232 (N_2232,N_1726,N_1681);
or U2233 (N_2233,N_1633,N_1593);
or U2234 (N_2234,N_1851,N_1797);
and U2235 (N_2235,N_1714,N_1621);
nand U2236 (N_2236,N_1838,N_1956);
nand U2237 (N_2237,N_1774,N_1669);
or U2238 (N_2238,N_1873,N_1981);
nand U2239 (N_2239,N_1886,N_1933);
nor U2240 (N_2240,N_1754,N_1722);
xnor U2241 (N_2241,N_1957,N_1631);
or U2242 (N_2242,N_1644,N_1561);
and U2243 (N_2243,N_1846,N_1877);
and U2244 (N_2244,N_1792,N_1967);
nor U2245 (N_2245,N_1953,N_1858);
or U2246 (N_2246,N_1713,N_1879);
or U2247 (N_2247,N_1626,N_1559);
nand U2248 (N_2248,N_1926,N_1789);
or U2249 (N_2249,N_1753,N_1962);
or U2250 (N_2250,N_1930,N_1876);
or U2251 (N_2251,N_1891,N_1923);
and U2252 (N_2252,N_1852,N_1712);
and U2253 (N_2253,N_1778,N_1583);
or U2254 (N_2254,N_1955,N_1657);
nor U2255 (N_2255,N_1962,N_1667);
nor U2256 (N_2256,N_1559,N_1967);
nand U2257 (N_2257,N_1581,N_1693);
nand U2258 (N_2258,N_1557,N_1784);
nor U2259 (N_2259,N_1904,N_1948);
and U2260 (N_2260,N_1685,N_1743);
nor U2261 (N_2261,N_1961,N_1737);
nand U2262 (N_2262,N_1794,N_1565);
nor U2263 (N_2263,N_1996,N_1684);
nor U2264 (N_2264,N_1905,N_1586);
nand U2265 (N_2265,N_1622,N_1887);
and U2266 (N_2266,N_1862,N_1819);
nor U2267 (N_2267,N_1667,N_1876);
nor U2268 (N_2268,N_1519,N_1921);
or U2269 (N_2269,N_1662,N_1984);
or U2270 (N_2270,N_1873,N_1730);
or U2271 (N_2271,N_1967,N_1740);
nor U2272 (N_2272,N_1541,N_1687);
nand U2273 (N_2273,N_1984,N_1922);
or U2274 (N_2274,N_1978,N_1668);
nand U2275 (N_2275,N_1795,N_1598);
nor U2276 (N_2276,N_1828,N_1506);
nand U2277 (N_2277,N_1580,N_1978);
nor U2278 (N_2278,N_1752,N_1887);
and U2279 (N_2279,N_1938,N_1517);
nor U2280 (N_2280,N_1525,N_1631);
and U2281 (N_2281,N_1752,N_1824);
nand U2282 (N_2282,N_1809,N_1909);
or U2283 (N_2283,N_1782,N_1955);
nand U2284 (N_2284,N_1725,N_1995);
and U2285 (N_2285,N_1932,N_1761);
nand U2286 (N_2286,N_1958,N_1733);
nor U2287 (N_2287,N_1715,N_1880);
or U2288 (N_2288,N_1813,N_1896);
nor U2289 (N_2289,N_1523,N_1804);
nor U2290 (N_2290,N_1848,N_1776);
and U2291 (N_2291,N_1658,N_1789);
nand U2292 (N_2292,N_1547,N_1847);
nand U2293 (N_2293,N_1614,N_1586);
nand U2294 (N_2294,N_1556,N_1638);
and U2295 (N_2295,N_1625,N_1572);
or U2296 (N_2296,N_1589,N_1744);
or U2297 (N_2297,N_1642,N_1793);
nand U2298 (N_2298,N_1970,N_1863);
nor U2299 (N_2299,N_1908,N_1516);
nor U2300 (N_2300,N_1986,N_1535);
nor U2301 (N_2301,N_1732,N_1979);
and U2302 (N_2302,N_1953,N_1817);
and U2303 (N_2303,N_1866,N_1814);
nand U2304 (N_2304,N_1692,N_1539);
and U2305 (N_2305,N_1727,N_1956);
and U2306 (N_2306,N_1785,N_1962);
nor U2307 (N_2307,N_1517,N_1646);
and U2308 (N_2308,N_1666,N_1591);
and U2309 (N_2309,N_1844,N_1669);
nand U2310 (N_2310,N_1503,N_1756);
or U2311 (N_2311,N_1991,N_1533);
or U2312 (N_2312,N_1549,N_1614);
and U2313 (N_2313,N_1792,N_1904);
nand U2314 (N_2314,N_1837,N_1612);
or U2315 (N_2315,N_1814,N_1570);
and U2316 (N_2316,N_1621,N_1746);
and U2317 (N_2317,N_1694,N_1855);
nand U2318 (N_2318,N_1947,N_1637);
or U2319 (N_2319,N_1690,N_1770);
nor U2320 (N_2320,N_1962,N_1937);
nor U2321 (N_2321,N_1529,N_1634);
or U2322 (N_2322,N_1904,N_1968);
nor U2323 (N_2323,N_1522,N_1610);
nand U2324 (N_2324,N_1949,N_1974);
nor U2325 (N_2325,N_1608,N_1848);
nand U2326 (N_2326,N_1685,N_1520);
nand U2327 (N_2327,N_1740,N_1757);
nand U2328 (N_2328,N_1851,N_1941);
nand U2329 (N_2329,N_1617,N_1881);
nand U2330 (N_2330,N_1897,N_1949);
xor U2331 (N_2331,N_1985,N_1761);
nor U2332 (N_2332,N_1877,N_1990);
nor U2333 (N_2333,N_1773,N_1634);
nor U2334 (N_2334,N_1889,N_1857);
and U2335 (N_2335,N_1674,N_1807);
and U2336 (N_2336,N_1906,N_1695);
and U2337 (N_2337,N_1810,N_1909);
nand U2338 (N_2338,N_1935,N_1954);
nand U2339 (N_2339,N_1691,N_1557);
and U2340 (N_2340,N_1784,N_1952);
or U2341 (N_2341,N_1885,N_1818);
and U2342 (N_2342,N_1719,N_1549);
or U2343 (N_2343,N_1557,N_1747);
or U2344 (N_2344,N_1785,N_1617);
nand U2345 (N_2345,N_1979,N_1528);
and U2346 (N_2346,N_1589,N_1551);
nand U2347 (N_2347,N_1646,N_1524);
nor U2348 (N_2348,N_1740,N_1501);
nand U2349 (N_2349,N_1605,N_1981);
nor U2350 (N_2350,N_1878,N_1547);
nor U2351 (N_2351,N_1960,N_1552);
nor U2352 (N_2352,N_1657,N_1675);
nand U2353 (N_2353,N_1856,N_1778);
xnor U2354 (N_2354,N_1937,N_1823);
or U2355 (N_2355,N_1595,N_1560);
nor U2356 (N_2356,N_1970,N_1545);
nand U2357 (N_2357,N_1925,N_1895);
nand U2358 (N_2358,N_1861,N_1893);
nor U2359 (N_2359,N_1647,N_1770);
nor U2360 (N_2360,N_1628,N_1755);
nand U2361 (N_2361,N_1583,N_1517);
and U2362 (N_2362,N_1774,N_1687);
nor U2363 (N_2363,N_1895,N_1821);
and U2364 (N_2364,N_1782,N_1708);
or U2365 (N_2365,N_1905,N_1902);
nand U2366 (N_2366,N_1913,N_1579);
nor U2367 (N_2367,N_1888,N_1727);
and U2368 (N_2368,N_1893,N_1630);
nor U2369 (N_2369,N_1638,N_1698);
nor U2370 (N_2370,N_1515,N_1609);
nand U2371 (N_2371,N_1676,N_1827);
and U2372 (N_2372,N_1993,N_1572);
and U2373 (N_2373,N_1944,N_1570);
and U2374 (N_2374,N_1657,N_1909);
nand U2375 (N_2375,N_1723,N_1547);
and U2376 (N_2376,N_1908,N_1789);
and U2377 (N_2377,N_1685,N_1938);
or U2378 (N_2378,N_1900,N_1973);
nand U2379 (N_2379,N_1855,N_1538);
nand U2380 (N_2380,N_1633,N_1728);
nand U2381 (N_2381,N_1737,N_1787);
nor U2382 (N_2382,N_1897,N_1951);
nand U2383 (N_2383,N_1729,N_1709);
and U2384 (N_2384,N_1882,N_1997);
nand U2385 (N_2385,N_1565,N_1601);
nor U2386 (N_2386,N_1923,N_1854);
nand U2387 (N_2387,N_1696,N_1786);
nand U2388 (N_2388,N_1543,N_1975);
and U2389 (N_2389,N_1571,N_1579);
nand U2390 (N_2390,N_1847,N_1505);
nor U2391 (N_2391,N_1974,N_1954);
or U2392 (N_2392,N_1599,N_1559);
xnor U2393 (N_2393,N_1683,N_1695);
nand U2394 (N_2394,N_1885,N_1581);
nor U2395 (N_2395,N_1565,N_1907);
or U2396 (N_2396,N_1702,N_1897);
and U2397 (N_2397,N_1643,N_1925);
and U2398 (N_2398,N_1680,N_1616);
nor U2399 (N_2399,N_1976,N_1768);
nand U2400 (N_2400,N_1767,N_1617);
nand U2401 (N_2401,N_1701,N_1536);
and U2402 (N_2402,N_1774,N_1570);
or U2403 (N_2403,N_1609,N_1966);
nand U2404 (N_2404,N_1696,N_1564);
nand U2405 (N_2405,N_1679,N_1885);
or U2406 (N_2406,N_1548,N_1664);
or U2407 (N_2407,N_1765,N_1923);
or U2408 (N_2408,N_1795,N_1526);
and U2409 (N_2409,N_1786,N_1742);
or U2410 (N_2410,N_1787,N_1664);
and U2411 (N_2411,N_1817,N_1797);
nor U2412 (N_2412,N_1993,N_1968);
or U2413 (N_2413,N_1820,N_1883);
and U2414 (N_2414,N_1969,N_1553);
or U2415 (N_2415,N_1570,N_1521);
and U2416 (N_2416,N_1613,N_1870);
nor U2417 (N_2417,N_1639,N_1968);
and U2418 (N_2418,N_1924,N_1759);
nand U2419 (N_2419,N_1512,N_1665);
nor U2420 (N_2420,N_1871,N_1701);
or U2421 (N_2421,N_1923,N_1825);
and U2422 (N_2422,N_1885,N_1523);
nor U2423 (N_2423,N_1567,N_1699);
or U2424 (N_2424,N_1939,N_1509);
and U2425 (N_2425,N_1647,N_1606);
and U2426 (N_2426,N_1699,N_1571);
nand U2427 (N_2427,N_1575,N_1581);
or U2428 (N_2428,N_1882,N_1748);
nor U2429 (N_2429,N_1944,N_1936);
and U2430 (N_2430,N_1676,N_1765);
nand U2431 (N_2431,N_1918,N_1646);
nand U2432 (N_2432,N_1887,N_1883);
or U2433 (N_2433,N_1985,N_1830);
nand U2434 (N_2434,N_1807,N_1723);
and U2435 (N_2435,N_1834,N_1580);
or U2436 (N_2436,N_1600,N_1502);
or U2437 (N_2437,N_1694,N_1612);
nor U2438 (N_2438,N_1571,N_1609);
or U2439 (N_2439,N_1612,N_1679);
and U2440 (N_2440,N_1968,N_1783);
nand U2441 (N_2441,N_1897,N_1647);
or U2442 (N_2442,N_1535,N_1932);
and U2443 (N_2443,N_1542,N_1956);
nor U2444 (N_2444,N_1510,N_1820);
and U2445 (N_2445,N_1504,N_1823);
and U2446 (N_2446,N_1799,N_1606);
nor U2447 (N_2447,N_1753,N_1666);
and U2448 (N_2448,N_1840,N_1907);
or U2449 (N_2449,N_1844,N_1810);
nand U2450 (N_2450,N_1952,N_1922);
nand U2451 (N_2451,N_1720,N_1918);
nand U2452 (N_2452,N_1694,N_1621);
or U2453 (N_2453,N_1627,N_1684);
and U2454 (N_2454,N_1833,N_1746);
nor U2455 (N_2455,N_1842,N_1949);
nand U2456 (N_2456,N_1817,N_1820);
nor U2457 (N_2457,N_1721,N_1765);
nand U2458 (N_2458,N_1580,N_1796);
xor U2459 (N_2459,N_1881,N_1612);
nand U2460 (N_2460,N_1596,N_1958);
nand U2461 (N_2461,N_1938,N_1686);
nor U2462 (N_2462,N_1545,N_1949);
or U2463 (N_2463,N_1564,N_1954);
or U2464 (N_2464,N_1578,N_1601);
and U2465 (N_2465,N_1884,N_1504);
nand U2466 (N_2466,N_1609,N_1998);
nand U2467 (N_2467,N_1521,N_1852);
nand U2468 (N_2468,N_1803,N_1951);
or U2469 (N_2469,N_1679,N_1653);
nor U2470 (N_2470,N_1514,N_1670);
nand U2471 (N_2471,N_1768,N_1733);
and U2472 (N_2472,N_1509,N_1738);
nor U2473 (N_2473,N_1705,N_1634);
or U2474 (N_2474,N_1659,N_1945);
and U2475 (N_2475,N_1537,N_1561);
nand U2476 (N_2476,N_1904,N_1503);
or U2477 (N_2477,N_1657,N_1663);
and U2478 (N_2478,N_1617,N_1825);
or U2479 (N_2479,N_1851,N_1648);
or U2480 (N_2480,N_1742,N_1916);
or U2481 (N_2481,N_1669,N_1573);
nand U2482 (N_2482,N_1665,N_1949);
nor U2483 (N_2483,N_1622,N_1837);
nand U2484 (N_2484,N_1546,N_1626);
or U2485 (N_2485,N_1566,N_1862);
nand U2486 (N_2486,N_1632,N_1883);
nor U2487 (N_2487,N_1657,N_1997);
and U2488 (N_2488,N_1961,N_1675);
nand U2489 (N_2489,N_1948,N_1665);
and U2490 (N_2490,N_1743,N_1680);
or U2491 (N_2491,N_1749,N_1892);
nor U2492 (N_2492,N_1904,N_1768);
nand U2493 (N_2493,N_1514,N_1777);
and U2494 (N_2494,N_1634,N_1684);
or U2495 (N_2495,N_1612,N_1801);
or U2496 (N_2496,N_1762,N_1991);
or U2497 (N_2497,N_1766,N_1683);
and U2498 (N_2498,N_1794,N_1513);
and U2499 (N_2499,N_1684,N_1743);
nor U2500 (N_2500,N_2329,N_2241);
nor U2501 (N_2501,N_2212,N_2416);
and U2502 (N_2502,N_2346,N_2439);
nor U2503 (N_2503,N_2195,N_2214);
nand U2504 (N_2504,N_2088,N_2394);
nand U2505 (N_2505,N_2110,N_2421);
and U2506 (N_2506,N_2288,N_2203);
and U2507 (N_2507,N_2048,N_2261);
nor U2508 (N_2508,N_2138,N_2001);
xor U2509 (N_2509,N_2226,N_2101);
or U2510 (N_2510,N_2236,N_2106);
xnor U2511 (N_2511,N_2426,N_2423);
or U2512 (N_2512,N_2130,N_2472);
and U2513 (N_2513,N_2420,N_2022);
and U2514 (N_2514,N_2114,N_2386);
nor U2515 (N_2515,N_2078,N_2289);
nand U2516 (N_2516,N_2186,N_2284);
or U2517 (N_2517,N_2403,N_2321);
nand U2518 (N_2518,N_2396,N_2330);
or U2519 (N_2519,N_2123,N_2467);
nor U2520 (N_2520,N_2466,N_2100);
nor U2521 (N_2521,N_2415,N_2332);
xnor U2522 (N_2522,N_2004,N_2308);
and U2523 (N_2523,N_2343,N_2377);
nand U2524 (N_2524,N_2266,N_2198);
and U2525 (N_2525,N_2052,N_2159);
or U2526 (N_2526,N_2071,N_2497);
and U2527 (N_2527,N_2325,N_2320);
nand U2528 (N_2528,N_2199,N_2446);
and U2529 (N_2529,N_2444,N_2194);
or U2530 (N_2530,N_2188,N_2135);
and U2531 (N_2531,N_2112,N_2306);
nor U2532 (N_2532,N_2147,N_2316);
or U2533 (N_2533,N_2014,N_2040);
nand U2534 (N_2534,N_2462,N_2141);
and U2535 (N_2535,N_2249,N_2077);
and U2536 (N_2536,N_2448,N_2218);
nor U2537 (N_2537,N_2428,N_2368);
nand U2538 (N_2538,N_2271,N_2066);
and U2539 (N_2539,N_2491,N_2438);
or U2540 (N_2540,N_2006,N_2397);
nor U2541 (N_2541,N_2156,N_2276);
nand U2542 (N_2542,N_2360,N_2470);
nor U2543 (N_2543,N_2399,N_2365);
nand U2544 (N_2544,N_2378,N_2176);
nor U2545 (N_2545,N_2418,N_2221);
nand U2546 (N_2546,N_2425,N_2207);
nand U2547 (N_2547,N_2158,N_2118);
and U2548 (N_2548,N_2098,N_2084);
and U2549 (N_2549,N_2015,N_2274);
and U2550 (N_2550,N_2155,N_2489);
or U2551 (N_2551,N_2171,N_2083);
nor U2552 (N_2552,N_2046,N_2452);
nand U2553 (N_2553,N_2460,N_2073);
nand U2554 (N_2554,N_2020,N_2181);
or U2555 (N_2555,N_2055,N_2002);
or U2556 (N_2556,N_2469,N_2069);
nand U2557 (N_2557,N_2028,N_2391);
nand U2558 (N_2558,N_2179,N_2036);
xnor U2559 (N_2559,N_2382,N_2016);
nor U2560 (N_2560,N_2344,N_2104);
and U2561 (N_2561,N_2119,N_2010);
or U2562 (N_2562,N_2349,N_2409);
or U2563 (N_2563,N_2196,N_2183);
or U2564 (N_2564,N_2304,N_2301);
or U2565 (N_2565,N_2383,N_2081);
and U2566 (N_2566,N_2051,N_2362);
nor U2567 (N_2567,N_2495,N_2471);
nand U2568 (N_2568,N_2305,N_2000);
or U2569 (N_2569,N_2092,N_2201);
nor U2570 (N_2570,N_2410,N_2458);
nand U2571 (N_2571,N_2042,N_2056);
or U2572 (N_2572,N_2313,N_2085);
or U2573 (N_2573,N_2030,N_2370);
nand U2574 (N_2574,N_2142,N_2224);
nor U2575 (N_2575,N_2486,N_2461);
or U2576 (N_2576,N_2244,N_2229);
or U2577 (N_2577,N_2075,N_2427);
or U2578 (N_2578,N_2189,N_2436);
nor U2579 (N_2579,N_2499,N_2095);
or U2580 (N_2580,N_2367,N_2352);
and U2581 (N_2581,N_2024,N_2220);
nor U2582 (N_2582,N_2240,N_2404);
nand U2583 (N_2583,N_2223,N_2034);
nor U2584 (N_2584,N_2414,N_2290);
and U2585 (N_2585,N_2480,N_2453);
or U2586 (N_2586,N_2139,N_2216);
nand U2587 (N_2587,N_2395,N_2173);
nor U2588 (N_2588,N_2468,N_2167);
nand U2589 (N_2589,N_2160,N_2253);
and U2590 (N_2590,N_2113,N_2294);
nor U2591 (N_2591,N_2099,N_2231);
or U2592 (N_2592,N_2376,N_2434);
nand U2593 (N_2593,N_2031,N_2317);
nor U2594 (N_2594,N_2437,N_2451);
nor U2595 (N_2595,N_2431,N_2125);
nand U2596 (N_2596,N_2232,N_2090);
or U2597 (N_2597,N_2282,N_2197);
xor U2598 (N_2598,N_2140,N_2337);
or U2599 (N_2599,N_2345,N_2277);
and U2600 (N_2600,N_2025,N_2127);
nand U2601 (N_2601,N_2251,N_2256);
and U2602 (N_2602,N_2496,N_2222);
or U2603 (N_2603,N_2029,N_2405);
nor U2604 (N_2604,N_2273,N_2485);
or U2605 (N_2605,N_2278,N_2260);
and U2606 (N_2606,N_2279,N_2348);
and U2607 (N_2607,N_2153,N_2300);
nor U2608 (N_2608,N_2474,N_2412);
nand U2609 (N_2609,N_2061,N_2169);
nand U2610 (N_2610,N_2192,N_2390);
and U2611 (N_2611,N_2298,N_2387);
or U2612 (N_2612,N_2108,N_2219);
and U2613 (N_2613,N_2182,N_2054);
nand U2614 (N_2614,N_2137,N_2144);
nand U2615 (N_2615,N_2287,N_2215);
or U2616 (N_2616,N_2152,N_2285);
nand U2617 (N_2617,N_2441,N_2356);
nor U2618 (N_2618,N_2359,N_2413);
or U2619 (N_2619,N_2033,N_2336);
or U2620 (N_2620,N_2432,N_2177);
or U2621 (N_2621,N_2191,N_2208);
nor U2622 (N_2622,N_2262,N_2115);
nand U2623 (N_2623,N_2038,N_2205);
or U2624 (N_2624,N_2082,N_2435);
or U2625 (N_2625,N_2018,N_2105);
nor U2626 (N_2626,N_2246,N_2148);
nor U2627 (N_2627,N_2258,N_2315);
or U2628 (N_2628,N_2267,N_2059);
nand U2629 (N_2629,N_2227,N_2264);
or U2630 (N_2630,N_2184,N_2166);
nor U2631 (N_2631,N_2398,N_2419);
and U2632 (N_2632,N_2126,N_2326);
nand U2633 (N_2633,N_2488,N_2479);
nand U2634 (N_2634,N_2079,N_2017);
or U2635 (N_2635,N_2297,N_2202);
or U2636 (N_2636,N_2185,N_2333);
nand U2637 (N_2637,N_2407,N_2060);
nand U2638 (N_2638,N_2465,N_2093);
and U2639 (N_2639,N_2373,N_2323);
or U2640 (N_2640,N_2097,N_2401);
nand U2641 (N_2641,N_2286,N_2358);
and U2642 (N_2642,N_2058,N_2178);
nand U2643 (N_2643,N_2041,N_2440);
nor U2644 (N_2644,N_2136,N_2131);
and U2645 (N_2645,N_2026,N_2089);
nor U2646 (N_2646,N_2193,N_2408);
nand U2647 (N_2647,N_2483,N_2340);
or U2648 (N_2648,N_2237,N_2165);
and U2649 (N_2649,N_2094,N_2442);
or U2650 (N_2650,N_2430,N_2049);
nand U2651 (N_2651,N_2257,N_2044);
nand U2652 (N_2652,N_2389,N_2250);
nand U2653 (N_2653,N_2080,N_2353);
and U2654 (N_2654,N_2291,N_2154);
or U2655 (N_2655,N_2037,N_2456);
nor U2656 (N_2656,N_2374,N_2023);
nand U2657 (N_2657,N_2380,N_2270);
and U2658 (N_2658,N_2375,N_2209);
or U2659 (N_2659,N_2050,N_2355);
or U2660 (N_2660,N_2369,N_2454);
nor U2661 (N_2661,N_2351,N_2045);
nand U2662 (N_2662,N_2005,N_2393);
and U2663 (N_2663,N_2269,N_2180);
or U2664 (N_2664,N_2494,N_2263);
or U2665 (N_2665,N_2233,N_2213);
nor U2666 (N_2666,N_2477,N_2011);
nand U2667 (N_2667,N_2062,N_2172);
and U2668 (N_2668,N_2357,N_2457);
nor U2669 (N_2669,N_2230,N_2475);
and U2670 (N_2670,N_2281,N_2076);
or U2671 (N_2671,N_2129,N_2449);
nor U2672 (N_2672,N_2007,N_2314);
nand U2673 (N_2673,N_2206,N_2299);
nor U2674 (N_2674,N_2309,N_2347);
nand U2675 (N_2675,N_2303,N_2255);
or U2676 (N_2676,N_2200,N_2107);
xnor U2677 (N_2677,N_2243,N_2068);
or U2678 (N_2678,N_2235,N_2265);
nor U2679 (N_2679,N_2162,N_2053);
nor U2680 (N_2680,N_2292,N_2161);
nor U2681 (N_2681,N_2063,N_2381);
or U2682 (N_2682,N_2259,N_2411);
and U2683 (N_2683,N_2476,N_2319);
or U2684 (N_2684,N_2372,N_2417);
nand U2685 (N_2685,N_2027,N_2064);
or U2686 (N_2686,N_2385,N_2328);
or U2687 (N_2687,N_2311,N_2482);
or U2688 (N_2688,N_2013,N_2217);
and U2689 (N_2689,N_2091,N_2283);
and U2690 (N_2690,N_2366,N_2361);
or U2691 (N_2691,N_2254,N_2481);
nor U2692 (N_2692,N_2490,N_2111);
nand U2693 (N_2693,N_2318,N_2478);
and U2694 (N_2694,N_2032,N_2145);
nand U2695 (N_2695,N_2245,N_2388);
or U2696 (N_2696,N_2331,N_2043);
nor U2697 (N_2697,N_2295,N_2150);
or U2698 (N_2698,N_2463,N_2109);
and U2699 (N_2699,N_2302,N_2324);
nand U2700 (N_2700,N_2455,N_2164);
and U2701 (N_2701,N_2341,N_2335);
or U2702 (N_2702,N_2350,N_2307);
nand U2703 (N_2703,N_2190,N_2143);
nor U2704 (N_2704,N_2146,N_2424);
nand U2705 (N_2705,N_2087,N_2492);
or U2706 (N_2706,N_2204,N_2242);
and U2707 (N_2707,N_2248,N_2354);
xnor U2708 (N_2708,N_2234,N_2252);
nand U2709 (N_2709,N_2116,N_2012);
and U2710 (N_2710,N_2065,N_2211);
and U2711 (N_2711,N_2338,N_2121);
and U2712 (N_2712,N_2443,N_2117);
nor U2713 (N_2713,N_2447,N_2272);
or U2714 (N_2714,N_2379,N_2371);
or U2715 (N_2715,N_2310,N_2384);
nor U2716 (N_2716,N_2035,N_2429);
or U2717 (N_2717,N_2296,N_2074);
and U2718 (N_2718,N_2342,N_2120);
and U2719 (N_2719,N_2280,N_2149);
and U2720 (N_2720,N_2473,N_2008);
nor U2721 (N_2721,N_2067,N_2493);
nor U2722 (N_2722,N_2163,N_2210);
nor U2723 (N_2723,N_2487,N_2433);
and U2724 (N_2724,N_2021,N_2392);
nand U2725 (N_2725,N_2247,N_2039);
or U2726 (N_2726,N_2459,N_2239);
or U2727 (N_2727,N_2134,N_2057);
nor U2728 (N_2728,N_2122,N_2187);
or U2729 (N_2729,N_2327,N_2406);
and U2730 (N_2730,N_2124,N_2103);
nor U2731 (N_2731,N_2498,N_2096);
or U2732 (N_2732,N_2072,N_2275);
and U2733 (N_2733,N_2019,N_2445);
nor U2734 (N_2734,N_2225,N_2450);
or U2735 (N_2735,N_2402,N_2132);
nor U2736 (N_2736,N_2268,N_2228);
or U2737 (N_2737,N_2174,N_2364);
nand U2738 (N_2738,N_2157,N_2400);
nor U2739 (N_2739,N_2047,N_2086);
nand U2740 (N_2740,N_2151,N_2312);
nand U2741 (N_2741,N_2363,N_2168);
and U2742 (N_2742,N_2293,N_2003);
and U2743 (N_2743,N_2322,N_2339);
and U2744 (N_2744,N_2102,N_2334);
or U2745 (N_2745,N_2128,N_2070);
nand U2746 (N_2746,N_2238,N_2133);
and U2747 (N_2747,N_2484,N_2422);
nor U2748 (N_2748,N_2009,N_2170);
nand U2749 (N_2749,N_2464,N_2175);
nand U2750 (N_2750,N_2079,N_2472);
or U2751 (N_2751,N_2004,N_2186);
and U2752 (N_2752,N_2135,N_2354);
or U2753 (N_2753,N_2191,N_2448);
nor U2754 (N_2754,N_2249,N_2041);
and U2755 (N_2755,N_2136,N_2303);
nand U2756 (N_2756,N_2314,N_2431);
and U2757 (N_2757,N_2080,N_2337);
nor U2758 (N_2758,N_2075,N_2341);
nand U2759 (N_2759,N_2300,N_2173);
nor U2760 (N_2760,N_2233,N_2195);
nor U2761 (N_2761,N_2226,N_2319);
or U2762 (N_2762,N_2041,N_2139);
and U2763 (N_2763,N_2042,N_2450);
nor U2764 (N_2764,N_2205,N_2218);
nand U2765 (N_2765,N_2376,N_2290);
and U2766 (N_2766,N_2036,N_2045);
nor U2767 (N_2767,N_2297,N_2162);
nand U2768 (N_2768,N_2174,N_2011);
and U2769 (N_2769,N_2299,N_2440);
nor U2770 (N_2770,N_2471,N_2059);
nand U2771 (N_2771,N_2268,N_2235);
and U2772 (N_2772,N_2016,N_2034);
nor U2773 (N_2773,N_2364,N_2458);
and U2774 (N_2774,N_2311,N_2261);
and U2775 (N_2775,N_2162,N_2124);
or U2776 (N_2776,N_2180,N_2188);
and U2777 (N_2777,N_2187,N_2127);
and U2778 (N_2778,N_2116,N_2263);
or U2779 (N_2779,N_2411,N_2393);
nand U2780 (N_2780,N_2124,N_2028);
or U2781 (N_2781,N_2219,N_2160);
nand U2782 (N_2782,N_2132,N_2343);
nor U2783 (N_2783,N_2250,N_2008);
nand U2784 (N_2784,N_2063,N_2035);
nand U2785 (N_2785,N_2041,N_2050);
and U2786 (N_2786,N_2299,N_2106);
nand U2787 (N_2787,N_2343,N_2401);
nor U2788 (N_2788,N_2088,N_2377);
and U2789 (N_2789,N_2008,N_2132);
nand U2790 (N_2790,N_2135,N_2189);
or U2791 (N_2791,N_2005,N_2197);
or U2792 (N_2792,N_2441,N_2345);
nor U2793 (N_2793,N_2242,N_2004);
nor U2794 (N_2794,N_2422,N_2168);
and U2795 (N_2795,N_2478,N_2403);
nand U2796 (N_2796,N_2488,N_2067);
or U2797 (N_2797,N_2350,N_2195);
nor U2798 (N_2798,N_2211,N_2099);
nor U2799 (N_2799,N_2210,N_2179);
or U2800 (N_2800,N_2440,N_2129);
nand U2801 (N_2801,N_2452,N_2474);
nand U2802 (N_2802,N_2476,N_2279);
or U2803 (N_2803,N_2050,N_2415);
nor U2804 (N_2804,N_2085,N_2253);
or U2805 (N_2805,N_2047,N_2331);
nand U2806 (N_2806,N_2485,N_2020);
nor U2807 (N_2807,N_2044,N_2006);
nand U2808 (N_2808,N_2283,N_2075);
and U2809 (N_2809,N_2291,N_2149);
and U2810 (N_2810,N_2391,N_2327);
and U2811 (N_2811,N_2301,N_2424);
or U2812 (N_2812,N_2366,N_2323);
nor U2813 (N_2813,N_2057,N_2163);
or U2814 (N_2814,N_2313,N_2253);
or U2815 (N_2815,N_2318,N_2388);
or U2816 (N_2816,N_2399,N_2253);
or U2817 (N_2817,N_2215,N_2114);
and U2818 (N_2818,N_2073,N_2385);
and U2819 (N_2819,N_2412,N_2036);
and U2820 (N_2820,N_2185,N_2419);
nand U2821 (N_2821,N_2473,N_2347);
nor U2822 (N_2822,N_2338,N_2149);
nor U2823 (N_2823,N_2471,N_2079);
or U2824 (N_2824,N_2146,N_2133);
and U2825 (N_2825,N_2181,N_2329);
and U2826 (N_2826,N_2161,N_2029);
and U2827 (N_2827,N_2441,N_2338);
nor U2828 (N_2828,N_2467,N_2097);
nand U2829 (N_2829,N_2424,N_2447);
or U2830 (N_2830,N_2186,N_2417);
nand U2831 (N_2831,N_2350,N_2391);
or U2832 (N_2832,N_2385,N_2197);
nor U2833 (N_2833,N_2190,N_2052);
nor U2834 (N_2834,N_2288,N_2117);
and U2835 (N_2835,N_2440,N_2145);
or U2836 (N_2836,N_2261,N_2184);
or U2837 (N_2837,N_2182,N_2193);
or U2838 (N_2838,N_2235,N_2369);
nand U2839 (N_2839,N_2184,N_2027);
and U2840 (N_2840,N_2230,N_2322);
and U2841 (N_2841,N_2042,N_2118);
nand U2842 (N_2842,N_2066,N_2138);
nand U2843 (N_2843,N_2018,N_2171);
nor U2844 (N_2844,N_2065,N_2054);
nor U2845 (N_2845,N_2039,N_2456);
or U2846 (N_2846,N_2318,N_2229);
xnor U2847 (N_2847,N_2455,N_2383);
nand U2848 (N_2848,N_2104,N_2385);
nor U2849 (N_2849,N_2356,N_2185);
or U2850 (N_2850,N_2228,N_2316);
nand U2851 (N_2851,N_2055,N_2067);
nand U2852 (N_2852,N_2499,N_2115);
and U2853 (N_2853,N_2226,N_2305);
or U2854 (N_2854,N_2345,N_2092);
and U2855 (N_2855,N_2070,N_2158);
and U2856 (N_2856,N_2278,N_2478);
and U2857 (N_2857,N_2393,N_2001);
and U2858 (N_2858,N_2391,N_2013);
nand U2859 (N_2859,N_2439,N_2185);
and U2860 (N_2860,N_2151,N_2318);
and U2861 (N_2861,N_2070,N_2053);
or U2862 (N_2862,N_2433,N_2326);
and U2863 (N_2863,N_2078,N_2002);
and U2864 (N_2864,N_2176,N_2055);
and U2865 (N_2865,N_2411,N_2324);
and U2866 (N_2866,N_2276,N_2077);
nand U2867 (N_2867,N_2378,N_2124);
or U2868 (N_2868,N_2372,N_2116);
nor U2869 (N_2869,N_2390,N_2256);
and U2870 (N_2870,N_2490,N_2084);
or U2871 (N_2871,N_2336,N_2365);
nand U2872 (N_2872,N_2173,N_2432);
or U2873 (N_2873,N_2309,N_2090);
or U2874 (N_2874,N_2279,N_2179);
and U2875 (N_2875,N_2354,N_2385);
nand U2876 (N_2876,N_2326,N_2068);
and U2877 (N_2877,N_2428,N_2306);
or U2878 (N_2878,N_2012,N_2337);
or U2879 (N_2879,N_2127,N_2288);
nand U2880 (N_2880,N_2026,N_2020);
nor U2881 (N_2881,N_2221,N_2252);
nand U2882 (N_2882,N_2183,N_2273);
nand U2883 (N_2883,N_2418,N_2045);
nand U2884 (N_2884,N_2234,N_2225);
and U2885 (N_2885,N_2115,N_2051);
and U2886 (N_2886,N_2199,N_2250);
nand U2887 (N_2887,N_2472,N_2289);
or U2888 (N_2888,N_2146,N_2409);
and U2889 (N_2889,N_2040,N_2298);
or U2890 (N_2890,N_2191,N_2279);
nor U2891 (N_2891,N_2197,N_2408);
nand U2892 (N_2892,N_2486,N_2135);
nor U2893 (N_2893,N_2210,N_2111);
and U2894 (N_2894,N_2268,N_2269);
and U2895 (N_2895,N_2190,N_2268);
nand U2896 (N_2896,N_2144,N_2088);
nand U2897 (N_2897,N_2030,N_2023);
or U2898 (N_2898,N_2441,N_2296);
and U2899 (N_2899,N_2140,N_2210);
or U2900 (N_2900,N_2409,N_2071);
and U2901 (N_2901,N_2192,N_2490);
nor U2902 (N_2902,N_2062,N_2196);
xnor U2903 (N_2903,N_2023,N_2432);
and U2904 (N_2904,N_2228,N_2073);
nand U2905 (N_2905,N_2438,N_2062);
nor U2906 (N_2906,N_2032,N_2319);
or U2907 (N_2907,N_2282,N_2259);
or U2908 (N_2908,N_2119,N_2295);
or U2909 (N_2909,N_2098,N_2143);
or U2910 (N_2910,N_2024,N_2456);
nor U2911 (N_2911,N_2335,N_2467);
and U2912 (N_2912,N_2094,N_2234);
and U2913 (N_2913,N_2476,N_2222);
and U2914 (N_2914,N_2336,N_2260);
and U2915 (N_2915,N_2441,N_2119);
and U2916 (N_2916,N_2086,N_2319);
nor U2917 (N_2917,N_2151,N_2280);
nand U2918 (N_2918,N_2204,N_2220);
nand U2919 (N_2919,N_2389,N_2326);
or U2920 (N_2920,N_2340,N_2361);
or U2921 (N_2921,N_2454,N_2355);
xor U2922 (N_2922,N_2259,N_2402);
nand U2923 (N_2923,N_2380,N_2231);
nand U2924 (N_2924,N_2196,N_2359);
or U2925 (N_2925,N_2232,N_2100);
nand U2926 (N_2926,N_2279,N_2148);
nor U2927 (N_2927,N_2356,N_2384);
and U2928 (N_2928,N_2022,N_2125);
or U2929 (N_2929,N_2304,N_2058);
nand U2930 (N_2930,N_2256,N_2078);
and U2931 (N_2931,N_2170,N_2428);
nor U2932 (N_2932,N_2064,N_2399);
and U2933 (N_2933,N_2312,N_2364);
nand U2934 (N_2934,N_2325,N_2152);
or U2935 (N_2935,N_2294,N_2209);
or U2936 (N_2936,N_2458,N_2237);
or U2937 (N_2937,N_2356,N_2165);
nand U2938 (N_2938,N_2377,N_2304);
or U2939 (N_2939,N_2064,N_2107);
and U2940 (N_2940,N_2319,N_2449);
or U2941 (N_2941,N_2212,N_2417);
and U2942 (N_2942,N_2475,N_2301);
and U2943 (N_2943,N_2187,N_2267);
nor U2944 (N_2944,N_2354,N_2420);
nor U2945 (N_2945,N_2181,N_2141);
and U2946 (N_2946,N_2302,N_2322);
or U2947 (N_2947,N_2233,N_2284);
and U2948 (N_2948,N_2422,N_2393);
and U2949 (N_2949,N_2102,N_2379);
nor U2950 (N_2950,N_2407,N_2036);
nor U2951 (N_2951,N_2232,N_2305);
and U2952 (N_2952,N_2363,N_2396);
or U2953 (N_2953,N_2234,N_2358);
nor U2954 (N_2954,N_2457,N_2348);
and U2955 (N_2955,N_2307,N_2484);
nor U2956 (N_2956,N_2456,N_2076);
nand U2957 (N_2957,N_2091,N_2437);
and U2958 (N_2958,N_2299,N_2131);
and U2959 (N_2959,N_2434,N_2287);
nor U2960 (N_2960,N_2318,N_2205);
or U2961 (N_2961,N_2091,N_2409);
and U2962 (N_2962,N_2360,N_2142);
or U2963 (N_2963,N_2408,N_2380);
and U2964 (N_2964,N_2142,N_2398);
or U2965 (N_2965,N_2192,N_2107);
and U2966 (N_2966,N_2197,N_2353);
or U2967 (N_2967,N_2106,N_2069);
nand U2968 (N_2968,N_2284,N_2315);
nand U2969 (N_2969,N_2336,N_2011);
or U2970 (N_2970,N_2470,N_2422);
nand U2971 (N_2971,N_2157,N_2374);
nor U2972 (N_2972,N_2017,N_2313);
nand U2973 (N_2973,N_2203,N_2312);
nand U2974 (N_2974,N_2434,N_2113);
or U2975 (N_2975,N_2186,N_2225);
nand U2976 (N_2976,N_2162,N_2385);
and U2977 (N_2977,N_2485,N_2122);
nor U2978 (N_2978,N_2377,N_2059);
nor U2979 (N_2979,N_2161,N_2250);
nand U2980 (N_2980,N_2070,N_2279);
and U2981 (N_2981,N_2366,N_2117);
and U2982 (N_2982,N_2089,N_2127);
nand U2983 (N_2983,N_2145,N_2033);
and U2984 (N_2984,N_2485,N_2079);
nor U2985 (N_2985,N_2373,N_2314);
nor U2986 (N_2986,N_2144,N_2107);
nand U2987 (N_2987,N_2444,N_2288);
and U2988 (N_2988,N_2056,N_2093);
or U2989 (N_2989,N_2364,N_2134);
or U2990 (N_2990,N_2385,N_2467);
and U2991 (N_2991,N_2129,N_2058);
or U2992 (N_2992,N_2087,N_2231);
or U2993 (N_2993,N_2304,N_2203);
nor U2994 (N_2994,N_2143,N_2019);
nor U2995 (N_2995,N_2331,N_2305);
or U2996 (N_2996,N_2219,N_2204);
nor U2997 (N_2997,N_2106,N_2470);
nand U2998 (N_2998,N_2267,N_2304);
nand U2999 (N_2999,N_2339,N_2344);
xor U3000 (N_3000,N_2539,N_2879);
nand U3001 (N_3001,N_2929,N_2795);
and U3002 (N_3002,N_2503,N_2570);
or U3003 (N_3003,N_2722,N_2869);
nand U3004 (N_3004,N_2985,N_2699);
nor U3005 (N_3005,N_2797,N_2993);
nand U3006 (N_3006,N_2639,N_2673);
nand U3007 (N_3007,N_2670,N_2995);
nand U3008 (N_3008,N_2712,N_2893);
nand U3009 (N_3009,N_2744,N_2844);
and U3010 (N_3010,N_2927,N_2936);
or U3011 (N_3011,N_2693,N_2585);
and U3012 (N_3012,N_2692,N_2983);
and U3013 (N_3013,N_2717,N_2875);
nand U3014 (N_3014,N_2773,N_2600);
nor U3015 (N_3015,N_2841,N_2633);
nand U3016 (N_3016,N_2534,N_2680);
or U3017 (N_3017,N_2897,N_2914);
xnor U3018 (N_3018,N_2952,N_2713);
nand U3019 (N_3019,N_2855,N_2672);
or U3020 (N_3020,N_2548,N_2991);
or U3021 (N_3021,N_2973,N_2965);
nor U3022 (N_3022,N_2777,N_2596);
nor U3023 (N_3023,N_2880,N_2960);
and U3024 (N_3024,N_2850,N_2611);
or U3025 (N_3025,N_2813,N_2878);
nand U3026 (N_3026,N_2975,N_2566);
nand U3027 (N_3027,N_2872,N_2899);
and U3028 (N_3028,N_2522,N_2691);
or U3029 (N_3029,N_2725,N_2829);
or U3030 (N_3030,N_2848,N_2513);
nor U3031 (N_3031,N_2967,N_2906);
nor U3032 (N_3032,N_2714,N_2977);
or U3033 (N_3033,N_2516,N_2601);
nand U3034 (N_3034,N_2833,N_2506);
or U3035 (N_3035,N_2599,N_2959);
or U3036 (N_3036,N_2902,N_2963);
nand U3037 (N_3037,N_2593,N_2726);
or U3038 (N_3038,N_2598,N_2812);
or U3039 (N_3039,N_2700,N_2647);
or U3040 (N_3040,N_2877,N_2703);
nand U3041 (N_3041,N_2937,N_2617);
nand U3042 (N_3042,N_2823,N_2769);
and U3043 (N_3043,N_2885,N_2940);
or U3044 (N_3044,N_2618,N_2884);
or U3045 (N_3045,N_2948,N_2849);
or U3046 (N_3046,N_2501,N_2721);
nor U3047 (N_3047,N_2631,N_2547);
or U3048 (N_3048,N_2730,N_2775);
or U3049 (N_3049,N_2792,N_2799);
nand U3050 (N_3050,N_2562,N_2784);
and U3051 (N_3051,N_2565,N_2741);
nor U3052 (N_3052,N_2542,N_2742);
and U3053 (N_3053,N_2745,N_2904);
or U3054 (N_3054,N_2577,N_2519);
and U3055 (N_3055,N_2932,N_2698);
or U3056 (N_3056,N_2626,N_2851);
nand U3057 (N_3057,N_2881,N_2671);
nor U3058 (N_3058,N_2933,N_2729);
nor U3059 (N_3059,N_2966,N_2941);
nand U3060 (N_3060,N_2718,N_2727);
nand U3061 (N_3061,N_2916,N_2835);
nor U3062 (N_3062,N_2989,N_2651);
and U3063 (N_3063,N_2980,N_2590);
and U3064 (N_3064,N_2676,N_2808);
or U3065 (N_3065,N_2694,N_2768);
nor U3066 (N_3066,N_2576,N_2535);
nand U3067 (N_3067,N_2707,N_2649);
or U3068 (N_3068,N_2752,N_2706);
or U3069 (N_3069,N_2669,N_2947);
nor U3070 (N_3070,N_2802,N_2635);
and U3071 (N_3071,N_2859,N_2822);
and U3072 (N_3072,N_2763,N_2650);
and U3073 (N_3073,N_2734,N_2976);
or U3074 (N_3074,N_2951,N_2846);
or U3075 (N_3075,N_2688,N_2824);
or U3076 (N_3076,N_2986,N_2908);
nand U3077 (N_3077,N_2946,N_2922);
or U3078 (N_3078,N_2774,N_2826);
and U3079 (N_3079,N_2756,N_2935);
or U3080 (N_3080,N_2701,N_2815);
nor U3081 (N_3081,N_2820,N_2955);
nand U3082 (N_3082,N_2876,N_2587);
nor U3083 (N_3083,N_2981,N_2594);
or U3084 (N_3084,N_2719,N_2920);
and U3085 (N_3085,N_2665,N_2549);
and U3086 (N_3086,N_2733,N_2910);
nor U3087 (N_3087,N_2818,N_2541);
and U3088 (N_3088,N_2751,N_2934);
or U3089 (N_3089,N_2810,N_2771);
or U3090 (N_3090,N_2529,N_2648);
nor U3091 (N_3091,N_2919,N_2766);
or U3092 (N_3092,N_2526,N_2903);
or U3093 (N_3093,N_2761,N_2753);
or U3094 (N_3094,N_2954,N_2858);
nand U3095 (N_3095,N_2504,N_2999);
nor U3096 (N_3096,N_2540,N_2597);
or U3097 (N_3097,N_2837,N_2956);
and U3098 (N_3098,N_2962,N_2575);
xor U3099 (N_3099,N_2931,N_2873);
nand U3100 (N_3100,N_2731,N_2687);
and U3101 (N_3101,N_2732,N_2621);
nor U3102 (N_3102,N_2690,N_2682);
nand U3103 (N_3103,N_2634,N_2895);
or U3104 (N_3104,N_2524,N_2567);
nor U3105 (N_3105,N_2588,N_2632);
or U3106 (N_3106,N_2595,N_2654);
xor U3107 (N_3107,N_2883,N_2847);
nor U3108 (N_3108,N_2968,N_2961);
and U3109 (N_3109,N_2544,N_2842);
nor U3110 (N_3110,N_2620,N_2554);
nand U3111 (N_3111,N_2867,N_2556);
or U3112 (N_3112,N_2759,N_2583);
nand U3113 (N_3113,N_2990,N_2652);
nand U3114 (N_3114,N_2572,N_2898);
nor U3115 (N_3115,N_2949,N_2923);
and U3116 (N_3116,N_2950,N_2560);
or U3117 (N_3117,N_2625,N_2992);
or U3118 (N_3118,N_2589,N_2553);
and U3119 (N_3119,N_2805,N_2638);
nor U3120 (N_3120,N_2735,N_2579);
or U3121 (N_3121,N_2508,N_2939);
or U3122 (N_3122,N_2798,N_2658);
nand U3123 (N_3123,N_2655,N_2748);
nor U3124 (N_3124,N_2646,N_2845);
and U3125 (N_3125,N_2907,N_2788);
or U3126 (N_3126,N_2653,N_2716);
and U3127 (N_3127,N_2584,N_2942);
or U3128 (N_3128,N_2558,N_2708);
and U3129 (N_3129,N_2723,N_2628);
nand U3130 (N_3130,N_2843,N_2533);
nor U3131 (N_3131,N_2557,N_2709);
or U3132 (N_3132,N_2945,N_2972);
nand U3133 (N_3133,N_2552,N_2607);
nand U3134 (N_3134,N_2586,N_2643);
and U3135 (N_3135,N_2988,N_2930);
nand U3136 (N_3136,N_2755,N_2537);
nand U3137 (N_3137,N_2657,N_2864);
nor U3138 (N_3138,N_2765,N_2715);
nand U3139 (N_3139,N_2978,N_2800);
nor U3140 (N_3140,N_2606,N_2677);
and U3141 (N_3141,N_2627,N_2695);
and U3142 (N_3142,N_2760,N_2604);
nand U3143 (N_3143,N_2518,N_2666);
and U3144 (N_3144,N_2912,N_2896);
nand U3145 (N_3145,N_2862,N_2832);
or U3146 (N_3146,N_2924,N_2834);
nor U3147 (N_3147,N_2664,N_2612);
nor U3148 (N_3148,N_2551,N_2659);
nor U3149 (N_3149,N_2816,N_2642);
or U3150 (N_3150,N_2783,N_2622);
and U3151 (N_3151,N_2790,N_2770);
or U3152 (N_3152,N_2809,N_2894);
nor U3153 (N_3153,N_2514,N_2982);
and U3154 (N_3154,N_2866,N_2569);
and U3155 (N_3155,N_2710,N_2683);
or U3156 (N_3156,N_2528,N_2602);
and U3157 (N_3157,N_2743,N_2979);
nor U3158 (N_3158,N_2758,N_2520);
nor U3159 (N_3159,N_2675,N_2772);
nor U3160 (N_3160,N_2679,N_2740);
nand U3161 (N_3161,N_2865,N_2891);
or U3162 (N_3162,N_2925,N_2724);
or U3163 (N_3163,N_2996,N_2668);
nand U3164 (N_3164,N_2767,N_2641);
or U3165 (N_3165,N_2509,N_2836);
or U3166 (N_3166,N_2616,N_2591);
or U3167 (N_3167,N_2791,N_2938);
or U3168 (N_3168,N_2871,N_2780);
nand U3169 (N_3169,N_2624,N_2856);
nor U3170 (N_3170,N_2559,N_2640);
nand U3171 (N_3171,N_2807,N_2505);
nand U3172 (N_3172,N_2971,N_2573);
nor U3173 (N_3173,N_2737,N_2702);
xnor U3174 (N_3174,N_2543,N_2811);
and U3175 (N_3175,N_2926,N_2689);
and U3176 (N_3176,N_2803,N_2974);
nand U3177 (N_3177,N_2747,N_2900);
or U3178 (N_3178,N_2997,N_2609);
or U3179 (N_3179,N_2913,N_2582);
nor U3180 (N_3180,N_2530,N_2874);
nor U3181 (N_3181,N_2605,N_2825);
or U3182 (N_3182,N_2521,N_2804);
or U3183 (N_3183,N_2515,N_2821);
and U3184 (N_3184,N_2512,N_2827);
and U3185 (N_3185,N_2746,N_2660);
nor U3186 (N_3186,N_2574,N_2704);
nor U3187 (N_3187,N_2613,N_2739);
and U3188 (N_3188,N_2564,N_2776);
or U3189 (N_3189,N_2987,N_2550);
nand U3190 (N_3190,N_2532,N_2667);
nor U3191 (N_3191,N_2629,N_2853);
nor U3192 (N_3192,N_2728,N_2500);
or U3193 (N_3193,N_2969,N_2568);
nand U3194 (N_3194,N_2678,N_2944);
nand U3195 (N_3195,N_2662,N_2828);
nand U3196 (N_3196,N_2786,N_2819);
nand U3197 (N_3197,N_2523,N_2531);
and U3198 (N_3198,N_2754,N_2830);
and U3199 (N_3199,N_2921,N_2536);
or U3200 (N_3200,N_2636,N_2905);
and U3201 (N_3201,N_2840,N_2854);
nand U3202 (N_3202,N_2909,N_2787);
or U3203 (N_3203,N_2661,N_2868);
nand U3204 (N_3204,N_2507,N_2546);
nor U3205 (N_3205,N_2538,N_2852);
or U3206 (N_3206,N_2592,N_2890);
or U3207 (N_3207,N_2749,N_2782);
and U3208 (N_3208,N_2831,N_2644);
nor U3209 (N_3209,N_2984,N_2958);
or U3210 (N_3210,N_2887,N_2762);
nand U3211 (N_3211,N_2738,N_2889);
nand U3212 (N_3212,N_2863,N_2711);
xor U3213 (N_3213,N_2861,N_2750);
nand U3214 (N_3214,N_2663,N_2794);
or U3215 (N_3215,N_2870,N_2764);
nor U3216 (N_3216,N_2517,N_2608);
nand U3217 (N_3217,N_2860,N_2892);
or U3218 (N_3218,N_2736,N_2806);
nand U3219 (N_3219,N_2901,N_2637);
and U3220 (N_3220,N_2511,N_2581);
xnor U3221 (N_3221,N_2757,N_2957);
nor U3222 (N_3222,N_2525,N_2502);
nand U3223 (N_3223,N_2779,N_2720);
nor U3224 (N_3224,N_2571,N_2814);
or U3225 (N_3225,N_2917,N_2561);
and U3226 (N_3226,N_2623,N_2778);
nand U3227 (N_3227,N_2882,N_2857);
or U3228 (N_3228,N_2686,N_2697);
or U3229 (N_3229,N_2796,N_2555);
and U3230 (N_3230,N_2696,N_2888);
nand U3231 (N_3231,N_2911,N_2580);
nor U3232 (N_3232,N_2527,N_2681);
and U3233 (N_3233,N_2839,N_2943);
nand U3234 (N_3234,N_2793,N_2970);
nand U3235 (N_3235,N_2603,N_2619);
and U3236 (N_3236,N_2886,N_2915);
and U3237 (N_3237,N_2674,N_2705);
nand U3238 (N_3238,N_2545,N_2817);
or U3239 (N_3239,N_2994,N_2656);
and U3240 (N_3240,N_2928,N_2563);
nor U3241 (N_3241,N_2801,N_2615);
xnor U3242 (N_3242,N_2964,N_2998);
and U3243 (N_3243,N_2838,N_2785);
nand U3244 (N_3244,N_2630,N_2789);
and U3245 (N_3245,N_2510,N_2685);
or U3246 (N_3246,N_2918,N_2684);
and U3247 (N_3247,N_2645,N_2578);
nand U3248 (N_3248,N_2614,N_2953);
xor U3249 (N_3249,N_2781,N_2610);
nor U3250 (N_3250,N_2904,N_2576);
nand U3251 (N_3251,N_2773,N_2623);
nor U3252 (N_3252,N_2645,N_2925);
and U3253 (N_3253,N_2536,N_2941);
xnor U3254 (N_3254,N_2603,N_2698);
and U3255 (N_3255,N_2579,N_2500);
nand U3256 (N_3256,N_2789,N_2762);
or U3257 (N_3257,N_2704,N_2564);
or U3258 (N_3258,N_2910,N_2822);
nor U3259 (N_3259,N_2702,N_2899);
or U3260 (N_3260,N_2678,N_2600);
nand U3261 (N_3261,N_2506,N_2639);
nand U3262 (N_3262,N_2821,N_2878);
nand U3263 (N_3263,N_2834,N_2626);
nand U3264 (N_3264,N_2890,N_2927);
nor U3265 (N_3265,N_2771,N_2526);
or U3266 (N_3266,N_2964,N_2538);
nor U3267 (N_3267,N_2592,N_2857);
nor U3268 (N_3268,N_2582,N_2851);
or U3269 (N_3269,N_2636,N_2732);
nand U3270 (N_3270,N_2850,N_2672);
and U3271 (N_3271,N_2505,N_2647);
nand U3272 (N_3272,N_2600,N_2727);
or U3273 (N_3273,N_2874,N_2743);
nand U3274 (N_3274,N_2538,N_2558);
or U3275 (N_3275,N_2936,N_2538);
or U3276 (N_3276,N_2751,N_2900);
nand U3277 (N_3277,N_2852,N_2707);
and U3278 (N_3278,N_2683,N_2848);
or U3279 (N_3279,N_2874,N_2591);
and U3280 (N_3280,N_2999,N_2909);
nor U3281 (N_3281,N_2754,N_2587);
and U3282 (N_3282,N_2826,N_2898);
nand U3283 (N_3283,N_2738,N_2942);
and U3284 (N_3284,N_2716,N_2875);
nand U3285 (N_3285,N_2543,N_2814);
nand U3286 (N_3286,N_2545,N_2982);
or U3287 (N_3287,N_2844,N_2718);
and U3288 (N_3288,N_2534,N_2900);
or U3289 (N_3289,N_2848,N_2787);
nor U3290 (N_3290,N_2787,N_2584);
nand U3291 (N_3291,N_2553,N_2941);
or U3292 (N_3292,N_2905,N_2796);
nor U3293 (N_3293,N_2793,N_2683);
or U3294 (N_3294,N_2606,N_2979);
and U3295 (N_3295,N_2977,N_2598);
or U3296 (N_3296,N_2811,N_2569);
or U3297 (N_3297,N_2617,N_2683);
or U3298 (N_3298,N_2801,N_2563);
or U3299 (N_3299,N_2923,N_2547);
nor U3300 (N_3300,N_2712,N_2895);
nor U3301 (N_3301,N_2817,N_2715);
and U3302 (N_3302,N_2613,N_2781);
and U3303 (N_3303,N_2817,N_2622);
nand U3304 (N_3304,N_2694,N_2720);
nand U3305 (N_3305,N_2803,N_2505);
nor U3306 (N_3306,N_2651,N_2616);
nand U3307 (N_3307,N_2810,N_2674);
nor U3308 (N_3308,N_2698,N_2706);
or U3309 (N_3309,N_2593,N_2851);
nor U3310 (N_3310,N_2773,N_2505);
or U3311 (N_3311,N_2699,N_2647);
nand U3312 (N_3312,N_2861,N_2538);
nor U3313 (N_3313,N_2907,N_2901);
and U3314 (N_3314,N_2652,N_2940);
nor U3315 (N_3315,N_2768,N_2952);
nand U3316 (N_3316,N_2647,N_2503);
nand U3317 (N_3317,N_2675,N_2690);
or U3318 (N_3318,N_2921,N_2835);
or U3319 (N_3319,N_2968,N_2883);
nor U3320 (N_3320,N_2848,N_2970);
or U3321 (N_3321,N_2534,N_2937);
and U3322 (N_3322,N_2601,N_2919);
and U3323 (N_3323,N_2706,N_2511);
and U3324 (N_3324,N_2789,N_2735);
or U3325 (N_3325,N_2615,N_2850);
and U3326 (N_3326,N_2779,N_2842);
or U3327 (N_3327,N_2916,N_2614);
and U3328 (N_3328,N_2963,N_2923);
or U3329 (N_3329,N_2749,N_2589);
nand U3330 (N_3330,N_2858,N_2847);
and U3331 (N_3331,N_2504,N_2831);
and U3332 (N_3332,N_2910,N_2525);
nor U3333 (N_3333,N_2804,N_2700);
nor U3334 (N_3334,N_2670,N_2713);
or U3335 (N_3335,N_2596,N_2984);
or U3336 (N_3336,N_2652,N_2686);
and U3337 (N_3337,N_2588,N_2549);
nor U3338 (N_3338,N_2619,N_2609);
nor U3339 (N_3339,N_2833,N_2643);
or U3340 (N_3340,N_2805,N_2706);
and U3341 (N_3341,N_2572,N_2720);
nor U3342 (N_3342,N_2689,N_2694);
nor U3343 (N_3343,N_2771,N_2854);
nor U3344 (N_3344,N_2974,N_2687);
xnor U3345 (N_3345,N_2896,N_2657);
nand U3346 (N_3346,N_2998,N_2742);
or U3347 (N_3347,N_2954,N_2809);
nand U3348 (N_3348,N_2502,N_2885);
nand U3349 (N_3349,N_2737,N_2626);
and U3350 (N_3350,N_2607,N_2848);
nor U3351 (N_3351,N_2658,N_2511);
or U3352 (N_3352,N_2961,N_2920);
or U3353 (N_3353,N_2667,N_2877);
nand U3354 (N_3354,N_2870,N_2806);
or U3355 (N_3355,N_2503,N_2604);
or U3356 (N_3356,N_2608,N_2858);
and U3357 (N_3357,N_2834,N_2698);
or U3358 (N_3358,N_2856,N_2878);
nor U3359 (N_3359,N_2554,N_2509);
nand U3360 (N_3360,N_2953,N_2715);
nor U3361 (N_3361,N_2673,N_2978);
nand U3362 (N_3362,N_2812,N_2591);
nand U3363 (N_3363,N_2607,N_2767);
nand U3364 (N_3364,N_2946,N_2568);
nand U3365 (N_3365,N_2671,N_2551);
or U3366 (N_3366,N_2654,N_2846);
or U3367 (N_3367,N_2681,N_2997);
or U3368 (N_3368,N_2723,N_2649);
and U3369 (N_3369,N_2532,N_2627);
or U3370 (N_3370,N_2637,N_2536);
nor U3371 (N_3371,N_2581,N_2541);
nand U3372 (N_3372,N_2830,N_2569);
and U3373 (N_3373,N_2566,N_2591);
nor U3374 (N_3374,N_2544,N_2844);
nor U3375 (N_3375,N_2895,N_2864);
and U3376 (N_3376,N_2779,N_2703);
nand U3377 (N_3377,N_2611,N_2596);
nor U3378 (N_3378,N_2663,N_2594);
or U3379 (N_3379,N_2914,N_2608);
nor U3380 (N_3380,N_2507,N_2615);
xor U3381 (N_3381,N_2761,N_2778);
and U3382 (N_3382,N_2708,N_2997);
nor U3383 (N_3383,N_2530,N_2645);
nand U3384 (N_3384,N_2754,N_2975);
and U3385 (N_3385,N_2695,N_2631);
nor U3386 (N_3386,N_2504,N_2625);
nor U3387 (N_3387,N_2554,N_2704);
or U3388 (N_3388,N_2902,N_2607);
nor U3389 (N_3389,N_2828,N_2564);
and U3390 (N_3390,N_2814,N_2899);
nand U3391 (N_3391,N_2855,N_2513);
nor U3392 (N_3392,N_2633,N_2765);
or U3393 (N_3393,N_2743,N_2637);
and U3394 (N_3394,N_2919,N_2938);
nor U3395 (N_3395,N_2688,N_2583);
xor U3396 (N_3396,N_2803,N_2729);
or U3397 (N_3397,N_2768,N_2577);
nor U3398 (N_3398,N_2801,N_2883);
or U3399 (N_3399,N_2619,N_2624);
and U3400 (N_3400,N_2907,N_2651);
or U3401 (N_3401,N_2569,N_2601);
xor U3402 (N_3402,N_2574,N_2841);
and U3403 (N_3403,N_2521,N_2682);
nand U3404 (N_3404,N_2623,N_2964);
nand U3405 (N_3405,N_2917,N_2908);
and U3406 (N_3406,N_2614,N_2788);
or U3407 (N_3407,N_2599,N_2621);
and U3408 (N_3408,N_2832,N_2541);
or U3409 (N_3409,N_2989,N_2730);
nand U3410 (N_3410,N_2624,N_2806);
nand U3411 (N_3411,N_2719,N_2808);
nor U3412 (N_3412,N_2950,N_2774);
or U3413 (N_3413,N_2797,N_2549);
and U3414 (N_3414,N_2978,N_2761);
nor U3415 (N_3415,N_2989,N_2922);
or U3416 (N_3416,N_2968,N_2534);
nand U3417 (N_3417,N_2649,N_2712);
nor U3418 (N_3418,N_2717,N_2964);
and U3419 (N_3419,N_2912,N_2760);
and U3420 (N_3420,N_2522,N_2834);
and U3421 (N_3421,N_2621,N_2644);
nor U3422 (N_3422,N_2632,N_2517);
and U3423 (N_3423,N_2903,N_2944);
nor U3424 (N_3424,N_2806,N_2588);
nand U3425 (N_3425,N_2519,N_2563);
and U3426 (N_3426,N_2528,N_2668);
or U3427 (N_3427,N_2632,N_2780);
nand U3428 (N_3428,N_2820,N_2599);
nor U3429 (N_3429,N_2885,N_2820);
xor U3430 (N_3430,N_2522,N_2820);
nand U3431 (N_3431,N_2729,N_2839);
nor U3432 (N_3432,N_2969,N_2701);
or U3433 (N_3433,N_2960,N_2862);
nor U3434 (N_3434,N_2746,N_2793);
nor U3435 (N_3435,N_2591,N_2884);
nand U3436 (N_3436,N_2721,N_2621);
or U3437 (N_3437,N_2694,N_2906);
and U3438 (N_3438,N_2701,N_2575);
nor U3439 (N_3439,N_2765,N_2712);
nand U3440 (N_3440,N_2728,N_2531);
and U3441 (N_3441,N_2925,N_2790);
nor U3442 (N_3442,N_2751,N_2609);
and U3443 (N_3443,N_2999,N_2682);
or U3444 (N_3444,N_2566,N_2526);
nor U3445 (N_3445,N_2679,N_2990);
or U3446 (N_3446,N_2864,N_2974);
nand U3447 (N_3447,N_2922,N_2612);
or U3448 (N_3448,N_2761,N_2691);
nor U3449 (N_3449,N_2517,N_2754);
nor U3450 (N_3450,N_2798,N_2823);
xor U3451 (N_3451,N_2888,N_2707);
and U3452 (N_3452,N_2500,N_2853);
and U3453 (N_3453,N_2882,N_2737);
and U3454 (N_3454,N_2671,N_2768);
nor U3455 (N_3455,N_2599,N_2691);
nand U3456 (N_3456,N_2756,N_2707);
nor U3457 (N_3457,N_2644,N_2563);
or U3458 (N_3458,N_2935,N_2735);
nor U3459 (N_3459,N_2543,N_2644);
or U3460 (N_3460,N_2872,N_2953);
nor U3461 (N_3461,N_2738,N_2878);
nand U3462 (N_3462,N_2939,N_2837);
and U3463 (N_3463,N_2993,N_2825);
and U3464 (N_3464,N_2869,N_2817);
and U3465 (N_3465,N_2760,N_2632);
or U3466 (N_3466,N_2531,N_2638);
and U3467 (N_3467,N_2703,N_2601);
nand U3468 (N_3468,N_2806,N_2694);
nand U3469 (N_3469,N_2999,N_2918);
nor U3470 (N_3470,N_2641,N_2658);
nand U3471 (N_3471,N_2608,N_2634);
or U3472 (N_3472,N_2992,N_2891);
nor U3473 (N_3473,N_2835,N_2704);
and U3474 (N_3474,N_2697,N_2831);
and U3475 (N_3475,N_2626,N_2968);
or U3476 (N_3476,N_2826,N_2879);
nand U3477 (N_3477,N_2662,N_2776);
and U3478 (N_3478,N_2922,N_2782);
and U3479 (N_3479,N_2772,N_2594);
or U3480 (N_3480,N_2507,N_2981);
nor U3481 (N_3481,N_2794,N_2555);
nand U3482 (N_3482,N_2856,N_2827);
nor U3483 (N_3483,N_2654,N_2587);
nor U3484 (N_3484,N_2937,N_2707);
or U3485 (N_3485,N_2536,N_2817);
and U3486 (N_3486,N_2707,N_2641);
and U3487 (N_3487,N_2910,N_2549);
or U3488 (N_3488,N_2801,N_2981);
or U3489 (N_3489,N_2715,N_2689);
and U3490 (N_3490,N_2940,N_2599);
or U3491 (N_3491,N_2741,N_2623);
nor U3492 (N_3492,N_2767,N_2667);
or U3493 (N_3493,N_2504,N_2840);
or U3494 (N_3494,N_2509,N_2786);
nand U3495 (N_3495,N_2859,N_2863);
nor U3496 (N_3496,N_2621,N_2631);
and U3497 (N_3497,N_2866,N_2579);
nor U3498 (N_3498,N_2550,N_2921);
and U3499 (N_3499,N_2502,N_2689);
and U3500 (N_3500,N_3197,N_3068);
and U3501 (N_3501,N_3282,N_3439);
nor U3502 (N_3502,N_3041,N_3373);
or U3503 (N_3503,N_3288,N_3492);
or U3504 (N_3504,N_3482,N_3372);
nand U3505 (N_3505,N_3094,N_3264);
and U3506 (N_3506,N_3452,N_3299);
nor U3507 (N_3507,N_3378,N_3255);
nand U3508 (N_3508,N_3143,N_3252);
and U3509 (N_3509,N_3029,N_3271);
nand U3510 (N_3510,N_3075,N_3474);
nor U3511 (N_3511,N_3384,N_3367);
and U3512 (N_3512,N_3345,N_3462);
nand U3513 (N_3513,N_3153,N_3332);
and U3514 (N_3514,N_3013,N_3025);
nand U3515 (N_3515,N_3289,N_3381);
and U3516 (N_3516,N_3359,N_3489);
nor U3517 (N_3517,N_3159,N_3021);
and U3518 (N_3518,N_3083,N_3225);
nor U3519 (N_3519,N_3443,N_3056);
nand U3520 (N_3520,N_3238,N_3376);
nand U3521 (N_3521,N_3044,N_3087);
and U3522 (N_3522,N_3101,N_3274);
or U3523 (N_3523,N_3123,N_3292);
and U3524 (N_3524,N_3458,N_3002);
or U3525 (N_3525,N_3106,N_3410);
nand U3526 (N_3526,N_3118,N_3163);
nor U3527 (N_3527,N_3471,N_3052);
and U3528 (N_3528,N_3177,N_3257);
or U3529 (N_3529,N_3450,N_3334);
or U3530 (N_3530,N_3221,N_3499);
and U3531 (N_3531,N_3497,N_3327);
nor U3532 (N_3532,N_3435,N_3108);
or U3533 (N_3533,N_3433,N_3201);
or U3534 (N_3534,N_3165,N_3098);
nor U3535 (N_3535,N_3166,N_3062);
or U3536 (N_3536,N_3297,N_3429);
and U3537 (N_3537,N_3230,N_3045);
or U3538 (N_3538,N_3486,N_3001);
or U3539 (N_3539,N_3063,N_3447);
nand U3540 (N_3540,N_3047,N_3493);
nor U3541 (N_3541,N_3409,N_3220);
and U3542 (N_3542,N_3321,N_3399);
nand U3543 (N_3543,N_3005,N_3065);
or U3544 (N_3544,N_3003,N_3107);
nand U3545 (N_3545,N_3024,N_3295);
nand U3546 (N_3546,N_3188,N_3310);
and U3547 (N_3547,N_3073,N_3317);
and U3548 (N_3548,N_3416,N_3226);
and U3549 (N_3549,N_3028,N_3020);
nor U3550 (N_3550,N_3357,N_3354);
nand U3551 (N_3551,N_3451,N_3015);
nand U3552 (N_3552,N_3174,N_3356);
or U3553 (N_3553,N_3389,N_3371);
and U3554 (N_3554,N_3401,N_3491);
and U3555 (N_3555,N_3016,N_3228);
or U3556 (N_3556,N_3358,N_3190);
or U3557 (N_3557,N_3404,N_3270);
and U3558 (N_3558,N_3322,N_3046);
and U3559 (N_3559,N_3239,N_3223);
nand U3560 (N_3560,N_3480,N_3302);
and U3561 (N_3561,N_3039,N_3360);
nor U3562 (N_3562,N_3275,N_3236);
and U3563 (N_3563,N_3078,N_3030);
and U3564 (N_3564,N_3432,N_3396);
nand U3565 (N_3565,N_3192,N_3428);
and U3566 (N_3566,N_3129,N_3348);
and U3567 (N_3567,N_3392,N_3048);
or U3568 (N_3568,N_3457,N_3448);
nor U3569 (N_3569,N_3350,N_3121);
nor U3570 (N_3570,N_3290,N_3180);
and U3571 (N_3571,N_3495,N_3351);
nor U3572 (N_3572,N_3314,N_3479);
and U3573 (N_3573,N_3060,N_3261);
nand U3574 (N_3574,N_3200,N_3242);
nand U3575 (N_3575,N_3011,N_3050);
nor U3576 (N_3576,N_3125,N_3249);
nand U3577 (N_3577,N_3481,N_3339);
nor U3578 (N_3578,N_3364,N_3391);
nor U3579 (N_3579,N_3244,N_3146);
nand U3580 (N_3580,N_3199,N_3250);
nand U3581 (N_3581,N_3109,N_3352);
or U3582 (N_3582,N_3059,N_3186);
nor U3583 (N_3583,N_3415,N_3012);
xor U3584 (N_3584,N_3164,N_3222);
or U3585 (N_3585,N_3444,N_3144);
nor U3586 (N_3586,N_3366,N_3086);
nand U3587 (N_3587,N_3139,N_3173);
nor U3588 (N_3588,N_3120,N_3379);
or U3589 (N_3589,N_3387,N_3193);
or U3590 (N_3590,N_3038,N_3124);
and U3591 (N_3591,N_3122,N_3467);
and U3592 (N_3592,N_3307,N_3110);
or U3593 (N_3593,N_3422,N_3229);
or U3594 (N_3594,N_3105,N_3394);
nor U3595 (N_3595,N_3294,N_3100);
and U3596 (N_3596,N_3427,N_3390);
and U3597 (N_3597,N_3276,N_3205);
and U3598 (N_3598,N_3331,N_3206);
nor U3599 (N_3599,N_3355,N_3018);
nand U3600 (N_3600,N_3218,N_3343);
nand U3601 (N_3601,N_3049,N_3070);
nand U3602 (N_3602,N_3248,N_3162);
and U3603 (N_3603,N_3328,N_3388);
and U3604 (N_3604,N_3277,N_3405);
or U3605 (N_3605,N_3459,N_3338);
and U3606 (N_3606,N_3082,N_3305);
or U3607 (N_3607,N_3287,N_3363);
nor U3608 (N_3608,N_3449,N_3187);
nand U3609 (N_3609,N_3134,N_3067);
nor U3610 (N_3610,N_3335,N_3279);
nor U3611 (N_3611,N_3209,N_3019);
or U3612 (N_3612,N_3051,N_3494);
nor U3613 (N_3613,N_3437,N_3240);
and U3614 (N_3614,N_3176,N_3420);
nand U3615 (N_3615,N_3496,N_3483);
or U3616 (N_3616,N_3325,N_3419);
or U3617 (N_3617,N_3140,N_3278);
nand U3618 (N_3618,N_3320,N_3233);
and U3619 (N_3619,N_3397,N_3333);
nor U3620 (N_3620,N_3074,N_3076);
or U3621 (N_3621,N_3145,N_3172);
nand U3622 (N_3622,N_3178,N_3008);
nor U3623 (N_3623,N_3303,N_3309);
nand U3624 (N_3624,N_3440,N_3114);
nand U3625 (N_3625,N_3217,N_3465);
nor U3626 (N_3626,N_3231,N_3402);
nor U3627 (N_3627,N_3202,N_3204);
nor U3628 (N_3628,N_3156,N_3254);
or U3629 (N_3629,N_3344,N_3263);
nor U3630 (N_3630,N_3215,N_3211);
or U3631 (N_3631,N_3301,N_3113);
nand U3632 (N_3632,N_3219,N_3417);
and U3633 (N_3633,N_3374,N_3132);
nor U3634 (N_3634,N_3088,N_3179);
nand U3635 (N_3635,N_3256,N_3407);
and U3636 (N_3636,N_3414,N_3365);
nand U3637 (N_3637,N_3247,N_3408);
and U3638 (N_3638,N_3484,N_3071);
and U3639 (N_3639,N_3403,N_3023);
and U3640 (N_3640,N_3085,N_3477);
and U3641 (N_3641,N_3473,N_3102);
nand U3642 (N_3642,N_3423,N_3099);
nor U3643 (N_3643,N_3418,N_3184);
or U3644 (N_3644,N_3269,N_3196);
nor U3645 (N_3645,N_3326,N_3042);
or U3646 (N_3646,N_3171,N_3235);
nand U3647 (N_3647,N_3412,N_3136);
nand U3648 (N_3648,N_3468,N_3490);
or U3649 (N_3649,N_3137,N_3293);
or U3650 (N_3650,N_3285,N_3434);
or U3651 (N_3651,N_3323,N_3361);
and U3652 (N_3652,N_3154,N_3266);
and U3653 (N_3653,N_3097,N_3111);
nor U3654 (N_3654,N_3488,N_3198);
and U3655 (N_3655,N_3259,N_3284);
nor U3656 (N_3656,N_3079,N_3161);
nand U3657 (N_3657,N_3368,N_3461);
nand U3658 (N_3658,N_3031,N_3445);
nand U3659 (N_3659,N_3470,N_3214);
nor U3660 (N_3660,N_3064,N_3426);
nand U3661 (N_3661,N_3128,N_3181);
nor U3662 (N_3662,N_3382,N_3095);
or U3663 (N_3663,N_3103,N_3246);
nand U3664 (N_3664,N_3112,N_3116);
nand U3665 (N_3665,N_3189,N_3195);
nor U3666 (N_3666,N_3476,N_3232);
xor U3667 (N_3667,N_3436,N_3340);
nand U3668 (N_3668,N_3010,N_3286);
nand U3669 (N_3669,N_3182,N_3130);
nand U3670 (N_3670,N_3273,N_3280);
and U3671 (N_3671,N_3329,N_3341);
or U3672 (N_3672,N_3478,N_3148);
nor U3673 (N_3673,N_3006,N_3370);
nand U3674 (N_3674,N_3265,N_3191);
nor U3675 (N_3675,N_3241,N_3253);
nand U3676 (N_3676,N_3258,N_3413);
nor U3677 (N_3677,N_3375,N_3089);
and U3678 (N_3678,N_3267,N_3066);
nand U3679 (N_3679,N_3315,N_3456);
or U3680 (N_3680,N_3152,N_3119);
nor U3681 (N_3681,N_3061,N_3243);
or U3682 (N_3682,N_3040,N_3306);
and U3683 (N_3683,N_3336,N_3393);
or U3684 (N_3684,N_3349,N_3210);
nand U3685 (N_3685,N_3069,N_3141);
nor U3686 (N_3686,N_3380,N_3212);
nand U3687 (N_3687,N_3469,N_3281);
nand U3688 (N_3688,N_3017,N_3183);
nand U3689 (N_3689,N_3117,N_3147);
nand U3690 (N_3690,N_3425,N_3245);
and U3691 (N_3691,N_3057,N_3460);
or U3692 (N_3692,N_3272,N_3055);
or U3693 (N_3693,N_3454,N_3369);
nor U3694 (N_3694,N_3167,N_3158);
and U3695 (N_3695,N_3026,N_3446);
nor U3696 (N_3696,N_3313,N_3395);
or U3697 (N_3697,N_3007,N_3421);
and U3698 (N_3698,N_3022,N_3090);
nor U3699 (N_3699,N_3438,N_3131);
or U3700 (N_3700,N_3169,N_3463);
nor U3701 (N_3701,N_3027,N_3308);
nand U3702 (N_3702,N_3466,N_3072);
nor U3703 (N_3703,N_3377,N_3298);
or U3704 (N_3704,N_3283,N_3155);
nor U3705 (N_3705,N_3092,N_3096);
nand U3706 (N_3706,N_3406,N_3054);
or U3707 (N_3707,N_3398,N_3033);
and U3708 (N_3708,N_3224,N_3431);
or U3709 (N_3709,N_3311,N_3160);
or U3710 (N_3710,N_3077,N_3442);
or U3711 (N_3711,N_3150,N_3135);
or U3712 (N_3712,N_3126,N_3138);
or U3713 (N_3713,N_3034,N_3216);
nor U3714 (N_3714,N_3081,N_3151);
or U3715 (N_3715,N_3170,N_3485);
nor U3716 (N_3716,N_3014,N_3262);
nor U3717 (N_3717,N_3227,N_3383);
nand U3718 (N_3718,N_3304,N_3487);
nor U3719 (N_3719,N_3342,N_3009);
nor U3720 (N_3720,N_3093,N_3453);
nor U3721 (N_3721,N_3175,N_3347);
and U3722 (N_3722,N_3208,N_3080);
and U3723 (N_3723,N_3157,N_3324);
or U3724 (N_3724,N_3203,N_3004);
nand U3725 (N_3725,N_3035,N_3316);
and U3726 (N_3726,N_3346,N_3260);
and U3727 (N_3727,N_3168,N_3115);
or U3728 (N_3728,N_3091,N_3237);
and U3729 (N_3729,N_3291,N_3475);
and U3730 (N_3730,N_3207,N_3185);
and U3731 (N_3731,N_3037,N_3213);
or U3732 (N_3732,N_3424,N_3053);
or U3733 (N_3733,N_3337,N_3441);
and U3734 (N_3734,N_3127,N_3300);
nor U3735 (N_3735,N_3455,N_3385);
nand U3736 (N_3736,N_3296,N_3036);
nand U3737 (N_3737,N_3430,N_3353);
nor U3738 (N_3738,N_3084,N_3318);
nand U3739 (N_3739,N_3194,N_3498);
xor U3740 (N_3740,N_3234,N_3472);
nand U3741 (N_3741,N_3319,N_3032);
or U3742 (N_3742,N_3268,N_3058);
nand U3743 (N_3743,N_3251,N_3362);
nor U3744 (N_3744,N_3464,N_3400);
nand U3745 (N_3745,N_3386,N_3133);
nor U3746 (N_3746,N_3312,N_3149);
or U3747 (N_3747,N_3000,N_3142);
or U3748 (N_3748,N_3043,N_3104);
or U3749 (N_3749,N_3411,N_3330);
nor U3750 (N_3750,N_3258,N_3390);
nand U3751 (N_3751,N_3459,N_3464);
nand U3752 (N_3752,N_3440,N_3007);
nand U3753 (N_3753,N_3219,N_3254);
nor U3754 (N_3754,N_3355,N_3443);
or U3755 (N_3755,N_3396,N_3487);
and U3756 (N_3756,N_3111,N_3121);
and U3757 (N_3757,N_3147,N_3144);
and U3758 (N_3758,N_3079,N_3498);
nor U3759 (N_3759,N_3103,N_3017);
and U3760 (N_3760,N_3266,N_3101);
or U3761 (N_3761,N_3383,N_3281);
nor U3762 (N_3762,N_3347,N_3096);
and U3763 (N_3763,N_3368,N_3415);
and U3764 (N_3764,N_3206,N_3454);
nor U3765 (N_3765,N_3372,N_3047);
or U3766 (N_3766,N_3044,N_3006);
nor U3767 (N_3767,N_3113,N_3407);
or U3768 (N_3768,N_3211,N_3352);
nor U3769 (N_3769,N_3471,N_3379);
or U3770 (N_3770,N_3090,N_3151);
nor U3771 (N_3771,N_3309,N_3327);
nor U3772 (N_3772,N_3158,N_3104);
nor U3773 (N_3773,N_3179,N_3028);
or U3774 (N_3774,N_3136,N_3285);
nand U3775 (N_3775,N_3171,N_3331);
and U3776 (N_3776,N_3206,N_3486);
nand U3777 (N_3777,N_3154,N_3319);
nand U3778 (N_3778,N_3003,N_3307);
and U3779 (N_3779,N_3145,N_3050);
nor U3780 (N_3780,N_3245,N_3243);
nor U3781 (N_3781,N_3058,N_3339);
nand U3782 (N_3782,N_3399,N_3288);
nor U3783 (N_3783,N_3424,N_3272);
nor U3784 (N_3784,N_3390,N_3188);
or U3785 (N_3785,N_3452,N_3345);
nand U3786 (N_3786,N_3475,N_3253);
or U3787 (N_3787,N_3183,N_3241);
or U3788 (N_3788,N_3471,N_3376);
or U3789 (N_3789,N_3157,N_3085);
or U3790 (N_3790,N_3258,N_3089);
nand U3791 (N_3791,N_3087,N_3226);
nand U3792 (N_3792,N_3476,N_3341);
or U3793 (N_3793,N_3116,N_3063);
or U3794 (N_3794,N_3300,N_3107);
and U3795 (N_3795,N_3275,N_3163);
nor U3796 (N_3796,N_3090,N_3005);
and U3797 (N_3797,N_3088,N_3173);
nand U3798 (N_3798,N_3256,N_3141);
nor U3799 (N_3799,N_3420,N_3363);
or U3800 (N_3800,N_3442,N_3404);
nor U3801 (N_3801,N_3424,N_3222);
xor U3802 (N_3802,N_3245,N_3431);
nand U3803 (N_3803,N_3071,N_3326);
or U3804 (N_3804,N_3462,N_3383);
nor U3805 (N_3805,N_3405,N_3090);
and U3806 (N_3806,N_3034,N_3443);
and U3807 (N_3807,N_3157,N_3138);
or U3808 (N_3808,N_3458,N_3202);
or U3809 (N_3809,N_3360,N_3361);
nand U3810 (N_3810,N_3450,N_3420);
nand U3811 (N_3811,N_3361,N_3417);
nor U3812 (N_3812,N_3485,N_3482);
and U3813 (N_3813,N_3050,N_3293);
nor U3814 (N_3814,N_3307,N_3005);
nor U3815 (N_3815,N_3062,N_3180);
nor U3816 (N_3816,N_3215,N_3120);
nand U3817 (N_3817,N_3203,N_3470);
and U3818 (N_3818,N_3173,N_3118);
nand U3819 (N_3819,N_3077,N_3096);
or U3820 (N_3820,N_3410,N_3355);
and U3821 (N_3821,N_3005,N_3189);
nand U3822 (N_3822,N_3246,N_3011);
and U3823 (N_3823,N_3410,N_3427);
nand U3824 (N_3824,N_3451,N_3222);
nand U3825 (N_3825,N_3453,N_3353);
nor U3826 (N_3826,N_3497,N_3093);
nor U3827 (N_3827,N_3299,N_3205);
or U3828 (N_3828,N_3205,N_3314);
and U3829 (N_3829,N_3062,N_3343);
or U3830 (N_3830,N_3033,N_3115);
and U3831 (N_3831,N_3450,N_3366);
or U3832 (N_3832,N_3232,N_3330);
or U3833 (N_3833,N_3095,N_3148);
and U3834 (N_3834,N_3109,N_3488);
or U3835 (N_3835,N_3015,N_3019);
or U3836 (N_3836,N_3170,N_3423);
and U3837 (N_3837,N_3490,N_3054);
nand U3838 (N_3838,N_3319,N_3024);
and U3839 (N_3839,N_3393,N_3409);
nand U3840 (N_3840,N_3027,N_3486);
nand U3841 (N_3841,N_3304,N_3363);
or U3842 (N_3842,N_3091,N_3376);
or U3843 (N_3843,N_3037,N_3022);
or U3844 (N_3844,N_3114,N_3200);
or U3845 (N_3845,N_3071,N_3358);
or U3846 (N_3846,N_3132,N_3337);
nor U3847 (N_3847,N_3245,N_3311);
and U3848 (N_3848,N_3123,N_3362);
or U3849 (N_3849,N_3057,N_3066);
nand U3850 (N_3850,N_3084,N_3090);
nor U3851 (N_3851,N_3376,N_3029);
or U3852 (N_3852,N_3427,N_3480);
and U3853 (N_3853,N_3244,N_3355);
and U3854 (N_3854,N_3199,N_3312);
or U3855 (N_3855,N_3374,N_3172);
or U3856 (N_3856,N_3499,N_3370);
nand U3857 (N_3857,N_3058,N_3342);
nand U3858 (N_3858,N_3369,N_3379);
nor U3859 (N_3859,N_3212,N_3355);
or U3860 (N_3860,N_3099,N_3308);
or U3861 (N_3861,N_3322,N_3190);
or U3862 (N_3862,N_3379,N_3171);
or U3863 (N_3863,N_3300,N_3147);
nand U3864 (N_3864,N_3239,N_3262);
and U3865 (N_3865,N_3421,N_3476);
nor U3866 (N_3866,N_3392,N_3490);
and U3867 (N_3867,N_3324,N_3469);
and U3868 (N_3868,N_3240,N_3012);
or U3869 (N_3869,N_3309,N_3497);
and U3870 (N_3870,N_3066,N_3131);
nand U3871 (N_3871,N_3230,N_3256);
nor U3872 (N_3872,N_3432,N_3047);
or U3873 (N_3873,N_3353,N_3420);
and U3874 (N_3874,N_3211,N_3401);
or U3875 (N_3875,N_3126,N_3388);
and U3876 (N_3876,N_3356,N_3349);
nor U3877 (N_3877,N_3472,N_3035);
and U3878 (N_3878,N_3405,N_3365);
nand U3879 (N_3879,N_3072,N_3211);
nor U3880 (N_3880,N_3170,N_3042);
nor U3881 (N_3881,N_3161,N_3267);
nand U3882 (N_3882,N_3301,N_3112);
nand U3883 (N_3883,N_3103,N_3327);
nor U3884 (N_3884,N_3373,N_3202);
or U3885 (N_3885,N_3204,N_3297);
nand U3886 (N_3886,N_3425,N_3057);
nor U3887 (N_3887,N_3340,N_3037);
or U3888 (N_3888,N_3479,N_3044);
or U3889 (N_3889,N_3307,N_3232);
or U3890 (N_3890,N_3091,N_3170);
nand U3891 (N_3891,N_3494,N_3232);
nand U3892 (N_3892,N_3100,N_3163);
nand U3893 (N_3893,N_3062,N_3146);
or U3894 (N_3894,N_3322,N_3490);
nand U3895 (N_3895,N_3042,N_3456);
or U3896 (N_3896,N_3303,N_3420);
nand U3897 (N_3897,N_3291,N_3338);
nand U3898 (N_3898,N_3032,N_3234);
nor U3899 (N_3899,N_3238,N_3477);
nor U3900 (N_3900,N_3478,N_3300);
nor U3901 (N_3901,N_3475,N_3157);
and U3902 (N_3902,N_3331,N_3378);
nand U3903 (N_3903,N_3208,N_3358);
nor U3904 (N_3904,N_3383,N_3280);
nor U3905 (N_3905,N_3256,N_3332);
and U3906 (N_3906,N_3104,N_3454);
or U3907 (N_3907,N_3468,N_3053);
and U3908 (N_3908,N_3408,N_3002);
nand U3909 (N_3909,N_3420,N_3406);
nand U3910 (N_3910,N_3276,N_3227);
nand U3911 (N_3911,N_3164,N_3413);
nand U3912 (N_3912,N_3125,N_3291);
and U3913 (N_3913,N_3276,N_3202);
or U3914 (N_3914,N_3436,N_3233);
nand U3915 (N_3915,N_3442,N_3448);
nor U3916 (N_3916,N_3353,N_3097);
nand U3917 (N_3917,N_3403,N_3266);
and U3918 (N_3918,N_3346,N_3088);
or U3919 (N_3919,N_3262,N_3486);
and U3920 (N_3920,N_3284,N_3497);
nand U3921 (N_3921,N_3452,N_3079);
or U3922 (N_3922,N_3114,N_3061);
or U3923 (N_3923,N_3339,N_3085);
or U3924 (N_3924,N_3327,N_3194);
and U3925 (N_3925,N_3188,N_3205);
nor U3926 (N_3926,N_3178,N_3317);
nor U3927 (N_3927,N_3398,N_3045);
and U3928 (N_3928,N_3006,N_3345);
or U3929 (N_3929,N_3376,N_3182);
or U3930 (N_3930,N_3407,N_3486);
nand U3931 (N_3931,N_3335,N_3452);
and U3932 (N_3932,N_3367,N_3325);
and U3933 (N_3933,N_3492,N_3250);
or U3934 (N_3934,N_3155,N_3187);
and U3935 (N_3935,N_3408,N_3202);
or U3936 (N_3936,N_3299,N_3227);
and U3937 (N_3937,N_3304,N_3131);
or U3938 (N_3938,N_3243,N_3117);
or U3939 (N_3939,N_3276,N_3316);
and U3940 (N_3940,N_3419,N_3407);
nor U3941 (N_3941,N_3415,N_3134);
nand U3942 (N_3942,N_3106,N_3232);
nor U3943 (N_3943,N_3073,N_3312);
or U3944 (N_3944,N_3005,N_3375);
or U3945 (N_3945,N_3258,N_3117);
or U3946 (N_3946,N_3216,N_3026);
or U3947 (N_3947,N_3196,N_3408);
and U3948 (N_3948,N_3460,N_3203);
nor U3949 (N_3949,N_3227,N_3151);
nor U3950 (N_3950,N_3035,N_3479);
and U3951 (N_3951,N_3477,N_3251);
nand U3952 (N_3952,N_3319,N_3487);
nand U3953 (N_3953,N_3215,N_3293);
or U3954 (N_3954,N_3315,N_3182);
or U3955 (N_3955,N_3022,N_3053);
nor U3956 (N_3956,N_3026,N_3233);
nor U3957 (N_3957,N_3220,N_3383);
and U3958 (N_3958,N_3167,N_3478);
or U3959 (N_3959,N_3268,N_3222);
nand U3960 (N_3960,N_3030,N_3443);
xnor U3961 (N_3961,N_3333,N_3077);
or U3962 (N_3962,N_3195,N_3059);
nand U3963 (N_3963,N_3015,N_3218);
or U3964 (N_3964,N_3076,N_3376);
or U3965 (N_3965,N_3016,N_3237);
nand U3966 (N_3966,N_3409,N_3309);
and U3967 (N_3967,N_3047,N_3266);
or U3968 (N_3968,N_3130,N_3423);
nand U3969 (N_3969,N_3145,N_3196);
nand U3970 (N_3970,N_3210,N_3203);
nand U3971 (N_3971,N_3262,N_3317);
nand U3972 (N_3972,N_3399,N_3298);
nand U3973 (N_3973,N_3363,N_3142);
nand U3974 (N_3974,N_3410,N_3306);
nor U3975 (N_3975,N_3425,N_3485);
or U3976 (N_3976,N_3418,N_3034);
nor U3977 (N_3977,N_3268,N_3351);
nand U3978 (N_3978,N_3002,N_3216);
and U3979 (N_3979,N_3420,N_3386);
and U3980 (N_3980,N_3157,N_3192);
and U3981 (N_3981,N_3208,N_3435);
nand U3982 (N_3982,N_3483,N_3406);
and U3983 (N_3983,N_3164,N_3332);
and U3984 (N_3984,N_3493,N_3464);
nand U3985 (N_3985,N_3484,N_3378);
nand U3986 (N_3986,N_3141,N_3331);
nand U3987 (N_3987,N_3362,N_3445);
nor U3988 (N_3988,N_3353,N_3196);
and U3989 (N_3989,N_3392,N_3416);
nand U3990 (N_3990,N_3061,N_3399);
nand U3991 (N_3991,N_3190,N_3077);
nor U3992 (N_3992,N_3489,N_3446);
nor U3993 (N_3993,N_3160,N_3113);
nor U3994 (N_3994,N_3432,N_3039);
nand U3995 (N_3995,N_3467,N_3110);
nor U3996 (N_3996,N_3017,N_3167);
xnor U3997 (N_3997,N_3026,N_3164);
nand U3998 (N_3998,N_3465,N_3192);
or U3999 (N_3999,N_3312,N_3390);
nand U4000 (N_4000,N_3918,N_3678);
or U4001 (N_4001,N_3848,N_3560);
and U4002 (N_4002,N_3594,N_3648);
or U4003 (N_4003,N_3994,N_3601);
or U4004 (N_4004,N_3725,N_3645);
nand U4005 (N_4005,N_3552,N_3523);
and U4006 (N_4006,N_3893,N_3957);
or U4007 (N_4007,N_3618,N_3781);
nand U4008 (N_4008,N_3865,N_3608);
or U4009 (N_4009,N_3586,N_3628);
nor U4010 (N_4010,N_3988,N_3640);
nor U4011 (N_4011,N_3903,N_3967);
nor U4012 (N_4012,N_3672,N_3683);
nor U4013 (N_4013,N_3923,N_3687);
nor U4014 (N_4014,N_3634,N_3636);
and U4015 (N_4015,N_3630,N_3774);
or U4016 (N_4016,N_3802,N_3579);
nand U4017 (N_4017,N_3732,N_3599);
and U4018 (N_4018,N_3713,N_3897);
nand U4019 (N_4019,N_3797,N_3717);
nand U4020 (N_4020,N_3724,N_3894);
nor U4021 (N_4021,N_3766,N_3712);
or U4022 (N_4022,N_3580,N_3547);
or U4023 (N_4023,N_3762,N_3696);
and U4024 (N_4024,N_3503,N_3790);
and U4025 (N_4025,N_3557,N_3595);
nor U4026 (N_4026,N_3705,N_3651);
nor U4027 (N_4027,N_3920,N_3829);
nor U4028 (N_4028,N_3597,N_3900);
and U4029 (N_4029,N_3864,N_3840);
or U4030 (N_4030,N_3937,N_3989);
and U4031 (N_4031,N_3824,N_3924);
and U4032 (N_4032,N_3615,N_3772);
or U4033 (N_4033,N_3735,N_3784);
nor U4034 (N_4034,N_3609,N_3926);
nor U4035 (N_4035,N_3853,N_3878);
nand U4036 (N_4036,N_3688,N_3767);
nor U4037 (N_4037,N_3568,N_3936);
or U4038 (N_4038,N_3838,N_3791);
nor U4039 (N_4039,N_3553,N_3941);
xnor U4040 (N_4040,N_3535,N_3642);
nor U4041 (N_4041,N_3583,N_3663);
and U4042 (N_4042,N_3916,N_3700);
or U4043 (N_4043,N_3985,N_3955);
or U4044 (N_4044,N_3549,N_3953);
nor U4045 (N_4045,N_3999,N_3668);
nor U4046 (N_4046,N_3904,N_3911);
nand U4047 (N_4047,N_3611,N_3525);
nor U4048 (N_4048,N_3795,N_3852);
nand U4049 (N_4049,N_3960,N_3973);
and U4050 (N_4050,N_3914,N_3565);
nand U4051 (N_4051,N_3971,N_3555);
nor U4052 (N_4052,N_3585,N_3970);
and U4053 (N_4053,N_3868,N_3661);
and U4054 (N_4054,N_3606,N_3607);
and U4055 (N_4055,N_3947,N_3785);
nor U4056 (N_4056,N_3563,N_3823);
or U4057 (N_4057,N_3614,N_3912);
and U4058 (N_4058,N_3892,N_3908);
and U4059 (N_4059,N_3910,N_3657);
nand U4060 (N_4060,N_3677,N_3812);
and U4061 (N_4061,N_3662,N_3980);
xor U4062 (N_4062,N_3819,N_3537);
nor U4063 (N_4063,N_3575,N_3899);
nor U4064 (N_4064,N_3898,N_3627);
nor U4065 (N_4065,N_3885,N_3682);
or U4066 (N_4066,N_3693,N_3629);
and U4067 (N_4067,N_3534,N_3993);
and U4068 (N_4068,N_3773,N_3799);
nand U4069 (N_4069,N_3620,N_3593);
nand U4070 (N_4070,N_3760,N_3942);
or U4071 (N_4071,N_3689,N_3741);
and U4072 (N_4072,N_3940,N_3654);
and U4073 (N_4073,N_3917,N_3604);
nor U4074 (N_4074,N_3851,N_3948);
and U4075 (N_4075,N_3979,N_3816);
or U4076 (N_4076,N_3850,N_3633);
or U4077 (N_4077,N_3887,N_3830);
or U4078 (N_4078,N_3703,N_3788);
nor U4079 (N_4079,N_3653,N_3721);
and U4080 (N_4080,N_3775,N_3745);
and U4081 (N_4081,N_3572,N_3965);
or U4082 (N_4082,N_3706,N_3810);
nand U4083 (N_4083,N_3617,N_3927);
nand U4084 (N_4084,N_3641,N_3876);
nand U4085 (N_4085,N_3938,N_3660);
nor U4086 (N_4086,N_3834,N_3991);
nor U4087 (N_4087,N_3872,N_3733);
nand U4088 (N_4088,N_3931,N_3747);
nor U4089 (N_4089,N_3859,N_3949);
nor U4090 (N_4090,N_3544,N_3727);
or U4091 (N_4091,N_3809,N_3820);
and U4092 (N_4092,N_3765,N_3612);
or U4093 (N_4093,N_3811,N_3891);
and U4094 (N_4094,N_3932,N_3956);
nand U4095 (N_4095,N_3977,N_3744);
and U4096 (N_4096,N_3909,N_3521);
nor U4097 (N_4097,N_3888,N_3874);
nand U4098 (N_4098,N_3519,N_3805);
nor U4099 (N_4099,N_3704,N_3800);
nor U4100 (N_4100,N_3846,N_3930);
or U4101 (N_4101,N_3778,N_3694);
nor U4102 (N_4102,N_3906,N_3798);
nand U4103 (N_4103,N_3610,N_3670);
and U4104 (N_4104,N_3709,N_3540);
nor U4105 (N_4105,N_3818,N_3839);
nor U4106 (N_4106,N_3626,N_3666);
nand U4107 (N_4107,N_3833,N_3987);
or U4108 (N_4108,N_3720,N_3964);
and U4109 (N_4109,N_3808,N_3777);
nand U4110 (N_4110,N_3982,N_3837);
or U4111 (N_4111,N_3913,N_3621);
nor U4112 (N_4112,N_3881,N_3718);
and U4113 (N_4113,N_3925,N_3889);
nor U4114 (N_4114,N_3740,N_3510);
nor U4115 (N_4115,N_3558,N_3751);
nor U4116 (N_4116,N_3602,N_3684);
and U4117 (N_4117,N_3961,N_3655);
and U4118 (N_4118,N_3590,N_3723);
nand U4119 (N_4119,N_3821,N_3841);
nor U4120 (N_4120,N_3992,N_3962);
nand U4121 (N_4121,N_3545,N_3532);
or U4122 (N_4122,N_3562,N_3815);
or U4123 (N_4123,N_3807,N_3637);
or U4124 (N_4124,N_3921,N_3543);
and U4125 (N_4125,N_3652,N_3857);
nand U4126 (N_4126,N_3755,N_3582);
and U4127 (N_4127,N_3915,N_3516);
and U4128 (N_4128,N_3561,N_3500);
and U4129 (N_4129,N_3571,N_3715);
nand U4130 (N_4130,N_3928,N_3929);
and U4131 (N_4131,N_3882,N_3554);
and U4132 (N_4132,N_3530,N_3714);
and U4133 (N_4133,N_3842,N_3761);
nand U4134 (N_4134,N_3613,N_3646);
and U4135 (N_4135,N_3573,N_3952);
nand U4136 (N_4136,N_3591,N_3729);
nand U4137 (N_4137,N_3763,N_3522);
or U4138 (N_4138,N_3528,N_3697);
and U4139 (N_4139,N_3849,N_3556);
nor U4140 (N_4140,N_3526,N_3538);
nand U4141 (N_4141,N_3509,N_3998);
nor U4142 (N_4142,N_3983,N_3650);
nor U4143 (N_4143,N_3665,N_3954);
and U4144 (N_4144,N_3875,N_3539);
and U4145 (N_4145,N_3708,N_3863);
nor U4146 (N_4146,N_3879,N_3787);
nand U4147 (N_4147,N_3649,N_3542);
and U4148 (N_4148,N_3736,N_3685);
nor U4149 (N_4149,N_3635,N_3782);
or U4150 (N_4150,N_3789,N_3548);
nor U4151 (N_4151,N_3935,N_3739);
or U4152 (N_4152,N_3623,N_3570);
or U4153 (N_4153,N_3513,N_3959);
nand U4154 (N_4154,N_3968,N_3944);
or U4155 (N_4155,N_3995,N_3581);
or U4156 (N_4156,N_3716,N_3836);
xor U4157 (N_4157,N_3862,N_3598);
and U4158 (N_4158,N_3576,N_3981);
nand U4159 (N_4159,N_3592,N_3691);
nor U4160 (N_4160,N_3858,N_3742);
nand U4161 (N_4161,N_3814,N_3754);
and U4162 (N_4162,N_3825,N_3536);
or U4163 (N_4163,N_3667,N_3669);
nand U4164 (N_4164,N_3531,N_3769);
and U4165 (N_4165,N_3871,N_3616);
and U4166 (N_4166,N_3806,N_3776);
or U4167 (N_4167,N_3647,N_3845);
and U4168 (N_4168,N_3564,N_3551);
or U4169 (N_4169,N_3946,N_3835);
nand U4170 (N_4170,N_3511,N_3905);
nor U4171 (N_4171,N_3753,N_3870);
nor U4172 (N_4172,N_3577,N_3867);
nand U4173 (N_4173,N_3675,N_3939);
and U4174 (N_4174,N_3951,N_3737);
or U4175 (N_4175,N_3780,N_3710);
nand U4176 (N_4176,N_3644,N_3746);
nor U4177 (N_4177,N_3786,N_3886);
nand U4178 (N_4178,N_3950,N_3728);
nand U4179 (N_4179,N_3984,N_3587);
nand U4180 (N_4180,N_3719,N_3707);
and U4181 (N_4181,N_3966,N_3877);
and U4182 (N_4182,N_3501,N_3958);
or U4183 (N_4183,N_3890,N_3758);
or U4184 (N_4184,N_3726,N_3550);
nor U4185 (N_4185,N_3731,N_3796);
nor U4186 (N_4186,N_3896,N_3673);
or U4187 (N_4187,N_3690,N_3686);
nor U4188 (N_4188,N_3856,N_3658);
and U4189 (N_4189,N_3515,N_3880);
or U4190 (N_4190,N_3996,N_3822);
nor U4191 (N_4191,N_3698,N_3801);
nor U4192 (N_4192,N_3794,N_3638);
or U4193 (N_4193,N_3679,N_3990);
and U4194 (N_4194,N_3533,N_3943);
or U4195 (N_4195,N_3699,N_3507);
or U4196 (N_4196,N_3559,N_3974);
nand U4197 (N_4197,N_3884,N_3596);
nor U4198 (N_4198,N_3768,N_3676);
or U4199 (N_4199,N_3907,N_3975);
or U4200 (N_4200,N_3631,N_3792);
and U4201 (N_4201,N_3963,N_3783);
and U4202 (N_4202,N_3681,N_3771);
nor U4203 (N_4203,N_3770,N_3695);
and U4204 (N_4204,N_3860,N_3529);
nor U4205 (N_4205,N_3828,N_3978);
or U4206 (N_4206,N_3643,N_3502);
and U4207 (N_4207,N_3517,N_3506);
or U4208 (N_4208,N_3748,N_3520);
and U4209 (N_4209,N_3831,N_3826);
or U4210 (N_4210,N_3674,N_3779);
nor U4211 (N_4211,N_3873,N_3622);
nand U4212 (N_4212,N_3969,N_3584);
nor U4213 (N_4213,N_3578,N_3569);
nand U4214 (N_4214,N_3813,N_3827);
nor U4215 (N_4215,N_3804,N_3750);
or U4216 (N_4216,N_3866,N_3701);
or U4217 (N_4217,N_3588,N_3605);
or U4218 (N_4218,N_3730,N_3844);
and U4219 (N_4219,N_3883,N_3832);
or U4220 (N_4220,N_3793,N_3803);
nand U4221 (N_4221,N_3817,N_3902);
nor U4222 (N_4222,N_3574,N_3976);
or U4223 (N_4223,N_3671,N_3738);
and U4224 (N_4224,N_3600,N_3512);
nor U4225 (N_4225,N_3518,N_3566);
and U4226 (N_4226,N_3734,N_3625);
nand U4227 (N_4227,N_3711,N_3847);
nand U4228 (N_4228,N_3702,N_3722);
nand U4229 (N_4229,N_3680,N_3546);
nor U4230 (N_4230,N_3986,N_3659);
nor U4231 (N_4231,N_3756,N_3919);
nand U4232 (N_4232,N_3997,N_3692);
nand U4233 (N_4233,N_3541,N_3759);
or U4234 (N_4234,N_3624,N_3639);
and U4235 (N_4235,N_3749,N_3854);
nand U4236 (N_4236,N_3524,N_3743);
nor U4237 (N_4237,N_3945,N_3895);
nand U4238 (N_4238,N_3603,N_3527);
nor U4239 (N_4239,N_3504,N_3934);
and U4240 (N_4240,N_3619,N_3843);
or U4241 (N_4241,N_3514,N_3861);
nor U4242 (N_4242,N_3933,N_3505);
nor U4243 (N_4243,N_3855,N_3764);
or U4244 (N_4244,N_3922,N_3757);
or U4245 (N_4245,N_3508,N_3656);
nand U4246 (N_4246,N_3567,N_3752);
nand U4247 (N_4247,N_3589,N_3664);
nor U4248 (N_4248,N_3632,N_3901);
nand U4249 (N_4249,N_3972,N_3869);
and U4250 (N_4250,N_3724,N_3516);
and U4251 (N_4251,N_3825,N_3931);
nor U4252 (N_4252,N_3894,N_3908);
nand U4253 (N_4253,N_3547,N_3771);
or U4254 (N_4254,N_3931,N_3691);
nor U4255 (N_4255,N_3535,N_3888);
nor U4256 (N_4256,N_3882,N_3632);
or U4257 (N_4257,N_3933,N_3789);
nand U4258 (N_4258,N_3744,N_3823);
nor U4259 (N_4259,N_3669,N_3502);
or U4260 (N_4260,N_3602,N_3946);
nor U4261 (N_4261,N_3515,N_3710);
nor U4262 (N_4262,N_3624,N_3961);
or U4263 (N_4263,N_3887,N_3743);
and U4264 (N_4264,N_3932,N_3677);
nor U4265 (N_4265,N_3900,N_3610);
or U4266 (N_4266,N_3569,N_3695);
nand U4267 (N_4267,N_3795,N_3880);
and U4268 (N_4268,N_3887,N_3557);
nor U4269 (N_4269,N_3700,N_3649);
nand U4270 (N_4270,N_3837,N_3836);
and U4271 (N_4271,N_3889,N_3862);
or U4272 (N_4272,N_3860,N_3547);
and U4273 (N_4273,N_3546,N_3768);
or U4274 (N_4274,N_3643,N_3776);
nand U4275 (N_4275,N_3671,N_3767);
nand U4276 (N_4276,N_3847,N_3899);
and U4277 (N_4277,N_3584,N_3994);
nor U4278 (N_4278,N_3578,N_3506);
nor U4279 (N_4279,N_3939,N_3918);
nor U4280 (N_4280,N_3629,N_3818);
nor U4281 (N_4281,N_3570,N_3730);
xor U4282 (N_4282,N_3927,N_3970);
nor U4283 (N_4283,N_3504,N_3571);
xor U4284 (N_4284,N_3964,N_3841);
nor U4285 (N_4285,N_3855,N_3859);
nand U4286 (N_4286,N_3784,N_3743);
nor U4287 (N_4287,N_3868,N_3633);
and U4288 (N_4288,N_3503,N_3928);
nand U4289 (N_4289,N_3934,N_3835);
nand U4290 (N_4290,N_3959,N_3629);
nand U4291 (N_4291,N_3938,N_3948);
or U4292 (N_4292,N_3900,N_3851);
and U4293 (N_4293,N_3818,N_3985);
or U4294 (N_4294,N_3779,N_3940);
or U4295 (N_4295,N_3508,N_3874);
nor U4296 (N_4296,N_3577,N_3694);
nand U4297 (N_4297,N_3968,N_3962);
or U4298 (N_4298,N_3510,N_3685);
or U4299 (N_4299,N_3783,N_3561);
nor U4300 (N_4300,N_3831,N_3825);
nor U4301 (N_4301,N_3920,N_3633);
and U4302 (N_4302,N_3944,N_3732);
xnor U4303 (N_4303,N_3686,N_3529);
and U4304 (N_4304,N_3719,N_3756);
or U4305 (N_4305,N_3521,N_3882);
nand U4306 (N_4306,N_3660,N_3900);
nor U4307 (N_4307,N_3948,N_3804);
and U4308 (N_4308,N_3649,N_3602);
and U4309 (N_4309,N_3690,N_3713);
nand U4310 (N_4310,N_3764,N_3680);
and U4311 (N_4311,N_3817,N_3775);
or U4312 (N_4312,N_3530,N_3773);
nor U4313 (N_4313,N_3871,N_3685);
or U4314 (N_4314,N_3719,N_3888);
nand U4315 (N_4315,N_3749,N_3722);
nor U4316 (N_4316,N_3867,N_3834);
or U4317 (N_4317,N_3733,N_3925);
nor U4318 (N_4318,N_3883,N_3704);
nand U4319 (N_4319,N_3568,N_3809);
nand U4320 (N_4320,N_3669,N_3692);
and U4321 (N_4321,N_3605,N_3880);
and U4322 (N_4322,N_3602,N_3623);
nor U4323 (N_4323,N_3752,N_3512);
and U4324 (N_4324,N_3988,N_3541);
nand U4325 (N_4325,N_3561,N_3695);
or U4326 (N_4326,N_3954,N_3727);
nor U4327 (N_4327,N_3654,N_3750);
nor U4328 (N_4328,N_3548,N_3720);
and U4329 (N_4329,N_3517,N_3728);
nor U4330 (N_4330,N_3767,N_3792);
or U4331 (N_4331,N_3814,N_3574);
and U4332 (N_4332,N_3733,N_3812);
nor U4333 (N_4333,N_3885,N_3739);
or U4334 (N_4334,N_3990,N_3946);
nand U4335 (N_4335,N_3968,N_3736);
nand U4336 (N_4336,N_3565,N_3842);
nor U4337 (N_4337,N_3539,N_3908);
or U4338 (N_4338,N_3627,N_3857);
nand U4339 (N_4339,N_3873,N_3765);
nor U4340 (N_4340,N_3643,N_3913);
or U4341 (N_4341,N_3740,N_3985);
or U4342 (N_4342,N_3962,N_3952);
nand U4343 (N_4343,N_3559,N_3605);
or U4344 (N_4344,N_3950,N_3800);
xnor U4345 (N_4345,N_3927,N_3813);
and U4346 (N_4346,N_3955,N_3820);
or U4347 (N_4347,N_3646,N_3633);
nand U4348 (N_4348,N_3522,N_3901);
or U4349 (N_4349,N_3983,N_3769);
or U4350 (N_4350,N_3617,N_3742);
nor U4351 (N_4351,N_3591,N_3792);
nor U4352 (N_4352,N_3943,N_3755);
or U4353 (N_4353,N_3825,N_3732);
and U4354 (N_4354,N_3607,N_3980);
or U4355 (N_4355,N_3664,N_3689);
nor U4356 (N_4356,N_3583,N_3525);
nor U4357 (N_4357,N_3729,N_3560);
nor U4358 (N_4358,N_3756,N_3538);
nand U4359 (N_4359,N_3695,N_3846);
or U4360 (N_4360,N_3778,N_3810);
nand U4361 (N_4361,N_3772,N_3595);
or U4362 (N_4362,N_3962,N_3706);
xnor U4363 (N_4363,N_3643,N_3549);
or U4364 (N_4364,N_3659,N_3584);
nand U4365 (N_4365,N_3898,N_3509);
and U4366 (N_4366,N_3506,N_3893);
or U4367 (N_4367,N_3725,N_3508);
and U4368 (N_4368,N_3636,N_3768);
and U4369 (N_4369,N_3990,N_3855);
nor U4370 (N_4370,N_3559,N_3777);
nor U4371 (N_4371,N_3931,N_3546);
nand U4372 (N_4372,N_3762,N_3744);
and U4373 (N_4373,N_3879,N_3537);
or U4374 (N_4374,N_3587,N_3584);
and U4375 (N_4375,N_3709,N_3699);
nand U4376 (N_4376,N_3791,N_3517);
nor U4377 (N_4377,N_3747,N_3671);
nand U4378 (N_4378,N_3606,N_3726);
and U4379 (N_4379,N_3535,N_3595);
and U4380 (N_4380,N_3968,N_3656);
or U4381 (N_4381,N_3793,N_3642);
or U4382 (N_4382,N_3981,N_3697);
nand U4383 (N_4383,N_3533,N_3590);
nand U4384 (N_4384,N_3853,N_3703);
nor U4385 (N_4385,N_3776,N_3762);
nand U4386 (N_4386,N_3552,N_3531);
and U4387 (N_4387,N_3871,N_3869);
and U4388 (N_4388,N_3631,N_3970);
nor U4389 (N_4389,N_3774,N_3833);
and U4390 (N_4390,N_3527,N_3786);
and U4391 (N_4391,N_3904,N_3541);
and U4392 (N_4392,N_3883,N_3567);
or U4393 (N_4393,N_3758,N_3986);
or U4394 (N_4394,N_3722,N_3920);
nor U4395 (N_4395,N_3852,N_3530);
nor U4396 (N_4396,N_3568,N_3876);
and U4397 (N_4397,N_3588,N_3729);
nand U4398 (N_4398,N_3947,N_3562);
or U4399 (N_4399,N_3782,N_3714);
nand U4400 (N_4400,N_3879,N_3734);
nand U4401 (N_4401,N_3646,N_3738);
nand U4402 (N_4402,N_3673,N_3602);
nor U4403 (N_4403,N_3584,N_3887);
or U4404 (N_4404,N_3791,N_3957);
nand U4405 (N_4405,N_3626,N_3902);
or U4406 (N_4406,N_3766,N_3641);
or U4407 (N_4407,N_3649,N_3834);
and U4408 (N_4408,N_3661,N_3722);
and U4409 (N_4409,N_3722,N_3560);
or U4410 (N_4410,N_3884,N_3975);
or U4411 (N_4411,N_3972,N_3525);
nand U4412 (N_4412,N_3671,N_3871);
or U4413 (N_4413,N_3695,N_3550);
nand U4414 (N_4414,N_3704,N_3695);
xor U4415 (N_4415,N_3948,N_3946);
nor U4416 (N_4416,N_3668,N_3757);
or U4417 (N_4417,N_3703,N_3696);
or U4418 (N_4418,N_3911,N_3933);
and U4419 (N_4419,N_3569,N_3812);
nor U4420 (N_4420,N_3886,N_3711);
or U4421 (N_4421,N_3545,N_3684);
and U4422 (N_4422,N_3662,N_3847);
or U4423 (N_4423,N_3643,N_3824);
nand U4424 (N_4424,N_3990,N_3676);
nand U4425 (N_4425,N_3920,N_3545);
nor U4426 (N_4426,N_3930,N_3985);
and U4427 (N_4427,N_3738,N_3975);
nor U4428 (N_4428,N_3606,N_3997);
and U4429 (N_4429,N_3528,N_3689);
and U4430 (N_4430,N_3623,N_3920);
and U4431 (N_4431,N_3674,N_3812);
nand U4432 (N_4432,N_3717,N_3824);
and U4433 (N_4433,N_3929,N_3564);
nor U4434 (N_4434,N_3701,N_3526);
and U4435 (N_4435,N_3992,N_3529);
or U4436 (N_4436,N_3664,N_3809);
nand U4437 (N_4437,N_3773,N_3973);
nand U4438 (N_4438,N_3646,N_3877);
and U4439 (N_4439,N_3535,N_3655);
nor U4440 (N_4440,N_3545,N_3541);
or U4441 (N_4441,N_3656,N_3987);
nand U4442 (N_4442,N_3972,N_3831);
nand U4443 (N_4443,N_3904,N_3975);
and U4444 (N_4444,N_3778,N_3843);
nor U4445 (N_4445,N_3932,N_3850);
nor U4446 (N_4446,N_3583,N_3672);
nor U4447 (N_4447,N_3985,N_3741);
nor U4448 (N_4448,N_3923,N_3783);
nand U4449 (N_4449,N_3803,N_3841);
and U4450 (N_4450,N_3880,N_3694);
or U4451 (N_4451,N_3588,N_3567);
or U4452 (N_4452,N_3558,N_3592);
or U4453 (N_4453,N_3827,N_3609);
and U4454 (N_4454,N_3524,N_3615);
and U4455 (N_4455,N_3979,N_3525);
and U4456 (N_4456,N_3971,N_3504);
nor U4457 (N_4457,N_3757,N_3509);
or U4458 (N_4458,N_3826,N_3772);
or U4459 (N_4459,N_3943,N_3791);
and U4460 (N_4460,N_3692,N_3918);
and U4461 (N_4461,N_3581,N_3732);
and U4462 (N_4462,N_3962,N_3645);
nor U4463 (N_4463,N_3833,N_3661);
nor U4464 (N_4464,N_3915,N_3747);
and U4465 (N_4465,N_3627,N_3909);
nor U4466 (N_4466,N_3556,N_3787);
or U4467 (N_4467,N_3795,N_3842);
nor U4468 (N_4468,N_3637,N_3911);
nor U4469 (N_4469,N_3886,N_3737);
nand U4470 (N_4470,N_3624,N_3670);
and U4471 (N_4471,N_3662,N_3603);
and U4472 (N_4472,N_3575,N_3935);
nor U4473 (N_4473,N_3943,N_3996);
nor U4474 (N_4474,N_3550,N_3937);
or U4475 (N_4475,N_3648,N_3646);
nand U4476 (N_4476,N_3724,N_3660);
and U4477 (N_4477,N_3521,N_3614);
nor U4478 (N_4478,N_3624,N_3630);
nand U4479 (N_4479,N_3554,N_3688);
nor U4480 (N_4480,N_3907,N_3510);
or U4481 (N_4481,N_3999,N_3708);
nor U4482 (N_4482,N_3995,N_3562);
nor U4483 (N_4483,N_3936,N_3811);
nand U4484 (N_4484,N_3758,N_3970);
nand U4485 (N_4485,N_3685,N_3590);
xor U4486 (N_4486,N_3542,N_3734);
or U4487 (N_4487,N_3561,N_3935);
and U4488 (N_4488,N_3773,N_3711);
nor U4489 (N_4489,N_3775,N_3864);
nor U4490 (N_4490,N_3744,N_3887);
or U4491 (N_4491,N_3820,N_3533);
and U4492 (N_4492,N_3636,N_3528);
nand U4493 (N_4493,N_3829,N_3688);
nand U4494 (N_4494,N_3647,N_3874);
nand U4495 (N_4495,N_3664,N_3746);
or U4496 (N_4496,N_3603,N_3899);
and U4497 (N_4497,N_3946,N_3589);
or U4498 (N_4498,N_3759,N_3874);
and U4499 (N_4499,N_3564,N_3901);
or U4500 (N_4500,N_4219,N_4126);
nand U4501 (N_4501,N_4214,N_4488);
or U4502 (N_4502,N_4484,N_4270);
and U4503 (N_4503,N_4168,N_4090);
nor U4504 (N_4504,N_4059,N_4338);
and U4505 (N_4505,N_4404,N_4436);
or U4506 (N_4506,N_4023,N_4200);
nor U4507 (N_4507,N_4376,N_4105);
nor U4508 (N_4508,N_4045,N_4055);
nor U4509 (N_4509,N_4493,N_4463);
nor U4510 (N_4510,N_4032,N_4448);
nand U4511 (N_4511,N_4497,N_4489);
and U4512 (N_4512,N_4442,N_4135);
nor U4513 (N_4513,N_4389,N_4157);
and U4514 (N_4514,N_4264,N_4085);
nor U4515 (N_4515,N_4426,N_4277);
nand U4516 (N_4516,N_4378,N_4445);
or U4517 (N_4517,N_4474,N_4349);
nand U4518 (N_4518,N_4464,N_4098);
nor U4519 (N_4519,N_4165,N_4314);
or U4520 (N_4520,N_4174,N_4281);
or U4521 (N_4521,N_4400,N_4272);
and U4522 (N_4522,N_4038,N_4225);
nor U4523 (N_4523,N_4242,N_4339);
or U4524 (N_4524,N_4235,N_4461);
nand U4525 (N_4525,N_4186,N_4382);
nand U4526 (N_4526,N_4472,N_4063);
nor U4527 (N_4527,N_4154,N_4030);
and U4528 (N_4528,N_4170,N_4124);
or U4529 (N_4529,N_4470,N_4097);
nand U4530 (N_4530,N_4304,N_4428);
or U4531 (N_4531,N_4251,N_4300);
nand U4532 (N_4532,N_4054,N_4106);
nor U4533 (N_4533,N_4273,N_4358);
or U4534 (N_4534,N_4469,N_4140);
nand U4535 (N_4535,N_4475,N_4401);
nand U4536 (N_4536,N_4323,N_4375);
or U4537 (N_4537,N_4341,N_4353);
and U4538 (N_4538,N_4485,N_4095);
nor U4539 (N_4539,N_4016,N_4333);
or U4540 (N_4540,N_4012,N_4262);
nor U4541 (N_4541,N_4177,N_4076);
or U4542 (N_4542,N_4245,N_4259);
and U4543 (N_4543,N_4418,N_4433);
and U4544 (N_4544,N_4176,N_4394);
nand U4545 (N_4545,N_4241,N_4355);
or U4546 (N_4546,N_4381,N_4018);
nor U4547 (N_4547,N_4388,N_4073);
nand U4548 (N_4548,N_4374,N_4123);
nand U4549 (N_4549,N_4197,N_4454);
nand U4550 (N_4550,N_4346,N_4396);
nor U4551 (N_4551,N_4002,N_4099);
nand U4552 (N_4552,N_4253,N_4222);
nor U4553 (N_4553,N_4424,N_4078);
nand U4554 (N_4554,N_4212,N_4194);
and U4555 (N_4555,N_4092,N_4319);
and U4556 (N_4556,N_4109,N_4243);
nor U4557 (N_4557,N_4004,N_4148);
nand U4558 (N_4558,N_4289,N_4334);
nand U4559 (N_4559,N_4008,N_4340);
nand U4560 (N_4560,N_4440,N_4216);
nand U4561 (N_4561,N_4064,N_4288);
nor U4562 (N_4562,N_4133,N_4482);
nand U4563 (N_4563,N_4301,N_4034);
nor U4564 (N_4564,N_4127,N_4129);
nor U4565 (N_4565,N_4258,N_4263);
nand U4566 (N_4566,N_4326,N_4081);
or U4567 (N_4567,N_4383,N_4450);
nor U4568 (N_4568,N_4083,N_4208);
and U4569 (N_4569,N_4217,N_4025);
or U4570 (N_4570,N_4006,N_4011);
or U4571 (N_4571,N_4101,N_4250);
nor U4572 (N_4572,N_4047,N_4000);
nor U4573 (N_4573,N_4211,N_4395);
and U4574 (N_4574,N_4456,N_4020);
nand U4575 (N_4575,N_4184,N_4466);
nor U4576 (N_4576,N_4439,N_4316);
nor U4577 (N_4577,N_4056,N_4185);
nand U4578 (N_4578,N_4048,N_4294);
nand U4579 (N_4579,N_4427,N_4136);
or U4580 (N_4580,N_4380,N_4271);
nand U4581 (N_4581,N_4192,N_4224);
or U4582 (N_4582,N_4147,N_4026);
or U4583 (N_4583,N_4213,N_4221);
and U4584 (N_4584,N_4368,N_4308);
or U4585 (N_4585,N_4286,N_4033);
nand U4586 (N_4586,N_4332,N_4142);
nand U4587 (N_4587,N_4207,N_4306);
and U4588 (N_4588,N_4416,N_4494);
nor U4589 (N_4589,N_4209,N_4202);
and U4590 (N_4590,N_4093,N_4462);
nand U4591 (N_4591,N_4255,N_4405);
or U4592 (N_4592,N_4287,N_4290);
and U4593 (N_4593,N_4188,N_4412);
nand U4594 (N_4594,N_4161,N_4166);
nor U4595 (N_4595,N_4422,N_4195);
or U4596 (N_4596,N_4429,N_4162);
nand U4597 (N_4597,N_4385,N_4490);
or U4598 (N_4598,N_4043,N_4163);
and U4599 (N_4599,N_4201,N_4317);
and U4600 (N_4600,N_4451,N_4116);
nor U4601 (N_4601,N_4069,N_4363);
and U4602 (N_4602,N_4228,N_4292);
nor U4603 (N_4603,N_4117,N_4402);
and U4604 (N_4604,N_4437,N_4128);
and U4605 (N_4605,N_4238,N_4397);
or U4606 (N_4606,N_4231,N_4313);
or U4607 (N_4607,N_4080,N_4110);
nand U4608 (N_4608,N_4421,N_4443);
and U4609 (N_4609,N_4114,N_4203);
and U4610 (N_4610,N_4041,N_4302);
or U4611 (N_4611,N_4199,N_4303);
and U4612 (N_4612,N_4060,N_4134);
nor U4613 (N_4613,N_4257,N_4392);
or U4614 (N_4614,N_4491,N_4345);
nor U4615 (N_4615,N_4122,N_4495);
or U4616 (N_4616,N_4321,N_4407);
nand U4617 (N_4617,N_4130,N_4252);
or U4618 (N_4618,N_4285,N_4434);
nor U4619 (N_4619,N_4236,N_4145);
and U4620 (N_4620,N_4307,N_4352);
nand U4621 (N_4621,N_4343,N_4296);
or U4622 (N_4622,N_4467,N_4248);
and U4623 (N_4623,N_4377,N_4379);
nand U4624 (N_4624,N_4137,N_4279);
nor U4625 (N_4625,N_4205,N_4246);
nand U4626 (N_4626,N_4138,N_4172);
nor U4627 (N_4627,N_4067,N_4232);
nor U4628 (N_4628,N_4113,N_4100);
or U4629 (N_4629,N_4373,N_4031);
nand U4630 (N_4630,N_4015,N_4473);
nand U4631 (N_4631,N_4049,N_4223);
nand U4632 (N_4632,N_4365,N_4075);
nand U4633 (N_4633,N_4053,N_4387);
nand U4634 (N_4634,N_4274,N_4447);
nor U4635 (N_4635,N_4087,N_4282);
nand U4636 (N_4636,N_4143,N_4438);
nand U4637 (N_4637,N_4149,N_4268);
nand U4638 (N_4638,N_4318,N_4329);
or U4639 (N_4639,N_4226,N_4362);
nand U4640 (N_4640,N_4039,N_4283);
nor U4641 (N_4641,N_4360,N_4139);
xnor U4642 (N_4642,N_4052,N_4249);
or U4643 (N_4643,N_4057,N_4411);
or U4644 (N_4644,N_4084,N_4210);
and U4645 (N_4645,N_4452,N_4417);
or U4646 (N_4646,N_4311,N_4029);
or U4647 (N_4647,N_4089,N_4435);
nand U4648 (N_4648,N_4327,N_4146);
nand U4649 (N_4649,N_4050,N_4071);
and U4650 (N_4650,N_4414,N_4091);
or U4651 (N_4651,N_4419,N_4423);
or U4652 (N_4652,N_4022,N_4441);
and U4653 (N_4653,N_4010,N_4372);
and U4654 (N_4654,N_4468,N_4309);
and U4655 (N_4655,N_4171,N_4390);
or U4656 (N_4656,N_4460,N_4028);
nor U4657 (N_4657,N_4481,N_4062);
nor U4658 (N_4658,N_4027,N_4183);
or U4659 (N_4659,N_4458,N_4112);
nor U4660 (N_4660,N_4167,N_4103);
or U4661 (N_4661,N_4227,N_4477);
or U4662 (N_4662,N_4320,N_4131);
and U4663 (N_4663,N_4266,N_4275);
nand U4664 (N_4664,N_4348,N_4393);
nor U4665 (N_4665,N_4189,N_4111);
or U4666 (N_4666,N_4361,N_4384);
and U4667 (N_4667,N_4061,N_4187);
nor U4668 (N_4668,N_4206,N_4230);
nor U4669 (N_4669,N_4449,N_4175);
or U4670 (N_4670,N_4074,N_4324);
nand U4671 (N_4671,N_4102,N_4386);
nor U4672 (N_4672,N_4001,N_4218);
nand U4673 (N_4673,N_4003,N_4325);
nor U4674 (N_4674,N_4121,N_4181);
or U4675 (N_4675,N_4337,N_4403);
and U4676 (N_4676,N_4009,N_4391);
or U4677 (N_4677,N_4088,N_4068);
and U4678 (N_4678,N_4237,N_4359);
nand U4679 (N_4679,N_4180,N_4369);
and U4680 (N_4680,N_4155,N_4005);
nor U4681 (N_4681,N_4125,N_4370);
and U4682 (N_4682,N_4420,N_4265);
and U4683 (N_4683,N_4159,N_4158);
nand U4684 (N_4684,N_4169,N_4364);
and U4685 (N_4685,N_4153,N_4107);
or U4686 (N_4686,N_4017,N_4179);
nor U4687 (N_4687,N_4086,N_4024);
or U4688 (N_4688,N_4471,N_4476);
and U4689 (N_4689,N_4310,N_4173);
and U4690 (N_4690,N_4492,N_4425);
and U4691 (N_4691,N_4079,N_4284);
or U4692 (N_4692,N_4409,N_4444);
and U4693 (N_4693,N_4351,N_4280);
nand U4694 (N_4694,N_4479,N_4036);
nand U4695 (N_4695,N_4058,N_4413);
and U4696 (N_4696,N_4120,N_4478);
or U4697 (N_4697,N_4335,N_4104);
and U4698 (N_4698,N_4406,N_4256);
nor U4699 (N_4699,N_4156,N_4164);
nor U4700 (N_4700,N_4051,N_4037);
nand U4701 (N_4701,N_4046,N_4261);
nand U4702 (N_4702,N_4328,N_4293);
or U4703 (N_4703,N_4215,N_4331);
or U4704 (N_4704,N_4042,N_4072);
or U4705 (N_4705,N_4496,N_4118);
nor U4706 (N_4706,N_4410,N_4141);
or U4707 (N_4707,N_4007,N_4070);
nand U4708 (N_4708,N_4269,N_4297);
nand U4709 (N_4709,N_4196,N_4182);
or U4710 (N_4710,N_4204,N_4193);
nor U4711 (N_4711,N_4298,N_4239);
or U4712 (N_4712,N_4066,N_4035);
nand U4713 (N_4713,N_4160,N_4299);
nor U4714 (N_4714,N_4019,N_4347);
nor U4715 (N_4715,N_4357,N_4350);
nand U4716 (N_4716,N_4498,N_4178);
nand U4717 (N_4717,N_4152,N_4480);
nor U4718 (N_4718,N_4446,N_4330);
nand U4719 (N_4719,N_4094,N_4014);
or U4720 (N_4720,N_4315,N_4233);
nor U4721 (N_4721,N_4432,N_4415);
or U4722 (N_4722,N_4244,N_4312);
nand U4723 (N_4723,N_4344,N_4198);
nor U4724 (N_4724,N_4096,N_4115);
nand U4725 (N_4725,N_4366,N_4234);
or U4726 (N_4726,N_4021,N_4291);
or U4727 (N_4727,N_4151,N_4254);
and U4728 (N_4728,N_4399,N_4431);
or U4729 (N_4729,N_4305,N_4220);
nor U4730 (N_4730,N_4336,N_4459);
nor U4731 (N_4731,N_4082,N_4371);
and U4732 (N_4732,N_4044,N_4077);
nor U4733 (N_4733,N_4267,N_4144);
or U4734 (N_4734,N_4150,N_4398);
nor U4735 (N_4735,N_4065,N_4276);
nor U4736 (N_4736,N_4408,N_4457);
nor U4737 (N_4737,N_4322,N_4455);
and U4738 (N_4738,N_4499,N_4486);
and U4739 (N_4739,N_4013,N_4040);
nor U4740 (N_4740,N_4132,N_4247);
xnor U4741 (N_4741,N_4229,N_4260);
nor U4742 (N_4742,N_4483,N_4465);
nand U4743 (N_4743,N_4430,N_4354);
nor U4744 (N_4744,N_4487,N_4191);
and U4745 (N_4745,N_4240,N_4453);
xor U4746 (N_4746,N_4278,N_4367);
nand U4747 (N_4747,N_4119,N_4342);
nor U4748 (N_4748,N_4295,N_4190);
nand U4749 (N_4749,N_4356,N_4108);
or U4750 (N_4750,N_4109,N_4433);
nand U4751 (N_4751,N_4179,N_4343);
or U4752 (N_4752,N_4097,N_4343);
and U4753 (N_4753,N_4418,N_4215);
nand U4754 (N_4754,N_4362,N_4304);
or U4755 (N_4755,N_4374,N_4499);
nand U4756 (N_4756,N_4449,N_4266);
nand U4757 (N_4757,N_4209,N_4207);
or U4758 (N_4758,N_4171,N_4463);
nor U4759 (N_4759,N_4042,N_4376);
nand U4760 (N_4760,N_4411,N_4040);
or U4761 (N_4761,N_4020,N_4089);
nor U4762 (N_4762,N_4191,N_4081);
nand U4763 (N_4763,N_4125,N_4434);
or U4764 (N_4764,N_4297,N_4017);
and U4765 (N_4765,N_4189,N_4166);
nor U4766 (N_4766,N_4177,N_4427);
and U4767 (N_4767,N_4119,N_4240);
nor U4768 (N_4768,N_4457,N_4029);
nor U4769 (N_4769,N_4268,N_4026);
and U4770 (N_4770,N_4497,N_4019);
or U4771 (N_4771,N_4417,N_4136);
and U4772 (N_4772,N_4138,N_4355);
and U4773 (N_4773,N_4000,N_4329);
nor U4774 (N_4774,N_4480,N_4030);
or U4775 (N_4775,N_4112,N_4421);
or U4776 (N_4776,N_4034,N_4384);
and U4777 (N_4777,N_4007,N_4117);
nand U4778 (N_4778,N_4036,N_4053);
or U4779 (N_4779,N_4432,N_4349);
nor U4780 (N_4780,N_4066,N_4111);
or U4781 (N_4781,N_4282,N_4278);
nor U4782 (N_4782,N_4124,N_4347);
and U4783 (N_4783,N_4076,N_4023);
and U4784 (N_4784,N_4211,N_4457);
nor U4785 (N_4785,N_4358,N_4241);
or U4786 (N_4786,N_4449,N_4427);
or U4787 (N_4787,N_4166,N_4091);
and U4788 (N_4788,N_4116,N_4255);
nand U4789 (N_4789,N_4380,N_4447);
nand U4790 (N_4790,N_4350,N_4329);
and U4791 (N_4791,N_4434,N_4010);
or U4792 (N_4792,N_4257,N_4296);
nor U4793 (N_4793,N_4455,N_4098);
and U4794 (N_4794,N_4214,N_4460);
nor U4795 (N_4795,N_4416,N_4277);
nor U4796 (N_4796,N_4466,N_4249);
nor U4797 (N_4797,N_4190,N_4216);
and U4798 (N_4798,N_4385,N_4232);
or U4799 (N_4799,N_4421,N_4392);
or U4800 (N_4800,N_4079,N_4215);
nand U4801 (N_4801,N_4311,N_4223);
or U4802 (N_4802,N_4085,N_4173);
and U4803 (N_4803,N_4337,N_4261);
or U4804 (N_4804,N_4330,N_4138);
nor U4805 (N_4805,N_4212,N_4101);
or U4806 (N_4806,N_4423,N_4208);
or U4807 (N_4807,N_4082,N_4499);
and U4808 (N_4808,N_4466,N_4337);
nand U4809 (N_4809,N_4010,N_4399);
nor U4810 (N_4810,N_4110,N_4353);
nor U4811 (N_4811,N_4062,N_4384);
nor U4812 (N_4812,N_4405,N_4316);
or U4813 (N_4813,N_4351,N_4440);
or U4814 (N_4814,N_4269,N_4307);
or U4815 (N_4815,N_4079,N_4267);
xnor U4816 (N_4816,N_4038,N_4265);
and U4817 (N_4817,N_4219,N_4164);
nor U4818 (N_4818,N_4369,N_4117);
nand U4819 (N_4819,N_4152,N_4120);
and U4820 (N_4820,N_4382,N_4180);
or U4821 (N_4821,N_4346,N_4452);
nor U4822 (N_4822,N_4386,N_4225);
or U4823 (N_4823,N_4063,N_4396);
or U4824 (N_4824,N_4193,N_4357);
or U4825 (N_4825,N_4218,N_4165);
nor U4826 (N_4826,N_4113,N_4460);
and U4827 (N_4827,N_4253,N_4244);
or U4828 (N_4828,N_4309,N_4378);
nor U4829 (N_4829,N_4045,N_4336);
or U4830 (N_4830,N_4397,N_4246);
nor U4831 (N_4831,N_4328,N_4294);
or U4832 (N_4832,N_4195,N_4206);
and U4833 (N_4833,N_4354,N_4093);
or U4834 (N_4834,N_4137,N_4159);
nand U4835 (N_4835,N_4041,N_4400);
nor U4836 (N_4836,N_4121,N_4064);
nor U4837 (N_4837,N_4487,N_4063);
and U4838 (N_4838,N_4215,N_4496);
xnor U4839 (N_4839,N_4231,N_4018);
nor U4840 (N_4840,N_4134,N_4496);
and U4841 (N_4841,N_4155,N_4109);
and U4842 (N_4842,N_4410,N_4333);
or U4843 (N_4843,N_4219,N_4141);
nor U4844 (N_4844,N_4274,N_4275);
nor U4845 (N_4845,N_4431,N_4366);
xor U4846 (N_4846,N_4098,N_4284);
nand U4847 (N_4847,N_4151,N_4380);
and U4848 (N_4848,N_4174,N_4475);
and U4849 (N_4849,N_4185,N_4496);
nand U4850 (N_4850,N_4389,N_4415);
nand U4851 (N_4851,N_4473,N_4132);
nand U4852 (N_4852,N_4323,N_4080);
and U4853 (N_4853,N_4319,N_4154);
or U4854 (N_4854,N_4239,N_4086);
nor U4855 (N_4855,N_4181,N_4162);
nand U4856 (N_4856,N_4369,N_4216);
and U4857 (N_4857,N_4089,N_4101);
or U4858 (N_4858,N_4140,N_4009);
and U4859 (N_4859,N_4446,N_4216);
nand U4860 (N_4860,N_4393,N_4249);
nor U4861 (N_4861,N_4290,N_4088);
nor U4862 (N_4862,N_4318,N_4117);
nand U4863 (N_4863,N_4035,N_4172);
nor U4864 (N_4864,N_4170,N_4095);
and U4865 (N_4865,N_4442,N_4238);
or U4866 (N_4866,N_4256,N_4113);
or U4867 (N_4867,N_4238,N_4347);
and U4868 (N_4868,N_4499,N_4026);
or U4869 (N_4869,N_4467,N_4136);
nor U4870 (N_4870,N_4415,N_4319);
or U4871 (N_4871,N_4130,N_4234);
or U4872 (N_4872,N_4210,N_4191);
nor U4873 (N_4873,N_4355,N_4050);
nor U4874 (N_4874,N_4170,N_4378);
and U4875 (N_4875,N_4461,N_4232);
or U4876 (N_4876,N_4367,N_4111);
or U4877 (N_4877,N_4170,N_4275);
or U4878 (N_4878,N_4205,N_4442);
nand U4879 (N_4879,N_4033,N_4411);
nor U4880 (N_4880,N_4023,N_4293);
and U4881 (N_4881,N_4233,N_4263);
nand U4882 (N_4882,N_4159,N_4352);
and U4883 (N_4883,N_4206,N_4225);
or U4884 (N_4884,N_4034,N_4209);
and U4885 (N_4885,N_4354,N_4002);
and U4886 (N_4886,N_4126,N_4422);
and U4887 (N_4887,N_4415,N_4004);
nor U4888 (N_4888,N_4148,N_4358);
nand U4889 (N_4889,N_4444,N_4264);
or U4890 (N_4890,N_4262,N_4071);
or U4891 (N_4891,N_4068,N_4312);
nand U4892 (N_4892,N_4447,N_4276);
or U4893 (N_4893,N_4411,N_4466);
and U4894 (N_4894,N_4477,N_4002);
and U4895 (N_4895,N_4342,N_4391);
and U4896 (N_4896,N_4433,N_4345);
or U4897 (N_4897,N_4324,N_4342);
and U4898 (N_4898,N_4267,N_4369);
nor U4899 (N_4899,N_4406,N_4195);
nand U4900 (N_4900,N_4249,N_4422);
nand U4901 (N_4901,N_4049,N_4083);
and U4902 (N_4902,N_4308,N_4349);
xnor U4903 (N_4903,N_4054,N_4132);
nand U4904 (N_4904,N_4365,N_4106);
and U4905 (N_4905,N_4243,N_4312);
nand U4906 (N_4906,N_4164,N_4064);
or U4907 (N_4907,N_4077,N_4076);
nor U4908 (N_4908,N_4428,N_4172);
nand U4909 (N_4909,N_4376,N_4322);
nand U4910 (N_4910,N_4187,N_4468);
and U4911 (N_4911,N_4269,N_4292);
nor U4912 (N_4912,N_4073,N_4466);
nor U4913 (N_4913,N_4031,N_4256);
or U4914 (N_4914,N_4162,N_4076);
and U4915 (N_4915,N_4210,N_4268);
and U4916 (N_4916,N_4308,N_4114);
nand U4917 (N_4917,N_4460,N_4156);
and U4918 (N_4918,N_4150,N_4187);
nand U4919 (N_4919,N_4287,N_4201);
nor U4920 (N_4920,N_4082,N_4099);
and U4921 (N_4921,N_4252,N_4285);
nand U4922 (N_4922,N_4026,N_4014);
and U4923 (N_4923,N_4153,N_4226);
and U4924 (N_4924,N_4138,N_4350);
nor U4925 (N_4925,N_4299,N_4227);
or U4926 (N_4926,N_4203,N_4497);
or U4927 (N_4927,N_4378,N_4355);
nand U4928 (N_4928,N_4361,N_4367);
and U4929 (N_4929,N_4468,N_4460);
nor U4930 (N_4930,N_4032,N_4088);
and U4931 (N_4931,N_4189,N_4036);
nor U4932 (N_4932,N_4185,N_4277);
nand U4933 (N_4933,N_4224,N_4328);
or U4934 (N_4934,N_4313,N_4331);
nor U4935 (N_4935,N_4355,N_4139);
and U4936 (N_4936,N_4388,N_4167);
nor U4937 (N_4937,N_4009,N_4453);
or U4938 (N_4938,N_4108,N_4079);
and U4939 (N_4939,N_4259,N_4098);
and U4940 (N_4940,N_4220,N_4140);
nand U4941 (N_4941,N_4127,N_4243);
or U4942 (N_4942,N_4109,N_4173);
nor U4943 (N_4943,N_4423,N_4273);
and U4944 (N_4944,N_4057,N_4249);
or U4945 (N_4945,N_4487,N_4199);
nor U4946 (N_4946,N_4478,N_4154);
xnor U4947 (N_4947,N_4414,N_4140);
and U4948 (N_4948,N_4107,N_4276);
or U4949 (N_4949,N_4414,N_4070);
and U4950 (N_4950,N_4050,N_4387);
nand U4951 (N_4951,N_4130,N_4175);
or U4952 (N_4952,N_4032,N_4432);
and U4953 (N_4953,N_4003,N_4240);
or U4954 (N_4954,N_4148,N_4171);
nand U4955 (N_4955,N_4252,N_4027);
nor U4956 (N_4956,N_4137,N_4140);
and U4957 (N_4957,N_4308,N_4077);
nor U4958 (N_4958,N_4444,N_4473);
nor U4959 (N_4959,N_4310,N_4047);
or U4960 (N_4960,N_4237,N_4432);
nor U4961 (N_4961,N_4446,N_4075);
nand U4962 (N_4962,N_4424,N_4296);
nand U4963 (N_4963,N_4027,N_4001);
nor U4964 (N_4964,N_4151,N_4416);
nand U4965 (N_4965,N_4448,N_4491);
and U4966 (N_4966,N_4060,N_4125);
and U4967 (N_4967,N_4284,N_4058);
or U4968 (N_4968,N_4012,N_4261);
or U4969 (N_4969,N_4217,N_4397);
or U4970 (N_4970,N_4101,N_4200);
nor U4971 (N_4971,N_4443,N_4203);
and U4972 (N_4972,N_4240,N_4176);
and U4973 (N_4973,N_4096,N_4221);
or U4974 (N_4974,N_4105,N_4418);
and U4975 (N_4975,N_4153,N_4013);
and U4976 (N_4976,N_4226,N_4003);
or U4977 (N_4977,N_4492,N_4347);
xor U4978 (N_4978,N_4015,N_4282);
nand U4979 (N_4979,N_4349,N_4009);
nor U4980 (N_4980,N_4219,N_4182);
nor U4981 (N_4981,N_4462,N_4297);
nand U4982 (N_4982,N_4022,N_4214);
or U4983 (N_4983,N_4029,N_4190);
and U4984 (N_4984,N_4059,N_4236);
nand U4985 (N_4985,N_4083,N_4074);
or U4986 (N_4986,N_4127,N_4232);
or U4987 (N_4987,N_4058,N_4056);
or U4988 (N_4988,N_4213,N_4376);
nor U4989 (N_4989,N_4321,N_4386);
nand U4990 (N_4990,N_4033,N_4250);
nor U4991 (N_4991,N_4100,N_4129);
and U4992 (N_4992,N_4279,N_4110);
nor U4993 (N_4993,N_4381,N_4039);
nand U4994 (N_4994,N_4399,N_4340);
nand U4995 (N_4995,N_4160,N_4342);
and U4996 (N_4996,N_4479,N_4403);
and U4997 (N_4997,N_4257,N_4065);
or U4998 (N_4998,N_4128,N_4384);
or U4999 (N_4999,N_4192,N_4137);
nand UO_0 (O_0,N_4680,N_4938);
nor UO_1 (O_1,N_4587,N_4775);
nand UO_2 (O_2,N_4980,N_4918);
nand UO_3 (O_3,N_4895,N_4771);
nor UO_4 (O_4,N_4612,N_4844);
and UO_5 (O_5,N_4764,N_4580);
or UO_6 (O_6,N_4576,N_4598);
nor UO_7 (O_7,N_4558,N_4990);
or UO_8 (O_8,N_4661,N_4744);
and UO_9 (O_9,N_4815,N_4782);
and UO_10 (O_10,N_4953,N_4541);
nor UO_11 (O_11,N_4684,N_4718);
or UO_12 (O_12,N_4685,N_4769);
nor UO_13 (O_13,N_4637,N_4523);
nand UO_14 (O_14,N_4968,N_4539);
nor UO_15 (O_15,N_4935,N_4682);
or UO_16 (O_16,N_4556,N_4912);
and UO_17 (O_17,N_4675,N_4843);
nand UO_18 (O_18,N_4588,N_4826);
or UO_19 (O_19,N_4616,N_4805);
nor UO_20 (O_20,N_4985,N_4631);
nand UO_21 (O_21,N_4821,N_4641);
or UO_22 (O_22,N_4544,N_4596);
or UO_23 (O_23,N_4929,N_4621);
and UO_24 (O_24,N_4960,N_4525);
nor UO_25 (O_25,N_4885,N_4836);
nand UO_26 (O_26,N_4794,N_4873);
or UO_27 (O_27,N_4638,N_4811);
and UO_28 (O_28,N_4984,N_4550);
or UO_29 (O_29,N_4948,N_4939);
and UO_30 (O_30,N_4973,N_4781);
nor UO_31 (O_31,N_4878,N_4795);
nand UO_32 (O_32,N_4609,N_4864);
nand UO_33 (O_33,N_4733,N_4704);
nor UO_34 (O_34,N_4942,N_4943);
nand UO_35 (O_35,N_4772,N_4709);
nand UO_36 (O_36,N_4854,N_4954);
nand UO_37 (O_37,N_4933,N_4664);
nand UO_38 (O_38,N_4650,N_4966);
and UO_39 (O_39,N_4894,N_4976);
or UO_40 (O_40,N_4725,N_4837);
and UO_41 (O_41,N_4698,N_4535);
and UO_42 (O_42,N_4803,N_4625);
or UO_43 (O_43,N_4762,N_4917);
and UO_44 (O_44,N_4571,N_4706);
nand UO_45 (O_45,N_4840,N_4770);
nor UO_46 (O_46,N_4613,N_4652);
nand UO_47 (O_47,N_4737,N_4947);
nor UO_48 (O_48,N_4866,N_4982);
and UO_49 (O_49,N_4622,N_4699);
nand UO_50 (O_50,N_4624,N_4869);
or UO_51 (O_51,N_4888,N_4986);
nand UO_52 (O_52,N_4841,N_4537);
xnor UO_53 (O_53,N_4785,N_4940);
or UO_54 (O_54,N_4883,N_4830);
or UO_55 (O_55,N_4790,N_4904);
and UO_56 (O_56,N_4767,N_4502);
nand UO_57 (O_57,N_4672,N_4657);
nor UO_58 (O_58,N_4521,N_4635);
or UO_59 (O_59,N_4529,N_4500);
nand UO_60 (O_60,N_4681,N_4530);
nand UO_61 (O_61,N_4879,N_4552);
nand UO_62 (O_62,N_4952,N_4505);
nand UO_63 (O_63,N_4582,N_4784);
nor UO_64 (O_64,N_4850,N_4755);
nand UO_65 (O_65,N_4645,N_4723);
nor UO_66 (O_66,N_4597,N_4632);
nand UO_67 (O_67,N_4633,N_4872);
or UO_68 (O_68,N_4881,N_4614);
nor UO_69 (O_69,N_4858,N_4579);
nor UO_70 (O_70,N_4691,N_4676);
and UO_71 (O_71,N_4687,N_4574);
or UO_72 (O_72,N_4860,N_4928);
nand UO_73 (O_73,N_4907,N_4729);
xnor UO_74 (O_74,N_4916,N_4651);
nor UO_75 (O_75,N_4848,N_4889);
or UO_76 (O_76,N_4833,N_4644);
xnor UO_77 (O_77,N_4604,N_4874);
and UO_78 (O_78,N_4668,N_4827);
and UO_79 (O_79,N_4893,N_4654);
nand UO_80 (O_80,N_4787,N_4665);
or UO_81 (O_81,N_4591,N_4886);
or UO_82 (O_82,N_4969,N_4822);
nand UO_83 (O_83,N_4835,N_4527);
nand UO_84 (O_84,N_4540,N_4802);
nand UO_85 (O_85,N_4719,N_4807);
nor UO_86 (O_86,N_4640,N_4825);
and UO_87 (O_87,N_4964,N_4583);
nor UO_88 (O_88,N_4518,N_4642);
nor UO_89 (O_89,N_4839,N_4511);
nand UO_90 (O_90,N_4779,N_4958);
nand UO_91 (O_91,N_4610,N_4615);
nor UO_92 (O_92,N_4573,N_4814);
or UO_93 (O_93,N_4504,N_4713);
and UO_94 (O_94,N_4568,N_4600);
and UO_95 (O_95,N_4849,N_4914);
nor UO_96 (O_96,N_4570,N_4546);
or UO_97 (O_97,N_4659,N_4910);
or UO_98 (O_98,N_4602,N_4962);
and UO_99 (O_99,N_4520,N_4722);
nor UO_100 (O_100,N_4920,N_4901);
or UO_101 (O_101,N_4512,N_4911);
or UO_102 (O_102,N_4798,N_4533);
nand UO_103 (O_103,N_4908,N_4710);
nand UO_104 (O_104,N_4741,N_4996);
nand UO_105 (O_105,N_4743,N_4619);
nand UO_106 (O_106,N_4561,N_4617);
nand UO_107 (O_107,N_4824,N_4995);
and UO_108 (O_108,N_4763,N_4788);
or UO_109 (O_109,N_4750,N_4845);
nor UO_110 (O_110,N_4847,N_4630);
nor UO_111 (O_111,N_4646,N_4834);
or UO_112 (O_112,N_4891,N_4581);
or UO_113 (O_113,N_4932,N_4892);
and UO_114 (O_114,N_4851,N_4700);
or UO_115 (O_115,N_4658,N_4522);
nor UO_116 (O_116,N_4753,N_4857);
nor UO_117 (O_117,N_4515,N_4590);
and UO_118 (O_118,N_4697,N_4934);
nand UO_119 (O_119,N_4946,N_4514);
nand UO_120 (O_120,N_4711,N_4890);
or UO_121 (O_121,N_4856,N_4909);
nor UO_122 (O_122,N_4993,N_4861);
or UO_123 (O_123,N_4792,N_4717);
nand UO_124 (O_124,N_4760,N_4662);
or UO_125 (O_125,N_4715,N_4905);
nor UO_126 (O_126,N_4673,N_4551);
nand UO_127 (O_127,N_4670,N_4941);
nor UO_128 (O_128,N_4585,N_4870);
nand UO_129 (O_129,N_4999,N_4705);
nor UO_130 (O_130,N_4859,N_4877);
or UO_131 (O_131,N_4620,N_4832);
nor UO_132 (O_132,N_4906,N_4693);
nand UO_133 (O_133,N_4863,N_4963);
or UO_134 (O_134,N_4897,N_4528);
or UO_135 (O_135,N_4746,N_4818);
nor UO_136 (O_136,N_4876,N_4749);
nor UO_137 (O_137,N_4677,N_4507);
and UO_138 (O_138,N_4970,N_4606);
nand UO_139 (O_139,N_4819,N_4936);
nand UO_140 (O_140,N_4768,N_4643);
and UO_141 (O_141,N_4738,N_4951);
nand UO_142 (O_142,N_4628,N_4971);
and UO_143 (O_143,N_4801,N_4660);
and UO_144 (O_144,N_4517,N_4816);
nand UO_145 (O_145,N_4708,N_4666);
nand UO_146 (O_146,N_4930,N_4862);
nand UO_147 (O_147,N_4742,N_4875);
or UO_148 (O_148,N_4577,N_4747);
and UO_149 (O_149,N_4967,N_4538);
nor UO_150 (O_150,N_4957,N_4601);
nand UO_151 (O_151,N_4789,N_4532);
and UO_152 (O_152,N_4689,N_4548);
nor UO_153 (O_153,N_4627,N_4842);
nand UO_154 (O_154,N_4989,N_4626);
nor UO_155 (O_155,N_4757,N_4567);
or UO_156 (O_156,N_4926,N_4956);
and UO_157 (O_157,N_4846,N_4900);
or UO_158 (O_158,N_4688,N_4778);
nand UO_159 (O_159,N_4994,N_4902);
and UO_160 (O_160,N_4783,N_4636);
nand UO_161 (O_161,N_4656,N_4503);
or UO_162 (O_162,N_4524,N_4671);
or UO_163 (O_163,N_4647,N_4707);
or UO_164 (O_164,N_4562,N_4578);
nor UO_165 (O_165,N_4748,N_4634);
nor UO_166 (O_166,N_4734,N_4828);
nand UO_167 (O_167,N_4542,N_4829);
nand UO_168 (O_168,N_4739,N_4509);
nand UO_169 (O_169,N_4800,N_4608);
or UO_170 (O_170,N_4751,N_4611);
or UO_171 (O_171,N_4547,N_4797);
nor UO_172 (O_172,N_4534,N_4761);
or UO_173 (O_173,N_4678,N_4865);
or UO_174 (O_174,N_4983,N_4721);
or UO_175 (O_175,N_4603,N_4720);
xnor UO_176 (O_176,N_4852,N_4786);
and UO_177 (O_177,N_4975,N_4868);
and UO_178 (O_178,N_4730,N_4959);
nand UO_179 (O_179,N_4736,N_4991);
nand UO_180 (O_180,N_4649,N_4855);
and UO_181 (O_181,N_4618,N_4988);
or UO_182 (O_182,N_4508,N_4607);
nand UO_183 (O_183,N_4766,N_4683);
nand UO_184 (O_184,N_4978,N_4882);
nor UO_185 (O_185,N_4648,N_4853);
nor UO_186 (O_186,N_4553,N_4732);
and UO_187 (O_187,N_4563,N_4997);
and UO_188 (O_188,N_4831,N_4667);
or UO_189 (O_189,N_4773,N_4549);
nor UO_190 (O_190,N_4961,N_4898);
nand UO_191 (O_191,N_4589,N_4663);
or UO_192 (O_192,N_4925,N_4728);
or UO_193 (O_193,N_4812,N_4545);
or UO_194 (O_194,N_4560,N_4922);
nand UO_195 (O_195,N_4896,N_4655);
or UO_196 (O_196,N_4595,N_4605);
and UO_197 (O_197,N_4526,N_4593);
nor UO_198 (O_198,N_4899,N_4793);
nor UO_199 (O_199,N_4931,N_4752);
nor UO_200 (O_200,N_4998,N_4565);
nand UO_201 (O_201,N_4726,N_4813);
nor UO_202 (O_202,N_4809,N_4927);
or UO_203 (O_203,N_4937,N_4838);
or UO_204 (O_204,N_4740,N_4731);
or UO_205 (O_205,N_4955,N_4759);
nand UO_206 (O_206,N_4880,N_4765);
nor UO_207 (O_207,N_4694,N_4594);
or UO_208 (O_208,N_4806,N_4965);
nand UO_209 (O_209,N_4913,N_4516);
or UO_210 (O_210,N_4592,N_4776);
nor UO_211 (O_211,N_4714,N_4695);
xnor UO_212 (O_212,N_4674,N_4745);
nand UO_213 (O_213,N_4777,N_4977);
or UO_214 (O_214,N_4510,N_4915);
nor UO_215 (O_215,N_4799,N_4629);
nand UO_216 (O_216,N_4808,N_4756);
or UO_217 (O_217,N_4690,N_4554);
and UO_218 (O_218,N_4944,N_4623);
nor UO_219 (O_219,N_4702,N_4557);
nand UO_220 (O_220,N_4653,N_4712);
and UO_221 (O_221,N_4919,N_4639);
and UO_222 (O_222,N_4584,N_4531);
nor UO_223 (O_223,N_4804,N_4735);
and UO_224 (O_224,N_4923,N_4513);
and UO_225 (O_225,N_4501,N_4586);
and UO_226 (O_226,N_4703,N_4903);
nor UO_227 (O_227,N_4754,N_4575);
nor UO_228 (O_228,N_4887,N_4987);
nor UO_229 (O_229,N_4572,N_4669);
or UO_230 (O_230,N_4823,N_4796);
and UO_231 (O_231,N_4724,N_4727);
nand UO_232 (O_232,N_4924,N_4810);
nor UO_233 (O_233,N_4679,N_4921);
and UO_234 (O_234,N_4701,N_4979);
nor UO_235 (O_235,N_4780,N_4506);
nand UO_236 (O_236,N_4555,N_4566);
and UO_237 (O_237,N_4974,N_4716);
and UO_238 (O_238,N_4519,N_4992);
and UO_239 (O_239,N_4950,N_4871);
and UO_240 (O_240,N_4972,N_4543);
or UO_241 (O_241,N_4949,N_4981);
and UO_242 (O_242,N_4599,N_4820);
nand UO_243 (O_243,N_4817,N_4536);
and UO_244 (O_244,N_4559,N_4696);
or UO_245 (O_245,N_4791,N_4945);
and UO_246 (O_246,N_4692,N_4774);
nor UO_247 (O_247,N_4686,N_4867);
nand UO_248 (O_248,N_4758,N_4569);
and UO_249 (O_249,N_4884,N_4564);
nand UO_250 (O_250,N_4593,N_4701);
or UO_251 (O_251,N_4936,N_4645);
nor UO_252 (O_252,N_4863,N_4781);
and UO_253 (O_253,N_4708,N_4888);
and UO_254 (O_254,N_4712,N_4565);
or UO_255 (O_255,N_4971,N_4612);
nor UO_256 (O_256,N_4997,N_4727);
nand UO_257 (O_257,N_4922,N_4927);
nor UO_258 (O_258,N_4772,N_4965);
or UO_259 (O_259,N_4881,N_4872);
or UO_260 (O_260,N_4565,N_4559);
nor UO_261 (O_261,N_4728,N_4790);
and UO_262 (O_262,N_4843,N_4633);
and UO_263 (O_263,N_4597,N_4824);
nor UO_264 (O_264,N_4974,N_4524);
and UO_265 (O_265,N_4517,N_4931);
or UO_266 (O_266,N_4933,N_4614);
nand UO_267 (O_267,N_4680,N_4660);
nor UO_268 (O_268,N_4659,N_4677);
or UO_269 (O_269,N_4702,N_4792);
and UO_270 (O_270,N_4813,N_4945);
nand UO_271 (O_271,N_4648,N_4594);
and UO_272 (O_272,N_4951,N_4665);
nand UO_273 (O_273,N_4634,N_4741);
nand UO_274 (O_274,N_4963,N_4658);
and UO_275 (O_275,N_4567,N_4700);
or UO_276 (O_276,N_4650,N_4976);
and UO_277 (O_277,N_4623,N_4874);
nand UO_278 (O_278,N_4910,N_4757);
xor UO_279 (O_279,N_4993,N_4560);
nand UO_280 (O_280,N_4794,N_4693);
and UO_281 (O_281,N_4726,N_4841);
or UO_282 (O_282,N_4740,N_4826);
and UO_283 (O_283,N_4731,N_4837);
or UO_284 (O_284,N_4969,N_4760);
nand UO_285 (O_285,N_4597,N_4979);
or UO_286 (O_286,N_4720,N_4894);
nand UO_287 (O_287,N_4681,N_4966);
and UO_288 (O_288,N_4715,N_4638);
and UO_289 (O_289,N_4955,N_4737);
or UO_290 (O_290,N_4649,N_4511);
nand UO_291 (O_291,N_4720,N_4724);
and UO_292 (O_292,N_4526,N_4578);
nor UO_293 (O_293,N_4626,N_4982);
nand UO_294 (O_294,N_4883,N_4727);
or UO_295 (O_295,N_4935,N_4591);
nor UO_296 (O_296,N_4808,N_4840);
and UO_297 (O_297,N_4882,N_4540);
and UO_298 (O_298,N_4777,N_4957);
nand UO_299 (O_299,N_4993,N_4828);
and UO_300 (O_300,N_4593,N_4976);
or UO_301 (O_301,N_4850,N_4862);
or UO_302 (O_302,N_4671,N_4592);
nand UO_303 (O_303,N_4673,N_4909);
nor UO_304 (O_304,N_4999,N_4538);
and UO_305 (O_305,N_4580,N_4802);
nor UO_306 (O_306,N_4632,N_4703);
and UO_307 (O_307,N_4741,N_4816);
and UO_308 (O_308,N_4754,N_4722);
nor UO_309 (O_309,N_4817,N_4878);
or UO_310 (O_310,N_4660,N_4739);
or UO_311 (O_311,N_4844,N_4790);
and UO_312 (O_312,N_4765,N_4551);
nor UO_313 (O_313,N_4895,N_4713);
and UO_314 (O_314,N_4506,N_4785);
or UO_315 (O_315,N_4989,N_4613);
and UO_316 (O_316,N_4981,N_4929);
nand UO_317 (O_317,N_4551,N_4541);
nor UO_318 (O_318,N_4591,N_4555);
and UO_319 (O_319,N_4744,N_4697);
nor UO_320 (O_320,N_4882,N_4866);
nand UO_321 (O_321,N_4900,N_4507);
nand UO_322 (O_322,N_4940,N_4606);
nand UO_323 (O_323,N_4644,N_4999);
and UO_324 (O_324,N_4953,N_4584);
nor UO_325 (O_325,N_4866,N_4920);
and UO_326 (O_326,N_4729,N_4637);
nand UO_327 (O_327,N_4932,N_4974);
and UO_328 (O_328,N_4878,N_4767);
or UO_329 (O_329,N_4948,N_4591);
or UO_330 (O_330,N_4748,N_4520);
nor UO_331 (O_331,N_4873,N_4744);
nand UO_332 (O_332,N_4929,N_4982);
nor UO_333 (O_333,N_4750,N_4815);
nor UO_334 (O_334,N_4689,N_4802);
and UO_335 (O_335,N_4593,N_4731);
nor UO_336 (O_336,N_4523,N_4900);
nor UO_337 (O_337,N_4810,N_4589);
or UO_338 (O_338,N_4633,N_4757);
or UO_339 (O_339,N_4774,N_4807);
nor UO_340 (O_340,N_4547,N_4645);
or UO_341 (O_341,N_4910,N_4847);
or UO_342 (O_342,N_4511,N_4983);
nand UO_343 (O_343,N_4800,N_4770);
and UO_344 (O_344,N_4883,N_4801);
nand UO_345 (O_345,N_4676,N_4704);
nand UO_346 (O_346,N_4650,N_4605);
nand UO_347 (O_347,N_4674,N_4871);
or UO_348 (O_348,N_4593,N_4648);
or UO_349 (O_349,N_4912,N_4522);
or UO_350 (O_350,N_4788,N_4808);
nor UO_351 (O_351,N_4725,N_4690);
nand UO_352 (O_352,N_4508,N_4655);
and UO_353 (O_353,N_4766,N_4541);
or UO_354 (O_354,N_4995,N_4575);
and UO_355 (O_355,N_4964,N_4681);
and UO_356 (O_356,N_4847,N_4959);
nor UO_357 (O_357,N_4704,N_4569);
nor UO_358 (O_358,N_4916,N_4769);
or UO_359 (O_359,N_4521,N_4652);
or UO_360 (O_360,N_4537,N_4605);
nand UO_361 (O_361,N_4696,N_4787);
nor UO_362 (O_362,N_4850,N_4967);
and UO_363 (O_363,N_4877,N_4719);
nand UO_364 (O_364,N_4500,N_4944);
and UO_365 (O_365,N_4912,N_4786);
nand UO_366 (O_366,N_4625,N_4694);
or UO_367 (O_367,N_4513,N_4616);
nor UO_368 (O_368,N_4504,N_4913);
nor UO_369 (O_369,N_4513,N_4966);
and UO_370 (O_370,N_4783,N_4984);
or UO_371 (O_371,N_4662,N_4868);
and UO_372 (O_372,N_4654,N_4562);
nand UO_373 (O_373,N_4510,N_4969);
or UO_374 (O_374,N_4947,N_4960);
and UO_375 (O_375,N_4901,N_4590);
and UO_376 (O_376,N_4800,N_4903);
nand UO_377 (O_377,N_4881,N_4710);
and UO_378 (O_378,N_4517,N_4737);
and UO_379 (O_379,N_4554,N_4873);
or UO_380 (O_380,N_4929,N_4998);
nor UO_381 (O_381,N_4639,N_4941);
nand UO_382 (O_382,N_4905,N_4552);
nor UO_383 (O_383,N_4994,N_4844);
nand UO_384 (O_384,N_4856,N_4987);
nor UO_385 (O_385,N_4715,N_4531);
nor UO_386 (O_386,N_4611,N_4527);
or UO_387 (O_387,N_4843,N_4963);
and UO_388 (O_388,N_4615,N_4916);
or UO_389 (O_389,N_4562,N_4509);
and UO_390 (O_390,N_4787,N_4517);
nand UO_391 (O_391,N_4853,N_4534);
and UO_392 (O_392,N_4661,N_4707);
and UO_393 (O_393,N_4575,N_4577);
nor UO_394 (O_394,N_4556,N_4859);
or UO_395 (O_395,N_4865,N_4563);
xnor UO_396 (O_396,N_4564,N_4987);
or UO_397 (O_397,N_4578,N_4618);
nor UO_398 (O_398,N_4560,N_4548);
nand UO_399 (O_399,N_4987,N_4888);
nand UO_400 (O_400,N_4651,N_4833);
xor UO_401 (O_401,N_4580,N_4534);
nand UO_402 (O_402,N_4619,N_4828);
and UO_403 (O_403,N_4636,N_4752);
or UO_404 (O_404,N_4933,N_4584);
nand UO_405 (O_405,N_4554,N_4995);
and UO_406 (O_406,N_4982,N_4546);
nor UO_407 (O_407,N_4647,N_4542);
nand UO_408 (O_408,N_4945,N_4907);
or UO_409 (O_409,N_4818,N_4863);
or UO_410 (O_410,N_4710,N_4961);
nor UO_411 (O_411,N_4930,N_4716);
and UO_412 (O_412,N_4872,N_4505);
and UO_413 (O_413,N_4733,N_4763);
and UO_414 (O_414,N_4526,N_4597);
nand UO_415 (O_415,N_4608,N_4579);
or UO_416 (O_416,N_4592,N_4947);
nor UO_417 (O_417,N_4994,N_4650);
nand UO_418 (O_418,N_4973,N_4551);
nor UO_419 (O_419,N_4506,N_4609);
or UO_420 (O_420,N_4638,N_4873);
and UO_421 (O_421,N_4899,N_4957);
nor UO_422 (O_422,N_4933,N_4644);
nor UO_423 (O_423,N_4676,N_4697);
or UO_424 (O_424,N_4516,N_4537);
nor UO_425 (O_425,N_4666,N_4939);
or UO_426 (O_426,N_4518,N_4616);
nor UO_427 (O_427,N_4793,N_4571);
nor UO_428 (O_428,N_4544,N_4648);
or UO_429 (O_429,N_4544,N_4689);
nor UO_430 (O_430,N_4635,N_4630);
nand UO_431 (O_431,N_4527,N_4860);
or UO_432 (O_432,N_4691,N_4776);
and UO_433 (O_433,N_4697,N_4856);
nor UO_434 (O_434,N_4886,N_4794);
nand UO_435 (O_435,N_4917,N_4542);
nand UO_436 (O_436,N_4646,N_4528);
nand UO_437 (O_437,N_4869,N_4990);
nor UO_438 (O_438,N_4909,N_4614);
and UO_439 (O_439,N_4981,N_4756);
nand UO_440 (O_440,N_4917,N_4500);
nand UO_441 (O_441,N_4931,N_4782);
or UO_442 (O_442,N_4541,N_4835);
nor UO_443 (O_443,N_4925,N_4533);
or UO_444 (O_444,N_4846,N_4517);
or UO_445 (O_445,N_4859,N_4534);
and UO_446 (O_446,N_4852,N_4964);
or UO_447 (O_447,N_4620,N_4665);
and UO_448 (O_448,N_4735,N_4722);
nand UO_449 (O_449,N_4682,N_4930);
or UO_450 (O_450,N_4804,N_4749);
or UO_451 (O_451,N_4991,N_4719);
nor UO_452 (O_452,N_4556,N_4684);
nand UO_453 (O_453,N_4687,N_4558);
nand UO_454 (O_454,N_4799,N_4651);
nor UO_455 (O_455,N_4566,N_4560);
or UO_456 (O_456,N_4708,N_4910);
and UO_457 (O_457,N_4712,N_4877);
or UO_458 (O_458,N_4782,N_4589);
nor UO_459 (O_459,N_4561,N_4863);
nand UO_460 (O_460,N_4958,N_4749);
nand UO_461 (O_461,N_4838,N_4962);
nor UO_462 (O_462,N_4826,N_4835);
xor UO_463 (O_463,N_4984,N_4585);
nor UO_464 (O_464,N_4794,N_4695);
nand UO_465 (O_465,N_4752,N_4854);
nand UO_466 (O_466,N_4659,N_4807);
or UO_467 (O_467,N_4901,N_4672);
nand UO_468 (O_468,N_4859,N_4664);
or UO_469 (O_469,N_4700,N_4989);
and UO_470 (O_470,N_4886,N_4593);
nand UO_471 (O_471,N_4770,N_4996);
nor UO_472 (O_472,N_4544,N_4826);
or UO_473 (O_473,N_4941,N_4537);
nor UO_474 (O_474,N_4556,N_4678);
nand UO_475 (O_475,N_4985,N_4989);
nor UO_476 (O_476,N_4934,N_4720);
nor UO_477 (O_477,N_4635,N_4899);
nor UO_478 (O_478,N_4634,N_4754);
nand UO_479 (O_479,N_4960,N_4884);
and UO_480 (O_480,N_4972,N_4915);
and UO_481 (O_481,N_4544,N_4538);
nand UO_482 (O_482,N_4996,N_4803);
nand UO_483 (O_483,N_4526,N_4552);
nor UO_484 (O_484,N_4730,N_4926);
and UO_485 (O_485,N_4873,N_4952);
or UO_486 (O_486,N_4728,N_4609);
nand UO_487 (O_487,N_4776,N_4987);
nor UO_488 (O_488,N_4640,N_4547);
and UO_489 (O_489,N_4529,N_4548);
or UO_490 (O_490,N_4957,N_4868);
nor UO_491 (O_491,N_4947,N_4525);
xnor UO_492 (O_492,N_4654,N_4688);
nor UO_493 (O_493,N_4911,N_4716);
nor UO_494 (O_494,N_4748,N_4829);
nand UO_495 (O_495,N_4855,N_4614);
nor UO_496 (O_496,N_4597,N_4787);
and UO_497 (O_497,N_4988,N_4926);
or UO_498 (O_498,N_4952,N_4991);
nor UO_499 (O_499,N_4584,N_4658);
nand UO_500 (O_500,N_4814,N_4586);
nand UO_501 (O_501,N_4762,N_4580);
or UO_502 (O_502,N_4806,N_4912);
or UO_503 (O_503,N_4582,N_4769);
nor UO_504 (O_504,N_4914,N_4885);
nor UO_505 (O_505,N_4846,N_4979);
nor UO_506 (O_506,N_4925,N_4604);
and UO_507 (O_507,N_4589,N_4623);
nor UO_508 (O_508,N_4989,N_4703);
or UO_509 (O_509,N_4890,N_4813);
and UO_510 (O_510,N_4584,N_4972);
and UO_511 (O_511,N_4923,N_4619);
nor UO_512 (O_512,N_4939,N_4759);
nor UO_513 (O_513,N_4614,N_4568);
nor UO_514 (O_514,N_4547,N_4578);
and UO_515 (O_515,N_4889,N_4989);
nor UO_516 (O_516,N_4885,N_4629);
and UO_517 (O_517,N_4892,N_4517);
nand UO_518 (O_518,N_4650,N_4525);
and UO_519 (O_519,N_4929,N_4927);
nor UO_520 (O_520,N_4880,N_4771);
nand UO_521 (O_521,N_4819,N_4664);
nor UO_522 (O_522,N_4857,N_4618);
nand UO_523 (O_523,N_4840,N_4978);
and UO_524 (O_524,N_4545,N_4897);
and UO_525 (O_525,N_4784,N_4968);
nand UO_526 (O_526,N_4908,N_4821);
nor UO_527 (O_527,N_4646,N_4996);
nand UO_528 (O_528,N_4509,N_4545);
nor UO_529 (O_529,N_4632,N_4651);
nor UO_530 (O_530,N_4798,N_4541);
nor UO_531 (O_531,N_4884,N_4834);
and UO_532 (O_532,N_4669,N_4523);
nand UO_533 (O_533,N_4705,N_4920);
nand UO_534 (O_534,N_4612,N_4559);
and UO_535 (O_535,N_4946,N_4850);
or UO_536 (O_536,N_4970,N_4909);
and UO_537 (O_537,N_4949,N_4778);
nand UO_538 (O_538,N_4525,N_4591);
nand UO_539 (O_539,N_4803,N_4650);
or UO_540 (O_540,N_4598,N_4678);
nor UO_541 (O_541,N_4796,N_4686);
or UO_542 (O_542,N_4613,N_4944);
or UO_543 (O_543,N_4659,N_4961);
nor UO_544 (O_544,N_4921,N_4647);
nor UO_545 (O_545,N_4862,N_4618);
or UO_546 (O_546,N_4948,N_4553);
nor UO_547 (O_547,N_4717,N_4850);
nand UO_548 (O_548,N_4575,N_4593);
and UO_549 (O_549,N_4870,N_4887);
or UO_550 (O_550,N_4896,N_4858);
nand UO_551 (O_551,N_4531,N_4664);
and UO_552 (O_552,N_4638,N_4903);
nor UO_553 (O_553,N_4681,N_4934);
and UO_554 (O_554,N_4590,N_4636);
and UO_555 (O_555,N_4771,N_4948);
and UO_556 (O_556,N_4551,N_4604);
or UO_557 (O_557,N_4542,N_4896);
or UO_558 (O_558,N_4845,N_4927);
nand UO_559 (O_559,N_4513,N_4712);
nor UO_560 (O_560,N_4981,N_4689);
nor UO_561 (O_561,N_4661,N_4566);
or UO_562 (O_562,N_4568,N_4965);
and UO_563 (O_563,N_4967,N_4877);
and UO_564 (O_564,N_4786,N_4526);
nor UO_565 (O_565,N_4670,N_4817);
or UO_566 (O_566,N_4583,N_4951);
nand UO_567 (O_567,N_4663,N_4522);
nor UO_568 (O_568,N_4594,N_4896);
nand UO_569 (O_569,N_4697,N_4737);
and UO_570 (O_570,N_4582,N_4890);
nand UO_571 (O_571,N_4940,N_4650);
nand UO_572 (O_572,N_4864,N_4513);
or UO_573 (O_573,N_4715,N_4825);
nor UO_574 (O_574,N_4769,N_4721);
nand UO_575 (O_575,N_4761,N_4549);
nor UO_576 (O_576,N_4913,N_4917);
and UO_577 (O_577,N_4589,N_4800);
nor UO_578 (O_578,N_4909,N_4874);
nand UO_579 (O_579,N_4752,N_4715);
and UO_580 (O_580,N_4548,N_4879);
nand UO_581 (O_581,N_4756,N_4609);
and UO_582 (O_582,N_4832,N_4674);
nor UO_583 (O_583,N_4796,N_4778);
and UO_584 (O_584,N_4902,N_4645);
and UO_585 (O_585,N_4686,N_4585);
or UO_586 (O_586,N_4991,N_4683);
nor UO_587 (O_587,N_4991,N_4799);
nand UO_588 (O_588,N_4766,N_4832);
nor UO_589 (O_589,N_4802,N_4813);
or UO_590 (O_590,N_4808,N_4878);
nor UO_591 (O_591,N_4920,N_4567);
nand UO_592 (O_592,N_4697,N_4707);
nor UO_593 (O_593,N_4617,N_4756);
or UO_594 (O_594,N_4669,N_4881);
nor UO_595 (O_595,N_4876,N_4679);
or UO_596 (O_596,N_4585,N_4550);
and UO_597 (O_597,N_4711,N_4906);
and UO_598 (O_598,N_4829,N_4819);
or UO_599 (O_599,N_4534,N_4753);
or UO_600 (O_600,N_4881,N_4531);
nand UO_601 (O_601,N_4955,N_4893);
and UO_602 (O_602,N_4561,N_4947);
or UO_603 (O_603,N_4691,N_4966);
or UO_604 (O_604,N_4821,N_4542);
and UO_605 (O_605,N_4640,N_4829);
nor UO_606 (O_606,N_4651,N_4737);
nand UO_607 (O_607,N_4536,N_4955);
or UO_608 (O_608,N_4781,N_4679);
nor UO_609 (O_609,N_4856,N_4668);
nor UO_610 (O_610,N_4909,N_4526);
or UO_611 (O_611,N_4844,N_4627);
nor UO_612 (O_612,N_4969,N_4620);
nor UO_613 (O_613,N_4590,N_4793);
xor UO_614 (O_614,N_4661,N_4676);
and UO_615 (O_615,N_4977,N_4981);
or UO_616 (O_616,N_4854,N_4669);
nor UO_617 (O_617,N_4735,N_4949);
nand UO_618 (O_618,N_4975,N_4702);
and UO_619 (O_619,N_4825,N_4796);
nand UO_620 (O_620,N_4801,N_4725);
nand UO_621 (O_621,N_4626,N_4802);
and UO_622 (O_622,N_4529,N_4883);
or UO_623 (O_623,N_4604,N_4653);
and UO_624 (O_624,N_4551,N_4593);
nand UO_625 (O_625,N_4947,N_4695);
nand UO_626 (O_626,N_4539,N_4578);
or UO_627 (O_627,N_4751,N_4828);
or UO_628 (O_628,N_4801,N_4698);
xnor UO_629 (O_629,N_4625,N_4681);
nor UO_630 (O_630,N_4695,N_4767);
or UO_631 (O_631,N_4621,N_4629);
or UO_632 (O_632,N_4715,N_4559);
nor UO_633 (O_633,N_4719,N_4995);
and UO_634 (O_634,N_4684,N_4809);
and UO_635 (O_635,N_4763,N_4648);
and UO_636 (O_636,N_4754,N_4692);
or UO_637 (O_637,N_4737,N_4740);
or UO_638 (O_638,N_4745,N_4823);
and UO_639 (O_639,N_4939,N_4603);
nor UO_640 (O_640,N_4617,N_4508);
or UO_641 (O_641,N_4616,N_4760);
or UO_642 (O_642,N_4511,N_4686);
or UO_643 (O_643,N_4651,N_4826);
nand UO_644 (O_644,N_4903,N_4996);
and UO_645 (O_645,N_4738,N_4810);
or UO_646 (O_646,N_4894,N_4711);
nor UO_647 (O_647,N_4770,N_4557);
nor UO_648 (O_648,N_4679,N_4890);
and UO_649 (O_649,N_4703,N_4866);
and UO_650 (O_650,N_4785,N_4587);
nor UO_651 (O_651,N_4727,N_4825);
and UO_652 (O_652,N_4593,N_4541);
nand UO_653 (O_653,N_4862,N_4927);
nor UO_654 (O_654,N_4953,N_4589);
nand UO_655 (O_655,N_4964,N_4634);
and UO_656 (O_656,N_4684,N_4638);
or UO_657 (O_657,N_4819,N_4828);
and UO_658 (O_658,N_4827,N_4685);
nor UO_659 (O_659,N_4787,N_4634);
nor UO_660 (O_660,N_4936,N_4744);
and UO_661 (O_661,N_4998,N_4789);
and UO_662 (O_662,N_4960,N_4571);
nand UO_663 (O_663,N_4738,N_4824);
or UO_664 (O_664,N_4511,N_4503);
nand UO_665 (O_665,N_4516,N_4933);
nor UO_666 (O_666,N_4529,N_4998);
nor UO_667 (O_667,N_4831,N_4841);
or UO_668 (O_668,N_4650,N_4670);
nand UO_669 (O_669,N_4574,N_4820);
or UO_670 (O_670,N_4709,N_4794);
and UO_671 (O_671,N_4746,N_4663);
and UO_672 (O_672,N_4846,N_4666);
and UO_673 (O_673,N_4976,N_4575);
or UO_674 (O_674,N_4509,N_4879);
nor UO_675 (O_675,N_4507,N_4684);
and UO_676 (O_676,N_4764,N_4886);
or UO_677 (O_677,N_4828,N_4989);
nand UO_678 (O_678,N_4788,N_4534);
and UO_679 (O_679,N_4615,N_4737);
nor UO_680 (O_680,N_4935,N_4597);
nand UO_681 (O_681,N_4843,N_4901);
or UO_682 (O_682,N_4805,N_4740);
or UO_683 (O_683,N_4654,N_4640);
and UO_684 (O_684,N_4596,N_4981);
nand UO_685 (O_685,N_4824,N_4857);
or UO_686 (O_686,N_4652,N_4794);
nand UO_687 (O_687,N_4658,N_4677);
or UO_688 (O_688,N_4812,N_4744);
xnor UO_689 (O_689,N_4601,N_4878);
or UO_690 (O_690,N_4580,N_4845);
and UO_691 (O_691,N_4831,N_4791);
or UO_692 (O_692,N_4811,N_4674);
or UO_693 (O_693,N_4573,N_4610);
or UO_694 (O_694,N_4531,N_4878);
or UO_695 (O_695,N_4594,N_4519);
nor UO_696 (O_696,N_4979,N_4753);
nand UO_697 (O_697,N_4610,N_4626);
and UO_698 (O_698,N_4565,N_4800);
or UO_699 (O_699,N_4589,N_4771);
and UO_700 (O_700,N_4941,N_4507);
nand UO_701 (O_701,N_4731,N_4641);
nor UO_702 (O_702,N_4611,N_4687);
nor UO_703 (O_703,N_4928,N_4880);
nand UO_704 (O_704,N_4934,N_4586);
nor UO_705 (O_705,N_4928,N_4604);
nor UO_706 (O_706,N_4598,N_4922);
and UO_707 (O_707,N_4608,N_4658);
nand UO_708 (O_708,N_4581,N_4628);
or UO_709 (O_709,N_4590,N_4568);
nand UO_710 (O_710,N_4504,N_4752);
nor UO_711 (O_711,N_4747,N_4536);
nor UO_712 (O_712,N_4642,N_4698);
or UO_713 (O_713,N_4933,N_4622);
and UO_714 (O_714,N_4935,N_4663);
or UO_715 (O_715,N_4585,N_4932);
nand UO_716 (O_716,N_4636,N_4851);
and UO_717 (O_717,N_4676,N_4693);
and UO_718 (O_718,N_4789,N_4741);
or UO_719 (O_719,N_4890,N_4753);
and UO_720 (O_720,N_4595,N_4598);
and UO_721 (O_721,N_4523,N_4618);
nor UO_722 (O_722,N_4878,N_4589);
nand UO_723 (O_723,N_4504,N_4893);
and UO_724 (O_724,N_4817,N_4698);
and UO_725 (O_725,N_4880,N_4702);
or UO_726 (O_726,N_4840,N_4565);
nor UO_727 (O_727,N_4721,N_4948);
nand UO_728 (O_728,N_4723,N_4815);
or UO_729 (O_729,N_4954,N_4827);
and UO_730 (O_730,N_4597,N_4649);
and UO_731 (O_731,N_4751,N_4680);
and UO_732 (O_732,N_4506,N_4755);
nand UO_733 (O_733,N_4870,N_4916);
nor UO_734 (O_734,N_4887,N_4687);
nand UO_735 (O_735,N_4699,N_4979);
or UO_736 (O_736,N_4685,N_4561);
and UO_737 (O_737,N_4796,N_4974);
or UO_738 (O_738,N_4525,N_4934);
and UO_739 (O_739,N_4988,N_4952);
nand UO_740 (O_740,N_4551,N_4811);
and UO_741 (O_741,N_4629,N_4778);
and UO_742 (O_742,N_4873,N_4800);
or UO_743 (O_743,N_4586,N_4767);
or UO_744 (O_744,N_4557,N_4608);
and UO_745 (O_745,N_4612,N_4503);
nand UO_746 (O_746,N_4978,N_4944);
nor UO_747 (O_747,N_4732,N_4626);
nor UO_748 (O_748,N_4755,N_4530);
nand UO_749 (O_749,N_4962,N_4905);
nand UO_750 (O_750,N_4538,N_4568);
and UO_751 (O_751,N_4539,N_4951);
nand UO_752 (O_752,N_4954,N_4566);
or UO_753 (O_753,N_4534,N_4777);
and UO_754 (O_754,N_4809,N_4907);
or UO_755 (O_755,N_4942,N_4535);
nand UO_756 (O_756,N_4822,N_4990);
nor UO_757 (O_757,N_4587,N_4655);
nor UO_758 (O_758,N_4796,N_4672);
nor UO_759 (O_759,N_4855,N_4547);
nand UO_760 (O_760,N_4852,N_4763);
nor UO_761 (O_761,N_4599,N_4769);
nand UO_762 (O_762,N_4500,N_4834);
and UO_763 (O_763,N_4793,N_4833);
or UO_764 (O_764,N_4794,N_4848);
nand UO_765 (O_765,N_4708,N_4611);
and UO_766 (O_766,N_4996,N_4610);
or UO_767 (O_767,N_4994,N_4864);
and UO_768 (O_768,N_4532,N_4586);
or UO_769 (O_769,N_4912,N_4524);
or UO_770 (O_770,N_4581,N_4580);
nand UO_771 (O_771,N_4873,N_4696);
nand UO_772 (O_772,N_4906,N_4689);
nor UO_773 (O_773,N_4700,N_4915);
nor UO_774 (O_774,N_4551,N_4978);
nand UO_775 (O_775,N_4685,N_4523);
or UO_776 (O_776,N_4668,N_4787);
nor UO_777 (O_777,N_4618,N_4682);
nand UO_778 (O_778,N_4926,N_4676);
or UO_779 (O_779,N_4714,N_4589);
and UO_780 (O_780,N_4667,N_4501);
and UO_781 (O_781,N_4553,N_4669);
nand UO_782 (O_782,N_4898,N_4854);
nor UO_783 (O_783,N_4921,N_4574);
and UO_784 (O_784,N_4863,N_4711);
and UO_785 (O_785,N_4500,N_4946);
or UO_786 (O_786,N_4713,N_4607);
or UO_787 (O_787,N_4525,N_4589);
or UO_788 (O_788,N_4559,N_4546);
nand UO_789 (O_789,N_4712,N_4700);
and UO_790 (O_790,N_4904,N_4676);
nor UO_791 (O_791,N_4980,N_4793);
and UO_792 (O_792,N_4678,N_4515);
and UO_793 (O_793,N_4701,N_4688);
or UO_794 (O_794,N_4802,N_4974);
nor UO_795 (O_795,N_4706,N_4694);
nor UO_796 (O_796,N_4838,N_4683);
nor UO_797 (O_797,N_4833,N_4692);
nor UO_798 (O_798,N_4768,N_4668);
nand UO_799 (O_799,N_4986,N_4873);
nand UO_800 (O_800,N_4780,N_4725);
nand UO_801 (O_801,N_4703,N_4882);
nand UO_802 (O_802,N_4555,N_4874);
nor UO_803 (O_803,N_4755,N_4847);
nor UO_804 (O_804,N_4824,N_4825);
nor UO_805 (O_805,N_4527,N_4957);
and UO_806 (O_806,N_4602,N_4800);
nand UO_807 (O_807,N_4849,N_4519);
or UO_808 (O_808,N_4576,N_4879);
nand UO_809 (O_809,N_4841,N_4798);
nand UO_810 (O_810,N_4896,N_4983);
nor UO_811 (O_811,N_4540,N_4548);
or UO_812 (O_812,N_4539,N_4749);
and UO_813 (O_813,N_4741,N_4697);
nor UO_814 (O_814,N_4501,N_4730);
or UO_815 (O_815,N_4545,N_4555);
and UO_816 (O_816,N_4875,N_4674);
nor UO_817 (O_817,N_4755,N_4891);
nor UO_818 (O_818,N_4825,N_4863);
or UO_819 (O_819,N_4804,N_4587);
or UO_820 (O_820,N_4649,N_4512);
nand UO_821 (O_821,N_4848,N_4765);
and UO_822 (O_822,N_4806,N_4909);
nand UO_823 (O_823,N_4760,N_4774);
nand UO_824 (O_824,N_4793,N_4821);
nand UO_825 (O_825,N_4849,N_4986);
nor UO_826 (O_826,N_4632,N_4922);
nor UO_827 (O_827,N_4554,N_4762);
nor UO_828 (O_828,N_4736,N_4724);
nor UO_829 (O_829,N_4895,N_4513);
nand UO_830 (O_830,N_4796,N_4532);
nand UO_831 (O_831,N_4831,N_4928);
or UO_832 (O_832,N_4739,N_4851);
and UO_833 (O_833,N_4988,N_4841);
nand UO_834 (O_834,N_4814,N_4822);
and UO_835 (O_835,N_4574,N_4639);
nand UO_836 (O_836,N_4859,N_4985);
and UO_837 (O_837,N_4892,N_4872);
and UO_838 (O_838,N_4881,N_4757);
and UO_839 (O_839,N_4913,N_4738);
nor UO_840 (O_840,N_4621,N_4695);
nand UO_841 (O_841,N_4965,N_4932);
nor UO_842 (O_842,N_4802,N_4864);
and UO_843 (O_843,N_4662,N_4909);
or UO_844 (O_844,N_4589,N_4836);
nor UO_845 (O_845,N_4520,N_4502);
nor UO_846 (O_846,N_4645,N_4877);
or UO_847 (O_847,N_4718,N_4985);
nand UO_848 (O_848,N_4600,N_4915);
nor UO_849 (O_849,N_4703,N_4699);
xor UO_850 (O_850,N_4809,N_4556);
or UO_851 (O_851,N_4534,N_4894);
nor UO_852 (O_852,N_4831,N_4798);
and UO_853 (O_853,N_4519,N_4667);
nand UO_854 (O_854,N_4902,N_4719);
nand UO_855 (O_855,N_4570,N_4555);
or UO_856 (O_856,N_4963,N_4623);
or UO_857 (O_857,N_4958,N_4833);
nand UO_858 (O_858,N_4714,N_4994);
nor UO_859 (O_859,N_4500,N_4758);
and UO_860 (O_860,N_4716,N_4532);
and UO_861 (O_861,N_4650,N_4841);
nor UO_862 (O_862,N_4683,N_4684);
and UO_863 (O_863,N_4591,N_4840);
or UO_864 (O_864,N_4995,N_4685);
or UO_865 (O_865,N_4513,N_4901);
nor UO_866 (O_866,N_4649,N_4678);
or UO_867 (O_867,N_4817,N_4755);
nand UO_868 (O_868,N_4563,N_4560);
nor UO_869 (O_869,N_4958,N_4948);
and UO_870 (O_870,N_4830,N_4870);
and UO_871 (O_871,N_4841,N_4870);
nand UO_872 (O_872,N_4668,N_4750);
nand UO_873 (O_873,N_4649,N_4742);
or UO_874 (O_874,N_4951,N_4679);
nor UO_875 (O_875,N_4979,N_4876);
and UO_876 (O_876,N_4844,N_4787);
nor UO_877 (O_877,N_4668,N_4736);
or UO_878 (O_878,N_4960,N_4558);
nor UO_879 (O_879,N_4884,N_4629);
nor UO_880 (O_880,N_4594,N_4966);
or UO_881 (O_881,N_4762,N_4908);
and UO_882 (O_882,N_4639,N_4657);
nand UO_883 (O_883,N_4692,N_4952);
nand UO_884 (O_884,N_4677,N_4565);
nor UO_885 (O_885,N_4915,N_4729);
and UO_886 (O_886,N_4998,N_4597);
nor UO_887 (O_887,N_4947,N_4844);
or UO_888 (O_888,N_4805,N_4721);
nand UO_889 (O_889,N_4731,N_4989);
or UO_890 (O_890,N_4731,N_4640);
or UO_891 (O_891,N_4790,N_4675);
nor UO_892 (O_892,N_4888,N_4729);
and UO_893 (O_893,N_4502,N_4660);
or UO_894 (O_894,N_4622,N_4919);
nand UO_895 (O_895,N_4682,N_4625);
xnor UO_896 (O_896,N_4835,N_4881);
nand UO_897 (O_897,N_4827,N_4556);
and UO_898 (O_898,N_4768,N_4914);
nand UO_899 (O_899,N_4932,N_4569);
nor UO_900 (O_900,N_4990,N_4918);
nor UO_901 (O_901,N_4936,N_4627);
and UO_902 (O_902,N_4857,N_4558);
or UO_903 (O_903,N_4881,N_4567);
nor UO_904 (O_904,N_4800,N_4967);
or UO_905 (O_905,N_4954,N_4662);
nand UO_906 (O_906,N_4919,N_4977);
nand UO_907 (O_907,N_4774,N_4824);
nand UO_908 (O_908,N_4673,N_4751);
and UO_909 (O_909,N_4907,N_4663);
nor UO_910 (O_910,N_4780,N_4750);
and UO_911 (O_911,N_4506,N_4772);
nand UO_912 (O_912,N_4646,N_4632);
or UO_913 (O_913,N_4734,N_4759);
nand UO_914 (O_914,N_4999,N_4687);
nand UO_915 (O_915,N_4582,N_4716);
and UO_916 (O_916,N_4897,N_4669);
nor UO_917 (O_917,N_4748,N_4603);
nor UO_918 (O_918,N_4675,N_4717);
or UO_919 (O_919,N_4919,N_4511);
and UO_920 (O_920,N_4792,N_4630);
and UO_921 (O_921,N_4979,N_4789);
nor UO_922 (O_922,N_4839,N_4797);
and UO_923 (O_923,N_4767,N_4707);
and UO_924 (O_924,N_4953,N_4979);
or UO_925 (O_925,N_4640,N_4721);
and UO_926 (O_926,N_4858,N_4818);
or UO_927 (O_927,N_4685,N_4792);
and UO_928 (O_928,N_4652,N_4854);
or UO_929 (O_929,N_4596,N_4957);
and UO_930 (O_930,N_4520,N_4785);
nand UO_931 (O_931,N_4543,N_4644);
nor UO_932 (O_932,N_4880,N_4918);
nand UO_933 (O_933,N_4974,N_4865);
nand UO_934 (O_934,N_4785,N_4600);
or UO_935 (O_935,N_4844,N_4818);
and UO_936 (O_936,N_4991,N_4912);
nor UO_937 (O_937,N_4708,N_4920);
nor UO_938 (O_938,N_4717,N_4729);
and UO_939 (O_939,N_4992,N_4931);
nor UO_940 (O_940,N_4811,N_4990);
and UO_941 (O_941,N_4517,N_4652);
nor UO_942 (O_942,N_4926,N_4815);
nand UO_943 (O_943,N_4854,N_4927);
or UO_944 (O_944,N_4503,N_4790);
nand UO_945 (O_945,N_4788,N_4596);
or UO_946 (O_946,N_4544,N_4608);
and UO_947 (O_947,N_4712,N_4922);
or UO_948 (O_948,N_4581,N_4815);
or UO_949 (O_949,N_4866,N_4719);
nor UO_950 (O_950,N_4723,N_4891);
nand UO_951 (O_951,N_4936,N_4884);
and UO_952 (O_952,N_4796,N_4907);
and UO_953 (O_953,N_4866,N_4540);
nor UO_954 (O_954,N_4740,N_4611);
or UO_955 (O_955,N_4955,N_4630);
nand UO_956 (O_956,N_4714,N_4896);
nand UO_957 (O_957,N_4758,N_4517);
or UO_958 (O_958,N_4981,N_4681);
nor UO_959 (O_959,N_4734,N_4708);
and UO_960 (O_960,N_4598,N_4772);
or UO_961 (O_961,N_4703,N_4545);
nand UO_962 (O_962,N_4885,N_4582);
nor UO_963 (O_963,N_4787,N_4951);
nor UO_964 (O_964,N_4616,N_4943);
nand UO_965 (O_965,N_4541,N_4651);
and UO_966 (O_966,N_4650,N_4955);
nand UO_967 (O_967,N_4889,N_4665);
or UO_968 (O_968,N_4743,N_4545);
nor UO_969 (O_969,N_4568,N_4813);
or UO_970 (O_970,N_4635,N_4729);
and UO_971 (O_971,N_4682,N_4884);
nand UO_972 (O_972,N_4729,N_4995);
and UO_973 (O_973,N_4577,N_4726);
or UO_974 (O_974,N_4609,N_4742);
and UO_975 (O_975,N_4534,N_4825);
or UO_976 (O_976,N_4686,N_4773);
nand UO_977 (O_977,N_4640,N_4927);
nand UO_978 (O_978,N_4800,N_4843);
nor UO_979 (O_979,N_4756,N_4857);
nand UO_980 (O_980,N_4885,N_4880);
and UO_981 (O_981,N_4935,N_4667);
and UO_982 (O_982,N_4599,N_4952);
and UO_983 (O_983,N_4855,N_4662);
or UO_984 (O_984,N_4833,N_4844);
nor UO_985 (O_985,N_4836,N_4692);
or UO_986 (O_986,N_4910,N_4848);
nand UO_987 (O_987,N_4919,N_4860);
nor UO_988 (O_988,N_4629,N_4789);
and UO_989 (O_989,N_4712,N_4617);
or UO_990 (O_990,N_4510,N_4624);
and UO_991 (O_991,N_4698,N_4978);
nand UO_992 (O_992,N_4618,N_4956);
and UO_993 (O_993,N_4651,N_4877);
and UO_994 (O_994,N_4646,N_4958);
and UO_995 (O_995,N_4831,N_4712);
and UO_996 (O_996,N_4918,N_4638);
nand UO_997 (O_997,N_4894,N_4758);
or UO_998 (O_998,N_4802,N_4708);
and UO_999 (O_999,N_4691,N_4810);
endmodule