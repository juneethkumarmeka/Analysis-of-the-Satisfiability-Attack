module basic_1000_10000_1500_5_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_833,In_756);
nor U1 (N_1,In_186,In_114);
nand U2 (N_2,In_256,In_282);
nor U3 (N_3,In_215,In_330);
and U4 (N_4,In_537,In_854);
and U5 (N_5,In_948,In_489);
nand U6 (N_6,In_83,In_661);
nor U7 (N_7,In_898,In_936);
nor U8 (N_8,In_824,In_320);
nand U9 (N_9,In_927,In_737);
nor U10 (N_10,In_87,In_490);
and U11 (N_11,In_356,In_352);
nand U12 (N_12,In_705,In_398);
and U13 (N_13,In_216,In_411);
xnor U14 (N_14,In_617,In_906);
and U15 (N_15,In_899,In_228);
or U16 (N_16,In_928,In_664);
or U17 (N_17,In_91,In_478);
and U18 (N_18,In_77,In_673);
or U19 (N_19,In_305,In_378);
nand U20 (N_20,In_389,In_280);
or U21 (N_21,In_197,In_979);
and U22 (N_22,In_657,In_415);
or U23 (N_23,In_968,In_417);
nor U24 (N_24,In_296,In_358);
or U25 (N_25,In_588,In_327);
xor U26 (N_26,In_602,In_525);
or U27 (N_27,In_867,In_696);
or U28 (N_28,In_33,In_106);
and U29 (N_29,In_628,In_800);
nand U30 (N_30,In_89,In_204);
nand U31 (N_31,In_691,In_420);
and U32 (N_32,In_193,In_307);
nor U33 (N_33,In_722,In_931);
nor U34 (N_34,In_865,In_316);
or U35 (N_35,In_333,In_68);
or U36 (N_36,In_183,In_759);
or U37 (N_37,In_714,In_128);
or U38 (N_38,In_450,In_483);
or U39 (N_39,In_96,In_26);
nor U40 (N_40,In_784,In_101);
and U41 (N_41,In_584,In_182);
nand U42 (N_42,In_880,In_404);
or U43 (N_43,In_773,In_125);
nor U44 (N_44,In_903,In_965);
and U45 (N_45,In_325,In_137);
nand U46 (N_46,In_403,In_142);
and U47 (N_47,In_765,In_422);
or U48 (N_48,In_630,In_921);
nor U49 (N_49,In_988,In_161);
and U50 (N_50,In_690,In_318);
nor U51 (N_51,In_19,In_958);
or U52 (N_52,In_946,In_158);
and U53 (N_53,In_603,In_729);
nor U54 (N_54,In_541,In_886);
nand U55 (N_55,In_48,In_770);
nand U56 (N_56,In_817,In_247);
nor U57 (N_57,In_973,In_526);
nor U58 (N_58,In_544,In_185);
nand U59 (N_59,In_970,In_976);
and U60 (N_60,In_834,In_530);
and U61 (N_61,In_589,In_510);
nand U62 (N_62,In_803,In_639);
nand U63 (N_63,In_313,In_146);
and U64 (N_64,In_223,In_295);
nand U65 (N_65,In_39,In_112);
nor U66 (N_66,In_306,In_935);
and U67 (N_67,In_311,In_576);
nor U68 (N_68,In_437,In_986);
nand U69 (N_69,In_761,In_943);
nand U70 (N_70,In_816,In_789);
or U71 (N_71,In_888,In_315);
nand U72 (N_72,In_346,In_753);
or U73 (N_73,In_799,In_907);
or U74 (N_74,In_259,In_942);
or U75 (N_75,In_231,In_500);
or U76 (N_76,In_262,In_874);
nand U77 (N_77,In_517,In_629);
and U78 (N_78,In_268,In_312);
or U79 (N_79,In_50,In_615);
nand U80 (N_80,In_975,In_364);
and U81 (N_81,In_459,In_441);
nand U82 (N_82,In_416,In_273);
nand U83 (N_83,In_766,In_395);
and U84 (N_84,In_872,In_613);
nand U85 (N_85,In_558,In_180);
nor U86 (N_86,In_631,In_245);
and U87 (N_87,In_751,In_987);
nand U88 (N_88,In_43,In_377);
nor U89 (N_89,In_202,In_226);
nor U90 (N_90,In_876,In_674);
or U91 (N_91,In_815,In_263);
or U92 (N_92,In_900,In_16);
and U93 (N_93,In_607,In_80);
or U94 (N_94,In_995,In_980);
nand U95 (N_95,In_782,In_902);
nand U96 (N_96,In_848,In_650);
nor U97 (N_97,In_741,In_731);
nor U98 (N_98,In_894,In_847);
nand U99 (N_99,In_805,In_791);
or U100 (N_100,In_331,In_619);
and U101 (N_101,In_69,In_439);
nand U102 (N_102,In_725,In_301);
nand U103 (N_103,In_961,In_353);
nand U104 (N_104,In_107,In_922);
or U105 (N_105,In_538,In_998);
nand U106 (N_106,In_695,In_655);
nand U107 (N_107,In_21,In_956);
or U108 (N_108,In_598,In_487);
nor U109 (N_109,In_924,In_337);
nor U110 (N_110,In_912,In_365);
nand U111 (N_111,In_555,In_762);
or U112 (N_112,In_14,In_804);
nor U113 (N_113,In_964,In_777);
and U114 (N_114,In_812,In_250);
or U115 (N_115,In_357,In_432);
nor U116 (N_116,In_65,In_474);
or U117 (N_117,In_78,In_425);
nand U118 (N_118,In_570,In_4);
or U119 (N_119,In_326,In_658);
and U120 (N_120,In_994,In_966);
nor U121 (N_121,In_72,In_191);
or U122 (N_122,In_119,In_93);
and U123 (N_123,In_620,In_997);
or U124 (N_124,In_739,In_689);
nor U125 (N_125,In_15,In_520);
nand U126 (N_126,In_669,In_608);
nand U127 (N_127,In_891,In_138);
nand U128 (N_128,In_755,In_497);
and U129 (N_129,In_572,In_379);
and U130 (N_130,In_345,In_332);
or U131 (N_131,In_122,In_594);
nor U132 (N_132,In_347,In_230);
or U133 (N_133,In_435,In_444);
nand U134 (N_134,In_179,In_261);
nor U135 (N_135,In_633,In_218);
nand U136 (N_136,In_303,In_289);
nor U137 (N_137,In_343,In_818);
nand U138 (N_138,In_982,In_473);
or U139 (N_139,In_536,In_727);
nand U140 (N_140,In_823,In_436);
nor U141 (N_141,In_13,In_496);
nor U142 (N_142,In_451,In_243);
nor U143 (N_143,In_317,In_322);
or U144 (N_144,In_11,In_719);
nor U145 (N_145,In_88,In_533);
nor U146 (N_146,In_144,In_49);
nand U147 (N_147,In_813,In_6);
nand U148 (N_148,In_232,In_479);
xnor U149 (N_149,In_857,In_290);
and U150 (N_150,In_267,In_351);
and U151 (N_151,In_644,In_989);
or U152 (N_152,In_29,In_760);
or U153 (N_153,In_844,In_199);
and U154 (N_154,In_985,In_192);
and U155 (N_155,In_699,In_920);
and U156 (N_156,In_772,In_505);
nor U157 (N_157,In_492,In_671);
and U158 (N_158,In_810,In_217);
nor U159 (N_159,In_150,In_362);
or U160 (N_160,In_999,In_391);
and U161 (N_161,In_700,In_592);
or U162 (N_162,In_667,In_646);
nor U163 (N_163,In_776,In_410);
nor U164 (N_164,In_92,In_786);
nor U165 (N_165,In_819,In_569);
nor U166 (N_166,In_654,In_368);
nor U167 (N_167,In_484,In_885);
nand U168 (N_168,In_960,In_471);
nand U169 (N_169,In_547,In_110);
and U170 (N_170,In_668,In_950);
nand U171 (N_171,In_535,In_22);
and U172 (N_172,In_895,In_40);
or U173 (N_173,In_10,In_213);
nand U174 (N_174,In_284,In_428);
or U175 (N_175,In_911,In_622);
or U176 (N_176,In_704,In_868);
or U177 (N_177,In_889,In_159);
nor U178 (N_178,In_480,In_390);
and U179 (N_179,In_923,In_18);
or U180 (N_180,In_58,In_926);
and U181 (N_181,In_531,In_752);
or U182 (N_182,In_76,In_798);
or U183 (N_183,In_913,In_567);
and U184 (N_184,In_328,In_723);
and U185 (N_185,In_399,In_148);
nor U186 (N_186,In_67,In_860);
and U187 (N_187,In_599,In_418);
nand U188 (N_188,In_581,In_853);
nand U189 (N_189,In_556,In_807);
or U190 (N_190,In_488,In_74);
nor U191 (N_191,In_653,In_693);
nor U192 (N_192,In_440,In_600);
nor U193 (N_193,In_394,In_339);
nor U194 (N_194,In_869,In_507);
nor U195 (N_195,In_575,In_111);
nand U196 (N_196,In_181,In_504);
or U197 (N_197,In_297,In_861);
and U198 (N_198,In_201,In_797);
nor U199 (N_199,In_694,In_219);
and U200 (N_200,In_996,In_837);
nor U201 (N_201,In_542,In_839);
nor U202 (N_202,In_468,In_879);
and U203 (N_203,In_171,In_430);
or U204 (N_204,In_601,In_858);
or U205 (N_205,In_338,In_512);
nor U206 (N_206,In_446,In_467);
nor U207 (N_207,In_904,In_363);
or U208 (N_208,In_453,In_165);
nor U209 (N_209,In_408,In_130);
or U210 (N_210,In_12,In_47);
or U211 (N_211,In_513,In_370);
nor U212 (N_212,In_822,In_291);
or U213 (N_213,In_421,In_702);
nand U214 (N_214,In_604,In_577);
and U215 (N_215,In_127,In_175);
or U216 (N_216,In_659,In_758);
and U217 (N_217,In_168,In_145);
nand U218 (N_218,In_277,In_454);
or U219 (N_219,In_384,In_24);
nor U220 (N_220,In_963,In_470);
nand U221 (N_221,In_35,In_220);
nand U222 (N_222,In_665,In_143);
and U223 (N_223,In_244,In_309);
and U224 (N_224,In_698,In_200);
nor U225 (N_225,In_257,In_910);
and U226 (N_226,In_552,In_503);
nor U227 (N_227,In_534,In_832);
and U228 (N_228,In_750,In_118);
nor U229 (N_229,In_627,In_222);
nor U230 (N_230,In_662,In_481);
nand U231 (N_231,In_258,In_407);
nand U232 (N_232,In_652,In_20);
nor U233 (N_233,In_778,In_445);
nand U234 (N_234,In_178,In_734);
or U235 (N_235,In_709,In_373);
or U236 (N_236,In_707,In_463);
and U237 (N_237,In_856,In_189);
nor U238 (N_238,In_551,In_710);
nand U239 (N_239,In_173,In_252);
nor U240 (N_240,In_177,In_897);
nor U241 (N_241,In_635,In_506);
or U242 (N_242,In_585,In_167);
or U243 (N_243,In_610,In_176);
nor U244 (N_244,In_745,In_383);
or U245 (N_245,In_457,In_701);
nand U246 (N_246,In_350,In_406);
nand U247 (N_247,In_529,In_540);
nand U248 (N_248,In_42,In_715);
or U249 (N_249,In_593,In_54);
and U250 (N_250,In_387,In_154);
xnor U251 (N_251,In_944,In_103);
nor U252 (N_252,In_388,In_224);
and U253 (N_253,In_366,In_571);
nand U254 (N_254,In_632,In_937);
nor U255 (N_255,In_787,In_207);
nand U256 (N_256,In_211,In_135);
or U257 (N_257,In_713,In_845);
nand U258 (N_258,In_342,In_426);
nand U259 (N_259,In_835,In_275);
nor U260 (N_260,In_742,In_855);
or U261 (N_261,In_153,In_302);
and U262 (N_262,In_254,In_401);
and U263 (N_263,In_870,In_249);
nand U264 (N_264,In_509,In_553);
nor U265 (N_265,In_683,In_233);
nand U266 (N_266,In_649,In_951);
or U267 (N_267,In_519,In_642);
and U268 (N_268,In_239,In_27);
and U269 (N_269,In_901,In_814);
nor U270 (N_270,In_184,In_744);
and U271 (N_271,In_152,In_666);
and U272 (N_272,In_246,In_266);
xnor U273 (N_273,In_2,In_79);
nand U274 (N_274,In_372,In_826);
and U275 (N_275,In_133,In_308);
nand U276 (N_276,In_574,In_638);
or U277 (N_277,In_925,In_851);
and U278 (N_278,In_785,In_166);
or U279 (N_279,In_283,In_579);
nand U280 (N_280,In_908,In_811);
nor U281 (N_281,In_203,In_136);
nor U282 (N_282,In_205,In_476);
nand U283 (N_283,In_893,In_708);
nor U284 (N_284,In_429,In_397);
nand U285 (N_285,In_933,In_304);
and U286 (N_286,In_121,In_482);
nand U287 (N_287,In_53,In_838);
xor U288 (N_288,In_836,In_7);
or U289 (N_289,In_8,In_413);
nand U290 (N_290,In_281,In_625);
nor U291 (N_291,In_809,In_566);
nand U292 (N_292,In_160,In_730);
nand U293 (N_293,In_286,In_335);
and U294 (N_294,In_196,In_369);
or U295 (N_295,In_323,In_796);
or U296 (N_296,In_458,In_157);
and U297 (N_297,In_596,In_149);
nand U298 (N_298,In_806,In_170);
or U299 (N_299,In_682,In_499);
or U300 (N_300,In_914,In_208);
nand U301 (N_301,In_747,In_918);
nor U302 (N_302,In_442,In_38);
nor U303 (N_303,In_539,In_692);
or U304 (N_304,In_916,In_462);
nor U305 (N_305,In_502,In_237);
nand U306 (N_306,In_801,In_508);
and U307 (N_307,In_623,In_23);
or U308 (N_308,In_528,In_381);
and U309 (N_309,In_991,In_711);
nand U310 (N_310,In_344,In_977);
nand U311 (N_311,In_456,In_882);
or U312 (N_312,In_0,In_134);
nor U313 (N_313,In_293,In_763);
nand U314 (N_314,In_45,In_896);
and U315 (N_315,In_890,In_721);
xnor U316 (N_316,In_324,In_543);
nand U317 (N_317,In_374,In_371);
or U318 (N_318,In_206,In_792);
and U319 (N_319,In_978,In_477);
or U320 (N_320,In_941,In_559);
nand U321 (N_321,In_828,In_591);
nor U322 (N_322,In_706,In_568);
nand U323 (N_323,In_276,In_367);
nand U324 (N_324,In_962,In_278);
or U325 (N_325,In_174,In_70);
nand U326 (N_326,In_427,In_685);
or U327 (N_327,In_808,In_597);
nand U328 (N_328,In_195,In_953);
and U329 (N_329,In_141,In_637);
or U330 (N_330,In_887,In_155);
nor U331 (N_331,In_983,In_63);
or U332 (N_332,In_939,In_340);
nor U333 (N_333,In_621,In_645);
nor U334 (N_334,In_279,In_272);
and U335 (N_335,In_561,In_788);
nor U336 (N_336,In_656,In_606);
nand U337 (N_337,In_647,In_210);
or U338 (N_338,In_321,In_64);
nand U339 (N_339,In_733,In_738);
or U340 (N_340,In_841,In_768);
nor U341 (N_341,In_984,In_686);
and U342 (N_342,In_866,In_423);
and U343 (N_343,In_299,In_892);
nor U344 (N_344,In_164,In_433);
nand U345 (N_345,In_959,In_562);
and U346 (N_346,In_115,In_843);
nor U347 (N_347,In_618,In_774);
nor U348 (N_348,In_287,In_329);
nand U349 (N_349,In_781,In_227);
or U350 (N_350,In_614,In_717);
and U351 (N_351,In_475,In_85);
or U352 (N_352,In_41,In_57);
and U353 (N_353,In_678,In_590);
or U354 (N_354,In_469,In_732);
or U355 (N_355,In_46,In_697);
and U356 (N_356,In_522,In_449);
or U357 (N_357,In_564,In_90);
or U358 (N_358,In_234,In_675);
and U359 (N_359,In_221,In_3);
nand U360 (N_360,In_932,In_188);
and U361 (N_361,In_466,In_151);
and U362 (N_362,In_793,In_414);
nand U363 (N_363,In_663,In_560);
nor U364 (N_364,In_846,In_105);
nor U365 (N_365,In_955,In_679);
nor U366 (N_366,In_424,In_992);
nand U367 (N_367,In_491,In_735);
and U368 (N_368,In_636,In_419);
or U369 (N_369,In_831,In_56);
and U370 (N_370,In_676,In_126);
nor U371 (N_371,In_236,In_523);
or U372 (N_372,In_156,In_494);
and U373 (N_373,In_550,In_871);
nor U374 (N_374,In_355,In_461);
nand U375 (N_375,In_957,In_465);
nand U376 (N_376,In_198,In_929);
nand U377 (N_377,In_66,In_163);
and U378 (N_378,In_298,In_726);
or U379 (N_379,In_820,In_75);
and U380 (N_380,In_452,In_36);
nand U381 (N_381,In_190,In_940);
or U382 (N_382,In_310,In_884);
nor U383 (N_383,In_749,In_486);
nand U384 (N_384,In_549,In_25);
nor U385 (N_385,In_716,In_881);
or U386 (N_386,In_34,In_648);
or U387 (N_387,In_253,In_612);
nor U388 (N_388,In_651,In_187);
nor U389 (N_389,In_840,In_949);
nor U390 (N_390,In_5,In_485);
and U391 (N_391,In_260,In_400);
nand U392 (N_392,In_455,In_640);
and U393 (N_393,In_229,In_514);
nand U394 (N_394,In_60,In_409);
nor U395 (N_395,In_162,In_687);
nor U396 (N_396,In_681,In_270);
and U397 (N_397,In_862,In_595);
nor U398 (N_398,In_532,In_132);
nand U399 (N_399,In_240,In_361);
nor U400 (N_400,In_194,In_393);
or U401 (N_401,In_117,In_255);
nand U402 (N_402,In_993,In_672);
nand U403 (N_403,In_875,In_341);
and U404 (N_404,In_274,In_109);
nand U405 (N_405,In_775,In_688);
nand U406 (N_406,In_31,In_974);
or U407 (N_407,In_938,In_52);
nand U408 (N_408,In_314,In_140);
nand U409 (N_409,In_934,In_81);
nand U410 (N_410,In_578,In_9);
nor U411 (N_411,In_17,In_336);
xor U412 (N_412,In_554,In_472);
nor U413 (N_413,In_780,In_269);
and U414 (N_414,In_95,In_385);
nor U415 (N_415,In_883,In_359);
or U416 (N_416,In_915,In_392);
or U417 (N_417,In_842,In_447);
or U418 (N_418,In_864,In_251);
nand U419 (N_419,In_794,In_241);
and U420 (N_420,In_412,In_557);
nor U421 (N_421,In_582,In_587);
nand U422 (N_422,In_396,In_740);
or U423 (N_423,In_82,In_294);
nand U424 (N_424,In_728,In_242);
nor U425 (N_425,In_873,In_501);
nor U426 (N_426,In_565,In_746);
nand U427 (N_427,In_626,In_108);
nand U428 (N_428,In_349,In_736);
nand U429 (N_429,In_863,In_967);
nand U430 (N_430,In_586,In_670);
nand U431 (N_431,In_905,In_764);
or U432 (N_432,In_757,In_172);
nor U433 (N_433,In_30,In_376);
and U434 (N_434,In_877,In_99);
nor U435 (N_435,In_431,In_852);
nand U436 (N_436,In_73,In_104);
and U437 (N_437,In_516,In_334);
nor U438 (N_438,In_545,In_609);
or U439 (N_439,In_285,In_769);
nand U440 (N_440,In_71,In_548);
and U441 (N_441,In_859,In_546);
nor U442 (N_442,In_59,In_300);
xor U443 (N_443,In_825,In_97);
nor U444 (N_444,In_28,In_634);
nand U445 (N_445,In_438,In_919);
and U446 (N_446,In_62,In_288);
nor U447 (N_447,In_643,In_790);
nand U448 (N_448,In_878,In_515);
nor U449 (N_449,In_795,In_386);
and U450 (N_450,In_498,In_743);
or U451 (N_451,In_55,In_680);
nor U452 (N_452,In_583,In_754);
nor U453 (N_453,In_720,In_225);
and U454 (N_454,In_100,In_1);
and U455 (N_455,In_402,In_292);
or U456 (N_456,In_518,In_493);
or U457 (N_457,In_116,In_660);
nand U458 (N_458,In_495,In_524);
nand U459 (N_459,In_616,In_32);
nand U460 (N_460,In_684,In_212);
and U461 (N_461,In_86,In_611);
or U462 (N_462,In_460,In_238);
or U463 (N_463,In_972,In_521);
nand U464 (N_464,In_98,In_718);
nor U465 (N_465,In_969,In_563);
or U466 (N_466,In_248,In_147);
and U467 (N_467,In_802,In_830);
nor U468 (N_468,In_971,In_61);
nor U469 (N_469,In_129,In_771);
and U470 (N_470,In_169,In_120);
and U471 (N_471,In_84,In_264);
and U472 (N_472,In_829,In_209);
nand U473 (N_473,In_319,In_945);
or U474 (N_474,In_265,In_102);
or U475 (N_475,In_952,In_909);
or U476 (N_476,In_767,In_113);
nand U477 (N_477,In_405,In_139);
and U478 (N_478,In_981,In_724);
nor U479 (N_479,In_677,In_783);
nand U480 (N_480,In_382,In_131);
or U481 (N_481,In_94,In_624);
nor U482 (N_482,In_712,In_947);
nor U483 (N_483,In_511,In_850);
or U484 (N_484,In_354,In_464);
and U485 (N_485,In_930,In_123);
nor U486 (N_486,In_527,In_573);
nor U487 (N_487,In_360,In_827);
and U488 (N_488,In_954,In_448);
nand U489 (N_489,In_703,In_917);
and U490 (N_490,In_271,In_348);
and U491 (N_491,In_124,In_605);
or U492 (N_492,In_37,In_580);
nor U493 (N_493,In_375,In_434);
or U494 (N_494,In_443,In_51);
and U495 (N_495,In_748,In_779);
nor U496 (N_496,In_235,In_849);
or U497 (N_497,In_214,In_821);
or U498 (N_498,In_380,In_44);
nand U499 (N_499,In_990,In_641);
and U500 (N_500,In_824,In_52);
and U501 (N_501,In_41,In_953);
nor U502 (N_502,In_395,In_313);
and U503 (N_503,In_403,In_439);
nor U504 (N_504,In_343,In_130);
or U505 (N_505,In_700,In_207);
xnor U506 (N_506,In_714,In_385);
or U507 (N_507,In_793,In_608);
and U508 (N_508,In_975,In_276);
or U509 (N_509,In_733,In_969);
nand U510 (N_510,In_832,In_481);
or U511 (N_511,In_734,In_636);
nand U512 (N_512,In_641,In_414);
or U513 (N_513,In_285,In_801);
and U514 (N_514,In_307,In_456);
and U515 (N_515,In_222,In_115);
or U516 (N_516,In_918,In_243);
nor U517 (N_517,In_499,In_296);
nor U518 (N_518,In_3,In_39);
and U519 (N_519,In_593,In_442);
nor U520 (N_520,In_167,In_998);
and U521 (N_521,In_159,In_947);
nor U522 (N_522,In_298,In_508);
nor U523 (N_523,In_680,In_131);
nor U524 (N_524,In_487,In_774);
and U525 (N_525,In_608,In_36);
nand U526 (N_526,In_630,In_730);
nor U527 (N_527,In_179,In_857);
or U528 (N_528,In_110,In_337);
nor U529 (N_529,In_535,In_744);
xor U530 (N_530,In_977,In_16);
nor U531 (N_531,In_351,In_96);
or U532 (N_532,In_509,In_217);
or U533 (N_533,In_656,In_564);
nand U534 (N_534,In_815,In_629);
nor U535 (N_535,In_256,In_660);
or U536 (N_536,In_667,In_382);
nand U537 (N_537,In_594,In_448);
nor U538 (N_538,In_346,In_527);
nand U539 (N_539,In_918,In_806);
or U540 (N_540,In_406,In_701);
or U541 (N_541,In_709,In_273);
nor U542 (N_542,In_386,In_40);
or U543 (N_543,In_98,In_92);
nor U544 (N_544,In_556,In_229);
and U545 (N_545,In_943,In_713);
or U546 (N_546,In_787,In_467);
nand U547 (N_547,In_879,In_706);
nor U548 (N_548,In_235,In_417);
nor U549 (N_549,In_516,In_307);
nor U550 (N_550,In_483,In_345);
and U551 (N_551,In_927,In_267);
nand U552 (N_552,In_36,In_763);
nor U553 (N_553,In_568,In_254);
nor U554 (N_554,In_181,In_450);
and U555 (N_555,In_915,In_837);
nand U556 (N_556,In_955,In_800);
and U557 (N_557,In_176,In_878);
or U558 (N_558,In_543,In_620);
nand U559 (N_559,In_314,In_360);
and U560 (N_560,In_183,In_697);
or U561 (N_561,In_856,In_544);
and U562 (N_562,In_516,In_666);
nor U563 (N_563,In_340,In_209);
and U564 (N_564,In_577,In_607);
and U565 (N_565,In_580,In_497);
nor U566 (N_566,In_238,In_210);
nand U567 (N_567,In_285,In_575);
nand U568 (N_568,In_739,In_433);
or U569 (N_569,In_3,In_539);
nand U570 (N_570,In_858,In_741);
and U571 (N_571,In_909,In_290);
nand U572 (N_572,In_770,In_488);
nor U573 (N_573,In_343,In_811);
nor U574 (N_574,In_702,In_536);
nand U575 (N_575,In_105,In_188);
or U576 (N_576,In_969,In_62);
and U577 (N_577,In_705,In_823);
nand U578 (N_578,In_609,In_946);
nand U579 (N_579,In_61,In_389);
nor U580 (N_580,In_163,In_404);
and U581 (N_581,In_280,In_797);
nand U582 (N_582,In_675,In_223);
and U583 (N_583,In_606,In_826);
nand U584 (N_584,In_469,In_176);
and U585 (N_585,In_169,In_720);
nand U586 (N_586,In_367,In_517);
nand U587 (N_587,In_370,In_607);
nand U588 (N_588,In_238,In_597);
nand U589 (N_589,In_239,In_807);
nand U590 (N_590,In_99,In_491);
nand U591 (N_591,In_753,In_809);
nand U592 (N_592,In_428,In_188);
or U593 (N_593,In_804,In_937);
or U594 (N_594,In_333,In_157);
nor U595 (N_595,In_549,In_675);
or U596 (N_596,In_117,In_684);
or U597 (N_597,In_564,In_242);
or U598 (N_598,In_454,In_153);
nand U599 (N_599,In_625,In_699);
and U600 (N_600,In_474,In_666);
nor U601 (N_601,In_23,In_977);
and U602 (N_602,In_556,In_929);
nand U603 (N_603,In_298,In_660);
and U604 (N_604,In_719,In_267);
or U605 (N_605,In_734,In_598);
and U606 (N_606,In_971,In_884);
nor U607 (N_607,In_130,In_500);
and U608 (N_608,In_277,In_715);
and U609 (N_609,In_885,In_193);
nand U610 (N_610,In_935,In_715);
or U611 (N_611,In_888,In_550);
nand U612 (N_612,In_284,In_996);
and U613 (N_613,In_144,In_524);
or U614 (N_614,In_991,In_832);
or U615 (N_615,In_990,In_683);
nand U616 (N_616,In_423,In_685);
or U617 (N_617,In_779,In_103);
nor U618 (N_618,In_847,In_534);
nor U619 (N_619,In_608,In_152);
nor U620 (N_620,In_5,In_472);
nand U621 (N_621,In_853,In_719);
nand U622 (N_622,In_479,In_820);
nand U623 (N_623,In_756,In_624);
nand U624 (N_624,In_899,In_709);
nor U625 (N_625,In_919,In_841);
nand U626 (N_626,In_534,In_453);
nand U627 (N_627,In_374,In_817);
nand U628 (N_628,In_860,In_660);
nor U629 (N_629,In_934,In_815);
and U630 (N_630,In_776,In_434);
and U631 (N_631,In_474,In_665);
and U632 (N_632,In_387,In_110);
and U633 (N_633,In_839,In_712);
and U634 (N_634,In_44,In_660);
or U635 (N_635,In_906,In_246);
and U636 (N_636,In_362,In_352);
nand U637 (N_637,In_475,In_247);
or U638 (N_638,In_812,In_895);
or U639 (N_639,In_740,In_728);
or U640 (N_640,In_1,In_264);
or U641 (N_641,In_136,In_38);
and U642 (N_642,In_790,In_58);
and U643 (N_643,In_574,In_479);
nor U644 (N_644,In_500,In_339);
nand U645 (N_645,In_714,In_191);
nand U646 (N_646,In_661,In_972);
and U647 (N_647,In_150,In_208);
or U648 (N_648,In_380,In_952);
and U649 (N_649,In_194,In_603);
or U650 (N_650,In_735,In_347);
or U651 (N_651,In_582,In_324);
or U652 (N_652,In_677,In_461);
xnor U653 (N_653,In_53,In_438);
or U654 (N_654,In_543,In_809);
or U655 (N_655,In_148,In_900);
nor U656 (N_656,In_836,In_245);
nor U657 (N_657,In_681,In_305);
or U658 (N_658,In_847,In_732);
or U659 (N_659,In_400,In_78);
nand U660 (N_660,In_177,In_204);
nor U661 (N_661,In_80,In_992);
and U662 (N_662,In_716,In_745);
nand U663 (N_663,In_604,In_705);
or U664 (N_664,In_608,In_947);
and U665 (N_665,In_351,In_845);
or U666 (N_666,In_998,In_436);
or U667 (N_667,In_532,In_11);
nor U668 (N_668,In_98,In_129);
nand U669 (N_669,In_481,In_251);
or U670 (N_670,In_323,In_272);
nand U671 (N_671,In_376,In_712);
or U672 (N_672,In_693,In_47);
and U673 (N_673,In_789,In_990);
or U674 (N_674,In_357,In_20);
nand U675 (N_675,In_481,In_943);
and U676 (N_676,In_129,In_999);
or U677 (N_677,In_483,In_904);
and U678 (N_678,In_414,In_39);
or U679 (N_679,In_943,In_361);
and U680 (N_680,In_312,In_266);
and U681 (N_681,In_215,In_667);
or U682 (N_682,In_475,In_822);
or U683 (N_683,In_715,In_61);
nand U684 (N_684,In_564,In_602);
nor U685 (N_685,In_883,In_193);
nand U686 (N_686,In_879,In_792);
nand U687 (N_687,In_126,In_951);
or U688 (N_688,In_875,In_49);
or U689 (N_689,In_4,In_400);
nor U690 (N_690,In_468,In_486);
nor U691 (N_691,In_784,In_140);
nor U692 (N_692,In_453,In_824);
nor U693 (N_693,In_127,In_884);
or U694 (N_694,In_926,In_769);
and U695 (N_695,In_851,In_481);
nand U696 (N_696,In_532,In_381);
nor U697 (N_697,In_706,In_992);
nand U698 (N_698,In_977,In_406);
nand U699 (N_699,In_53,In_942);
and U700 (N_700,In_176,In_384);
nor U701 (N_701,In_800,In_894);
and U702 (N_702,In_491,In_570);
and U703 (N_703,In_162,In_917);
nor U704 (N_704,In_972,In_771);
nand U705 (N_705,In_876,In_675);
or U706 (N_706,In_936,In_506);
nor U707 (N_707,In_427,In_730);
nand U708 (N_708,In_632,In_357);
nand U709 (N_709,In_943,In_336);
nand U710 (N_710,In_468,In_152);
nand U711 (N_711,In_415,In_697);
and U712 (N_712,In_311,In_991);
nand U713 (N_713,In_262,In_296);
nor U714 (N_714,In_125,In_861);
nand U715 (N_715,In_440,In_906);
or U716 (N_716,In_323,In_470);
and U717 (N_717,In_468,In_401);
and U718 (N_718,In_195,In_878);
nand U719 (N_719,In_144,In_104);
or U720 (N_720,In_212,In_70);
nor U721 (N_721,In_984,In_171);
or U722 (N_722,In_337,In_954);
nor U723 (N_723,In_72,In_6);
nand U724 (N_724,In_893,In_17);
or U725 (N_725,In_714,In_754);
or U726 (N_726,In_949,In_824);
nand U727 (N_727,In_360,In_363);
nor U728 (N_728,In_232,In_810);
nor U729 (N_729,In_74,In_470);
nor U730 (N_730,In_29,In_465);
xnor U731 (N_731,In_541,In_952);
and U732 (N_732,In_403,In_554);
nand U733 (N_733,In_182,In_726);
or U734 (N_734,In_922,In_137);
nor U735 (N_735,In_577,In_305);
or U736 (N_736,In_995,In_688);
or U737 (N_737,In_639,In_507);
nor U738 (N_738,In_37,In_464);
or U739 (N_739,In_699,In_272);
or U740 (N_740,In_454,In_210);
or U741 (N_741,In_653,In_277);
nand U742 (N_742,In_758,In_3);
nor U743 (N_743,In_651,In_871);
nand U744 (N_744,In_423,In_202);
nand U745 (N_745,In_431,In_611);
and U746 (N_746,In_954,In_373);
nand U747 (N_747,In_346,In_149);
nor U748 (N_748,In_413,In_836);
nor U749 (N_749,In_288,In_798);
or U750 (N_750,In_179,In_431);
and U751 (N_751,In_341,In_736);
or U752 (N_752,In_73,In_267);
nor U753 (N_753,In_104,In_983);
and U754 (N_754,In_942,In_586);
or U755 (N_755,In_392,In_206);
nand U756 (N_756,In_788,In_631);
nor U757 (N_757,In_596,In_739);
nor U758 (N_758,In_114,In_699);
and U759 (N_759,In_516,In_760);
and U760 (N_760,In_348,In_919);
or U761 (N_761,In_898,In_592);
nor U762 (N_762,In_248,In_770);
or U763 (N_763,In_794,In_496);
and U764 (N_764,In_717,In_15);
nor U765 (N_765,In_118,In_625);
nand U766 (N_766,In_723,In_90);
or U767 (N_767,In_326,In_859);
or U768 (N_768,In_66,In_391);
and U769 (N_769,In_926,In_798);
nand U770 (N_770,In_267,In_206);
nand U771 (N_771,In_541,In_821);
nand U772 (N_772,In_440,In_388);
nor U773 (N_773,In_676,In_421);
nor U774 (N_774,In_894,In_464);
or U775 (N_775,In_636,In_515);
nor U776 (N_776,In_508,In_214);
nor U777 (N_777,In_325,In_169);
or U778 (N_778,In_951,In_754);
or U779 (N_779,In_77,In_850);
and U780 (N_780,In_733,In_668);
nand U781 (N_781,In_834,In_91);
nor U782 (N_782,In_347,In_993);
or U783 (N_783,In_675,In_856);
nor U784 (N_784,In_453,In_433);
nor U785 (N_785,In_840,In_125);
xor U786 (N_786,In_684,In_706);
and U787 (N_787,In_148,In_947);
nand U788 (N_788,In_613,In_490);
or U789 (N_789,In_930,In_611);
and U790 (N_790,In_985,In_805);
nor U791 (N_791,In_384,In_440);
or U792 (N_792,In_966,In_815);
nand U793 (N_793,In_569,In_154);
and U794 (N_794,In_879,In_723);
nor U795 (N_795,In_874,In_649);
or U796 (N_796,In_881,In_944);
or U797 (N_797,In_199,In_782);
and U798 (N_798,In_567,In_695);
nand U799 (N_799,In_429,In_95);
and U800 (N_800,In_177,In_223);
or U801 (N_801,In_89,In_112);
nand U802 (N_802,In_814,In_451);
nand U803 (N_803,In_134,In_786);
and U804 (N_804,In_793,In_370);
and U805 (N_805,In_822,In_152);
and U806 (N_806,In_92,In_392);
nand U807 (N_807,In_825,In_402);
nand U808 (N_808,In_535,In_921);
nor U809 (N_809,In_771,In_134);
nand U810 (N_810,In_41,In_37);
nor U811 (N_811,In_885,In_307);
and U812 (N_812,In_342,In_712);
nor U813 (N_813,In_563,In_682);
nand U814 (N_814,In_290,In_52);
and U815 (N_815,In_732,In_617);
nor U816 (N_816,In_125,In_737);
nor U817 (N_817,In_495,In_44);
or U818 (N_818,In_746,In_987);
and U819 (N_819,In_205,In_659);
nand U820 (N_820,In_712,In_119);
or U821 (N_821,In_27,In_598);
nor U822 (N_822,In_515,In_214);
or U823 (N_823,In_786,In_640);
and U824 (N_824,In_352,In_687);
nor U825 (N_825,In_971,In_575);
nor U826 (N_826,In_719,In_221);
and U827 (N_827,In_485,In_798);
nor U828 (N_828,In_956,In_381);
or U829 (N_829,In_527,In_546);
nand U830 (N_830,In_457,In_393);
or U831 (N_831,In_444,In_521);
and U832 (N_832,In_843,In_299);
and U833 (N_833,In_121,In_290);
or U834 (N_834,In_759,In_608);
or U835 (N_835,In_425,In_410);
and U836 (N_836,In_0,In_687);
and U837 (N_837,In_421,In_390);
and U838 (N_838,In_227,In_210);
nor U839 (N_839,In_650,In_27);
or U840 (N_840,In_754,In_742);
and U841 (N_841,In_331,In_134);
nor U842 (N_842,In_71,In_867);
or U843 (N_843,In_558,In_898);
and U844 (N_844,In_715,In_243);
nand U845 (N_845,In_878,In_158);
and U846 (N_846,In_279,In_646);
nand U847 (N_847,In_746,In_293);
nand U848 (N_848,In_479,In_406);
and U849 (N_849,In_63,In_369);
or U850 (N_850,In_499,In_20);
or U851 (N_851,In_607,In_255);
or U852 (N_852,In_339,In_378);
nand U853 (N_853,In_458,In_858);
or U854 (N_854,In_323,In_222);
xnor U855 (N_855,In_725,In_608);
or U856 (N_856,In_146,In_772);
and U857 (N_857,In_371,In_485);
and U858 (N_858,In_769,In_161);
and U859 (N_859,In_872,In_316);
or U860 (N_860,In_485,In_612);
nand U861 (N_861,In_645,In_889);
nand U862 (N_862,In_427,In_64);
and U863 (N_863,In_476,In_498);
or U864 (N_864,In_227,In_348);
or U865 (N_865,In_288,In_25);
nand U866 (N_866,In_931,In_220);
and U867 (N_867,In_497,In_225);
and U868 (N_868,In_617,In_711);
and U869 (N_869,In_123,In_811);
nand U870 (N_870,In_495,In_232);
nor U871 (N_871,In_876,In_425);
or U872 (N_872,In_656,In_147);
or U873 (N_873,In_346,In_626);
and U874 (N_874,In_668,In_332);
and U875 (N_875,In_825,In_464);
or U876 (N_876,In_151,In_378);
nor U877 (N_877,In_265,In_321);
nand U878 (N_878,In_702,In_447);
xor U879 (N_879,In_263,In_810);
or U880 (N_880,In_436,In_805);
and U881 (N_881,In_483,In_744);
and U882 (N_882,In_673,In_395);
nand U883 (N_883,In_159,In_205);
nand U884 (N_884,In_276,In_830);
and U885 (N_885,In_268,In_166);
nor U886 (N_886,In_19,In_794);
nor U887 (N_887,In_845,In_333);
nand U888 (N_888,In_914,In_879);
nand U889 (N_889,In_635,In_840);
and U890 (N_890,In_834,In_579);
or U891 (N_891,In_127,In_434);
and U892 (N_892,In_110,In_847);
nand U893 (N_893,In_807,In_406);
and U894 (N_894,In_744,In_845);
nor U895 (N_895,In_914,In_745);
nand U896 (N_896,In_380,In_891);
and U897 (N_897,In_995,In_240);
and U898 (N_898,In_757,In_667);
nor U899 (N_899,In_53,In_552);
or U900 (N_900,In_499,In_581);
and U901 (N_901,In_536,In_360);
and U902 (N_902,In_50,In_483);
nand U903 (N_903,In_851,In_120);
and U904 (N_904,In_542,In_923);
and U905 (N_905,In_543,In_106);
and U906 (N_906,In_889,In_213);
nand U907 (N_907,In_802,In_94);
and U908 (N_908,In_719,In_422);
or U909 (N_909,In_670,In_551);
nand U910 (N_910,In_913,In_696);
and U911 (N_911,In_759,In_974);
and U912 (N_912,In_571,In_424);
nand U913 (N_913,In_215,In_869);
or U914 (N_914,In_279,In_529);
and U915 (N_915,In_37,In_971);
nand U916 (N_916,In_753,In_814);
and U917 (N_917,In_851,In_884);
or U918 (N_918,In_31,In_97);
or U919 (N_919,In_561,In_523);
nand U920 (N_920,In_715,In_480);
nor U921 (N_921,In_591,In_312);
xor U922 (N_922,In_593,In_880);
or U923 (N_923,In_39,In_838);
or U924 (N_924,In_409,In_633);
and U925 (N_925,In_529,In_246);
and U926 (N_926,In_901,In_250);
nor U927 (N_927,In_648,In_429);
or U928 (N_928,In_278,In_909);
nor U929 (N_929,In_202,In_162);
nor U930 (N_930,In_960,In_861);
and U931 (N_931,In_74,In_979);
nor U932 (N_932,In_91,In_578);
nor U933 (N_933,In_821,In_170);
and U934 (N_934,In_839,In_593);
or U935 (N_935,In_34,In_209);
and U936 (N_936,In_242,In_357);
and U937 (N_937,In_999,In_67);
nand U938 (N_938,In_514,In_579);
nor U939 (N_939,In_6,In_934);
nor U940 (N_940,In_432,In_100);
nor U941 (N_941,In_419,In_98);
or U942 (N_942,In_804,In_526);
or U943 (N_943,In_440,In_526);
nand U944 (N_944,In_634,In_730);
or U945 (N_945,In_713,In_464);
and U946 (N_946,In_569,In_71);
nand U947 (N_947,In_346,In_300);
and U948 (N_948,In_133,In_138);
and U949 (N_949,In_128,In_638);
nor U950 (N_950,In_695,In_766);
nor U951 (N_951,In_647,In_247);
or U952 (N_952,In_204,In_670);
nand U953 (N_953,In_162,In_76);
nor U954 (N_954,In_478,In_882);
and U955 (N_955,In_221,In_219);
nor U956 (N_956,In_710,In_624);
nand U957 (N_957,In_184,In_589);
and U958 (N_958,In_825,In_684);
nand U959 (N_959,In_945,In_574);
and U960 (N_960,In_445,In_855);
and U961 (N_961,In_244,In_293);
or U962 (N_962,In_689,In_391);
and U963 (N_963,In_416,In_533);
nand U964 (N_964,In_763,In_878);
nor U965 (N_965,In_572,In_517);
xnor U966 (N_966,In_608,In_797);
or U967 (N_967,In_422,In_508);
nand U968 (N_968,In_724,In_907);
or U969 (N_969,In_620,In_895);
or U970 (N_970,In_529,In_899);
nand U971 (N_971,In_914,In_229);
nor U972 (N_972,In_676,In_828);
nand U973 (N_973,In_704,In_93);
nand U974 (N_974,In_780,In_888);
nand U975 (N_975,In_524,In_834);
nor U976 (N_976,In_536,In_565);
and U977 (N_977,In_352,In_179);
nor U978 (N_978,In_795,In_801);
nor U979 (N_979,In_891,In_393);
and U980 (N_980,In_48,In_199);
or U981 (N_981,In_773,In_699);
nand U982 (N_982,In_12,In_56);
or U983 (N_983,In_143,In_635);
nand U984 (N_984,In_749,In_606);
or U985 (N_985,In_275,In_480);
or U986 (N_986,In_991,In_509);
or U987 (N_987,In_630,In_110);
and U988 (N_988,In_181,In_175);
nor U989 (N_989,In_395,In_577);
nor U990 (N_990,In_325,In_869);
and U991 (N_991,In_827,In_436);
nor U992 (N_992,In_327,In_862);
and U993 (N_993,In_327,In_844);
and U994 (N_994,In_45,In_970);
nor U995 (N_995,In_376,In_467);
or U996 (N_996,In_504,In_988);
nand U997 (N_997,In_406,In_5);
nand U998 (N_998,In_285,In_660);
nand U999 (N_999,In_791,In_624);
and U1000 (N_1000,In_281,In_743);
nand U1001 (N_1001,In_660,In_896);
or U1002 (N_1002,In_17,In_522);
nand U1003 (N_1003,In_127,In_629);
nand U1004 (N_1004,In_170,In_135);
nor U1005 (N_1005,In_317,In_882);
or U1006 (N_1006,In_955,In_792);
and U1007 (N_1007,In_296,In_901);
nor U1008 (N_1008,In_710,In_513);
and U1009 (N_1009,In_133,In_215);
nor U1010 (N_1010,In_821,In_513);
nand U1011 (N_1011,In_923,In_264);
nand U1012 (N_1012,In_834,In_818);
and U1013 (N_1013,In_361,In_536);
nand U1014 (N_1014,In_648,In_567);
or U1015 (N_1015,In_729,In_757);
and U1016 (N_1016,In_534,In_350);
or U1017 (N_1017,In_337,In_147);
and U1018 (N_1018,In_198,In_392);
nor U1019 (N_1019,In_630,In_100);
and U1020 (N_1020,In_800,In_661);
and U1021 (N_1021,In_859,In_576);
and U1022 (N_1022,In_998,In_584);
nand U1023 (N_1023,In_791,In_846);
nor U1024 (N_1024,In_87,In_245);
or U1025 (N_1025,In_311,In_207);
or U1026 (N_1026,In_291,In_935);
and U1027 (N_1027,In_257,In_104);
nand U1028 (N_1028,In_84,In_298);
or U1029 (N_1029,In_924,In_426);
nor U1030 (N_1030,In_668,In_352);
or U1031 (N_1031,In_963,In_842);
nand U1032 (N_1032,In_22,In_613);
or U1033 (N_1033,In_139,In_368);
or U1034 (N_1034,In_79,In_543);
or U1035 (N_1035,In_102,In_330);
or U1036 (N_1036,In_199,In_134);
nand U1037 (N_1037,In_701,In_264);
and U1038 (N_1038,In_403,In_416);
nand U1039 (N_1039,In_525,In_961);
nor U1040 (N_1040,In_525,In_114);
nor U1041 (N_1041,In_574,In_120);
and U1042 (N_1042,In_151,In_392);
nand U1043 (N_1043,In_239,In_245);
nand U1044 (N_1044,In_777,In_100);
or U1045 (N_1045,In_276,In_920);
nand U1046 (N_1046,In_841,In_68);
nand U1047 (N_1047,In_511,In_79);
nand U1048 (N_1048,In_494,In_134);
and U1049 (N_1049,In_353,In_596);
nand U1050 (N_1050,In_466,In_212);
or U1051 (N_1051,In_273,In_646);
or U1052 (N_1052,In_83,In_614);
and U1053 (N_1053,In_378,In_683);
and U1054 (N_1054,In_667,In_944);
or U1055 (N_1055,In_657,In_562);
nor U1056 (N_1056,In_680,In_727);
nand U1057 (N_1057,In_290,In_940);
or U1058 (N_1058,In_806,In_223);
nand U1059 (N_1059,In_742,In_250);
and U1060 (N_1060,In_533,In_11);
and U1061 (N_1061,In_485,In_460);
or U1062 (N_1062,In_82,In_783);
or U1063 (N_1063,In_340,In_482);
nand U1064 (N_1064,In_537,In_20);
and U1065 (N_1065,In_949,In_689);
and U1066 (N_1066,In_979,In_736);
nand U1067 (N_1067,In_127,In_130);
nand U1068 (N_1068,In_565,In_137);
nand U1069 (N_1069,In_154,In_485);
nand U1070 (N_1070,In_382,In_409);
nand U1071 (N_1071,In_591,In_587);
and U1072 (N_1072,In_232,In_571);
nand U1073 (N_1073,In_489,In_123);
nor U1074 (N_1074,In_907,In_403);
nand U1075 (N_1075,In_25,In_105);
nor U1076 (N_1076,In_512,In_728);
or U1077 (N_1077,In_164,In_97);
nor U1078 (N_1078,In_771,In_686);
and U1079 (N_1079,In_483,In_265);
nor U1080 (N_1080,In_800,In_946);
nor U1081 (N_1081,In_135,In_563);
and U1082 (N_1082,In_284,In_740);
nand U1083 (N_1083,In_954,In_365);
and U1084 (N_1084,In_708,In_735);
and U1085 (N_1085,In_203,In_879);
nor U1086 (N_1086,In_182,In_1);
or U1087 (N_1087,In_594,In_64);
and U1088 (N_1088,In_265,In_983);
or U1089 (N_1089,In_2,In_703);
and U1090 (N_1090,In_917,In_977);
and U1091 (N_1091,In_211,In_789);
nor U1092 (N_1092,In_313,In_344);
and U1093 (N_1093,In_400,In_597);
nor U1094 (N_1094,In_375,In_59);
nor U1095 (N_1095,In_463,In_573);
and U1096 (N_1096,In_582,In_477);
nand U1097 (N_1097,In_86,In_62);
or U1098 (N_1098,In_325,In_720);
or U1099 (N_1099,In_687,In_635);
and U1100 (N_1100,In_425,In_682);
nand U1101 (N_1101,In_434,In_271);
nor U1102 (N_1102,In_348,In_577);
nor U1103 (N_1103,In_283,In_770);
nand U1104 (N_1104,In_641,In_829);
and U1105 (N_1105,In_508,In_565);
nor U1106 (N_1106,In_119,In_140);
and U1107 (N_1107,In_650,In_765);
nand U1108 (N_1108,In_267,In_724);
and U1109 (N_1109,In_139,In_594);
nor U1110 (N_1110,In_327,In_491);
nand U1111 (N_1111,In_496,In_155);
or U1112 (N_1112,In_425,In_992);
nor U1113 (N_1113,In_275,In_231);
and U1114 (N_1114,In_590,In_184);
and U1115 (N_1115,In_944,In_192);
or U1116 (N_1116,In_222,In_733);
or U1117 (N_1117,In_235,In_559);
nand U1118 (N_1118,In_668,In_448);
nand U1119 (N_1119,In_577,In_991);
nor U1120 (N_1120,In_988,In_73);
and U1121 (N_1121,In_250,In_77);
nor U1122 (N_1122,In_318,In_917);
or U1123 (N_1123,In_921,In_703);
nor U1124 (N_1124,In_898,In_681);
nand U1125 (N_1125,In_194,In_179);
or U1126 (N_1126,In_956,In_859);
and U1127 (N_1127,In_256,In_957);
or U1128 (N_1128,In_389,In_895);
and U1129 (N_1129,In_130,In_156);
nand U1130 (N_1130,In_320,In_885);
nand U1131 (N_1131,In_992,In_548);
or U1132 (N_1132,In_206,In_347);
or U1133 (N_1133,In_546,In_586);
nand U1134 (N_1134,In_551,In_856);
or U1135 (N_1135,In_678,In_396);
or U1136 (N_1136,In_656,In_710);
nor U1137 (N_1137,In_196,In_140);
nand U1138 (N_1138,In_410,In_687);
nor U1139 (N_1139,In_608,In_271);
or U1140 (N_1140,In_926,In_912);
nor U1141 (N_1141,In_555,In_443);
and U1142 (N_1142,In_791,In_567);
or U1143 (N_1143,In_436,In_734);
and U1144 (N_1144,In_953,In_443);
nor U1145 (N_1145,In_411,In_178);
nand U1146 (N_1146,In_22,In_202);
nor U1147 (N_1147,In_135,In_927);
nor U1148 (N_1148,In_493,In_66);
nor U1149 (N_1149,In_290,In_808);
nand U1150 (N_1150,In_496,In_452);
nand U1151 (N_1151,In_894,In_769);
nand U1152 (N_1152,In_801,In_710);
or U1153 (N_1153,In_801,In_544);
nand U1154 (N_1154,In_362,In_702);
and U1155 (N_1155,In_711,In_680);
or U1156 (N_1156,In_265,In_765);
nor U1157 (N_1157,In_484,In_386);
or U1158 (N_1158,In_991,In_657);
and U1159 (N_1159,In_356,In_169);
nor U1160 (N_1160,In_960,In_820);
nand U1161 (N_1161,In_878,In_524);
nand U1162 (N_1162,In_201,In_602);
nor U1163 (N_1163,In_702,In_16);
xor U1164 (N_1164,In_341,In_991);
nor U1165 (N_1165,In_707,In_860);
nor U1166 (N_1166,In_140,In_398);
or U1167 (N_1167,In_598,In_143);
and U1168 (N_1168,In_733,In_130);
nor U1169 (N_1169,In_547,In_68);
nor U1170 (N_1170,In_203,In_428);
and U1171 (N_1171,In_269,In_214);
or U1172 (N_1172,In_348,In_232);
or U1173 (N_1173,In_634,In_333);
nand U1174 (N_1174,In_644,In_414);
or U1175 (N_1175,In_580,In_369);
nand U1176 (N_1176,In_651,In_230);
and U1177 (N_1177,In_877,In_945);
nand U1178 (N_1178,In_222,In_289);
nor U1179 (N_1179,In_844,In_207);
and U1180 (N_1180,In_333,In_318);
nand U1181 (N_1181,In_877,In_20);
and U1182 (N_1182,In_292,In_932);
or U1183 (N_1183,In_817,In_570);
and U1184 (N_1184,In_69,In_99);
and U1185 (N_1185,In_476,In_22);
and U1186 (N_1186,In_834,In_512);
nor U1187 (N_1187,In_601,In_709);
and U1188 (N_1188,In_778,In_126);
or U1189 (N_1189,In_383,In_572);
nand U1190 (N_1190,In_995,In_194);
or U1191 (N_1191,In_376,In_942);
nand U1192 (N_1192,In_139,In_926);
nor U1193 (N_1193,In_598,In_294);
or U1194 (N_1194,In_615,In_85);
or U1195 (N_1195,In_210,In_593);
nand U1196 (N_1196,In_26,In_878);
nand U1197 (N_1197,In_483,In_437);
nand U1198 (N_1198,In_643,In_264);
or U1199 (N_1199,In_481,In_766);
nand U1200 (N_1200,In_895,In_829);
nand U1201 (N_1201,In_753,In_475);
xor U1202 (N_1202,In_30,In_855);
and U1203 (N_1203,In_318,In_567);
or U1204 (N_1204,In_83,In_55);
nor U1205 (N_1205,In_577,In_573);
nor U1206 (N_1206,In_378,In_579);
nand U1207 (N_1207,In_504,In_222);
nand U1208 (N_1208,In_551,In_330);
nand U1209 (N_1209,In_1,In_436);
nand U1210 (N_1210,In_900,In_747);
nand U1211 (N_1211,In_63,In_15);
nand U1212 (N_1212,In_453,In_386);
and U1213 (N_1213,In_289,In_879);
or U1214 (N_1214,In_228,In_69);
or U1215 (N_1215,In_809,In_482);
nor U1216 (N_1216,In_331,In_194);
nand U1217 (N_1217,In_246,In_847);
and U1218 (N_1218,In_152,In_272);
nor U1219 (N_1219,In_119,In_22);
nand U1220 (N_1220,In_249,In_366);
nand U1221 (N_1221,In_947,In_914);
nor U1222 (N_1222,In_229,In_825);
nor U1223 (N_1223,In_112,In_58);
nor U1224 (N_1224,In_760,In_535);
or U1225 (N_1225,In_58,In_260);
nor U1226 (N_1226,In_843,In_298);
nor U1227 (N_1227,In_209,In_690);
or U1228 (N_1228,In_572,In_580);
or U1229 (N_1229,In_56,In_487);
nor U1230 (N_1230,In_503,In_492);
or U1231 (N_1231,In_208,In_472);
xnor U1232 (N_1232,In_249,In_946);
or U1233 (N_1233,In_300,In_251);
or U1234 (N_1234,In_193,In_147);
nor U1235 (N_1235,In_711,In_367);
or U1236 (N_1236,In_598,In_841);
or U1237 (N_1237,In_265,In_784);
xor U1238 (N_1238,In_190,In_520);
nand U1239 (N_1239,In_941,In_274);
and U1240 (N_1240,In_443,In_309);
or U1241 (N_1241,In_329,In_295);
and U1242 (N_1242,In_114,In_591);
nand U1243 (N_1243,In_57,In_724);
nand U1244 (N_1244,In_137,In_819);
and U1245 (N_1245,In_265,In_979);
and U1246 (N_1246,In_195,In_836);
and U1247 (N_1247,In_178,In_446);
and U1248 (N_1248,In_255,In_109);
and U1249 (N_1249,In_122,In_198);
nor U1250 (N_1250,In_621,In_477);
nor U1251 (N_1251,In_232,In_968);
and U1252 (N_1252,In_274,In_90);
nand U1253 (N_1253,In_457,In_148);
and U1254 (N_1254,In_595,In_195);
or U1255 (N_1255,In_430,In_309);
or U1256 (N_1256,In_462,In_713);
or U1257 (N_1257,In_507,In_327);
nor U1258 (N_1258,In_973,In_527);
or U1259 (N_1259,In_629,In_454);
nand U1260 (N_1260,In_88,In_724);
and U1261 (N_1261,In_701,In_517);
or U1262 (N_1262,In_905,In_308);
nor U1263 (N_1263,In_228,In_369);
nor U1264 (N_1264,In_42,In_921);
or U1265 (N_1265,In_609,In_861);
nand U1266 (N_1266,In_554,In_490);
nand U1267 (N_1267,In_145,In_612);
nor U1268 (N_1268,In_422,In_918);
nor U1269 (N_1269,In_326,In_321);
nor U1270 (N_1270,In_389,In_777);
or U1271 (N_1271,In_231,In_732);
nor U1272 (N_1272,In_384,In_491);
nand U1273 (N_1273,In_855,In_556);
nand U1274 (N_1274,In_125,In_283);
or U1275 (N_1275,In_711,In_313);
or U1276 (N_1276,In_182,In_874);
or U1277 (N_1277,In_165,In_101);
nor U1278 (N_1278,In_348,In_422);
or U1279 (N_1279,In_89,In_307);
nor U1280 (N_1280,In_287,In_984);
and U1281 (N_1281,In_681,In_0);
nand U1282 (N_1282,In_61,In_431);
or U1283 (N_1283,In_243,In_941);
nor U1284 (N_1284,In_952,In_450);
nand U1285 (N_1285,In_149,In_284);
nor U1286 (N_1286,In_486,In_436);
and U1287 (N_1287,In_304,In_402);
nand U1288 (N_1288,In_5,In_134);
and U1289 (N_1289,In_51,In_783);
or U1290 (N_1290,In_886,In_270);
or U1291 (N_1291,In_929,In_631);
nand U1292 (N_1292,In_306,In_631);
and U1293 (N_1293,In_110,In_449);
nor U1294 (N_1294,In_585,In_6);
nor U1295 (N_1295,In_494,In_287);
nor U1296 (N_1296,In_385,In_22);
and U1297 (N_1297,In_461,In_797);
nor U1298 (N_1298,In_672,In_61);
nor U1299 (N_1299,In_562,In_387);
or U1300 (N_1300,In_462,In_960);
nand U1301 (N_1301,In_305,In_407);
and U1302 (N_1302,In_988,In_200);
nand U1303 (N_1303,In_593,In_230);
and U1304 (N_1304,In_177,In_778);
nand U1305 (N_1305,In_771,In_783);
nand U1306 (N_1306,In_357,In_546);
nor U1307 (N_1307,In_422,In_216);
nand U1308 (N_1308,In_942,In_886);
nand U1309 (N_1309,In_45,In_14);
nor U1310 (N_1310,In_310,In_948);
nand U1311 (N_1311,In_192,In_792);
and U1312 (N_1312,In_408,In_37);
nand U1313 (N_1313,In_68,In_745);
nor U1314 (N_1314,In_41,In_421);
or U1315 (N_1315,In_209,In_52);
or U1316 (N_1316,In_558,In_383);
or U1317 (N_1317,In_609,In_162);
or U1318 (N_1318,In_622,In_74);
and U1319 (N_1319,In_979,In_338);
nand U1320 (N_1320,In_963,In_636);
and U1321 (N_1321,In_655,In_455);
nor U1322 (N_1322,In_710,In_863);
nor U1323 (N_1323,In_685,In_800);
nand U1324 (N_1324,In_414,In_385);
nand U1325 (N_1325,In_896,In_478);
nand U1326 (N_1326,In_216,In_979);
nor U1327 (N_1327,In_130,In_510);
xor U1328 (N_1328,In_590,In_918);
nor U1329 (N_1329,In_895,In_665);
nand U1330 (N_1330,In_578,In_150);
nor U1331 (N_1331,In_432,In_99);
nand U1332 (N_1332,In_242,In_675);
and U1333 (N_1333,In_359,In_383);
nor U1334 (N_1334,In_2,In_211);
nor U1335 (N_1335,In_53,In_902);
and U1336 (N_1336,In_871,In_41);
nor U1337 (N_1337,In_351,In_777);
nand U1338 (N_1338,In_800,In_918);
nor U1339 (N_1339,In_759,In_516);
and U1340 (N_1340,In_356,In_177);
or U1341 (N_1341,In_975,In_734);
or U1342 (N_1342,In_811,In_919);
or U1343 (N_1343,In_968,In_439);
nand U1344 (N_1344,In_94,In_272);
or U1345 (N_1345,In_226,In_354);
nor U1346 (N_1346,In_949,In_914);
nand U1347 (N_1347,In_225,In_584);
and U1348 (N_1348,In_79,In_550);
nor U1349 (N_1349,In_499,In_723);
nor U1350 (N_1350,In_393,In_85);
or U1351 (N_1351,In_726,In_713);
and U1352 (N_1352,In_352,In_249);
or U1353 (N_1353,In_827,In_449);
nor U1354 (N_1354,In_171,In_803);
nor U1355 (N_1355,In_361,In_592);
or U1356 (N_1356,In_538,In_235);
or U1357 (N_1357,In_235,In_899);
and U1358 (N_1358,In_418,In_585);
and U1359 (N_1359,In_484,In_165);
nand U1360 (N_1360,In_943,In_650);
and U1361 (N_1361,In_63,In_673);
nand U1362 (N_1362,In_931,In_980);
or U1363 (N_1363,In_209,In_856);
or U1364 (N_1364,In_679,In_897);
nor U1365 (N_1365,In_319,In_198);
and U1366 (N_1366,In_889,In_749);
nor U1367 (N_1367,In_159,In_316);
and U1368 (N_1368,In_315,In_1);
nand U1369 (N_1369,In_513,In_941);
nand U1370 (N_1370,In_765,In_651);
and U1371 (N_1371,In_150,In_36);
nand U1372 (N_1372,In_404,In_474);
nor U1373 (N_1373,In_143,In_556);
nand U1374 (N_1374,In_129,In_340);
nand U1375 (N_1375,In_995,In_521);
or U1376 (N_1376,In_777,In_463);
nand U1377 (N_1377,In_660,In_642);
or U1378 (N_1378,In_989,In_749);
and U1379 (N_1379,In_800,In_412);
nand U1380 (N_1380,In_270,In_892);
nand U1381 (N_1381,In_996,In_367);
nand U1382 (N_1382,In_965,In_703);
or U1383 (N_1383,In_558,In_538);
nor U1384 (N_1384,In_130,In_180);
and U1385 (N_1385,In_321,In_589);
and U1386 (N_1386,In_290,In_105);
nand U1387 (N_1387,In_51,In_282);
nor U1388 (N_1388,In_354,In_616);
and U1389 (N_1389,In_821,In_568);
and U1390 (N_1390,In_587,In_252);
nor U1391 (N_1391,In_707,In_354);
or U1392 (N_1392,In_501,In_390);
nand U1393 (N_1393,In_198,In_211);
or U1394 (N_1394,In_262,In_495);
or U1395 (N_1395,In_314,In_73);
and U1396 (N_1396,In_105,In_405);
and U1397 (N_1397,In_693,In_60);
xor U1398 (N_1398,In_417,In_743);
nor U1399 (N_1399,In_117,In_760);
nor U1400 (N_1400,In_382,In_256);
nand U1401 (N_1401,In_130,In_192);
nor U1402 (N_1402,In_246,In_900);
and U1403 (N_1403,In_204,In_910);
nor U1404 (N_1404,In_777,In_3);
nor U1405 (N_1405,In_796,In_758);
or U1406 (N_1406,In_264,In_457);
or U1407 (N_1407,In_55,In_542);
nand U1408 (N_1408,In_135,In_367);
and U1409 (N_1409,In_556,In_271);
or U1410 (N_1410,In_737,In_566);
nor U1411 (N_1411,In_598,In_662);
nand U1412 (N_1412,In_79,In_739);
or U1413 (N_1413,In_980,In_662);
nand U1414 (N_1414,In_239,In_930);
and U1415 (N_1415,In_464,In_493);
nand U1416 (N_1416,In_247,In_740);
nor U1417 (N_1417,In_978,In_760);
nor U1418 (N_1418,In_475,In_128);
nand U1419 (N_1419,In_738,In_804);
nor U1420 (N_1420,In_639,In_377);
nand U1421 (N_1421,In_273,In_203);
nand U1422 (N_1422,In_286,In_677);
nor U1423 (N_1423,In_110,In_314);
and U1424 (N_1424,In_715,In_884);
or U1425 (N_1425,In_327,In_544);
and U1426 (N_1426,In_387,In_627);
or U1427 (N_1427,In_78,In_211);
nand U1428 (N_1428,In_230,In_423);
nor U1429 (N_1429,In_231,In_505);
and U1430 (N_1430,In_796,In_946);
nand U1431 (N_1431,In_543,In_814);
and U1432 (N_1432,In_68,In_894);
nor U1433 (N_1433,In_699,In_131);
or U1434 (N_1434,In_5,In_404);
or U1435 (N_1435,In_506,In_892);
or U1436 (N_1436,In_565,In_419);
and U1437 (N_1437,In_681,In_982);
nor U1438 (N_1438,In_634,In_257);
and U1439 (N_1439,In_57,In_895);
or U1440 (N_1440,In_921,In_442);
and U1441 (N_1441,In_388,In_307);
nand U1442 (N_1442,In_315,In_528);
or U1443 (N_1443,In_234,In_64);
nand U1444 (N_1444,In_840,In_341);
and U1445 (N_1445,In_208,In_439);
nand U1446 (N_1446,In_836,In_783);
and U1447 (N_1447,In_792,In_716);
or U1448 (N_1448,In_420,In_683);
nand U1449 (N_1449,In_299,In_764);
nand U1450 (N_1450,In_972,In_180);
and U1451 (N_1451,In_80,In_325);
and U1452 (N_1452,In_569,In_790);
nand U1453 (N_1453,In_0,In_106);
nor U1454 (N_1454,In_663,In_18);
nor U1455 (N_1455,In_527,In_97);
xnor U1456 (N_1456,In_994,In_639);
and U1457 (N_1457,In_88,In_740);
and U1458 (N_1458,In_937,In_406);
nor U1459 (N_1459,In_252,In_755);
xnor U1460 (N_1460,In_800,In_508);
nor U1461 (N_1461,In_765,In_141);
or U1462 (N_1462,In_875,In_227);
nand U1463 (N_1463,In_616,In_17);
and U1464 (N_1464,In_67,In_47);
nor U1465 (N_1465,In_720,In_416);
nand U1466 (N_1466,In_576,In_372);
nand U1467 (N_1467,In_973,In_478);
nor U1468 (N_1468,In_255,In_791);
nand U1469 (N_1469,In_630,In_276);
nand U1470 (N_1470,In_824,In_494);
or U1471 (N_1471,In_825,In_618);
nor U1472 (N_1472,In_435,In_613);
nand U1473 (N_1473,In_257,In_699);
and U1474 (N_1474,In_685,In_376);
nand U1475 (N_1475,In_164,In_834);
nor U1476 (N_1476,In_600,In_894);
or U1477 (N_1477,In_798,In_615);
and U1478 (N_1478,In_457,In_996);
nand U1479 (N_1479,In_441,In_88);
or U1480 (N_1480,In_766,In_916);
or U1481 (N_1481,In_139,In_74);
and U1482 (N_1482,In_710,In_39);
or U1483 (N_1483,In_562,In_713);
or U1484 (N_1484,In_245,In_931);
nor U1485 (N_1485,In_704,In_958);
nor U1486 (N_1486,In_173,In_971);
nor U1487 (N_1487,In_864,In_256);
and U1488 (N_1488,In_804,In_308);
nor U1489 (N_1489,In_613,In_400);
nor U1490 (N_1490,In_202,In_188);
nor U1491 (N_1491,In_840,In_35);
or U1492 (N_1492,In_982,In_380);
and U1493 (N_1493,In_143,In_798);
xor U1494 (N_1494,In_979,In_255);
nand U1495 (N_1495,In_769,In_231);
nand U1496 (N_1496,In_576,In_660);
and U1497 (N_1497,In_113,In_79);
nand U1498 (N_1498,In_155,In_130);
or U1499 (N_1499,In_382,In_915);
nor U1500 (N_1500,In_259,In_966);
and U1501 (N_1501,In_197,In_396);
nand U1502 (N_1502,In_829,In_645);
and U1503 (N_1503,In_555,In_142);
or U1504 (N_1504,In_189,In_651);
and U1505 (N_1505,In_453,In_679);
nand U1506 (N_1506,In_11,In_406);
nor U1507 (N_1507,In_299,In_384);
and U1508 (N_1508,In_330,In_378);
nor U1509 (N_1509,In_380,In_372);
or U1510 (N_1510,In_641,In_484);
nand U1511 (N_1511,In_729,In_998);
nor U1512 (N_1512,In_286,In_532);
or U1513 (N_1513,In_510,In_251);
nand U1514 (N_1514,In_452,In_9);
or U1515 (N_1515,In_910,In_703);
or U1516 (N_1516,In_442,In_825);
and U1517 (N_1517,In_439,In_262);
or U1518 (N_1518,In_891,In_599);
nand U1519 (N_1519,In_591,In_204);
and U1520 (N_1520,In_100,In_235);
nand U1521 (N_1521,In_525,In_776);
or U1522 (N_1522,In_140,In_679);
or U1523 (N_1523,In_452,In_975);
and U1524 (N_1524,In_459,In_457);
nor U1525 (N_1525,In_520,In_855);
nand U1526 (N_1526,In_889,In_415);
nor U1527 (N_1527,In_398,In_303);
nand U1528 (N_1528,In_844,In_264);
nor U1529 (N_1529,In_23,In_299);
nand U1530 (N_1530,In_567,In_135);
and U1531 (N_1531,In_54,In_177);
or U1532 (N_1532,In_74,In_450);
nor U1533 (N_1533,In_251,In_305);
and U1534 (N_1534,In_351,In_345);
or U1535 (N_1535,In_817,In_473);
nor U1536 (N_1536,In_423,In_407);
or U1537 (N_1537,In_219,In_330);
and U1538 (N_1538,In_650,In_58);
and U1539 (N_1539,In_662,In_505);
nand U1540 (N_1540,In_818,In_33);
or U1541 (N_1541,In_117,In_537);
nor U1542 (N_1542,In_529,In_940);
and U1543 (N_1543,In_684,In_535);
and U1544 (N_1544,In_483,In_251);
and U1545 (N_1545,In_909,In_600);
nand U1546 (N_1546,In_724,In_459);
and U1547 (N_1547,In_79,In_671);
and U1548 (N_1548,In_191,In_140);
or U1549 (N_1549,In_773,In_844);
nor U1550 (N_1550,In_290,In_935);
nand U1551 (N_1551,In_335,In_987);
or U1552 (N_1552,In_145,In_660);
and U1553 (N_1553,In_7,In_452);
nor U1554 (N_1554,In_930,In_658);
nor U1555 (N_1555,In_548,In_241);
and U1556 (N_1556,In_603,In_669);
and U1557 (N_1557,In_683,In_56);
nand U1558 (N_1558,In_25,In_410);
nor U1559 (N_1559,In_288,In_386);
or U1560 (N_1560,In_326,In_942);
and U1561 (N_1561,In_109,In_850);
nand U1562 (N_1562,In_646,In_855);
nand U1563 (N_1563,In_357,In_901);
or U1564 (N_1564,In_760,In_233);
and U1565 (N_1565,In_389,In_650);
and U1566 (N_1566,In_712,In_366);
nor U1567 (N_1567,In_891,In_784);
nor U1568 (N_1568,In_529,In_562);
nor U1569 (N_1569,In_233,In_593);
nor U1570 (N_1570,In_763,In_722);
nor U1571 (N_1571,In_781,In_132);
nand U1572 (N_1572,In_622,In_817);
or U1573 (N_1573,In_52,In_672);
nor U1574 (N_1574,In_212,In_542);
or U1575 (N_1575,In_391,In_778);
or U1576 (N_1576,In_839,In_440);
nand U1577 (N_1577,In_545,In_373);
nand U1578 (N_1578,In_858,In_77);
or U1579 (N_1579,In_30,In_822);
nand U1580 (N_1580,In_79,In_554);
or U1581 (N_1581,In_677,In_52);
nand U1582 (N_1582,In_463,In_277);
and U1583 (N_1583,In_43,In_259);
nand U1584 (N_1584,In_290,In_668);
nand U1585 (N_1585,In_97,In_388);
nor U1586 (N_1586,In_58,In_110);
xnor U1587 (N_1587,In_392,In_340);
nor U1588 (N_1588,In_41,In_211);
nor U1589 (N_1589,In_156,In_110);
nor U1590 (N_1590,In_435,In_524);
nand U1591 (N_1591,In_857,In_254);
nand U1592 (N_1592,In_916,In_826);
and U1593 (N_1593,In_372,In_528);
nor U1594 (N_1594,In_465,In_83);
and U1595 (N_1595,In_324,In_290);
or U1596 (N_1596,In_573,In_746);
or U1597 (N_1597,In_192,In_835);
nor U1598 (N_1598,In_316,In_214);
nor U1599 (N_1599,In_91,In_961);
or U1600 (N_1600,In_713,In_138);
and U1601 (N_1601,In_592,In_617);
and U1602 (N_1602,In_285,In_73);
nand U1603 (N_1603,In_803,In_825);
nand U1604 (N_1604,In_386,In_812);
and U1605 (N_1605,In_650,In_474);
nor U1606 (N_1606,In_343,In_127);
nand U1607 (N_1607,In_250,In_199);
or U1608 (N_1608,In_238,In_3);
nor U1609 (N_1609,In_498,In_762);
nand U1610 (N_1610,In_358,In_583);
and U1611 (N_1611,In_559,In_819);
and U1612 (N_1612,In_30,In_853);
nand U1613 (N_1613,In_93,In_395);
nor U1614 (N_1614,In_815,In_974);
nor U1615 (N_1615,In_331,In_416);
nor U1616 (N_1616,In_50,In_427);
nor U1617 (N_1617,In_587,In_900);
and U1618 (N_1618,In_434,In_96);
and U1619 (N_1619,In_551,In_556);
or U1620 (N_1620,In_655,In_466);
or U1621 (N_1621,In_50,In_291);
nand U1622 (N_1622,In_375,In_588);
or U1623 (N_1623,In_222,In_403);
nor U1624 (N_1624,In_229,In_546);
and U1625 (N_1625,In_959,In_531);
nor U1626 (N_1626,In_309,In_944);
or U1627 (N_1627,In_544,In_970);
and U1628 (N_1628,In_340,In_824);
nand U1629 (N_1629,In_738,In_529);
nor U1630 (N_1630,In_231,In_722);
or U1631 (N_1631,In_159,In_908);
or U1632 (N_1632,In_299,In_751);
nor U1633 (N_1633,In_132,In_492);
and U1634 (N_1634,In_417,In_678);
and U1635 (N_1635,In_35,In_662);
and U1636 (N_1636,In_30,In_395);
nand U1637 (N_1637,In_590,In_426);
nor U1638 (N_1638,In_966,In_770);
and U1639 (N_1639,In_275,In_627);
nand U1640 (N_1640,In_432,In_178);
or U1641 (N_1641,In_460,In_374);
nand U1642 (N_1642,In_574,In_774);
and U1643 (N_1643,In_904,In_947);
nor U1644 (N_1644,In_417,In_654);
or U1645 (N_1645,In_169,In_485);
nand U1646 (N_1646,In_446,In_785);
and U1647 (N_1647,In_55,In_559);
and U1648 (N_1648,In_648,In_496);
nor U1649 (N_1649,In_108,In_795);
nor U1650 (N_1650,In_958,In_966);
nand U1651 (N_1651,In_501,In_806);
or U1652 (N_1652,In_664,In_571);
and U1653 (N_1653,In_545,In_81);
nor U1654 (N_1654,In_989,In_760);
and U1655 (N_1655,In_495,In_338);
nor U1656 (N_1656,In_24,In_554);
nor U1657 (N_1657,In_597,In_91);
and U1658 (N_1658,In_511,In_493);
and U1659 (N_1659,In_462,In_51);
or U1660 (N_1660,In_148,In_127);
nand U1661 (N_1661,In_707,In_640);
nor U1662 (N_1662,In_264,In_589);
or U1663 (N_1663,In_530,In_150);
nor U1664 (N_1664,In_815,In_683);
or U1665 (N_1665,In_695,In_741);
nor U1666 (N_1666,In_322,In_753);
nand U1667 (N_1667,In_952,In_515);
nand U1668 (N_1668,In_616,In_357);
nand U1669 (N_1669,In_863,In_264);
nand U1670 (N_1670,In_773,In_680);
nor U1671 (N_1671,In_478,In_634);
and U1672 (N_1672,In_505,In_716);
or U1673 (N_1673,In_641,In_115);
nand U1674 (N_1674,In_787,In_100);
nand U1675 (N_1675,In_926,In_35);
or U1676 (N_1676,In_963,In_982);
and U1677 (N_1677,In_989,In_940);
or U1678 (N_1678,In_949,In_872);
nor U1679 (N_1679,In_378,In_512);
nand U1680 (N_1680,In_644,In_156);
or U1681 (N_1681,In_263,In_76);
and U1682 (N_1682,In_42,In_570);
nor U1683 (N_1683,In_314,In_421);
and U1684 (N_1684,In_741,In_682);
and U1685 (N_1685,In_193,In_529);
nand U1686 (N_1686,In_478,In_152);
and U1687 (N_1687,In_594,In_562);
nor U1688 (N_1688,In_707,In_819);
nor U1689 (N_1689,In_739,In_558);
nor U1690 (N_1690,In_840,In_276);
or U1691 (N_1691,In_258,In_676);
nor U1692 (N_1692,In_26,In_481);
nand U1693 (N_1693,In_454,In_27);
nor U1694 (N_1694,In_661,In_155);
or U1695 (N_1695,In_3,In_652);
and U1696 (N_1696,In_602,In_213);
and U1697 (N_1697,In_707,In_955);
or U1698 (N_1698,In_348,In_990);
nor U1699 (N_1699,In_971,In_449);
and U1700 (N_1700,In_870,In_627);
or U1701 (N_1701,In_452,In_936);
nand U1702 (N_1702,In_278,In_682);
and U1703 (N_1703,In_333,In_663);
nor U1704 (N_1704,In_547,In_267);
or U1705 (N_1705,In_238,In_0);
nand U1706 (N_1706,In_65,In_198);
or U1707 (N_1707,In_820,In_333);
nand U1708 (N_1708,In_727,In_975);
nand U1709 (N_1709,In_207,In_376);
nand U1710 (N_1710,In_533,In_237);
nand U1711 (N_1711,In_165,In_377);
nor U1712 (N_1712,In_76,In_706);
nor U1713 (N_1713,In_10,In_456);
nand U1714 (N_1714,In_214,In_551);
nor U1715 (N_1715,In_36,In_34);
and U1716 (N_1716,In_188,In_242);
nand U1717 (N_1717,In_701,In_195);
and U1718 (N_1718,In_807,In_860);
or U1719 (N_1719,In_956,In_810);
or U1720 (N_1720,In_149,In_105);
and U1721 (N_1721,In_62,In_23);
or U1722 (N_1722,In_425,In_886);
nor U1723 (N_1723,In_233,In_323);
or U1724 (N_1724,In_225,In_730);
or U1725 (N_1725,In_398,In_726);
nor U1726 (N_1726,In_161,In_209);
or U1727 (N_1727,In_518,In_664);
and U1728 (N_1728,In_617,In_78);
xor U1729 (N_1729,In_345,In_115);
xor U1730 (N_1730,In_804,In_270);
nand U1731 (N_1731,In_620,In_397);
or U1732 (N_1732,In_457,In_898);
or U1733 (N_1733,In_593,In_278);
and U1734 (N_1734,In_215,In_593);
nand U1735 (N_1735,In_405,In_219);
nor U1736 (N_1736,In_385,In_517);
nand U1737 (N_1737,In_710,In_615);
nand U1738 (N_1738,In_215,In_272);
nor U1739 (N_1739,In_617,In_589);
nand U1740 (N_1740,In_837,In_45);
nor U1741 (N_1741,In_282,In_412);
nor U1742 (N_1742,In_604,In_770);
nand U1743 (N_1743,In_192,In_134);
and U1744 (N_1744,In_387,In_889);
and U1745 (N_1745,In_35,In_560);
nand U1746 (N_1746,In_850,In_249);
nor U1747 (N_1747,In_31,In_105);
nor U1748 (N_1748,In_517,In_318);
and U1749 (N_1749,In_337,In_457);
or U1750 (N_1750,In_284,In_204);
and U1751 (N_1751,In_614,In_576);
or U1752 (N_1752,In_632,In_810);
nand U1753 (N_1753,In_371,In_239);
nand U1754 (N_1754,In_779,In_98);
nand U1755 (N_1755,In_813,In_714);
or U1756 (N_1756,In_310,In_865);
and U1757 (N_1757,In_843,In_570);
nand U1758 (N_1758,In_738,In_339);
nand U1759 (N_1759,In_35,In_156);
xnor U1760 (N_1760,In_69,In_637);
or U1761 (N_1761,In_548,In_635);
or U1762 (N_1762,In_790,In_955);
or U1763 (N_1763,In_641,In_26);
and U1764 (N_1764,In_998,In_73);
xnor U1765 (N_1765,In_107,In_447);
nand U1766 (N_1766,In_342,In_267);
or U1767 (N_1767,In_879,In_509);
nand U1768 (N_1768,In_30,In_607);
nand U1769 (N_1769,In_554,In_514);
and U1770 (N_1770,In_286,In_495);
and U1771 (N_1771,In_721,In_989);
nor U1772 (N_1772,In_68,In_886);
or U1773 (N_1773,In_872,In_809);
and U1774 (N_1774,In_31,In_590);
nor U1775 (N_1775,In_595,In_746);
nand U1776 (N_1776,In_169,In_118);
nor U1777 (N_1777,In_307,In_720);
and U1778 (N_1778,In_459,In_971);
or U1779 (N_1779,In_531,In_309);
and U1780 (N_1780,In_581,In_530);
nor U1781 (N_1781,In_374,In_443);
and U1782 (N_1782,In_292,In_465);
or U1783 (N_1783,In_742,In_78);
or U1784 (N_1784,In_440,In_424);
nor U1785 (N_1785,In_738,In_492);
nand U1786 (N_1786,In_907,In_286);
nand U1787 (N_1787,In_126,In_809);
nand U1788 (N_1788,In_72,In_479);
nor U1789 (N_1789,In_148,In_851);
or U1790 (N_1790,In_622,In_896);
and U1791 (N_1791,In_367,In_443);
and U1792 (N_1792,In_575,In_23);
or U1793 (N_1793,In_279,In_481);
or U1794 (N_1794,In_108,In_894);
and U1795 (N_1795,In_773,In_208);
and U1796 (N_1796,In_256,In_913);
and U1797 (N_1797,In_914,In_283);
or U1798 (N_1798,In_219,In_970);
nor U1799 (N_1799,In_403,In_671);
and U1800 (N_1800,In_488,In_215);
nor U1801 (N_1801,In_892,In_166);
and U1802 (N_1802,In_504,In_959);
or U1803 (N_1803,In_894,In_651);
nor U1804 (N_1804,In_614,In_366);
nand U1805 (N_1805,In_797,In_874);
nor U1806 (N_1806,In_953,In_420);
and U1807 (N_1807,In_408,In_401);
nor U1808 (N_1808,In_90,In_205);
nand U1809 (N_1809,In_71,In_674);
nor U1810 (N_1810,In_733,In_726);
nand U1811 (N_1811,In_945,In_357);
nand U1812 (N_1812,In_97,In_198);
and U1813 (N_1813,In_522,In_22);
nand U1814 (N_1814,In_609,In_915);
and U1815 (N_1815,In_416,In_184);
or U1816 (N_1816,In_703,In_766);
nand U1817 (N_1817,In_633,In_896);
or U1818 (N_1818,In_482,In_575);
nor U1819 (N_1819,In_348,In_807);
nor U1820 (N_1820,In_481,In_550);
nand U1821 (N_1821,In_396,In_273);
nor U1822 (N_1822,In_542,In_489);
or U1823 (N_1823,In_197,In_273);
and U1824 (N_1824,In_960,In_221);
nor U1825 (N_1825,In_956,In_722);
or U1826 (N_1826,In_852,In_69);
nor U1827 (N_1827,In_767,In_634);
and U1828 (N_1828,In_765,In_107);
and U1829 (N_1829,In_554,In_92);
nor U1830 (N_1830,In_772,In_382);
and U1831 (N_1831,In_733,In_399);
or U1832 (N_1832,In_878,In_862);
or U1833 (N_1833,In_508,In_206);
nand U1834 (N_1834,In_214,In_442);
and U1835 (N_1835,In_215,In_792);
nor U1836 (N_1836,In_327,In_38);
or U1837 (N_1837,In_97,In_371);
nor U1838 (N_1838,In_549,In_331);
or U1839 (N_1839,In_638,In_399);
nand U1840 (N_1840,In_903,In_725);
nand U1841 (N_1841,In_545,In_26);
nor U1842 (N_1842,In_202,In_186);
and U1843 (N_1843,In_104,In_832);
nor U1844 (N_1844,In_932,In_413);
nor U1845 (N_1845,In_537,In_953);
and U1846 (N_1846,In_349,In_97);
or U1847 (N_1847,In_33,In_105);
and U1848 (N_1848,In_216,In_734);
nand U1849 (N_1849,In_810,In_708);
nand U1850 (N_1850,In_64,In_90);
or U1851 (N_1851,In_354,In_408);
nand U1852 (N_1852,In_227,In_975);
and U1853 (N_1853,In_643,In_641);
and U1854 (N_1854,In_371,In_619);
nand U1855 (N_1855,In_295,In_555);
and U1856 (N_1856,In_152,In_335);
and U1857 (N_1857,In_838,In_75);
nand U1858 (N_1858,In_156,In_333);
nand U1859 (N_1859,In_795,In_412);
or U1860 (N_1860,In_163,In_347);
nand U1861 (N_1861,In_752,In_992);
or U1862 (N_1862,In_207,In_276);
or U1863 (N_1863,In_352,In_407);
nand U1864 (N_1864,In_998,In_326);
nor U1865 (N_1865,In_166,In_320);
nand U1866 (N_1866,In_452,In_177);
nor U1867 (N_1867,In_142,In_502);
nand U1868 (N_1868,In_464,In_958);
nand U1869 (N_1869,In_377,In_114);
or U1870 (N_1870,In_189,In_431);
nor U1871 (N_1871,In_425,In_952);
and U1872 (N_1872,In_252,In_448);
or U1873 (N_1873,In_417,In_383);
and U1874 (N_1874,In_204,In_507);
nor U1875 (N_1875,In_49,In_285);
and U1876 (N_1876,In_330,In_295);
and U1877 (N_1877,In_494,In_532);
nand U1878 (N_1878,In_839,In_96);
nand U1879 (N_1879,In_306,In_732);
or U1880 (N_1880,In_418,In_298);
and U1881 (N_1881,In_419,In_633);
or U1882 (N_1882,In_345,In_610);
or U1883 (N_1883,In_279,In_792);
and U1884 (N_1884,In_506,In_667);
and U1885 (N_1885,In_363,In_825);
nand U1886 (N_1886,In_122,In_406);
and U1887 (N_1887,In_513,In_833);
nand U1888 (N_1888,In_659,In_302);
nand U1889 (N_1889,In_534,In_463);
nor U1890 (N_1890,In_239,In_76);
or U1891 (N_1891,In_766,In_547);
nor U1892 (N_1892,In_656,In_91);
nand U1893 (N_1893,In_811,In_494);
and U1894 (N_1894,In_698,In_454);
and U1895 (N_1895,In_112,In_884);
or U1896 (N_1896,In_24,In_103);
or U1897 (N_1897,In_606,In_3);
and U1898 (N_1898,In_491,In_138);
and U1899 (N_1899,In_961,In_574);
nand U1900 (N_1900,In_355,In_921);
nand U1901 (N_1901,In_867,In_721);
or U1902 (N_1902,In_247,In_989);
and U1903 (N_1903,In_938,In_300);
nor U1904 (N_1904,In_505,In_265);
or U1905 (N_1905,In_233,In_600);
or U1906 (N_1906,In_253,In_185);
nand U1907 (N_1907,In_944,In_374);
xnor U1908 (N_1908,In_787,In_435);
and U1909 (N_1909,In_948,In_568);
xor U1910 (N_1910,In_148,In_117);
and U1911 (N_1911,In_208,In_58);
nand U1912 (N_1912,In_998,In_823);
and U1913 (N_1913,In_223,In_746);
and U1914 (N_1914,In_986,In_299);
nand U1915 (N_1915,In_363,In_219);
nand U1916 (N_1916,In_225,In_762);
or U1917 (N_1917,In_652,In_173);
nand U1918 (N_1918,In_461,In_38);
and U1919 (N_1919,In_139,In_349);
and U1920 (N_1920,In_611,In_202);
nand U1921 (N_1921,In_428,In_841);
and U1922 (N_1922,In_602,In_23);
and U1923 (N_1923,In_63,In_925);
nor U1924 (N_1924,In_31,In_420);
nand U1925 (N_1925,In_72,In_289);
nand U1926 (N_1926,In_499,In_351);
nor U1927 (N_1927,In_254,In_452);
or U1928 (N_1928,In_971,In_705);
or U1929 (N_1929,In_356,In_946);
and U1930 (N_1930,In_212,In_387);
and U1931 (N_1931,In_150,In_900);
nand U1932 (N_1932,In_673,In_679);
or U1933 (N_1933,In_162,In_471);
nand U1934 (N_1934,In_129,In_650);
nand U1935 (N_1935,In_481,In_980);
or U1936 (N_1936,In_659,In_202);
nand U1937 (N_1937,In_415,In_541);
and U1938 (N_1938,In_370,In_13);
nor U1939 (N_1939,In_289,In_102);
or U1940 (N_1940,In_785,In_651);
nor U1941 (N_1941,In_362,In_441);
nor U1942 (N_1942,In_383,In_20);
or U1943 (N_1943,In_466,In_700);
nor U1944 (N_1944,In_759,In_434);
and U1945 (N_1945,In_400,In_937);
xnor U1946 (N_1946,In_695,In_598);
nand U1947 (N_1947,In_469,In_613);
nand U1948 (N_1948,In_436,In_990);
and U1949 (N_1949,In_189,In_960);
and U1950 (N_1950,In_79,In_540);
or U1951 (N_1951,In_590,In_21);
nor U1952 (N_1952,In_280,In_343);
and U1953 (N_1953,In_920,In_636);
or U1954 (N_1954,In_200,In_748);
nand U1955 (N_1955,In_270,In_264);
xor U1956 (N_1956,In_787,In_381);
nor U1957 (N_1957,In_963,In_212);
and U1958 (N_1958,In_61,In_870);
or U1959 (N_1959,In_205,In_776);
and U1960 (N_1960,In_261,In_915);
and U1961 (N_1961,In_3,In_478);
or U1962 (N_1962,In_391,In_179);
or U1963 (N_1963,In_901,In_542);
and U1964 (N_1964,In_460,In_499);
and U1965 (N_1965,In_714,In_984);
or U1966 (N_1966,In_160,In_215);
and U1967 (N_1967,In_267,In_94);
or U1968 (N_1968,In_787,In_20);
and U1969 (N_1969,In_309,In_562);
or U1970 (N_1970,In_440,In_168);
nor U1971 (N_1971,In_453,In_380);
or U1972 (N_1972,In_25,In_728);
nor U1973 (N_1973,In_574,In_889);
nor U1974 (N_1974,In_185,In_718);
xor U1975 (N_1975,In_702,In_418);
or U1976 (N_1976,In_583,In_45);
nor U1977 (N_1977,In_572,In_876);
nor U1978 (N_1978,In_964,In_950);
or U1979 (N_1979,In_374,In_91);
and U1980 (N_1980,In_974,In_908);
or U1981 (N_1981,In_812,In_704);
or U1982 (N_1982,In_550,In_154);
nand U1983 (N_1983,In_848,In_457);
nand U1984 (N_1984,In_95,In_497);
nor U1985 (N_1985,In_141,In_95);
nand U1986 (N_1986,In_899,In_729);
and U1987 (N_1987,In_729,In_336);
nand U1988 (N_1988,In_146,In_736);
nand U1989 (N_1989,In_660,In_11);
nor U1990 (N_1990,In_950,In_834);
nor U1991 (N_1991,In_319,In_43);
nor U1992 (N_1992,In_422,In_226);
nor U1993 (N_1993,In_288,In_83);
and U1994 (N_1994,In_99,In_463);
or U1995 (N_1995,In_509,In_193);
nand U1996 (N_1996,In_167,In_683);
nand U1997 (N_1997,In_525,In_173);
nor U1998 (N_1998,In_734,In_527);
or U1999 (N_1999,In_893,In_714);
and U2000 (N_2000,N_1789,N_45);
nor U2001 (N_2001,N_1281,N_403);
nand U2002 (N_2002,N_878,N_542);
nand U2003 (N_2003,N_31,N_11);
nand U2004 (N_2004,N_1106,N_1068);
and U2005 (N_2005,N_381,N_423);
and U2006 (N_2006,N_226,N_605);
nor U2007 (N_2007,N_1684,N_813);
and U2008 (N_2008,N_360,N_39);
or U2009 (N_2009,N_201,N_74);
or U2010 (N_2010,N_728,N_1774);
and U2011 (N_2011,N_438,N_629);
or U2012 (N_2012,N_1412,N_1022);
nor U2013 (N_2013,N_1333,N_168);
nor U2014 (N_2014,N_1012,N_1960);
or U2015 (N_2015,N_1053,N_1058);
and U2016 (N_2016,N_1201,N_348);
and U2017 (N_2017,N_1753,N_1628);
nand U2018 (N_2018,N_318,N_746);
and U2019 (N_2019,N_1839,N_1922);
or U2020 (N_2020,N_169,N_1406);
nor U2021 (N_2021,N_800,N_328);
nor U2022 (N_2022,N_1108,N_1315);
nand U2023 (N_2023,N_1984,N_1651);
nand U2024 (N_2024,N_339,N_1205);
and U2025 (N_2025,N_1302,N_1078);
nand U2026 (N_2026,N_286,N_1366);
and U2027 (N_2027,N_1314,N_1511);
nand U2028 (N_2028,N_1507,N_1580);
or U2029 (N_2029,N_1608,N_87);
nor U2030 (N_2030,N_937,N_128);
nor U2031 (N_2031,N_698,N_171);
nand U2032 (N_2032,N_1141,N_1597);
and U2033 (N_2033,N_1599,N_1893);
or U2034 (N_2034,N_1750,N_1988);
nor U2035 (N_2035,N_81,N_1242);
nor U2036 (N_2036,N_1697,N_998);
nor U2037 (N_2037,N_13,N_1279);
nand U2038 (N_2038,N_176,N_1531);
and U2039 (N_2039,N_1060,N_1342);
and U2040 (N_2040,N_1257,N_1883);
and U2041 (N_2041,N_492,N_1876);
and U2042 (N_2042,N_1429,N_1648);
nand U2043 (N_2043,N_662,N_118);
nand U2044 (N_2044,N_270,N_1128);
and U2045 (N_2045,N_1027,N_1488);
and U2046 (N_2046,N_915,N_1170);
nand U2047 (N_2047,N_557,N_1555);
nor U2048 (N_2048,N_60,N_1017);
nand U2049 (N_2049,N_56,N_988);
or U2050 (N_2050,N_1030,N_723);
or U2051 (N_2051,N_1588,N_1325);
or U2052 (N_2052,N_603,N_479);
and U2053 (N_2053,N_1211,N_1400);
xnor U2054 (N_2054,N_209,N_734);
and U2055 (N_2055,N_1755,N_535);
or U2056 (N_2056,N_566,N_591);
or U2057 (N_2057,N_643,N_616);
or U2058 (N_2058,N_92,N_1891);
and U2059 (N_2059,N_1538,N_1807);
xor U2060 (N_2060,N_1417,N_185);
and U2061 (N_2061,N_1031,N_1163);
nor U2062 (N_2062,N_1390,N_1035);
nor U2063 (N_2063,N_71,N_249);
nand U2064 (N_2064,N_753,N_1716);
nand U2065 (N_2065,N_1259,N_214);
nand U2066 (N_2066,N_1808,N_1143);
nand U2067 (N_2067,N_1380,N_613);
nor U2068 (N_2068,N_1700,N_795);
or U2069 (N_2069,N_906,N_920);
nor U2070 (N_2070,N_511,N_1975);
and U2071 (N_2071,N_383,N_1646);
nand U2072 (N_2072,N_1356,N_556);
or U2073 (N_2073,N_1742,N_1419);
nor U2074 (N_2074,N_294,N_1041);
nand U2075 (N_2075,N_1777,N_330);
nor U2076 (N_2076,N_830,N_1731);
or U2077 (N_2077,N_9,N_792);
and U2078 (N_2078,N_1806,N_1393);
nand U2079 (N_2079,N_869,N_1675);
nand U2080 (N_2080,N_415,N_1452);
nor U2081 (N_2081,N_458,N_1404);
nand U2082 (N_2082,N_1265,N_430);
nor U2083 (N_2083,N_1887,N_400);
and U2084 (N_2084,N_1728,N_1207);
nor U2085 (N_2085,N_1440,N_720);
xnor U2086 (N_2086,N_326,N_633);
or U2087 (N_2087,N_1190,N_773);
or U2088 (N_2088,N_1647,N_628);
or U2089 (N_2089,N_929,N_136);
nand U2090 (N_2090,N_206,N_861);
or U2091 (N_2091,N_1252,N_963);
and U2092 (N_2092,N_1187,N_1218);
and U2093 (N_2093,N_1316,N_1309);
nor U2094 (N_2094,N_1306,N_1153);
xnor U2095 (N_2095,N_623,N_1310);
or U2096 (N_2096,N_1104,N_562);
nor U2097 (N_2097,N_585,N_778);
nand U2098 (N_2098,N_1475,N_303);
or U2099 (N_2099,N_1363,N_1465);
and U2100 (N_2100,N_1087,N_1308);
xnor U2101 (N_2101,N_677,N_35);
or U2102 (N_2102,N_1947,N_1147);
and U2103 (N_2103,N_112,N_1896);
nor U2104 (N_2104,N_429,N_212);
nor U2105 (N_2105,N_1998,N_109);
nor U2106 (N_2106,N_1392,N_1900);
or U2107 (N_2107,N_626,N_1243);
nand U2108 (N_2108,N_150,N_42);
nand U2109 (N_2109,N_1819,N_460);
nor U2110 (N_2110,N_1083,N_283);
or U2111 (N_2111,N_1817,N_964);
or U2112 (N_2112,N_1919,N_829);
and U2113 (N_2113,N_1957,N_1722);
and U2114 (N_2114,N_395,N_984);
and U2115 (N_2115,N_1358,N_1156);
or U2116 (N_2116,N_1081,N_1842);
nor U2117 (N_2117,N_621,N_1369);
and U2118 (N_2118,N_587,N_772);
nand U2119 (N_2119,N_292,N_1816);
and U2120 (N_2120,N_1550,N_1881);
nor U2121 (N_2121,N_908,N_27);
or U2122 (N_2122,N_1296,N_1101);
and U2123 (N_2123,N_1735,N_1815);
and U2124 (N_2124,N_102,N_363);
nand U2125 (N_2125,N_853,N_922);
and U2126 (N_2126,N_198,N_1091);
nor U2127 (N_2127,N_611,N_285);
nand U2128 (N_2128,N_533,N_174);
nor U2129 (N_2129,N_748,N_1561);
or U2130 (N_2130,N_1189,N_192);
nor U2131 (N_2131,N_1095,N_1791);
nand U2132 (N_2132,N_268,N_1952);
and U2133 (N_2133,N_565,N_1518);
nor U2134 (N_2134,N_186,N_692);
or U2135 (N_2135,N_468,N_49);
nand U2136 (N_2136,N_1051,N_439);
nand U2137 (N_2137,N_1523,N_1300);
nor U2138 (N_2138,N_1196,N_1470);
nand U2139 (N_2139,N_1332,N_287);
or U2140 (N_2140,N_1226,N_582);
nand U2141 (N_2141,N_491,N_1371);
and U2142 (N_2142,N_965,N_1779);
nand U2143 (N_2143,N_1831,N_1076);
nor U2144 (N_2144,N_450,N_505);
and U2145 (N_2145,N_1782,N_1403);
nand U2146 (N_2146,N_1540,N_1373);
nand U2147 (N_2147,N_1705,N_131);
nor U2148 (N_2148,N_227,N_173);
nor U2149 (N_2149,N_1563,N_986);
nor U2150 (N_2150,N_968,N_817);
or U2151 (N_2151,N_14,N_1948);
and U2152 (N_2152,N_1469,N_612);
nand U2153 (N_2153,N_1803,N_251);
and U2154 (N_2154,N_1418,N_705);
nand U2155 (N_2155,N_596,N_104);
nand U2156 (N_2156,N_989,N_321);
and U2157 (N_2157,N_1630,N_253);
or U2158 (N_2158,N_1943,N_604);
nor U2159 (N_2159,N_534,N_1422);
nor U2160 (N_2160,N_1554,N_1216);
and U2161 (N_2161,N_1394,N_1622);
nand U2162 (N_2162,N_1365,N_64);
or U2163 (N_2163,N_1926,N_1640);
nand U2164 (N_2164,N_1913,N_580);
and U2165 (N_2165,N_1672,N_1024);
or U2166 (N_2166,N_1154,N_806);
nor U2167 (N_2167,N_432,N_702);
or U2168 (N_2168,N_632,N_546);
nor U2169 (N_2169,N_1991,N_180);
or U2170 (N_2170,N_1945,N_729);
and U2171 (N_2171,N_759,N_5);
nor U2172 (N_2172,N_271,N_838);
nand U2173 (N_2173,N_1951,N_1486);
nor U2174 (N_2174,N_870,N_1754);
and U2175 (N_2175,N_1157,N_1214);
nor U2176 (N_2176,N_379,N_1834);
nand U2177 (N_2177,N_1547,N_1125);
or U2178 (N_2178,N_1906,N_1005);
and U2179 (N_2179,N_222,N_12);
nor U2180 (N_2180,N_1769,N_1276);
or U2181 (N_2181,N_356,N_519);
or U2182 (N_2182,N_0,N_467);
nor U2183 (N_2183,N_1927,N_548);
nor U2184 (N_2184,N_133,N_687);
or U2185 (N_2185,N_19,N_143);
or U2186 (N_2186,N_1911,N_962);
and U2187 (N_2187,N_899,N_1349);
nor U2188 (N_2188,N_1225,N_1983);
nor U2189 (N_2189,N_1822,N_857);
or U2190 (N_2190,N_375,N_1097);
or U2191 (N_2191,N_428,N_1982);
nand U2192 (N_2192,N_398,N_1649);
and U2193 (N_2193,N_1908,N_865);
and U2194 (N_2194,N_1884,N_1286);
or U2195 (N_2195,N_1758,N_799);
and U2196 (N_2196,N_950,N_106);
nor U2197 (N_2197,N_418,N_655);
or U2198 (N_2198,N_296,N_1541);
or U2199 (N_2199,N_1474,N_1334);
or U2200 (N_2200,N_127,N_1075);
or U2201 (N_2201,N_371,N_1036);
or U2202 (N_2202,N_1503,N_1338);
or U2203 (N_2203,N_1650,N_495);
and U2204 (N_2204,N_854,N_1639);
nand U2205 (N_2205,N_1450,N_724);
nor U2206 (N_2206,N_1551,N_1160);
and U2207 (N_2207,N_62,N_1423);
nand U2208 (N_2208,N_16,N_125);
nand U2209 (N_2209,N_1532,N_1443);
nor U2210 (N_2210,N_1268,N_1577);
or U2211 (N_2211,N_502,N_581);
and U2212 (N_2212,N_1484,N_1631);
and U2213 (N_2213,N_298,N_170);
or U2214 (N_2214,N_1074,N_847);
or U2215 (N_2215,N_137,N_1433);
xor U2216 (N_2216,N_1458,N_1456);
or U2217 (N_2217,N_455,N_1910);
nor U2218 (N_2218,N_837,N_284);
nand U2219 (N_2219,N_1290,N_1341);
nand U2220 (N_2220,N_1120,N_153);
nand U2221 (N_2221,N_665,N_1050);
or U2222 (N_2222,N_1621,N_1335);
nand U2223 (N_2223,N_664,N_392);
nand U2224 (N_2224,N_615,N_1064);
and U2225 (N_2225,N_480,N_1402);
and U2226 (N_2226,N_1123,N_789);
and U2227 (N_2227,N_866,N_788);
and U2228 (N_2228,N_441,N_1837);
and U2229 (N_2229,N_116,N_1864);
nor U2230 (N_2230,N_1641,N_203);
nor U2231 (N_2231,N_1627,N_1212);
or U2232 (N_2232,N_1294,N_179);
nor U2233 (N_2233,N_1105,N_952);
and U2234 (N_2234,N_1553,N_333);
nor U2235 (N_2235,N_297,N_175);
and U2236 (N_2236,N_641,N_992);
nand U2237 (N_2237,N_618,N_1655);
nand U2238 (N_2238,N_999,N_259);
nand U2239 (N_2239,N_1263,N_1133);
nand U2240 (N_2240,N_888,N_1144);
nand U2241 (N_2241,N_835,N_1751);
or U2242 (N_2242,N_916,N_1925);
nand U2243 (N_2243,N_17,N_549);
nor U2244 (N_2244,N_931,N_316);
nand U2245 (N_2245,N_500,N_1330);
nand U2246 (N_2246,N_1854,N_1770);
or U2247 (N_2247,N_1931,N_1015);
nor U2248 (N_2248,N_684,N_1937);
nor U2249 (N_2249,N_1367,N_782);
nor U2250 (N_2250,N_1915,N_1969);
and U2251 (N_2251,N_1388,N_1185);
and U2252 (N_2252,N_466,N_1763);
or U2253 (N_2253,N_1601,N_364);
and U2254 (N_2254,N_384,N_1016);
and U2255 (N_2255,N_1084,N_1796);
and U2256 (N_2256,N_1351,N_1583);
nor U2257 (N_2257,N_1549,N_661);
nor U2258 (N_2258,N_1132,N_1914);
nand U2259 (N_2259,N_1353,N_204);
nand U2260 (N_2260,N_402,N_1326);
nand U2261 (N_2261,N_528,N_636);
xnor U2262 (N_2262,N_1570,N_541);
or U2263 (N_2263,N_974,N_293);
nand U2264 (N_2264,N_544,N_38);
nand U2265 (N_2265,N_1814,N_673);
and U2266 (N_2266,N_1451,N_193);
and U2267 (N_2267,N_58,N_719);
and U2268 (N_2268,N_1061,N_927);
or U2269 (N_2269,N_84,N_889);
nor U2270 (N_2270,N_68,N_1544);
nand U2271 (N_2271,N_928,N_163);
nand U2272 (N_2272,N_833,N_1637);
nand U2273 (N_2273,N_1985,N_602);
and U2274 (N_2274,N_1527,N_1029);
and U2275 (N_2275,N_1855,N_158);
or U2276 (N_2276,N_783,N_1530);
nor U2277 (N_2277,N_306,N_561);
nand U2278 (N_2278,N_1956,N_211);
and U2279 (N_2279,N_678,N_564);
nor U2280 (N_2280,N_417,N_786);
nor U2281 (N_2281,N_738,N_697);
and U2282 (N_2282,N_1245,N_1677);
nand U2283 (N_2283,N_1692,N_766);
or U2284 (N_2284,N_1683,N_1589);
or U2285 (N_2285,N_91,N_448);
and U2286 (N_2286,N_1841,N_787);
and U2287 (N_2287,N_836,N_820);
nand U2288 (N_2288,N_1206,N_237);
or U2289 (N_2289,N_224,N_1929);
and U2290 (N_2290,N_1849,N_1065);
nor U2291 (N_2291,N_779,N_26);
nand U2292 (N_2292,N_290,N_461);
nand U2293 (N_2293,N_508,N_159);
or U2294 (N_2294,N_944,N_1227);
nor U2295 (N_2295,N_691,N_1699);
and U2296 (N_2296,N_1591,N_197);
or U2297 (N_2297,N_905,N_101);
nor U2298 (N_2298,N_1711,N_440);
and U2299 (N_2299,N_957,N_1992);
nand U2300 (N_2300,N_1460,N_1886);
or U2301 (N_2301,N_1278,N_396);
or U2302 (N_2302,N_1890,N_246);
or U2303 (N_2303,N_1823,N_443);
xor U2304 (N_2304,N_1961,N_1493);
nor U2305 (N_2305,N_1395,N_1034);
and U2306 (N_2306,N_907,N_1139);
or U2307 (N_2307,N_1044,N_529);
nand U2308 (N_2308,N_1192,N_785);
or U2309 (N_2309,N_183,N_105);
or U2310 (N_2310,N_1520,N_1501);
xor U2311 (N_2311,N_1569,N_1739);
and U2312 (N_2312,N_353,N_1892);
nor U2313 (N_2313,N_1566,N_311);
nor U2314 (N_2314,N_1668,N_1416);
or U2315 (N_2315,N_1071,N_243);
nand U2316 (N_2316,N_97,N_1603);
nor U2317 (N_2317,N_1466,N_841);
nor U2318 (N_2318,N_953,N_649);
nor U2319 (N_2319,N_1197,N_737);
and U2320 (N_2320,N_1669,N_498);
nor U2321 (N_2321,N_313,N_1571);
nor U2322 (N_2322,N_1611,N_1783);
nor U2323 (N_2323,N_1399,N_1000);
and U2324 (N_2324,N_1923,N_1730);
or U2325 (N_2325,N_345,N_1293);
and U2326 (N_2326,N_1134,N_901);
nor U2327 (N_2327,N_1378,N_302);
nor U2328 (N_2328,N_1933,N_412);
or U2329 (N_2329,N_1489,N_512);
nor U2330 (N_2330,N_996,N_754);
or U2331 (N_2331,N_1069,N_1155);
nand U2332 (N_2332,N_877,N_257);
nor U2333 (N_2333,N_1496,N_1347);
or U2334 (N_2334,N_1159,N_1498);
or U2335 (N_2335,N_1271,N_1250);
or U2336 (N_2336,N_149,N_474);
nand U2337 (N_2337,N_1826,N_653);
and U2338 (N_2338,N_1678,N_1584);
and U2339 (N_2339,N_1836,N_555);
xnor U2340 (N_2340,N_213,N_1409);
or U2341 (N_2341,N_427,N_1100);
nor U2342 (N_2342,N_1209,N_409);
nor U2343 (N_2343,N_1327,N_1632);
nand U2344 (N_2344,N_1478,N_413);
nand U2345 (N_2345,N_1413,N_1901);
nand U2346 (N_2346,N_744,N_951);
and U2347 (N_2347,N_497,N_1537);
and U2348 (N_2348,N_791,N_609);
and U2349 (N_2349,N_242,N_1512);
nor U2350 (N_2350,N_588,N_863);
nor U2351 (N_2351,N_368,N_681);
and U2352 (N_2352,N_682,N_1319);
nand U2353 (N_2353,N_516,N_1624);
nor U2354 (N_2354,N_1936,N_851);
nor U2355 (N_2355,N_1479,N_732);
nor U2356 (N_2356,N_282,N_571);
and U2357 (N_2357,N_524,N_642);
nand U2358 (N_2358,N_995,N_1536);
nand U2359 (N_2359,N_1810,N_775);
and U2360 (N_2360,N_501,N_1447);
nor U2361 (N_2361,N_1989,N_597);
nand U2362 (N_2362,N_390,N_736);
or U2363 (N_2363,N_485,N_1918);
or U2364 (N_2364,N_1695,N_1467);
or U2365 (N_2365,N_827,N_80);
nor U2366 (N_2366,N_416,N_453);
nor U2367 (N_2367,N_1348,N_651);
or U2368 (N_2368,N_1248,N_1485);
and U2369 (N_2369,N_86,N_1008);
or U2370 (N_2370,N_1636,N_247);
nand U2371 (N_2371,N_666,N_1436);
nand U2372 (N_2372,N_1321,N_1618);
and U2373 (N_2373,N_327,N_1519);
nand U2374 (N_2374,N_199,N_66);
or U2375 (N_2375,N_1165,N_776);
or U2376 (N_2376,N_1964,N_140);
nor U2377 (N_2377,N_599,N_1558);
nor U2378 (N_2378,N_966,N_1747);
and U2379 (N_2379,N_221,N_1950);
nand U2380 (N_2380,N_1202,N_164);
and U2381 (N_2381,N_1152,N_1217);
nor U2382 (N_2382,N_2,N_1829);
nand U2383 (N_2383,N_157,N_1021);
nor U2384 (N_2384,N_489,N_796);
and U2385 (N_2385,N_1492,N_1346);
xnor U2386 (N_2386,N_1938,N_1067);
nor U2387 (N_2387,N_1904,N_939);
nand U2388 (N_2388,N_231,N_1360);
nand U2389 (N_2389,N_579,N_15);
nand U2390 (N_2390,N_601,N_469);
and U2391 (N_2391,N_1800,N_538);
nor U2392 (N_2392,N_1194,N_55);
nor U2393 (N_2393,N_1203,N_1233);
nor U2394 (N_2394,N_1173,N_210);
or U2395 (N_2395,N_1515,N_446);
and U2396 (N_2396,N_525,N_1255);
and U2397 (N_2397,N_295,N_1019);
or U2398 (N_2398,N_1247,N_289);
and U2399 (N_2399,N_1934,N_1652);
and U2400 (N_2400,N_73,N_454);
nor U2401 (N_2401,N_1568,N_471);
and U2402 (N_2402,N_144,N_864);
nand U2403 (N_2403,N_1978,N_933);
nor U2404 (N_2404,N_1759,N_1052);
nand U2405 (N_2405,N_1917,N_1744);
nor U2406 (N_2406,N_1131,N_167);
nand U2407 (N_2407,N_223,N_1781);
or U2408 (N_2408,N_1838,N_1273);
or U2409 (N_2409,N_510,N_627);
and U2410 (N_2410,N_1798,N_1113);
nor U2411 (N_2411,N_804,N_425);
nor U2412 (N_2412,N_1521,N_1843);
nor U2413 (N_2413,N_1797,N_419);
and U2414 (N_2414,N_818,N_32);
nand U2415 (N_2415,N_794,N_261);
or U2416 (N_2416,N_83,N_1606);
and U2417 (N_2417,N_1653,N_954);
and U2418 (N_2418,N_380,N_188);
and U2419 (N_2419,N_156,N_648);
nand U2420 (N_2420,N_1320,N_452);
or U2421 (N_2421,N_1262,N_1946);
nand U2422 (N_2422,N_756,N_1355);
or U2423 (N_2423,N_693,N_1665);
nand U2424 (N_2424,N_1230,N_1736);
and U2425 (N_2425,N_1572,N_1118);
nand U2426 (N_2426,N_1374,N_914);
or U2427 (N_2427,N_595,N_1193);
and U2428 (N_2428,N_1556,N_22);
and U2429 (N_2429,N_1965,N_631);
or U2430 (N_2430,N_85,N_1701);
nand U2431 (N_2431,N_570,N_926);
nand U2432 (N_2432,N_1088,N_1720);
nor U2433 (N_2433,N_743,N_1459);
and U2434 (N_2434,N_1623,N_695);
or U2435 (N_2435,N_1018,N_1787);
or U2436 (N_2436,N_522,N_1146);
nand U2437 (N_2437,N_1949,N_1240);
or U2438 (N_2438,N_1862,N_671);
or U2439 (N_2439,N_1654,N_713);
nand U2440 (N_2440,N_437,N_1851);
nand U2441 (N_2441,N_1004,N_146);
and U2442 (N_2442,N_372,N_1283);
and U2443 (N_2443,N_1013,N_1275);
nor U2444 (N_2444,N_955,N_36);
or U2445 (N_2445,N_336,N_278);
or U2446 (N_2446,N_7,N_28);
nor U2447 (N_2447,N_1704,N_1344);
or U2448 (N_2448,N_184,N_378);
nor U2449 (N_2449,N_1574,N_828);
or U2450 (N_2450,N_96,N_1103);
nor U2451 (N_2451,N_1733,N_859);
nand U2452 (N_2452,N_917,N_904);
nand U2453 (N_2453,N_1732,N_1629);
or U2454 (N_2454,N_1298,N_521);
nand U2455 (N_2455,N_803,N_393);
or U2456 (N_2456,N_919,N_1702);
nand U2457 (N_2457,N_1685,N_1329);
nand U2458 (N_2458,N_658,N_1014);
and U2459 (N_2459,N_1375,N_1506);
nor U2460 (N_2460,N_1661,N_54);
or U2461 (N_2461,N_1726,N_1136);
nand U2462 (N_2462,N_1644,N_886);
and U2463 (N_2463,N_1368,N_1059);
and U2464 (N_2464,N_879,N_431);
or U2465 (N_2465,N_774,N_987);
or U2466 (N_2466,N_1181,N_1533);
nor U2467 (N_2467,N_559,N_1534);
and U2468 (N_2468,N_1743,N_921);
and U2469 (N_2469,N_1545,N_281);
and U2470 (N_2470,N_1072,N_1020);
nand U2471 (N_2471,N_645,N_802);
and U2472 (N_2472,N_1438,N_1172);
or U2473 (N_2473,N_1727,N_1437);
nand U2474 (N_2474,N_232,N_319);
and U2475 (N_2475,N_1425,N_82);
or U2476 (N_2476,N_476,N_1408);
and U2477 (N_2477,N_52,N_1856);
nor U2478 (N_2478,N_1057,N_1713);
nor U2479 (N_2479,N_332,N_758);
or U2480 (N_2480,N_1508,N_1039);
or U2481 (N_2481,N_255,N_536);
or U2482 (N_2482,N_1266,N_1182);
and U2483 (N_2483,N_1424,N_1613);
nand U2484 (N_2484,N_76,N_166);
xnor U2485 (N_2485,N_1526,N_250);
xnor U2486 (N_2486,N_1888,N_690);
or U2487 (N_2487,N_1176,N_1038);
nor U2488 (N_2488,N_1494,N_1959);
nand U2489 (N_2489,N_236,N_749);
and U2490 (N_2490,N_1323,N_1878);
and U2491 (N_2491,N_590,N_1706);
nand U2492 (N_2492,N_735,N_189);
and U2493 (N_2493,N_1169,N_1213);
and U2494 (N_2494,N_1756,N_1110);
nor U2495 (N_2495,N_811,N_1757);
and U2496 (N_2496,N_463,N_1096);
nor U2497 (N_2497,N_477,N_47);
nor U2498 (N_2498,N_1663,N_1619);
nand U2499 (N_2499,N_1431,N_93);
and U2500 (N_2500,N_483,N_1142);
or U2501 (N_2501,N_1215,N_1037);
nor U2502 (N_2502,N_1303,N_1301);
nor U2503 (N_2503,N_1517,N_1411);
nand U2504 (N_2504,N_1307,N_1481);
nor U2505 (N_2505,N_1620,N_320);
nand U2506 (N_2506,N_718,N_537);
and U2507 (N_2507,N_205,N_424);
and U2508 (N_2508,N_1381,N_1175);
nand U2509 (N_2509,N_1604,N_624);
nand U2510 (N_2510,N_620,N_196);
nor U2511 (N_2511,N_470,N_1174);
and U2512 (N_2512,N_1625,N_1578);
and U2513 (N_2513,N_161,N_993);
or U2514 (N_2514,N_385,N_961);
nand U2515 (N_2515,N_110,N_586);
nor U2516 (N_2516,N_387,N_540);
nor U2517 (N_2517,N_312,N_801);
nand U2518 (N_2518,N_1339,N_1126);
and U2519 (N_2519,N_714,N_1434);
nand U2520 (N_2520,N_761,N_852);
nand U2521 (N_2521,N_1869,N_975);
nand U2522 (N_2522,N_858,N_433);
and U2523 (N_2523,N_1898,N_239);
nor U2524 (N_2524,N_350,N_1528);
nor U2525 (N_2525,N_1396,N_1682);
nand U2526 (N_2526,N_194,N_1239);
and U2527 (N_2527,N_1738,N_1428);
nand U2528 (N_2528,N_1760,N_493);
xor U2529 (N_2529,N_1430,N_1043);
nor U2530 (N_2530,N_1382,N_674);
nor U2531 (N_2531,N_299,N_1092);
or U2532 (N_2532,N_1612,N_1107);
and U2533 (N_2533,N_948,N_969);
or U2534 (N_2534,N_1567,N_637);
and U2535 (N_2535,N_280,N_78);
nand U2536 (N_2536,N_569,N_1195);
and U2537 (N_2537,N_1444,N_1102);
nand U2538 (N_2538,N_575,N_750);
or U2539 (N_2539,N_1026,N_1510);
or U2540 (N_2540,N_217,N_366);
and U2541 (N_2541,N_457,N_1935);
nand U2542 (N_2542,N_960,N_1564);
nor U2543 (N_2543,N_1762,N_1859);
and U2544 (N_2544,N_1383,N_1483);
and U2545 (N_2545,N_1670,N_1993);
nand U2546 (N_2546,N_1524,N_1228);
and U2547 (N_2547,N_1966,N_347);
nand U2548 (N_2548,N_1799,N_607);
and U2549 (N_2549,N_819,N_1282);
or U2550 (N_2550,N_238,N_1151);
nor U2551 (N_2551,N_475,N_890);
or U2552 (N_2552,N_1609,N_435);
nand U2553 (N_2553,N_1994,N_1865);
or U2554 (N_2554,N_1680,N_1274);
nand U2555 (N_2555,N_530,N_343);
nand U2556 (N_2556,N_1331,N_1179);
or U2557 (N_2557,N_370,N_531);
and U2558 (N_2558,N_1099,N_499);
or U2559 (N_2559,N_181,N_1063);
or U2560 (N_2560,N_404,N_1903);
or U2561 (N_2561,N_1224,N_1860);
and U2562 (N_2562,N_1009,N_1171);
nand U2563 (N_2563,N_1291,N_1539);
or U2564 (N_2564,N_129,N_1658);
nor U2565 (N_2565,N_100,N_43);
and U2566 (N_2566,N_814,N_980);
nor U2567 (N_2567,N_589,N_1184);
and U2568 (N_2568,N_970,N_24);
xnor U2569 (N_2569,N_739,N_335);
nor U2570 (N_2570,N_1186,N_1696);
nand U2571 (N_2571,N_77,N_1385);
nand U2572 (N_2572,N_593,N_1721);
and U2573 (N_2573,N_504,N_1924);
nand U2574 (N_2574,N_924,N_598);
and U2575 (N_2575,N_672,N_1772);
or U2576 (N_2576,N_1812,N_1766);
nor U2577 (N_2577,N_997,N_288);
nor U2578 (N_2578,N_709,N_860);
nor U2579 (N_2579,N_509,N_138);
or U2580 (N_2580,N_1850,N_1028);
or U2581 (N_2581,N_177,N_765);
nor U2582 (N_2582,N_1804,N_1288);
and U2583 (N_2583,N_1222,N_1150);
and U2584 (N_2584,N_490,N_1734);
and U2585 (N_2585,N_1077,N_1477);
and U2586 (N_2586,N_563,N_1045);
nand U2587 (N_2587,N_1280,N_816);
or U2588 (N_2588,N_600,N_1006);
nand U2589 (N_2589,N_1761,N_912);
or U2590 (N_2590,N_1482,N_1776);
nor U2591 (N_2591,N_369,N_1698);
nand U2592 (N_2592,N_1880,N_1897);
and U2593 (N_2593,N_1236,N_777);
and U2594 (N_2594,N_1905,N_887);
xor U2595 (N_2595,N_862,N_63);
and U2596 (N_2596,N_1707,N_61);
and U2597 (N_2597,N_1500,N_981);
nor U2598 (N_2598,N_1548,N_1600);
and U2599 (N_2599,N_1594,N_619);
and U2600 (N_2600,N_898,N_871);
or U2601 (N_2601,N_338,N_1180);
or U2602 (N_2602,N_160,N_1198);
nor U2603 (N_2603,N_1188,N_1710);
or U2604 (N_2604,N_59,N_694);
nor U2605 (N_2605,N_848,N_376);
nor U2606 (N_2606,N_1912,N_930);
or U2607 (N_2607,N_1802,N_34);
nor U2608 (N_2608,N_307,N_503);
nand U2609 (N_2609,N_208,N_844);
or U2610 (N_2610,N_1260,N_1562);
or U2611 (N_2611,N_1112,N_1970);
nand U2612 (N_2612,N_1049,N_1514);
nor U2613 (N_2613,N_108,N_721);
or U2614 (N_2614,N_868,N_1879);
or U2615 (N_2615,N_639,N_1962);
nand U2616 (N_2616,N_1830,N_805);
nor U2617 (N_2617,N_1846,N_708);
nor U2618 (N_2618,N_1305,N_770);
nor U2619 (N_2619,N_1939,N_824);
nand U2620 (N_2620,N_883,N_1073);
and U2621 (N_2621,N_578,N_355);
nor U2622 (N_2622,N_977,N_1313);
and U2623 (N_2623,N_1656,N_545);
or U2624 (N_2624,N_1853,N_148);
and U2625 (N_2625,N_1312,N_526);
nand U2626 (N_2626,N_374,N_660);
nor U2627 (N_2627,N_365,N_315);
nand U2628 (N_2628,N_763,N_527);
or U2629 (N_2629,N_506,N_594);
nor U2630 (N_2630,N_1835,N_554);
nor U2631 (N_2631,N_1,N_659);
nor U2632 (N_2632,N_696,N_855);
nand U2633 (N_2633,N_932,N_715);
nand U2634 (N_2634,N_434,N_940);
nand U2635 (N_2635,N_1177,N_1161);
nor U2636 (N_2636,N_88,N_1085);
and U2637 (N_2637,N_1135,N_1867);
nor U2638 (N_2638,N_1979,N_1449);
or U2639 (N_2639,N_1328,N_1119);
or U2640 (N_2640,N_346,N_342);
nand U2641 (N_2641,N_876,N_1256);
xnor U2642 (N_2642,N_822,N_1138);
or U2643 (N_2643,N_1741,N_892);
nor U2644 (N_2644,N_1253,N_1219);
nor U2645 (N_2645,N_334,N_1254);
nand U2646 (N_2646,N_680,N_1748);
nor U2647 (N_2647,N_1267,N_414);
and U2648 (N_2648,N_277,N_391);
nand U2649 (N_2649,N_885,N_683);
nor U2650 (N_2650,N_147,N_1241);
or U2651 (N_2651,N_3,N_991);
and U2652 (N_2652,N_230,N_1746);
or U2653 (N_2653,N_507,N_567);
or U2654 (N_2654,N_1920,N_98);
nand U2655 (N_2655,N_1350,N_162);
and U2656 (N_2656,N_711,N_1414);
nor U2657 (N_2657,N_134,N_1208);
or U2658 (N_2658,N_1055,N_831);
and U2659 (N_2659,N_676,N_1398);
and U2660 (N_2660,N_382,N_971);
or U2661 (N_2661,N_103,N_1048);
nor U2662 (N_2662,N_1158,N_1638);
and U2663 (N_2663,N_1795,N_1780);
or U2664 (N_2664,N_1295,N_1805);
and U2665 (N_2665,N_1832,N_4);
or U2666 (N_2666,N_742,N_784);
nand U2667 (N_2667,N_275,N_1011);
nor U2668 (N_2668,N_1928,N_165);
nand U2669 (N_2669,N_229,N_1304);
nand U2670 (N_2670,N_154,N_654);
nor U2671 (N_2671,N_421,N_717);
nand U2672 (N_2672,N_207,N_1575);
nor U2673 (N_2673,N_1054,N_1809);
or U2674 (N_2674,N_1066,N_614);
and U2675 (N_2675,N_872,N_132);
or U2676 (N_2676,N_1535,N_1565);
or U2677 (N_2677,N_79,N_310);
or U2678 (N_2678,N_925,N_688);
nor U2679 (N_2679,N_331,N_1792);
nor U2680 (N_2680,N_1497,N_1667);
nand U2681 (N_2681,N_1542,N_1930);
and U2682 (N_2682,N_464,N_200);
and U2683 (N_2683,N_638,N_1405);
or U2684 (N_2684,N_494,N_1042);
and U2685 (N_2685,N_1464,N_1093);
nand U2686 (N_2686,N_1686,N_1079);
nor U2687 (N_2687,N_248,N_1117);
nor U2688 (N_2688,N_880,N_1902);
or U2689 (N_2689,N_1752,N_20);
and U2690 (N_2690,N_1786,N_1788);
nor U2691 (N_2691,N_608,N_967);
nand U2692 (N_2692,N_934,N_1237);
or U2693 (N_2693,N_976,N_979);
or U2694 (N_2694,N_913,N_834);
nand U2695 (N_2695,N_123,N_1062);
nand U2696 (N_2696,N_1820,N_405);
nand U2697 (N_2697,N_354,N_644);
and U2698 (N_2698,N_1137,N_1056);
nor U2699 (N_2699,N_1875,N_1703);
or U2700 (N_2700,N_647,N_263);
nand U2701 (N_2701,N_340,N_911);
or U2702 (N_2702,N_1086,N_1824);
nor U2703 (N_2703,N_1972,N_1605);
and U2704 (N_2704,N_1689,N_1657);
nand U2705 (N_2705,N_1445,N_1167);
nor U2706 (N_2706,N_1468,N_1094);
nand U2707 (N_2707,N_918,N_305);
or U2708 (N_2708,N_51,N_324);
nand U2709 (N_2709,N_1124,N_244);
nor U2710 (N_2710,N_1958,N_1415);
nor U2711 (N_2711,N_1676,N_1617);
nor U2712 (N_2712,N_946,N_436);
and U2713 (N_2713,N_1585,N_361);
or U2714 (N_2714,N_1121,N_1635);
or U2715 (N_2715,N_1397,N_94);
nor U2716 (N_2716,N_1420,N_1111);
nand U2717 (N_2717,N_1432,N_1040);
or U2718 (N_2718,N_72,N_1932);
or U2719 (N_2719,N_606,N_1340);
and U2720 (N_2720,N_426,N_1223);
or U2721 (N_2721,N_1980,N_228);
or U2722 (N_2722,N_1708,N_406);
and U2723 (N_2723,N_1848,N_517);
nand U2724 (N_2724,N_139,N_1318);
nand U2725 (N_2725,N_947,N_553);
or U2726 (N_2726,N_625,N_769);
nor U2727 (N_2727,N_1098,N_1688);
or U2728 (N_2728,N_269,N_573);
and U2729 (N_2729,N_240,N_513);
nor U2730 (N_2730,N_1709,N_1082);
nand U2731 (N_2731,N_1874,N_202);
and U2732 (N_2732,N_1940,N_1909);
nor U2733 (N_2733,N_826,N_1793);
nor U2734 (N_2734,N_1357,N_1235);
nor U2735 (N_2735,N_1372,N_1794);
or U2736 (N_2736,N_191,N_543);
nand U2737 (N_2737,N_456,N_685);
and U2738 (N_2738,N_135,N_107);
or U2739 (N_2739,N_710,N_1457);
nor U2740 (N_2740,N_634,N_771);
and U2741 (N_2741,N_121,N_1974);
or U2742 (N_2742,N_1127,N_1882);
nor U2743 (N_2743,N_1522,N_357);
and U2744 (N_2744,N_1899,N_1999);
nand U2745 (N_2745,N_1967,N_1873);
nand U2746 (N_2746,N_1987,N_576);
or U2747 (N_2747,N_1130,N_111);
or U2748 (N_2748,N_584,N_234);
nor U2749 (N_2749,N_1191,N_943);
nand U2750 (N_2750,N_1889,N_1343);
nand U2751 (N_2751,N_1513,N_1895);
or U2752 (N_2752,N_1299,N_514);
nor U2753 (N_2753,N_1954,N_839);
nor U2754 (N_2754,N_1246,N_1659);
xor U2755 (N_2755,N_1285,N_856);
and U2756 (N_2756,N_1324,N_1023);
and U2757 (N_2757,N_539,N_178);
nor U2758 (N_2758,N_793,N_329);
nand U2759 (N_2759,N_1953,N_6);
nor U2760 (N_2760,N_1345,N_1487);
nor U2761 (N_2761,N_126,N_1070);
and U2762 (N_2762,N_622,N_1626);
and U2763 (N_2763,N_235,N_1080);
nor U2764 (N_2764,N_1109,N_1579);
or U2765 (N_2765,N_1813,N_532);
nor U2766 (N_2766,N_323,N_399);
and U2767 (N_2767,N_1337,N_1200);
and U2768 (N_2768,N_956,N_1129);
and U2769 (N_2769,N_903,N_1505);
nand U2770 (N_2770,N_1364,N_1463);
nand U2771 (N_2771,N_1007,N_1712);
and U2772 (N_2772,N_1811,N_1354);
nand U2773 (N_2773,N_95,N_1003);
nor U2774 (N_2774,N_1955,N_881);
nor U2775 (N_2775,N_1386,N_1586);
nand U2776 (N_2776,N_1687,N_1261);
nand U2777 (N_2777,N_1990,N_577);
nand U2778 (N_2778,N_444,N_1765);
nor U2779 (N_2779,N_1941,N_1921);
nand U2780 (N_2780,N_1529,N_1166);
nor U2781 (N_2781,N_547,N_1775);
nand U2782 (N_2782,N_337,N_652);
nor U2783 (N_2783,N_151,N_1145);
nand U2784 (N_2784,N_1204,N_1871);
or U2785 (N_2785,N_1289,N_1968);
nor U2786 (N_2786,N_389,N_1352);
nor U2787 (N_2787,N_472,N_1502);
or U2788 (N_2788,N_115,N_910);
and U2789 (N_2789,N_449,N_1546);
nand U2790 (N_2790,N_520,N_1499);
and U2791 (N_2791,N_1840,N_1690);
nor U2792 (N_2792,N_117,N_701);
and U2793 (N_2793,N_1461,N_938);
nand U2794 (N_2794,N_1322,N_1047);
and U2795 (N_2795,N_1582,N_767);
or U2796 (N_2796,N_893,N_990);
nand U2797 (N_2797,N_65,N_635);
or U2798 (N_2798,N_760,N_195);
or U2799 (N_2799,N_1877,N_1472);
and U2800 (N_2800,N_1453,N_670);
or U2801 (N_2801,N_909,N_1614);
nand U2802 (N_2802,N_10,N_845);
nor U2803 (N_2803,N_959,N_1764);
nor U2804 (N_2804,N_982,N_1825);
or U2805 (N_2805,N_1148,N_496);
nand U2806 (N_2806,N_1495,N_1616);
nor U2807 (N_2807,N_875,N_465);
nand U2808 (N_2808,N_712,N_1595);
nand U2809 (N_2809,N_1238,N_57);
nand U2810 (N_2810,N_764,N_473);
or U2811 (N_2811,N_1377,N_1581);
or U2812 (N_2812,N_120,N_18);
or U2813 (N_2813,N_276,N_994);
nand U2814 (N_2814,N_1596,N_1391);
nor U2815 (N_2815,N_1963,N_1719);
nand U2816 (N_2816,N_1410,N_843);
nand U2817 (N_2817,N_1439,N_40);
nand U2818 (N_2818,N_44,N_1001);
or U2819 (N_2819,N_973,N_245);
or U2820 (N_2820,N_699,N_730);
nand U2821 (N_2821,N_727,N_215);
and U2822 (N_2822,N_942,N_668);
or U2823 (N_2823,N_484,N_640);
nand U2824 (N_2824,N_344,N_1401);
and U2825 (N_2825,N_1662,N_1297);
nand U2826 (N_2826,N_808,N_362);
or U2827 (N_2827,N_1446,N_842);
nor U2828 (N_2828,N_1916,N_1361);
nand U2829 (N_2829,N_1724,N_1183);
or U2830 (N_2830,N_1114,N_481);
or U2831 (N_2831,N_897,N_972);
and U2832 (N_2832,N_1694,N_1767);
and U2833 (N_2833,N_351,N_1642);
nand U2834 (N_2834,N_958,N_1480);
and U2835 (N_2835,N_442,N_30);
and U2836 (N_2836,N_1660,N_1389);
nand U2837 (N_2837,N_486,N_1971);
nand U2838 (N_2838,N_1162,N_985);
nor U2839 (N_2839,N_155,N_873);
nor U2840 (N_2840,N_704,N_141);
or U2841 (N_2841,N_523,N_89);
nand U2842 (N_2842,N_462,N_1633);
and U2843 (N_2843,N_124,N_1277);
or U2844 (N_2844,N_849,N_1116);
or U2845 (N_2845,N_1387,N_23);
or U2846 (N_2846,N_896,N_1973);
and U2847 (N_2847,N_304,N_716);
and U2848 (N_2848,N_1723,N_1768);
nand U2849 (N_2849,N_1229,N_790);
nor U2850 (N_2850,N_265,N_274);
and U2851 (N_2851,N_1643,N_1745);
or U2852 (N_2852,N_29,N_359);
nand U2853 (N_2853,N_190,N_488);
or U2854 (N_2854,N_325,N_1336);
or U2855 (N_2855,N_1210,N_407);
nand U2856 (N_2856,N_825,N_1234);
nand U2857 (N_2857,N_1863,N_583);
nor U2858 (N_2858,N_309,N_1525);
nor U2859 (N_2859,N_768,N_341);
and U2860 (N_2860,N_1442,N_1269);
or U2861 (N_2861,N_75,N_1010);
or U2862 (N_2862,N_1249,N_1857);
or U2863 (N_2863,N_1376,N_21);
and U2864 (N_2864,N_722,N_122);
nor U2865 (N_2865,N_1090,N_1679);
and U2866 (N_2866,N_731,N_1462);
nand U2867 (N_2867,N_1749,N_936);
nor U2868 (N_2868,N_552,N_1995);
and U2869 (N_2869,N_747,N_1718);
xor U2870 (N_2870,N_119,N_386);
nor U2871 (N_2871,N_408,N_264);
nand U2872 (N_2872,N_50,N_300);
or U2873 (N_2873,N_233,N_1244);
and U2874 (N_2874,N_1046,N_1421);
and U2875 (N_2875,N_1674,N_1634);
nor U2876 (N_2876,N_145,N_1251);
nor U2877 (N_2877,N_1491,N_923);
nand U2878 (N_2878,N_1996,N_1559);
nand U2879 (N_2879,N_1740,N_902);
nand U2880 (N_2880,N_218,N_610);
or U2881 (N_2881,N_273,N_1592);
and U2882 (N_2882,N_515,N_459);
and U2883 (N_2883,N_679,N_945);
nand U2884 (N_2884,N_978,N_1818);
and U2885 (N_2885,N_900,N_895);
and U2886 (N_2886,N_1359,N_99);
nor U2887 (N_2887,N_884,N_797);
or U2888 (N_2888,N_1866,N_422);
or U2889 (N_2889,N_1976,N_322);
and U2890 (N_2890,N_741,N_46);
and U2891 (N_2891,N_894,N_941);
nand U2892 (N_2892,N_451,N_241);
or U2893 (N_2893,N_518,N_812);
nand U2894 (N_2894,N_1448,N_733);
and U2895 (N_2895,N_1801,N_703);
and U2896 (N_2896,N_1778,N_301);
and U2897 (N_2897,N_551,N_267);
or U2898 (N_2898,N_1221,N_1140);
and U2899 (N_2899,N_706,N_707);
nand U2900 (N_2900,N_1370,N_367);
and U2901 (N_2901,N_675,N_689);
and U2902 (N_2902,N_1362,N_1593);
xnor U2903 (N_2903,N_8,N_1942);
nand U2904 (N_2904,N_1784,N_1435);
and U2905 (N_2905,N_48,N_1149);
nand U2906 (N_2906,N_1615,N_807);
and U2907 (N_2907,N_1122,N_1509);
or U2908 (N_2908,N_1693,N_751);
and U2909 (N_2909,N_41,N_1264);
nor U2910 (N_2910,N_810,N_254);
nand U2911 (N_2911,N_1426,N_1645);
nand U2912 (N_2912,N_1476,N_755);
nor U2913 (N_2913,N_172,N_1833);
or U2914 (N_2914,N_114,N_752);
or U2915 (N_2915,N_1790,N_219);
nor U2916 (N_2916,N_1894,N_1771);
xnor U2917 (N_2917,N_397,N_823);
or U2918 (N_2918,N_1560,N_252);
nor U2919 (N_2919,N_867,N_37);
and U2920 (N_2920,N_815,N_1164);
and U2921 (N_2921,N_142,N_663);
and U2922 (N_2922,N_130,N_1168);
or U2923 (N_2923,N_850,N_1986);
nand U2924 (N_2924,N_686,N_1607);
nand U2925 (N_2925,N_1427,N_67);
or U2926 (N_2926,N_272,N_1317);
or U2927 (N_2927,N_1178,N_182);
and U2928 (N_2928,N_1666,N_447);
or U2929 (N_2929,N_317,N_657);
or U2930 (N_2930,N_256,N_667);
or U2931 (N_2931,N_949,N_1610);
or U2932 (N_2932,N_487,N_1199);
nor U2933 (N_2933,N_1032,N_821);
or U2934 (N_2934,N_617,N_1828);
or U2935 (N_2935,N_1270,N_314);
nor U2936 (N_2936,N_669,N_291);
and U2937 (N_2937,N_592,N_725);
and U2938 (N_2938,N_1576,N_1997);
nor U2939 (N_2939,N_1907,N_420);
and U2940 (N_2940,N_25,N_840);
and U2941 (N_2941,N_1858,N_1590);
nand U2942 (N_2942,N_832,N_745);
and U2943 (N_2943,N_891,N_1587);
or U2944 (N_2944,N_1981,N_780);
or U2945 (N_2945,N_1002,N_33);
or U2946 (N_2946,N_70,N_700);
or U2947 (N_2947,N_1292,N_574);
nor U2948 (N_2948,N_1455,N_411);
nor U2949 (N_2949,N_740,N_1311);
nand U2950 (N_2950,N_1231,N_630);
nor U2951 (N_2951,N_558,N_220);
nand U2952 (N_2952,N_1573,N_1454);
or U2953 (N_2953,N_1773,N_1598);
and U2954 (N_2954,N_262,N_568);
nand U2955 (N_2955,N_1785,N_1407);
xor U2956 (N_2956,N_1870,N_1272);
nand U2957 (N_2957,N_798,N_1033);
and U2958 (N_2958,N_1490,N_410);
nand U2959 (N_2959,N_377,N_358);
nand U2960 (N_2960,N_394,N_1557);
and U2961 (N_2961,N_1552,N_1232);
and U2962 (N_2962,N_1220,N_1543);
and U2963 (N_2963,N_762,N_260);
nor U2964 (N_2964,N_1473,N_90);
and U2965 (N_2965,N_1681,N_560);
nor U2966 (N_2966,N_650,N_1115);
nor U2967 (N_2967,N_1827,N_1847);
nand U2968 (N_2968,N_1664,N_1471);
nand U2969 (N_2969,N_216,N_1944);
nand U2970 (N_2970,N_279,N_478);
nand U2971 (N_2971,N_1845,N_1725);
nand U2972 (N_2972,N_1715,N_1737);
nand U2973 (N_2973,N_646,N_258);
and U2974 (N_2974,N_352,N_1729);
and U2975 (N_2975,N_1861,N_874);
nand U2976 (N_2976,N_1977,N_1868);
nor U2977 (N_2977,N_809,N_1516);
or U2978 (N_2978,N_1821,N_308);
and U2979 (N_2979,N_1844,N_225);
nor U2980 (N_2980,N_572,N_69);
nand U2981 (N_2981,N_1258,N_482);
nor U2982 (N_2982,N_373,N_983);
nor U2983 (N_2983,N_550,N_1602);
nor U2984 (N_2984,N_726,N_1852);
or U2985 (N_2985,N_1717,N_1384);
or U2986 (N_2986,N_1441,N_1885);
nand U2987 (N_2987,N_846,N_53);
and U2988 (N_2988,N_1379,N_1025);
and U2989 (N_2989,N_266,N_935);
nor U2990 (N_2990,N_757,N_1284);
and U2991 (N_2991,N_1714,N_152);
nand U2992 (N_2992,N_1504,N_401);
nor U2993 (N_2993,N_349,N_1691);
nor U2994 (N_2994,N_1872,N_388);
and U2995 (N_2995,N_882,N_1089);
and U2996 (N_2996,N_1671,N_1287);
and U2997 (N_2997,N_656,N_187);
or U2998 (N_2998,N_445,N_113);
nor U2999 (N_2999,N_781,N_1673);
or U3000 (N_3000,N_775,N_173);
nor U3001 (N_3001,N_360,N_1666);
nand U3002 (N_3002,N_913,N_1178);
and U3003 (N_3003,N_63,N_1347);
nor U3004 (N_3004,N_396,N_1571);
or U3005 (N_3005,N_1621,N_1744);
and U3006 (N_3006,N_649,N_1401);
nor U3007 (N_3007,N_182,N_960);
nand U3008 (N_3008,N_1429,N_1137);
nand U3009 (N_3009,N_813,N_1445);
or U3010 (N_3010,N_1047,N_361);
nor U3011 (N_3011,N_1845,N_1899);
nor U3012 (N_3012,N_1769,N_921);
or U3013 (N_3013,N_1888,N_828);
or U3014 (N_3014,N_718,N_1454);
and U3015 (N_3015,N_55,N_1863);
and U3016 (N_3016,N_1148,N_845);
or U3017 (N_3017,N_1415,N_1157);
nor U3018 (N_3018,N_1140,N_246);
nor U3019 (N_3019,N_295,N_728);
nor U3020 (N_3020,N_1286,N_160);
nor U3021 (N_3021,N_410,N_1685);
or U3022 (N_3022,N_904,N_188);
and U3023 (N_3023,N_1302,N_1876);
or U3024 (N_3024,N_1503,N_1641);
nor U3025 (N_3025,N_483,N_1384);
and U3026 (N_3026,N_1324,N_1655);
or U3027 (N_3027,N_1399,N_763);
and U3028 (N_3028,N_936,N_1026);
and U3029 (N_3029,N_1355,N_1842);
and U3030 (N_3030,N_360,N_1257);
nor U3031 (N_3031,N_686,N_239);
xnor U3032 (N_3032,N_443,N_471);
xnor U3033 (N_3033,N_214,N_1384);
or U3034 (N_3034,N_865,N_240);
or U3035 (N_3035,N_1241,N_1580);
nand U3036 (N_3036,N_1886,N_1296);
nor U3037 (N_3037,N_880,N_1285);
and U3038 (N_3038,N_1538,N_21);
nand U3039 (N_3039,N_645,N_158);
or U3040 (N_3040,N_1829,N_1399);
nand U3041 (N_3041,N_952,N_1916);
or U3042 (N_3042,N_551,N_1635);
and U3043 (N_3043,N_135,N_1761);
nand U3044 (N_3044,N_306,N_791);
or U3045 (N_3045,N_942,N_835);
nand U3046 (N_3046,N_816,N_805);
or U3047 (N_3047,N_1440,N_1507);
nand U3048 (N_3048,N_1528,N_1708);
nor U3049 (N_3049,N_924,N_1305);
nor U3050 (N_3050,N_1232,N_1546);
or U3051 (N_3051,N_603,N_1469);
nor U3052 (N_3052,N_1463,N_663);
or U3053 (N_3053,N_1866,N_538);
nor U3054 (N_3054,N_1863,N_806);
or U3055 (N_3055,N_1164,N_147);
nand U3056 (N_3056,N_79,N_802);
xnor U3057 (N_3057,N_1250,N_94);
or U3058 (N_3058,N_1694,N_1192);
nand U3059 (N_3059,N_1741,N_1961);
or U3060 (N_3060,N_203,N_1386);
and U3061 (N_3061,N_1605,N_814);
or U3062 (N_3062,N_371,N_154);
and U3063 (N_3063,N_62,N_93);
or U3064 (N_3064,N_1697,N_1286);
nand U3065 (N_3065,N_1868,N_877);
nand U3066 (N_3066,N_1153,N_1033);
nor U3067 (N_3067,N_1304,N_452);
or U3068 (N_3068,N_28,N_1886);
or U3069 (N_3069,N_1543,N_866);
nor U3070 (N_3070,N_1961,N_1297);
and U3071 (N_3071,N_945,N_983);
and U3072 (N_3072,N_1623,N_1700);
and U3073 (N_3073,N_794,N_1921);
nor U3074 (N_3074,N_1462,N_351);
and U3075 (N_3075,N_36,N_117);
nor U3076 (N_3076,N_26,N_1275);
and U3077 (N_3077,N_1372,N_396);
nor U3078 (N_3078,N_618,N_499);
nor U3079 (N_3079,N_144,N_666);
xor U3080 (N_3080,N_1382,N_695);
or U3081 (N_3081,N_764,N_931);
and U3082 (N_3082,N_1533,N_580);
nor U3083 (N_3083,N_435,N_1296);
and U3084 (N_3084,N_680,N_426);
or U3085 (N_3085,N_952,N_1663);
or U3086 (N_3086,N_1540,N_495);
nand U3087 (N_3087,N_1192,N_258);
and U3088 (N_3088,N_1942,N_1622);
nand U3089 (N_3089,N_904,N_1103);
and U3090 (N_3090,N_532,N_215);
nand U3091 (N_3091,N_1122,N_169);
and U3092 (N_3092,N_277,N_1201);
or U3093 (N_3093,N_765,N_1675);
nor U3094 (N_3094,N_265,N_125);
or U3095 (N_3095,N_397,N_1934);
xnor U3096 (N_3096,N_1752,N_779);
and U3097 (N_3097,N_163,N_409);
nand U3098 (N_3098,N_518,N_2);
nor U3099 (N_3099,N_403,N_1851);
and U3100 (N_3100,N_875,N_691);
nor U3101 (N_3101,N_328,N_978);
nand U3102 (N_3102,N_1189,N_1374);
and U3103 (N_3103,N_916,N_634);
nand U3104 (N_3104,N_62,N_454);
nor U3105 (N_3105,N_757,N_1131);
nor U3106 (N_3106,N_803,N_1885);
or U3107 (N_3107,N_450,N_1218);
or U3108 (N_3108,N_495,N_1346);
and U3109 (N_3109,N_1726,N_193);
nor U3110 (N_3110,N_1291,N_1580);
xnor U3111 (N_3111,N_1091,N_1796);
nand U3112 (N_3112,N_1179,N_1287);
nand U3113 (N_3113,N_248,N_523);
nor U3114 (N_3114,N_587,N_250);
or U3115 (N_3115,N_1566,N_943);
nor U3116 (N_3116,N_701,N_1040);
and U3117 (N_3117,N_208,N_62);
or U3118 (N_3118,N_918,N_1450);
and U3119 (N_3119,N_881,N_674);
nor U3120 (N_3120,N_370,N_1884);
nand U3121 (N_3121,N_912,N_1434);
or U3122 (N_3122,N_1705,N_1858);
nand U3123 (N_3123,N_951,N_75);
nand U3124 (N_3124,N_990,N_597);
and U3125 (N_3125,N_97,N_1000);
or U3126 (N_3126,N_1966,N_1359);
or U3127 (N_3127,N_554,N_1841);
nor U3128 (N_3128,N_871,N_1689);
nand U3129 (N_3129,N_1927,N_531);
nand U3130 (N_3130,N_1253,N_620);
nor U3131 (N_3131,N_745,N_1116);
and U3132 (N_3132,N_159,N_1696);
or U3133 (N_3133,N_188,N_1372);
or U3134 (N_3134,N_504,N_594);
or U3135 (N_3135,N_420,N_484);
nand U3136 (N_3136,N_1505,N_1124);
nor U3137 (N_3137,N_1063,N_656);
nand U3138 (N_3138,N_727,N_1550);
nand U3139 (N_3139,N_1571,N_1293);
and U3140 (N_3140,N_960,N_1483);
and U3141 (N_3141,N_1140,N_1145);
and U3142 (N_3142,N_1934,N_1805);
nand U3143 (N_3143,N_589,N_234);
nor U3144 (N_3144,N_1970,N_1731);
nor U3145 (N_3145,N_1671,N_643);
nor U3146 (N_3146,N_1963,N_1586);
or U3147 (N_3147,N_937,N_547);
nor U3148 (N_3148,N_1495,N_1212);
nor U3149 (N_3149,N_564,N_1973);
nand U3150 (N_3150,N_513,N_832);
nand U3151 (N_3151,N_1167,N_1223);
nand U3152 (N_3152,N_650,N_1202);
and U3153 (N_3153,N_1745,N_538);
nand U3154 (N_3154,N_1800,N_1029);
or U3155 (N_3155,N_910,N_1375);
nor U3156 (N_3156,N_494,N_1491);
and U3157 (N_3157,N_269,N_1059);
nor U3158 (N_3158,N_258,N_1675);
and U3159 (N_3159,N_1170,N_1994);
nand U3160 (N_3160,N_1880,N_707);
nand U3161 (N_3161,N_604,N_1024);
nand U3162 (N_3162,N_450,N_359);
and U3163 (N_3163,N_1764,N_1111);
nand U3164 (N_3164,N_525,N_265);
or U3165 (N_3165,N_271,N_814);
and U3166 (N_3166,N_268,N_892);
and U3167 (N_3167,N_52,N_1008);
nor U3168 (N_3168,N_1706,N_195);
nand U3169 (N_3169,N_1803,N_1226);
nand U3170 (N_3170,N_1845,N_997);
nor U3171 (N_3171,N_1881,N_1915);
nor U3172 (N_3172,N_746,N_329);
and U3173 (N_3173,N_80,N_1377);
nor U3174 (N_3174,N_1918,N_463);
nand U3175 (N_3175,N_650,N_671);
nor U3176 (N_3176,N_350,N_939);
nand U3177 (N_3177,N_835,N_462);
and U3178 (N_3178,N_1956,N_1301);
or U3179 (N_3179,N_293,N_1010);
and U3180 (N_3180,N_916,N_1049);
or U3181 (N_3181,N_815,N_345);
and U3182 (N_3182,N_905,N_1455);
nand U3183 (N_3183,N_10,N_582);
nand U3184 (N_3184,N_871,N_441);
or U3185 (N_3185,N_117,N_1111);
nor U3186 (N_3186,N_1272,N_1025);
or U3187 (N_3187,N_1415,N_1408);
and U3188 (N_3188,N_626,N_102);
nor U3189 (N_3189,N_220,N_1624);
or U3190 (N_3190,N_96,N_752);
and U3191 (N_3191,N_1540,N_1486);
nand U3192 (N_3192,N_1379,N_1408);
nand U3193 (N_3193,N_1457,N_974);
nor U3194 (N_3194,N_1673,N_983);
or U3195 (N_3195,N_115,N_236);
and U3196 (N_3196,N_1318,N_271);
nand U3197 (N_3197,N_880,N_728);
nor U3198 (N_3198,N_259,N_1968);
or U3199 (N_3199,N_616,N_1772);
nand U3200 (N_3200,N_1334,N_109);
or U3201 (N_3201,N_604,N_1534);
and U3202 (N_3202,N_876,N_1536);
or U3203 (N_3203,N_670,N_42);
nand U3204 (N_3204,N_1287,N_1748);
nor U3205 (N_3205,N_1866,N_1611);
and U3206 (N_3206,N_1880,N_347);
or U3207 (N_3207,N_690,N_1005);
nor U3208 (N_3208,N_862,N_175);
nand U3209 (N_3209,N_1360,N_1952);
xnor U3210 (N_3210,N_1844,N_836);
or U3211 (N_3211,N_1021,N_1029);
nor U3212 (N_3212,N_1495,N_1230);
and U3213 (N_3213,N_144,N_675);
and U3214 (N_3214,N_111,N_596);
nor U3215 (N_3215,N_420,N_1989);
nand U3216 (N_3216,N_1313,N_457);
nor U3217 (N_3217,N_1015,N_1896);
nand U3218 (N_3218,N_761,N_826);
nand U3219 (N_3219,N_651,N_1152);
nor U3220 (N_3220,N_868,N_30);
and U3221 (N_3221,N_1246,N_1086);
nor U3222 (N_3222,N_121,N_1033);
and U3223 (N_3223,N_1798,N_709);
nand U3224 (N_3224,N_405,N_196);
or U3225 (N_3225,N_1357,N_1989);
nand U3226 (N_3226,N_829,N_1061);
nor U3227 (N_3227,N_1240,N_1062);
or U3228 (N_3228,N_1967,N_1162);
nor U3229 (N_3229,N_437,N_542);
or U3230 (N_3230,N_1985,N_801);
nand U3231 (N_3231,N_1222,N_1480);
nand U3232 (N_3232,N_1798,N_269);
nand U3233 (N_3233,N_1286,N_949);
and U3234 (N_3234,N_923,N_1461);
and U3235 (N_3235,N_474,N_1711);
xnor U3236 (N_3236,N_1579,N_130);
xnor U3237 (N_3237,N_852,N_1728);
or U3238 (N_3238,N_869,N_1003);
nor U3239 (N_3239,N_38,N_1966);
nor U3240 (N_3240,N_264,N_143);
and U3241 (N_3241,N_1781,N_698);
or U3242 (N_3242,N_234,N_1532);
or U3243 (N_3243,N_1879,N_745);
and U3244 (N_3244,N_265,N_354);
nor U3245 (N_3245,N_1236,N_255);
or U3246 (N_3246,N_347,N_187);
nor U3247 (N_3247,N_1415,N_1173);
or U3248 (N_3248,N_1984,N_1850);
nor U3249 (N_3249,N_1661,N_1010);
nor U3250 (N_3250,N_742,N_217);
xor U3251 (N_3251,N_986,N_503);
nor U3252 (N_3252,N_1351,N_1541);
nor U3253 (N_3253,N_1078,N_244);
or U3254 (N_3254,N_97,N_1935);
nor U3255 (N_3255,N_806,N_864);
or U3256 (N_3256,N_474,N_120);
nor U3257 (N_3257,N_1534,N_1377);
nand U3258 (N_3258,N_532,N_1469);
nand U3259 (N_3259,N_1085,N_264);
nand U3260 (N_3260,N_92,N_1239);
nand U3261 (N_3261,N_1713,N_1882);
nand U3262 (N_3262,N_1448,N_351);
nor U3263 (N_3263,N_1094,N_860);
nand U3264 (N_3264,N_943,N_366);
nor U3265 (N_3265,N_6,N_513);
and U3266 (N_3266,N_133,N_1956);
and U3267 (N_3267,N_799,N_450);
nor U3268 (N_3268,N_193,N_1208);
and U3269 (N_3269,N_295,N_846);
and U3270 (N_3270,N_832,N_1327);
or U3271 (N_3271,N_907,N_1093);
or U3272 (N_3272,N_82,N_436);
nor U3273 (N_3273,N_217,N_725);
nor U3274 (N_3274,N_726,N_1305);
nand U3275 (N_3275,N_1820,N_130);
nor U3276 (N_3276,N_758,N_297);
or U3277 (N_3277,N_1712,N_1083);
and U3278 (N_3278,N_670,N_1874);
nand U3279 (N_3279,N_737,N_1167);
nand U3280 (N_3280,N_565,N_1762);
and U3281 (N_3281,N_652,N_1672);
nand U3282 (N_3282,N_1728,N_663);
nor U3283 (N_3283,N_1695,N_757);
and U3284 (N_3284,N_1663,N_258);
nor U3285 (N_3285,N_282,N_1371);
and U3286 (N_3286,N_1379,N_335);
or U3287 (N_3287,N_399,N_1844);
nor U3288 (N_3288,N_1538,N_25);
or U3289 (N_3289,N_681,N_83);
nand U3290 (N_3290,N_1525,N_1141);
and U3291 (N_3291,N_1328,N_1596);
nor U3292 (N_3292,N_592,N_1108);
nor U3293 (N_3293,N_1259,N_1944);
nor U3294 (N_3294,N_271,N_951);
or U3295 (N_3295,N_279,N_1258);
nor U3296 (N_3296,N_1200,N_612);
or U3297 (N_3297,N_1048,N_1721);
and U3298 (N_3298,N_1402,N_1149);
and U3299 (N_3299,N_614,N_443);
or U3300 (N_3300,N_1438,N_1457);
and U3301 (N_3301,N_1996,N_27);
nor U3302 (N_3302,N_493,N_1527);
and U3303 (N_3303,N_1371,N_1460);
nor U3304 (N_3304,N_983,N_1801);
nor U3305 (N_3305,N_1420,N_48);
or U3306 (N_3306,N_1314,N_1106);
and U3307 (N_3307,N_797,N_98);
or U3308 (N_3308,N_655,N_1935);
xor U3309 (N_3309,N_1058,N_234);
and U3310 (N_3310,N_1680,N_1454);
nor U3311 (N_3311,N_307,N_105);
or U3312 (N_3312,N_1856,N_463);
nand U3313 (N_3313,N_1673,N_309);
nor U3314 (N_3314,N_1707,N_147);
nand U3315 (N_3315,N_512,N_1752);
and U3316 (N_3316,N_561,N_647);
nor U3317 (N_3317,N_1522,N_1128);
nor U3318 (N_3318,N_1123,N_230);
xor U3319 (N_3319,N_1959,N_1249);
and U3320 (N_3320,N_1879,N_760);
or U3321 (N_3321,N_578,N_1645);
and U3322 (N_3322,N_1244,N_251);
or U3323 (N_3323,N_829,N_178);
nor U3324 (N_3324,N_922,N_459);
and U3325 (N_3325,N_1086,N_1394);
and U3326 (N_3326,N_1619,N_1001);
or U3327 (N_3327,N_866,N_1337);
nand U3328 (N_3328,N_949,N_78);
nor U3329 (N_3329,N_1892,N_399);
nand U3330 (N_3330,N_1831,N_1989);
or U3331 (N_3331,N_318,N_940);
nand U3332 (N_3332,N_1888,N_640);
nor U3333 (N_3333,N_11,N_543);
or U3334 (N_3334,N_1975,N_1466);
or U3335 (N_3335,N_1946,N_133);
and U3336 (N_3336,N_301,N_380);
nand U3337 (N_3337,N_602,N_909);
or U3338 (N_3338,N_40,N_1291);
nor U3339 (N_3339,N_599,N_1547);
nor U3340 (N_3340,N_1234,N_810);
or U3341 (N_3341,N_702,N_781);
nor U3342 (N_3342,N_704,N_1403);
or U3343 (N_3343,N_1618,N_147);
nand U3344 (N_3344,N_657,N_1844);
and U3345 (N_3345,N_581,N_1897);
nand U3346 (N_3346,N_1250,N_1751);
and U3347 (N_3347,N_1328,N_788);
or U3348 (N_3348,N_1788,N_1096);
nor U3349 (N_3349,N_1490,N_1294);
nor U3350 (N_3350,N_1848,N_1463);
nand U3351 (N_3351,N_413,N_1220);
and U3352 (N_3352,N_1108,N_330);
nand U3353 (N_3353,N_738,N_127);
nor U3354 (N_3354,N_1123,N_1116);
and U3355 (N_3355,N_1269,N_982);
nor U3356 (N_3356,N_508,N_1649);
and U3357 (N_3357,N_896,N_326);
or U3358 (N_3358,N_904,N_760);
nand U3359 (N_3359,N_1242,N_1844);
nor U3360 (N_3360,N_757,N_240);
and U3361 (N_3361,N_741,N_1310);
and U3362 (N_3362,N_43,N_1052);
and U3363 (N_3363,N_529,N_992);
and U3364 (N_3364,N_677,N_1614);
nand U3365 (N_3365,N_1225,N_1557);
or U3366 (N_3366,N_1365,N_861);
and U3367 (N_3367,N_1475,N_373);
and U3368 (N_3368,N_1969,N_546);
or U3369 (N_3369,N_1995,N_1993);
and U3370 (N_3370,N_1105,N_49);
nor U3371 (N_3371,N_926,N_1964);
nor U3372 (N_3372,N_530,N_995);
nand U3373 (N_3373,N_334,N_602);
or U3374 (N_3374,N_256,N_535);
nand U3375 (N_3375,N_1000,N_1620);
and U3376 (N_3376,N_1343,N_1006);
nor U3377 (N_3377,N_1104,N_908);
or U3378 (N_3378,N_1658,N_239);
nor U3379 (N_3379,N_1737,N_79);
nor U3380 (N_3380,N_1782,N_622);
nor U3381 (N_3381,N_784,N_1367);
and U3382 (N_3382,N_850,N_1181);
nand U3383 (N_3383,N_1352,N_1544);
nor U3384 (N_3384,N_1605,N_880);
nand U3385 (N_3385,N_1966,N_1214);
or U3386 (N_3386,N_322,N_1892);
or U3387 (N_3387,N_1042,N_1089);
nor U3388 (N_3388,N_908,N_1243);
nor U3389 (N_3389,N_748,N_1834);
and U3390 (N_3390,N_1719,N_1112);
nand U3391 (N_3391,N_177,N_96);
or U3392 (N_3392,N_756,N_740);
nand U3393 (N_3393,N_787,N_288);
nor U3394 (N_3394,N_649,N_1750);
xnor U3395 (N_3395,N_544,N_502);
and U3396 (N_3396,N_853,N_25);
nor U3397 (N_3397,N_1243,N_1666);
nand U3398 (N_3398,N_1789,N_1468);
and U3399 (N_3399,N_1163,N_1412);
nand U3400 (N_3400,N_1810,N_820);
nand U3401 (N_3401,N_135,N_1523);
or U3402 (N_3402,N_716,N_1329);
nor U3403 (N_3403,N_745,N_354);
and U3404 (N_3404,N_1421,N_1414);
or U3405 (N_3405,N_1032,N_1177);
and U3406 (N_3406,N_587,N_524);
nor U3407 (N_3407,N_104,N_1828);
or U3408 (N_3408,N_1233,N_645);
nand U3409 (N_3409,N_16,N_400);
and U3410 (N_3410,N_1512,N_354);
or U3411 (N_3411,N_238,N_1060);
nand U3412 (N_3412,N_1252,N_1977);
nand U3413 (N_3413,N_27,N_1889);
and U3414 (N_3414,N_1137,N_1559);
xnor U3415 (N_3415,N_1737,N_1341);
nand U3416 (N_3416,N_1799,N_1895);
nand U3417 (N_3417,N_379,N_878);
nor U3418 (N_3418,N_1365,N_536);
nor U3419 (N_3419,N_1793,N_1018);
nor U3420 (N_3420,N_508,N_1628);
and U3421 (N_3421,N_306,N_1830);
nor U3422 (N_3422,N_712,N_543);
or U3423 (N_3423,N_496,N_580);
nor U3424 (N_3424,N_41,N_285);
nand U3425 (N_3425,N_34,N_1156);
or U3426 (N_3426,N_237,N_1436);
nor U3427 (N_3427,N_183,N_391);
and U3428 (N_3428,N_32,N_225);
nand U3429 (N_3429,N_1111,N_1760);
nor U3430 (N_3430,N_636,N_567);
nor U3431 (N_3431,N_691,N_360);
or U3432 (N_3432,N_1690,N_363);
nand U3433 (N_3433,N_321,N_1537);
and U3434 (N_3434,N_233,N_588);
nor U3435 (N_3435,N_1225,N_729);
and U3436 (N_3436,N_830,N_1830);
and U3437 (N_3437,N_1469,N_1940);
nor U3438 (N_3438,N_1901,N_1879);
nor U3439 (N_3439,N_604,N_8);
or U3440 (N_3440,N_1021,N_1193);
or U3441 (N_3441,N_721,N_280);
nand U3442 (N_3442,N_644,N_752);
and U3443 (N_3443,N_1962,N_1096);
or U3444 (N_3444,N_921,N_892);
or U3445 (N_3445,N_1420,N_431);
nor U3446 (N_3446,N_1710,N_1038);
or U3447 (N_3447,N_1006,N_1568);
nand U3448 (N_3448,N_1476,N_818);
nor U3449 (N_3449,N_1105,N_119);
nor U3450 (N_3450,N_1735,N_1570);
nor U3451 (N_3451,N_608,N_1242);
or U3452 (N_3452,N_693,N_140);
or U3453 (N_3453,N_828,N_1644);
nor U3454 (N_3454,N_866,N_1041);
nand U3455 (N_3455,N_1026,N_95);
nand U3456 (N_3456,N_1309,N_1579);
nand U3457 (N_3457,N_247,N_1827);
nand U3458 (N_3458,N_1913,N_304);
or U3459 (N_3459,N_713,N_1003);
nor U3460 (N_3460,N_1560,N_1254);
xnor U3461 (N_3461,N_1569,N_1525);
nor U3462 (N_3462,N_1285,N_924);
nand U3463 (N_3463,N_564,N_1886);
or U3464 (N_3464,N_776,N_1243);
or U3465 (N_3465,N_499,N_1973);
and U3466 (N_3466,N_1525,N_1600);
or U3467 (N_3467,N_1369,N_1900);
nand U3468 (N_3468,N_311,N_540);
nor U3469 (N_3469,N_1236,N_647);
nor U3470 (N_3470,N_340,N_1574);
or U3471 (N_3471,N_1440,N_122);
nand U3472 (N_3472,N_562,N_1560);
nor U3473 (N_3473,N_981,N_1973);
nand U3474 (N_3474,N_620,N_708);
nand U3475 (N_3475,N_1107,N_1507);
nor U3476 (N_3476,N_1627,N_439);
nand U3477 (N_3477,N_1917,N_259);
or U3478 (N_3478,N_42,N_1922);
nor U3479 (N_3479,N_1431,N_534);
and U3480 (N_3480,N_210,N_363);
nand U3481 (N_3481,N_1656,N_772);
nand U3482 (N_3482,N_623,N_700);
nand U3483 (N_3483,N_1327,N_300);
xor U3484 (N_3484,N_1369,N_468);
or U3485 (N_3485,N_1988,N_1368);
or U3486 (N_3486,N_104,N_1433);
nand U3487 (N_3487,N_1881,N_1180);
nand U3488 (N_3488,N_921,N_1114);
or U3489 (N_3489,N_1503,N_1836);
nor U3490 (N_3490,N_1530,N_788);
nand U3491 (N_3491,N_1902,N_695);
or U3492 (N_3492,N_404,N_517);
nand U3493 (N_3493,N_809,N_1151);
or U3494 (N_3494,N_1572,N_1139);
or U3495 (N_3495,N_1194,N_275);
nand U3496 (N_3496,N_1856,N_1200);
nor U3497 (N_3497,N_647,N_1889);
and U3498 (N_3498,N_1421,N_1537);
or U3499 (N_3499,N_1014,N_1829);
nand U3500 (N_3500,N_567,N_1530);
nor U3501 (N_3501,N_1663,N_220);
and U3502 (N_3502,N_934,N_702);
xnor U3503 (N_3503,N_727,N_1700);
or U3504 (N_3504,N_461,N_1667);
xor U3505 (N_3505,N_1859,N_543);
and U3506 (N_3506,N_421,N_1585);
or U3507 (N_3507,N_1586,N_74);
and U3508 (N_3508,N_1748,N_1244);
and U3509 (N_3509,N_1758,N_341);
or U3510 (N_3510,N_147,N_834);
nand U3511 (N_3511,N_1473,N_613);
nand U3512 (N_3512,N_789,N_1205);
and U3513 (N_3513,N_1140,N_179);
nand U3514 (N_3514,N_1563,N_961);
nand U3515 (N_3515,N_1419,N_929);
and U3516 (N_3516,N_421,N_1359);
or U3517 (N_3517,N_213,N_1533);
nand U3518 (N_3518,N_1673,N_1697);
nand U3519 (N_3519,N_1355,N_214);
nor U3520 (N_3520,N_1651,N_876);
nor U3521 (N_3521,N_1261,N_618);
nor U3522 (N_3522,N_413,N_23);
or U3523 (N_3523,N_882,N_209);
nand U3524 (N_3524,N_1014,N_771);
nand U3525 (N_3525,N_1015,N_1484);
nand U3526 (N_3526,N_99,N_1935);
nand U3527 (N_3527,N_1755,N_1045);
nor U3528 (N_3528,N_715,N_426);
and U3529 (N_3529,N_1630,N_203);
nor U3530 (N_3530,N_841,N_1746);
and U3531 (N_3531,N_646,N_1273);
nor U3532 (N_3532,N_790,N_370);
or U3533 (N_3533,N_1427,N_1050);
and U3534 (N_3534,N_1660,N_740);
or U3535 (N_3535,N_1100,N_659);
nand U3536 (N_3536,N_818,N_416);
and U3537 (N_3537,N_938,N_1118);
or U3538 (N_3538,N_3,N_728);
nand U3539 (N_3539,N_291,N_1806);
nor U3540 (N_3540,N_1475,N_1999);
and U3541 (N_3541,N_91,N_573);
and U3542 (N_3542,N_879,N_234);
nor U3543 (N_3543,N_1099,N_1426);
and U3544 (N_3544,N_35,N_140);
nor U3545 (N_3545,N_1091,N_121);
nor U3546 (N_3546,N_1439,N_407);
nand U3547 (N_3547,N_539,N_710);
nor U3548 (N_3548,N_1632,N_1833);
and U3549 (N_3549,N_654,N_13);
nand U3550 (N_3550,N_1807,N_1960);
or U3551 (N_3551,N_1759,N_1039);
nor U3552 (N_3552,N_1432,N_1496);
or U3553 (N_3553,N_732,N_1624);
or U3554 (N_3554,N_543,N_1286);
and U3555 (N_3555,N_461,N_163);
nand U3556 (N_3556,N_532,N_645);
nand U3557 (N_3557,N_395,N_916);
or U3558 (N_3558,N_1544,N_1942);
and U3559 (N_3559,N_977,N_1395);
nor U3560 (N_3560,N_1069,N_309);
nor U3561 (N_3561,N_1465,N_536);
and U3562 (N_3562,N_1902,N_756);
nand U3563 (N_3563,N_1789,N_527);
and U3564 (N_3564,N_1347,N_211);
nor U3565 (N_3565,N_746,N_849);
nor U3566 (N_3566,N_1860,N_1050);
nand U3567 (N_3567,N_790,N_114);
nor U3568 (N_3568,N_1640,N_599);
or U3569 (N_3569,N_246,N_362);
nor U3570 (N_3570,N_793,N_195);
nand U3571 (N_3571,N_689,N_792);
or U3572 (N_3572,N_819,N_1112);
and U3573 (N_3573,N_1973,N_802);
and U3574 (N_3574,N_1831,N_1142);
nand U3575 (N_3575,N_793,N_1593);
nor U3576 (N_3576,N_1274,N_365);
or U3577 (N_3577,N_691,N_1678);
or U3578 (N_3578,N_884,N_1197);
or U3579 (N_3579,N_1530,N_468);
xnor U3580 (N_3580,N_385,N_1153);
nand U3581 (N_3581,N_76,N_358);
and U3582 (N_3582,N_1188,N_431);
nand U3583 (N_3583,N_1703,N_372);
nor U3584 (N_3584,N_1738,N_482);
and U3585 (N_3585,N_1732,N_955);
or U3586 (N_3586,N_1329,N_343);
nor U3587 (N_3587,N_1361,N_1502);
and U3588 (N_3588,N_1298,N_1565);
or U3589 (N_3589,N_1885,N_1282);
and U3590 (N_3590,N_383,N_1419);
nand U3591 (N_3591,N_1827,N_115);
nand U3592 (N_3592,N_1547,N_797);
and U3593 (N_3593,N_926,N_733);
nor U3594 (N_3594,N_1207,N_1429);
nor U3595 (N_3595,N_1976,N_1645);
nand U3596 (N_3596,N_1636,N_1388);
and U3597 (N_3597,N_1434,N_735);
or U3598 (N_3598,N_1033,N_797);
and U3599 (N_3599,N_1155,N_1482);
nor U3600 (N_3600,N_55,N_568);
nand U3601 (N_3601,N_1030,N_1240);
or U3602 (N_3602,N_84,N_1105);
nor U3603 (N_3603,N_1417,N_325);
and U3604 (N_3604,N_1661,N_819);
nand U3605 (N_3605,N_1358,N_730);
nor U3606 (N_3606,N_1526,N_1819);
or U3607 (N_3607,N_317,N_1593);
and U3608 (N_3608,N_913,N_1908);
and U3609 (N_3609,N_1506,N_1408);
or U3610 (N_3610,N_223,N_384);
nor U3611 (N_3611,N_404,N_122);
and U3612 (N_3612,N_394,N_1224);
nand U3613 (N_3613,N_1826,N_418);
nand U3614 (N_3614,N_1563,N_903);
nand U3615 (N_3615,N_1551,N_1483);
nor U3616 (N_3616,N_677,N_826);
nand U3617 (N_3617,N_514,N_1833);
nand U3618 (N_3618,N_1085,N_1585);
nand U3619 (N_3619,N_936,N_1497);
nor U3620 (N_3620,N_132,N_684);
nor U3621 (N_3621,N_619,N_969);
nor U3622 (N_3622,N_1387,N_688);
and U3623 (N_3623,N_1292,N_1341);
nand U3624 (N_3624,N_1272,N_97);
and U3625 (N_3625,N_1168,N_1664);
and U3626 (N_3626,N_427,N_230);
nor U3627 (N_3627,N_1928,N_1166);
or U3628 (N_3628,N_755,N_1015);
or U3629 (N_3629,N_1695,N_169);
or U3630 (N_3630,N_1468,N_1217);
nor U3631 (N_3631,N_1736,N_1497);
nor U3632 (N_3632,N_1663,N_1834);
and U3633 (N_3633,N_1045,N_1946);
or U3634 (N_3634,N_1543,N_711);
or U3635 (N_3635,N_1392,N_1517);
nor U3636 (N_3636,N_740,N_1228);
nor U3637 (N_3637,N_257,N_864);
and U3638 (N_3638,N_1919,N_1581);
nand U3639 (N_3639,N_1473,N_1838);
and U3640 (N_3640,N_1075,N_1313);
and U3641 (N_3641,N_899,N_442);
or U3642 (N_3642,N_1759,N_665);
and U3643 (N_3643,N_1574,N_1340);
nor U3644 (N_3644,N_1296,N_1519);
or U3645 (N_3645,N_1008,N_1000);
nand U3646 (N_3646,N_1385,N_824);
nand U3647 (N_3647,N_817,N_846);
or U3648 (N_3648,N_1358,N_36);
nand U3649 (N_3649,N_283,N_1931);
or U3650 (N_3650,N_825,N_98);
nor U3651 (N_3651,N_1760,N_1764);
and U3652 (N_3652,N_1988,N_36);
or U3653 (N_3653,N_874,N_820);
nand U3654 (N_3654,N_785,N_761);
and U3655 (N_3655,N_683,N_1620);
or U3656 (N_3656,N_1496,N_953);
nand U3657 (N_3657,N_1855,N_941);
nand U3658 (N_3658,N_577,N_420);
nand U3659 (N_3659,N_1424,N_1252);
nor U3660 (N_3660,N_1604,N_665);
and U3661 (N_3661,N_957,N_1326);
nand U3662 (N_3662,N_1717,N_327);
and U3663 (N_3663,N_340,N_1043);
nand U3664 (N_3664,N_742,N_988);
and U3665 (N_3665,N_180,N_623);
nor U3666 (N_3666,N_550,N_543);
and U3667 (N_3667,N_565,N_408);
nor U3668 (N_3668,N_234,N_19);
nand U3669 (N_3669,N_614,N_1335);
nand U3670 (N_3670,N_360,N_259);
or U3671 (N_3671,N_1149,N_1397);
nor U3672 (N_3672,N_487,N_814);
or U3673 (N_3673,N_1604,N_853);
nand U3674 (N_3674,N_1510,N_1743);
nand U3675 (N_3675,N_536,N_1939);
and U3676 (N_3676,N_1886,N_614);
or U3677 (N_3677,N_1625,N_243);
nand U3678 (N_3678,N_505,N_1550);
nor U3679 (N_3679,N_817,N_1554);
xor U3680 (N_3680,N_1520,N_1704);
nor U3681 (N_3681,N_1374,N_1311);
nand U3682 (N_3682,N_1046,N_928);
nor U3683 (N_3683,N_1275,N_263);
or U3684 (N_3684,N_406,N_27);
nor U3685 (N_3685,N_92,N_1331);
or U3686 (N_3686,N_1911,N_63);
or U3687 (N_3687,N_1595,N_1302);
or U3688 (N_3688,N_900,N_1471);
nor U3689 (N_3689,N_827,N_833);
nor U3690 (N_3690,N_392,N_928);
or U3691 (N_3691,N_48,N_1740);
and U3692 (N_3692,N_137,N_1077);
or U3693 (N_3693,N_670,N_1970);
or U3694 (N_3694,N_1774,N_359);
nor U3695 (N_3695,N_1580,N_22);
and U3696 (N_3696,N_810,N_1142);
or U3697 (N_3697,N_464,N_1923);
and U3698 (N_3698,N_1709,N_205);
nand U3699 (N_3699,N_1244,N_577);
and U3700 (N_3700,N_709,N_1781);
or U3701 (N_3701,N_1979,N_1227);
nand U3702 (N_3702,N_1231,N_542);
and U3703 (N_3703,N_764,N_995);
nand U3704 (N_3704,N_1175,N_691);
and U3705 (N_3705,N_370,N_992);
and U3706 (N_3706,N_1029,N_1244);
nand U3707 (N_3707,N_917,N_1319);
and U3708 (N_3708,N_1620,N_964);
or U3709 (N_3709,N_1374,N_1233);
or U3710 (N_3710,N_289,N_1569);
or U3711 (N_3711,N_1403,N_112);
nand U3712 (N_3712,N_295,N_1702);
nor U3713 (N_3713,N_1929,N_192);
nand U3714 (N_3714,N_1583,N_797);
or U3715 (N_3715,N_772,N_1109);
or U3716 (N_3716,N_443,N_1777);
and U3717 (N_3717,N_1136,N_1573);
nor U3718 (N_3718,N_1074,N_1320);
nand U3719 (N_3719,N_841,N_1559);
or U3720 (N_3720,N_842,N_1661);
nor U3721 (N_3721,N_1658,N_53);
and U3722 (N_3722,N_1607,N_297);
nor U3723 (N_3723,N_1173,N_1202);
nand U3724 (N_3724,N_1860,N_961);
or U3725 (N_3725,N_1591,N_1255);
and U3726 (N_3726,N_1806,N_1007);
nand U3727 (N_3727,N_285,N_1719);
and U3728 (N_3728,N_1554,N_989);
nand U3729 (N_3729,N_1743,N_1414);
and U3730 (N_3730,N_314,N_816);
nor U3731 (N_3731,N_601,N_1103);
or U3732 (N_3732,N_1562,N_580);
and U3733 (N_3733,N_1239,N_1269);
nand U3734 (N_3734,N_1097,N_1218);
nand U3735 (N_3735,N_310,N_1391);
nor U3736 (N_3736,N_1487,N_1235);
and U3737 (N_3737,N_1707,N_1643);
and U3738 (N_3738,N_1848,N_1049);
or U3739 (N_3739,N_421,N_942);
or U3740 (N_3740,N_1676,N_1266);
and U3741 (N_3741,N_278,N_1578);
or U3742 (N_3742,N_89,N_1372);
xor U3743 (N_3743,N_1553,N_32);
nor U3744 (N_3744,N_1426,N_1971);
or U3745 (N_3745,N_1953,N_996);
and U3746 (N_3746,N_178,N_534);
or U3747 (N_3747,N_813,N_549);
nor U3748 (N_3748,N_506,N_1535);
and U3749 (N_3749,N_1906,N_1003);
or U3750 (N_3750,N_282,N_1946);
and U3751 (N_3751,N_1108,N_669);
or U3752 (N_3752,N_1085,N_1042);
nor U3753 (N_3753,N_1656,N_1175);
nor U3754 (N_3754,N_1600,N_1007);
or U3755 (N_3755,N_1689,N_670);
nor U3756 (N_3756,N_26,N_30);
or U3757 (N_3757,N_1602,N_1943);
xnor U3758 (N_3758,N_544,N_264);
nand U3759 (N_3759,N_1250,N_104);
nor U3760 (N_3760,N_1885,N_1991);
nand U3761 (N_3761,N_810,N_1195);
and U3762 (N_3762,N_1990,N_34);
and U3763 (N_3763,N_1406,N_18);
nor U3764 (N_3764,N_986,N_441);
and U3765 (N_3765,N_1335,N_1177);
or U3766 (N_3766,N_1832,N_1289);
or U3767 (N_3767,N_848,N_1980);
and U3768 (N_3768,N_1837,N_1357);
nor U3769 (N_3769,N_1714,N_200);
nor U3770 (N_3770,N_701,N_854);
or U3771 (N_3771,N_1612,N_600);
nor U3772 (N_3772,N_703,N_1181);
nand U3773 (N_3773,N_1401,N_1382);
nand U3774 (N_3774,N_1898,N_1287);
and U3775 (N_3775,N_1471,N_650);
and U3776 (N_3776,N_1244,N_6);
and U3777 (N_3777,N_345,N_868);
and U3778 (N_3778,N_1809,N_1592);
and U3779 (N_3779,N_1222,N_1381);
nand U3780 (N_3780,N_1653,N_1113);
or U3781 (N_3781,N_670,N_1244);
and U3782 (N_3782,N_768,N_1809);
and U3783 (N_3783,N_817,N_636);
nand U3784 (N_3784,N_1561,N_342);
nand U3785 (N_3785,N_1391,N_1404);
nor U3786 (N_3786,N_852,N_1299);
or U3787 (N_3787,N_1916,N_1688);
and U3788 (N_3788,N_1500,N_5);
nand U3789 (N_3789,N_1062,N_307);
or U3790 (N_3790,N_748,N_10);
nor U3791 (N_3791,N_1418,N_1443);
or U3792 (N_3792,N_219,N_75);
nand U3793 (N_3793,N_1572,N_1219);
or U3794 (N_3794,N_478,N_1639);
or U3795 (N_3795,N_1843,N_441);
or U3796 (N_3796,N_1556,N_919);
or U3797 (N_3797,N_1602,N_347);
or U3798 (N_3798,N_239,N_1870);
or U3799 (N_3799,N_1765,N_1157);
nand U3800 (N_3800,N_600,N_1064);
and U3801 (N_3801,N_191,N_1960);
or U3802 (N_3802,N_1938,N_511);
nand U3803 (N_3803,N_1523,N_1749);
or U3804 (N_3804,N_1006,N_436);
nor U3805 (N_3805,N_874,N_1576);
and U3806 (N_3806,N_1672,N_1094);
and U3807 (N_3807,N_325,N_791);
and U3808 (N_3808,N_1834,N_1863);
nor U3809 (N_3809,N_1411,N_1363);
and U3810 (N_3810,N_1067,N_1827);
nor U3811 (N_3811,N_1843,N_1735);
nor U3812 (N_3812,N_432,N_1562);
nor U3813 (N_3813,N_540,N_1356);
or U3814 (N_3814,N_1331,N_1599);
or U3815 (N_3815,N_1650,N_960);
or U3816 (N_3816,N_1044,N_1216);
nand U3817 (N_3817,N_1709,N_1037);
or U3818 (N_3818,N_1684,N_409);
nand U3819 (N_3819,N_31,N_1408);
and U3820 (N_3820,N_552,N_1522);
nor U3821 (N_3821,N_1131,N_602);
nor U3822 (N_3822,N_488,N_575);
and U3823 (N_3823,N_1170,N_1797);
and U3824 (N_3824,N_300,N_455);
nand U3825 (N_3825,N_29,N_537);
nand U3826 (N_3826,N_1107,N_1139);
and U3827 (N_3827,N_272,N_1960);
nor U3828 (N_3828,N_1495,N_761);
nor U3829 (N_3829,N_682,N_936);
or U3830 (N_3830,N_1688,N_1433);
and U3831 (N_3831,N_1012,N_93);
nor U3832 (N_3832,N_558,N_405);
and U3833 (N_3833,N_1930,N_1996);
or U3834 (N_3834,N_1535,N_444);
or U3835 (N_3835,N_206,N_1568);
and U3836 (N_3836,N_1244,N_764);
nand U3837 (N_3837,N_409,N_1782);
nor U3838 (N_3838,N_1525,N_615);
or U3839 (N_3839,N_1443,N_337);
nor U3840 (N_3840,N_253,N_1822);
and U3841 (N_3841,N_783,N_188);
nor U3842 (N_3842,N_492,N_722);
nor U3843 (N_3843,N_1523,N_343);
nand U3844 (N_3844,N_1450,N_1361);
and U3845 (N_3845,N_1915,N_390);
nand U3846 (N_3846,N_295,N_580);
nor U3847 (N_3847,N_1243,N_385);
or U3848 (N_3848,N_1609,N_419);
nor U3849 (N_3849,N_1690,N_1739);
or U3850 (N_3850,N_270,N_449);
nand U3851 (N_3851,N_1033,N_1986);
or U3852 (N_3852,N_1806,N_1560);
nor U3853 (N_3853,N_1739,N_742);
nor U3854 (N_3854,N_1339,N_1413);
and U3855 (N_3855,N_494,N_1957);
and U3856 (N_3856,N_1613,N_141);
or U3857 (N_3857,N_817,N_1949);
and U3858 (N_3858,N_1018,N_1092);
nand U3859 (N_3859,N_980,N_832);
or U3860 (N_3860,N_1565,N_1157);
nand U3861 (N_3861,N_246,N_932);
nand U3862 (N_3862,N_831,N_111);
or U3863 (N_3863,N_252,N_1917);
or U3864 (N_3864,N_1417,N_1661);
nor U3865 (N_3865,N_655,N_784);
nand U3866 (N_3866,N_221,N_286);
nor U3867 (N_3867,N_209,N_794);
nor U3868 (N_3868,N_112,N_1846);
and U3869 (N_3869,N_711,N_59);
nand U3870 (N_3870,N_1400,N_1928);
nor U3871 (N_3871,N_1141,N_362);
nor U3872 (N_3872,N_1277,N_111);
nand U3873 (N_3873,N_174,N_761);
nand U3874 (N_3874,N_544,N_1449);
nor U3875 (N_3875,N_963,N_148);
nor U3876 (N_3876,N_1625,N_754);
and U3877 (N_3877,N_520,N_25);
and U3878 (N_3878,N_550,N_1288);
nand U3879 (N_3879,N_714,N_1764);
or U3880 (N_3880,N_1659,N_700);
nand U3881 (N_3881,N_1360,N_671);
and U3882 (N_3882,N_22,N_1175);
and U3883 (N_3883,N_452,N_1738);
nand U3884 (N_3884,N_365,N_481);
nand U3885 (N_3885,N_13,N_101);
nor U3886 (N_3886,N_564,N_659);
nor U3887 (N_3887,N_588,N_755);
and U3888 (N_3888,N_454,N_1592);
nand U3889 (N_3889,N_1704,N_1640);
or U3890 (N_3890,N_804,N_1900);
nor U3891 (N_3891,N_1295,N_124);
and U3892 (N_3892,N_151,N_1067);
or U3893 (N_3893,N_1232,N_840);
and U3894 (N_3894,N_463,N_1967);
nand U3895 (N_3895,N_991,N_224);
and U3896 (N_3896,N_1144,N_160);
nand U3897 (N_3897,N_299,N_266);
and U3898 (N_3898,N_1668,N_347);
nor U3899 (N_3899,N_1909,N_523);
nor U3900 (N_3900,N_1606,N_1123);
nor U3901 (N_3901,N_1958,N_672);
and U3902 (N_3902,N_1465,N_1238);
or U3903 (N_3903,N_866,N_1531);
or U3904 (N_3904,N_27,N_1314);
or U3905 (N_3905,N_1287,N_1498);
or U3906 (N_3906,N_336,N_1800);
or U3907 (N_3907,N_880,N_1860);
nor U3908 (N_3908,N_1853,N_943);
or U3909 (N_3909,N_293,N_1896);
nand U3910 (N_3910,N_1760,N_881);
nand U3911 (N_3911,N_986,N_631);
and U3912 (N_3912,N_473,N_1708);
nand U3913 (N_3913,N_1078,N_271);
nor U3914 (N_3914,N_877,N_1290);
and U3915 (N_3915,N_1656,N_743);
or U3916 (N_3916,N_1264,N_1587);
nor U3917 (N_3917,N_624,N_397);
nand U3918 (N_3918,N_287,N_1827);
or U3919 (N_3919,N_223,N_14);
and U3920 (N_3920,N_1933,N_1905);
nand U3921 (N_3921,N_1795,N_371);
or U3922 (N_3922,N_1726,N_1146);
nand U3923 (N_3923,N_1137,N_1642);
nand U3924 (N_3924,N_373,N_787);
and U3925 (N_3925,N_588,N_934);
nand U3926 (N_3926,N_255,N_1972);
and U3927 (N_3927,N_1085,N_380);
nor U3928 (N_3928,N_396,N_349);
nand U3929 (N_3929,N_1466,N_1317);
xor U3930 (N_3930,N_713,N_1219);
nand U3931 (N_3931,N_917,N_1490);
nor U3932 (N_3932,N_1573,N_338);
xnor U3933 (N_3933,N_556,N_764);
nand U3934 (N_3934,N_126,N_1564);
and U3935 (N_3935,N_1974,N_1130);
nor U3936 (N_3936,N_800,N_1599);
nand U3937 (N_3937,N_1187,N_765);
nor U3938 (N_3938,N_1107,N_1512);
nand U3939 (N_3939,N_334,N_66);
and U3940 (N_3940,N_1545,N_1965);
nor U3941 (N_3941,N_1094,N_1441);
or U3942 (N_3942,N_1451,N_1900);
nand U3943 (N_3943,N_181,N_1313);
nor U3944 (N_3944,N_1024,N_966);
or U3945 (N_3945,N_432,N_1004);
nor U3946 (N_3946,N_1754,N_1470);
or U3947 (N_3947,N_240,N_62);
nand U3948 (N_3948,N_320,N_67);
nor U3949 (N_3949,N_321,N_179);
and U3950 (N_3950,N_909,N_1061);
nand U3951 (N_3951,N_302,N_364);
or U3952 (N_3952,N_523,N_338);
and U3953 (N_3953,N_1062,N_947);
nand U3954 (N_3954,N_1743,N_1842);
and U3955 (N_3955,N_986,N_1303);
xnor U3956 (N_3956,N_1710,N_955);
and U3957 (N_3957,N_854,N_408);
or U3958 (N_3958,N_1865,N_1268);
nor U3959 (N_3959,N_701,N_655);
or U3960 (N_3960,N_10,N_1442);
nand U3961 (N_3961,N_1484,N_1156);
or U3962 (N_3962,N_380,N_912);
nand U3963 (N_3963,N_1778,N_440);
or U3964 (N_3964,N_1267,N_571);
nor U3965 (N_3965,N_1344,N_1934);
or U3966 (N_3966,N_1090,N_891);
or U3967 (N_3967,N_625,N_1543);
nor U3968 (N_3968,N_1842,N_1670);
nand U3969 (N_3969,N_1065,N_246);
and U3970 (N_3970,N_1215,N_1752);
xor U3971 (N_3971,N_845,N_375);
nor U3972 (N_3972,N_288,N_938);
nand U3973 (N_3973,N_1055,N_570);
and U3974 (N_3974,N_1430,N_1030);
nand U3975 (N_3975,N_820,N_629);
nand U3976 (N_3976,N_1800,N_761);
nand U3977 (N_3977,N_233,N_1922);
or U3978 (N_3978,N_1398,N_1204);
nor U3979 (N_3979,N_1965,N_1061);
or U3980 (N_3980,N_453,N_1369);
nand U3981 (N_3981,N_1947,N_640);
and U3982 (N_3982,N_1992,N_1711);
nand U3983 (N_3983,N_1771,N_238);
nand U3984 (N_3984,N_1522,N_576);
nand U3985 (N_3985,N_1647,N_139);
nand U3986 (N_3986,N_607,N_1576);
and U3987 (N_3987,N_1607,N_986);
or U3988 (N_3988,N_463,N_228);
and U3989 (N_3989,N_444,N_248);
or U3990 (N_3990,N_1125,N_1520);
nor U3991 (N_3991,N_1373,N_329);
nand U3992 (N_3992,N_433,N_1667);
and U3993 (N_3993,N_1237,N_154);
nor U3994 (N_3994,N_1242,N_1519);
or U3995 (N_3995,N_900,N_1395);
or U3996 (N_3996,N_1558,N_1597);
nor U3997 (N_3997,N_586,N_984);
nand U3998 (N_3998,N_321,N_1665);
and U3999 (N_3999,N_1745,N_1579);
nor U4000 (N_4000,N_3385,N_2815);
nor U4001 (N_4001,N_3541,N_2335);
nor U4002 (N_4002,N_3967,N_3804);
or U4003 (N_4003,N_3260,N_3783);
nand U4004 (N_4004,N_2210,N_2889);
nand U4005 (N_4005,N_3686,N_3203);
nor U4006 (N_4006,N_2022,N_3728);
nor U4007 (N_4007,N_3162,N_2908);
nor U4008 (N_4008,N_2409,N_3999);
nand U4009 (N_4009,N_3193,N_3188);
nor U4010 (N_4010,N_3475,N_2885);
nor U4011 (N_4011,N_3125,N_3230);
and U4012 (N_4012,N_3298,N_3714);
and U4013 (N_4013,N_2485,N_3735);
and U4014 (N_4014,N_2006,N_3764);
nand U4015 (N_4015,N_3722,N_2924);
nand U4016 (N_4016,N_2611,N_3987);
or U4017 (N_4017,N_2187,N_3587);
or U4018 (N_4018,N_2715,N_2248);
or U4019 (N_4019,N_3430,N_2476);
or U4020 (N_4020,N_2422,N_3194);
or U4021 (N_4021,N_3647,N_3350);
nand U4022 (N_4022,N_3052,N_2141);
or U4023 (N_4023,N_3198,N_2111);
or U4024 (N_4024,N_3152,N_3304);
nor U4025 (N_4025,N_3551,N_2457);
nand U4026 (N_4026,N_3671,N_2710);
and U4027 (N_4027,N_2453,N_2559);
nor U4028 (N_4028,N_2250,N_2847);
or U4029 (N_4029,N_2594,N_3779);
and U4030 (N_4030,N_2202,N_2403);
and U4031 (N_4031,N_2155,N_2145);
or U4032 (N_4032,N_3993,N_3703);
and U4033 (N_4033,N_3894,N_3909);
or U4034 (N_4034,N_2382,N_3892);
nand U4035 (N_4035,N_3536,N_3013);
and U4036 (N_4036,N_3928,N_3268);
or U4037 (N_4037,N_3219,N_3449);
and U4038 (N_4038,N_2685,N_2851);
nor U4039 (N_4039,N_3835,N_3064);
nand U4040 (N_4040,N_3661,N_2993);
and U4041 (N_4041,N_2821,N_2814);
and U4042 (N_4042,N_3994,N_3591);
and U4043 (N_4043,N_2163,N_2305);
and U4044 (N_4044,N_3720,N_3960);
nand U4045 (N_4045,N_3159,N_3971);
nor U4046 (N_4046,N_3858,N_3412);
nor U4047 (N_4047,N_2070,N_3984);
nor U4048 (N_4048,N_2966,N_3086);
nor U4049 (N_4049,N_2200,N_3290);
nor U4050 (N_4050,N_2373,N_3017);
or U4051 (N_4051,N_3269,N_2791);
nand U4052 (N_4052,N_2819,N_2365);
nor U4053 (N_4053,N_3459,N_2771);
nand U4054 (N_4054,N_3090,N_3594);
or U4055 (N_4055,N_3970,N_3483);
nand U4056 (N_4056,N_2096,N_3990);
and U4057 (N_4057,N_2560,N_2109);
nor U4058 (N_4058,N_3905,N_3254);
or U4059 (N_4059,N_2033,N_3733);
and U4060 (N_4060,N_2462,N_3698);
and U4061 (N_4061,N_2002,N_2666);
nor U4062 (N_4062,N_3539,N_3983);
nor U4063 (N_4063,N_3360,N_2190);
and U4064 (N_4064,N_2739,N_2029);
and U4065 (N_4065,N_2314,N_3362);
and U4066 (N_4066,N_3220,N_2989);
or U4067 (N_4067,N_3570,N_3942);
or U4068 (N_4068,N_3514,N_2215);
nand U4069 (N_4069,N_3370,N_2824);
nor U4070 (N_4070,N_2711,N_3511);
and U4071 (N_4071,N_2927,N_2933);
and U4072 (N_4072,N_2510,N_2825);
nor U4073 (N_4073,N_2579,N_3618);
nand U4074 (N_4074,N_3453,N_2923);
nor U4075 (N_4075,N_2965,N_3561);
or U4076 (N_4076,N_3082,N_3129);
or U4077 (N_4077,N_3431,N_2631);
or U4078 (N_4078,N_2508,N_2533);
and U4079 (N_4079,N_2165,N_2073);
nor U4080 (N_4080,N_3363,N_2001);
and U4081 (N_4081,N_2188,N_2865);
or U4082 (N_4082,N_2057,N_2333);
or U4083 (N_4083,N_2385,N_2737);
nand U4084 (N_4084,N_2998,N_2479);
and U4085 (N_4085,N_2468,N_3712);
xnor U4086 (N_4086,N_2375,N_2044);
nand U4087 (N_4087,N_3955,N_3436);
nor U4088 (N_4088,N_3098,N_3816);
or U4089 (N_4089,N_3284,N_3118);
or U4090 (N_4090,N_3818,N_3359);
and U4091 (N_4091,N_2366,N_3390);
nor U4092 (N_4092,N_3989,N_2123);
and U4093 (N_4093,N_2499,N_2871);
and U4094 (N_4094,N_2266,N_3531);
nor U4095 (N_4095,N_2629,N_3935);
nor U4096 (N_4096,N_3176,N_2331);
or U4097 (N_4097,N_2224,N_3902);
and U4098 (N_4098,N_2034,N_3228);
nand U4099 (N_4099,N_3919,N_2676);
nand U4100 (N_4100,N_3236,N_2026);
nor U4101 (N_4101,N_3426,N_3206);
or U4102 (N_4102,N_2590,N_2564);
or U4103 (N_4103,N_2869,N_3336);
or U4104 (N_4104,N_2370,N_2286);
and U4105 (N_4105,N_3883,N_3774);
or U4106 (N_4106,N_3624,N_2838);
nand U4107 (N_4107,N_3001,N_2613);
and U4108 (N_4108,N_3634,N_3307);
and U4109 (N_4109,N_2903,N_2780);
or U4110 (N_4110,N_3031,N_2856);
and U4111 (N_4111,N_3903,N_2696);
nand U4112 (N_4112,N_2291,N_3326);
nand U4113 (N_4113,N_3223,N_3553);
nor U4114 (N_4114,N_2405,N_2466);
and U4115 (N_4115,N_2374,N_3628);
xor U4116 (N_4116,N_3180,N_2731);
and U4117 (N_4117,N_3812,N_3866);
or U4118 (N_4118,N_2263,N_3943);
nand U4119 (N_4119,N_2999,N_2521);
and U4120 (N_4120,N_3213,N_2035);
and U4121 (N_4121,N_3339,N_3301);
or U4122 (N_4122,N_3857,N_3771);
and U4123 (N_4123,N_2194,N_2108);
and U4124 (N_4124,N_3292,N_2164);
or U4125 (N_4125,N_2640,N_2706);
nor U4126 (N_4126,N_2239,N_3755);
nand U4127 (N_4127,N_2399,N_2496);
or U4128 (N_4128,N_2955,N_3470);
and U4129 (N_4129,N_3043,N_3906);
and U4130 (N_4130,N_2032,N_3968);
nand U4131 (N_4131,N_3007,N_2555);
nand U4132 (N_4132,N_2960,N_2284);
or U4133 (N_4133,N_3338,N_2772);
and U4134 (N_4134,N_2605,N_2980);
nor U4135 (N_4135,N_2655,N_3309);
nor U4136 (N_4136,N_3524,N_2487);
nand U4137 (N_4137,N_3966,N_3973);
and U4138 (N_4138,N_2297,N_2943);
nand U4139 (N_4139,N_2671,N_2099);
nor U4140 (N_4140,N_3833,N_2475);
nand U4141 (N_4141,N_2642,N_2738);
and U4142 (N_4142,N_3543,N_2336);
or U4143 (N_4143,N_2502,N_2665);
or U4144 (N_4144,N_3873,N_2151);
nand U4145 (N_4145,N_3956,N_3692);
nand U4146 (N_4146,N_3654,N_3663);
nand U4147 (N_4147,N_2622,N_2095);
nor U4148 (N_4148,N_3940,N_2830);
or U4149 (N_4149,N_3177,N_3952);
nand U4150 (N_4150,N_3060,N_3274);
or U4151 (N_4151,N_3695,N_2883);
nor U4152 (N_4152,N_3854,N_2222);
and U4153 (N_4153,N_2074,N_3044);
nand U4154 (N_4154,N_2818,N_2509);
or U4155 (N_4155,N_3104,N_3155);
or U4156 (N_4156,N_2065,N_3329);
and U4157 (N_4157,N_3235,N_2736);
nor U4158 (N_4158,N_2437,N_2808);
and U4159 (N_4159,N_2971,N_3716);
nor U4160 (N_4160,N_3102,N_2803);
nand U4161 (N_4161,N_3679,N_2234);
or U4162 (N_4162,N_3314,N_2486);
nand U4163 (N_4163,N_3502,N_2441);
or U4164 (N_4164,N_3417,N_3391);
and U4165 (N_4165,N_2528,N_3185);
or U4166 (N_4166,N_3912,N_2567);
nand U4167 (N_4167,N_3322,N_2352);
or U4168 (N_4168,N_2388,N_3070);
nand U4169 (N_4169,N_3766,N_2969);
and U4170 (N_4170,N_2673,N_2784);
xor U4171 (N_4171,N_3374,N_3335);
nor U4172 (N_4172,N_3782,N_2782);
or U4173 (N_4173,N_3174,N_2678);
and U4174 (N_4174,N_2831,N_3058);
and U4175 (N_4175,N_2727,N_3564);
nor U4176 (N_4176,N_3798,N_3303);
and U4177 (N_4177,N_3160,N_3781);
nor U4178 (N_4178,N_3710,N_2191);
nor U4179 (N_4179,N_3035,N_2970);
and U4180 (N_4180,N_2227,N_2419);
or U4181 (N_4181,N_2037,N_2454);
and U4182 (N_4182,N_3724,N_3186);
or U4183 (N_4183,N_2277,N_3075);
and U4184 (N_4184,N_2907,N_3709);
nand U4185 (N_4185,N_2758,N_2828);
and U4186 (N_4186,N_3232,N_2843);
or U4187 (N_4187,N_2411,N_2730);
xnor U4188 (N_4188,N_2635,N_3879);
or U4189 (N_4189,N_3595,N_2931);
nand U4190 (N_4190,N_3183,N_2338);
and U4191 (N_4191,N_2554,N_3584);
and U4192 (N_4192,N_3821,N_2058);
nor U4193 (N_4193,N_3582,N_3773);
nand U4194 (N_4194,N_2645,N_3667);
and U4195 (N_4195,N_3615,N_3776);
and U4196 (N_4196,N_3717,N_2625);
nand U4197 (N_4197,N_3910,N_2773);
nand U4198 (N_4198,N_2376,N_2060);
and U4199 (N_4199,N_3738,N_3754);
or U4200 (N_4200,N_2805,N_3132);
and U4201 (N_4201,N_2361,N_3355);
or U4202 (N_4202,N_3332,N_2093);
and U4203 (N_4203,N_2402,N_2106);
nor U4204 (N_4204,N_3196,N_2763);
nand U4205 (N_4205,N_2523,N_2469);
and U4206 (N_4206,N_2174,N_3830);
or U4207 (N_4207,N_2588,N_3736);
nand U4208 (N_4208,N_2862,N_3337);
and U4209 (N_4209,N_3827,N_3682);
or U4210 (N_4210,N_3440,N_3522);
and U4211 (N_4211,N_3218,N_2514);
nand U4212 (N_4212,N_3424,N_3158);
or U4213 (N_4213,N_2801,N_2294);
nor U4214 (N_4214,N_2327,N_3597);
nor U4215 (N_4215,N_3382,N_3500);
nand U4216 (N_4216,N_2343,N_3498);
or U4217 (N_4217,N_3049,N_3974);
or U4218 (N_4218,N_2104,N_3255);
and U4219 (N_4219,N_3101,N_2094);
xor U4220 (N_4220,N_3383,N_3611);
nor U4221 (N_4221,N_3165,N_2794);
or U4222 (N_4222,N_3538,N_2707);
nand U4223 (N_4223,N_3747,N_3884);
and U4224 (N_4224,N_3042,N_2332);
nor U4225 (N_4225,N_2986,N_2247);
and U4226 (N_4226,N_2872,N_2085);
and U4227 (N_4227,N_3084,N_2348);
and U4228 (N_4228,N_3111,N_2130);
and U4229 (N_4229,N_3120,N_2648);
xor U4230 (N_4230,N_3146,N_3019);
or U4231 (N_4231,N_3923,N_3533);
and U4232 (N_4232,N_3809,N_2015);
nor U4233 (N_4233,N_2786,N_2922);
or U4234 (N_4234,N_2604,N_3088);
and U4235 (N_4235,N_3109,N_2283);
nor U4236 (N_4236,N_2860,N_2792);
and U4237 (N_4237,N_2593,N_2765);
and U4238 (N_4238,N_3458,N_3216);
nand U4239 (N_4239,N_3068,N_2627);
nor U4240 (N_4240,N_3488,N_2734);
nand U4241 (N_4241,N_3026,N_3113);
nor U4242 (N_4242,N_2072,N_2692);
and U4243 (N_4243,N_3127,N_3652);
and U4244 (N_4244,N_2699,N_3881);
or U4245 (N_4245,N_2062,N_3550);
nand U4246 (N_4246,N_2974,N_2483);
or U4247 (N_4247,N_3921,N_2039);
or U4248 (N_4248,N_2020,N_3768);
and U4249 (N_4249,N_2281,N_2303);
or U4250 (N_4250,N_3843,N_2103);
nand U4251 (N_4251,N_3168,N_2116);
and U4252 (N_4252,N_2480,N_2478);
nor U4253 (N_4253,N_2396,N_3893);
nand U4254 (N_4254,N_3794,N_3876);
nand U4255 (N_4255,N_3321,N_2682);
nand U4256 (N_4256,N_3706,N_2578);
or U4257 (N_4257,N_2204,N_2649);
nor U4258 (N_4258,N_3263,N_2054);
xor U4259 (N_4259,N_2539,N_2262);
and U4260 (N_4260,N_2958,N_2557);
nor U4261 (N_4261,N_2364,N_2901);
and U4262 (N_4262,N_3108,N_3758);
and U4263 (N_4263,N_2290,N_3869);
and U4264 (N_4264,N_2313,N_2356);
nand U4265 (N_4265,N_2008,N_3778);
xnor U4266 (N_4266,N_2158,N_3140);
and U4267 (N_4267,N_2232,N_3369);
nand U4268 (N_4268,N_2410,N_3191);
nand U4269 (N_4269,N_3750,N_2688);
nand U4270 (N_4270,N_2205,N_3405);
nor U4271 (N_4271,N_2017,N_3341);
and U4272 (N_4272,N_2119,N_2280);
xor U4273 (N_4273,N_3559,N_2064);
and U4274 (N_4274,N_3046,N_2684);
nor U4275 (N_4275,N_2630,N_3549);
nor U4276 (N_4276,N_2850,N_3691);
nand U4277 (N_4277,N_2372,N_3051);
nor U4278 (N_4278,N_3091,N_2783);
or U4279 (N_4279,N_3266,N_3985);
nor U4280 (N_4280,N_2185,N_2620);
nor U4281 (N_4281,N_3081,N_2747);
xor U4282 (N_4282,N_3788,N_2906);
or U4283 (N_4283,N_2669,N_2392);
or U4284 (N_4284,N_2249,N_2458);
or U4285 (N_4285,N_2324,N_3351);
or U4286 (N_4286,N_3563,N_2681);
or U4287 (N_4287,N_2051,N_3422);
nand U4288 (N_4288,N_2025,N_2701);
nand U4289 (N_4289,N_2724,N_3711);
nand U4290 (N_4290,N_3354,N_3664);
nand U4291 (N_4291,N_2391,N_2694);
nor U4292 (N_4292,N_2349,N_3689);
or U4293 (N_4293,N_3889,N_3586);
nand U4294 (N_4294,N_3285,N_3838);
and U4295 (N_4295,N_3775,N_3650);
and U4296 (N_4296,N_2873,N_3271);
and U4297 (N_4297,N_3767,N_2654);
nor U4298 (N_4298,N_3904,N_3143);
or U4299 (N_4299,N_3721,N_2769);
or U4300 (N_4300,N_2552,N_3467);
nor U4301 (N_4301,N_3100,N_2316);
or U4302 (N_4302,N_2144,N_2602);
nor U4303 (N_4303,N_3694,N_2414);
or U4304 (N_4304,N_2870,N_3862);
nand U4305 (N_4305,N_2122,N_2518);
and U4306 (N_4306,N_3006,N_3518);
and U4307 (N_4307,N_2279,N_3085);
nand U4308 (N_4308,N_3130,N_3197);
xor U4309 (N_4309,N_3240,N_3673);
nor U4310 (N_4310,N_2633,N_2686);
nor U4311 (N_4311,N_3908,N_3872);
and U4312 (N_4312,N_2914,N_3455);
nor U4313 (N_4313,N_2482,N_2050);
or U4314 (N_4314,N_3525,N_2031);
nor U4315 (N_4315,N_3510,N_2964);
nand U4316 (N_4316,N_3425,N_2426);
and U4317 (N_4317,N_3267,N_3485);
nor U4318 (N_4318,N_2810,N_3115);
nor U4319 (N_4319,N_3464,N_2255);
and U4320 (N_4320,N_2695,N_3361);
nor U4321 (N_4321,N_2363,N_3151);
nor U4322 (N_4322,N_3730,N_3402);
nor U4323 (N_4323,N_3953,N_3420);
and U4324 (N_4324,N_2340,N_3708);
nor U4325 (N_4325,N_2131,N_3701);
and U4326 (N_4326,N_2726,N_2162);
nand U4327 (N_4327,N_3173,N_2059);
or U4328 (N_4328,N_3713,N_3726);
nor U4329 (N_4329,N_2206,N_3373);
nand U4330 (N_4330,N_2646,N_2369);
and U4331 (N_4331,N_2735,N_3039);
and U4332 (N_4332,N_3045,N_3117);
nor U4333 (N_4333,N_2744,N_2799);
nand U4334 (N_4334,N_2916,N_3528);
nand U4335 (N_4335,N_3947,N_2325);
nor U4336 (N_4336,N_2498,N_2941);
or U4337 (N_4337,N_3787,N_3157);
and U4338 (N_4338,N_3831,N_3150);
nand U4339 (N_4339,N_3975,N_2504);
and U4340 (N_4340,N_3318,N_3010);
nor U4341 (N_4341,N_2817,N_2473);
nand U4342 (N_4342,N_3477,N_2957);
and U4343 (N_4343,N_3327,N_2788);
or U4344 (N_4344,N_3937,N_3154);
nor U4345 (N_4345,N_3471,N_3565);
or U4346 (N_4346,N_2570,N_2910);
nand U4347 (N_4347,N_3763,N_2027);
nand U4348 (N_4348,N_3080,N_2987);
or U4349 (N_4349,N_2056,N_2619);
nand U4350 (N_4350,N_3796,N_2456);
nand U4351 (N_4351,N_3258,N_2751);
nor U4352 (N_4352,N_2705,N_3891);
and U4353 (N_4353,N_2952,N_2220);
or U4354 (N_4354,N_2143,N_2770);
nand U4355 (N_4355,N_2544,N_2086);
nor U4356 (N_4356,N_2595,N_2028);
and U4357 (N_4357,N_3317,N_2089);
nor U4358 (N_4358,N_2585,N_3495);
nor U4359 (N_4359,N_3486,N_2767);
and U4360 (N_4360,N_3447,N_2354);
and U4361 (N_4361,N_2192,N_2530);
nor U4362 (N_4362,N_2937,N_2946);
and U4363 (N_4363,N_3599,N_3182);
nor U4364 (N_4364,N_3861,N_2992);
or U4365 (N_4365,N_2083,N_3573);
and U4366 (N_4366,N_3614,N_2413);
nand U4367 (N_4367,N_2603,N_2785);
nand U4368 (N_4368,N_3604,N_2836);
nand U4369 (N_4369,N_3334,N_2079);
nor U4370 (N_4370,N_2230,N_3110);
or U4371 (N_4371,N_3503,N_2729);
nor U4372 (N_4372,N_2047,N_3256);
or U4373 (N_4373,N_3548,N_3875);
or U4374 (N_4374,N_3959,N_2442);
nand U4375 (N_4375,N_3655,N_2218);
or U4376 (N_4376,N_3294,N_3037);
nor U4377 (N_4377,N_3592,N_3069);
nand U4378 (N_4378,N_3209,N_2626);
and U4379 (N_4379,N_3920,N_2421);
and U4380 (N_4380,N_3946,N_3609);
nor U4381 (N_4381,N_3590,N_2121);
or U4382 (N_4382,N_2347,N_3397);
and U4383 (N_4383,N_3023,N_2844);
and U4384 (N_4384,N_3642,N_3576);
nand U4385 (N_4385,N_2975,N_3452);
and U4386 (N_4386,N_3786,N_2556);
and U4387 (N_4387,N_3648,N_2193);
or U4388 (N_4388,N_2754,N_3596);
and U4389 (N_4389,N_3015,N_3684);
nand U4390 (N_4390,N_2489,N_3676);
nor U4391 (N_4391,N_3653,N_3179);
and U4392 (N_4392,N_3311,N_2935);
or U4393 (N_4393,N_2319,N_2076);
nor U4394 (N_4394,N_3333,N_3171);
nor U4395 (N_4395,N_3319,N_2996);
nor U4396 (N_4396,N_3980,N_2139);
nand U4397 (N_4397,N_2634,N_3008);
or U4398 (N_4398,N_3633,N_3434);
nand U4399 (N_4399,N_2494,N_3742);
nand U4400 (N_4400,N_3372,N_2092);
nor U4401 (N_4401,N_3867,N_2078);
nand U4402 (N_4402,N_3546,N_2928);
and U4403 (N_4403,N_2542,N_3612);
nand U4404 (N_4404,N_3096,N_3649);
nor U4405 (N_4405,N_3242,N_3808);
nor U4406 (N_4406,N_3446,N_2126);
and U4407 (N_4407,N_2124,N_2623);
nor U4408 (N_4408,N_2238,N_2439);
or U4409 (N_4409,N_2691,N_3913);
nor U4410 (N_4410,N_3041,N_2282);
nand U4411 (N_4411,N_2713,N_2149);
or U4412 (N_4412,N_2849,N_2826);
or U4413 (N_4413,N_3670,N_3674);
nand U4414 (N_4414,N_2425,N_3797);
nor U4415 (N_4415,N_3344,N_3253);
nor U4416 (N_4416,N_3662,N_2837);
or U4417 (N_4417,N_2863,N_2795);
nor U4418 (N_4418,N_2379,N_2904);
or U4419 (N_4419,N_3247,N_3442);
nand U4420 (N_4420,N_3958,N_2460);
nand U4421 (N_4421,N_2179,N_3126);
and U4422 (N_4422,N_2875,N_3448);
nor U4423 (N_4423,N_2512,N_2806);
or U4424 (N_4424,N_2972,N_3700);
nand U4425 (N_4425,N_3375,N_2477);
or U4426 (N_4426,N_3419,N_2199);
or U4427 (N_4427,N_2068,N_2446);
or U4428 (N_4428,N_2293,N_3342);
and U4429 (N_4429,N_2156,N_2175);
or U4430 (N_4430,N_3018,N_3976);
or U4431 (N_4431,N_2697,N_3400);
or U4432 (N_4432,N_2178,N_2979);
or U4433 (N_4433,N_3699,N_2451);
or U4434 (N_4434,N_3462,N_3312);
nor U4435 (N_4435,N_3169,N_2326);
nand U4436 (N_4436,N_3749,N_2398);
nor U4437 (N_4437,N_2142,N_2265);
nand U4438 (N_4438,N_2323,N_3792);
nor U4439 (N_4439,N_2624,N_2617);
and U4440 (N_4440,N_2071,N_3600);
nor U4441 (N_4441,N_3626,N_3687);
and U4442 (N_4442,N_3261,N_2168);
or U4443 (N_4443,N_2353,N_3469);
nand U4444 (N_4444,N_2687,N_2540);
nor U4445 (N_4445,N_2471,N_3443);
and U4446 (N_4446,N_2522,N_2704);
or U4447 (N_4447,N_2896,N_3033);
and U4448 (N_4448,N_3793,N_3895);
xor U4449 (N_4449,N_3074,N_3265);
nand U4450 (N_4450,N_2030,N_2968);
or U4451 (N_4451,N_3392,N_2947);
nand U4452 (N_4452,N_2147,N_3588);
nand U4453 (N_4453,N_2113,N_3629);
and U4454 (N_4454,N_2925,N_2926);
nor U4455 (N_4455,N_3142,N_3799);
nor U4456 (N_4456,N_2052,N_3731);
or U4457 (N_4457,N_3660,N_3380);
and U4458 (N_4458,N_2587,N_2644);
nor U4459 (N_4459,N_2527,N_2661);
nand U4460 (N_4460,N_3316,N_2535);
and U4461 (N_4461,N_3320,N_3535);
or U4462 (N_4462,N_2445,N_3746);
and U4463 (N_4463,N_3190,N_3501);
or U4464 (N_4464,N_2725,N_2488);
and U4465 (N_4465,N_2606,N_2018);
nor U4466 (N_4466,N_2983,N_2362);
nand U4467 (N_4467,N_2420,N_2911);
and U4468 (N_4468,N_3523,N_2455);
nor U4469 (N_4469,N_2228,N_2082);
and U4470 (N_4470,N_3677,N_2913);
or U4471 (N_4471,N_2448,N_2272);
xor U4472 (N_4472,N_2990,N_3529);
or U4473 (N_4473,N_2917,N_3249);
and U4474 (N_4474,N_2967,N_2643);
nand U4475 (N_4475,N_2720,N_3364);
and U4476 (N_4476,N_2306,N_2041);
nand U4477 (N_4477,N_3246,N_2534);
nand U4478 (N_4478,N_3534,N_2915);
nor U4479 (N_4479,N_2670,N_3264);
nor U4480 (N_4480,N_3050,N_2137);
nor U4481 (N_4481,N_3991,N_3437);
and U4482 (N_4482,N_2097,N_2524);
nand U4483 (N_4483,N_3852,N_3558);
nand U4484 (N_4484,N_3393,N_2171);
or U4485 (N_4485,N_2401,N_2884);
and U4486 (N_4486,N_3878,N_3156);
nor U4487 (N_4487,N_2921,N_2939);
nand U4488 (N_4488,N_2236,N_2895);
nor U4489 (N_4489,N_3083,N_2301);
nor U4490 (N_4490,N_2797,N_2355);
nand U4491 (N_4491,N_2621,N_2219);
or U4492 (N_4492,N_3489,N_2812);
and U4493 (N_4493,N_2507,N_2214);
or U4494 (N_4494,N_2444,N_3103);
or U4495 (N_4495,N_2351,N_2383);
or U4496 (N_4496,N_2173,N_3308);
nand U4497 (N_4497,N_3574,N_3805);
and U4498 (N_4498,N_2598,N_2016);
nand U4499 (N_4499,N_3250,N_3651);
and U4500 (N_4500,N_3791,N_3438);
nor U4501 (N_4501,N_3961,N_2450);
nor U4502 (N_4502,N_3814,N_2984);
nor U4503 (N_4503,N_3868,N_3067);
nand U4504 (N_4504,N_3887,N_2107);
nor U4505 (N_4505,N_3856,N_3640);
and U4506 (N_4506,N_2288,N_3832);
nand U4507 (N_4507,N_2386,N_2212);
and U4508 (N_4508,N_3890,N_3252);
and U4509 (N_4509,N_3986,N_3610);
nand U4510 (N_4510,N_3461,N_2994);
or U4511 (N_4511,N_3021,N_3938);
or U4512 (N_4512,N_2289,N_3916);
nor U4513 (N_4513,N_2599,N_2547);
nand U4514 (N_4514,N_3849,N_3825);
or U4515 (N_4515,N_2934,N_2668);
or U4516 (N_4516,N_2615,N_2612);
nor U4517 (N_4517,N_3520,N_3071);
or U4518 (N_4518,N_2345,N_3617);
nand U4519 (N_4519,N_2418,N_2584);
or U4520 (N_4520,N_2246,N_2600);
or U4521 (N_4521,N_3352,N_2525);
or U4522 (N_4522,N_3657,N_2577);
nand U4523 (N_4523,N_2894,N_3855);
nor U4524 (N_4524,N_2723,N_3537);
nor U4525 (N_4525,N_3589,N_3433);
and U4526 (N_4526,N_2607,N_2464);
or U4527 (N_4527,N_2395,N_3944);
nand U4528 (N_4528,N_2991,N_2430);
and U4529 (N_4529,N_2647,N_2846);
and U4530 (N_4530,N_2197,N_2069);
nor U4531 (N_4531,N_2492,N_2427);
and U4532 (N_4532,N_2519,N_3480);
nand U4533 (N_4533,N_3519,N_3998);
or U4534 (N_4534,N_3262,N_3208);
or U4535 (N_4535,N_2253,N_2732);
or U4536 (N_4536,N_3214,N_2912);
nand U4537 (N_4537,N_3291,N_2461);
and U4538 (N_4538,N_2436,N_3065);
nand U4539 (N_4539,N_3801,N_3493);
and U4540 (N_4540,N_2330,N_2302);
or U4541 (N_4541,N_2133,N_3388);
and U4542 (N_4542,N_2861,N_2679);
and U4543 (N_4543,N_2452,N_3607);
or U4544 (N_4544,N_3226,N_2787);
or U4545 (N_4545,N_3672,N_2066);
or U4546 (N_4546,N_3598,N_2742);
nand U4547 (N_4547,N_2154,N_3411);
or U4548 (N_4548,N_3325,N_2435);
nand U4549 (N_4549,N_3406,N_3515);
nor U4550 (N_4550,N_2537,N_2745);
nand U4551 (N_4551,N_3384,N_3231);
or U4552 (N_4552,N_2244,N_2148);
and U4553 (N_4553,N_2371,N_3259);
nor U4554 (N_4554,N_3079,N_2024);
and U4555 (N_4555,N_3073,N_3439);
and U4556 (N_4556,N_3167,N_2878);
nand U4557 (N_4557,N_3739,N_3931);
or U4558 (N_4558,N_3000,N_2759);
nor U4559 (N_4559,N_3136,N_3295);
or U4560 (N_4560,N_3072,N_2802);
and U4561 (N_4561,N_2346,N_3769);
and U4562 (N_4562,N_3105,N_2406);
or U4563 (N_4563,N_2905,N_2043);
or U4564 (N_4564,N_2274,N_3358);
nand U4565 (N_4565,N_3207,N_2254);
nor U4566 (N_4566,N_3988,N_2198);
and U4567 (N_4567,N_3847,N_3340);
xor U4568 (N_4568,N_2942,N_3497);
nor U4569 (N_4569,N_2760,N_2881);
or U4570 (N_4570,N_3435,N_2309);
nand U4571 (N_4571,N_2639,N_2918);
or U4572 (N_4572,N_3837,N_2513);
nor U4573 (N_4573,N_3727,N_3820);
and U4574 (N_4574,N_3668,N_2474);
or U4575 (N_4575,N_2463,N_3807);
nand U4576 (N_4576,N_3560,N_3950);
or U4577 (N_4577,N_3737,N_3760);
or U4578 (N_4578,N_3450,N_3800);
nor U4579 (N_4579,N_2201,N_3119);
and U4580 (N_4580,N_3225,N_3934);
or U4581 (N_4581,N_2891,N_2848);
and U4582 (N_4582,N_3819,N_3472);
or U4583 (N_4583,N_2258,N_3283);
or U4584 (N_4584,N_2211,N_3897);
or U4585 (N_4585,N_2310,N_3665);
and U4586 (N_4586,N_2161,N_3398);
or U4587 (N_4587,N_3927,N_2189);
or U4588 (N_4588,N_3428,N_2813);
nand U4589 (N_4589,N_3211,N_3785);
nor U4590 (N_4590,N_3696,N_3885);
and U4591 (N_4591,N_2235,N_3865);
nor U4592 (N_4592,N_2636,N_2733);
nand U4593 (N_4593,N_3656,N_3659);
nor U4594 (N_4594,N_3145,N_3941);
or U4595 (N_4595,N_2134,N_3978);
or U4596 (N_4596,N_2115,N_2674);
nor U4597 (N_4597,N_2260,N_2412);
and U4598 (N_4598,N_3077,N_2841);
nand U4599 (N_4599,N_2378,N_2750);
and U4600 (N_4600,N_2882,N_2546);
and U4601 (N_4601,N_2013,N_2500);
nand U4602 (N_4602,N_2221,N_3772);
nand U4603 (N_4603,N_3099,N_2764);
nor U4604 (N_4604,N_2601,N_2459);
nand U4605 (N_4605,N_2261,N_2664);
or U4606 (N_4606,N_2110,N_2888);
nor U4607 (N_4607,N_2334,N_2663);
nor U4608 (N_4608,N_3245,N_3874);
xnor U4609 (N_4609,N_3053,N_3466);
nand U4610 (N_4610,N_2075,N_2088);
nand U4611 (N_4611,N_3882,N_3569);
nand U4612 (N_4612,N_2000,N_3756);
nand U4613 (N_4613,N_2811,N_2529);
nand U4614 (N_4614,N_3557,N_2899);
nand U4615 (N_4615,N_3568,N_2367);
nand U4616 (N_4616,N_3745,N_2793);
nand U4617 (N_4617,N_2798,N_3513);
nor U4618 (N_4618,N_3841,N_3925);
or U4619 (N_4619,N_2098,N_2589);
and U4620 (N_4620,N_3637,N_3257);
nand U4621 (N_4621,N_2576,N_3556);
nor U4622 (N_4622,N_2768,N_2118);
nand U4623 (N_4623,N_3829,N_3404);
nor U4624 (N_4624,N_3826,N_3957);
and U4625 (N_4625,N_2938,N_3378);
and U4626 (N_4626,N_2879,N_3636);
nor U4627 (N_4627,N_3124,N_3484);
nand U4628 (N_4628,N_2781,N_2565);
and U4629 (N_4629,N_3123,N_3022);
or U4630 (N_4630,N_3817,N_2857);
and U4631 (N_4631,N_2011,N_2890);
nand U4632 (N_4632,N_3996,N_2112);
or U4633 (N_4633,N_3898,N_2827);
or U4634 (N_4634,N_2003,N_2287);
and U4635 (N_4635,N_3057,N_3945);
nand U4636 (N_4636,N_3273,N_2186);
or U4637 (N_4637,N_2558,N_2761);
nor U4638 (N_4638,N_3850,N_2709);
and U4639 (N_4639,N_3572,N_2491);
nand U4640 (N_4640,N_3296,N_3705);
nand U4641 (N_4641,N_3227,N_3575);
nand U4642 (N_4642,N_2566,N_2055);
nand U4643 (N_4643,N_2160,N_3396);
nand U4644 (N_4644,N_2536,N_3287);
nor U4645 (N_4645,N_3566,N_3842);
nor U4646 (N_4646,N_2299,N_2359);
and U4647 (N_4647,N_3963,N_3248);
nand U4648 (N_4648,N_3929,N_3087);
or U4649 (N_4649,N_3202,N_2423);
or U4650 (N_4650,N_2583,N_2835);
nand U4651 (N_4651,N_3040,N_3187);
nor U4652 (N_4652,N_3016,N_3602);
and U4653 (N_4653,N_2381,N_3277);
and U4654 (N_4654,N_3144,N_2693);
or U4655 (N_4655,N_3275,N_3137);
and U4656 (N_4656,N_2776,N_3540);
nand U4657 (N_4657,N_3416,N_2752);
nand U4658 (N_4658,N_3324,N_3544);
and U4659 (N_4659,N_2961,N_2779);
nand U4660 (N_4660,N_3859,N_2019);
nand U4661 (N_4661,N_3784,N_3593);
and U4662 (N_4662,N_3504,N_3606);
nand U4663 (N_4663,N_2384,N_2120);
nand U4664 (N_4664,N_3147,N_3752);
nor U4665 (N_4665,N_2874,N_3639);
nor U4666 (N_4666,N_2434,N_3106);
nand U4667 (N_4667,N_3962,N_3719);
nor U4668 (N_4668,N_3122,N_3715);
and U4669 (N_4669,N_3394,N_2241);
nor U4670 (N_4670,N_3297,N_3478);
nor U4671 (N_4671,N_2948,N_2440);
nor U4672 (N_4672,N_2628,N_3795);
nand U4673 (N_4673,N_3401,N_2067);
or U4674 (N_4674,N_2650,N_3482);
nor U4675 (N_4675,N_3770,N_2569);
nor U4676 (N_4676,N_3761,N_2177);
nor U4677 (N_4677,N_3844,N_2839);
and U4678 (N_4678,N_3494,N_2641);
or U4679 (N_4679,N_3054,N_3305);
and U4680 (N_4680,N_3181,N_2080);
and U4681 (N_4681,N_2531,N_2859);
or U4682 (N_4682,N_3474,N_2503);
or U4683 (N_4683,N_3062,N_3846);
nand U4684 (N_4684,N_3930,N_2484);
nor U4685 (N_4685,N_3680,N_2574);
nand U4686 (N_4686,N_2614,N_2823);
or U4687 (N_4687,N_3951,N_3212);
and U4688 (N_4688,N_3896,N_2892);
or U4689 (N_4689,N_3444,N_2978);
nand U4690 (N_4690,N_2501,N_2703);
or U4691 (N_4691,N_2140,N_3577);
or U4692 (N_4692,N_2900,N_2582);
or U4693 (N_4693,N_2256,N_2358);
nand U4694 (N_4694,N_3379,N_2315);
nand U4695 (N_4695,N_2495,N_3097);
nand U4696 (N_4696,N_2545,N_3315);
or U4697 (N_4697,N_3408,N_3166);
nand U4698 (N_4698,N_2944,N_3056);
nor U4699 (N_4699,N_2181,N_2897);
or U4700 (N_4700,N_3302,N_2114);
nor U4701 (N_4701,N_2909,N_3454);
and U4702 (N_4702,N_2962,N_3407);
or U4703 (N_4703,N_3251,N_2716);
nor U4704 (N_4704,N_2307,N_2740);
nand U4705 (N_4705,N_3585,N_2563);
or U4706 (N_4706,N_2864,N_3900);
and U4707 (N_4707,N_2743,N_3418);
nand U4708 (N_4708,N_2311,N_2796);
and U4709 (N_4709,N_2719,N_3977);
and U4710 (N_4710,N_2497,N_2789);
or U4711 (N_4711,N_2610,N_3580);
or U4712 (N_4712,N_2063,N_2728);
or U4713 (N_4713,N_2428,N_3063);
nor U4714 (N_4714,N_2341,N_2756);
or U4715 (N_4715,N_2950,N_3744);
or U4716 (N_4716,N_3005,N_3395);
nor U4717 (N_4717,N_2775,N_2213);
or U4718 (N_4718,N_2700,N_3204);
nor U4719 (N_4719,N_3289,N_3221);
nand U4720 (N_4720,N_3748,N_2273);
or U4721 (N_4721,N_3627,N_2209);
nor U4722 (N_4722,N_2893,N_2562);
nand U4723 (N_4723,N_2973,N_2505);
nand U4724 (N_4724,N_2397,N_3555);
and U4725 (N_4725,N_2132,N_3845);
and U4726 (N_4726,N_3014,N_3205);
and U4727 (N_4727,N_3034,N_2251);
or U4728 (N_4728,N_2138,N_2902);
nand U4729 (N_4729,N_3270,N_2226);
or U4730 (N_4730,N_3377,N_3389);
and U4731 (N_4731,N_3293,N_3463);
nor U4732 (N_4732,N_2976,N_2573);
and U4733 (N_4733,N_3527,N_2853);
or U4734 (N_4734,N_2511,N_3836);
nor U4735 (N_4735,N_2651,N_2616);
nand U4736 (N_4736,N_3004,N_3490);
nor U4737 (N_4737,N_2102,N_2159);
and U4738 (N_4738,N_3762,N_3516);
or U4739 (N_4739,N_3547,N_3840);
and U4740 (N_4740,N_2240,N_3815);
or U4741 (N_4741,N_3765,N_2465);
nor U4742 (N_4742,N_2829,N_3545);
or U4743 (N_4743,N_2766,N_3032);
and U4744 (N_4744,N_2959,N_3693);
or U4745 (N_4745,N_3028,N_3286);
nor U4746 (N_4746,N_2653,N_2312);
or U4747 (N_4747,N_2252,N_2081);
nand U4748 (N_4748,N_2541,N_3282);
nand U4749 (N_4749,N_2127,N_3581);
nand U4750 (N_4750,N_3571,N_2919);
nor U4751 (N_4751,N_2166,N_3201);
and U4752 (N_4752,N_3310,N_3457);
nand U4753 (N_4753,N_2045,N_2840);
and U4754 (N_4754,N_3734,N_3922);
and U4755 (N_4755,N_3161,N_3743);
nand U4756 (N_4756,N_2169,N_2090);
nand U4757 (N_4757,N_3367,N_3200);
or U4758 (N_4758,N_3759,N_2285);
or U4759 (N_4759,N_3810,N_3365);
nor U4760 (N_4760,N_3479,N_2009);
and U4761 (N_4761,N_3403,N_3210);
nor U4762 (N_4762,N_2932,N_2608);
nor U4763 (N_4763,N_3681,N_3932);
nor U4764 (N_4764,N_3330,N_3658);
nand U4765 (N_4765,N_3707,N_2267);
nand U4766 (N_4766,N_3002,N_2004);
or U4767 (N_4767,N_2007,N_2985);
or U4768 (N_4768,N_2278,N_2053);
or U4769 (N_4769,N_3992,N_2855);
and U4770 (N_4770,N_3481,N_2515);
or U4771 (N_4771,N_3092,N_3011);
and U4772 (N_4772,N_2183,N_2543);
nor U4773 (N_4773,N_3414,N_3972);
nor U4774 (N_4774,N_2433,N_3924);
or U4775 (N_4775,N_2656,N_3613);
nor U4776 (N_4776,N_3112,N_3704);
and U4777 (N_4777,N_2834,N_3729);
and U4778 (N_4778,N_3583,N_2380);
nor U4779 (N_4779,N_2493,N_3554);
or U4780 (N_4780,N_3357,N_3027);
nor U4781 (N_4781,N_2517,N_2820);
nor U4782 (N_4782,N_2195,N_3508);
nand U4783 (N_4783,N_2317,N_3911);
nand U4784 (N_4784,N_2295,N_2845);
or U4785 (N_4785,N_3532,N_2717);
and U4786 (N_4786,N_3178,N_2216);
nor U4787 (N_4787,N_2680,N_2152);
or U4788 (N_4788,N_2982,N_2561);
nand U4789 (N_4789,N_2415,N_3445);
nor U4790 (N_4790,N_3877,N_3899);
nor U4791 (N_4791,N_2337,N_2344);
nor U4792 (N_4792,N_3153,N_2963);
and U4793 (N_4793,N_3189,N_3288);
nand U4794 (N_4794,N_3870,N_2551);
and U4795 (N_4795,N_3643,N_3690);
nor U4796 (N_4796,N_2276,N_3496);
and U4797 (N_4797,N_3195,N_3623);
nand U4798 (N_4798,N_2268,N_3244);
nand U4799 (N_4799,N_2526,N_3229);
and U4800 (N_4800,N_2936,N_2549);
xor U4801 (N_4801,N_2898,N_3003);
nand U4802 (N_4802,N_3116,N_2675);
or U4803 (N_4803,N_3323,N_3499);
nor U4804 (N_4804,N_3024,N_3751);
nand U4805 (N_4805,N_3066,N_2231);
nand U4806 (N_4806,N_3410,N_3954);
nor U4807 (N_4807,N_2125,N_3828);
or U4808 (N_4808,N_2757,N_2659);
nor U4809 (N_4809,N_3813,N_3685);
nor U4810 (N_4810,N_3409,N_3644);
nor U4811 (N_4811,N_2949,N_2269);
nand U4812 (N_4812,N_2822,N_3757);
and U4813 (N_4813,N_3886,N_2852);
and U4814 (N_4814,N_2407,N_2753);
or U4815 (N_4815,N_2807,N_2658);
nand U4816 (N_4816,N_2432,N_2580);
and U4817 (N_4817,N_3366,N_2449);
or U4818 (N_4818,N_2550,N_3949);
and U4819 (N_4819,N_2712,N_3089);
nand U4820 (N_4820,N_3777,N_2049);
nand U4821 (N_4821,N_2538,N_2176);
nand U4822 (N_4822,N_3901,N_3718);
nor U4823 (N_4823,N_3824,N_3399);
or U4824 (N_4824,N_3048,N_3163);
and U4825 (N_4825,N_3306,N_2091);
or U4826 (N_4826,N_3386,N_3641);
or U4827 (N_4827,N_3917,N_3530);
nand U4828 (N_4828,N_3135,N_3601);
or U4829 (N_4829,N_2638,N_3345);
and U4830 (N_4830,N_2292,N_3451);
nand U4831 (N_4831,N_2242,N_2774);
or U4832 (N_4832,N_2005,N_2977);
xor U4833 (N_4833,N_3969,N_2718);
or U4834 (N_4834,N_3915,N_2223);
or U4835 (N_4835,N_2790,N_3918);
or U4836 (N_4836,N_2877,N_3346);
or U4837 (N_4837,N_2532,N_2954);
nor U4838 (N_4838,N_3473,N_2866);
or U4839 (N_4839,N_2467,N_2077);
nand U4840 (N_4840,N_3141,N_3371);
nand U4841 (N_4841,N_2225,N_2182);
nor U4842 (N_4842,N_2318,N_3939);
or U4843 (N_4843,N_3936,N_2394);
or U4844 (N_4844,N_2997,N_3638);
and U4845 (N_4845,N_3780,N_2390);
nand U4846 (N_4846,N_2233,N_3095);
nor U4847 (N_4847,N_3376,N_3678);
nand U4848 (N_4848,N_2520,N_3562);
nor U4849 (N_4849,N_3688,N_3184);
nor U4850 (N_4850,N_2568,N_3888);
nor U4851 (N_4851,N_2553,N_3948);
nand U4852 (N_4852,N_2778,N_2084);
or U4853 (N_4853,N_3914,N_2951);
and U4854 (N_4854,N_2417,N_2438);
nor U4855 (N_4855,N_3441,N_3300);
nor U4856 (N_4856,N_3272,N_2800);
nor U4857 (N_4857,N_2328,N_3012);
and U4858 (N_4858,N_3860,N_2749);
nor U4859 (N_4859,N_3029,N_3061);
nor U4860 (N_4860,N_3237,N_3505);
nor U4861 (N_4861,N_3241,N_2609);
or U4862 (N_4862,N_2360,N_2408);
nor U4863 (N_4863,N_3552,N_2014);
and U4864 (N_4864,N_3725,N_3851);
and U4865 (N_4865,N_3507,N_2597);
nor U4866 (N_4866,N_3094,N_2867);
and U4867 (N_4867,N_2393,N_3164);
or U4868 (N_4868,N_2275,N_3645);
xnor U4869 (N_4869,N_2389,N_2714);
nor U4870 (N_4870,N_3278,N_2038);
nor U4871 (N_4871,N_3995,N_2571);
xnor U4872 (N_4872,N_2804,N_2506);
or U4873 (N_4873,N_3476,N_2816);
nand U4874 (N_4874,N_2581,N_2683);
nand U4875 (N_4875,N_2322,N_2672);
or U4876 (N_4876,N_2722,N_3343);
or U4877 (N_4877,N_3848,N_3353);
nor U4878 (N_4878,N_3456,N_2995);
nand U4879 (N_4879,N_2637,N_2575);
and U4880 (N_4880,N_2702,N_3093);
nand U4881 (N_4881,N_3215,N_3347);
and U4882 (N_4882,N_3009,N_3630);
nor U4883 (N_4883,N_3631,N_2721);
or U4884 (N_4884,N_2618,N_2217);
and U4885 (N_4885,N_3238,N_2443);
nor U4886 (N_4886,N_3131,N_2061);
nand U4887 (N_4887,N_3413,N_3175);
or U4888 (N_4888,N_3632,N_2339);
nand U4889 (N_4889,N_3427,N_3863);
and U4890 (N_4890,N_2012,N_3133);
and U4891 (N_4891,N_2321,N_3823);
nor U4892 (N_4892,N_3128,N_2172);
or U4893 (N_4893,N_3880,N_2167);
nand U4894 (N_4894,N_3170,N_2447);
nand U4895 (N_4895,N_3036,N_2842);
xnor U4896 (N_4896,N_2400,N_3512);
or U4897 (N_4897,N_3224,N_2981);
and U4898 (N_4898,N_2196,N_2105);
or U4899 (N_4899,N_3666,N_3619);
nor U4900 (N_4900,N_2298,N_2548);
and U4901 (N_4901,N_2329,N_2404);
nand U4902 (N_4902,N_3429,N_2387);
and U4903 (N_4903,N_2257,N_3871);
or U4904 (N_4904,N_3368,N_3834);
or U4905 (N_4905,N_2170,N_2157);
or U4906 (N_4906,N_2490,N_2146);
and U4907 (N_4907,N_2876,N_2259);
or U4908 (N_4908,N_3622,N_3243);
or U4909 (N_4909,N_2592,N_2698);
nor U4910 (N_4910,N_2887,N_2136);
or U4911 (N_4911,N_3822,N_3349);
xnor U4912 (N_4912,N_3076,N_2868);
nor U4913 (N_4913,N_3542,N_2662);
nor U4914 (N_4914,N_3025,N_3806);
and U4915 (N_4915,N_2930,N_2652);
nand U4916 (N_4916,N_3811,N_3222);
or U4917 (N_4917,N_3603,N_3965);
nor U4918 (N_4918,N_3517,N_2135);
nand U4919 (N_4919,N_3933,N_3521);
nand U4920 (N_4920,N_2596,N_2516);
nor U4921 (N_4921,N_2021,N_3635);
nand U4922 (N_4922,N_3981,N_2270);
nor U4923 (N_4923,N_2690,N_3683);
and U4924 (N_4924,N_2741,N_2929);
nand U4925 (N_4925,N_2657,N_2100);
or U4926 (N_4926,N_2207,N_3234);
or U4927 (N_4927,N_3279,N_2832);
nand U4928 (N_4928,N_3646,N_3331);
nand U4929 (N_4929,N_2023,N_3199);
or U4930 (N_4930,N_2586,N_3280);
or U4931 (N_4931,N_2748,N_3139);
or U4932 (N_4932,N_3038,N_3616);
and U4933 (N_4933,N_2809,N_2377);
and U4934 (N_4934,N_3387,N_3864);
nor U4935 (N_4935,N_2208,N_2667);
or U4936 (N_4936,N_2591,N_3149);
nand U4937 (N_4937,N_3620,N_2296);
and U4938 (N_4938,N_2040,N_2956);
xor U4939 (N_4939,N_3491,N_3675);
and U4940 (N_4940,N_2087,N_3492);
nor U4941 (N_4941,N_2129,N_3753);
nand U4942 (N_4942,N_2858,N_3625);
and U4943 (N_4943,N_3526,N_3020);
and U4944 (N_4944,N_3299,N_2677);
and U4945 (N_4945,N_3217,N_3030);
nand U4946 (N_4946,N_2746,N_2203);
nand U4947 (N_4947,N_3421,N_3579);
nor U4948 (N_4948,N_3134,N_2320);
and U4949 (N_4949,N_3926,N_3982);
nor U4950 (N_4950,N_3669,N_2424);
nand U4951 (N_4951,N_3381,N_3839);
or U4952 (N_4952,N_2472,N_2229);
nand U4953 (N_4953,N_3276,N_2572);
and U4954 (N_4954,N_3802,N_3732);
or U4955 (N_4955,N_2264,N_3121);
and U4956 (N_4956,N_2048,N_3790);
or U4957 (N_4957,N_3697,N_2042);
nand U4958 (N_4958,N_3078,N_2429);
and U4959 (N_4959,N_3432,N_2046);
nor U4960 (N_4960,N_3055,N_2368);
nand U4961 (N_4961,N_3348,N_2243);
nor U4962 (N_4962,N_3468,N_2101);
and U4963 (N_4963,N_2117,N_3997);
nand U4964 (N_4964,N_2833,N_3723);
and U4965 (N_4965,N_3460,N_3415);
nand U4966 (N_4966,N_2854,N_2308);
nor U4967 (N_4967,N_3621,N_2945);
nor U4968 (N_4968,N_3740,N_3578);
nor U4969 (N_4969,N_2036,N_3608);
and U4970 (N_4970,N_3506,N_3907);
nand U4971 (N_4971,N_3487,N_3233);
nor U4972 (N_4972,N_2940,N_3114);
nor U4973 (N_4973,N_2237,N_3702);
and U4974 (N_4974,N_3356,N_2762);
and U4975 (N_4975,N_3138,N_3192);
and U4976 (N_4976,N_2689,N_2777);
nor U4977 (N_4977,N_3803,N_2180);
nor U4978 (N_4978,N_2880,N_2271);
nor U4979 (N_4979,N_3047,N_2755);
nor U4980 (N_4980,N_3789,N_2886);
and U4981 (N_4981,N_2350,N_3741);
nand U4982 (N_4982,N_2660,N_3059);
and U4983 (N_4983,N_3313,N_2988);
and U4984 (N_4984,N_2184,N_3172);
xor U4985 (N_4985,N_3328,N_2300);
or U4986 (N_4986,N_2153,N_2708);
nor U4987 (N_4987,N_2416,N_2128);
and U4988 (N_4988,N_3465,N_3605);
nand U4989 (N_4989,N_3964,N_2150);
xnor U4990 (N_4990,N_3509,N_3281);
nand U4991 (N_4991,N_2245,N_2010);
nor U4992 (N_4992,N_3148,N_3567);
nor U4993 (N_4993,N_2357,N_2470);
xnor U4994 (N_4994,N_3107,N_2342);
or U4995 (N_4995,N_2304,N_3423);
nor U4996 (N_4996,N_2431,N_2953);
nand U4997 (N_4997,N_3853,N_3979);
or U4998 (N_4998,N_2920,N_2481);
or U4999 (N_4999,N_2632,N_3239);
nor U5000 (N_5000,N_3576,N_3262);
or U5001 (N_5001,N_3819,N_3217);
and U5002 (N_5002,N_3025,N_2108);
nand U5003 (N_5003,N_2682,N_3425);
or U5004 (N_5004,N_3242,N_3803);
nor U5005 (N_5005,N_2176,N_3297);
and U5006 (N_5006,N_2468,N_3336);
nand U5007 (N_5007,N_2964,N_2202);
nor U5008 (N_5008,N_3546,N_2844);
and U5009 (N_5009,N_2804,N_2308);
xnor U5010 (N_5010,N_2194,N_3060);
and U5011 (N_5011,N_2145,N_3032);
nor U5012 (N_5012,N_3002,N_3941);
or U5013 (N_5013,N_3750,N_2761);
and U5014 (N_5014,N_3839,N_3820);
nor U5015 (N_5015,N_2405,N_2427);
or U5016 (N_5016,N_3817,N_2182);
or U5017 (N_5017,N_3534,N_2854);
nand U5018 (N_5018,N_2568,N_3979);
nor U5019 (N_5019,N_2470,N_2800);
nor U5020 (N_5020,N_3977,N_3589);
nor U5021 (N_5021,N_2230,N_2328);
nand U5022 (N_5022,N_2069,N_3555);
nand U5023 (N_5023,N_2554,N_3704);
nor U5024 (N_5024,N_2036,N_3353);
and U5025 (N_5025,N_2630,N_2892);
or U5026 (N_5026,N_2928,N_2699);
nor U5027 (N_5027,N_3208,N_3978);
and U5028 (N_5028,N_3736,N_3711);
and U5029 (N_5029,N_3204,N_2346);
and U5030 (N_5030,N_3042,N_2451);
nor U5031 (N_5031,N_3883,N_3766);
or U5032 (N_5032,N_3636,N_3951);
nand U5033 (N_5033,N_3137,N_3473);
nand U5034 (N_5034,N_3955,N_2354);
and U5035 (N_5035,N_2130,N_2527);
or U5036 (N_5036,N_2983,N_2324);
and U5037 (N_5037,N_3923,N_2997);
or U5038 (N_5038,N_2923,N_2955);
nor U5039 (N_5039,N_2898,N_3224);
or U5040 (N_5040,N_2290,N_3656);
nand U5041 (N_5041,N_3941,N_3042);
and U5042 (N_5042,N_2445,N_2285);
and U5043 (N_5043,N_2004,N_3567);
nor U5044 (N_5044,N_2617,N_3593);
nand U5045 (N_5045,N_2605,N_2239);
and U5046 (N_5046,N_2781,N_2188);
or U5047 (N_5047,N_3890,N_2837);
nand U5048 (N_5048,N_2529,N_2629);
or U5049 (N_5049,N_3541,N_2531);
nor U5050 (N_5050,N_3087,N_2765);
nand U5051 (N_5051,N_2917,N_3079);
and U5052 (N_5052,N_2904,N_3068);
or U5053 (N_5053,N_2548,N_3723);
and U5054 (N_5054,N_3473,N_3302);
nand U5055 (N_5055,N_2982,N_2610);
nand U5056 (N_5056,N_3677,N_2269);
nor U5057 (N_5057,N_2075,N_2963);
nand U5058 (N_5058,N_2683,N_2154);
nor U5059 (N_5059,N_3055,N_2996);
nor U5060 (N_5060,N_2107,N_3826);
nand U5061 (N_5061,N_3403,N_3873);
or U5062 (N_5062,N_2294,N_3539);
and U5063 (N_5063,N_3564,N_3462);
or U5064 (N_5064,N_3068,N_3782);
or U5065 (N_5065,N_3955,N_2635);
or U5066 (N_5066,N_2254,N_2008);
and U5067 (N_5067,N_3339,N_3430);
and U5068 (N_5068,N_3734,N_3267);
or U5069 (N_5069,N_2318,N_2398);
nor U5070 (N_5070,N_3700,N_3969);
nor U5071 (N_5071,N_3960,N_3468);
and U5072 (N_5072,N_3103,N_2375);
or U5073 (N_5073,N_3129,N_2279);
and U5074 (N_5074,N_2751,N_2232);
or U5075 (N_5075,N_3874,N_2397);
or U5076 (N_5076,N_3859,N_2745);
or U5077 (N_5077,N_2110,N_3871);
and U5078 (N_5078,N_3925,N_3887);
xnor U5079 (N_5079,N_3863,N_2521);
nand U5080 (N_5080,N_3724,N_3302);
or U5081 (N_5081,N_2570,N_2176);
or U5082 (N_5082,N_3482,N_3732);
and U5083 (N_5083,N_2887,N_2663);
or U5084 (N_5084,N_3656,N_2165);
and U5085 (N_5085,N_3808,N_2459);
and U5086 (N_5086,N_2589,N_2486);
or U5087 (N_5087,N_3853,N_2853);
and U5088 (N_5088,N_2247,N_3425);
or U5089 (N_5089,N_3364,N_3842);
xnor U5090 (N_5090,N_2652,N_3671);
or U5091 (N_5091,N_2610,N_2758);
or U5092 (N_5092,N_3078,N_2586);
nand U5093 (N_5093,N_3782,N_2546);
or U5094 (N_5094,N_3347,N_2405);
nand U5095 (N_5095,N_3558,N_2587);
and U5096 (N_5096,N_3086,N_3103);
or U5097 (N_5097,N_2556,N_2504);
nor U5098 (N_5098,N_2616,N_3137);
nor U5099 (N_5099,N_2836,N_2176);
or U5100 (N_5100,N_2850,N_3210);
and U5101 (N_5101,N_2634,N_3568);
nor U5102 (N_5102,N_2091,N_3695);
nor U5103 (N_5103,N_2805,N_3120);
or U5104 (N_5104,N_2803,N_3751);
nand U5105 (N_5105,N_2693,N_2014);
or U5106 (N_5106,N_2313,N_2437);
nor U5107 (N_5107,N_3568,N_3065);
and U5108 (N_5108,N_2841,N_3737);
nor U5109 (N_5109,N_2192,N_2310);
and U5110 (N_5110,N_3321,N_2475);
nor U5111 (N_5111,N_3992,N_2404);
nor U5112 (N_5112,N_2731,N_2889);
or U5113 (N_5113,N_2031,N_3211);
or U5114 (N_5114,N_2633,N_3961);
or U5115 (N_5115,N_2486,N_3112);
and U5116 (N_5116,N_3884,N_2561);
nand U5117 (N_5117,N_2421,N_3512);
and U5118 (N_5118,N_2665,N_2640);
nand U5119 (N_5119,N_2524,N_3879);
and U5120 (N_5120,N_2211,N_3529);
nand U5121 (N_5121,N_2480,N_3436);
nand U5122 (N_5122,N_2684,N_3943);
nor U5123 (N_5123,N_2922,N_2812);
nand U5124 (N_5124,N_3186,N_3132);
nor U5125 (N_5125,N_2509,N_3643);
nand U5126 (N_5126,N_3792,N_2689);
or U5127 (N_5127,N_3852,N_2686);
nor U5128 (N_5128,N_3691,N_3317);
or U5129 (N_5129,N_2268,N_3253);
and U5130 (N_5130,N_2448,N_3331);
nor U5131 (N_5131,N_3685,N_2729);
nand U5132 (N_5132,N_3055,N_2717);
nor U5133 (N_5133,N_3251,N_3673);
and U5134 (N_5134,N_3465,N_3805);
and U5135 (N_5135,N_3008,N_2557);
nand U5136 (N_5136,N_2206,N_2984);
nor U5137 (N_5137,N_2346,N_3591);
nand U5138 (N_5138,N_3160,N_2349);
xor U5139 (N_5139,N_3407,N_2416);
nand U5140 (N_5140,N_2225,N_3105);
nand U5141 (N_5141,N_3017,N_3398);
nand U5142 (N_5142,N_2423,N_2406);
nand U5143 (N_5143,N_2348,N_3846);
or U5144 (N_5144,N_2019,N_2047);
nand U5145 (N_5145,N_2650,N_3462);
nor U5146 (N_5146,N_3111,N_2997);
xnor U5147 (N_5147,N_3261,N_3219);
and U5148 (N_5148,N_2408,N_3742);
nor U5149 (N_5149,N_3308,N_2422);
or U5150 (N_5150,N_3897,N_3528);
nand U5151 (N_5151,N_3533,N_2455);
nand U5152 (N_5152,N_3998,N_3444);
or U5153 (N_5153,N_2789,N_2592);
or U5154 (N_5154,N_2713,N_3986);
nand U5155 (N_5155,N_3671,N_2186);
nand U5156 (N_5156,N_3311,N_3864);
and U5157 (N_5157,N_2534,N_2233);
and U5158 (N_5158,N_2263,N_2378);
and U5159 (N_5159,N_2178,N_2648);
nor U5160 (N_5160,N_3657,N_2791);
or U5161 (N_5161,N_2876,N_3688);
or U5162 (N_5162,N_3626,N_2198);
and U5163 (N_5163,N_2034,N_3912);
and U5164 (N_5164,N_2490,N_2640);
and U5165 (N_5165,N_3651,N_2705);
nor U5166 (N_5166,N_3832,N_3549);
nor U5167 (N_5167,N_3200,N_3291);
nand U5168 (N_5168,N_2294,N_2398);
nor U5169 (N_5169,N_3813,N_3353);
nand U5170 (N_5170,N_2648,N_2208);
nand U5171 (N_5171,N_3421,N_2818);
and U5172 (N_5172,N_2258,N_3382);
and U5173 (N_5173,N_3410,N_2092);
nor U5174 (N_5174,N_3393,N_2407);
nor U5175 (N_5175,N_3760,N_2212);
nor U5176 (N_5176,N_3320,N_2038);
nand U5177 (N_5177,N_3864,N_3496);
or U5178 (N_5178,N_3033,N_2788);
nand U5179 (N_5179,N_2080,N_2671);
and U5180 (N_5180,N_3791,N_2246);
nand U5181 (N_5181,N_3769,N_2496);
or U5182 (N_5182,N_3306,N_3257);
nand U5183 (N_5183,N_3073,N_3574);
or U5184 (N_5184,N_3871,N_2749);
or U5185 (N_5185,N_2606,N_2869);
and U5186 (N_5186,N_3866,N_2637);
or U5187 (N_5187,N_2746,N_3818);
nor U5188 (N_5188,N_3169,N_2725);
nand U5189 (N_5189,N_3869,N_3881);
or U5190 (N_5190,N_3993,N_2322);
nor U5191 (N_5191,N_2309,N_2424);
nor U5192 (N_5192,N_2979,N_2905);
and U5193 (N_5193,N_2283,N_2153);
or U5194 (N_5194,N_3621,N_3746);
nand U5195 (N_5195,N_3329,N_2407);
nor U5196 (N_5196,N_2735,N_2860);
nand U5197 (N_5197,N_2738,N_2475);
or U5198 (N_5198,N_2575,N_3097);
nor U5199 (N_5199,N_3073,N_2133);
and U5200 (N_5200,N_2820,N_3818);
and U5201 (N_5201,N_3786,N_3479);
and U5202 (N_5202,N_3072,N_3582);
or U5203 (N_5203,N_2738,N_2396);
nor U5204 (N_5204,N_2691,N_3041);
nand U5205 (N_5205,N_2023,N_3121);
and U5206 (N_5206,N_2337,N_3070);
nor U5207 (N_5207,N_3205,N_3033);
and U5208 (N_5208,N_3758,N_2508);
nor U5209 (N_5209,N_2928,N_3667);
or U5210 (N_5210,N_3512,N_3390);
nand U5211 (N_5211,N_3686,N_3996);
or U5212 (N_5212,N_3074,N_3273);
or U5213 (N_5213,N_2283,N_3018);
and U5214 (N_5214,N_3021,N_3730);
and U5215 (N_5215,N_2947,N_2811);
or U5216 (N_5216,N_2783,N_2307);
nand U5217 (N_5217,N_2134,N_2898);
nand U5218 (N_5218,N_3722,N_2624);
and U5219 (N_5219,N_3528,N_2375);
nor U5220 (N_5220,N_2760,N_2006);
nor U5221 (N_5221,N_2926,N_3622);
or U5222 (N_5222,N_3428,N_3647);
nand U5223 (N_5223,N_3710,N_2183);
or U5224 (N_5224,N_2328,N_2958);
or U5225 (N_5225,N_2994,N_3575);
or U5226 (N_5226,N_3172,N_2450);
nand U5227 (N_5227,N_3032,N_3060);
or U5228 (N_5228,N_2289,N_2381);
and U5229 (N_5229,N_3172,N_2920);
and U5230 (N_5230,N_2640,N_2509);
and U5231 (N_5231,N_3262,N_2988);
or U5232 (N_5232,N_2261,N_2974);
or U5233 (N_5233,N_3860,N_2326);
nand U5234 (N_5234,N_2934,N_2391);
or U5235 (N_5235,N_2769,N_2971);
and U5236 (N_5236,N_3942,N_3245);
or U5237 (N_5237,N_2054,N_3140);
xnor U5238 (N_5238,N_2782,N_2909);
nor U5239 (N_5239,N_2887,N_2691);
or U5240 (N_5240,N_3574,N_2093);
and U5241 (N_5241,N_2816,N_3021);
and U5242 (N_5242,N_3603,N_2561);
or U5243 (N_5243,N_2869,N_3080);
nand U5244 (N_5244,N_3322,N_3132);
and U5245 (N_5245,N_2786,N_2504);
and U5246 (N_5246,N_2665,N_2589);
nor U5247 (N_5247,N_2305,N_3175);
nand U5248 (N_5248,N_3566,N_2244);
or U5249 (N_5249,N_3979,N_2622);
and U5250 (N_5250,N_2783,N_2056);
and U5251 (N_5251,N_2539,N_2037);
or U5252 (N_5252,N_3950,N_2321);
nor U5253 (N_5253,N_2920,N_3543);
nand U5254 (N_5254,N_3353,N_3737);
or U5255 (N_5255,N_2581,N_2650);
nand U5256 (N_5256,N_2829,N_2675);
or U5257 (N_5257,N_2266,N_2063);
nand U5258 (N_5258,N_2849,N_3952);
and U5259 (N_5259,N_3101,N_3243);
and U5260 (N_5260,N_3686,N_2030);
and U5261 (N_5261,N_2443,N_3395);
or U5262 (N_5262,N_3391,N_2818);
nor U5263 (N_5263,N_3374,N_2814);
nor U5264 (N_5264,N_3021,N_3532);
and U5265 (N_5265,N_3776,N_2915);
xor U5266 (N_5266,N_2835,N_3222);
or U5267 (N_5267,N_2847,N_3220);
or U5268 (N_5268,N_3919,N_2591);
or U5269 (N_5269,N_3866,N_3128);
nand U5270 (N_5270,N_3412,N_2702);
or U5271 (N_5271,N_3363,N_2479);
and U5272 (N_5272,N_3761,N_3196);
or U5273 (N_5273,N_3766,N_3451);
nand U5274 (N_5274,N_2928,N_2521);
nor U5275 (N_5275,N_3365,N_2537);
nor U5276 (N_5276,N_2461,N_2735);
nor U5277 (N_5277,N_2224,N_2781);
or U5278 (N_5278,N_2650,N_3991);
nand U5279 (N_5279,N_3066,N_3272);
or U5280 (N_5280,N_2972,N_3525);
nor U5281 (N_5281,N_3097,N_3117);
nand U5282 (N_5282,N_3757,N_2720);
and U5283 (N_5283,N_2801,N_3313);
nor U5284 (N_5284,N_3712,N_3812);
or U5285 (N_5285,N_3846,N_2878);
nor U5286 (N_5286,N_3614,N_2407);
nor U5287 (N_5287,N_3786,N_2372);
nor U5288 (N_5288,N_3339,N_3743);
or U5289 (N_5289,N_3488,N_3373);
and U5290 (N_5290,N_3354,N_2868);
nand U5291 (N_5291,N_2208,N_3444);
nand U5292 (N_5292,N_2402,N_2737);
and U5293 (N_5293,N_2983,N_3313);
or U5294 (N_5294,N_2885,N_3953);
nor U5295 (N_5295,N_3368,N_3615);
and U5296 (N_5296,N_2316,N_3489);
or U5297 (N_5297,N_2290,N_3493);
nor U5298 (N_5298,N_2093,N_2150);
nand U5299 (N_5299,N_3449,N_2171);
nand U5300 (N_5300,N_2556,N_2506);
and U5301 (N_5301,N_3099,N_2636);
or U5302 (N_5302,N_3439,N_2801);
nand U5303 (N_5303,N_3388,N_2154);
nor U5304 (N_5304,N_2409,N_2316);
and U5305 (N_5305,N_3167,N_2501);
nand U5306 (N_5306,N_2118,N_3688);
or U5307 (N_5307,N_3259,N_3431);
nor U5308 (N_5308,N_2692,N_2562);
nand U5309 (N_5309,N_2092,N_2745);
nand U5310 (N_5310,N_2781,N_2349);
and U5311 (N_5311,N_3226,N_3111);
nand U5312 (N_5312,N_2794,N_3301);
or U5313 (N_5313,N_2108,N_3006);
nor U5314 (N_5314,N_2726,N_2190);
nor U5315 (N_5315,N_3104,N_2336);
nor U5316 (N_5316,N_3474,N_3028);
nor U5317 (N_5317,N_2021,N_2392);
nor U5318 (N_5318,N_2266,N_2335);
and U5319 (N_5319,N_3408,N_2265);
or U5320 (N_5320,N_3469,N_3729);
nor U5321 (N_5321,N_2809,N_2579);
and U5322 (N_5322,N_2431,N_3928);
and U5323 (N_5323,N_2387,N_3735);
and U5324 (N_5324,N_2688,N_3234);
nand U5325 (N_5325,N_3357,N_3963);
nand U5326 (N_5326,N_3791,N_3916);
nor U5327 (N_5327,N_3103,N_2329);
nor U5328 (N_5328,N_3506,N_2590);
nand U5329 (N_5329,N_2761,N_3184);
and U5330 (N_5330,N_3122,N_3039);
nor U5331 (N_5331,N_3474,N_3773);
nand U5332 (N_5332,N_3250,N_3629);
or U5333 (N_5333,N_2257,N_3396);
xor U5334 (N_5334,N_3528,N_2522);
or U5335 (N_5335,N_2899,N_2010);
nand U5336 (N_5336,N_3793,N_3588);
and U5337 (N_5337,N_2854,N_3704);
and U5338 (N_5338,N_3646,N_2226);
or U5339 (N_5339,N_3200,N_2988);
and U5340 (N_5340,N_2148,N_3866);
nand U5341 (N_5341,N_2528,N_3476);
and U5342 (N_5342,N_2356,N_3315);
or U5343 (N_5343,N_2462,N_3093);
and U5344 (N_5344,N_2180,N_3426);
and U5345 (N_5345,N_2874,N_3587);
nor U5346 (N_5346,N_3131,N_3703);
nor U5347 (N_5347,N_2029,N_3211);
or U5348 (N_5348,N_2038,N_3125);
nand U5349 (N_5349,N_2462,N_2166);
and U5350 (N_5350,N_2141,N_2064);
or U5351 (N_5351,N_3672,N_2107);
or U5352 (N_5352,N_3736,N_3994);
nand U5353 (N_5353,N_3691,N_3527);
or U5354 (N_5354,N_2935,N_3342);
and U5355 (N_5355,N_2953,N_2758);
or U5356 (N_5356,N_2665,N_2728);
and U5357 (N_5357,N_3154,N_3881);
or U5358 (N_5358,N_3638,N_3917);
and U5359 (N_5359,N_3199,N_3478);
or U5360 (N_5360,N_2991,N_2752);
nor U5361 (N_5361,N_2178,N_3561);
and U5362 (N_5362,N_2010,N_3629);
nand U5363 (N_5363,N_2311,N_2595);
nand U5364 (N_5364,N_2486,N_3306);
nand U5365 (N_5365,N_3658,N_3692);
nor U5366 (N_5366,N_3329,N_3170);
nand U5367 (N_5367,N_3778,N_3699);
nor U5368 (N_5368,N_3865,N_3856);
or U5369 (N_5369,N_2418,N_2129);
or U5370 (N_5370,N_2903,N_2662);
and U5371 (N_5371,N_3881,N_3666);
nand U5372 (N_5372,N_2502,N_3157);
nor U5373 (N_5373,N_2075,N_3088);
or U5374 (N_5374,N_3755,N_3811);
or U5375 (N_5375,N_2755,N_2609);
nor U5376 (N_5376,N_2571,N_2066);
nand U5377 (N_5377,N_2225,N_2755);
and U5378 (N_5378,N_3444,N_2012);
or U5379 (N_5379,N_3880,N_3993);
nor U5380 (N_5380,N_2688,N_2649);
or U5381 (N_5381,N_3307,N_2455);
or U5382 (N_5382,N_3747,N_3090);
or U5383 (N_5383,N_2481,N_3789);
nor U5384 (N_5384,N_2750,N_3685);
nand U5385 (N_5385,N_2863,N_3534);
nor U5386 (N_5386,N_2000,N_3176);
nor U5387 (N_5387,N_3904,N_2303);
nor U5388 (N_5388,N_3946,N_2105);
or U5389 (N_5389,N_3812,N_2136);
nand U5390 (N_5390,N_3943,N_3811);
and U5391 (N_5391,N_3563,N_3405);
nand U5392 (N_5392,N_2268,N_3551);
nand U5393 (N_5393,N_3438,N_3395);
or U5394 (N_5394,N_3247,N_3487);
nand U5395 (N_5395,N_2395,N_3257);
nor U5396 (N_5396,N_2132,N_2344);
or U5397 (N_5397,N_3727,N_3088);
and U5398 (N_5398,N_2588,N_3790);
or U5399 (N_5399,N_2706,N_2528);
or U5400 (N_5400,N_2600,N_2807);
nand U5401 (N_5401,N_3601,N_3023);
nor U5402 (N_5402,N_2755,N_2378);
nor U5403 (N_5403,N_3700,N_2160);
and U5404 (N_5404,N_2736,N_3805);
nand U5405 (N_5405,N_3065,N_2655);
nand U5406 (N_5406,N_2692,N_2289);
nor U5407 (N_5407,N_2078,N_3069);
nor U5408 (N_5408,N_2275,N_3364);
or U5409 (N_5409,N_2066,N_3542);
or U5410 (N_5410,N_2858,N_2083);
nor U5411 (N_5411,N_2898,N_2719);
and U5412 (N_5412,N_2563,N_3743);
nor U5413 (N_5413,N_2065,N_2333);
nor U5414 (N_5414,N_3244,N_3698);
nor U5415 (N_5415,N_2481,N_3058);
or U5416 (N_5416,N_2843,N_3604);
nand U5417 (N_5417,N_2067,N_2293);
and U5418 (N_5418,N_3708,N_3184);
and U5419 (N_5419,N_3181,N_3175);
nor U5420 (N_5420,N_3934,N_2147);
nand U5421 (N_5421,N_2516,N_2954);
nand U5422 (N_5422,N_3065,N_2915);
nand U5423 (N_5423,N_3410,N_3432);
or U5424 (N_5424,N_2841,N_2205);
nor U5425 (N_5425,N_3903,N_3418);
nor U5426 (N_5426,N_3209,N_2639);
or U5427 (N_5427,N_3184,N_2678);
nor U5428 (N_5428,N_2479,N_3610);
nor U5429 (N_5429,N_2078,N_3847);
or U5430 (N_5430,N_3081,N_3062);
and U5431 (N_5431,N_3108,N_2494);
nor U5432 (N_5432,N_3592,N_3566);
nor U5433 (N_5433,N_2559,N_2926);
nor U5434 (N_5434,N_3634,N_2581);
and U5435 (N_5435,N_3531,N_2263);
nand U5436 (N_5436,N_2818,N_2947);
nor U5437 (N_5437,N_3559,N_3025);
and U5438 (N_5438,N_3263,N_3987);
xnor U5439 (N_5439,N_3981,N_3320);
nand U5440 (N_5440,N_2369,N_2874);
or U5441 (N_5441,N_2371,N_2289);
or U5442 (N_5442,N_3993,N_2461);
and U5443 (N_5443,N_3278,N_3428);
nand U5444 (N_5444,N_2240,N_2083);
nor U5445 (N_5445,N_2573,N_2793);
nand U5446 (N_5446,N_2739,N_3328);
or U5447 (N_5447,N_2805,N_3488);
or U5448 (N_5448,N_3745,N_3017);
nand U5449 (N_5449,N_3665,N_3190);
and U5450 (N_5450,N_2248,N_2239);
and U5451 (N_5451,N_2877,N_3274);
xor U5452 (N_5452,N_3381,N_2897);
and U5453 (N_5453,N_2273,N_3790);
or U5454 (N_5454,N_2703,N_3450);
nand U5455 (N_5455,N_2289,N_2915);
nand U5456 (N_5456,N_2194,N_3742);
or U5457 (N_5457,N_3559,N_2368);
nand U5458 (N_5458,N_2505,N_2090);
and U5459 (N_5459,N_2313,N_2367);
or U5460 (N_5460,N_2335,N_3298);
xor U5461 (N_5461,N_2293,N_2933);
nor U5462 (N_5462,N_2298,N_2837);
and U5463 (N_5463,N_3696,N_3206);
or U5464 (N_5464,N_2790,N_3541);
xor U5465 (N_5465,N_3655,N_3437);
or U5466 (N_5466,N_2114,N_3544);
nor U5467 (N_5467,N_3731,N_2116);
nor U5468 (N_5468,N_3218,N_3855);
nand U5469 (N_5469,N_3862,N_2818);
nor U5470 (N_5470,N_2733,N_3673);
and U5471 (N_5471,N_3771,N_2429);
nor U5472 (N_5472,N_2279,N_3712);
or U5473 (N_5473,N_3954,N_3551);
nand U5474 (N_5474,N_3400,N_3769);
nor U5475 (N_5475,N_2331,N_2572);
nor U5476 (N_5476,N_3858,N_3040);
nand U5477 (N_5477,N_3623,N_2708);
and U5478 (N_5478,N_3703,N_3932);
and U5479 (N_5479,N_3232,N_3661);
nand U5480 (N_5480,N_3516,N_3174);
or U5481 (N_5481,N_2258,N_3898);
nand U5482 (N_5482,N_3195,N_3729);
or U5483 (N_5483,N_2921,N_2857);
xnor U5484 (N_5484,N_3840,N_3193);
nor U5485 (N_5485,N_3348,N_3586);
and U5486 (N_5486,N_3339,N_3283);
nand U5487 (N_5487,N_2623,N_3457);
nand U5488 (N_5488,N_2239,N_3986);
nor U5489 (N_5489,N_3144,N_3164);
and U5490 (N_5490,N_2483,N_3616);
or U5491 (N_5491,N_2735,N_2808);
and U5492 (N_5492,N_3701,N_2898);
nand U5493 (N_5493,N_2714,N_2461);
or U5494 (N_5494,N_2722,N_2019);
nand U5495 (N_5495,N_3703,N_2098);
and U5496 (N_5496,N_2988,N_3747);
and U5497 (N_5497,N_3788,N_3467);
or U5498 (N_5498,N_2991,N_3528);
or U5499 (N_5499,N_2851,N_2247);
or U5500 (N_5500,N_3159,N_3864);
nand U5501 (N_5501,N_3707,N_3527);
or U5502 (N_5502,N_2118,N_3159);
nand U5503 (N_5503,N_3619,N_3368);
nor U5504 (N_5504,N_2827,N_2679);
or U5505 (N_5505,N_3594,N_2768);
or U5506 (N_5506,N_3251,N_3725);
nand U5507 (N_5507,N_2081,N_3058);
nor U5508 (N_5508,N_2457,N_2239);
nand U5509 (N_5509,N_3908,N_3955);
and U5510 (N_5510,N_2185,N_3767);
nand U5511 (N_5511,N_2442,N_3143);
nor U5512 (N_5512,N_3616,N_3081);
nor U5513 (N_5513,N_3303,N_2140);
nand U5514 (N_5514,N_2711,N_3119);
nand U5515 (N_5515,N_3388,N_2375);
nor U5516 (N_5516,N_3371,N_3010);
or U5517 (N_5517,N_2372,N_2583);
or U5518 (N_5518,N_2990,N_2040);
and U5519 (N_5519,N_2349,N_3183);
nor U5520 (N_5520,N_3122,N_2732);
nand U5521 (N_5521,N_2753,N_2215);
nor U5522 (N_5522,N_2856,N_2130);
nor U5523 (N_5523,N_2703,N_2487);
or U5524 (N_5524,N_2529,N_2251);
or U5525 (N_5525,N_2960,N_3370);
nor U5526 (N_5526,N_2335,N_2854);
and U5527 (N_5527,N_3333,N_2586);
and U5528 (N_5528,N_3187,N_3222);
or U5529 (N_5529,N_2774,N_3633);
nor U5530 (N_5530,N_3460,N_3456);
or U5531 (N_5531,N_2229,N_3755);
nor U5532 (N_5532,N_3530,N_3204);
and U5533 (N_5533,N_2854,N_2152);
and U5534 (N_5534,N_3111,N_3097);
nor U5535 (N_5535,N_2969,N_2298);
and U5536 (N_5536,N_3446,N_2991);
nor U5537 (N_5537,N_3501,N_3871);
nor U5538 (N_5538,N_2212,N_2872);
or U5539 (N_5539,N_2517,N_3844);
and U5540 (N_5540,N_3846,N_3360);
and U5541 (N_5541,N_3151,N_2037);
or U5542 (N_5542,N_3448,N_3237);
and U5543 (N_5543,N_3054,N_3470);
and U5544 (N_5544,N_2488,N_3126);
nand U5545 (N_5545,N_3112,N_2358);
nand U5546 (N_5546,N_2902,N_3161);
nor U5547 (N_5547,N_3205,N_3722);
nor U5548 (N_5548,N_2982,N_2473);
or U5549 (N_5549,N_2414,N_3312);
nor U5550 (N_5550,N_3208,N_2432);
nor U5551 (N_5551,N_2647,N_2868);
nor U5552 (N_5552,N_2509,N_3128);
or U5553 (N_5553,N_3098,N_2737);
or U5554 (N_5554,N_3675,N_3990);
or U5555 (N_5555,N_3589,N_2316);
and U5556 (N_5556,N_2345,N_2740);
nor U5557 (N_5557,N_2163,N_2026);
nor U5558 (N_5558,N_2934,N_2158);
nor U5559 (N_5559,N_3419,N_2713);
nand U5560 (N_5560,N_2745,N_3716);
or U5561 (N_5561,N_3820,N_3195);
and U5562 (N_5562,N_2670,N_3940);
and U5563 (N_5563,N_2175,N_3885);
nand U5564 (N_5564,N_3297,N_2692);
or U5565 (N_5565,N_3126,N_2890);
and U5566 (N_5566,N_3332,N_2252);
nand U5567 (N_5567,N_3415,N_3318);
or U5568 (N_5568,N_2376,N_3025);
and U5569 (N_5569,N_2285,N_2880);
and U5570 (N_5570,N_3876,N_2866);
or U5571 (N_5571,N_3729,N_3981);
or U5572 (N_5572,N_3163,N_2097);
nor U5573 (N_5573,N_2452,N_2850);
and U5574 (N_5574,N_2450,N_3634);
xor U5575 (N_5575,N_3409,N_2671);
nand U5576 (N_5576,N_3840,N_3084);
or U5577 (N_5577,N_2322,N_2424);
or U5578 (N_5578,N_3414,N_2167);
and U5579 (N_5579,N_3297,N_2712);
nor U5580 (N_5580,N_2699,N_2686);
nand U5581 (N_5581,N_2796,N_2443);
or U5582 (N_5582,N_2144,N_2549);
nor U5583 (N_5583,N_2823,N_2897);
nand U5584 (N_5584,N_3706,N_3743);
nor U5585 (N_5585,N_2356,N_3268);
and U5586 (N_5586,N_2942,N_3662);
xor U5587 (N_5587,N_2475,N_3639);
and U5588 (N_5588,N_2635,N_3251);
and U5589 (N_5589,N_2927,N_2891);
or U5590 (N_5590,N_3992,N_3344);
and U5591 (N_5591,N_2220,N_2136);
or U5592 (N_5592,N_3525,N_3218);
nand U5593 (N_5593,N_2807,N_3260);
nand U5594 (N_5594,N_3346,N_2620);
nand U5595 (N_5595,N_3241,N_3461);
nor U5596 (N_5596,N_3574,N_3367);
nand U5597 (N_5597,N_3127,N_2398);
nor U5598 (N_5598,N_3299,N_2475);
and U5599 (N_5599,N_3411,N_2734);
nor U5600 (N_5600,N_2981,N_2055);
nand U5601 (N_5601,N_2204,N_3504);
or U5602 (N_5602,N_3098,N_3031);
nand U5603 (N_5603,N_3708,N_3605);
nor U5604 (N_5604,N_2197,N_2275);
nand U5605 (N_5605,N_3358,N_2469);
or U5606 (N_5606,N_3686,N_2058);
or U5607 (N_5607,N_2263,N_2535);
nor U5608 (N_5608,N_3207,N_2403);
nor U5609 (N_5609,N_2444,N_3708);
nand U5610 (N_5610,N_2779,N_3041);
nor U5611 (N_5611,N_2284,N_2791);
or U5612 (N_5612,N_2233,N_2770);
nand U5613 (N_5613,N_3993,N_3442);
nand U5614 (N_5614,N_3860,N_3578);
or U5615 (N_5615,N_3078,N_3067);
nor U5616 (N_5616,N_2705,N_2220);
nand U5617 (N_5617,N_3337,N_3092);
nor U5618 (N_5618,N_3847,N_3217);
xnor U5619 (N_5619,N_2897,N_3693);
and U5620 (N_5620,N_2721,N_2264);
or U5621 (N_5621,N_2371,N_2391);
nor U5622 (N_5622,N_2924,N_2278);
nand U5623 (N_5623,N_2543,N_2552);
and U5624 (N_5624,N_3189,N_3352);
and U5625 (N_5625,N_2351,N_3679);
nor U5626 (N_5626,N_2380,N_3431);
or U5627 (N_5627,N_2866,N_2777);
nand U5628 (N_5628,N_2846,N_2101);
nor U5629 (N_5629,N_2744,N_3620);
nor U5630 (N_5630,N_3441,N_2079);
and U5631 (N_5631,N_3309,N_3573);
nand U5632 (N_5632,N_3449,N_3088);
or U5633 (N_5633,N_3295,N_2660);
nor U5634 (N_5634,N_3677,N_2539);
or U5635 (N_5635,N_2050,N_3656);
nand U5636 (N_5636,N_2884,N_2054);
nand U5637 (N_5637,N_3997,N_3855);
and U5638 (N_5638,N_3320,N_3597);
and U5639 (N_5639,N_2562,N_2427);
nor U5640 (N_5640,N_3421,N_2423);
nand U5641 (N_5641,N_2885,N_2755);
or U5642 (N_5642,N_2324,N_3059);
and U5643 (N_5643,N_3248,N_2355);
nand U5644 (N_5644,N_3248,N_2057);
or U5645 (N_5645,N_2794,N_3245);
nor U5646 (N_5646,N_3615,N_3924);
and U5647 (N_5647,N_2669,N_3464);
or U5648 (N_5648,N_2925,N_3939);
or U5649 (N_5649,N_3166,N_2736);
nand U5650 (N_5650,N_2412,N_3380);
and U5651 (N_5651,N_3344,N_3209);
and U5652 (N_5652,N_3063,N_2157);
nor U5653 (N_5653,N_2138,N_3483);
and U5654 (N_5654,N_2995,N_3678);
nor U5655 (N_5655,N_3293,N_2325);
nand U5656 (N_5656,N_3709,N_2169);
and U5657 (N_5657,N_3902,N_3188);
or U5658 (N_5658,N_3689,N_3098);
or U5659 (N_5659,N_3943,N_3062);
nor U5660 (N_5660,N_2856,N_3370);
or U5661 (N_5661,N_3711,N_3013);
nor U5662 (N_5662,N_3368,N_3181);
or U5663 (N_5663,N_3370,N_3130);
nand U5664 (N_5664,N_3187,N_3004);
and U5665 (N_5665,N_3657,N_3870);
or U5666 (N_5666,N_3088,N_2267);
nor U5667 (N_5667,N_2165,N_2747);
nor U5668 (N_5668,N_2084,N_2322);
or U5669 (N_5669,N_3502,N_2795);
nand U5670 (N_5670,N_3449,N_2633);
xnor U5671 (N_5671,N_3364,N_3702);
or U5672 (N_5672,N_3759,N_2144);
nand U5673 (N_5673,N_2910,N_3733);
or U5674 (N_5674,N_2927,N_2651);
nand U5675 (N_5675,N_2178,N_2816);
nor U5676 (N_5676,N_3309,N_3092);
nor U5677 (N_5677,N_3746,N_2193);
or U5678 (N_5678,N_2463,N_2588);
nor U5679 (N_5679,N_3759,N_2794);
nor U5680 (N_5680,N_3640,N_2647);
nand U5681 (N_5681,N_3790,N_2600);
or U5682 (N_5682,N_2171,N_2960);
nor U5683 (N_5683,N_3366,N_3718);
or U5684 (N_5684,N_3837,N_2859);
and U5685 (N_5685,N_2569,N_3043);
nor U5686 (N_5686,N_3662,N_2180);
or U5687 (N_5687,N_3256,N_3964);
nand U5688 (N_5688,N_2706,N_3119);
nor U5689 (N_5689,N_3538,N_2985);
and U5690 (N_5690,N_3754,N_3099);
nand U5691 (N_5691,N_3214,N_2373);
nand U5692 (N_5692,N_3225,N_2830);
nor U5693 (N_5693,N_2911,N_3766);
nand U5694 (N_5694,N_3127,N_2609);
and U5695 (N_5695,N_2119,N_3946);
and U5696 (N_5696,N_3401,N_3651);
nor U5697 (N_5697,N_2068,N_3925);
nor U5698 (N_5698,N_2739,N_2630);
or U5699 (N_5699,N_3501,N_2763);
nor U5700 (N_5700,N_3003,N_3381);
and U5701 (N_5701,N_3912,N_2638);
or U5702 (N_5702,N_3978,N_3524);
nand U5703 (N_5703,N_3289,N_3174);
nor U5704 (N_5704,N_2154,N_3648);
nor U5705 (N_5705,N_2487,N_3849);
or U5706 (N_5706,N_3925,N_2583);
and U5707 (N_5707,N_3629,N_2801);
and U5708 (N_5708,N_3697,N_3132);
nand U5709 (N_5709,N_2314,N_2623);
nor U5710 (N_5710,N_2062,N_2860);
xnor U5711 (N_5711,N_3909,N_3525);
or U5712 (N_5712,N_3631,N_2028);
nand U5713 (N_5713,N_2419,N_3400);
nor U5714 (N_5714,N_2605,N_3213);
and U5715 (N_5715,N_3843,N_2342);
or U5716 (N_5716,N_2672,N_2229);
nand U5717 (N_5717,N_2234,N_2370);
and U5718 (N_5718,N_3438,N_2278);
nand U5719 (N_5719,N_3122,N_2308);
nor U5720 (N_5720,N_3370,N_2517);
nand U5721 (N_5721,N_3694,N_2079);
nand U5722 (N_5722,N_2546,N_3017);
nand U5723 (N_5723,N_3306,N_3160);
or U5724 (N_5724,N_3922,N_2341);
nor U5725 (N_5725,N_3206,N_2731);
and U5726 (N_5726,N_2579,N_2922);
and U5727 (N_5727,N_3862,N_2649);
nand U5728 (N_5728,N_3641,N_2351);
and U5729 (N_5729,N_2792,N_3963);
or U5730 (N_5730,N_3617,N_3805);
and U5731 (N_5731,N_2201,N_3651);
nor U5732 (N_5732,N_2705,N_3166);
or U5733 (N_5733,N_2063,N_2693);
or U5734 (N_5734,N_3088,N_3765);
nor U5735 (N_5735,N_3152,N_3883);
and U5736 (N_5736,N_3304,N_3418);
and U5737 (N_5737,N_2186,N_2670);
nand U5738 (N_5738,N_2002,N_2082);
nand U5739 (N_5739,N_3476,N_2526);
or U5740 (N_5740,N_2390,N_3837);
nand U5741 (N_5741,N_3171,N_2253);
or U5742 (N_5742,N_3351,N_3405);
or U5743 (N_5743,N_2422,N_3891);
nor U5744 (N_5744,N_3527,N_2087);
nand U5745 (N_5745,N_3317,N_2325);
nand U5746 (N_5746,N_3584,N_2708);
nor U5747 (N_5747,N_3248,N_2237);
nand U5748 (N_5748,N_2665,N_3233);
xnor U5749 (N_5749,N_2649,N_3466);
nand U5750 (N_5750,N_2765,N_3131);
nand U5751 (N_5751,N_2706,N_3432);
or U5752 (N_5752,N_2069,N_3401);
nand U5753 (N_5753,N_2241,N_3689);
or U5754 (N_5754,N_3444,N_3073);
or U5755 (N_5755,N_2905,N_2699);
and U5756 (N_5756,N_2238,N_3681);
and U5757 (N_5757,N_3573,N_3458);
and U5758 (N_5758,N_3940,N_3318);
nor U5759 (N_5759,N_3200,N_2702);
nor U5760 (N_5760,N_3121,N_3789);
and U5761 (N_5761,N_3165,N_2807);
nor U5762 (N_5762,N_3712,N_3903);
nand U5763 (N_5763,N_3079,N_2388);
or U5764 (N_5764,N_3231,N_3764);
nor U5765 (N_5765,N_3112,N_3876);
nor U5766 (N_5766,N_3827,N_2575);
or U5767 (N_5767,N_2897,N_3875);
nand U5768 (N_5768,N_3447,N_3234);
and U5769 (N_5769,N_2783,N_3827);
and U5770 (N_5770,N_3977,N_2950);
and U5771 (N_5771,N_2988,N_3615);
nor U5772 (N_5772,N_2422,N_3205);
nor U5773 (N_5773,N_2451,N_2847);
nand U5774 (N_5774,N_3466,N_3467);
nor U5775 (N_5775,N_2029,N_3043);
and U5776 (N_5776,N_3626,N_2203);
or U5777 (N_5777,N_3819,N_3629);
nand U5778 (N_5778,N_2659,N_2057);
nor U5779 (N_5779,N_3783,N_3163);
and U5780 (N_5780,N_2431,N_2465);
or U5781 (N_5781,N_2553,N_3235);
or U5782 (N_5782,N_3230,N_2715);
and U5783 (N_5783,N_2766,N_2534);
nor U5784 (N_5784,N_2383,N_3514);
or U5785 (N_5785,N_2424,N_3918);
nand U5786 (N_5786,N_3049,N_2708);
and U5787 (N_5787,N_3286,N_2003);
nor U5788 (N_5788,N_2930,N_3294);
or U5789 (N_5789,N_2900,N_2563);
and U5790 (N_5790,N_2614,N_3924);
nor U5791 (N_5791,N_3981,N_2624);
and U5792 (N_5792,N_2375,N_3998);
or U5793 (N_5793,N_3752,N_3465);
nand U5794 (N_5794,N_2495,N_2291);
and U5795 (N_5795,N_2040,N_2985);
nor U5796 (N_5796,N_2144,N_2315);
nor U5797 (N_5797,N_3187,N_2342);
nand U5798 (N_5798,N_3209,N_3501);
or U5799 (N_5799,N_3503,N_3007);
xnor U5800 (N_5800,N_3865,N_2010);
or U5801 (N_5801,N_3122,N_3210);
nor U5802 (N_5802,N_2273,N_3538);
and U5803 (N_5803,N_2066,N_2605);
and U5804 (N_5804,N_2323,N_3316);
nand U5805 (N_5805,N_3965,N_3487);
nand U5806 (N_5806,N_2896,N_3692);
and U5807 (N_5807,N_2920,N_3654);
nand U5808 (N_5808,N_2575,N_2193);
nor U5809 (N_5809,N_2500,N_2009);
nand U5810 (N_5810,N_2464,N_2228);
nor U5811 (N_5811,N_3425,N_2388);
nand U5812 (N_5812,N_2601,N_2011);
and U5813 (N_5813,N_3899,N_3861);
nor U5814 (N_5814,N_2827,N_3424);
nand U5815 (N_5815,N_3905,N_3798);
or U5816 (N_5816,N_2554,N_3976);
or U5817 (N_5817,N_2247,N_2544);
and U5818 (N_5818,N_2386,N_3114);
nor U5819 (N_5819,N_3291,N_2344);
nand U5820 (N_5820,N_3293,N_3913);
and U5821 (N_5821,N_2135,N_3894);
or U5822 (N_5822,N_3513,N_3301);
nand U5823 (N_5823,N_2695,N_2617);
nor U5824 (N_5824,N_2706,N_3224);
nor U5825 (N_5825,N_2790,N_2013);
nor U5826 (N_5826,N_3349,N_3040);
nand U5827 (N_5827,N_2883,N_3534);
and U5828 (N_5828,N_3366,N_2779);
or U5829 (N_5829,N_2277,N_3136);
or U5830 (N_5830,N_2134,N_2110);
or U5831 (N_5831,N_3045,N_3964);
nor U5832 (N_5832,N_2219,N_3450);
and U5833 (N_5833,N_3070,N_3802);
nand U5834 (N_5834,N_3258,N_3252);
nand U5835 (N_5835,N_3089,N_2247);
and U5836 (N_5836,N_3667,N_2403);
nand U5837 (N_5837,N_3258,N_3893);
nor U5838 (N_5838,N_3266,N_2835);
nor U5839 (N_5839,N_3480,N_3234);
or U5840 (N_5840,N_2264,N_3791);
xor U5841 (N_5841,N_2272,N_3708);
and U5842 (N_5842,N_3932,N_2409);
and U5843 (N_5843,N_3807,N_3387);
nor U5844 (N_5844,N_2155,N_3137);
and U5845 (N_5845,N_3382,N_3282);
or U5846 (N_5846,N_2840,N_2554);
nand U5847 (N_5847,N_2960,N_3362);
nand U5848 (N_5848,N_2586,N_2641);
nor U5849 (N_5849,N_3288,N_2506);
nand U5850 (N_5850,N_3797,N_2493);
nand U5851 (N_5851,N_3495,N_2465);
and U5852 (N_5852,N_3682,N_3859);
nor U5853 (N_5853,N_2227,N_3730);
and U5854 (N_5854,N_3100,N_3612);
or U5855 (N_5855,N_2908,N_3241);
nor U5856 (N_5856,N_2835,N_3020);
or U5857 (N_5857,N_2086,N_2557);
nand U5858 (N_5858,N_2699,N_2812);
nor U5859 (N_5859,N_2256,N_3999);
nand U5860 (N_5860,N_3141,N_3459);
and U5861 (N_5861,N_2780,N_3520);
nor U5862 (N_5862,N_3326,N_3507);
nor U5863 (N_5863,N_3828,N_2668);
or U5864 (N_5864,N_2959,N_2991);
nor U5865 (N_5865,N_2475,N_2217);
nor U5866 (N_5866,N_3672,N_2691);
or U5867 (N_5867,N_2139,N_3392);
and U5868 (N_5868,N_2490,N_3617);
and U5869 (N_5869,N_3786,N_3118);
nor U5870 (N_5870,N_3485,N_3152);
and U5871 (N_5871,N_2283,N_3992);
nor U5872 (N_5872,N_2065,N_2902);
nand U5873 (N_5873,N_2782,N_2037);
nor U5874 (N_5874,N_3507,N_3977);
xor U5875 (N_5875,N_3192,N_2131);
and U5876 (N_5876,N_2223,N_3185);
and U5877 (N_5877,N_3192,N_2451);
and U5878 (N_5878,N_3616,N_3855);
and U5879 (N_5879,N_3894,N_2227);
nand U5880 (N_5880,N_3090,N_2081);
nor U5881 (N_5881,N_2199,N_2555);
and U5882 (N_5882,N_3061,N_3391);
or U5883 (N_5883,N_3994,N_2561);
nand U5884 (N_5884,N_2982,N_3786);
and U5885 (N_5885,N_3919,N_2449);
nand U5886 (N_5886,N_3543,N_3023);
nand U5887 (N_5887,N_3927,N_3906);
or U5888 (N_5888,N_3157,N_3769);
or U5889 (N_5889,N_3867,N_2843);
nand U5890 (N_5890,N_3023,N_2724);
and U5891 (N_5891,N_3675,N_2838);
and U5892 (N_5892,N_2910,N_3172);
and U5893 (N_5893,N_2961,N_3166);
nand U5894 (N_5894,N_2669,N_2449);
nor U5895 (N_5895,N_2592,N_2347);
nor U5896 (N_5896,N_3750,N_2890);
nor U5897 (N_5897,N_2640,N_2992);
nand U5898 (N_5898,N_2791,N_2334);
or U5899 (N_5899,N_3004,N_2044);
nand U5900 (N_5900,N_3514,N_3556);
xnor U5901 (N_5901,N_3713,N_3658);
nor U5902 (N_5902,N_3331,N_3602);
nand U5903 (N_5903,N_3605,N_2025);
or U5904 (N_5904,N_3848,N_2137);
nand U5905 (N_5905,N_2964,N_3994);
or U5906 (N_5906,N_2280,N_3732);
nand U5907 (N_5907,N_2327,N_3278);
nand U5908 (N_5908,N_2603,N_2760);
nor U5909 (N_5909,N_2993,N_2622);
nor U5910 (N_5910,N_3047,N_3038);
or U5911 (N_5911,N_3522,N_2018);
nand U5912 (N_5912,N_3303,N_3340);
nor U5913 (N_5913,N_2097,N_3089);
or U5914 (N_5914,N_2315,N_2827);
or U5915 (N_5915,N_2802,N_2280);
nor U5916 (N_5916,N_2194,N_2236);
and U5917 (N_5917,N_3559,N_2290);
and U5918 (N_5918,N_2459,N_3261);
nand U5919 (N_5919,N_3818,N_2587);
nor U5920 (N_5920,N_2766,N_2368);
or U5921 (N_5921,N_2604,N_3744);
or U5922 (N_5922,N_2449,N_2429);
or U5923 (N_5923,N_2003,N_3357);
nand U5924 (N_5924,N_3742,N_2986);
nand U5925 (N_5925,N_2684,N_3665);
or U5926 (N_5926,N_3075,N_3718);
or U5927 (N_5927,N_3665,N_2807);
nor U5928 (N_5928,N_3932,N_3731);
and U5929 (N_5929,N_2255,N_3107);
or U5930 (N_5930,N_3374,N_2169);
or U5931 (N_5931,N_2354,N_2739);
or U5932 (N_5932,N_3411,N_3886);
nor U5933 (N_5933,N_2338,N_2004);
or U5934 (N_5934,N_3150,N_3402);
nand U5935 (N_5935,N_3018,N_3049);
and U5936 (N_5936,N_2996,N_3869);
xor U5937 (N_5937,N_2613,N_3524);
nor U5938 (N_5938,N_2412,N_3940);
or U5939 (N_5939,N_3836,N_3546);
nand U5940 (N_5940,N_2968,N_2609);
nor U5941 (N_5941,N_2886,N_2157);
nor U5942 (N_5942,N_2950,N_3047);
or U5943 (N_5943,N_2916,N_2393);
nand U5944 (N_5944,N_3705,N_3513);
or U5945 (N_5945,N_2279,N_2395);
nor U5946 (N_5946,N_3252,N_2065);
and U5947 (N_5947,N_3018,N_3980);
and U5948 (N_5948,N_2580,N_3268);
or U5949 (N_5949,N_2394,N_3291);
and U5950 (N_5950,N_3609,N_2846);
or U5951 (N_5951,N_2895,N_2323);
nor U5952 (N_5952,N_3562,N_3791);
nor U5953 (N_5953,N_3843,N_3133);
nor U5954 (N_5954,N_3880,N_2346);
nand U5955 (N_5955,N_3797,N_3245);
nor U5956 (N_5956,N_3255,N_2141);
and U5957 (N_5957,N_3874,N_2398);
or U5958 (N_5958,N_2544,N_3576);
or U5959 (N_5959,N_3919,N_3131);
nor U5960 (N_5960,N_2400,N_2688);
nand U5961 (N_5961,N_2274,N_2769);
or U5962 (N_5962,N_2680,N_3693);
nor U5963 (N_5963,N_2809,N_2711);
nand U5964 (N_5964,N_2470,N_2637);
or U5965 (N_5965,N_3887,N_2409);
nand U5966 (N_5966,N_2065,N_3455);
and U5967 (N_5967,N_3951,N_3233);
and U5968 (N_5968,N_3502,N_2122);
nand U5969 (N_5969,N_3873,N_2893);
nand U5970 (N_5970,N_3615,N_2130);
nor U5971 (N_5971,N_3918,N_2999);
or U5972 (N_5972,N_3117,N_2882);
nand U5973 (N_5973,N_2284,N_3672);
or U5974 (N_5974,N_2265,N_2694);
or U5975 (N_5975,N_2594,N_3331);
and U5976 (N_5976,N_2031,N_2148);
nor U5977 (N_5977,N_2546,N_3315);
or U5978 (N_5978,N_2583,N_2892);
nor U5979 (N_5979,N_2969,N_2345);
nand U5980 (N_5980,N_2516,N_2855);
nand U5981 (N_5981,N_2445,N_3846);
xor U5982 (N_5982,N_3469,N_3636);
nor U5983 (N_5983,N_3754,N_2247);
nand U5984 (N_5984,N_3396,N_3186);
nor U5985 (N_5985,N_2667,N_2524);
nand U5986 (N_5986,N_3587,N_3647);
nor U5987 (N_5987,N_3800,N_2044);
nor U5988 (N_5988,N_3362,N_3048);
and U5989 (N_5989,N_2344,N_3751);
nor U5990 (N_5990,N_3296,N_3663);
nand U5991 (N_5991,N_2679,N_2863);
nand U5992 (N_5992,N_2443,N_3989);
nand U5993 (N_5993,N_3976,N_3853);
nor U5994 (N_5994,N_2019,N_2251);
nor U5995 (N_5995,N_2851,N_2513);
or U5996 (N_5996,N_2184,N_2219);
nand U5997 (N_5997,N_2693,N_3059);
and U5998 (N_5998,N_2285,N_2997);
or U5999 (N_5999,N_2136,N_3932);
or U6000 (N_6000,N_4454,N_5351);
or U6001 (N_6001,N_5319,N_4635);
nand U6002 (N_6002,N_5111,N_4701);
nand U6003 (N_6003,N_4231,N_5030);
or U6004 (N_6004,N_5214,N_4978);
and U6005 (N_6005,N_5082,N_5017);
nor U6006 (N_6006,N_5307,N_4673);
and U6007 (N_6007,N_5436,N_5930);
and U6008 (N_6008,N_5672,N_5509);
or U6009 (N_6009,N_5777,N_5589);
and U6010 (N_6010,N_5202,N_5572);
or U6011 (N_6011,N_4941,N_5187);
nand U6012 (N_6012,N_5485,N_5142);
nor U6013 (N_6013,N_5624,N_4090);
nor U6014 (N_6014,N_5028,N_4161);
or U6015 (N_6015,N_5300,N_5648);
or U6016 (N_6016,N_5623,N_5954);
nor U6017 (N_6017,N_4572,N_4399);
nor U6018 (N_6018,N_4733,N_4084);
and U6019 (N_6019,N_5877,N_4292);
nor U6020 (N_6020,N_5942,N_4177);
nand U6021 (N_6021,N_5128,N_5796);
or U6022 (N_6022,N_4983,N_4883);
nand U6023 (N_6023,N_4312,N_5217);
and U6024 (N_6024,N_4957,N_5753);
nand U6025 (N_6025,N_4287,N_4439);
nand U6026 (N_6026,N_4366,N_4588);
or U6027 (N_6027,N_4008,N_5715);
nor U6028 (N_6028,N_5906,N_4894);
and U6029 (N_6029,N_5296,N_4972);
and U6030 (N_6030,N_4882,N_5940);
nand U6031 (N_6031,N_4423,N_5646);
or U6032 (N_6032,N_4469,N_4269);
nand U6033 (N_6033,N_4089,N_4553);
or U6034 (N_6034,N_5054,N_5491);
and U6035 (N_6035,N_5250,N_5806);
nand U6036 (N_6036,N_4738,N_5680);
or U6037 (N_6037,N_4647,N_5123);
nor U6038 (N_6038,N_4163,N_5075);
or U6039 (N_6039,N_4664,N_4666);
nand U6040 (N_6040,N_5014,N_5630);
nor U6041 (N_6041,N_5546,N_4582);
nor U6042 (N_6042,N_4461,N_4318);
nor U6043 (N_6043,N_4601,N_4911);
nand U6044 (N_6044,N_4115,N_4800);
nand U6045 (N_6045,N_5809,N_4552);
nand U6046 (N_6046,N_4913,N_4153);
nor U6047 (N_6047,N_5769,N_5064);
nand U6048 (N_6048,N_4612,N_4729);
nor U6049 (N_6049,N_5227,N_5074);
nor U6050 (N_6050,N_4736,N_4675);
and U6051 (N_6051,N_5905,N_5944);
nor U6052 (N_6052,N_4880,N_5783);
nand U6053 (N_6053,N_4766,N_4056);
and U6054 (N_6054,N_4573,N_4965);
and U6055 (N_6055,N_4508,N_5695);
nor U6056 (N_6056,N_5342,N_4904);
or U6057 (N_6057,N_5448,N_4191);
nand U6058 (N_6058,N_4719,N_5883);
nor U6059 (N_6059,N_4500,N_5698);
nor U6060 (N_6060,N_5803,N_4422);
nor U6061 (N_6061,N_4174,N_5601);
nor U6062 (N_6062,N_4046,N_5279);
and U6063 (N_6063,N_5941,N_4782);
and U6064 (N_6064,N_4218,N_4967);
nor U6065 (N_6065,N_5470,N_5165);
and U6066 (N_6066,N_5513,N_4614);
nor U6067 (N_6067,N_4406,N_4049);
or U6068 (N_6068,N_4820,N_5405);
nand U6069 (N_6069,N_4827,N_5627);
or U6070 (N_6070,N_5482,N_4328);
or U6071 (N_6071,N_5970,N_5324);
and U6072 (N_6072,N_5357,N_4768);
or U6073 (N_6073,N_5321,N_4438);
and U6074 (N_6074,N_5125,N_5688);
and U6075 (N_6075,N_5552,N_4711);
and U6076 (N_6076,N_4680,N_4309);
nor U6077 (N_6077,N_4129,N_4688);
and U6078 (N_6078,N_5486,N_5330);
nand U6079 (N_6079,N_4630,N_5257);
or U6080 (N_6080,N_4307,N_5558);
nor U6081 (N_6081,N_4565,N_4844);
or U6082 (N_6082,N_4826,N_5718);
or U6083 (N_6083,N_5000,N_5246);
nand U6084 (N_6084,N_5745,N_5443);
and U6085 (N_6085,N_5723,N_4662);
nor U6086 (N_6086,N_5046,N_4367);
nor U6087 (N_6087,N_5761,N_4035);
or U6088 (N_6088,N_4576,N_4808);
nand U6089 (N_6089,N_4502,N_5929);
nor U6090 (N_6090,N_4257,N_5216);
xnor U6091 (N_6091,N_5422,N_5189);
nand U6092 (N_6092,N_5355,N_4943);
and U6093 (N_6093,N_4950,N_5302);
or U6094 (N_6094,N_5754,N_4110);
nand U6095 (N_6095,N_4154,N_4798);
or U6096 (N_6096,N_5069,N_5298);
nor U6097 (N_6097,N_5711,N_5800);
and U6098 (N_6098,N_5099,N_5913);
and U6099 (N_6099,N_4634,N_5760);
or U6100 (N_6100,N_4770,N_5729);
and U6101 (N_6101,N_4494,N_5925);
xnor U6102 (N_6102,N_5036,N_4443);
and U6103 (N_6103,N_4092,N_5713);
nand U6104 (N_6104,N_4258,N_5797);
and U6105 (N_6105,N_5714,N_4044);
and U6106 (N_6106,N_5370,N_4263);
nand U6107 (N_6107,N_5595,N_5038);
nor U6108 (N_6108,N_5466,N_4790);
or U6109 (N_6109,N_5990,N_5684);
and U6110 (N_6110,N_4003,N_4503);
or U6111 (N_6111,N_4128,N_4986);
or U6112 (N_6112,N_5223,N_5742);
nor U6113 (N_6113,N_5037,N_4535);
nor U6114 (N_6114,N_4100,N_5136);
or U6115 (N_6115,N_5040,N_5410);
nand U6116 (N_6116,N_4636,N_5984);
or U6117 (N_6117,N_5171,N_4350);
and U6118 (N_6118,N_4223,N_5577);
nor U6119 (N_6119,N_4984,N_5852);
nor U6120 (N_6120,N_5198,N_5946);
or U6121 (N_6121,N_5219,N_4839);
and U6122 (N_6122,N_5560,N_4465);
or U6123 (N_6123,N_5763,N_5186);
or U6124 (N_6124,N_4294,N_4561);
and U6125 (N_6125,N_5935,N_4053);
nand U6126 (N_6126,N_5519,N_4916);
nand U6127 (N_6127,N_5840,N_4495);
nor U6128 (N_6128,N_4448,N_4834);
or U6129 (N_6129,N_4080,N_4047);
nor U6130 (N_6130,N_4705,N_4183);
nor U6131 (N_6131,N_5467,N_5656);
nor U6132 (N_6132,N_4869,N_5350);
and U6133 (N_6133,N_4681,N_5493);
or U6134 (N_6134,N_5266,N_5620);
or U6135 (N_6135,N_4813,N_4797);
nor U6136 (N_6136,N_5140,N_5662);
nand U6137 (N_6137,N_4109,N_5106);
and U6138 (N_6138,N_4375,N_4382);
nand U6139 (N_6139,N_4818,N_5550);
or U6140 (N_6140,N_5641,N_5093);
or U6141 (N_6141,N_4881,N_4915);
nor U6142 (N_6142,N_4404,N_4173);
nand U6143 (N_6143,N_5559,N_5902);
nand U6144 (N_6144,N_5555,N_4855);
or U6145 (N_6145,N_4569,N_5317);
nand U6146 (N_6146,N_5245,N_4857);
or U6147 (N_6147,N_5933,N_4171);
nor U6148 (N_6148,N_5706,N_4322);
and U6149 (N_6149,N_5308,N_5969);
nand U6150 (N_6150,N_4145,N_5389);
or U6151 (N_6151,N_4156,N_4440);
or U6152 (N_6152,N_4139,N_4268);
nand U6153 (N_6153,N_5091,N_4244);
nor U6154 (N_6154,N_5751,N_4851);
nor U6155 (N_6155,N_5903,N_4725);
nor U6156 (N_6156,N_4335,N_5583);
nand U6157 (N_6157,N_4707,N_4632);
or U6158 (N_6158,N_5653,N_5563);
and U6159 (N_6159,N_5013,N_5599);
or U6160 (N_6160,N_5503,N_5109);
or U6161 (N_6161,N_5784,N_4430);
and U6162 (N_6162,N_4018,N_4906);
nor U6163 (N_6163,N_4302,N_4394);
and U6164 (N_6164,N_5776,N_4124);
or U6165 (N_6165,N_4994,N_5501);
or U6166 (N_6166,N_4274,N_5476);
and U6167 (N_6167,N_4538,N_5561);
nor U6168 (N_6168,N_5158,N_5587);
nor U6169 (N_6169,N_5735,N_5932);
or U6170 (N_6170,N_4026,N_5051);
nand U6171 (N_6171,N_5786,N_5462);
nand U6172 (N_6172,N_4743,N_4284);
nand U6173 (N_6173,N_4849,N_5739);
nor U6174 (N_6174,N_5295,N_5256);
nor U6175 (N_6175,N_4618,N_4695);
nand U6176 (N_6176,N_5766,N_4871);
nand U6177 (N_6177,N_4400,N_4932);
or U6178 (N_6178,N_4667,N_5135);
and U6179 (N_6179,N_5384,N_5269);
or U6180 (N_6180,N_4720,N_4956);
nor U6181 (N_6181,N_5849,N_4980);
nor U6182 (N_6182,N_4964,N_4151);
and U6183 (N_6183,N_5669,N_5965);
and U6184 (N_6184,N_5282,N_5149);
nor U6185 (N_6185,N_4353,N_4391);
nand U6186 (N_6186,N_4023,N_4126);
and U6187 (N_6187,N_5886,N_4387);
or U6188 (N_6188,N_4106,N_4165);
nor U6189 (N_6189,N_4504,N_4989);
and U6190 (N_6190,N_4401,N_4337);
nor U6191 (N_6191,N_5571,N_5248);
nor U6192 (N_6192,N_5237,N_5768);
nand U6193 (N_6193,N_4144,N_4352);
nor U6194 (N_6194,N_5170,N_4033);
or U6195 (N_6195,N_5178,N_5318);
nor U6196 (N_6196,N_5221,N_4160);
and U6197 (N_6197,N_5566,N_5438);
or U6198 (N_6198,N_4641,N_4928);
nor U6199 (N_6199,N_5774,N_5162);
nor U6200 (N_6200,N_5673,N_5831);
or U6201 (N_6201,N_5041,N_5077);
nand U6202 (N_6202,N_4922,N_4319);
nand U6203 (N_6203,N_4425,N_5072);
or U6204 (N_6204,N_4193,N_5353);
or U6205 (N_6205,N_5825,N_4088);
nand U6206 (N_6206,N_4606,N_5594);
or U6207 (N_6207,N_4463,N_4396);
and U6208 (N_6208,N_4010,N_4246);
nor U6209 (N_6209,N_4131,N_4655);
nand U6210 (N_6210,N_5144,N_4155);
and U6211 (N_6211,N_4096,N_5474);
nor U6212 (N_6212,N_4537,N_5525);
and U6213 (N_6213,N_4359,N_4093);
and U6214 (N_6214,N_5315,N_4698);
or U6215 (N_6215,N_5376,N_4806);
nand U6216 (N_6216,N_4361,N_5987);
nor U6217 (N_6217,N_4501,N_5968);
or U6218 (N_6218,N_4686,N_4764);
and U6219 (N_6219,N_4013,N_4188);
or U6220 (N_6220,N_4012,N_5701);
and U6221 (N_6221,N_4543,N_5081);
nor U6222 (N_6222,N_5161,N_4933);
nand U6223 (N_6223,N_5616,N_5471);
nor U6224 (N_6224,N_4282,N_4142);
and U6225 (N_6225,N_5327,N_4479);
and U6226 (N_6226,N_4817,N_5129);
nand U6227 (N_6227,N_5749,N_4584);
and U6228 (N_6228,N_5048,N_4771);
and U6229 (N_6229,N_5110,N_5844);
and U6230 (N_6230,N_5868,N_4952);
or U6231 (N_6231,N_5645,N_4509);
nand U6232 (N_6232,N_5116,N_5687);
or U6233 (N_6233,N_5131,N_5240);
xnor U6234 (N_6234,N_4838,N_4371);
or U6235 (N_6235,N_4311,N_5105);
and U6236 (N_6236,N_5640,N_5365);
nand U6237 (N_6237,N_5708,N_5450);
nor U6238 (N_6238,N_4549,N_5272);
or U6239 (N_6239,N_4276,N_5615);
or U6240 (N_6240,N_5455,N_5130);
nand U6241 (N_6241,N_4671,N_5948);
nand U6242 (N_6242,N_5591,N_5690);
nor U6243 (N_6243,N_4007,N_4592);
nor U6244 (N_6244,N_4973,N_4858);
nor U6245 (N_6245,N_5702,N_5409);
nand U6246 (N_6246,N_5311,N_4819);
and U6247 (N_6247,N_5132,N_4583);
nand U6248 (N_6248,N_5988,N_5523);
nor U6249 (N_6249,N_5704,N_5372);
and U6250 (N_6250,N_5452,N_5277);
or U6251 (N_6251,N_5460,N_4296);
and U6252 (N_6252,N_4714,N_5520);
nor U6253 (N_6253,N_4314,N_5085);
or U6254 (N_6254,N_5575,N_4365);
or U6255 (N_6255,N_4853,N_5312);
nor U6256 (N_6256,N_4393,N_4867);
and U6257 (N_6257,N_5710,N_5526);
or U6258 (N_6258,N_5992,N_4987);
or U6259 (N_6259,N_4531,N_4214);
or U6260 (N_6260,N_5395,N_5454);
nand U6261 (N_6261,N_5562,N_4321);
nor U6262 (N_6262,N_4968,N_4014);
xnor U6263 (N_6263,N_4364,N_4703);
nand U6264 (N_6264,N_5744,N_5117);
nor U6265 (N_6265,N_5169,N_4187);
and U6266 (N_6266,N_4640,N_4863);
nand U6267 (N_6267,N_4101,N_5795);
nand U6268 (N_6268,N_4105,N_4997);
or U6269 (N_6269,N_4574,N_4029);
or U6270 (N_6270,N_5088,N_4992);
or U6271 (N_6271,N_5733,N_4324);
or U6272 (N_6272,N_5408,N_4488);
or U6273 (N_6273,N_4578,N_5604);
or U6274 (N_6274,N_4402,N_4937);
nand U6275 (N_6275,N_5549,N_4643);
and U6276 (N_6276,N_4716,N_5943);
nor U6277 (N_6277,N_4250,N_5107);
or U6278 (N_6278,N_4134,N_4814);
nor U6279 (N_6279,N_5885,N_4642);
nand U6280 (N_6280,N_5811,N_4627);
and U6281 (N_6281,N_4985,N_5382);
or U6282 (N_6282,N_5752,N_5524);
nand U6283 (N_6283,N_5586,N_5507);
nand U6284 (N_6284,N_5606,N_5912);
and U6285 (N_6285,N_5412,N_5021);
nor U6286 (N_6286,N_4095,N_5530);
and U6287 (N_6287,N_4613,N_4555);
nand U6288 (N_6288,N_5071,N_5204);
or U6289 (N_6289,N_5334,N_5755);
or U6290 (N_6290,N_4830,N_4498);
and U6291 (N_6291,N_5705,N_4718);
nor U6292 (N_6292,N_4854,N_4953);
and U6293 (N_6293,N_5335,N_5757);
nand U6294 (N_6294,N_4758,N_5445);
and U6295 (N_6295,N_4433,N_4521);
or U6296 (N_6296,N_4021,N_5772);
nand U6297 (N_6297,N_5537,N_5114);
or U6298 (N_6298,N_4836,N_5540);
nand U6299 (N_6299,N_5226,N_4037);
nor U6300 (N_6300,N_4386,N_5638);
or U6301 (N_6301,N_5456,N_4575);
nor U6302 (N_6302,N_4694,N_4082);
nor U6303 (N_6303,N_4807,N_5398);
and U6304 (N_6304,N_4467,N_5090);
or U6305 (N_6305,N_5590,N_4777);
and U6306 (N_6306,N_4330,N_5995);
nor U6307 (N_6307,N_4947,N_4946);
and U6308 (N_6308,N_5846,N_5926);
nor U6309 (N_6309,N_4708,N_5593);
or U6310 (N_6310,N_4672,N_5344);
nand U6311 (N_6311,N_4757,N_4068);
nor U6312 (N_6312,N_4169,N_4377);
nor U6313 (N_6313,N_5481,N_5651);
or U6314 (N_6314,N_4840,N_4484);
nand U6315 (N_6315,N_5104,N_4852);
or U6316 (N_6316,N_4270,N_4510);
or U6317 (N_6317,N_5251,N_5238);
and U6318 (N_6318,N_4963,N_4259);
and U6319 (N_6319,N_5665,N_4186);
and U6320 (N_6320,N_5893,N_4629);
nand U6321 (N_6321,N_5841,N_5862);
nand U6322 (N_6322,N_5889,N_5773);
nand U6323 (N_6323,N_5832,N_5947);
or U6324 (N_6324,N_4991,N_4735);
nand U6325 (N_6325,N_4104,N_4256);
nor U6326 (N_6326,N_4437,N_4000);
nand U6327 (N_6327,N_4842,N_4114);
nand U6328 (N_6328,N_4823,N_4480);
and U6329 (N_6329,N_5386,N_5057);
and U6330 (N_6330,N_4083,N_5998);
or U6331 (N_6331,N_4924,N_5492);
and U6332 (N_6332,N_5961,N_4732);
or U6333 (N_6333,N_4248,N_4179);
or U6334 (N_6334,N_4076,N_4930);
or U6335 (N_6335,N_4125,N_4526);
and U6336 (N_6336,N_5950,N_4455);
nand U6337 (N_6337,N_5053,N_4310);
or U6338 (N_6338,N_4597,N_5336);
and U6339 (N_6339,N_5819,N_5290);
nand U6340 (N_6340,N_4625,N_4682);
nand U6341 (N_6341,N_4513,N_4519);
nand U6342 (N_6342,N_4477,N_5024);
and U6343 (N_6343,N_5461,N_5789);
nand U6344 (N_6344,N_4816,N_4317);
and U6345 (N_6345,N_4343,N_5956);
or U6346 (N_6346,N_4648,N_4334);
nand U6347 (N_6347,N_4988,N_5346);
nand U6348 (N_6348,N_4559,N_5477);
or U6349 (N_6349,N_4293,N_4656);
and U6350 (N_6350,N_4492,N_5010);
nor U6351 (N_6351,N_4301,N_5859);
nor U6352 (N_6352,N_4219,N_4379);
or U6353 (N_6353,N_4976,N_5876);
and U6354 (N_6354,N_5804,N_4031);
nand U6355 (N_6355,N_4247,N_5097);
nor U6356 (N_6356,N_5428,N_5576);
and U6357 (N_6357,N_5887,N_5531);
nor U6358 (N_6358,N_5514,N_5029);
nand U6359 (N_6359,N_4590,N_4347);
or U6360 (N_6360,N_4748,N_5447);
or U6361 (N_6361,N_5817,N_5741);
and U6362 (N_6362,N_5652,N_4299);
and U6363 (N_6363,N_4547,N_5660);
and U6364 (N_6364,N_4271,N_5830);
or U6365 (N_6365,N_5378,N_4692);
nand U6366 (N_6366,N_5360,N_4679);
and U6367 (N_6367,N_5532,N_4772);
and U6368 (N_6368,N_4658,N_5195);
nor U6369 (N_6369,N_4742,N_4897);
nor U6370 (N_6370,N_4579,N_4712);
nand U6371 (N_6371,N_5473,N_5855);
and U6372 (N_6372,N_5596,N_5047);
or U6373 (N_6373,N_4593,N_5115);
or U6374 (N_6374,N_5921,N_5100);
or U6375 (N_6375,N_5442,N_4570);
and U6376 (N_6376,N_4344,N_4390);
nand U6377 (N_6377,N_4661,N_5818);
nor U6378 (N_6378,N_4039,N_4810);
nor U6379 (N_6379,N_5904,N_5626);
or U6380 (N_6380,N_4229,N_4357);
nor U6381 (N_6381,N_5260,N_4087);
nand U6382 (N_6382,N_4620,N_4242);
and U6383 (N_6383,N_4690,N_4192);
nor U6384 (N_6384,N_4870,N_5345);
or U6385 (N_6385,N_4385,N_4407);
or U6386 (N_6386,N_4801,N_4704);
nand U6387 (N_6387,N_4336,N_5391);
nand U6388 (N_6388,N_4607,N_4460);
or U6389 (N_6389,N_5668,N_4949);
nor U6390 (N_6390,N_5720,N_5693);
nand U6391 (N_6391,N_4812,N_4907);
nor U6392 (N_6392,N_5083,N_4756);
nand U6393 (N_6393,N_5339,N_4594);
nand U6394 (N_6394,N_5895,N_5553);
and U6395 (N_6395,N_4760,N_5610);
or U6396 (N_6396,N_4048,N_4489);
or U6397 (N_6397,N_4684,N_4064);
nand U6398 (N_6398,N_4241,N_4623);
and U6399 (N_6399,N_4700,N_4558);
and U6400 (N_6400,N_4586,N_4527);
nor U6401 (N_6401,N_4159,N_5018);
nand U6402 (N_6402,N_5647,N_5670);
nor U6403 (N_6403,N_4138,N_5451);
or U6404 (N_6404,N_5247,N_5043);
or U6405 (N_6405,N_4787,N_4468);
or U6406 (N_6406,N_5617,N_5964);
and U6407 (N_6407,N_5896,N_5120);
and U6408 (N_6408,N_5612,N_4472);
and U6409 (N_6409,N_4740,N_4283);
nand U6410 (N_6410,N_5898,N_5025);
nor U6411 (N_6411,N_4753,N_4079);
or U6412 (N_6412,N_4539,N_4912);
and U6413 (N_6413,N_4333,N_5629);
nor U6414 (N_6414,N_4659,N_5813);
nor U6415 (N_6415,N_4195,N_4428);
nand U6416 (N_6416,N_4966,N_5242);
xnor U6417 (N_6417,N_4074,N_5827);
or U6418 (N_6418,N_4075,N_5609);
nor U6419 (N_6419,N_5799,N_4567);
nor U6420 (N_6420,N_4320,N_5347);
nor U6421 (N_6421,N_5001,N_5417);
nand U6422 (N_6422,N_5363,N_4773);
and U6423 (N_6423,N_5967,N_4544);
or U6424 (N_6424,N_4693,N_4602);
and U6425 (N_6425,N_4493,N_4427);
or U6426 (N_6426,N_4847,N_4297);
and U6427 (N_6427,N_4751,N_4774);
or U6428 (N_6428,N_5991,N_5368);
and U6429 (N_6429,N_5325,N_4197);
nor U6430 (N_6430,N_5249,N_4358);
and U6431 (N_6431,N_4085,N_4470);
nand U6432 (N_6432,N_4696,N_4435);
or U6433 (N_6433,N_5734,N_5802);
or U6434 (N_6434,N_4646,N_4122);
or U6435 (N_6435,N_5848,N_4886);
nand U6436 (N_6436,N_4132,N_4875);
and U6437 (N_6437,N_5654,N_5557);
or U6438 (N_6438,N_5139,N_4215);
and U6439 (N_6439,N_4009,N_4341);
nor U6440 (N_6440,N_4081,N_5194);
or U6441 (N_6441,N_5015,N_5483);
or U6442 (N_6442,N_5413,N_4563);
nor U6443 (N_6443,N_4568,N_5999);
and U6444 (N_6444,N_4890,N_4405);
or U6445 (N_6445,N_4354,N_4133);
nand U6446 (N_6446,N_4529,N_4554);
nor U6447 (N_6447,N_4449,N_4213);
and U6448 (N_6448,N_4644,N_4058);
nand U6449 (N_6449,N_4560,N_4731);
or U6450 (N_6450,N_4859,N_5027);
nand U6451 (N_6451,N_5419,N_5108);
and U6452 (N_6452,N_5243,N_5996);
or U6453 (N_6453,N_4415,N_5976);
and U6454 (N_6454,N_5966,N_5686);
nand U6455 (N_6455,N_4117,N_5529);
and U6456 (N_6456,N_4522,N_5955);
nand U6457 (N_6457,N_5890,N_4065);
and U6458 (N_6458,N_5078,N_5499);
or U6459 (N_6459,N_4184,N_4212);
or U6460 (N_6460,N_4650,N_4887);
nor U6461 (N_6461,N_5369,N_5439);
or U6462 (N_6462,N_4196,N_5565);
nand U6463 (N_6463,N_4868,N_5835);
nor U6464 (N_6464,N_4776,N_4622);
and U6465 (N_6465,N_5118,N_4045);
or U6466 (N_6466,N_5418,N_5922);
nand U6467 (N_6467,N_5758,N_4715);
nand U6468 (N_6468,N_5354,N_5518);
or U6469 (N_6469,N_4861,N_5607);
nand U6470 (N_6470,N_5914,N_5547);
or U6471 (N_6471,N_5821,N_5511);
nand U6472 (N_6472,N_5127,N_5124);
or U6473 (N_6473,N_4811,N_4363);
or U6474 (N_6474,N_5387,N_5842);
and U6475 (N_6475,N_5393,N_5231);
or U6476 (N_6476,N_5736,N_5023);
nor U6477 (N_6477,N_4279,N_5193);
or U6478 (N_6478,N_5502,N_4392);
nor U6479 (N_6479,N_5756,N_4119);
and U6480 (N_6480,N_5801,N_5103);
nor U6481 (N_6481,N_5267,N_5009);
and U6482 (N_6482,N_4471,N_4030);
and U6483 (N_6483,N_5039,N_5810);
and U6484 (N_6484,N_4864,N_5314);
and U6485 (N_6485,N_5084,N_5978);
or U6486 (N_6486,N_5602,N_5423);
or U6487 (N_6487,N_5605,N_4541);
nand U6488 (N_6488,N_4595,N_4638);
nand U6489 (N_6489,N_5878,N_4918);
and U6490 (N_6490,N_4621,N_5076);
nand U6491 (N_6491,N_5006,N_5092);
and U6492 (N_6492,N_4243,N_4238);
xnor U6493 (N_6493,N_5847,N_4722);
or U6494 (N_6494,N_5642,N_4403);
nand U6495 (N_6495,N_5164,N_5993);
or U6496 (N_6496,N_5068,N_5960);
nand U6497 (N_6497,N_4608,N_5425);
or U6498 (N_6498,N_5341,N_4452);
nor U6499 (N_6499,N_5121,N_5934);
nand U6500 (N_6500,N_4977,N_4042);
nand U6501 (N_6501,N_5407,N_5163);
and U6502 (N_6502,N_5233,N_4931);
nand U6503 (N_6503,N_5899,N_4099);
or U6504 (N_6504,N_4604,N_4762);
nand U6505 (N_6505,N_5578,N_5432);
nand U6506 (N_6506,N_4028,N_4670);
or U6507 (N_6507,N_4668,N_5181);
or U6508 (N_6508,N_5853,N_5177);
nand U6509 (N_6509,N_5263,N_4611);
and U6510 (N_6510,N_5618,N_5138);
or U6511 (N_6511,N_5176,N_5230);
nand U6512 (N_6512,N_4262,N_4216);
and U6513 (N_6513,N_5707,N_5264);
nor U6514 (N_6514,N_4167,N_5157);
and U6515 (N_6515,N_4895,N_4550);
or U6516 (N_6516,N_5820,N_5147);
or U6517 (N_6517,N_5725,N_4038);
nand U6518 (N_6518,N_4744,N_4410);
or U6519 (N_6519,N_5065,N_5206);
nand U6520 (N_6520,N_4252,N_4856);
xor U6521 (N_6521,N_5180,N_4888);
and U6522 (N_6522,N_5936,N_4442);
or U6523 (N_6523,N_4524,N_4874);
and U6524 (N_6524,N_5611,N_5495);
nand U6525 (N_6525,N_4893,N_5631);
nor U6526 (N_6526,N_4118,N_4198);
nand U6527 (N_6527,N_5528,N_4837);
nand U6528 (N_6528,N_5380,N_4860);
nor U6529 (N_6529,N_5457,N_4032);
nor U6530 (N_6530,N_4349,N_5244);
nand U6531 (N_6531,N_5910,N_4373);
nand U6532 (N_6532,N_4203,N_5854);
nand U6533 (N_6533,N_5567,N_4290);
nor U6534 (N_6534,N_4954,N_4723);
and U6535 (N_6535,N_4665,N_5861);
nor U6536 (N_6536,N_5086,N_5340);
xor U6537 (N_6537,N_4057,N_4829);
and U6538 (N_6538,N_5649,N_4233);
nor U6539 (N_6539,N_4749,N_5621);
or U6540 (N_6540,N_5717,N_4441);
or U6541 (N_6541,N_5167,N_5112);
and U6542 (N_6542,N_4228,N_4651);
or U6543 (N_6543,N_4189,N_4657);
or U6544 (N_6544,N_5031,N_4609);
nand U6545 (N_6545,N_4157,N_5468);
or U6546 (N_6546,N_5287,N_4355);
nor U6547 (N_6547,N_5915,N_5533);
and U6548 (N_6548,N_5371,N_4434);
and U6549 (N_6549,N_4424,N_4591);
nand U6550 (N_6550,N_4793,N_4306);
and U6551 (N_6551,N_4205,N_5401);
nor U6552 (N_6552,N_4767,N_4927);
nor U6553 (N_6553,N_4945,N_4209);
or U6554 (N_6554,N_4398,N_4780);
nand U6555 (N_6555,N_5728,N_4211);
nand U6556 (N_6556,N_4958,N_4451);
and U6557 (N_6557,N_5446,N_5814);
nand U6558 (N_6558,N_5431,N_5488);
and U6559 (N_6559,N_5681,N_4974);
and U6560 (N_6560,N_4962,N_4063);
and U6561 (N_6561,N_5002,N_4397);
or U6562 (N_6562,N_5900,N_5016);
xnor U6563 (N_6563,N_5603,N_4687);
nand U6564 (N_6564,N_4530,N_4898);
nor U6565 (N_6565,N_5663,N_5433);
or U6566 (N_6566,N_5174,N_5959);
and U6567 (N_6567,N_5166,N_5962);
and U6568 (N_6568,N_5892,N_4796);
or U6569 (N_6569,N_5592,N_4896);
and U6570 (N_6570,N_4017,N_4717);
or U6571 (N_6571,N_5538,N_5726);
and U6572 (N_6572,N_5880,N_5866);
and U6573 (N_6573,N_4548,N_5367);
nand U6574 (N_6574,N_4135,N_5437);
nand U6575 (N_6575,N_4411,N_5032);
and U6576 (N_6576,N_5326,N_5207);
or U6577 (N_6577,N_4605,N_5508);
or U6578 (N_6578,N_4990,N_5301);
nor U6579 (N_6579,N_5544,N_5348);
nand U6580 (N_6580,N_4305,N_5600);
or U6581 (N_6581,N_5148,N_4123);
nand U6582 (N_6582,N_5424,N_5985);
nor U6583 (N_6583,N_5496,N_4027);
and U6584 (N_6584,N_4267,N_5160);
or U6585 (N_6585,N_4475,N_4878);
xnor U6586 (N_6586,N_5211,N_4523);
or U6587 (N_6587,N_4417,N_5285);
and U6588 (N_6588,N_5958,N_4781);
nor U6589 (N_6589,N_4281,N_4051);
nor U6590 (N_6590,N_5977,N_5535);
nor U6591 (N_6591,N_5812,N_4254);
or U6592 (N_6592,N_5901,N_4204);
nor U6593 (N_6593,N_5050,N_5919);
nand U6594 (N_6594,N_4727,N_4077);
nor U6595 (N_6595,N_4086,N_4208);
nor U6596 (N_6596,N_4520,N_4217);
and U6597 (N_6597,N_4409,N_5404);
nor U6598 (N_6598,N_4663,N_5212);
and U6599 (N_6599,N_4815,N_5504);
nor U6600 (N_6600,N_5435,N_4865);
nand U6601 (N_6601,N_5808,N_5657);
nor U6602 (N_6602,N_5034,N_4413);
or U6603 (N_6603,N_5062,N_4936);
nand U6604 (N_6604,N_5270,N_5983);
and U6605 (N_6605,N_5044,N_5570);
and U6606 (N_6606,N_4226,N_5724);
nor U6607 (N_6607,N_4062,N_4395);
or U6608 (N_6608,N_4778,N_4164);
or U6609 (N_6609,N_4070,N_4466);
nand U6610 (N_6610,N_5542,N_5971);
and U6611 (N_6611,N_5719,N_4802);
and U6612 (N_6612,N_5597,N_4002);
or U6613 (N_6613,N_4408,N_5505);
nor U6614 (N_6614,N_5920,N_5218);
or U6615 (N_6615,N_5882,N_5056);
and U6616 (N_6616,N_5699,N_4737);
and U6617 (N_6617,N_5033,N_4649);
or U6618 (N_6618,N_4289,N_4069);
nand U6619 (N_6619,N_5215,N_4342);
or U6620 (N_6620,N_5273,N_5779);
and U6621 (N_6621,N_5917,N_5639);
nor U6622 (N_6622,N_4619,N_4514);
and U6623 (N_6623,N_4181,N_5667);
nand U6624 (N_6624,N_5727,N_4224);
nor U6625 (N_6625,N_4674,N_4929);
or U6626 (N_6626,N_5888,N_4516);
nor U6627 (N_6627,N_5781,N_4239);
nor U6628 (N_6628,N_5323,N_5986);
or U6629 (N_6629,N_5721,N_4506);
and U6630 (N_6630,N_4872,N_4710);
nand U6631 (N_6631,N_4534,N_5487);
nor U6632 (N_6632,N_5328,N_5585);
nor U6633 (N_6633,N_5937,N_5343);
and U6634 (N_6634,N_5337,N_5201);
nand U6635 (N_6635,N_4482,N_4066);
or U6636 (N_6636,N_5792,N_5373);
and U6637 (N_6637,N_4308,N_5952);
and U6638 (N_6638,N_5145,N_4459);
nand U6639 (N_6639,N_4825,N_5356);
or U6640 (N_6640,N_5239,N_5304);
or U6641 (N_6641,N_5703,N_5767);
nor U6642 (N_6642,N_5512,N_5891);
nor U6643 (N_6643,N_5333,N_5635);
and U6644 (N_6644,N_5510,N_4022);
and U6645 (N_6645,N_5632,N_5659);
nor U6646 (N_6646,N_4331,N_5498);
or U6647 (N_6647,N_4730,N_4295);
nand U6648 (N_6648,N_4136,N_4709);
nor U6649 (N_6649,N_5063,N_4901);
nand U6650 (N_6650,N_4446,N_5141);
nor U6651 (N_6651,N_4788,N_5869);
nand U6652 (N_6652,N_4277,N_4822);
and U6653 (N_6653,N_5478,N_5780);
and U6654 (N_6654,N_4420,N_5856);
nand U6655 (N_6655,N_5625,N_5923);
nor U6656 (N_6656,N_5283,N_5358);
nand U6657 (N_6657,N_5782,N_5850);
nand U6658 (N_6658,N_5884,N_4143);
and U6659 (N_6659,N_5143,N_4304);
and U6660 (N_6660,N_4345,N_4381);
nand U6661 (N_6661,N_5822,N_5951);
and U6662 (N_6662,N_4848,N_4168);
nand U6663 (N_6663,N_5793,N_5516);
and U6664 (N_6664,N_5008,N_5716);
nor U6665 (N_6665,N_4982,N_5490);
or U6666 (N_6666,N_5975,N_4564);
nand U6667 (N_6667,N_4585,N_5070);
or U6668 (N_6668,N_4706,N_5205);
and U6669 (N_6669,N_4789,N_4598);
nor U6670 (N_6670,N_5989,N_5305);
nand U6671 (N_6671,N_5329,N_5838);
or U6672 (N_6672,N_4036,N_5402);
or U6673 (N_6673,N_5133,N_5479);
nor U6674 (N_6674,N_5865,N_5541);
nand U6675 (N_6675,N_4795,N_5210);
and U6676 (N_6676,N_4517,N_4255);
nand U6677 (N_6677,N_4511,N_5430);
nor U6678 (N_6678,N_4019,N_5153);
and U6679 (N_6679,N_4747,N_5388);
and U6680 (N_6680,N_4266,N_5361);
nor U6681 (N_6681,N_5527,N_4016);
or U6682 (N_6682,N_4006,N_5172);
nor U6683 (N_6683,N_4097,N_4914);
and U6684 (N_6684,N_4616,N_5192);
xnor U6685 (N_6685,N_5750,N_4889);
and U6686 (N_6686,N_4626,N_4236);
nor U6687 (N_6687,N_5472,N_4562);
nor U6688 (N_6688,N_4993,N_4102);
and U6689 (N_6689,N_4505,N_5894);
nor U6690 (N_6690,N_4478,N_5582);
nor U6691 (N_6691,N_4877,N_4275);
nand U6692 (N_6692,N_4199,N_5175);
nand U6693 (N_6693,N_4995,N_4999);
nor U6694 (N_6694,N_5199,N_5643);
nor U6695 (N_6695,N_4338,N_4507);
and U6696 (N_6696,N_4546,N_4923);
and U6697 (N_6697,N_4291,N_5834);
nand U6698 (N_6698,N_5152,N_4955);
nand U6699 (N_6699,N_5857,N_5564);
nor U6700 (N_6700,N_5265,N_5685);
nand U6701 (N_6701,N_4152,N_5924);
or U6702 (N_6702,N_5291,N_5377);
nor U6703 (N_6703,N_5297,N_5982);
nand U6704 (N_6704,N_5870,N_5981);
and U6705 (N_6705,N_4975,N_5183);
or U6706 (N_6706,N_4261,N_4805);
nand U6707 (N_6707,N_4685,N_5522);
nor U6708 (N_6708,N_5286,N_4542);
nor U6709 (N_6709,N_5119,N_4792);
nor U6710 (N_6710,N_5155,N_5458);
and U6711 (N_6711,N_5484,N_5190);
nand U6712 (N_6712,N_4754,N_5689);
and U6713 (N_6713,N_5449,N_5633);
nand U6714 (N_6714,N_5255,N_4775);
nand U6715 (N_6715,N_4491,N_5258);
or U6716 (N_6716,N_4245,N_5200);
or U6717 (N_6717,N_4264,N_4628);
or U6718 (N_6718,N_5203,N_4515);
nand U6719 (N_6719,N_5332,N_4368);
or U6720 (N_6720,N_4746,N_5765);
nand U6721 (N_6721,N_4525,N_4934);
nand U6722 (N_6722,N_5634,N_4721);
or U6723 (N_6723,N_5262,N_4416);
nor U6724 (N_6724,N_5775,N_4610);
or U6725 (N_6725,N_5785,N_4024);
or U6726 (N_6726,N_5979,N_4702);
or U6727 (N_6727,N_5379,N_4112);
xor U6728 (N_6728,N_4447,N_5274);
nor U6729 (N_6729,N_4938,N_5494);
or U6730 (N_6730,N_5052,N_4220);
or U6731 (N_6731,N_5534,N_5939);
nor U6732 (N_6732,N_5392,N_5588);
or U6733 (N_6733,N_5289,N_4456);
nand U6734 (N_6734,N_5220,N_5364);
and U6735 (N_6735,N_5731,N_4175);
or U6736 (N_6736,N_5427,N_4786);
and U6737 (N_6737,N_4374,N_4388);
nand U6738 (N_6738,N_4348,N_4891);
and U6739 (N_6739,N_4221,N_4919);
nand U6740 (N_6740,N_5692,N_4326);
xor U6741 (N_6741,N_4551,N_5788);
nor U6742 (N_6742,N_4278,N_5661);
nor U6743 (N_6743,N_4828,N_5837);
and U6744 (N_6744,N_4652,N_4900);
or U6745 (N_6745,N_5875,N_4249);
and U6746 (N_6746,N_5349,N_4998);
nor U6747 (N_6747,N_4288,N_4925);
nand U6748 (N_6748,N_5310,N_4020);
or U6749 (N_6749,N_5464,N_4235);
or U6750 (N_6750,N_5916,N_4948);
and U6751 (N_6751,N_4362,N_5580);
nand U6752 (N_6752,N_4908,N_5581);
and U6753 (N_6753,N_5406,N_5738);
and U6754 (N_6754,N_4265,N_4540);
and U6755 (N_6755,N_4879,N_4779);
nor U6756 (N_6756,N_5399,N_4824);
or U6757 (N_6757,N_4108,N_5396);
and U6758 (N_6758,N_5536,N_4316);
and U6759 (N_6759,N_5909,N_5949);
nor U6760 (N_6760,N_4713,N_4436);
nor U6761 (N_6761,N_4060,N_5826);
nand U6762 (N_6762,N_5026,N_5927);
nand U6763 (N_6763,N_5222,N_4981);
nand U6764 (N_6764,N_4785,N_5058);
nand U6765 (N_6765,N_4745,N_5864);
nor U6766 (N_6766,N_4286,N_5208);
nand U6767 (N_6767,N_4496,N_4166);
or U6768 (N_6768,N_5622,N_5500);
nor U6769 (N_6769,N_5957,N_5150);
or U6770 (N_6770,N_5292,N_4315);
nor U6771 (N_6771,N_5415,N_4412);
and U6772 (N_6772,N_5762,N_5235);
or U6773 (N_6773,N_5213,N_4130);
nand U6774 (N_6774,N_4873,N_4835);
nand U6775 (N_6775,N_4346,N_4884);
or U6776 (N_6776,N_5911,N_4536);
nand U6777 (N_6777,N_4182,N_5815);
nand U6778 (N_6778,N_5280,N_5453);
or U6779 (N_6779,N_5322,N_4426);
nand U6780 (N_6780,N_5366,N_4617);
nand U6781 (N_6781,N_5677,N_5381);
or U6782 (N_6782,N_5628,N_5126);
and U6783 (N_6783,N_5022,N_4728);
or U6784 (N_6784,N_4285,N_5778);
nor U6785 (N_6785,N_5113,N_4841);
nor U6786 (N_6786,N_4765,N_5020);
nand U6787 (N_6787,N_4926,N_4909);
nand U6788 (N_6788,N_5918,N_5012);
nor U6789 (N_6789,N_5475,N_5066);
nor U6790 (N_6790,N_5151,N_4678);
nor U6791 (N_6791,N_4432,N_5182);
or U6792 (N_6792,N_4783,N_4339);
and U6793 (N_6793,N_5805,N_4951);
or U6794 (N_6794,N_5790,N_4624);
xor U6795 (N_6795,N_4116,N_5374);
nand U6796 (N_6796,N_5569,N_5228);
and U6797 (N_6797,N_5650,N_5055);
and U6798 (N_6798,N_5049,N_5209);
and U6799 (N_6799,N_5241,N_4207);
and U6800 (N_6800,N_5907,N_5421);
and U6801 (N_6801,N_5737,N_4935);
and U6802 (N_6802,N_5764,N_4303);
or U6803 (N_6803,N_5463,N_5675);
nand U6804 (N_6804,N_4683,N_4921);
nand U6805 (N_6805,N_5945,N_5871);
nor U6806 (N_6806,N_4149,N_5833);
or U6807 (N_6807,N_5824,N_4111);
nor U6808 (N_6808,N_4577,N_5191);
nor U6809 (N_6809,N_4959,N_5096);
nor U6810 (N_6810,N_5881,N_4799);
or U6811 (N_6811,N_4944,N_4232);
nor U6812 (N_6812,N_4653,N_4376);
nand U6813 (N_6813,N_5574,N_4571);
nand U6814 (N_6814,N_4689,N_4004);
nor U6815 (N_6815,N_4759,N_5694);
nand U6816 (N_6816,N_4676,N_5791);
and U6817 (N_6817,N_4699,N_4421);
and U6818 (N_6818,N_5679,N_4589);
or U6819 (N_6819,N_4025,N_5288);
or U6820 (N_6820,N_4141,N_4078);
nand U6821 (N_6821,N_5007,N_4091);
nand U6822 (N_6822,N_4389,N_4833);
and U6823 (N_6823,N_5568,N_4137);
and U6824 (N_6824,N_4098,N_4862);
and U6825 (N_6825,N_5179,N_5188);
nor U6826 (N_6826,N_4015,N_5953);
or U6827 (N_6827,N_4356,N_5963);
and U6828 (N_6828,N_5658,N_4061);
nand U6829 (N_6829,N_5746,N_5271);
and U6830 (N_6830,N_4158,N_4180);
nand U6831 (N_6831,N_5416,N_5444);
and U6832 (N_6832,N_5845,N_5434);
or U6833 (N_6833,N_4190,N_5497);
or U6834 (N_6834,N_5489,N_4474);
or U6835 (N_6835,N_4639,N_4734);
nor U6836 (N_6836,N_5042,N_4327);
and U6837 (N_6837,N_4240,N_5506);
and U6838 (N_6838,N_4418,N_5816);
nand U6839 (N_6839,N_4486,N_4121);
and U6840 (N_6840,N_5173,N_5275);
or U6841 (N_6841,N_5515,N_4444);
and U6842 (N_6842,N_4910,N_5732);
nor U6843 (N_6843,N_5197,N_5863);
nor U6844 (N_6844,N_5697,N_4794);
or U6845 (N_6845,N_5666,N_5712);
nor U6846 (N_6846,N_4654,N_4809);
or U6847 (N_6847,N_5281,N_5897);
nand U6848 (N_6848,N_5928,N_5383);
nor U6849 (N_6849,N_5872,N_5168);
nor U6850 (N_6850,N_4059,N_4615);
nor U6851 (N_6851,N_4481,N_5067);
nand U6852 (N_6852,N_4172,N_4940);
nand U6853 (N_6853,N_5159,N_4313);
and U6854 (N_6854,N_5759,N_4769);
nand U6855 (N_6855,N_4969,N_4939);
nor U6856 (N_6856,N_4581,N_4419);
nand U6857 (N_6857,N_5545,N_5613);
and U6858 (N_6858,N_4556,N_4846);
nor U6859 (N_6859,N_4518,N_4580);
or U6860 (N_6860,N_5730,N_5974);
or U6861 (N_6861,N_5655,N_5134);
nand U6862 (N_6862,N_5309,N_4724);
or U6863 (N_6863,N_5867,N_4073);
and U6864 (N_6864,N_5060,N_5259);
or U6865 (N_6865,N_5122,N_5644);
nand U6866 (N_6866,N_5299,N_4763);
nor U6867 (N_6867,N_4378,N_4148);
nand U6868 (N_6868,N_4761,N_4476);
nand U6869 (N_6869,N_5554,N_5843);
nand U6870 (N_6870,N_5860,N_4041);
nor U6871 (N_6871,N_5087,N_4512);
or U6872 (N_6872,N_4210,N_5671);
nand U6873 (N_6873,N_4885,N_5254);
nor U6874 (N_6874,N_4201,N_5441);
and U6875 (N_6875,N_4850,N_5858);
nand U6876 (N_6876,N_4637,N_4034);
and U6877 (N_6877,N_5798,N_4237);
nand U6878 (N_6878,N_4821,N_4660);
or U6879 (N_6879,N_4113,N_5614);
and U6880 (N_6880,N_5411,N_5480);
nand U6881 (N_6881,N_5154,N_4831);
and U6882 (N_6882,N_5787,N_5839);
nand U6883 (N_6883,N_5094,N_4645);
nor U6884 (N_6884,N_4633,N_4323);
nand U6885 (N_6885,N_4431,N_4260);
nor U6886 (N_6886,N_4001,N_5390);
and U6887 (N_6887,N_5972,N_5224);
and U6888 (N_6888,N_5338,N_5551);
and U6889 (N_6889,N_4631,N_5873);
nand U6890 (N_6890,N_4380,N_5185);
nor U6891 (N_6891,N_5080,N_5584);
nand U6892 (N_6892,N_5823,N_5696);
and U6893 (N_6893,N_4445,N_5747);
nor U6894 (N_6894,N_5836,N_4803);
nor U6895 (N_6895,N_4600,N_5748);
or U6896 (N_6896,N_4603,N_4230);
and U6897 (N_6897,N_5019,N_4325);
nor U6898 (N_6898,N_4369,N_5556);
nand U6899 (N_6899,N_4253,N_4845);
and U6900 (N_6900,N_4804,N_5973);
or U6901 (N_6901,N_5543,N_4464);
or U6902 (N_6902,N_5980,N_4457);
or U6903 (N_6903,N_5252,N_4185);
nor U6904 (N_6904,N_5517,N_5579);
nor U6905 (N_6905,N_5306,N_4566);
nor U6906 (N_6906,N_5003,N_5059);
or U6907 (N_6907,N_5521,N_4202);
or U6908 (N_6908,N_4429,N_4052);
or U6909 (N_6909,N_4485,N_4227);
or U6910 (N_6910,N_4458,N_5011);
nand U6911 (N_6911,N_5851,N_4146);
nor U6912 (N_6912,N_4487,N_5362);
and U6913 (N_6913,N_5375,N_5938);
nand U6914 (N_6914,N_4194,N_5089);
and U6915 (N_6915,N_5225,N_4739);
nor U6916 (N_6916,N_5229,N_4866);
or U6917 (N_6917,N_4979,N_4750);
nor U6918 (N_6918,N_4120,N_5156);
nand U6919 (N_6919,N_4370,N_4726);
and U6920 (N_6920,N_5676,N_4905);
nand U6921 (N_6921,N_4225,N_5740);
nor U6922 (N_6922,N_4040,N_5102);
nor U6923 (N_6923,N_4162,N_5548);
and U6924 (N_6924,N_5459,N_5722);
nand U6925 (N_6925,N_5637,N_4055);
or U6926 (N_6926,N_4483,N_4072);
nor U6927 (N_6927,N_5709,N_5619);
or U6928 (N_6928,N_5931,N_4340);
nor U6929 (N_6929,N_4067,N_5440);
or U6930 (N_6930,N_5268,N_4222);
and U6931 (N_6931,N_5146,N_5828);
or U6932 (N_6932,N_5400,N_4054);
nand U6933 (N_6933,N_5469,N_4043);
nor U6934 (N_6934,N_4587,N_4942);
nor U6935 (N_6935,N_4533,N_4677);
and U6936 (N_6936,N_5184,N_4791);
and U6937 (N_6937,N_4329,N_5294);
nor U6938 (N_6938,N_5874,N_4920);
nor U6939 (N_6939,N_5278,N_5101);
and U6940 (N_6940,N_4752,N_4545);
and U6941 (N_6941,N_4251,N_5004);
nor U6942 (N_6942,N_5682,N_4497);
or U6943 (N_6943,N_5683,N_5829);
and U6944 (N_6944,N_4273,N_5770);
nor U6945 (N_6945,N_5079,N_4383);
nor U6946 (N_6946,N_4050,N_4917);
nand U6947 (N_6947,N_5994,N_4970);
nand U6948 (N_6948,N_5234,N_4170);
nor U6949 (N_6949,N_4200,N_5261);
and U6950 (N_6950,N_5678,N_5539);
nand U6951 (N_6951,N_4490,N_4902);
nor U6952 (N_6952,N_5807,N_4669);
nand U6953 (N_6953,N_5385,N_5232);
nor U6954 (N_6954,N_5331,N_4961);
nand U6955 (N_6955,N_5313,N_4094);
nor U6956 (N_6956,N_4103,N_5664);
nand U6957 (N_6957,N_5303,N_4532);
and U6958 (N_6958,N_5293,N_5253);
nand U6959 (N_6959,N_5397,N_4450);
and U6960 (N_6960,N_4755,N_5691);
nand U6961 (N_6961,N_5394,N_5236);
nor U6962 (N_6962,N_4372,N_5061);
and U6963 (N_6963,N_5196,N_4005);
nand U6964 (N_6964,N_4599,N_4899);
nand U6965 (N_6965,N_4697,N_5997);
nor U6966 (N_6966,N_4360,N_4499);
nand U6967 (N_6967,N_5045,N_5879);
nor U6968 (N_6968,N_4528,N_5403);
and U6969 (N_6969,N_4272,N_5573);
nand U6970 (N_6970,N_5794,N_4298);
and U6971 (N_6971,N_5095,N_4107);
nand U6972 (N_6972,N_4234,N_5420);
nand U6973 (N_6973,N_5465,N_5598);
nor U6974 (N_6974,N_5137,N_4453);
nor U6975 (N_6975,N_4903,N_4876);
or U6976 (N_6976,N_4332,N_4206);
nand U6977 (N_6977,N_4741,N_4960);
and U6978 (N_6978,N_4140,N_5284);
nand U6979 (N_6979,N_4971,N_5414);
or U6980 (N_6980,N_4280,N_4071);
nor U6981 (N_6981,N_5359,N_5700);
and U6982 (N_6982,N_5035,N_4127);
nor U6983 (N_6983,N_4178,N_4011);
and U6984 (N_6984,N_4176,N_4147);
nor U6985 (N_6985,N_4892,N_5908);
nand U6986 (N_6986,N_4832,N_5276);
and U6987 (N_6987,N_4596,N_4557);
nand U6988 (N_6988,N_5674,N_4462);
or U6989 (N_6989,N_5098,N_5316);
and U6990 (N_6990,N_5743,N_5608);
nand U6991 (N_6991,N_4351,N_4300);
nor U6992 (N_6992,N_5005,N_5426);
nor U6993 (N_6993,N_4414,N_4784);
and U6994 (N_6994,N_5429,N_5771);
and U6995 (N_6995,N_4384,N_4996);
and U6996 (N_6996,N_5320,N_4150);
nor U6997 (N_6997,N_4843,N_4473);
nand U6998 (N_6998,N_5073,N_4691);
or U6999 (N_6999,N_5636,N_5352);
or U7000 (N_7000,N_4804,N_5817);
and U7001 (N_7001,N_5911,N_4821);
nor U7002 (N_7002,N_5630,N_4797);
and U7003 (N_7003,N_5406,N_5694);
nor U7004 (N_7004,N_5415,N_5324);
nor U7005 (N_7005,N_5036,N_5321);
nor U7006 (N_7006,N_5578,N_4110);
or U7007 (N_7007,N_4151,N_4434);
nor U7008 (N_7008,N_4124,N_5308);
or U7009 (N_7009,N_5803,N_5697);
nand U7010 (N_7010,N_4483,N_4933);
or U7011 (N_7011,N_5165,N_5818);
and U7012 (N_7012,N_4587,N_5277);
and U7013 (N_7013,N_4593,N_4565);
and U7014 (N_7014,N_5622,N_4172);
or U7015 (N_7015,N_4237,N_4455);
nand U7016 (N_7016,N_4767,N_4678);
nor U7017 (N_7017,N_4657,N_4087);
or U7018 (N_7018,N_5597,N_4057);
or U7019 (N_7019,N_4794,N_4529);
or U7020 (N_7020,N_4833,N_5142);
nand U7021 (N_7021,N_5443,N_5656);
nand U7022 (N_7022,N_4957,N_5340);
nand U7023 (N_7023,N_4635,N_5556);
nor U7024 (N_7024,N_5061,N_4294);
and U7025 (N_7025,N_5315,N_5557);
and U7026 (N_7026,N_5697,N_5912);
nor U7027 (N_7027,N_4177,N_4245);
nand U7028 (N_7028,N_4474,N_4031);
and U7029 (N_7029,N_4126,N_4746);
and U7030 (N_7030,N_4569,N_4662);
or U7031 (N_7031,N_4799,N_5453);
or U7032 (N_7032,N_4478,N_5103);
and U7033 (N_7033,N_4086,N_5030);
nand U7034 (N_7034,N_5078,N_5645);
or U7035 (N_7035,N_5456,N_5803);
nor U7036 (N_7036,N_5875,N_4373);
nand U7037 (N_7037,N_4761,N_4154);
nand U7038 (N_7038,N_5637,N_5974);
or U7039 (N_7039,N_5888,N_5141);
and U7040 (N_7040,N_4823,N_5816);
or U7041 (N_7041,N_4914,N_5480);
nor U7042 (N_7042,N_5271,N_5750);
or U7043 (N_7043,N_4870,N_4858);
nand U7044 (N_7044,N_5583,N_5858);
and U7045 (N_7045,N_4860,N_4726);
and U7046 (N_7046,N_4332,N_5692);
nand U7047 (N_7047,N_5286,N_4321);
or U7048 (N_7048,N_4256,N_4093);
or U7049 (N_7049,N_5189,N_4004);
or U7050 (N_7050,N_5713,N_4692);
and U7051 (N_7051,N_4232,N_5798);
nand U7052 (N_7052,N_5667,N_4173);
and U7053 (N_7053,N_4797,N_5887);
or U7054 (N_7054,N_4230,N_4857);
nor U7055 (N_7055,N_4114,N_4392);
and U7056 (N_7056,N_5720,N_4911);
and U7057 (N_7057,N_4195,N_5615);
nand U7058 (N_7058,N_4648,N_5235);
and U7059 (N_7059,N_5983,N_5681);
nand U7060 (N_7060,N_5600,N_5427);
nand U7061 (N_7061,N_5801,N_4661);
nor U7062 (N_7062,N_5698,N_5408);
and U7063 (N_7063,N_4620,N_5686);
and U7064 (N_7064,N_5653,N_5844);
nand U7065 (N_7065,N_4823,N_5284);
or U7066 (N_7066,N_5601,N_4055);
xor U7067 (N_7067,N_5703,N_4461);
nand U7068 (N_7068,N_4053,N_4756);
nand U7069 (N_7069,N_5716,N_4724);
nor U7070 (N_7070,N_4196,N_5090);
nand U7071 (N_7071,N_5342,N_5812);
and U7072 (N_7072,N_4459,N_5641);
or U7073 (N_7073,N_5570,N_5479);
or U7074 (N_7074,N_5182,N_5117);
and U7075 (N_7075,N_5547,N_4132);
and U7076 (N_7076,N_4820,N_4718);
nand U7077 (N_7077,N_5060,N_5751);
nand U7078 (N_7078,N_5860,N_4075);
nor U7079 (N_7079,N_5846,N_4703);
or U7080 (N_7080,N_5693,N_4249);
nand U7081 (N_7081,N_4261,N_4260);
nor U7082 (N_7082,N_5718,N_5724);
and U7083 (N_7083,N_4681,N_4407);
nor U7084 (N_7084,N_4172,N_4517);
nor U7085 (N_7085,N_5102,N_4024);
and U7086 (N_7086,N_5711,N_5004);
nor U7087 (N_7087,N_4824,N_4382);
nor U7088 (N_7088,N_5456,N_4009);
nor U7089 (N_7089,N_4669,N_5645);
nor U7090 (N_7090,N_4121,N_4186);
nand U7091 (N_7091,N_5069,N_4733);
or U7092 (N_7092,N_4331,N_4042);
or U7093 (N_7093,N_5677,N_4529);
nand U7094 (N_7094,N_4332,N_4215);
and U7095 (N_7095,N_4855,N_5283);
and U7096 (N_7096,N_4760,N_5197);
and U7097 (N_7097,N_4973,N_5913);
and U7098 (N_7098,N_4423,N_4656);
nor U7099 (N_7099,N_5633,N_5131);
nand U7100 (N_7100,N_5103,N_4161);
or U7101 (N_7101,N_4729,N_4272);
and U7102 (N_7102,N_5673,N_5213);
xor U7103 (N_7103,N_4632,N_5234);
nand U7104 (N_7104,N_5067,N_5996);
nor U7105 (N_7105,N_5299,N_4579);
or U7106 (N_7106,N_5839,N_4234);
nor U7107 (N_7107,N_4033,N_4715);
nor U7108 (N_7108,N_5829,N_4888);
or U7109 (N_7109,N_4326,N_4242);
nor U7110 (N_7110,N_5207,N_4922);
and U7111 (N_7111,N_4688,N_4951);
and U7112 (N_7112,N_4705,N_5774);
nor U7113 (N_7113,N_4814,N_4149);
nand U7114 (N_7114,N_4972,N_4221);
or U7115 (N_7115,N_4695,N_5570);
nor U7116 (N_7116,N_5985,N_5958);
and U7117 (N_7117,N_5593,N_5242);
and U7118 (N_7118,N_4371,N_4125);
or U7119 (N_7119,N_5283,N_5745);
nor U7120 (N_7120,N_5455,N_5968);
or U7121 (N_7121,N_4214,N_4974);
or U7122 (N_7122,N_4019,N_5750);
nand U7123 (N_7123,N_5525,N_5656);
nand U7124 (N_7124,N_4808,N_5172);
and U7125 (N_7125,N_5146,N_4697);
and U7126 (N_7126,N_4323,N_4522);
nand U7127 (N_7127,N_4106,N_5680);
nand U7128 (N_7128,N_4830,N_5184);
nor U7129 (N_7129,N_4274,N_5710);
nand U7130 (N_7130,N_4968,N_4466);
nand U7131 (N_7131,N_4083,N_5340);
nand U7132 (N_7132,N_5756,N_4417);
and U7133 (N_7133,N_5920,N_4639);
nand U7134 (N_7134,N_5552,N_5784);
nand U7135 (N_7135,N_5134,N_5021);
or U7136 (N_7136,N_4561,N_4486);
or U7137 (N_7137,N_5918,N_5741);
or U7138 (N_7138,N_4304,N_5836);
and U7139 (N_7139,N_5107,N_5434);
xnor U7140 (N_7140,N_5897,N_5501);
nand U7141 (N_7141,N_5343,N_4301);
nor U7142 (N_7142,N_5105,N_4916);
nor U7143 (N_7143,N_5609,N_5503);
and U7144 (N_7144,N_4720,N_4113);
or U7145 (N_7145,N_5376,N_5311);
and U7146 (N_7146,N_5620,N_4153);
nor U7147 (N_7147,N_5633,N_4705);
xnor U7148 (N_7148,N_5908,N_4142);
or U7149 (N_7149,N_4577,N_5944);
nand U7150 (N_7150,N_5035,N_5571);
nor U7151 (N_7151,N_5294,N_5595);
nand U7152 (N_7152,N_5502,N_4073);
or U7153 (N_7153,N_4437,N_4941);
or U7154 (N_7154,N_5985,N_5709);
or U7155 (N_7155,N_4895,N_5359);
nand U7156 (N_7156,N_4732,N_5446);
and U7157 (N_7157,N_5250,N_4211);
and U7158 (N_7158,N_5622,N_4825);
or U7159 (N_7159,N_4630,N_4491);
and U7160 (N_7160,N_4447,N_5648);
and U7161 (N_7161,N_4802,N_4810);
or U7162 (N_7162,N_5661,N_4406);
and U7163 (N_7163,N_5408,N_5361);
or U7164 (N_7164,N_4297,N_4054);
nor U7165 (N_7165,N_4575,N_5591);
or U7166 (N_7166,N_4755,N_5751);
or U7167 (N_7167,N_4985,N_5162);
nor U7168 (N_7168,N_4309,N_5017);
nor U7169 (N_7169,N_4785,N_4351);
nand U7170 (N_7170,N_5880,N_4290);
or U7171 (N_7171,N_4455,N_5662);
nor U7172 (N_7172,N_4067,N_5370);
or U7173 (N_7173,N_4983,N_4276);
or U7174 (N_7174,N_4667,N_4341);
nor U7175 (N_7175,N_5207,N_4118);
or U7176 (N_7176,N_4593,N_4159);
or U7177 (N_7177,N_4712,N_4499);
or U7178 (N_7178,N_5964,N_4493);
or U7179 (N_7179,N_5235,N_4417);
nand U7180 (N_7180,N_4451,N_5171);
or U7181 (N_7181,N_5757,N_5506);
or U7182 (N_7182,N_4236,N_4927);
nand U7183 (N_7183,N_5589,N_5535);
nor U7184 (N_7184,N_5582,N_5319);
nand U7185 (N_7185,N_4308,N_4009);
nand U7186 (N_7186,N_5055,N_4035);
nor U7187 (N_7187,N_5852,N_5355);
nand U7188 (N_7188,N_5693,N_5100);
and U7189 (N_7189,N_4642,N_4539);
and U7190 (N_7190,N_5936,N_5947);
nor U7191 (N_7191,N_4596,N_5322);
or U7192 (N_7192,N_5035,N_5505);
nand U7193 (N_7193,N_5258,N_4084);
and U7194 (N_7194,N_5591,N_4593);
nor U7195 (N_7195,N_4857,N_4696);
nor U7196 (N_7196,N_5799,N_4036);
or U7197 (N_7197,N_5427,N_5036);
and U7198 (N_7198,N_4319,N_5157);
nand U7199 (N_7199,N_5255,N_4522);
nand U7200 (N_7200,N_4199,N_4876);
or U7201 (N_7201,N_5291,N_5927);
nor U7202 (N_7202,N_5342,N_4097);
or U7203 (N_7203,N_5632,N_5239);
nand U7204 (N_7204,N_5817,N_4924);
or U7205 (N_7205,N_4272,N_5974);
nand U7206 (N_7206,N_5851,N_4835);
nand U7207 (N_7207,N_5336,N_4751);
and U7208 (N_7208,N_5540,N_4208);
nand U7209 (N_7209,N_5957,N_4029);
nand U7210 (N_7210,N_4151,N_5853);
nor U7211 (N_7211,N_5174,N_5590);
nor U7212 (N_7212,N_5223,N_5563);
nor U7213 (N_7213,N_4912,N_4998);
nor U7214 (N_7214,N_4024,N_4149);
or U7215 (N_7215,N_5671,N_4297);
nand U7216 (N_7216,N_4704,N_4545);
or U7217 (N_7217,N_4577,N_5254);
or U7218 (N_7218,N_5705,N_4971);
nand U7219 (N_7219,N_5067,N_4473);
nand U7220 (N_7220,N_4432,N_5902);
nand U7221 (N_7221,N_5758,N_5772);
nor U7222 (N_7222,N_5562,N_5639);
nor U7223 (N_7223,N_5494,N_5929);
nor U7224 (N_7224,N_5763,N_4233);
nand U7225 (N_7225,N_5159,N_5363);
and U7226 (N_7226,N_4635,N_4526);
and U7227 (N_7227,N_5497,N_5603);
or U7228 (N_7228,N_5000,N_4239);
and U7229 (N_7229,N_5054,N_5252);
or U7230 (N_7230,N_5327,N_5156);
nand U7231 (N_7231,N_4461,N_4402);
nand U7232 (N_7232,N_5811,N_5986);
nand U7233 (N_7233,N_5999,N_4116);
and U7234 (N_7234,N_5344,N_4317);
or U7235 (N_7235,N_5462,N_4267);
xnor U7236 (N_7236,N_5597,N_5412);
or U7237 (N_7237,N_4903,N_4685);
and U7238 (N_7238,N_4369,N_4852);
or U7239 (N_7239,N_5402,N_4781);
nand U7240 (N_7240,N_5663,N_4769);
nand U7241 (N_7241,N_5845,N_5397);
nor U7242 (N_7242,N_4331,N_4792);
or U7243 (N_7243,N_5521,N_5894);
nor U7244 (N_7244,N_4702,N_4640);
nand U7245 (N_7245,N_5501,N_5982);
or U7246 (N_7246,N_4953,N_5932);
or U7247 (N_7247,N_4806,N_4100);
nor U7248 (N_7248,N_4472,N_5574);
or U7249 (N_7249,N_4802,N_4177);
nor U7250 (N_7250,N_5420,N_5585);
and U7251 (N_7251,N_4857,N_4034);
nand U7252 (N_7252,N_4210,N_5141);
and U7253 (N_7253,N_5223,N_4799);
nor U7254 (N_7254,N_5004,N_4747);
or U7255 (N_7255,N_5077,N_5342);
and U7256 (N_7256,N_5141,N_4882);
and U7257 (N_7257,N_4560,N_5749);
and U7258 (N_7258,N_4890,N_5109);
and U7259 (N_7259,N_5390,N_5460);
nor U7260 (N_7260,N_5972,N_5713);
nand U7261 (N_7261,N_5851,N_5573);
nor U7262 (N_7262,N_5801,N_5751);
nor U7263 (N_7263,N_5663,N_5395);
nand U7264 (N_7264,N_5365,N_5785);
nand U7265 (N_7265,N_4517,N_5507);
or U7266 (N_7266,N_5182,N_4721);
nor U7267 (N_7267,N_5805,N_5150);
nand U7268 (N_7268,N_4571,N_4876);
nand U7269 (N_7269,N_4379,N_4083);
nor U7270 (N_7270,N_4740,N_4960);
nor U7271 (N_7271,N_4804,N_5111);
and U7272 (N_7272,N_5062,N_5036);
or U7273 (N_7273,N_4998,N_5340);
or U7274 (N_7274,N_5750,N_4740);
nor U7275 (N_7275,N_5116,N_5182);
or U7276 (N_7276,N_4255,N_4708);
and U7277 (N_7277,N_4127,N_4640);
nand U7278 (N_7278,N_5176,N_5408);
nand U7279 (N_7279,N_5281,N_5567);
or U7280 (N_7280,N_4342,N_4929);
nor U7281 (N_7281,N_5593,N_4010);
and U7282 (N_7282,N_5017,N_4124);
or U7283 (N_7283,N_4498,N_5278);
nor U7284 (N_7284,N_4931,N_5350);
nand U7285 (N_7285,N_4100,N_5194);
nand U7286 (N_7286,N_5874,N_5677);
and U7287 (N_7287,N_4079,N_4994);
nand U7288 (N_7288,N_4689,N_5414);
or U7289 (N_7289,N_4699,N_4455);
nor U7290 (N_7290,N_5381,N_5000);
and U7291 (N_7291,N_4873,N_5359);
nor U7292 (N_7292,N_4649,N_5750);
nor U7293 (N_7293,N_5342,N_5326);
and U7294 (N_7294,N_4530,N_5480);
and U7295 (N_7295,N_4453,N_5879);
nor U7296 (N_7296,N_5537,N_5338);
nand U7297 (N_7297,N_5671,N_5035);
nand U7298 (N_7298,N_4173,N_5946);
and U7299 (N_7299,N_5875,N_5043);
nor U7300 (N_7300,N_4191,N_5198);
or U7301 (N_7301,N_4892,N_4158);
nand U7302 (N_7302,N_4936,N_4617);
or U7303 (N_7303,N_5487,N_4503);
nand U7304 (N_7304,N_5527,N_4823);
nor U7305 (N_7305,N_5809,N_5142);
nand U7306 (N_7306,N_4445,N_4302);
or U7307 (N_7307,N_5397,N_4340);
or U7308 (N_7308,N_4811,N_4180);
or U7309 (N_7309,N_5240,N_5860);
or U7310 (N_7310,N_5804,N_4382);
or U7311 (N_7311,N_5358,N_4946);
and U7312 (N_7312,N_4501,N_5497);
nor U7313 (N_7313,N_5896,N_5521);
and U7314 (N_7314,N_5121,N_5267);
nor U7315 (N_7315,N_5905,N_5051);
nand U7316 (N_7316,N_5959,N_4923);
nor U7317 (N_7317,N_4606,N_4494);
nor U7318 (N_7318,N_4127,N_5762);
and U7319 (N_7319,N_4739,N_5449);
and U7320 (N_7320,N_5148,N_5414);
nand U7321 (N_7321,N_4584,N_4645);
nor U7322 (N_7322,N_5173,N_5918);
nand U7323 (N_7323,N_5588,N_5476);
nor U7324 (N_7324,N_5169,N_5973);
nor U7325 (N_7325,N_5765,N_4766);
or U7326 (N_7326,N_4849,N_4344);
nor U7327 (N_7327,N_4261,N_4364);
nor U7328 (N_7328,N_5033,N_5324);
or U7329 (N_7329,N_5216,N_5780);
and U7330 (N_7330,N_5836,N_5043);
nor U7331 (N_7331,N_5931,N_5914);
nand U7332 (N_7332,N_5154,N_5391);
nand U7333 (N_7333,N_5331,N_5929);
and U7334 (N_7334,N_5027,N_5739);
and U7335 (N_7335,N_4928,N_4880);
or U7336 (N_7336,N_4029,N_5111);
nor U7337 (N_7337,N_4381,N_4707);
and U7338 (N_7338,N_4036,N_4454);
nor U7339 (N_7339,N_4790,N_4113);
and U7340 (N_7340,N_5703,N_5823);
nor U7341 (N_7341,N_5755,N_5560);
or U7342 (N_7342,N_5287,N_4518);
nor U7343 (N_7343,N_4075,N_4453);
nand U7344 (N_7344,N_4050,N_5015);
nor U7345 (N_7345,N_5243,N_5718);
or U7346 (N_7346,N_5307,N_5667);
and U7347 (N_7347,N_4499,N_5805);
nor U7348 (N_7348,N_5430,N_4066);
and U7349 (N_7349,N_4230,N_5398);
and U7350 (N_7350,N_4045,N_5465);
nand U7351 (N_7351,N_4361,N_4319);
and U7352 (N_7352,N_5592,N_5223);
and U7353 (N_7353,N_4511,N_4605);
nand U7354 (N_7354,N_5815,N_4222);
nor U7355 (N_7355,N_4660,N_5205);
or U7356 (N_7356,N_5975,N_4355);
xor U7357 (N_7357,N_5317,N_4295);
or U7358 (N_7358,N_4619,N_4845);
and U7359 (N_7359,N_4725,N_5596);
nand U7360 (N_7360,N_5967,N_4989);
nand U7361 (N_7361,N_5938,N_4016);
and U7362 (N_7362,N_4896,N_5886);
and U7363 (N_7363,N_4044,N_5788);
nand U7364 (N_7364,N_4184,N_5925);
nand U7365 (N_7365,N_4597,N_4221);
or U7366 (N_7366,N_5726,N_4170);
nor U7367 (N_7367,N_4048,N_4031);
or U7368 (N_7368,N_5417,N_5916);
or U7369 (N_7369,N_5460,N_4564);
nand U7370 (N_7370,N_5019,N_4969);
nand U7371 (N_7371,N_4072,N_4001);
nand U7372 (N_7372,N_5895,N_4067);
or U7373 (N_7373,N_5323,N_5488);
or U7374 (N_7374,N_4513,N_4174);
nand U7375 (N_7375,N_5431,N_5444);
and U7376 (N_7376,N_5216,N_5213);
or U7377 (N_7377,N_5389,N_4103);
nor U7378 (N_7378,N_4041,N_4101);
and U7379 (N_7379,N_4780,N_4746);
nand U7380 (N_7380,N_5600,N_5099);
nand U7381 (N_7381,N_5053,N_5776);
or U7382 (N_7382,N_5436,N_5466);
nand U7383 (N_7383,N_5975,N_5004);
nand U7384 (N_7384,N_5165,N_4758);
nor U7385 (N_7385,N_5206,N_5302);
nand U7386 (N_7386,N_4969,N_5962);
nand U7387 (N_7387,N_4183,N_4808);
nand U7388 (N_7388,N_4733,N_4277);
nor U7389 (N_7389,N_4067,N_4811);
nand U7390 (N_7390,N_4389,N_5306);
and U7391 (N_7391,N_4207,N_5100);
and U7392 (N_7392,N_4281,N_5826);
or U7393 (N_7393,N_5375,N_5336);
nor U7394 (N_7394,N_5615,N_4426);
or U7395 (N_7395,N_5864,N_4666);
nor U7396 (N_7396,N_5562,N_5039);
nor U7397 (N_7397,N_5279,N_5428);
or U7398 (N_7398,N_4142,N_5929);
and U7399 (N_7399,N_4903,N_5354);
or U7400 (N_7400,N_4292,N_5415);
and U7401 (N_7401,N_4413,N_4504);
nand U7402 (N_7402,N_4068,N_4155);
or U7403 (N_7403,N_4534,N_5762);
nand U7404 (N_7404,N_5351,N_4634);
or U7405 (N_7405,N_4783,N_5397);
and U7406 (N_7406,N_5663,N_5363);
and U7407 (N_7407,N_4739,N_4208);
nand U7408 (N_7408,N_4507,N_4511);
or U7409 (N_7409,N_4105,N_5282);
and U7410 (N_7410,N_4595,N_5195);
or U7411 (N_7411,N_5289,N_4679);
xnor U7412 (N_7412,N_4558,N_5769);
nor U7413 (N_7413,N_5322,N_5605);
nand U7414 (N_7414,N_4058,N_4498);
and U7415 (N_7415,N_5658,N_4155);
nand U7416 (N_7416,N_4546,N_5987);
nor U7417 (N_7417,N_4559,N_5390);
nor U7418 (N_7418,N_5830,N_4423);
and U7419 (N_7419,N_4709,N_4372);
nor U7420 (N_7420,N_5231,N_5743);
nor U7421 (N_7421,N_5188,N_4436);
nand U7422 (N_7422,N_4807,N_5769);
or U7423 (N_7423,N_4471,N_4476);
and U7424 (N_7424,N_5224,N_5703);
or U7425 (N_7425,N_5869,N_5053);
and U7426 (N_7426,N_4592,N_5386);
nand U7427 (N_7427,N_5441,N_5911);
nand U7428 (N_7428,N_4067,N_4204);
and U7429 (N_7429,N_5694,N_4051);
nand U7430 (N_7430,N_5100,N_4730);
xnor U7431 (N_7431,N_4068,N_5178);
nor U7432 (N_7432,N_5614,N_4198);
and U7433 (N_7433,N_4688,N_4228);
or U7434 (N_7434,N_5404,N_4372);
or U7435 (N_7435,N_4706,N_4100);
and U7436 (N_7436,N_4492,N_4173);
or U7437 (N_7437,N_4648,N_5924);
nor U7438 (N_7438,N_4381,N_5215);
and U7439 (N_7439,N_4452,N_5024);
or U7440 (N_7440,N_5679,N_5834);
nor U7441 (N_7441,N_5189,N_5997);
and U7442 (N_7442,N_4681,N_4511);
nand U7443 (N_7443,N_5946,N_4911);
or U7444 (N_7444,N_4061,N_4103);
and U7445 (N_7445,N_5535,N_4737);
or U7446 (N_7446,N_4027,N_5788);
nand U7447 (N_7447,N_5305,N_5323);
nand U7448 (N_7448,N_4373,N_4662);
nor U7449 (N_7449,N_4586,N_4839);
nand U7450 (N_7450,N_4992,N_5635);
nand U7451 (N_7451,N_5602,N_5198);
and U7452 (N_7452,N_5525,N_5559);
nor U7453 (N_7453,N_5502,N_4055);
and U7454 (N_7454,N_5410,N_5216);
nand U7455 (N_7455,N_4700,N_5911);
nand U7456 (N_7456,N_4591,N_5934);
nor U7457 (N_7457,N_4107,N_4649);
nor U7458 (N_7458,N_5701,N_5237);
nor U7459 (N_7459,N_5791,N_4198);
nand U7460 (N_7460,N_5354,N_5964);
or U7461 (N_7461,N_4245,N_4949);
nand U7462 (N_7462,N_4106,N_5181);
nand U7463 (N_7463,N_4627,N_4620);
and U7464 (N_7464,N_5412,N_4066);
and U7465 (N_7465,N_4853,N_5175);
and U7466 (N_7466,N_4680,N_5639);
nand U7467 (N_7467,N_4785,N_4721);
nor U7468 (N_7468,N_5580,N_5254);
xor U7469 (N_7469,N_5308,N_4169);
nand U7470 (N_7470,N_5526,N_4939);
nor U7471 (N_7471,N_4848,N_5719);
nor U7472 (N_7472,N_4516,N_5816);
nor U7473 (N_7473,N_5283,N_5732);
nand U7474 (N_7474,N_5025,N_4502);
and U7475 (N_7475,N_4933,N_4672);
nor U7476 (N_7476,N_4420,N_5133);
nand U7477 (N_7477,N_4529,N_4601);
and U7478 (N_7478,N_5788,N_4453);
nor U7479 (N_7479,N_4359,N_5427);
nand U7480 (N_7480,N_5381,N_5241);
or U7481 (N_7481,N_4808,N_5975);
or U7482 (N_7482,N_5910,N_4247);
nand U7483 (N_7483,N_5045,N_4718);
nor U7484 (N_7484,N_5143,N_4581);
nand U7485 (N_7485,N_5691,N_5942);
nand U7486 (N_7486,N_4089,N_4339);
nand U7487 (N_7487,N_5273,N_4703);
and U7488 (N_7488,N_5386,N_5460);
and U7489 (N_7489,N_5181,N_5802);
nor U7490 (N_7490,N_5759,N_5861);
or U7491 (N_7491,N_4122,N_4363);
nor U7492 (N_7492,N_4868,N_4585);
nand U7493 (N_7493,N_5187,N_5983);
nand U7494 (N_7494,N_5283,N_5584);
or U7495 (N_7495,N_5780,N_4377);
nand U7496 (N_7496,N_5314,N_4122);
and U7497 (N_7497,N_4234,N_4151);
and U7498 (N_7498,N_5578,N_4094);
nor U7499 (N_7499,N_5767,N_5660);
and U7500 (N_7500,N_4369,N_4301);
nand U7501 (N_7501,N_5458,N_4930);
nand U7502 (N_7502,N_4890,N_4075);
nor U7503 (N_7503,N_4962,N_4560);
or U7504 (N_7504,N_5636,N_5119);
nand U7505 (N_7505,N_4464,N_4610);
and U7506 (N_7506,N_5499,N_4368);
or U7507 (N_7507,N_4804,N_5352);
or U7508 (N_7508,N_4932,N_4491);
nor U7509 (N_7509,N_5922,N_4460);
or U7510 (N_7510,N_4839,N_4538);
and U7511 (N_7511,N_4536,N_5693);
nand U7512 (N_7512,N_4072,N_4114);
or U7513 (N_7513,N_5030,N_4186);
or U7514 (N_7514,N_4291,N_4018);
or U7515 (N_7515,N_4073,N_5220);
nor U7516 (N_7516,N_5915,N_5159);
or U7517 (N_7517,N_5001,N_4523);
nand U7518 (N_7518,N_4437,N_5419);
or U7519 (N_7519,N_4576,N_5939);
or U7520 (N_7520,N_4794,N_4327);
and U7521 (N_7521,N_5910,N_4928);
or U7522 (N_7522,N_4853,N_4169);
and U7523 (N_7523,N_4780,N_5882);
or U7524 (N_7524,N_5145,N_5047);
and U7525 (N_7525,N_5524,N_5605);
nor U7526 (N_7526,N_5474,N_5177);
and U7527 (N_7527,N_4228,N_5744);
and U7528 (N_7528,N_4149,N_4417);
or U7529 (N_7529,N_5557,N_5011);
nor U7530 (N_7530,N_4621,N_4727);
and U7531 (N_7531,N_5988,N_5540);
and U7532 (N_7532,N_4418,N_5135);
or U7533 (N_7533,N_4667,N_4833);
and U7534 (N_7534,N_4224,N_5772);
nor U7535 (N_7535,N_4152,N_5874);
nand U7536 (N_7536,N_5907,N_4931);
or U7537 (N_7537,N_4361,N_4362);
nand U7538 (N_7538,N_4849,N_4183);
and U7539 (N_7539,N_4729,N_5121);
nor U7540 (N_7540,N_5464,N_4572);
nor U7541 (N_7541,N_5458,N_5224);
nor U7542 (N_7542,N_4642,N_4728);
or U7543 (N_7543,N_4742,N_5036);
nor U7544 (N_7544,N_5862,N_5461);
nor U7545 (N_7545,N_4231,N_5043);
or U7546 (N_7546,N_5239,N_5852);
nor U7547 (N_7547,N_4691,N_4002);
and U7548 (N_7548,N_5752,N_5049);
nor U7549 (N_7549,N_5465,N_5389);
or U7550 (N_7550,N_4316,N_5721);
and U7551 (N_7551,N_4442,N_5595);
nand U7552 (N_7552,N_5469,N_4691);
or U7553 (N_7553,N_4734,N_5409);
or U7554 (N_7554,N_5226,N_4796);
or U7555 (N_7555,N_5065,N_5637);
nand U7556 (N_7556,N_5903,N_4678);
nor U7557 (N_7557,N_4458,N_5059);
xnor U7558 (N_7558,N_4590,N_5964);
nor U7559 (N_7559,N_4791,N_4128);
nor U7560 (N_7560,N_4210,N_4881);
and U7561 (N_7561,N_5395,N_4387);
or U7562 (N_7562,N_5749,N_4603);
nand U7563 (N_7563,N_4607,N_4873);
nand U7564 (N_7564,N_5574,N_5558);
or U7565 (N_7565,N_4587,N_5933);
or U7566 (N_7566,N_5211,N_4191);
and U7567 (N_7567,N_5110,N_4416);
xor U7568 (N_7568,N_4595,N_5839);
or U7569 (N_7569,N_4691,N_4948);
and U7570 (N_7570,N_5022,N_5453);
nand U7571 (N_7571,N_4578,N_4484);
nand U7572 (N_7572,N_5293,N_5590);
or U7573 (N_7573,N_4434,N_5298);
nor U7574 (N_7574,N_4066,N_4015);
or U7575 (N_7575,N_5717,N_5460);
or U7576 (N_7576,N_5214,N_4069);
nor U7577 (N_7577,N_4620,N_5095);
nand U7578 (N_7578,N_4462,N_4541);
or U7579 (N_7579,N_5895,N_5315);
nand U7580 (N_7580,N_4284,N_5175);
nand U7581 (N_7581,N_4614,N_4100);
or U7582 (N_7582,N_4592,N_5298);
and U7583 (N_7583,N_4212,N_4747);
nand U7584 (N_7584,N_5903,N_5992);
and U7585 (N_7585,N_4667,N_4710);
or U7586 (N_7586,N_5058,N_5669);
nor U7587 (N_7587,N_5182,N_5611);
and U7588 (N_7588,N_4549,N_5001);
nand U7589 (N_7589,N_5034,N_4686);
nor U7590 (N_7590,N_4533,N_4024);
or U7591 (N_7591,N_5559,N_4877);
nand U7592 (N_7592,N_5849,N_5190);
nand U7593 (N_7593,N_5445,N_5527);
or U7594 (N_7594,N_4659,N_4665);
nand U7595 (N_7595,N_4002,N_4135);
nor U7596 (N_7596,N_5073,N_4912);
or U7597 (N_7597,N_5793,N_5362);
xor U7598 (N_7598,N_5055,N_5875);
nor U7599 (N_7599,N_5655,N_5047);
nor U7600 (N_7600,N_5704,N_4818);
or U7601 (N_7601,N_4355,N_5158);
nor U7602 (N_7602,N_4169,N_4062);
nand U7603 (N_7603,N_5570,N_4651);
or U7604 (N_7604,N_5877,N_5069);
and U7605 (N_7605,N_4290,N_4955);
or U7606 (N_7606,N_5097,N_5730);
and U7607 (N_7607,N_5999,N_5157);
nor U7608 (N_7608,N_5077,N_4077);
nor U7609 (N_7609,N_4335,N_5197);
nor U7610 (N_7610,N_5373,N_4706);
nor U7611 (N_7611,N_4222,N_4964);
nor U7612 (N_7612,N_5062,N_4193);
and U7613 (N_7613,N_5261,N_4238);
nor U7614 (N_7614,N_5845,N_5027);
and U7615 (N_7615,N_4043,N_5820);
or U7616 (N_7616,N_4805,N_5130);
nor U7617 (N_7617,N_4200,N_5072);
and U7618 (N_7618,N_4355,N_5849);
nand U7619 (N_7619,N_4162,N_4963);
nor U7620 (N_7620,N_5056,N_5980);
and U7621 (N_7621,N_4495,N_5418);
or U7622 (N_7622,N_5885,N_4607);
nand U7623 (N_7623,N_4861,N_5502);
and U7624 (N_7624,N_4039,N_4166);
and U7625 (N_7625,N_5273,N_5420);
and U7626 (N_7626,N_5274,N_5598);
nand U7627 (N_7627,N_4269,N_4343);
nor U7628 (N_7628,N_5327,N_4628);
and U7629 (N_7629,N_5196,N_4731);
nor U7630 (N_7630,N_4108,N_5902);
nand U7631 (N_7631,N_5423,N_4443);
nand U7632 (N_7632,N_5464,N_5610);
nand U7633 (N_7633,N_4109,N_5282);
or U7634 (N_7634,N_4219,N_5752);
and U7635 (N_7635,N_4956,N_4678);
or U7636 (N_7636,N_4700,N_5992);
nor U7637 (N_7637,N_4923,N_5278);
nand U7638 (N_7638,N_4842,N_5375);
nand U7639 (N_7639,N_5328,N_5577);
or U7640 (N_7640,N_4441,N_5505);
nand U7641 (N_7641,N_4988,N_5420);
or U7642 (N_7642,N_5084,N_4256);
nor U7643 (N_7643,N_5512,N_5479);
and U7644 (N_7644,N_5550,N_4724);
and U7645 (N_7645,N_5715,N_5475);
nand U7646 (N_7646,N_4172,N_5512);
and U7647 (N_7647,N_4099,N_5894);
or U7648 (N_7648,N_4264,N_4036);
nor U7649 (N_7649,N_5552,N_5064);
and U7650 (N_7650,N_5876,N_5176);
nor U7651 (N_7651,N_4501,N_4885);
nor U7652 (N_7652,N_5720,N_4912);
or U7653 (N_7653,N_4895,N_4460);
and U7654 (N_7654,N_4228,N_4854);
or U7655 (N_7655,N_5506,N_4319);
xnor U7656 (N_7656,N_5668,N_5140);
or U7657 (N_7657,N_5782,N_5448);
nor U7658 (N_7658,N_5156,N_5980);
and U7659 (N_7659,N_4267,N_4314);
nor U7660 (N_7660,N_4893,N_4810);
nand U7661 (N_7661,N_5326,N_4610);
or U7662 (N_7662,N_4621,N_4557);
nand U7663 (N_7663,N_5310,N_4663);
or U7664 (N_7664,N_4145,N_4771);
or U7665 (N_7665,N_5402,N_4389);
nand U7666 (N_7666,N_4043,N_5775);
nand U7667 (N_7667,N_4817,N_5906);
nand U7668 (N_7668,N_4003,N_4191);
nand U7669 (N_7669,N_4105,N_5092);
nand U7670 (N_7670,N_5568,N_4358);
nor U7671 (N_7671,N_4674,N_5491);
nand U7672 (N_7672,N_4933,N_5436);
or U7673 (N_7673,N_5880,N_5464);
or U7674 (N_7674,N_5609,N_4019);
nand U7675 (N_7675,N_4822,N_5905);
nand U7676 (N_7676,N_5592,N_5619);
or U7677 (N_7677,N_4506,N_4179);
and U7678 (N_7678,N_4720,N_5913);
nor U7679 (N_7679,N_5995,N_4001);
nor U7680 (N_7680,N_4680,N_4459);
nor U7681 (N_7681,N_5990,N_4790);
nand U7682 (N_7682,N_4431,N_4805);
nand U7683 (N_7683,N_4178,N_4469);
nor U7684 (N_7684,N_4744,N_5698);
and U7685 (N_7685,N_5971,N_5415);
or U7686 (N_7686,N_5557,N_5154);
nor U7687 (N_7687,N_4613,N_4283);
nor U7688 (N_7688,N_4351,N_5347);
nor U7689 (N_7689,N_5200,N_4136);
nand U7690 (N_7690,N_4621,N_4117);
or U7691 (N_7691,N_5052,N_4448);
and U7692 (N_7692,N_4122,N_4421);
and U7693 (N_7693,N_5046,N_5054);
or U7694 (N_7694,N_5726,N_5316);
nor U7695 (N_7695,N_5509,N_5164);
or U7696 (N_7696,N_5570,N_5021);
or U7697 (N_7697,N_4748,N_5322);
or U7698 (N_7698,N_4031,N_4763);
or U7699 (N_7699,N_4370,N_4676);
and U7700 (N_7700,N_5058,N_5235);
nand U7701 (N_7701,N_5415,N_4255);
nor U7702 (N_7702,N_5465,N_5210);
nor U7703 (N_7703,N_4343,N_4563);
nor U7704 (N_7704,N_4042,N_4733);
nand U7705 (N_7705,N_4927,N_5138);
nor U7706 (N_7706,N_5285,N_4669);
nor U7707 (N_7707,N_5187,N_5188);
and U7708 (N_7708,N_4359,N_5235);
nand U7709 (N_7709,N_4886,N_5809);
and U7710 (N_7710,N_4201,N_4799);
and U7711 (N_7711,N_5052,N_5123);
xnor U7712 (N_7712,N_5281,N_5289);
or U7713 (N_7713,N_5377,N_4787);
nor U7714 (N_7714,N_5724,N_4634);
and U7715 (N_7715,N_4788,N_4068);
nand U7716 (N_7716,N_4626,N_5547);
or U7717 (N_7717,N_5712,N_4811);
nor U7718 (N_7718,N_4693,N_4879);
or U7719 (N_7719,N_5522,N_4591);
and U7720 (N_7720,N_4438,N_4970);
nand U7721 (N_7721,N_5598,N_5911);
and U7722 (N_7722,N_5311,N_4919);
or U7723 (N_7723,N_4885,N_4390);
and U7724 (N_7724,N_4187,N_4470);
or U7725 (N_7725,N_4736,N_5885);
nor U7726 (N_7726,N_5333,N_4820);
xor U7727 (N_7727,N_4475,N_4431);
nand U7728 (N_7728,N_4764,N_4200);
nand U7729 (N_7729,N_4719,N_5918);
and U7730 (N_7730,N_5744,N_5837);
nand U7731 (N_7731,N_4113,N_5217);
and U7732 (N_7732,N_5755,N_5558);
nand U7733 (N_7733,N_5251,N_5109);
and U7734 (N_7734,N_4465,N_4315);
nor U7735 (N_7735,N_5831,N_5111);
and U7736 (N_7736,N_4979,N_4989);
or U7737 (N_7737,N_4554,N_5545);
nand U7738 (N_7738,N_5023,N_5739);
nor U7739 (N_7739,N_5736,N_4941);
and U7740 (N_7740,N_5626,N_5571);
or U7741 (N_7741,N_5378,N_5881);
and U7742 (N_7742,N_5442,N_5181);
or U7743 (N_7743,N_5723,N_4944);
nand U7744 (N_7744,N_5637,N_4154);
nand U7745 (N_7745,N_4334,N_5920);
and U7746 (N_7746,N_5562,N_5970);
nor U7747 (N_7747,N_4855,N_4763);
and U7748 (N_7748,N_5050,N_5811);
or U7749 (N_7749,N_4423,N_5535);
nor U7750 (N_7750,N_5252,N_5195);
and U7751 (N_7751,N_4767,N_4265);
or U7752 (N_7752,N_5760,N_5201);
nor U7753 (N_7753,N_5710,N_4102);
nor U7754 (N_7754,N_5629,N_4660);
or U7755 (N_7755,N_5355,N_4354);
nand U7756 (N_7756,N_5015,N_5413);
or U7757 (N_7757,N_4943,N_5509);
and U7758 (N_7758,N_5539,N_5558);
nor U7759 (N_7759,N_4216,N_5221);
nand U7760 (N_7760,N_5240,N_5265);
and U7761 (N_7761,N_5011,N_5416);
and U7762 (N_7762,N_4906,N_5228);
nand U7763 (N_7763,N_4687,N_5089);
or U7764 (N_7764,N_5899,N_5376);
nor U7765 (N_7765,N_4473,N_5647);
nand U7766 (N_7766,N_4717,N_5971);
nand U7767 (N_7767,N_5662,N_5411);
nor U7768 (N_7768,N_5369,N_4315);
or U7769 (N_7769,N_5508,N_5306);
nor U7770 (N_7770,N_5198,N_5065);
or U7771 (N_7771,N_4491,N_4283);
and U7772 (N_7772,N_4763,N_4175);
nor U7773 (N_7773,N_4962,N_5139);
and U7774 (N_7774,N_4258,N_5527);
and U7775 (N_7775,N_5944,N_4809);
nand U7776 (N_7776,N_4730,N_4408);
nor U7777 (N_7777,N_4294,N_5628);
nor U7778 (N_7778,N_5035,N_4616);
or U7779 (N_7779,N_4439,N_4958);
and U7780 (N_7780,N_4840,N_5170);
nor U7781 (N_7781,N_5408,N_5089);
or U7782 (N_7782,N_5072,N_5720);
nand U7783 (N_7783,N_4377,N_5432);
or U7784 (N_7784,N_4470,N_5479);
and U7785 (N_7785,N_4065,N_5881);
nand U7786 (N_7786,N_4073,N_5486);
xor U7787 (N_7787,N_4457,N_5478);
or U7788 (N_7788,N_4894,N_4178);
or U7789 (N_7789,N_5076,N_5906);
nor U7790 (N_7790,N_4840,N_4842);
nor U7791 (N_7791,N_5930,N_5521);
or U7792 (N_7792,N_4240,N_5534);
nand U7793 (N_7793,N_5832,N_4668);
nand U7794 (N_7794,N_4790,N_4766);
or U7795 (N_7795,N_5584,N_5959);
nor U7796 (N_7796,N_5830,N_5407);
or U7797 (N_7797,N_5185,N_5157);
and U7798 (N_7798,N_4691,N_4051);
and U7799 (N_7799,N_5584,N_4253);
or U7800 (N_7800,N_5911,N_4522);
nand U7801 (N_7801,N_5103,N_4994);
nand U7802 (N_7802,N_4826,N_5077);
nand U7803 (N_7803,N_4477,N_5718);
nor U7804 (N_7804,N_4398,N_4830);
nand U7805 (N_7805,N_4754,N_5723);
nand U7806 (N_7806,N_5508,N_4850);
nand U7807 (N_7807,N_4613,N_5428);
nor U7808 (N_7808,N_4348,N_4920);
or U7809 (N_7809,N_4447,N_5965);
nand U7810 (N_7810,N_5051,N_4024);
nand U7811 (N_7811,N_4685,N_4146);
nor U7812 (N_7812,N_4864,N_4723);
nand U7813 (N_7813,N_4388,N_5735);
nand U7814 (N_7814,N_4541,N_5125);
xor U7815 (N_7815,N_5972,N_5930);
or U7816 (N_7816,N_4156,N_5918);
nand U7817 (N_7817,N_5542,N_4712);
nand U7818 (N_7818,N_5027,N_4615);
or U7819 (N_7819,N_5312,N_4422);
and U7820 (N_7820,N_4980,N_5121);
nor U7821 (N_7821,N_5613,N_4765);
nand U7822 (N_7822,N_5959,N_4945);
nor U7823 (N_7823,N_4213,N_4807);
nand U7824 (N_7824,N_5121,N_5436);
nor U7825 (N_7825,N_4263,N_4564);
nand U7826 (N_7826,N_4712,N_5769);
or U7827 (N_7827,N_5037,N_4031);
or U7828 (N_7828,N_4280,N_5955);
nand U7829 (N_7829,N_5874,N_5635);
nand U7830 (N_7830,N_4063,N_5986);
or U7831 (N_7831,N_4526,N_5544);
or U7832 (N_7832,N_4164,N_5890);
nor U7833 (N_7833,N_4888,N_4850);
nor U7834 (N_7834,N_5828,N_4825);
nand U7835 (N_7835,N_5748,N_4149);
nor U7836 (N_7836,N_5915,N_5546);
or U7837 (N_7837,N_4043,N_5592);
or U7838 (N_7838,N_4285,N_5824);
and U7839 (N_7839,N_4371,N_5538);
nand U7840 (N_7840,N_4627,N_4230);
nor U7841 (N_7841,N_4499,N_5009);
and U7842 (N_7842,N_5058,N_4320);
nand U7843 (N_7843,N_5948,N_4107);
nor U7844 (N_7844,N_4373,N_5140);
and U7845 (N_7845,N_4283,N_5547);
and U7846 (N_7846,N_4864,N_4016);
nand U7847 (N_7847,N_4949,N_5174);
and U7848 (N_7848,N_4921,N_5160);
and U7849 (N_7849,N_4019,N_5058);
nor U7850 (N_7850,N_5332,N_4469);
nor U7851 (N_7851,N_4793,N_5813);
nor U7852 (N_7852,N_4573,N_5555);
or U7853 (N_7853,N_5686,N_4773);
and U7854 (N_7854,N_5863,N_4682);
or U7855 (N_7855,N_5120,N_4437);
or U7856 (N_7856,N_5695,N_5182);
or U7857 (N_7857,N_4663,N_5975);
nand U7858 (N_7858,N_4688,N_4047);
or U7859 (N_7859,N_4344,N_5741);
or U7860 (N_7860,N_4363,N_5576);
and U7861 (N_7861,N_5840,N_5789);
and U7862 (N_7862,N_4562,N_4163);
or U7863 (N_7863,N_5874,N_4078);
nand U7864 (N_7864,N_4089,N_5719);
and U7865 (N_7865,N_4820,N_4929);
and U7866 (N_7866,N_5457,N_4378);
xnor U7867 (N_7867,N_4167,N_5020);
nor U7868 (N_7868,N_5233,N_4322);
nand U7869 (N_7869,N_5107,N_5953);
and U7870 (N_7870,N_4369,N_5890);
nor U7871 (N_7871,N_5070,N_5356);
and U7872 (N_7872,N_4025,N_4122);
nor U7873 (N_7873,N_4391,N_4314);
or U7874 (N_7874,N_4494,N_5662);
and U7875 (N_7875,N_4848,N_4576);
nand U7876 (N_7876,N_4421,N_4705);
or U7877 (N_7877,N_4972,N_4040);
nor U7878 (N_7878,N_5775,N_5408);
nand U7879 (N_7879,N_5326,N_5147);
or U7880 (N_7880,N_4184,N_4968);
nand U7881 (N_7881,N_5762,N_4909);
nor U7882 (N_7882,N_5148,N_4543);
nand U7883 (N_7883,N_4740,N_5024);
or U7884 (N_7884,N_5327,N_5644);
and U7885 (N_7885,N_5830,N_4417);
or U7886 (N_7886,N_5602,N_5324);
and U7887 (N_7887,N_5095,N_5177);
and U7888 (N_7888,N_5865,N_4018);
or U7889 (N_7889,N_4762,N_5814);
and U7890 (N_7890,N_4916,N_5134);
or U7891 (N_7891,N_5936,N_4003);
nor U7892 (N_7892,N_5614,N_4353);
or U7893 (N_7893,N_5251,N_4451);
nor U7894 (N_7894,N_5289,N_5564);
nor U7895 (N_7895,N_4352,N_5031);
nor U7896 (N_7896,N_4531,N_5585);
nand U7897 (N_7897,N_4025,N_4015);
nand U7898 (N_7898,N_4045,N_5485);
nor U7899 (N_7899,N_5244,N_4169);
nor U7900 (N_7900,N_4122,N_5242);
and U7901 (N_7901,N_5780,N_5659);
nor U7902 (N_7902,N_4383,N_5395);
and U7903 (N_7903,N_5030,N_5256);
or U7904 (N_7904,N_4249,N_5793);
or U7905 (N_7905,N_5940,N_4834);
nor U7906 (N_7906,N_4627,N_4438);
or U7907 (N_7907,N_5918,N_4136);
nand U7908 (N_7908,N_5654,N_4115);
nor U7909 (N_7909,N_5703,N_4633);
nand U7910 (N_7910,N_5582,N_4749);
nor U7911 (N_7911,N_5534,N_5989);
or U7912 (N_7912,N_4508,N_4542);
or U7913 (N_7913,N_4666,N_4572);
or U7914 (N_7914,N_5309,N_4435);
nand U7915 (N_7915,N_5835,N_4563);
nor U7916 (N_7916,N_4146,N_5811);
or U7917 (N_7917,N_4116,N_4683);
nor U7918 (N_7918,N_4451,N_5367);
and U7919 (N_7919,N_4957,N_4010);
nor U7920 (N_7920,N_4312,N_4186);
nor U7921 (N_7921,N_5140,N_5885);
or U7922 (N_7922,N_5461,N_5665);
and U7923 (N_7923,N_5884,N_4017);
nor U7924 (N_7924,N_5491,N_5753);
or U7925 (N_7925,N_4503,N_5205);
xor U7926 (N_7926,N_5202,N_4658);
xor U7927 (N_7927,N_5669,N_4522);
nand U7928 (N_7928,N_5677,N_4048);
nand U7929 (N_7929,N_5395,N_4911);
nor U7930 (N_7930,N_5589,N_5857);
nand U7931 (N_7931,N_5686,N_5303);
nand U7932 (N_7932,N_5072,N_4131);
and U7933 (N_7933,N_4265,N_5258);
and U7934 (N_7934,N_4983,N_4591);
nand U7935 (N_7935,N_4797,N_5848);
nor U7936 (N_7936,N_4079,N_4223);
or U7937 (N_7937,N_4271,N_5310);
and U7938 (N_7938,N_4414,N_4034);
nor U7939 (N_7939,N_5271,N_5353);
nor U7940 (N_7940,N_4780,N_4611);
nor U7941 (N_7941,N_5989,N_5229);
nand U7942 (N_7942,N_4790,N_4092);
or U7943 (N_7943,N_5921,N_5285);
nand U7944 (N_7944,N_5402,N_5923);
and U7945 (N_7945,N_4910,N_5008);
or U7946 (N_7946,N_5460,N_5242);
nor U7947 (N_7947,N_4360,N_5968);
nand U7948 (N_7948,N_5944,N_4794);
nor U7949 (N_7949,N_5585,N_4053);
nor U7950 (N_7950,N_5841,N_4914);
or U7951 (N_7951,N_5451,N_4510);
and U7952 (N_7952,N_5893,N_4982);
nor U7953 (N_7953,N_5391,N_5680);
nand U7954 (N_7954,N_5335,N_5216);
nor U7955 (N_7955,N_5639,N_5850);
and U7956 (N_7956,N_5889,N_4371);
or U7957 (N_7957,N_5343,N_4023);
and U7958 (N_7958,N_5075,N_4718);
and U7959 (N_7959,N_5035,N_5926);
and U7960 (N_7960,N_4384,N_5127);
nor U7961 (N_7961,N_4844,N_4861);
nor U7962 (N_7962,N_5652,N_5649);
or U7963 (N_7963,N_4879,N_5600);
and U7964 (N_7964,N_4117,N_5759);
nand U7965 (N_7965,N_4381,N_5030);
nand U7966 (N_7966,N_4701,N_5076);
nor U7967 (N_7967,N_4200,N_5984);
and U7968 (N_7968,N_4055,N_4314);
and U7969 (N_7969,N_5038,N_4072);
nand U7970 (N_7970,N_5829,N_4059);
or U7971 (N_7971,N_5613,N_4397);
or U7972 (N_7972,N_5814,N_4652);
and U7973 (N_7973,N_5329,N_5358);
or U7974 (N_7974,N_5219,N_5609);
or U7975 (N_7975,N_4922,N_4351);
and U7976 (N_7976,N_5616,N_5512);
and U7977 (N_7977,N_4140,N_5169);
and U7978 (N_7978,N_5065,N_5360);
nand U7979 (N_7979,N_4818,N_4010);
nor U7980 (N_7980,N_4221,N_5527);
nor U7981 (N_7981,N_4225,N_5551);
nor U7982 (N_7982,N_4030,N_4735);
nand U7983 (N_7983,N_4370,N_4087);
xor U7984 (N_7984,N_5348,N_5703);
or U7985 (N_7985,N_5821,N_5324);
nor U7986 (N_7986,N_4137,N_5648);
nand U7987 (N_7987,N_4117,N_5575);
nor U7988 (N_7988,N_4714,N_4366);
nand U7989 (N_7989,N_4743,N_4874);
nor U7990 (N_7990,N_5529,N_5381);
or U7991 (N_7991,N_4605,N_5873);
nand U7992 (N_7992,N_5859,N_4442);
nand U7993 (N_7993,N_5122,N_5661);
nand U7994 (N_7994,N_5794,N_5495);
nor U7995 (N_7995,N_5126,N_4528);
and U7996 (N_7996,N_4455,N_5958);
nor U7997 (N_7997,N_5389,N_4450);
and U7998 (N_7998,N_5644,N_4665);
nor U7999 (N_7999,N_5118,N_5653);
nor U8000 (N_8000,N_7099,N_7986);
nand U8001 (N_8001,N_6779,N_7589);
or U8002 (N_8002,N_6841,N_7610);
nand U8003 (N_8003,N_6972,N_6023);
nor U8004 (N_8004,N_7495,N_6766);
or U8005 (N_8005,N_7643,N_6606);
or U8006 (N_8006,N_7288,N_6134);
nand U8007 (N_8007,N_7568,N_7575);
nand U8008 (N_8008,N_7714,N_7534);
or U8009 (N_8009,N_7595,N_7564);
or U8010 (N_8010,N_7444,N_6494);
nand U8011 (N_8011,N_7787,N_7142);
nand U8012 (N_8012,N_7699,N_7219);
nand U8013 (N_8013,N_7826,N_7007);
and U8014 (N_8014,N_6338,N_6179);
or U8015 (N_8015,N_6824,N_7549);
nand U8016 (N_8016,N_6409,N_6844);
nand U8017 (N_8017,N_6503,N_7899);
or U8018 (N_8018,N_6658,N_7279);
nor U8019 (N_8019,N_6519,N_7351);
and U8020 (N_8020,N_6545,N_6860);
nor U8021 (N_8021,N_7242,N_6383);
nand U8022 (N_8022,N_7200,N_7260);
and U8023 (N_8023,N_7003,N_6728);
and U8024 (N_8024,N_6852,N_6075);
nand U8025 (N_8025,N_6129,N_6774);
and U8026 (N_8026,N_7909,N_7335);
nand U8027 (N_8027,N_7488,N_7792);
xor U8028 (N_8028,N_6107,N_6120);
nor U8029 (N_8029,N_6450,N_6556);
and U8030 (N_8030,N_7319,N_6663);
nor U8031 (N_8031,N_6033,N_7516);
or U8032 (N_8032,N_7720,N_7538);
or U8033 (N_8033,N_6891,N_6276);
nand U8034 (N_8034,N_6289,N_6470);
and U8035 (N_8035,N_6196,N_7917);
nand U8036 (N_8036,N_7911,N_7834);
nand U8037 (N_8037,N_6133,N_7703);
nor U8038 (N_8038,N_6329,N_6536);
and U8039 (N_8039,N_7565,N_7827);
nor U8040 (N_8040,N_7330,N_7512);
and U8041 (N_8041,N_6359,N_6219);
nor U8042 (N_8042,N_7076,N_6523);
and U8043 (N_8043,N_7008,N_7881);
nor U8044 (N_8044,N_7181,N_6006);
or U8045 (N_8045,N_6933,N_7172);
nand U8046 (N_8046,N_7506,N_6853);
and U8047 (N_8047,N_7618,N_6427);
and U8048 (N_8048,N_7135,N_7047);
nand U8049 (N_8049,N_7615,N_7851);
and U8050 (N_8050,N_6305,N_6081);
nor U8051 (N_8051,N_6594,N_6445);
nand U8052 (N_8052,N_7119,N_6463);
nor U8053 (N_8053,N_6464,N_7405);
nand U8054 (N_8054,N_7663,N_7887);
or U8055 (N_8055,N_6121,N_7111);
nor U8056 (N_8056,N_7636,N_7277);
and U8057 (N_8057,N_7089,N_6428);
nor U8058 (N_8058,N_7088,N_7372);
or U8059 (N_8059,N_6690,N_7596);
nor U8060 (N_8060,N_6735,N_6817);
and U8061 (N_8061,N_7964,N_6015);
and U8062 (N_8062,N_6508,N_7841);
nand U8063 (N_8063,N_6652,N_7650);
nor U8064 (N_8064,N_7418,N_7745);
nor U8065 (N_8065,N_6813,N_7144);
or U8066 (N_8066,N_6991,N_6723);
nand U8067 (N_8067,N_6716,N_6603);
or U8068 (N_8068,N_7670,N_7872);
or U8069 (N_8069,N_7107,N_6249);
nor U8070 (N_8070,N_7868,N_7258);
nand U8071 (N_8071,N_6098,N_7863);
nand U8072 (N_8072,N_6632,N_6402);
nor U8073 (N_8073,N_6783,N_6765);
nand U8074 (N_8074,N_6665,N_6253);
nand U8075 (N_8075,N_6158,N_7073);
nor U8076 (N_8076,N_6586,N_6234);
or U8077 (N_8077,N_6221,N_7097);
or U8078 (N_8078,N_7379,N_6283);
or U8079 (N_8079,N_7748,N_6975);
nor U8080 (N_8080,N_7044,N_6004);
or U8081 (N_8081,N_6713,N_6589);
or U8082 (N_8082,N_7944,N_7769);
or U8083 (N_8083,N_6225,N_6397);
nand U8084 (N_8084,N_6073,N_6250);
and U8085 (N_8085,N_7083,N_7197);
and U8086 (N_8086,N_7919,N_7475);
and U8087 (N_8087,N_6188,N_7025);
nand U8088 (N_8088,N_6672,N_6164);
or U8089 (N_8089,N_6647,N_7451);
or U8090 (N_8090,N_6016,N_7598);
nor U8091 (N_8091,N_7293,N_6432);
nor U8092 (N_8092,N_7424,N_7173);
or U8093 (N_8093,N_7949,N_6264);
or U8094 (N_8094,N_7784,N_6104);
or U8095 (N_8095,N_6823,N_7676);
and U8096 (N_8096,N_6487,N_7693);
or U8097 (N_8097,N_7168,N_6115);
or U8098 (N_8098,N_6204,N_7491);
nand U8099 (N_8099,N_6590,N_7873);
or U8100 (N_8100,N_6857,N_7979);
and U8101 (N_8101,N_6983,N_6879);
or U8102 (N_8102,N_6855,N_6867);
nor U8103 (N_8103,N_7735,N_6695);
nand U8104 (N_8104,N_7672,N_7952);
nor U8105 (N_8105,N_7519,N_6802);
and U8106 (N_8106,N_6419,N_7668);
nand U8107 (N_8107,N_7347,N_7913);
nor U8108 (N_8108,N_7785,N_7509);
nand U8109 (N_8109,N_6822,N_7696);
or U8110 (N_8110,N_7145,N_7018);
or U8111 (N_8111,N_6872,N_7716);
or U8112 (N_8112,N_6831,N_7381);
or U8113 (N_8113,N_7114,N_7504);
nand U8114 (N_8114,N_6273,N_7551);
and U8115 (N_8115,N_7946,N_6166);
nand U8116 (N_8116,N_6980,N_6581);
or U8117 (N_8117,N_7485,N_7717);
nor U8118 (N_8118,N_7477,N_6465);
or U8119 (N_8119,N_6788,N_7532);
and U8120 (N_8120,N_6638,N_7830);
nor U8121 (N_8121,N_7373,N_6531);
or U8122 (N_8122,N_6616,N_7237);
nand U8123 (N_8123,N_7022,N_7907);
and U8124 (N_8124,N_6185,N_7581);
and U8125 (N_8125,N_6694,N_6296);
or U8126 (N_8126,N_7726,N_7484);
and U8127 (N_8127,N_6248,N_7098);
or U8128 (N_8128,N_7426,N_7198);
or U8129 (N_8129,N_7705,N_7371);
or U8130 (N_8130,N_6335,N_7240);
and U8131 (N_8131,N_6314,N_7791);
nor U8132 (N_8132,N_7162,N_7065);
and U8133 (N_8133,N_6350,N_6444);
xor U8134 (N_8134,N_7657,N_7442);
nor U8135 (N_8135,N_7280,N_6082);
and U8136 (N_8136,N_6052,N_7563);
or U8137 (N_8137,N_6377,N_6769);
and U8138 (N_8138,N_6024,N_6733);
nand U8139 (N_8139,N_6436,N_7202);
or U8140 (N_8140,N_7447,N_7973);
nand U8141 (N_8141,N_7051,N_7250);
nor U8142 (N_8142,N_6984,N_6136);
nor U8143 (N_8143,N_6398,N_6643);
nand U8144 (N_8144,N_6348,N_6132);
nand U8145 (N_8145,N_7223,N_6499);
nor U8146 (N_8146,N_6753,N_6969);
nand U8147 (N_8147,N_7191,N_6563);
and U8148 (N_8148,N_7457,N_6598);
nor U8149 (N_8149,N_6080,N_7631);
nand U8150 (N_8150,N_7077,N_7421);
xnor U8151 (N_8151,N_7734,N_7861);
or U8152 (N_8152,N_7230,N_6256);
or U8153 (N_8153,N_7729,N_7039);
xor U8154 (N_8154,N_6722,N_7313);
and U8155 (N_8155,N_7943,N_6315);
nor U8156 (N_8156,N_7486,N_7758);
or U8157 (N_8157,N_7196,N_6391);
or U8158 (N_8158,N_6119,N_6462);
or U8159 (N_8159,N_6372,N_7993);
and U8160 (N_8160,N_6801,N_6193);
nand U8161 (N_8161,N_6306,N_6534);
nor U8162 (N_8162,N_6698,N_7015);
and U8163 (N_8163,N_7637,N_7527);
nor U8164 (N_8164,N_6094,N_7072);
and U8165 (N_8165,N_6384,N_6259);
nand U8166 (N_8166,N_7679,N_7209);
and U8167 (N_8167,N_7883,N_7174);
or U8168 (N_8168,N_7744,N_6020);
nor U8169 (N_8169,N_6954,N_6945);
nor U8170 (N_8170,N_6684,N_6689);
or U8171 (N_8171,N_7606,N_6803);
or U8172 (N_8172,N_7924,N_7317);
and U8173 (N_8173,N_6692,N_6005);
nand U8174 (N_8174,N_6940,N_7776);
nor U8175 (N_8175,N_6997,N_7754);
or U8176 (N_8176,N_6175,N_7374);
nor U8177 (N_8177,N_6067,N_6168);
or U8178 (N_8178,N_7803,N_6555);
or U8179 (N_8179,N_7594,N_7328);
nor U8180 (N_8180,N_7865,N_6217);
nand U8181 (N_8181,N_6008,N_7284);
nand U8182 (N_8182,N_7244,N_7882);
or U8183 (N_8183,N_6622,N_7265);
and U8184 (N_8184,N_7904,N_7462);
nand U8185 (N_8185,N_6302,N_6209);
or U8186 (N_8186,N_7613,N_6591);
nand U8187 (N_8187,N_6439,N_7027);
nand U8188 (N_8188,N_6559,N_7722);
or U8189 (N_8189,N_7701,N_6725);
and U8190 (N_8190,N_6513,N_6554);
nand U8191 (N_8191,N_7742,N_7248);
and U8192 (N_8192,N_7439,N_7297);
nor U8193 (N_8193,N_6916,N_7468);
nor U8194 (N_8194,N_7091,N_6349);
nor U8195 (N_8195,N_7109,N_7523);
and U8196 (N_8196,N_6245,N_6345);
and U8197 (N_8197,N_7796,N_6207);
xnor U8198 (N_8198,N_6744,N_7988);
and U8199 (N_8199,N_7286,N_6657);
nand U8200 (N_8200,N_6490,N_7361);
and U8201 (N_8201,N_6892,N_7362);
nor U8202 (N_8202,N_6573,N_6058);
nand U8203 (N_8203,N_6608,N_7306);
nand U8204 (N_8204,N_7352,N_6671);
nor U8205 (N_8205,N_6437,N_7525);
or U8206 (N_8206,N_7315,N_7471);
and U8207 (N_8207,N_7947,N_6660);
or U8208 (N_8208,N_7389,N_6840);
nor U8209 (N_8209,N_7228,N_7053);
nand U8210 (N_8210,N_6039,N_6491);
nor U8211 (N_8211,N_7945,N_6192);
and U8212 (N_8212,N_7210,N_7357);
nand U8213 (N_8213,N_7460,N_6010);
and U8214 (N_8214,N_6732,N_7817);
and U8215 (N_8215,N_6048,N_6325);
nand U8216 (N_8216,N_7948,N_7725);
or U8217 (N_8217,N_6995,N_7422);
nor U8218 (N_8218,N_7682,N_7493);
nor U8219 (N_8219,N_6927,N_7329);
or U8220 (N_8220,N_7354,N_7113);
and U8221 (N_8221,N_7648,N_6829);
or U8222 (N_8222,N_6908,N_7490);
nor U8223 (N_8223,N_7247,N_6926);
nor U8224 (N_8224,N_6510,N_7296);
xnor U8225 (N_8225,N_7399,N_6739);
nor U8226 (N_8226,N_6550,N_6291);
nand U8227 (N_8227,N_7012,N_7910);
and U8228 (N_8228,N_6165,N_6928);
nand U8229 (N_8229,N_6992,N_6096);
or U8230 (N_8230,N_6496,N_7128);
and U8231 (N_8231,N_6308,N_6903);
nor U8232 (N_8232,N_6833,N_6157);
and U8233 (N_8233,N_7252,N_7343);
nand U8234 (N_8234,N_6546,N_6205);
nand U8235 (N_8235,N_7987,N_6621);
nand U8236 (N_8236,N_6213,N_7544);
nor U8237 (N_8237,N_7915,N_7875);
nor U8238 (N_8238,N_7804,N_7190);
or U8239 (N_8239,N_6862,N_6569);
and U8240 (N_8240,N_7178,N_7625);
nand U8241 (N_8241,N_7478,N_7344);
nor U8242 (N_8242,N_7878,N_6812);
nand U8243 (N_8243,N_6049,N_6644);
nand U8244 (N_8244,N_7667,N_7423);
nand U8245 (N_8245,N_6442,N_6731);
or U8246 (N_8246,N_6413,N_7753);
nand U8247 (N_8247,N_6270,N_6599);
or U8248 (N_8248,N_6288,N_6474);
and U8249 (N_8249,N_7176,N_7188);
nor U8250 (N_8250,N_6105,N_6497);
nand U8251 (N_8251,N_7542,N_6810);
nor U8252 (N_8252,N_6395,N_7342);
nand U8253 (N_8253,N_7459,N_6422);
xnor U8254 (N_8254,N_7844,N_6155);
and U8255 (N_8255,N_7350,N_7182);
and U8256 (N_8256,N_6635,N_6246);
nor U8257 (N_8257,N_6012,N_7566);
nor U8258 (N_8258,N_7673,N_6939);
or U8259 (N_8259,N_6751,N_6214);
or U8260 (N_8260,N_6904,N_6141);
nor U8261 (N_8261,N_6382,N_7002);
or U8262 (N_8262,N_6304,N_6455);
nand U8263 (N_8263,N_7123,N_7583);
and U8264 (N_8264,N_7125,N_6650);
nor U8265 (N_8265,N_6285,N_6784);
nor U8266 (N_8266,N_7068,N_7724);
and U8267 (N_8267,N_6896,N_7074);
or U8268 (N_8268,N_6022,N_7063);
and U8269 (N_8269,N_7169,N_7760);
or U8270 (N_8270,N_7750,N_7243);
xnor U8271 (N_8271,N_6717,N_7283);
nor U8272 (N_8272,N_6292,N_7794);
nand U8273 (N_8273,N_7740,N_6267);
nor U8274 (N_8274,N_7756,N_6623);
and U8275 (N_8275,N_6887,N_7552);
or U8276 (N_8276,N_6173,N_6092);
and U8277 (N_8277,N_7553,N_7028);
and U8278 (N_8278,N_7404,N_7939);
and U8279 (N_8279,N_6243,N_7446);
nand U8280 (N_8280,N_6522,N_6056);
nand U8281 (N_8281,N_6232,N_7384);
or U8282 (N_8282,N_6152,N_6000);
or U8283 (N_8283,N_7236,N_7871);
nor U8284 (N_8284,N_7120,N_7082);
nor U8285 (N_8285,N_6262,N_6930);
or U8286 (N_8286,N_6147,N_7500);
nand U8287 (N_8287,N_7896,N_7307);
nand U8288 (N_8288,N_7560,N_7320);
and U8289 (N_8289,N_6483,N_7658);
nand U8290 (N_8290,N_7383,N_7189);
nand U8291 (N_8291,N_7062,N_7472);
or U8292 (N_8292,N_7194,N_6019);
nor U8293 (N_8293,N_7678,N_6620);
nor U8294 (N_8294,N_6361,N_7266);
and U8295 (N_8295,N_7840,N_7152);
nor U8296 (N_8296,N_7518,N_6985);
or U8297 (N_8297,N_6832,N_7254);
nor U8298 (N_8298,N_7390,N_7709);
nand U8299 (N_8299,N_7430,N_7517);
nand U8300 (N_8300,N_7936,N_6336);
or U8301 (N_8301,N_6626,N_7836);
nand U8302 (N_8302,N_7095,N_6913);
nor U8303 (N_8303,N_7121,N_7134);
nand U8304 (N_8304,N_6431,N_7337);
nor U8305 (N_8305,N_6678,N_7604);
nor U8306 (N_8306,N_7118,N_7775);
or U8307 (N_8307,N_6169,N_6202);
or U8308 (N_8308,N_7163,N_7316);
or U8309 (N_8309,N_6777,N_7149);
or U8310 (N_8310,N_7626,N_6894);
nand U8311 (N_8311,N_7129,N_7960);
nand U8312 (N_8312,N_7810,N_6322);
nand U8313 (N_8313,N_7327,N_6212);
and U8314 (N_8314,N_7481,N_7522);
and U8315 (N_8315,N_6047,N_7751);
nand U8316 (N_8316,N_6401,N_7353);
nor U8317 (N_8317,N_7434,N_6025);
nand U8318 (N_8318,N_7938,N_6977);
or U8319 (N_8319,N_7016,N_7749);
nor U8320 (N_8320,N_6543,N_6344);
and U8321 (N_8321,N_7999,N_6691);
xnor U8322 (N_8322,N_7591,N_7617);
nand U8323 (N_8323,N_7427,N_7757);
nand U8324 (N_8324,N_6925,N_6181);
nor U8325 (N_8325,N_6138,N_7257);
and U8326 (N_8326,N_7852,N_6309);
nand U8327 (N_8327,N_6634,N_6414);
nand U8328 (N_8328,N_6352,N_7982);
and U8329 (N_8329,N_6031,N_7180);
xnor U8330 (N_8330,N_7386,N_7815);
xor U8331 (N_8331,N_6963,N_6438);
nor U8332 (N_8332,N_7203,N_7133);
or U8333 (N_8333,N_6337,N_6710);
nand U8334 (N_8334,N_7922,N_7620);
or U8335 (N_8335,N_6389,N_6077);
nand U8336 (N_8336,N_6949,N_6957);
nor U8337 (N_8337,N_7880,N_7160);
or U8338 (N_8338,N_6441,N_6495);
and U8339 (N_8339,N_7239,N_6533);
nor U8340 (N_8340,N_7023,N_6737);
or U8341 (N_8341,N_6596,N_7037);
nor U8342 (N_8342,N_7743,N_7147);
nand U8343 (N_8343,N_7238,N_7417);
nand U8344 (N_8344,N_6918,N_7245);
and U8345 (N_8345,N_7452,N_6567);
and U8346 (N_8346,N_7848,N_6756);
nand U8347 (N_8347,N_6339,N_6680);
nor U8348 (N_8348,N_6210,N_7453);
nor U8349 (N_8349,N_6360,N_7829);
and U8350 (N_8350,N_7295,N_6501);
nand U8351 (N_8351,N_7420,N_6548);
nand U8352 (N_8352,N_6354,N_6869);
nor U8353 (N_8353,N_6353,N_6961);
or U8354 (N_8354,N_6342,N_7438);
nand U8355 (N_8355,N_6069,N_6907);
or U8356 (N_8356,N_7440,N_7043);
or U8357 (N_8357,N_6745,N_7660);
nor U8358 (N_8358,N_7687,N_6617);
nor U8359 (N_8359,N_6775,N_7856);
nand U8360 (N_8360,N_7222,N_7186);
nor U8361 (N_8361,N_7941,N_6525);
nor U8362 (N_8362,N_7229,N_6816);
xor U8363 (N_8363,N_7862,N_7094);
nor U8364 (N_8364,N_7850,N_6582);
nor U8365 (N_8365,N_6358,N_6102);
nand U8366 (N_8366,N_6043,N_6489);
or U8367 (N_8367,N_6661,N_6641);
nor U8368 (N_8368,N_7360,N_7268);
nand U8369 (N_8369,N_6114,N_6889);
nand U8370 (N_8370,N_7983,N_6109);
and U8371 (N_8371,N_7302,N_7020);
nand U8372 (N_8372,N_7912,N_6989);
and U8373 (N_8373,N_6203,N_7702);
nor U8374 (N_8374,N_7539,N_6378);
nor U8375 (N_8375,N_7771,N_6294);
nand U8376 (N_8376,N_7326,N_6757);
nor U8377 (N_8377,N_7482,N_7824);
and U8378 (N_8378,N_7814,N_6687);
nor U8379 (N_8379,N_6729,N_7788);
or U8380 (N_8380,N_7641,N_6041);
nor U8381 (N_8381,N_7718,N_7846);
nand U8382 (N_8382,N_7489,N_6333);
nor U8383 (N_8383,N_7392,N_7436);
nor U8384 (N_8384,N_7723,N_7175);
xnor U8385 (N_8385,N_7557,N_7078);
nor U8386 (N_8386,N_6231,N_7126);
or U8387 (N_8387,N_6628,N_6484);
nand U8388 (N_8388,N_6953,N_6746);
and U8389 (N_8389,N_7503,N_6355);
and U8390 (N_8390,N_6125,N_7689);
or U8391 (N_8391,N_6649,N_7762);
or U8392 (N_8392,N_6478,N_7727);
nand U8393 (N_8393,N_7502,N_7414);
or U8394 (N_8394,N_7640,N_7093);
or U8395 (N_8395,N_7808,N_6541);
xnor U8396 (N_8396,N_7707,N_7463);
and U8397 (N_8397,N_7321,N_6864);
or U8398 (N_8398,N_6321,N_6705);
nand U8399 (N_8399,N_7927,N_7487);
and U8400 (N_8400,N_7981,N_7621);
and U8401 (N_8401,N_7483,N_6226);
and U8402 (N_8402,N_6973,N_7665);
and U8403 (N_8403,N_6659,N_6874);
nor U8404 (N_8404,N_7780,N_7550);
xor U8405 (N_8405,N_7536,N_6269);
nand U8406 (N_8406,N_7050,N_7666);
nand U8407 (N_8407,N_7032,N_6197);
nand U8408 (N_8408,N_6280,N_7890);
and U8409 (N_8409,N_6265,N_7408);
nand U8410 (N_8410,N_6702,N_7324);
nand U8411 (N_8411,N_7556,N_6310);
or U8412 (N_8412,N_7821,N_6200);
nor U8413 (N_8413,N_7376,N_7639);
nor U8414 (N_8414,N_7739,N_6089);
nand U8415 (N_8415,N_6845,N_7545);
and U8416 (N_8416,N_7064,N_7234);
nand U8417 (N_8417,N_6178,N_6798);
nor U8418 (N_8418,N_7737,N_7406);
nor U8419 (N_8419,N_7644,N_7933);
nor U8420 (N_8420,N_7341,N_7600);
nand U8421 (N_8421,N_7274,N_7976);
or U8422 (N_8422,N_7363,N_6776);
or U8423 (N_8423,N_7645,N_7586);
nand U8424 (N_8424,N_6194,N_6014);
and U8425 (N_8425,N_6394,N_7956);
and U8426 (N_8426,N_7908,N_7412);
or U8427 (N_8427,N_6381,N_6611);
or U8428 (N_8428,N_6859,N_6911);
and U8429 (N_8429,N_6091,N_6459);
and U8430 (N_8430,N_6920,N_7634);
nor U8431 (N_8431,N_7470,N_7261);
nor U8432 (N_8432,N_6003,N_7071);
nand U8433 (N_8433,N_6106,N_6176);
and U8434 (N_8434,N_6607,N_7597);
nor U8435 (N_8435,N_6946,N_6718);
nor U8436 (N_8436,N_6180,N_7199);
nor U8437 (N_8437,N_7692,N_6547);
nand U8438 (N_8438,N_7377,N_6070);
nand U8439 (N_8439,N_6367,N_7662);
nand U8440 (N_8440,N_7096,N_6905);
nor U8441 (N_8441,N_7774,N_7958);
or U8442 (N_8442,N_6063,N_7358);
nor U8443 (N_8443,N_7388,N_6863);
or U8444 (N_8444,N_6252,N_6584);
and U8445 (N_8445,N_7278,N_6341);
nor U8446 (N_8446,N_7588,N_7339);
or U8447 (N_8447,N_6848,N_7079);
nor U8448 (N_8448,N_6524,N_6942);
nor U8449 (N_8449,N_6704,N_7603);
or U8450 (N_8450,N_6362,N_7393);
nand U8451 (N_8451,N_7797,N_7346);
nand U8452 (N_8452,N_7066,N_7712);
and U8453 (N_8453,N_7048,N_6492);
nand U8454 (N_8454,N_7496,N_6981);
nor U8455 (N_8455,N_7131,N_6509);
and U8456 (N_8456,N_7996,N_6222);
nor U8457 (N_8457,N_6423,N_6473);
and U8458 (N_8458,N_7259,N_6668);
and U8459 (N_8459,N_6208,N_6399);
nand U8460 (N_8460,N_6506,N_7289);
nor U8461 (N_8461,N_7100,N_7860);
nand U8462 (N_8462,N_6935,N_6258);
or U8463 (N_8463,N_7322,N_6759);
or U8464 (N_8464,N_6572,N_7501);
and U8465 (N_8465,N_6922,N_6493);
and U8466 (N_8466,N_7396,N_6415);
or U8467 (N_8467,N_6642,N_7014);
nand U8468 (N_8468,N_7975,N_6861);
and U8469 (N_8469,N_7494,N_6849);
and U8470 (N_8470,N_6417,N_7654);
nor U8471 (N_8471,N_7208,N_7579);
or U8472 (N_8472,N_6959,N_6171);
or U8473 (N_8473,N_7281,N_6293);
and U8474 (N_8474,N_6266,N_7906);
and U8475 (N_8475,N_6066,N_6677);
and U8476 (N_8476,N_7736,N_7164);
and U8477 (N_8477,N_7920,N_6486);
nor U8478 (N_8478,N_6738,N_6365);
xnor U8479 (N_8479,N_6055,N_6363);
or U8480 (N_8480,N_6696,N_7700);
or U8481 (N_8481,N_7193,N_7409);
nand U8482 (N_8482,N_7299,N_7599);
or U8483 (N_8483,N_7303,N_7783);
and U8484 (N_8484,N_6577,N_6426);
or U8485 (N_8485,N_6805,N_7675);
nand U8486 (N_8486,N_7526,N_6327);
and U8487 (N_8487,N_7171,N_6471);
or U8488 (N_8488,N_6469,N_7942);
and U8489 (N_8489,N_6866,N_6078);
nor U8490 (N_8490,N_7767,N_7998);
nor U8491 (N_8491,N_7391,N_6159);
nor U8492 (N_8492,N_6122,N_6885);
nand U8493 (N_8493,N_6346,N_7955);
or U8494 (N_8494,N_7355,N_6615);
nor U8495 (N_8495,N_7117,N_7772);
nor U8496 (N_8496,N_7019,N_6386);
xnor U8497 (N_8497,N_6609,N_6449);
or U8498 (N_8498,N_6742,N_7086);
nor U8499 (N_8499,N_6170,N_6387);
nor U8500 (N_8500,N_6369,N_6917);
or U8501 (N_8501,N_7578,N_7158);
xnor U8502 (N_8502,N_7157,N_6135);
nor U8503 (N_8503,N_6518,N_7761);
xor U8504 (N_8504,N_6271,N_6808);
or U8505 (N_8505,N_6924,N_7820);
and U8506 (N_8506,N_6433,N_7445);
nand U8507 (N_8507,N_6646,N_6950);
nand U8508 (N_8508,N_6182,N_7795);
and U8509 (N_8509,N_7653,N_7800);
and U8510 (N_8510,N_6839,N_6686);
nand U8511 (N_8511,N_6190,N_6084);
and U8512 (N_8512,N_6126,N_7994);
and U8513 (N_8513,N_6298,N_7825);
and U8514 (N_8514,N_6446,N_7253);
nor U8515 (N_8515,N_6500,N_6807);
or U8516 (N_8516,N_6111,N_6842);
and U8517 (N_8517,N_7479,N_7609);
nand U8518 (N_8518,N_6943,N_7055);
or U8519 (N_8519,N_7923,N_7590);
or U8520 (N_8520,N_6743,N_6477);
nor U8521 (N_8521,N_7161,N_7980);
nand U8522 (N_8522,N_6050,N_7205);
or U8523 (N_8523,N_6893,N_7467);
and U8524 (N_8524,N_6576,N_7546);
nor U8525 (N_8525,N_6110,N_7985);
and U8526 (N_8526,N_7897,N_6544);
nand U8527 (N_8527,N_6053,N_7204);
nor U8528 (N_8528,N_6850,N_6639);
nor U8529 (N_8529,N_7690,N_6787);
nand U8530 (N_8530,N_7647,N_7437);
or U8531 (N_8531,N_6206,N_6631);
nand U8532 (N_8532,N_7510,N_7349);
nand U8533 (N_8533,N_6565,N_6715);
and U8534 (N_8534,N_6488,N_7688);
nand U8535 (N_8535,N_7891,N_7458);
nor U8536 (N_8536,N_6085,N_6130);
or U8537 (N_8537,N_7535,N_7965);
nand U8538 (N_8538,N_6153,N_7410);
xnor U8539 (N_8539,N_6029,N_7507);
nand U8540 (N_8540,N_6674,N_6097);
nand U8541 (N_8541,N_7809,N_7642);
nor U8542 (N_8542,N_6828,N_6229);
or U8543 (N_8543,N_6870,N_7953);
nor U8544 (N_8544,N_7270,N_6366);
and U8545 (N_8545,N_7892,N_6163);
nor U8546 (N_8546,N_7456,N_7874);
or U8547 (N_8547,N_7148,N_7151);
nand U8548 (N_8548,N_7802,N_7789);
nand U8549 (N_8549,N_7378,N_7585);
nand U8550 (N_8550,N_7992,N_7380);
nor U8551 (N_8551,N_7183,N_6662);
nand U8552 (N_8552,N_6741,N_6574);
and U8553 (N_8553,N_6434,N_6770);
nand U8554 (N_8554,N_7232,N_7777);
or U8555 (N_8555,N_7831,N_6340);
or U8556 (N_8556,N_6318,N_6272);
or U8557 (N_8557,N_6086,N_7607);
and U8558 (N_8558,N_7040,N_6653);
or U8559 (N_8559,N_6976,N_7419);
nand U8560 (N_8560,N_7046,N_7515);
and U8561 (N_8561,N_6140,N_6815);
nand U8562 (N_8562,N_6326,N_6797);
and U8563 (N_8563,N_7674,N_7184);
nand U8564 (N_8564,N_7165,N_7370);
nand U8565 (N_8565,N_6669,N_7573);
and U8566 (N_8566,N_7466,N_7677);
and U8567 (N_8567,N_6316,N_6139);
xor U8568 (N_8568,N_7798,N_7632);
or U8569 (N_8569,N_7966,N_6792);
nand U8570 (N_8570,N_7167,N_7338);
and U8571 (N_8571,N_7847,N_7839);
or U8572 (N_8572,N_6244,N_7990);
or U8573 (N_8573,N_7227,N_7984);
nor U8574 (N_8574,N_6685,N_6682);
nor U8575 (N_8575,N_7115,N_6282);
nor U8576 (N_8576,N_7932,N_7513);
and U8577 (N_8577,N_6587,N_6035);
or U8578 (N_8578,N_6790,N_6755);
nor U8579 (N_8579,N_7323,N_6676);
and U8580 (N_8580,N_6027,N_7146);
or U8581 (N_8581,N_6748,N_6379);
and U8582 (N_8582,N_6794,N_6532);
nand U8583 (N_8583,N_6952,N_6558);
or U8584 (N_8584,N_7721,N_7058);
nor U8585 (N_8585,N_6312,N_7000);
or U8586 (N_8586,N_6410,N_6502);
and U8587 (N_8587,N_6364,N_6847);
nor U8588 (N_8588,N_6295,N_7004);
nor U8589 (N_8589,N_6151,N_7715);
nor U8590 (N_8590,N_6146,N_6430);
nand U8591 (N_8591,N_7474,N_6960);
and U8592 (N_8592,N_6625,N_6971);
or U8593 (N_8593,N_6937,N_7225);
nand U8594 (N_8594,N_6996,N_7766);
or U8595 (N_8595,N_7627,N_6982);
and U8596 (N_8596,N_6278,N_6145);
or U8597 (N_8597,N_6724,N_7562);
and U8598 (N_8598,N_6277,N_6651);
or U8599 (N_8599,N_6699,N_7646);
xor U8600 (N_8600,N_7070,N_7433);
nor U8601 (N_8601,N_6127,N_6116);
or U8602 (N_8602,N_6233,N_6238);
and U8603 (N_8603,N_7622,N_6970);
nor U8604 (N_8604,N_7903,N_6313);
nand U8605 (N_8605,N_6420,N_6895);
or U8606 (N_8606,N_6780,N_6380);
and U8607 (N_8607,N_6411,N_7385);
nand U8608 (N_8608,N_7567,N_7968);
nor U8609 (N_8609,N_7628,N_7367);
and U8610 (N_8610,N_6148,N_6656);
or U8611 (N_8611,N_7806,N_7132);
nor U8612 (N_8612,N_7611,N_6303);
nand U8613 (N_8613,N_7166,N_6461);
nor U8614 (N_8614,N_7312,N_6257);
nand U8615 (N_8615,N_7967,N_6886);
nor U8616 (N_8616,N_7858,N_6124);
or U8617 (N_8617,N_6079,N_6311);
or U8618 (N_8618,N_6406,N_6752);
or U8619 (N_8619,N_6076,N_6466);
or U8620 (N_8620,N_7914,N_7311);
nor U8621 (N_8621,N_7009,N_7429);
nand U8622 (N_8622,N_7450,N_7300);
and U8623 (N_8623,N_6480,N_7569);
and U8624 (N_8624,N_6909,N_7140);
and U8625 (N_8625,N_6938,N_6001);
nand U8626 (N_8626,N_6834,N_6396);
and U8627 (N_8627,N_6011,N_7963);
nand U8628 (N_8628,N_6216,N_6516);
nand U8629 (N_8629,N_7304,N_7574);
nor U8630 (N_8630,N_6421,N_6034);
or U8631 (N_8631,N_7170,N_7395);
nand U8632 (N_8632,N_7746,N_7601);
nor U8633 (N_8633,N_6675,N_6177);
nand U8634 (N_8634,N_7659,N_6404);
and U8635 (N_8635,N_7835,N_6370);
nand U8636 (N_8636,N_6588,N_6883);
or U8637 (N_8637,N_7110,N_7671);
or U8638 (N_8638,N_7572,N_6290);
and U8639 (N_8639,N_7995,N_6530);
and U8640 (N_8640,N_6251,N_6343);
nor U8641 (N_8641,N_7561,N_6912);
and U8642 (N_8642,N_7428,N_6592);
and U8643 (N_8643,N_6059,N_7741);
nor U8644 (N_8644,N_6602,N_6405);
nand U8645 (N_8645,N_7368,N_6224);
nand U8646 (N_8646,N_6186,N_7877);
nor U8647 (N_8647,N_7733,N_6054);
nand U8648 (N_8648,N_6062,N_7138);
or U8649 (N_8649,N_6373,N_7461);
nor U8650 (N_8650,N_6230,N_6629);
nor U8651 (N_8651,N_7263,N_7697);
nand U8652 (N_8652,N_6103,N_6630);
or U8653 (N_8653,N_6539,N_7680);
nand U8654 (N_8654,N_6324,N_7770);
and U8655 (N_8655,N_6460,N_7201);
nor U8656 (N_8656,N_6479,N_6655);
nor U8657 (N_8657,N_7013,N_6929);
or U8658 (N_8658,N_7069,N_6032);
and U8659 (N_8659,N_6906,N_7038);
nand U8660 (N_8660,N_6773,N_6601);
nand U8661 (N_8661,N_6553,N_6512);
and U8662 (N_8662,N_7041,N_7332);
nand U8663 (N_8663,N_6838,N_6772);
nand U8664 (N_8664,N_6375,N_7264);
nor U8665 (N_8665,N_7540,N_7081);
nand U8666 (N_8666,N_6931,N_6028);
and U8667 (N_8667,N_7763,N_7105);
nor U8668 (N_8668,N_6408,N_7045);
and U8669 (N_8669,N_6237,N_7291);
or U8670 (N_8670,N_7267,N_6174);
or U8671 (N_8671,N_7818,N_7214);
and U8672 (N_8672,N_7684,N_7137);
or U8673 (N_8673,N_7781,N_7686);
and U8674 (N_8674,N_7991,N_7959);
or U8675 (N_8675,N_6149,N_7226);
and U8676 (N_8676,N_6527,N_7087);
and U8677 (N_8677,N_6683,N_6167);
nand U8678 (N_8678,N_6915,N_7402);
or U8679 (N_8679,N_7977,N_6681);
nand U8680 (N_8680,N_6720,N_7473);
nor U8681 (N_8681,N_7558,N_7116);
and U8682 (N_8682,N_7582,N_7251);
nor U8683 (N_8683,N_6966,N_6921);
or U8684 (N_8684,N_7359,N_7143);
nor U8685 (N_8685,N_7533,N_6934);
nand U8686 (N_8686,N_7570,N_7918);
or U8687 (N_8687,N_7832,N_6357);
or U8688 (N_8688,N_7614,N_6978);
nor U8689 (N_8689,N_7001,N_6319);
nand U8690 (N_8690,N_6583,N_7813);
nand U8691 (N_8691,N_6542,N_6888);
or U8692 (N_8692,N_7833,N_7136);
nor U8693 (N_8693,N_6526,N_6948);
nor U8694 (N_8694,N_7755,N_7972);
or U8695 (N_8695,N_7819,N_7635);
or U8696 (N_8696,N_6038,N_6858);
nand U8697 (N_8697,N_6274,N_6965);
nor U8698 (N_8698,N_7630,N_6242);
nor U8699 (N_8699,N_6570,N_7623);
and U8700 (N_8700,N_6236,N_7413);
and U8701 (N_8701,N_6578,N_7454);
nor U8702 (N_8702,N_6825,N_6468);
nor U8703 (N_8703,N_6837,N_6637);
and U8704 (N_8704,N_7271,N_7902);
nor U8705 (N_8705,N_6240,N_7059);
and U8706 (N_8706,N_6719,N_7285);
and U8707 (N_8707,N_7448,N_7366);
nor U8708 (N_8708,N_6711,N_6990);
and U8709 (N_8709,N_7857,N_7521);
and U8710 (N_8710,N_6958,N_6108);
nor U8711 (N_8711,N_6400,N_6897);
or U8712 (N_8712,N_6263,N_7708);
or U8713 (N_8713,N_6819,N_7407);
nor U8714 (N_8714,N_6688,N_6568);
and U8715 (N_8715,N_7282,N_7195);
nand U8716 (N_8716,N_7711,N_7443);
and U8717 (N_8717,N_6551,N_6820);
and U8718 (N_8718,N_6968,N_7811);
nor U8719 (N_8719,N_7102,N_6944);
nor U8720 (N_8720,N_6880,N_7212);
and U8721 (N_8721,N_7345,N_7122);
or U8722 (N_8722,N_7394,N_6789);
or U8723 (N_8723,N_7864,N_6585);
nor U8724 (N_8724,N_6750,N_6123);
nor U8725 (N_8725,N_6951,N_6902);
nand U8726 (N_8726,N_7269,N_6162);
and U8727 (N_8727,N_6613,N_6161);
or U8728 (N_8728,N_7185,N_7782);
nand U8729 (N_8729,N_6806,N_6846);
nand U8730 (N_8730,N_7056,N_7218);
nor U8731 (N_8731,N_7492,N_6851);
nand U8732 (N_8732,N_6013,N_7416);
nor U8733 (N_8733,N_6899,N_6443);
nor U8734 (N_8734,N_7694,N_6932);
nor U8735 (N_8735,N_7531,N_7765);
nand U8736 (N_8736,N_6046,N_6520);
or U8737 (N_8737,N_6955,N_7633);
and U8738 (N_8738,N_6060,N_6600);
and U8739 (N_8739,N_7978,N_6456);
and U8740 (N_8740,N_6068,N_6268);
nand U8741 (N_8741,N_7206,N_7217);
or U8742 (N_8742,N_6830,N_6627);
nor U8743 (N_8743,N_7778,N_7017);
nor U8744 (N_8744,N_6307,N_7934);
or U8745 (N_8745,N_6580,N_7759);
and U8746 (N_8746,N_7619,N_7432);
and U8747 (N_8747,N_7719,N_6334);
nor U8748 (N_8748,N_7112,N_7843);
nor U8749 (N_8749,N_6201,N_6009);
or U8750 (N_8750,N_6754,N_7529);
nor U8751 (N_8751,N_7104,N_6156);
or U8752 (N_8752,N_6679,N_6901);
and U8753 (N_8753,N_6919,N_6083);
nor U8754 (N_8754,N_6017,N_6640);
nand U8755 (N_8755,N_6549,N_7656);
and U8756 (N_8756,N_6771,N_6826);
or U8757 (N_8757,N_6300,N_6452);
nor U8758 (N_8758,N_7807,N_6065);
or U8759 (N_8759,N_6100,N_7127);
and U8760 (N_8760,N_7156,N_7231);
nand U8761 (N_8761,N_7681,N_6809);
and U8762 (N_8762,N_6763,N_6514);
and U8763 (N_8763,N_7612,N_6071);
and U8764 (N_8764,N_6299,N_6988);
nand U8765 (N_8765,N_7106,N_7369);
nor U8766 (N_8766,N_6564,N_7221);
and U8767 (N_8767,N_7159,N_7005);
and U8768 (N_8768,N_6447,N_6454);
and U8769 (N_8769,N_6198,N_7340);
nor U8770 (N_8770,N_6749,N_6137);
and U8771 (N_8771,N_6037,N_7962);
nor U8772 (N_8772,N_6818,N_6701);
or U8773 (N_8773,N_7822,N_6796);
and U8774 (N_8774,N_7930,N_7889);
or U8775 (N_8775,N_7130,N_6425);
nor U8776 (N_8776,N_6974,N_6727);
and U8777 (N_8777,N_6557,N_7356);
nand U8778 (N_8778,N_6317,N_6786);
nor U8779 (N_8779,N_7153,N_6645);
nand U8780 (N_8780,N_6941,N_6368);
nor U8781 (N_8781,N_7052,N_6910);
and U8782 (N_8782,N_6287,N_7318);
and U8783 (N_8783,N_6112,N_7885);
or U8784 (N_8784,N_7520,N_7211);
or U8785 (N_8785,N_7262,N_7336);
nor U8786 (N_8786,N_6700,N_6504);
and U8787 (N_8787,N_6301,N_6467);
nand U8788 (N_8788,N_6072,N_7731);
or U8789 (N_8789,N_7006,N_6868);
or U8790 (N_8790,N_7192,N_6057);
nor U8791 (N_8791,N_7333,N_6154);
xor U8792 (N_8792,N_6215,N_6876);
nand U8793 (N_8793,N_7124,N_6762);
nand U8794 (N_8794,N_6881,N_6255);
nor U8795 (N_8795,N_7997,N_6374);
and U8796 (N_8796,N_7541,N_7382);
nand U8797 (N_8797,N_7849,N_7090);
nor U8798 (N_8798,N_7576,N_6535);
or U8799 (N_8799,N_6597,N_7901);
nor U8800 (N_8800,N_7031,N_6767);
and U8801 (N_8801,N_6498,N_6515);
nand U8802 (N_8802,N_6191,N_7387);
or U8803 (N_8803,N_6044,N_7465);
or U8804 (N_8804,N_6882,N_6351);
nand U8805 (N_8805,N_6087,N_6836);
and U8806 (N_8806,N_7314,N_7411);
nor U8807 (N_8807,N_7638,N_6654);
and U8808 (N_8808,N_6827,N_7812);
and U8809 (N_8809,N_6260,N_6618);
nand U8810 (N_8810,N_6785,N_6612);
or U8811 (N_8811,N_6002,N_6730);
nor U8812 (N_8812,N_7241,N_6800);
or U8813 (N_8813,N_6228,N_6878);
nand U8814 (N_8814,N_6051,N_7530);
nor U8815 (N_8815,N_6195,N_7926);
and U8816 (N_8816,N_7584,N_7869);
and U8817 (N_8817,N_7853,N_7925);
nor U8818 (N_8818,N_6566,N_6323);
nor U8819 (N_8819,N_6761,N_6987);
nor U8820 (N_8820,N_7888,N_7177);
nand U8821 (N_8821,N_6448,N_7559);
or U8822 (N_8822,N_7215,N_6747);
nand U8823 (N_8823,N_7049,N_6042);
nor U8824 (N_8824,N_6172,N_7931);
nor U8825 (N_8825,N_7629,N_6562);
nor U8826 (N_8826,N_6297,N_7108);
or U8827 (N_8827,N_7698,N_7928);
and U8828 (N_8828,N_7577,N_7790);
nand U8829 (N_8829,N_7415,N_7728);
and U8830 (N_8830,N_7498,N_7916);
nand U8831 (N_8831,N_6331,N_7894);
nand U8832 (N_8832,N_7275,N_7593);
xnor U8833 (N_8833,N_6709,N_7431);
and U8834 (N_8834,N_7524,N_7616);
and U8835 (N_8835,N_7605,N_6199);
and U8836 (N_8836,N_6142,N_7842);
xor U8837 (N_8837,N_6521,N_7691);
nor U8838 (N_8838,N_6964,N_6429);
nand U8839 (N_8839,N_6241,N_6593);
nor U8840 (N_8840,N_6664,N_6993);
nand U8841 (N_8841,N_7608,N_7970);
or U8842 (N_8842,N_7937,N_6768);
or U8843 (N_8843,N_6007,N_6254);
nand U8844 (N_8844,N_6736,N_6220);
nor U8845 (N_8845,N_6275,N_6998);
nand U8846 (N_8846,N_6956,N_6475);
and U8847 (N_8847,N_6393,N_7710);
or U8848 (N_8848,N_7256,N_6781);
or U8849 (N_8849,N_6407,N_7067);
nand U8850 (N_8850,N_7905,N_6099);
and U8851 (N_8851,N_6328,N_6804);
or U8852 (N_8852,N_7505,N_7305);
or U8853 (N_8853,N_6764,N_7235);
or U8854 (N_8854,N_6614,N_7290);
nor U8855 (N_8855,N_7704,N_6356);
nand U8856 (N_8856,N_6610,N_6703);
nor U8857 (N_8857,N_6854,N_6511);
and U8858 (N_8858,N_7375,N_7348);
nand U8859 (N_8859,N_6390,N_7139);
nor U8860 (N_8860,N_7828,N_6636);
and U8861 (N_8861,N_7024,N_7497);
nor U8862 (N_8862,N_7974,N_7554);
nor U8863 (N_8863,N_7021,N_6693);
xor U8864 (N_8864,N_7921,N_7730);
nand U8865 (N_8865,N_6223,N_6579);
or U8866 (N_8866,N_7401,N_7866);
nor U8867 (N_8867,N_6923,N_6795);
or U8868 (N_8868,N_7706,N_6385);
or U8869 (N_8869,N_7365,N_7224);
nor U8870 (N_8870,N_6714,N_6835);
or U8871 (N_8871,N_6575,N_6814);
nand U8872 (N_8872,N_7476,N_7057);
or U8873 (N_8873,N_7249,N_6435);
nand U8874 (N_8874,N_6538,N_7957);
and U8875 (N_8875,N_7738,N_6284);
nor U8876 (N_8876,N_6388,N_7425);
or U8877 (N_8877,N_7592,N_7961);
nor U8878 (N_8878,N_6440,N_6505);
or U8879 (N_8879,N_7571,N_6183);
nand U8880 (N_8880,N_7854,N_7398);
nand U8881 (N_8881,N_7084,N_6286);
and U8882 (N_8882,N_6947,N_7292);
and U8883 (N_8883,N_7364,N_6128);
and U8884 (N_8884,N_6799,N_6760);
or U8885 (N_8885,N_7103,N_6619);
and U8886 (N_8886,N_7602,N_6453);
nor U8887 (N_8887,N_7537,N_6734);
nand U8888 (N_8888,N_6697,N_7464);
or U8889 (N_8889,N_7870,N_7499);
and U8890 (N_8890,N_7779,N_7029);
and U8891 (N_8891,N_7845,N_7895);
or U8892 (N_8892,N_7951,N_6843);
nor U8893 (N_8893,N_6793,N_6239);
nand U8894 (N_8894,N_6472,N_6113);
and U8895 (N_8895,N_7092,N_7950);
or U8896 (N_8896,N_6507,N_7207);
nand U8897 (N_8897,N_6095,N_7768);
nand U8898 (N_8898,N_7514,N_6540);
nor U8899 (N_8899,N_6898,N_7528);
nand U8900 (N_8900,N_6090,N_6332);
nor U8901 (N_8901,N_7036,N_7054);
nor U8902 (N_8902,N_7898,N_7838);
nor U8903 (N_8903,N_6778,N_6890);
nand U8904 (N_8904,N_6045,N_7580);
and U8905 (N_8905,N_6712,N_7823);
nand U8906 (N_8906,N_6552,N_7651);
and U8907 (N_8907,N_6707,N_6184);
or U8908 (N_8908,N_6877,N_6666);
or U8909 (N_8909,N_7035,N_6561);
nand U8910 (N_8910,N_7655,N_6482);
nand U8911 (N_8911,N_6604,N_6528);
and U8912 (N_8912,N_7294,N_6994);
and U8913 (N_8913,N_7403,N_6667);
and U8914 (N_8914,N_6330,N_7033);
nor U8915 (N_8915,N_6403,N_7801);
nand U8916 (N_8916,N_7334,N_7455);
and U8917 (N_8917,N_7042,N_6457);
nand U8918 (N_8918,N_6347,N_6458);
and U8919 (N_8919,N_6451,N_7255);
nand U8920 (N_8920,N_7773,N_6392);
or U8921 (N_8921,N_6529,N_6873);
or U8922 (N_8922,N_7855,N_6030);
and U8923 (N_8923,N_6227,N_7884);
nor U8924 (N_8924,N_7309,N_6064);
or U8925 (N_8925,N_7233,N_7664);
nor U8926 (N_8926,N_6648,N_6026);
nor U8927 (N_8927,N_6101,N_7298);
and U8928 (N_8928,N_7669,N_7548);
and U8929 (N_8929,N_6320,N_6235);
or U8930 (N_8930,N_6865,N_7816);
or U8931 (N_8931,N_6093,N_6633);
and U8932 (N_8932,N_7325,N_7308);
and U8933 (N_8933,N_6605,N_6884);
and U8934 (N_8934,N_7276,N_7154);
nor U8935 (N_8935,N_7397,N_7893);
or U8936 (N_8936,N_7683,N_6595);
or U8937 (N_8937,N_7469,N_7940);
or U8938 (N_8938,N_7969,N_6247);
nor U8939 (N_8939,N_6189,N_7026);
and U8940 (N_8940,N_6875,N_6673);
nand U8941 (N_8941,N_6418,N_7187);
and U8942 (N_8942,N_6871,N_6560);
nand U8943 (N_8943,N_7216,N_7859);
nor U8944 (N_8944,N_7661,N_7287);
and U8945 (N_8945,N_7075,N_7150);
nand U8946 (N_8946,N_6160,N_7246);
nor U8947 (N_8947,N_6481,N_7624);
nor U8948 (N_8948,N_6811,N_6708);
or U8949 (N_8949,N_6218,N_6706);
nor U8950 (N_8950,N_6740,N_6782);
or U8951 (N_8951,N_7101,N_7649);
and U8952 (N_8952,N_7272,N_6036);
and U8953 (N_8953,N_6979,N_7034);
nand U8954 (N_8954,N_7010,N_7799);
nand U8955 (N_8955,N_7747,N_7547);
nor U8956 (N_8956,N_6821,N_7011);
and U8957 (N_8957,N_7480,N_6517);
nor U8958 (N_8958,N_7867,N_6143);
nor U8959 (N_8959,N_6412,N_7935);
nand U8960 (N_8960,N_7155,N_7876);
nor U8961 (N_8961,N_6118,N_7331);
and U8962 (N_8962,N_7971,N_7060);
nor U8963 (N_8963,N_7449,N_6999);
or U8964 (N_8964,N_7508,N_7301);
nor U8965 (N_8965,N_6416,N_7435);
nand U8966 (N_8966,N_7273,N_6131);
and U8967 (N_8967,N_7587,N_7543);
and U8968 (N_8968,N_6624,N_7511);
nand U8969 (N_8969,N_7900,N_6537);
or U8970 (N_8970,N_6856,N_7080);
or U8971 (N_8971,N_7141,N_6376);
nand U8972 (N_8972,N_6900,N_6485);
nor U8973 (N_8973,N_7441,N_6721);
nand U8974 (N_8974,N_6476,N_7764);
nand U8975 (N_8975,N_6261,N_7310);
or U8976 (N_8976,N_7929,N_6021);
or U8977 (N_8977,N_6967,N_7989);
nor U8978 (N_8978,N_7213,N_6150);
or U8979 (N_8979,N_7685,N_7400);
nor U8980 (N_8980,N_6424,N_6986);
or U8981 (N_8981,N_6279,N_6117);
nand U8982 (N_8982,N_7805,N_6187);
or U8983 (N_8983,N_7085,N_7061);
or U8984 (N_8984,N_7030,N_7695);
nor U8985 (N_8985,N_7713,N_6758);
or U8986 (N_8986,N_6281,N_6936);
or U8987 (N_8987,N_6144,N_6371);
nor U8988 (N_8988,N_7220,N_6726);
and U8989 (N_8989,N_6061,N_6018);
or U8990 (N_8990,N_7886,N_7652);
and U8991 (N_8991,N_7555,N_6670);
and U8992 (N_8992,N_6040,N_7954);
or U8993 (N_8993,N_6088,N_7837);
and U8994 (N_8994,N_6074,N_7752);
or U8995 (N_8995,N_7793,N_6211);
or U8996 (N_8996,N_6914,N_7179);
nand U8997 (N_8997,N_6571,N_6962);
nor U8998 (N_8998,N_6791,N_7786);
and U8999 (N_8999,N_7879,N_7732);
nand U9000 (N_9000,N_6804,N_6338);
nor U9001 (N_9001,N_6974,N_6747);
or U9002 (N_9002,N_7885,N_6710);
nand U9003 (N_9003,N_7463,N_7901);
nor U9004 (N_9004,N_7086,N_7360);
nand U9005 (N_9005,N_6062,N_6648);
nor U9006 (N_9006,N_6441,N_6184);
or U9007 (N_9007,N_6085,N_6260);
nand U9008 (N_9008,N_6412,N_7856);
or U9009 (N_9009,N_7863,N_6330);
nand U9010 (N_9010,N_7903,N_6936);
nand U9011 (N_9011,N_7555,N_6390);
or U9012 (N_9012,N_7661,N_7473);
and U9013 (N_9013,N_7187,N_6326);
nor U9014 (N_9014,N_6878,N_7258);
nor U9015 (N_9015,N_6499,N_7795);
nand U9016 (N_9016,N_6308,N_7437);
nor U9017 (N_9017,N_6125,N_6623);
nor U9018 (N_9018,N_7792,N_7114);
or U9019 (N_9019,N_7153,N_7767);
xnor U9020 (N_9020,N_6441,N_7162);
or U9021 (N_9021,N_6582,N_6806);
or U9022 (N_9022,N_6800,N_7428);
or U9023 (N_9023,N_7881,N_6793);
and U9024 (N_9024,N_6744,N_7538);
and U9025 (N_9025,N_7672,N_6710);
nor U9026 (N_9026,N_6008,N_7025);
nand U9027 (N_9027,N_7369,N_6693);
nor U9028 (N_9028,N_7373,N_6213);
nor U9029 (N_9029,N_6157,N_7079);
and U9030 (N_9030,N_6350,N_6977);
nand U9031 (N_9031,N_6704,N_6534);
nand U9032 (N_9032,N_6767,N_7264);
or U9033 (N_9033,N_6337,N_7073);
nand U9034 (N_9034,N_7399,N_7360);
nand U9035 (N_9035,N_6575,N_6317);
or U9036 (N_9036,N_6301,N_7544);
nand U9037 (N_9037,N_6821,N_6855);
or U9038 (N_9038,N_6038,N_6556);
or U9039 (N_9039,N_6088,N_6886);
and U9040 (N_9040,N_6890,N_7977);
nand U9041 (N_9041,N_6618,N_7429);
and U9042 (N_9042,N_7727,N_7640);
and U9043 (N_9043,N_6086,N_6580);
or U9044 (N_9044,N_6757,N_7960);
or U9045 (N_9045,N_7299,N_7190);
nand U9046 (N_9046,N_6221,N_6832);
nor U9047 (N_9047,N_6653,N_6426);
nor U9048 (N_9048,N_7160,N_6930);
nand U9049 (N_9049,N_6613,N_7168);
and U9050 (N_9050,N_6904,N_6071);
or U9051 (N_9051,N_6008,N_6283);
nand U9052 (N_9052,N_7676,N_7007);
nor U9053 (N_9053,N_6624,N_7458);
and U9054 (N_9054,N_7559,N_6753);
nand U9055 (N_9055,N_7624,N_7532);
or U9056 (N_9056,N_7658,N_7115);
or U9057 (N_9057,N_6928,N_7975);
nor U9058 (N_9058,N_7653,N_7901);
nor U9059 (N_9059,N_6113,N_7799);
nand U9060 (N_9060,N_7540,N_7303);
nor U9061 (N_9061,N_7696,N_6394);
nand U9062 (N_9062,N_6713,N_7961);
nor U9063 (N_9063,N_7070,N_6731);
nand U9064 (N_9064,N_7280,N_6115);
and U9065 (N_9065,N_7114,N_7418);
or U9066 (N_9066,N_6817,N_6704);
or U9067 (N_9067,N_7895,N_7301);
nor U9068 (N_9068,N_7211,N_6102);
nor U9069 (N_9069,N_7064,N_7553);
or U9070 (N_9070,N_6773,N_6613);
nand U9071 (N_9071,N_7129,N_6881);
and U9072 (N_9072,N_6710,N_6763);
nand U9073 (N_9073,N_6764,N_7576);
and U9074 (N_9074,N_6318,N_6589);
nor U9075 (N_9075,N_6909,N_7097);
nor U9076 (N_9076,N_6288,N_7077);
nor U9077 (N_9077,N_7326,N_6099);
or U9078 (N_9078,N_7718,N_7645);
or U9079 (N_9079,N_6437,N_6407);
nand U9080 (N_9080,N_6620,N_6313);
and U9081 (N_9081,N_6622,N_7935);
nand U9082 (N_9082,N_7201,N_6699);
or U9083 (N_9083,N_6554,N_7808);
nand U9084 (N_9084,N_6556,N_6791);
or U9085 (N_9085,N_6991,N_6705);
or U9086 (N_9086,N_6778,N_6148);
or U9087 (N_9087,N_7077,N_6122);
and U9088 (N_9088,N_6810,N_6803);
and U9089 (N_9089,N_7881,N_6863);
and U9090 (N_9090,N_7269,N_7294);
nor U9091 (N_9091,N_7702,N_7480);
and U9092 (N_9092,N_7067,N_7312);
and U9093 (N_9093,N_7275,N_7082);
nor U9094 (N_9094,N_7499,N_7707);
nand U9095 (N_9095,N_6875,N_6301);
or U9096 (N_9096,N_6837,N_6282);
nor U9097 (N_9097,N_7818,N_7649);
and U9098 (N_9098,N_7508,N_6266);
and U9099 (N_9099,N_6205,N_7126);
and U9100 (N_9100,N_7921,N_7314);
nor U9101 (N_9101,N_6938,N_7829);
and U9102 (N_9102,N_7397,N_6007);
or U9103 (N_9103,N_7383,N_7435);
nor U9104 (N_9104,N_7711,N_7318);
or U9105 (N_9105,N_7660,N_6215);
or U9106 (N_9106,N_6852,N_6249);
nor U9107 (N_9107,N_6820,N_6429);
or U9108 (N_9108,N_6916,N_6754);
nand U9109 (N_9109,N_7590,N_6570);
and U9110 (N_9110,N_6511,N_7273);
or U9111 (N_9111,N_6684,N_6693);
or U9112 (N_9112,N_6018,N_6657);
nand U9113 (N_9113,N_6709,N_6411);
and U9114 (N_9114,N_6182,N_7196);
nand U9115 (N_9115,N_6942,N_6076);
or U9116 (N_9116,N_6035,N_7491);
or U9117 (N_9117,N_6814,N_6106);
nor U9118 (N_9118,N_6819,N_7672);
and U9119 (N_9119,N_6553,N_7386);
nand U9120 (N_9120,N_6751,N_6732);
nor U9121 (N_9121,N_6783,N_7396);
or U9122 (N_9122,N_7984,N_7494);
xor U9123 (N_9123,N_7990,N_6230);
and U9124 (N_9124,N_7354,N_7972);
or U9125 (N_9125,N_7091,N_7230);
nand U9126 (N_9126,N_7458,N_6960);
and U9127 (N_9127,N_6485,N_7406);
nor U9128 (N_9128,N_7087,N_6777);
nand U9129 (N_9129,N_6146,N_6440);
or U9130 (N_9130,N_7229,N_6210);
nand U9131 (N_9131,N_7026,N_6715);
or U9132 (N_9132,N_7652,N_6396);
and U9133 (N_9133,N_6424,N_6755);
or U9134 (N_9134,N_6542,N_7832);
and U9135 (N_9135,N_6057,N_6933);
or U9136 (N_9136,N_7696,N_6760);
or U9137 (N_9137,N_7021,N_7621);
nand U9138 (N_9138,N_7172,N_6148);
xor U9139 (N_9139,N_6896,N_7903);
or U9140 (N_9140,N_6938,N_7440);
and U9141 (N_9141,N_7272,N_7066);
nand U9142 (N_9142,N_6249,N_7595);
or U9143 (N_9143,N_6663,N_6347);
or U9144 (N_9144,N_7263,N_7264);
and U9145 (N_9145,N_7724,N_7768);
and U9146 (N_9146,N_6472,N_6135);
or U9147 (N_9147,N_6634,N_7566);
and U9148 (N_9148,N_7977,N_7806);
or U9149 (N_9149,N_7696,N_6020);
and U9150 (N_9150,N_6555,N_7000);
or U9151 (N_9151,N_7148,N_7378);
nor U9152 (N_9152,N_6171,N_6531);
nor U9153 (N_9153,N_6681,N_7343);
nor U9154 (N_9154,N_6178,N_6254);
or U9155 (N_9155,N_7972,N_7611);
nand U9156 (N_9156,N_6864,N_6457);
or U9157 (N_9157,N_6026,N_6881);
nand U9158 (N_9158,N_6018,N_7631);
xnor U9159 (N_9159,N_6154,N_7917);
xnor U9160 (N_9160,N_7325,N_6083);
and U9161 (N_9161,N_7136,N_6984);
or U9162 (N_9162,N_6464,N_7145);
or U9163 (N_9163,N_6896,N_6774);
nand U9164 (N_9164,N_6101,N_6047);
and U9165 (N_9165,N_6911,N_6085);
nand U9166 (N_9166,N_7491,N_7246);
nand U9167 (N_9167,N_7809,N_7840);
and U9168 (N_9168,N_7645,N_7501);
and U9169 (N_9169,N_6396,N_7255);
or U9170 (N_9170,N_7176,N_7918);
and U9171 (N_9171,N_6833,N_6388);
nor U9172 (N_9172,N_7583,N_6924);
nor U9173 (N_9173,N_6717,N_7273);
and U9174 (N_9174,N_7978,N_6826);
or U9175 (N_9175,N_6437,N_7763);
and U9176 (N_9176,N_7023,N_7750);
and U9177 (N_9177,N_7903,N_6150);
or U9178 (N_9178,N_6512,N_7405);
nand U9179 (N_9179,N_7021,N_6018);
or U9180 (N_9180,N_7188,N_7994);
or U9181 (N_9181,N_6466,N_6015);
nor U9182 (N_9182,N_7770,N_6499);
or U9183 (N_9183,N_6822,N_6777);
and U9184 (N_9184,N_6592,N_6927);
nand U9185 (N_9185,N_7603,N_6482);
nand U9186 (N_9186,N_7375,N_6896);
nand U9187 (N_9187,N_6854,N_7512);
nand U9188 (N_9188,N_7746,N_7815);
nor U9189 (N_9189,N_7573,N_7581);
nor U9190 (N_9190,N_7113,N_6826);
or U9191 (N_9191,N_7665,N_7393);
nand U9192 (N_9192,N_7559,N_7157);
nand U9193 (N_9193,N_6882,N_7862);
nand U9194 (N_9194,N_6611,N_6508);
nor U9195 (N_9195,N_6016,N_7755);
nand U9196 (N_9196,N_6374,N_7201);
nor U9197 (N_9197,N_7234,N_7235);
or U9198 (N_9198,N_6596,N_7650);
nor U9199 (N_9199,N_6814,N_7989);
and U9200 (N_9200,N_6825,N_6767);
nor U9201 (N_9201,N_7636,N_6353);
nand U9202 (N_9202,N_6508,N_6043);
nand U9203 (N_9203,N_6076,N_7381);
nor U9204 (N_9204,N_7482,N_6144);
and U9205 (N_9205,N_7750,N_6929);
nand U9206 (N_9206,N_7461,N_7520);
nand U9207 (N_9207,N_6544,N_6528);
nand U9208 (N_9208,N_7496,N_6878);
and U9209 (N_9209,N_6327,N_6641);
or U9210 (N_9210,N_6315,N_7936);
nand U9211 (N_9211,N_7224,N_6900);
and U9212 (N_9212,N_6707,N_7897);
nand U9213 (N_9213,N_6600,N_6866);
nor U9214 (N_9214,N_7303,N_7167);
nor U9215 (N_9215,N_6531,N_6332);
and U9216 (N_9216,N_6301,N_7569);
and U9217 (N_9217,N_6582,N_6526);
and U9218 (N_9218,N_7333,N_6295);
or U9219 (N_9219,N_6565,N_7373);
nand U9220 (N_9220,N_7303,N_6595);
nor U9221 (N_9221,N_7519,N_7341);
nor U9222 (N_9222,N_6583,N_7830);
nand U9223 (N_9223,N_6240,N_6347);
or U9224 (N_9224,N_6787,N_6577);
and U9225 (N_9225,N_6877,N_6573);
and U9226 (N_9226,N_7045,N_7922);
or U9227 (N_9227,N_6655,N_7825);
nor U9228 (N_9228,N_7183,N_7255);
or U9229 (N_9229,N_7166,N_7175);
and U9230 (N_9230,N_6116,N_6967);
nor U9231 (N_9231,N_6287,N_6234);
xnor U9232 (N_9232,N_6613,N_7503);
or U9233 (N_9233,N_6321,N_6116);
and U9234 (N_9234,N_6819,N_7083);
nand U9235 (N_9235,N_7167,N_6435);
or U9236 (N_9236,N_6210,N_7141);
or U9237 (N_9237,N_6109,N_6821);
and U9238 (N_9238,N_7084,N_7766);
nor U9239 (N_9239,N_7488,N_7431);
nand U9240 (N_9240,N_6602,N_7595);
nor U9241 (N_9241,N_6024,N_7923);
or U9242 (N_9242,N_7596,N_6469);
nor U9243 (N_9243,N_6136,N_7268);
nand U9244 (N_9244,N_6111,N_6843);
or U9245 (N_9245,N_6994,N_6466);
nand U9246 (N_9246,N_7290,N_7285);
nor U9247 (N_9247,N_7633,N_7555);
nand U9248 (N_9248,N_6599,N_7543);
nand U9249 (N_9249,N_7694,N_7807);
or U9250 (N_9250,N_6059,N_7209);
nor U9251 (N_9251,N_7081,N_7401);
nand U9252 (N_9252,N_7664,N_7151);
nand U9253 (N_9253,N_6419,N_7939);
or U9254 (N_9254,N_7960,N_6083);
nor U9255 (N_9255,N_6478,N_6840);
nor U9256 (N_9256,N_7312,N_6439);
nor U9257 (N_9257,N_6075,N_7638);
xnor U9258 (N_9258,N_7104,N_6415);
nor U9259 (N_9259,N_7206,N_7976);
nand U9260 (N_9260,N_6292,N_7030);
and U9261 (N_9261,N_7828,N_7683);
nor U9262 (N_9262,N_7676,N_7170);
nand U9263 (N_9263,N_7774,N_6899);
nand U9264 (N_9264,N_7058,N_7757);
and U9265 (N_9265,N_6331,N_7541);
or U9266 (N_9266,N_7178,N_7626);
nor U9267 (N_9267,N_7405,N_6294);
nand U9268 (N_9268,N_6707,N_7257);
nand U9269 (N_9269,N_6803,N_6725);
nor U9270 (N_9270,N_7196,N_7560);
nor U9271 (N_9271,N_7783,N_7580);
or U9272 (N_9272,N_7655,N_6407);
and U9273 (N_9273,N_6946,N_7382);
or U9274 (N_9274,N_7099,N_6797);
nor U9275 (N_9275,N_6183,N_6364);
or U9276 (N_9276,N_6204,N_6947);
nor U9277 (N_9277,N_7932,N_7131);
and U9278 (N_9278,N_6137,N_7707);
or U9279 (N_9279,N_6701,N_7236);
or U9280 (N_9280,N_6091,N_7058);
nor U9281 (N_9281,N_6300,N_7274);
nor U9282 (N_9282,N_6721,N_6090);
and U9283 (N_9283,N_6689,N_6497);
nand U9284 (N_9284,N_6570,N_7030);
nand U9285 (N_9285,N_6756,N_6246);
or U9286 (N_9286,N_7329,N_7803);
or U9287 (N_9287,N_6213,N_6196);
nor U9288 (N_9288,N_6329,N_6771);
nand U9289 (N_9289,N_7907,N_6052);
nand U9290 (N_9290,N_7841,N_6141);
nor U9291 (N_9291,N_7844,N_6953);
or U9292 (N_9292,N_7987,N_7468);
and U9293 (N_9293,N_6211,N_7320);
nor U9294 (N_9294,N_7281,N_6469);
and U9295 (N_9295,N_7539,N_7315);
or U9296 (N_9296,N_6854,N_6961);
or U9297 (N_9297,N_6901,N_6340);
or U9298 (N_9298,N_6697,N_6296);
and U9299 (N_9299,N_6076,N_7646);
and U9300 (N_9300,N_6434,N_7656);
and U9301 (N_9301,N_7411,N_7052);
nand U9302 (N_9302,N_7823,N_7644);
or U9303 (N_9303,N_7859,N_7648);
and U9304 (N_9304,N_7498,N_7961);
nand U9305 (N_9305,N_6366,N_6259);
or U9306 (N_9306,N_7886,N_6915);
or U9307 (N_9307,N_7449,N_7145);
nand U9308 (N_9308,N_6811,N_6629);
or U9309 (N_9309,N_7258,N_6628);
or U9310 (N_9310,N_7627,N_6992);
nor U9311 (N_9311,N_6854,N_7488);
and U9312 (N_9312,N_7834,N_6380);
nor U9313 (N_9313,N_6757,N_7903);
nand U9314 (N_9314,N_6002,N_6444);
nor U9315 (N_9315,N_7797,N_7239);
and U9316 (N_9316,N_6037,N_6873);
and U9317 (N_9317,N_6192,N_7878);
and U9318 (N_9318,N_7418,N_6632);
and U9319 (N_9319,N_7714,N_6942);
nand U9320 (N_9320,N_7693,N_7075);
nand U9321 (N_9321,N_7354,N_6959);
or U9322 (N_9322,N_7268,N_7466);
or U9323 (N_9323,N_7904,N_7780);
or U9324 (N_9324,N_7139,N_6695);
or U9325 (N_9325,N_6219,N_6246);
or U9326 (N_9326,N_6101,N_7853);
nor U9327 (N_9327,N_7085,N_7580);
nand U9328 (N_9328,N_6145,N_7445);
or U9329 (N_9329,N_6818,N_6323);
and U9330 (N_9330,N_6081,N_7062);
and U9331 (N_9331,N_7280,N_6059);
or U9332 (N_9332,N_7930,N_6543);
and U9333 (N_9333,N_7768,N_6667);
and U9334 (N_9334,N_7663,N_6338);
nor U9335 (N_9335,N_7199,N_7462);
nand U9336 (N_9336,N_6823,N_6290);
and U9337 (N_9337,N_7179,N_6128);
and U9338 (N_9338,N_6842,N_7808);
and U9339 (N_9339,N_7096,N_7623);
nand U9340 (N_9340,N_7034,N_6367);
or U9341 (N_9341,N_7518,N_6965);
nor U9342 (N_9342,N_6030,N_7016);
nor U9343 (N_9343,N_7121,N_7011);
nor U9344 (N_9344,N_6836,N_6023);
and U9345 (N_9345,N_6049,N_7743);
or U9346 (N_9346,N_7969,N_6430);
nand U9347 (N_9347,N_6561,N_7171);
and U9348 (N_9348,N_6647,N_7740);
and U9349 (N_9349,N_6259,N_6838);
nor U9350 (N_9350,N_6579,N_6984);
and U9351 (N_9351,N_6741,N_7905);
or U9352 (N_9352,N_6649,N_7106);
nand U9353 (N_9353,N_6568,N_6731);
nor U9354 (N_9354,N_7753,N_7144);
nor U9355 (N_9355,N_7591,N_6654);
or U9356 (N_9356,N_7498,N_6060);
nand U9357 (N_9357,N_7139,N_6850);
nor U9358 (N_9358,N_7370,N_6040);
nand U9359 (N_9359,N_7622,N_7632);
and U9360 (N_9360,N_7932,N_6542);
and U9361 (N_9361,N_7009,N_7079);
nor U9362 (N_9362,N_7425,N_7648);
and U9363 (N_9363,N_7007,N_7708);
and U9364 (N_9364,N_7846,N_6658);
nand U9365 (N_9365,N_7237,N_7970);
nand U9366 (N_9366,N_6209,N_7349);
and U9367 (N_9367,N_7142,N_7483);
nand U9368 (N_9368,N_6722,N_6142);
nor U9369 (N_9369,N_6360,N_6216);
and U9370 (N_9370,N_6170,N_7492);
nor U9371 (N_9371,N_6872,N_7431);
nor U9372 (N_9372,N_6598,N_6149);
nand U9373 (N_9373,N_7378,N_6753);
nor U9374 (N_9374,N_7392,N_7405);
or U9375 (N_9375,N_6311,N_7777);
and U9376 (N_9376,N_6228,N_6616);
nand U9377 (N_9377,N_7319,N_7007);
or U9378 (N_9378,N_6793,N_6576);
or U9379 (N_9379,N_6066,N_7024);
and U9380 (N_9380,N_6644,N_6512);
and U9381 (N_9381,N_6542,N_7726);
and U9382 (N_9382,N_6880,N_6454);
nor U9383 (N_9383,N_7810,N_6130);
or U9384 (N_9384,N_7965,N_7803);
and U9385 (N_9385,N_7995,N_7663);
nor U9386 (N_9386,N_7372,N_6684);
or U9387 (N_9387,N_7022,N_7249);
nor U9388 (N_9388,N_7737,N_6943);
and U9389 (N_9389,N_7896,N_7421);
and U9390 (N_9390,N_7223,N_6959);
nand U9391 (N_9391,N_7794,N_7149);
nand U9392 (N_9392,N_7516,N_7633);
nand U9393 (N_9393,N_6858,N_7579);
and U9394 (N_9394,N_7403,N_6510);
and U9395 (N_9395,N_7767,N_6997);
or U9396 (N_9396,N_7015,N_7064);
or U9397 (N_9397,N_7466,N_7352);
nor U9398 (N_9398,N_7652,N_7534);
and U9399 (N_9399,N_7992,N_7590);
nor U9400 (N_9400,N_6717,N_7488);
nor U9401 (N_9401,N_7413,N_6582);
and U9402 (N_9402,N_7594,N_6918);
or U9403 (N_9403,N_7364,N_6960);
or U9404 (N_9404,N_7241,N_6242);
nor U9405 (N_9405,N_6455,N_6067);
or U9406 (N_9406,N_7097,N_7461);
and U9407 (N_9407,N_7034,N_6500);
nand U9408 (N_9408,N_6651,N_6946);
nand U9409 (N_9409,N_7901,N_6427);
and U9410 (N_9410,N_7417,N_7007);
and U9411 (N_9411,N_7674,N_6972);
or U9412 (N_9412,N_6429,N_6524);
or U9413 (N_9413,N_7694,N_6416);
nand U9414 (N_9414,N_7209,N_6930);
nor U9415 (N_9415,N_7523,N_7468);
and U9416 (N_9416,N_6470,N_7470);
and U9417 (N_9417,N_7623,N_7912);
nor U9418 (N_9418,N_7531,N_6937);
nor U9419 (N_9419,N_7786,N_7810);
nand U9420 (N_9420,N_6020,N_7714);
and U9421 (N_9421,N_6658,N_6300);
nor U9422 (N_9422,N_6784,N_6775);
nand U9423 (N_9423,N_7208,N_7741);
nor U9424 (N_9424,N_6196,N_6270);
nand U9425 (N_9425,N_7667,N_6642);
nor U9426 (N_9426,N_7349,N_6127);
nand U9427 (N_9427,N_6819,N_7545);
nor U9428 (N_9428,N_6914,N_7237);
and U9429 (N_9429,N_6447,N_7214);
and U9430 (N_9430,N_6333,N_6403);
nor U9431 (N_9431,N_7707,N_6005);
nor U9432 (N_9432,N_6417,N_7019);
nor U9433 (N_9433,N_7295,N_7347);
nor U9434 (N_9434,N_6145,N_7306);
and U9435 (N_9435,N_6768,N_6823);
nor U9436 (N_9436,N_7340,N_7834);
or U9437 (N_9437,N_7795,N_7855);
or U9438 (N_9438,N_7525,N_6235);
and U9439 (N_9439,N_7021,N_7253);
or U9440 (N_9440,N_6933,N_6617);
nor U9441 (N_9441,N_7316,N_7955);
and U9442 (N_9442,N_7119,N_7785);
and U9443 (N_9443,N_7712,N_7874);
and U9444 (N_9444,N_6483,N_6997);
nor U9445 (N_9445,N_6898,N_7438);
nor U9446 (N_9446,N_6041,N_7924);
and U9447 (N_9447,N_6042,N_7490);
nor U9448 (N_9448,N_6314,N_6245);
nand U9449 (N_9449,N_7938,N_6922);
nor U9450 (N_9450,N_6002,N_6970);
and U9451 (N_9451,N_6448,N_7396);
nor U9452 (N_9452,N_7195,N_6974);
nor U9453 (N_9453,N_6327,N_7385);
or U9454 (N_9454,N_7688,N_6685);
nor U9455 (N_9455,N_7804,N_6212);
and U9456 (N_9456,N_7736,N_6696);
nor U9457 (N_9457,N_6941,N_7732);
nand U9458 (N_9458,N_7419,N_7689);
or U9459 (N_9459,N_7649,N_6588);
xor U9460 (N_9460,N_6289,N_6876);
or U9461 (N_9461,N_6704,N_6497);
or U9462 (N_9462,N_6860,N_7759);
nand U9463 (N_9463,N_7623,N_7586);
nand U9464 (N_9464,N_6659,N_6858);
nor U9465 (N_9465,N_6711,N_7165);
or U9466 (N_9466,N_7315,N_7915);
and U9467 (N_9467,N_7290,N_7305);
or U9468 (N_9468,N_6618,N_6493);
nor U9469 (N_9469,N_6141,N_7296);
nor U9470 (N_9470,N_6124,N_7082);
and U9471 (N_9471,N_7801,N_7424);
xor U9472 (N_9472,N_7608,N_7532);
or U9473 (N_9473,N_7996,N_6735);
and U9474 (N_9474,N_7044,N_7791);
nor U9475 (N_9475,N_7116,N_6307);
and U9476 (N_9476,N_7387,N_7534);
nor U9477 (N_9477,N_6694,N_6309);
nor U9478 (N_9478,N_6306,N_6790);
or U9479 (N_9479,N_6249,N_7285);
xor U9480 (N_9480,N_6369,N_7579);
or U9481 (N_9481,N_7893,N_7987);
nor U9482 (N_9482,N_6802,N_7591);
nand U9483 (N_9483,N_7432,N_7046);
and U9484 (N_9484,N_7795,N_7680);
or U9485 (N_9485,N_7672,N_7681);
nand U9486 (N_9486,N_7804,N_6916);
and U9487 (N_9487,N_7274,N_7300);
and U9488 (N_9488,N_7188,N_7417);
nor U9489 (N_9489,N_7582,N_7004);
and U9490 (N_9490,N_7648,N_7845);
nor U9491 (N_9491,N_7357,N_7568);
or U9492 (N_9492,N_6963,N_6873);
or U9493 (N_9493,N_7500,N_7315);
or U9494 (N_9494,N_7028,N_7320);
nor U9495 (N_9495,N_7333,N_7860);
nor U9496 (N_9496,N_6991,N_7750);
and U9497 (N_9497,N_6003,N_6116);
nor U9498 (N_9498,N_7266,N_6163);
nor U9499 (N_9499,N_6241,N_6608);
or U9500 (N_9500,N_7059,N_7571);
nor U9501 (N_9501,N_6101,N_6213);
nor U9502 (N_9502,N_7477,N_7268);
or U9503 (N_9503,N_7118,N_6658);
and U9504 (N_9504,N_6957,N_7777);
nand U9505 (N_9505,N_7368,N_6771);
and U9506 (N_9506,N_7530,N_7761);
or U9507 (N_9507,N_6593,N_6319);
nor U9508 (N_9508,N_7950,N_7317);
nand U9509 (N_9509,N_6334,N_7656);
or U9510 (N_9510,N_6711,N_6077);
and U9511 (N_9511,N_6562,N_6406);
or U9512 (N_9512,N_6333,N_7050);
or U9513 (N_9513,N_7063,N_6125);
nor U9514 (N_9514,N_6146,N_7508);
nor U9515 (N_9515,N_7859,N_6372);
or U9516 (N_9516,N_6245,N_7653);
or U9517 (N_9517,N_6956,N_6663);
and U9518 (N_9518,N_7356,N_6332);
nand U9519 (N_9519,N_6145,N_6889);
nand U9520 (N_9520,N_6763,N_7817);
or U9521 (N_9521,N_6867,N_6440);
nand U9522 (N_9522,N_6155,N_6761);
nor U9523 (N_9523,N_6227,N_6622);
nor U9524 (N_9524,N_6496,N_6325);
nand U9525 (N_9525,N_7928,N_7882);
or U9526 (N_9526,N_7780,N_7409);
nor U9527 (N_9527,N_7458,N_7637);
and U9528 (N_9528,N_6309,N_6822);
nand U9529 (N_9529,N_7560,N_6595);
and U9530 (N_9530,N_6766,N_7496);
nor U9531 (N_9531,N_6721,N_7586);
nor U9532 (N_9532,N_6531,N_7954);
nand U9533 (N_9533,N_6956,N_7919);
nor U9534 (N_9534,N_7234,N_6940);
nand U9535 (N_9535,N_7924,N_6595);
nor U9536 (N_9536,N_7022,N_7963);
nor U9537 (N_9537,N_6833,N_7441);
or U9538 (N_9538,N_6878,N_6661);
or U9539 (N_9539,N_7395,N_7501);
or U9540 (N_9540,N_6626,N_7783);
or U9541 (N_9541,N_7370,N_6620);
nor U9542 (N_9542,N_6882,N_6722);
nor U9543 (N_9543,N_6684,N_6375);
or U9544 (N_9544,N_7200,N_6762);
or U9545 (N_9545,N_7212,N_6853);
nand U9546 (N_9546,N_7312,N_7158);
and U9547 (N_9547,N_7139,N_7199);
nand U9548 (N_9548,N_7097,N_7564);
nor U9549 (N_9549,N_6103,N_7053);
or U9550 (N_9550,N_7435,N_7672);
nand U9551 (N_9551,N_7671,N_7887);
nor U9552 (N_9552,N_6896,N_6658);
and U9553 (N_9553,N_6392,N_6058);
or U9554 (N_9554,N_6139,N_6392);
nand U9555 (N_9555,N_6245,N_6281);
and U9556 (N_9556,N_7474,N_6260);
nand U9557 (N_9557,N_6999,N_7355);
nor U9558 (N_9558,N_7099,N_7538);
or U9559 (N_9559,N_7414,N_6761);
nand U9560 (N_9560,N_6409,N_6642);
and U9561 (N_9561,N_7064,N_6144);
or U9562 (N_9562,N_7522,N_6711);
nor U9563 (N_9563,N_7220,N_6924);
and U9564 (N_9564,N_6396,N_7743);
and U9565 (N_9565,N_6324,N_6209);
or U9566 (N_9566,N_6295,N_6195);
or U9567 (N_9567,N_6698,N_6263);
or U9568 (N_9568,N_6202,N_6606);
nand U9569 (N_9569,N_6274,N_6299);
nor U9570 (N_9570,N_7153,N_6618);
and U9571 (N_9571,N_7286,N_6624);
and U9572 (N_9572,N_6510,N_6875);
and U9573 (N_9573,N_6969,N_7777);
or U9574 (N_9574,N_6599,N_7317);
or U9575 (N_9575,N_6848,N_7203);
nand U9576 (N_9576,N_6470,N_7176);
and U9577 (N_9577,N_7679,N_7869);
or U9578 (N_9578,N_7112,N_7715);
and U9579 (N_9579,N_7667,N_7559);
nand U9580 (N_9580,N_7774,N_6172);
nand U9581 (N_9581,N_7658,N_6691);
nor U9582 (N_9582,N_6632,N_7013);
nor U9583 (N_9583,N_6708,N_6181);
nor U9584 (N_9584,N_7766,N_7040);
nand U9585 (N_9585,N_7660,N_7165);
nor U9586 (N_9586,N_6971,N_6700);
or U9587 (N_9587,N_6953,N_6202);
xor U9588 (N_9588,N_6548,N_6987);
nand U9589 (N_9589,N_7762,N_6461);
or U9590 (N_9590,N_7091,N_7905);
nor U9591 (N_9591,N_6953,N_6948);
and U9592 (N_9592,N_6896,N_7389);
nor U9593 (N_9593,N_6445,N_7712);
nor U9594 (N_9594,N_6022,N_7093);
and U9595 (N_9595,N_7925,N_7819);
nand U9596 (N_9596,N_6268,N_7703);
or U9597 (N_9597,N_6402,N_7949);
and U9598 (N_9598,N_7996,N_7980);
or U9599 (N_9599,N_7385,N_6744);
or U9600 (N_9600,N_7503,N_6779);
nor U9601 (N_9601,N_7697,N_6641);
nor U9602 (N_9602,N_7083,N_7572);
nor U9603 (N_9603,N_7287,N_7862);
nand U9604 (N_9604,N_7561,N_6080);
and U9605 (N_9605,N_6184,N_6929);
nor U9606 (N_9606,N_7616,N_7357);
nor U9607 (N_9607,N_7079,N_7810);
or U9608 (N_9608,N_7384,N_7444);
and U9609 (N_9609,N_7809,N_7211);
or U9610 (N_9610,N_7451,N_7576);
or U9611 (N_9611,N_7805,N_7215);
nand U9612 (N_9612,N_7242,N_6015);
or U9613 (N_9613,N_6269,N_7962);
nor U9614 (N_9614,N_6558,N_7540);
and U9615 (N_9615,N_6221,N_6668);
or U9616 (N_9616,N_7228,N_6072);
or U9617 (N_9617,N_7712,N_7872);
xor U9618 (N_9618,N_7939,N_7518);
xor U9619 (N_9619,N_7000,N_6826);
nor U9620 (N_9620,N_7178,N_7978);
nand U9621 (N_9621,N_6924,N_7727);
nand U9622 (N_9622,N_7213,N_6980);
and U9623 (N_9623,N_6192,N_7722);
or U9624 (N_9624,N_7662,N_7420);
and U9625 (N_9625,N_7548,N_7812);
or U9626 (N_9626,N_7658,N_6219);
nor U9627 (N_9627,N_6757,N_7140);
and U9628 (N_9628,N_6520,N_7841);
and U9629 (N_9629,N_7541,N_7424);
or U9630 (N_9630,N_7626,N_7416);
nor U9631 (N_9631,N_6131,N_7343);
nor U9632 (N_9632,N_6243,N_7482);
and U9633 (N_9633,N_7123,N_6045);
nand U9634 (N_9634,N_7921,N_7196);
nor U9635 (N_9635,N_6285,N_6072);
and U9636 (N_9636,N_6737,N_7763);
and U9637 (N_9637,N_6615,N_7373);
or U9638 (N_9638,N_6739,N_6660);
nor U9639 (N_9639,N_7656,N_6066);
or U9640 (N_9640,N_7873,N_6972);
and U9641 (N_9641,N_6740,N_6086);
nor U9642 (N_9642,N_7656,N_6584);
nand U9643 (N_9643,N_6028,N_6269);
or U9644 (N_9644,N_7273,N_6744);
and U9645 (N_9645,N_6218,N_7422);
nor U9646 (N_9646,N_6687,N_6337);
nand U9647 (N_9647,N_6549,N_7633);
and U9648 (N_9648,N_7655,N_7250);
nor U9649 (N_9649,N_7476,N_7992);
or U9650 (N_9650,N_7614,N_6849);
and U9651 (N_9651,N_7241,N_7083);
nand U9652 (N_9652,N_7045,N_6830);
nor U9653 (N_9653,N_6006,N_7549);
nor U9654 (N_9654,N_7018,N_7425);
or U9655 (N_9655,N_6482,N_7310);
nand U9656 (N_9656,N_6214,N_7325);
nor U9657 (N_9657,N_7842,N_7158);
nor U9658 (N_9658,N_6428,N_6663);
or U9659 (N_9659,N_6557,N_7355);
and U9660 (N_9660,N_7955,N_7852);
nor U9661 (N_9661,N_6497,N_7893);
or U9662 (N_9662,N_7027,N_6872);
and U9663 (N_9663,N_7156,N_6691);
or U9664 (N_9664,N_6681,N_6078);
and U9665 (N_9665,N_7146,N_6086);
or U9666 (N_9666,N_6427,N_6018);
nor U9667 (N_9667,N_6556,N_7453);
nor U9668 (N_9668,N_7471,N_6225);
or U9669 (N_9669,N_7854,N_7128);
and U9670 (N_9670,N_7550,N_7052);
nor U9671 (N_9671,N_6017,N_6900);
or U9672 (N_9672,N_6631,N_6849);
nor U9673 (N_9673,N_6768,N_7192);
nand U9674 (N_9674,N_7963,N_6021);
and U9675 (N_9675,N_6374,N_7847);
or U9676 (N_9676,N_6565,N_7128);
and U9677 (N_9677,N_6923,N_6689);
nand U9678 (N_9678,N_6508,N_6418);
and U9679 (N_9679,N_6676,N_7631);
and U9680 (N_9680,N_7437,N_6941);
nor U9681 (N_9681,N_7256,N_6744);
or U9682 (N_9682,N_7328,N_7962);
nor U9683 (N_9683,N_7418,N_6095);
or U9684 (N_9684,N_7186,N_6169);
or U9685 (N_9685,N_6490,N_6021);
or U9686 (N_9686,N_7816,N_6795);
nor U9687 (N_9687,N_7222,N_7233);
nor U9688 (N_9688,N_6939,N_7572);
nand U9689 (N_9689,N_6454,N_7277);
and U9690 (N_9690,N_6355,N_6946);
nor U9691 (N_9691,N_6444,N_6425);
nand U9692 (N_9692,N_6995,N_7551);
and U9693 (N_9693,N_7873,N_7121);
or U9694 (N_9694,N_7980,N_6730);
nand U9695 (N_9695,N_7711,N_7391);
or U9696 (N_9696,N_7136,N_6726);
nor U9697 (N_9697,N_6738,N_6931);
nand U9698 (N_9698,N_7441,N_7775);
and U9699 (N_9699,N_6270,N_7264);
or U9700 (N_9700,N_6734,N_7601);
nor U9701 (N_9701,N_6636,N_6916);
and U9702 (N_9702,N_7683,N_6691);
xnor U9703 (N_9703,N_6089,N_6020);
nand U9704 (N_9704,N_7497,N_7459);
nor U9705 (N_9705,N_6880,N_6644);
nand U9706 (N_9706,N_7174,N_6414);
and U9707 (N_9707,N_7861,N_7724);
and U9708 (N_9708,N_6910,N_7859);
nor U9709 (N_9709,N_6176,N_7798);
or U9710 (N_9710,N_7210,N_7065);
and U9711 (N_9711,N_7949,N_6258);
or U9712 (N_9712,N_7482,N_6047);
nor U9713 (N_9713,N_6504,N_7409);
and U9714 (N_9714,N_6913,N_6924);
nor U9715 (N_9715,N_7839,N_7228);
nand U9716 (N_9716,N_6508,N_7781);
nand U9717 (N_9717,N_6117,N_7592);
nor U9718 (N_9718,N_6389,N_6537);
nand U9719 (N_9719,N_6025,N_6269);
nand U9720 (N_9720,N_7970,N_7418);
or U9721 (N_9721,N_6313,N_6488);
or U9722 (N_9722,N_6321,N_7511);
and U9723 (N_9723,N_6252,N_7406);
or U9724 (N_9724,N_7598,N_7078);
and U9725 (N_9725,N_7850,N_7778);
nor U9726 (N_9726,N_6112,N_7534);
or U9727 (N_9727,N_6978,N_6485);
nand U9728 (N_9728,N_6240,N_6472);
or U9729 (N_9729,N_6385,N_7375);
nor U9730 (N_9730,N_7454,N_7662);
nand U9731 (N_9731,N_7004,N_7620);
nor U9732 (N_9732,N_6282,N_7734);
nor U9733 (N_9733,N_6541,N_7526);
nor U9734 (N_9734,N_7721,N_7223);
nor U9735 (N_9735,N_7676,N_7198);
and U9736 (N_9736,N_6103,N_7954);
and U9737 (N_9737,N_6771,N_6767);
nand U9738 (N_9738,N_7037,N_6200);
and U9739 (N_9739,N_7172,N_6370);
and U9740 (N_9740,N_7583,N_7137);
or U9741 (N_9741,N_7343,N_6415);
nor U9742 (N_9742,N_7159,N_6968);
and U9743 (N_9743,N_7950,N_6291);
and U9744 (N_9744,N_7246,N_7313);
and U9745 (N_9745,N_6348,N_7710);
nand U9746 (N_9746,N_6388,N_6481);
nor U9747 (N_9747,N_6825,N_7863);
or U9748 (N_9748,N_7685,N_7617);
and U9749 (N_9749,N_6558,N_6097);
nor U9750 (N_9750,N_6328,N_6499);
or U9751 (N_9751,N_6918,N_6499);
or U9752 (N_9752,N_6901,N_6346);
and U9753 (N_9753,N_6960,N_7324);
nor U9754 (N_9754,N_6673,N_6192);
and U9755 (N_9755,N_6796,N_7999);
or U9756 (N_9756,N_7010,N_6655);
or U9757 (N_9757,N_6946,N_6283);
or U9758 (N_9758,N_7469,N_7820);
and U9759 (N_9759,N_7003,N_7774);
nand U9760 (N_9760,N_7031,N_6354);
and U9761 (N_9761,N_7679,N_7949);
nand U9762 (N_9762,N_7892,N_7288);
or U9763 (N_9763,N_7475,N_6313);
nand U9764 (N_9764,N_7400,N_6922);
or U9765 (N_9765,N_6445,N_7827);
and U9766 (N_9766,N_7390,N_6163);
and U9767 (N_9767,N_7124,N_6936);
and U9768 (N_9768,N_7584,N_6057);
and U9769 (N_9769,N_7247,N_7900);
nand U9770 (N_9770,N_7158,N_7819);
nor U9771 (N_9771,N_6656,N_7531);
and U9772 (N_9772,N_6123,N_6026);
and U9773 (N_9773,N_6895,N_7431);
or U9774 (N_9774,N_6079,N_7809);
nor U9775 (N_9775,N_7763,N_6001);
nor U9776 (N_9776,N_7493,N_6210);
or U9777 (N_9777,N_6833,N_6988);
nor U9778 (N_9778,N_7926,N_6180);
or U9779 (N_9779,N_6765,N_7914);
nor U9780 (N_9780,N_6640,N_7521);
nor U9781 (N_9781,N_6521,N_6188);
or U9782 (N_9782,N_6419,N_7526);
and U9783 (N_9783,N_7060,N_7394);
nor U9784 (N_9784,N_6947,N_7533);
nor U9785 (N_9785,N_6827,N_7493);
nor U9786 (N_9786,N_6074,N_7846);
or U9787 (N_9787,N_6741,N_6158);
or U9788 (N_9788,N_7106,N_6833);
and U9789 (N_9789,N_6186,N_7950);
or U9790 (N_9790,N_7129,N_7072);
nor U9791 (N_9791,N_7132,N_6510);
nor U9792 (N_9792,N_6068,N_7103);
or U9793 (N_9793,N_6270,N_6426);
nand U9794 (N_9794,N_6752,N_7689);
nor U9795 (N_9795,N_6077,N_6014);
and U9796 (N_9796,N_6191,N_7321);
nor U9797 (N_9797,N_7231,N_6808);
nor U9798 (N_9798,N_6338,N_7450);
or U9799 (N_9799,N_6231,N_7059);
and U9800 (N_9800,N_7507,N_6493);
nor U9801 (N_9801,N_6894,N_7766);
or U9802 (N_9802,N_6398,N_6892);
or U9803 (N_9803,N_7672,N_7168);
nor U9804 (N_9804,N_7903,N_7547);
nand U9805 (N_9805,N_6013,N_6374);
nor U9806 (N_9806,N_7613,N_7358);
or U9807 (N_9807,N_7196,N_7170);
or U9808 (N_9808,N_7638,N_6034);
and U9809 (N_9809,N_7590,N_6569);
and U9810 (N_9810,N_6088,N_6941);
nand U9811 (N_9811,N_6320,N_7396);
and U9812 (N_9812,N_6853,N_6109);
nor U9813 (N_9813,N_7715,N_6994);
or U9814 (N_9814,N_6879,N_6963);
nor U9815 (N_9815,N_7986,N_6615);
nand U9816 (N_9816,N_6630,N_6904);
or U9817 (N_9817,N_6054,N_7147);
and U9818 (N_9818,N_6246,N_7676);
and U9819 (N_9819,N_7484,N_7677);
or U9820 (N_9820,N_6608,N_6627);
and U9821 (N_9821,N_6382,N_7405);
or U9822 (N_9822,N_7611,N_6918);
and U9823 (N_9823,N_6193,N_6611);
nor U9824 (N_9824,N_6784,N_7568);
nand U9825 (N_9825,N_7740,N_7124);
and U9826 (N_9826,N_7499,N_6650);
nand U9827 (N_9827,N_7276,N_7880);
or U9828 (N_9828,N_7474,N_7868);
or U9829 (N_9829,N_6279,N_7911);
nand U9830 (N_9830,N_7702,N_6996);
and U9831 (N_9831,N_7329,N_7871);
nand U9832 (N_9832,N_6488,N_6364);
or U9833 (N_9833,N_7212,N_7756);
nor U9834 (N_9834,N_6580,N_6547);
or U9835 (N_9835,N_6712,N_6691);
nand U9836 (N_9836,N_7218,N_7800);
or U9837 (N_9837,N_6872,N_7491);
nand U9838 (N_9838,N_7435,N_7577);
and U9839 (N_9839,N_6009,N_7362);
nand U9840 (N_9840,N_7564,N_7445);
or U9841 (N_9841,N_6523,N_6586);
nand U9842 (N_9842,N_6184,N_7324);
nor U9843 (N_9843,N_7315,N_6970);
nand U9844 (N_9844,N_6647,N_6618);
and U9845 (N_9845,N_6254,N_7491);
or U9846 (N_9846,N_6222,N_7588);
nor U9847 (N_9847,N_7070,N_7842);
nor U9848 (N_9848,N_7625,N_6403);
or U9849 (N_9849,N_7921,N_7112);
and U9850 (N_9850,N_6053,N_6439);
nor U9851 (N_9851,N_7277,N_6865);
nand U9852 (N_9852,N_6908,N_6227);
nor U9853 (N_9853,N_7660,N_7445);
nand U9854 (N_9854,N_7679,N_6883);
or U9855 (N_9855,N_6237,N_6376);
and U9856 (N_9856,N_6627,N_7284);
nor U9857 (N_9857,N_6602,N_7298);
nor U9858 (N_9858,N_6556,N_6369);
or U9859 (N_9859,N_7356,N_7653);
nand U9860 (N_9860,N_7281,N_6615);
or U9861 (N_9861,N_6919,N_7086);
and U9862 (N_9862,N_7890,N_6386);
or U9863 (N_9863,N_7674,N_6835);
or U9864 (N_9864,N_6780,N_6170);
or U9865 (N_9865,N_6296,N_6859);
or U9866 (N_9866,N_6971,N_7052);
or U9867 (N_9867,N_7216,N_6562);
xor U9868 (N_9868,N_7061,N_6045);
and U9869 (N_9869,N_6786,N_7053);
or U9870 (N_9870,N_6410,N_7286);
nor U9871 (N_9871,N_6500,N_6480);
nand U9872 (N_9872,N_6927,N_7943);
nand U9873 (N_9873,N_6941,N_6731);
and U9874 (N_9874,N_7389,N_7708);
or U9875 (N_9875,N_6021,N_6584);
or U9876 (N_9876,N_7700,N_6968);
xor U9877 (N_9877,N_7509,N_7879);
nand U9878 (N_9878,N_7763,N_7230);
nor U9879 (N_9879,N_6270,N_6525);
nand U9880 (N_9880,N_7011,N_6541);
or U9881 (N_9881,N_6078,N_6052);
and U9882 (N_9882,N_7486,N_7279);
and U9883 (N_9883,N_7043,N_6880);
nor U9884 (N_9884,N_7789,N_7886);
nand U9885 (N_9885,N_6249,N_6572);
or U9886 (N_9886,N_6002,N_7299);
nor U9887 (N_9887,N_7387,N_7193);
and U9888 (N_9888,N_7708,N_6319);
and U9889 (N_9889,N_7600,N_6775);
and U9890 (N_9890,N_7574,N_7678);
nor U9891 (N_9891,N_6336,N_6209);
and U9892 (N_9892,N_7928,N_6817);
nor U9893 (N_9893,N_7119,N_6602);
and U9894 (N_9894,N_6519,N_7551);
and U9895 (N_9895,N_7617,N_7007);
nand U9896 (N_9896,N_6647,N_6512);
nor U9897 (N_9897,N_6570,N_7854);
and U9898 (N_9898,N_6288,N_7553);
nor U9899 (N_9899,N_6756,N_7757);
nand U9900 (N_9900,N_7701,N_6746);
nand U9901 (N_9901,N_6079,N_6174);
nand U9902 (N_9902,N_6257,N_7392);
and U9903 (N_9903,N_6665,N_6622);
and U9904 (N_9904,N_7852,N_6390);
nor U9905 (N_9905,N_7068,N_7087);
nand U9906 (N_9906,N_6517,N_7685);
or U9907 (N_9907,N_6702,N_6057);
nand U9908 (N_9908,N_6507,N_7431);
nor U9909 (N_9909,N_7188,N_6890);
xnor U9910 (N_9910,N_6989,N_7807);
nor U9911 (N_9911,N_6116,N_6315);
or U9912 (N_9912,N_6355,N_6465);
nor U9913 (N_9913,N_7598,N_6707);
and U9914 (N_9914,N_6030,N_7416);
and U9915 (N_9915,N_7834,N_7062);
and U9916 (N_9916,N_6349,N_6444);
or U9917 (N_9917,N_6782,N_7590);
and U9918 (N_9918,N_6685,N_7080);
or U9919 (N_9919,N_6764,N_6632);
or U9920 (N_9920,N_7259,N_7629);
nor U9921 (N_9921,N_7972,N_6405);
nor U9922 (N_9922,N_6987,N_7274);
nand U9923 (N_9923,N_6051,N_7721);
nor U9924 (N_9924,N_6931,N_7468);
nor U9925 (N_9925,N_7472,N_6037);
or U9926 (N_9926,N_7680,N_7261);
xnor U9927 (N_9927,N_6826,N_7400);
nand U9928 (N_9928,N_6307,N_6118);
nor U9929 (N_9929,N_6416,N_7241);
nor U9930 (N_9930,N_6747,N_7417);
nand U9931 (N_9931,N_7904,N_7874);
or U9932 (N_9932,N_7406,N_6066);
nor U9933 (N_9933,N_7065,N_6896);
nand U9934 (N_9934,N_7711,N_7118);
nor U9935 (N_9935,N_7467,N_7056);
and U9936 (N_9936,N_7795,N_7796);
or U9937 (N_9937,N_7031,N_7473);
or U9938 (N_9938,N_7693,N_6565);
and U9939 (N_9939,N_7309,N_7961);
nand U9940 (N_9940,N_6379,N_7917);
and U9941 (N_9941,N_6231,N_6400);
or U9942 (N_9942,N_7882,N_7242);
or U9943 (N_9943,N_7639,N_7631);
nor U9944 (N_9944,N_7500,N_7750);
nand U9945 (N_9945,N_7609,N_6551);
nand U9946 (N_9946,N_6999,N_7621);
or U9947 (N_9947,N_6482,N_6955);
and U9948 (N_9948,N_6155,N_7254);
or U9949 (N_9949,N_7182,N_6905);
nand U9950 (N_9950,N_6831,N_7995);
nor U9951 (N_9951,N_7541,N_6843);
nand U9952 (N_9952,N_7842,N_7836);
or U9953 (N_9953,N_7301,N_6774);
nor U9954 (N_9954,N_6372,N_7050);
nand U9955 (N_9955,N_6831,N_6629);
or U9956 (N_9956,N_6583,N_6834);
nor U9957 (N_9957,N_7274,N_6198);
and U9958 (N_9958,N_7196,N_7002);
nand U9959 (N_9959,N_7457,N_7196);
nand U9960 (N_9960,N_7235,N_6508);
and U9961 (N_9961,N_7958,N_6020);
or U9962 (N_9962,N_6975,N_6194);
and U9963 (N_9963,N_6241,N_7983);
and U9964 (N_9964,N_7130,N_7150);
and U9965 (N_9965,N_6787,N_6710);
nor U9966 (N_9966,N_7832,N_7979);
nor U9967 (N_9967,N_6550,N_6168);
or U9968 (N_9968,N_7386,N_6061);
and U9969 (N_9969,N_6572,N_7861);
nand U9970 (N_9970,N_7118,N_7082);
nor U9971 (N_9971,N_6601,N_6376);
or U9972 (N_9972,N_6649,N_7159);
nand U9973 (N_9973,N_6702,N_6637);
nor U9974 (N_9974,N_7101,N_7241);
and U9975 (N_9975,N_7119,N_6144);
and U9976 (N_9976,N_6461,N_7674);
or U9977 (N_9977,N_7222,N_7653);
nor U9978 (N_9978,N_7856,N_6815);
nor U9979 (N_9979,N_6376,N_7666);
nor U9980 (N_9980,N_7154,N_7100);
or U9981 (N_9981,N_6851,N_7235);
and U9982 (N_9982,N_7495,N_6520);
nor U9983 (N_9983,N_7514,N_7923);
nand U9984 (N_9984,N_6888,N_7726);
or U9985 (N_9985,N_6494,N_7931);
or U9986 (N_9986,N_6397,N_7237);
nand U9987 (N_9987,N_6285,N_7587);
and U9988 (N_9988,N_6589,N_6367);
nand U9989 (N_9989,N_7860,N_7709);
nor U9990 (N_9990,N_6172,N_7757);
or U9991 (N_9991,N_7472,N_7760);
nand U9992 (N_9992,N_6023,N_7175);
nand U9993 (N_9993,N_6556,N_6462);
nor U9994 (N_9994,N_7051,N_7803);
and U9995 (N_9995,N_7478,N_6429);
or U9996 (N_9996,N_6808,N_7813);
nor U9997 (N_9997,N_7837,N_6080);
or U9998 (N_9998,N_7072,N_6527);
nand U9999 (N_9999,N_7215,N_7691);
nand UO_0 (O_0,N_9361,N_9154);
or UO_1 (O_1,N_8466,N_8587);
nor UO_2 (O_2,N_8120,N_8874);
nor UO_3 (O_3,N_9371,N_9937);
or UO_4 (O_4,N_8658,N_8056);
or UO_5 (O_5,N_9811,N_9313);
nand UO_6 (O_6,N_9933,N_9574);
and UO_7 (O_7,N_8212,N_9172);
nand UO_8 (O_8,N_9387,N_8049);
and UO_9 (O_9,N_9695,N_9722);
or UO_10 (O_10,N_8945,N_9943);
nand UO_11 (O_11,N_9061,N_9660);
or UO_12 (O_12,N_8485,N_8821);
nand UO_13 (O_13,N_9346,N_9806);
xor UO_14 (O_14,N_8743,N_8002);
and UO_15 (O_15,N_9985,N_9597);
nand UO_16 (O_16,N_9487,N_9883);
xor UO_17 (O_17,N_9393,N_8293);
xnor UO_18 (O_18,N_8184,N_9657);
and UO_19 (O_19,N_9714,N_8629);
or UO_20 (O_20,N_9339,N_8584);
nand UO_21 (O_21,N_8304,N_9939);
or UO_22 (O_22,N_9818,N_8104);
nor UO_23 (O_23,N_8324,N_8146);
nand UO_24 (O_24,N_9631,N_8240);
nor UO_25 (O_25,N_9262,N_8286);
and UO_26 (O_26,N_9424,N_9456);
nor UO_27 (O_27,N_8110,N_8676);
nor UO_28 (O_28,N_9591,N_9754);
or UO_29 (O_29,N_8913,N_8115);
nand UO_30 (O_30,N_9435,N_9412);
and UO_31 (O_31,N_8158,N_9664);
or UO_32 (O_32,N_9954,N_9064);
xor UO_33 (O_33,N_9453,N_9922);
nor UO_34 (O_34,N_8238,N_9469);
nor UO_35 (O_35,N_9282,N_8458);
nand UO_36 (O_36,N_8457,N_9108);
or UO_37 (O_37,N_8926,N_9237);
nand UO_38 (O_38,N_9963,N_9659);
nand UO_39 (O_39,N_9827,N_9202);
and UO_40 (O_40,N_8174,N_8768);
and UO_41 (O_41,N_9198,N_9117);
or UO_42 (O_42,N_8614,N_8948);
nand UO_43 (O_43,N_8160,N_8532);
nand UO_44 (O_44,N_8495,N_8034);
nor UO_45 (O_45,N_9782,N_9715);
and UO_46 (O_46,N_8953,N_9304);
nor UO_47 (O_47,N_8771,N_8252);
and UO_48 (O_48,N_8351,N_9529);
or UO_49 (O_49,N_9952,N_8917);
and UO_50 (O_50,N_8352,N_8535);
or UO_51 (O_51,N_8521,N_9175);
and UO_52 (O_52,N_9966,N_9372);
nand UO_53 (O_53,N_8029,N_9964);
or UO_54 (O_54,N_8605,N_8973);
nand UO_55 (O_55,N_9614,N_8717);
or UO_56 (O_56,N_9792,N_9155);
nand UO_57 (O_57,N_9316,N_9137);
nor UO_58 (O_58,N_9377,N_8003);
nand UO_59 (O_59,N_8026,N_9809);
and UO_60 (O_60,N_8607,N_9897);
and UO_61 (O_61,N_9600,N_9975);
nand UO_62 (O_62,N_9936,N_9105);
or UO_63 (O_63,N_8401,N_9348);
and UO_64 (O_64,N_9696,N_9192);
or UO_65 (O_65,N_8559,N_9189);
or UO_66 (O_66,N_8877,N_9912);
nor UO_67 (O_67,N_9463,N_9395);
nand UO_68 (O_68,N_9716,N_8523);
and UO_69 (O_69,N_9701,N_8085);
nor UO_70 (O_70,N_9708,N_8490);
or UO_71 (O_71,N_8190,N_8317);
or UO_72 (O_72,N_8407,N_9088);
nand UO_73 (O_73,N_9434,N_9812);
and UO_74 (O_74,N_8388,N_9533);
and UO_75 (O_75,N_8140,N_9725);
nand UO_76 (O_76,N_9541,N_8161);
nand UO_77 (O_77,N_9444,N_8939);
or UO_78 (O_78,N_9068,N_9586);
nor UO_79 (O_79,N_9635,N_8928);
and UO_80 (O_80,N_8599,N_9143);
nand UO_81 (O_81,N_8764,N_8534);
or UO_82 (O_82,N_8012,N_8342);
nor UO_83 (O_83,N_8338,N_9568);
nor UO_84 (O_84,N_8994,N_8969);
nand UO_85 (O_85,N_9563,N_9113);
or UO_86 (O_86,N_9133,N_9232);
and UO_87 (O_87,N_9284,N_9881);
or UO_88 (O_88,N_8492,N_9810);
nand UO_89 (O_89,N_8859,N_8399);
nand UO_90 (O_90,N_9641,N_8009);
and UO_91 (O_91,N_9446,N_9616);
nor UO_92 (O_92,N_9879,N_9106);
or UO_93 (O_93,N_9242,N_9526);
and UO_94 (O_94,N_8751,N_8738);
nor UO_95 (O_95,N_8947,N_8270);
nor UO_96 (O_96,N_8977,N_8498);
or UO_97 (O_97,N_8779,N_9023);
and UO_98 (O_98,N_8542,N_8047);
and UO_99 (O_99,N_9235,N_9638);
or UO_100 (O_100,N_9968,N_9392);
nand UO_101 (O_101,N_9458,N_9190);
nor UO_102 (O_102,N_8289,N_8512);
nor UO_103 (O_103,N_8669,N_8907);
nor UO_104 (O_104,N_9479,N_9314);
or UO_105 (O_105,N_8220,N_8133);
nor UO_106 (O_106,N_8387,N_9405);
nand UO_107 (O_107,N_8437,N_8856);
nand UO_108 (O_108,N_9542,N_8265);
nor UO_109 (O_109,N_9762,N_8530);
or UO_110 (O_110,N_9970,N_9658);
or UO_111 (O_111,N_8068,N_9678);
and UO_112 (O_112,N_9560,N_9514);
nand UO_113 (O_113,N_8912,N_9000);
or UO_114 (O_114,N_8185,N_9025);
nand UO_115 (O_115,N_9866,N_8311);
nand UO_116 (O_116,N_9868,N_8908);
nand UO_117 (O_117,N_9502,N_9864);
nor UO_118 (O_118,N_9276,N_8063);
or UO_119 (O_119,N_9732,N_9623);
nor UO_120 (O_120,N_9473,N_8233);
or UO_121 (O_121,N_9146,N_9665);
xnor UO_122 (O_122,N_8232,N_9071);
nor UO_123 (O_123,N_8765,N_9628);
nor UO_124 (O_124,N_8054,N_9019);
nor UO_125 (O_125,N_9005,N_8130);
nand UO_126 (O_126,N_9383,N_9612);
nor UO_127 (O_127,N_8577,N_9196);
nand UO_128 (O_128,N_9437,N_9800);
or UO_129 (O_129,N_8038,N_8013);
or UO_130 (O_130,N_9858,N_9850);
nand UO_131 (O_131,N_8702,N_9540);
and UO_132 (O_132,N_8671,N_9150);
nand UO_133 (O_133,N_8760,N_9863);
and UO_134 (O_134,N_9211,N_9278);
nand UO_135 (O_135,N_9849,N_8114);
and UO_136 (O_136,N_8483,N_9305);
nor UO_137 (O_137,N_8596,N_8478);
and UO_138 (O_138,N_9666,N_9281);
nand UO_139 (O_139,N_8739,N_8718);
and UO_140 (O_140,N_9279,N_8082);
and UO_141 (O_141,N_9587,N_8119);
nor UO_142 (O_142,N_8960,N_8021);
nor UO_143 (O_143,N_8354,N_8621);
nand UO_144 (O_144,N_8789,N_9303);
nand UO_145 (O_145,N_8173,N_8080);
and UO_146 (O_146,N_8419,N_9216);
nand UO_147 (O_147,N_9918,N_9698);
nor UO_148 (O_148,N_9451,N_8198);
nor UO_149 (O_149,N_9249,N_8213);
nor UO_150 (O_150,N_8242,N_9063);
nand UO_151 (O_151,N_8321,N_9488);
nand UO_152 (O_152,N_9772,N_9191);
nand UO_153 (O_153,N_9325,N_8582);
and UO_154 (O_154,N_8776,N_9608);
nor UO_155 (O_155,N_9517,N_8566);
or UO_156 (O_156,N_9798,N_9466);
or UO_157 (O_157,N_8844,N_9275);
nand UO_158 (O_158,N_9752,N_8862);
or UO_159 (O_159,N_8217,N_9687);
nor UO_160 (O_160,N_9839,N_9861);
nor UO_161 (O_161,N_9930,N_9788);
nor UO_162 (O_162,N_8602,N_8520);
or UO_163 (O_163,N_9072,N_8744);
nor UO_164 (O_164,N_8793,N_9915);
nor UO_165 (O_165,N_9256,N_8235);
and UO_166 (O_166,N_9416,N_9382);
or UO_167 (O_167,N_9241,N_8272);
or UO_168 (O_168,N_9343,N_9536);
nor UO_169 (O_169,N_9047,N_9477);
and UO_170 (O_170,N_8803,N_8134);
or UO_171 (O_171,N_8590,N_9627);
or UO_172 (O_172,N_8097,N_9822);
nor UO_173 (O_173,N_8667,N_8550);
nand UO_174 (O_174,N_8285,N_8755);
nor UO_175 (O_175,N_8288,N_8326);
and UO_176 (O_176,N_9156,N_9662);
xnor UO_177 (O_177,N_8378,N_8347);
and UO_178 (O_178,N_9904,N_9669);
and UO_179 (O_179,N_8567,N_8456);
and UO_180 (O_180,N_8269,N_9356);
and UO_181 (O_181,N_8522,N_9969);
nand UO_182 (O_182,N_9765,N_9259);
nor UO_183 (O_183,N_9229,N_8704);
nand UO_184 (O_184,N_9595,N_9652);
nor UO_185 (O_185,N_8098,N_9130);
nand UO_186 (O_186,N_9280,N_9365);
nor UO_187 (O_187,N_8811,N_9821);
and UO_188 (O_188,N_8052,N_9869);
or UO_189 (O_189,N_8886,N_8872);
nor UO_190 (O_190,N_9097,N_9751);
or UO_191 (O_191,N_9168,N_9848);
or UO_192 (O_192,N_9690,N_9615);
or UO_193 (O_193,N_9508,N_8984);
and UO_194 (O_194,N_8782,N_9317);
or UO_195 (O_195,N_9749,N_9796);
and UO_196 (O_196,N_8683,N_8979);
or UO_197 (O_197,N_9484,N_9777);
and UO_198 (O_198,N_9993,N_9637);
or UO_199 (O_199,N_8087,N_8095);
or UO_200 (O_200,N_8817,N_9543);
nor UO_201 (O_201,N_8143,N_8619);
or UO_202 (O_202,N_9018,N_8788);
nor UO_203 (O_203,N_8147,N_8251);
nor UO_204 (O_204,N_8224,N_9029);
nand UO_205 (O_205,N_9425,N_8677);
nand UO_206 (O_206,N_8518,N_8888);
or UO_207 (O_207,N_8547,N_9187);
nand UO_208 (O_208,N_8613,N_8941);
or UO_209 (O_209,N_8835,N_8792);
and UO_210 (O_210,N_8215,N_9999);
nand UO_211 (O_211,N_9116,N_8340);
nand UO_212 (O_212,N_9925,N_8377);
or UO_213 (O_213,N_8059,N_9297);
nor UO_214 (O_214,N_9212,N_9758);
nand UO_215 (O_215,N_8894,N_8965);
and UO_216 (O_216,N_9221,N_8710);
or UO_217 (O_217,N_9033,N_8900);
nand UO_218 (O_218,N_8244,N_8164);
and UO_219 (O_219,N_8829,N_9344);
nor UO_220 (O_220,N_9441,N_8693);
nor UO_221 (O_221,N_9039,N_8039);
or UO_222 (O_222,N_8195,N_9406);
or UO_223 (O_223,N_8418,N_8306);
nor UO_224 (O_224,N_9285,N_8438);
nand UO_225 (O_225,N_9028,N_8362);
nand UO_226 (O_226,N_8804,N_9609);
nand UO_227 (O_227,N_9100,N_8543);
and UO_228 (O_228,N_9101,N_8774);
nand UO_229 (O_229,N_9823,N_9750);
nor UO_230 (O_230,N_9076,N_9693);
xor UO_231 (O_231,N_9567,N_9449);
nor UO_232 (O_232,N_9877,N_8830);
and UO_233 (O_233,N_8833,N_8129);
and UO_234 (O_234,N_9386,N_9862);
nand UO_235 (O_235,N_8564,N_9296);
nand UO_236 (O_236,N_9559,N_9480);
and UO_237 (O_237,N_8783,N_9509);
nand UO_238 (O_238,N_9647,N_9720);
nand UO_239 (O_239,N_8183,N_8366);
nor UO_240 (O_240,N_9495,N_8132);
nand UO_241 (O_241,N_8794,N_8665);
and UO_242 (O_242,N_9218,N_9397);
nor UO_243 (O_243,N_8452,N_8612);
nor UO_244 (O_244,N_9350,N_8513);
and UO_245 (O_245,N_8245,N_9006);
nor UO_246 (O_246,N_8486,N_8007);
nand UO_247 (O_247,N_9467,N_8692);
nor UO_248 (O_248,N_9555,N_9287);
nand UO_249 (O_249,N_8025,N_9905);
or UO_250 (O_250,N_9685,N_8089);
nand UO_251 (O_251,N_8943,N_9404);
nor UO_252 (O_252,N_9733,N_8509);
or UO_253 (O_253,N_8077,N_9209);
and UO_254 (O_254,N_8654,N_9704);
nand UO_255 (O_255,N_9620,N_8247);
nor UO_256 (O_256,N_9947,N_8946);
nor UO_257 (O_257,N_9825,N_8412);
and UO_258 (O_258,N_9181,N_8008);
nor UO_259 (O_259,N_9938,N_9083);
nor UO_260 (O_260,N_9926,N_8254);
or UO_261 (O_261,N_8046,N_8681);
and UO_262 (O_262,N_9889,N_8074);
nor UO_263 (O_263,N_9138,N_9024);
or UO_264 (O_264,N_9433,N_8927);
or UO_265 (O_265,N_9043,N_9056);
or UO_266 (O_266,N_9873,N_9428);
or UO_267 (O_267,N_9445,N_8929);
nor UO_268 (O_268,N_8345,N_9385);
and UO_269 (O_269,N_8379,N_9699);
or UO_270 (O_270,N_9440,N_8957);
nor UO_271 (O_271,N_9021,N_8241);
or UO_272 (O_272,N_8493,N_9478);
or UO_273 (O_273,N_8655,N_9914);
nand UO_274 (O_274,N_9817,N_9626);
and UO_275 (O_275,N_9258,N_9735);
nor UO_276 (O_276,N_9429,N_8799);
nor UO_277 (O_277,N_8186,N_8301);
or UO_278 (O_278,N_8514,N_9255);
or UO_279 (O_279,N_8227,N_9163);
and UO_280 (O_280,N_9675,N_8709);
nor UO_281 (O_281,N_8527,N_8404);
nor UO_282 (O_282,N_9394,N_8182);
nor UO_283 (O_283,N_8431,N_9320);
nand UO_284 (O_284,N_8515,N_9408);
or UO_285 (O_285,N_8219,N_9483);
nor UO_286 (O_286,N_9984,N_8924);
and UO_287 (O_287,N_8762,N_9413);
or UO_288 (O_288,N_8623,N_8944);
nor UO_289 (O_289,N_9173,N_8191);
nor UO_290 (O_290,N_8526,N_8053);
nor UO_291 (O_291,N_8450,N_9012);
and UO_292 (O_292,N_8290,N_8266);
nand UO_293 (O_293,N_8145,N_9624);
and UO_294 (O_294,N_8309,N_8178);
and UO_295 (O_295,N_8015,N_8787);
or UO_296 (O_296,N_8841,N_8958);
nand UO_297 (O_297,N_9578,N_8349);
and UO_298 (O_298,N_8127,N_8358);
nand UO_299 (O_299,N_8281,N_8597);
or UO_300 (O_300,N_9055,N_8346);
nor UO_301 (O_301,N_9236,N_9741);
and UO_302 (O_302,N_8696,N_8898);
or UO_303 (O_303,N_9575,N_9327);
and UO_304 (O_304,N_9503,N_9569);
nand UO_305 (O_305,N_8876,N_8428);
and UO_306 (O_306,N_8725,N_9731);
nand UO_307 (O_307,N_8375,N_8121);
nor UO_308 (O_308,N_8302,N_9805);
nor UO_309 (O_309,N_8642,N_8391);
or UO_310 (O_310,N_9058,N_8066);
or UO_311 (O_311,N_9894,N_8915);
and UO_312 (O_312,N_9921,N_9885);
nor UO_313 (O_313,N_8959,N_8636);
or UO_314 (O_314,N_9067,N_8703);
or UO_315 (O_315,N_9771,N_9328);
and UO_316 (O_316,N_8548,N_8987);
and UO_317 (O_317,N_9131,N_9794);
or UO_318 (O_318,N_9677,N_9188);
and UO_319 (O_319,N_9161,N_9786);
or UO_320 (O_320,N_8583,N_8570);
or UO_321 (O_321,N_8750,N_8851);
or UO_322 (O_322,N_8785,N_8761);
nand UO_323 (O_323,N_9919,N_8258);
nand UO_324 (O_324,N_9110,N_9579);
nand UO_325 (O_325,N_9847,N_8275);
and UO_326 (O_326,N_9095,N_8004);
nand UO_327 (O_327,N_9364,N_9228);
and UO_328 (O_328,N_8210,N_8933);
nor UO_329 (O_329,N_9472,N_9457);
nand UO_330 (O_330,N_9481,N_9051);
nor UO_331 (O_331,N_9410,N_8579);
nor UO_332 (O_332,N_8073,N_9745);
and UO_333 (O_333,N_8745,N_8749);
nor UO_334 (O_334,N_8307,N_9944);
nor UO_335 (O_335,N_8040,N_8594);
nand UO_336 (O_336,N_8263,N_9801);
nor UO_337 (O_337,N_8574,N_8474);
nand UO_338 (O_338,N_8069,N_8051);
or UO_339 (O_339,N_9124,N_9831);
nand UO_340 (O_340,N_9134,N_8967);
nor UO_341 (O_341,N_8268,N_9136);
nand UO_342 (O_342,N_9162,N_8990);
nand UO_343 (O_343,N_8386,N_9976);
and UO_344 (O_344,N_9780,N_8488);
or UO_345 (O_345,N_9081,N_9997);
or UO_346 (O_346,N_8648,N_9544);
or UO_347 (O_347,N_8413,N_9987);
and UO_348 (O_348,N_9485,N_8852);
and UO_349 (O_349,N_9375,N_9252);
nor UO_350 (O_350,N_9942,N_9605);
nand UO_351 (O_351,N_8814,N_9135);
or UO_352 (O_352,N_8062,N_9057);
or UO_353 (O_353,N_8650,N_9723);
and UO_354 (O_354,N_9760,N_9744);
and UO_355 (O_355,N_8157,N_9791);
nand UO_356 (O_356,N_9602,N_9353);
nor UO_357 (O_357,N_8261,N_9910);
or UO_358 (O_358,N_9515,N_8962);
nand UO_359 (O_359,N_9132,N_8432);
or UO_360 (O_360,N_9953,N_8017);
nand UO_361 (O_361,N_9774,N_9053);
and UO_362 (O_362,N_9703,N_9713);
or UO_363 (O_363,N_9512,N_9778);
nor UO_364 (O_364,N_9764,N_9443);
nand UO_365 (O_365,N_8328,N_8014);
or UO_366 (O_366,N_9442,N_8443);
nor UO_367 (O_367,N_8531,N_9253);
or UO_368 (O_368,N_8138,N_8964);
and UO_369 (O_369,N_9468,N_9802);
or UO_370 (O_370,N_9644,N_9008);
nand UO_371 (O_371,N_8628,N_8727);
nor UO_372 (O_372,N_9044,N_9245);
nor UO_373 (O_373,N_8497,N_9743);
nor UO_374 (O_374,N_9369,N_8234);
or UO_375 (O_375,N_8151,N_9414);
nand UO_376 (O_376,N_8341,N_8372);
and UO_377 (O_377,N_8336,N_9427);
nand UO_378 (O_378,N_8715,N_9739);
xor UO_379 (O_379,N_9349,N_9838);
and UO_380 (O_380,N_8769,N_8637);
nor UO_381 (O_381,N_9234,N_9389);
or UO_382 (O_382,N_8131,N_8961);
nor UO_383 (O_383,N_8858,N_9846);
nand UO_384 (O_384,N_8300,N_9391);
nand UO_385 (O_385,N_9300,N_8555);
and UO_386 (O_386,N_8823,N_9048);
and UO_387 (O_387,N_8154,N_9940);
and UO_388 (O_388,N_9426,N_9298);
nand UO_389 (O_389,N_9781,N_9002);
or UO_390 (O_390,N_9570,N_8397);
nor UO_391 (O_391,N_9826,N_9080);
nor UO_392 (O_392,N_9403,N_9576);
and UO_393 (O_393,N_9549,N_8554);
or UO_394 (O_394,N_8417,N_9840);
and UO_395 (O_395,N_8722,N_9972);
and UO_396 (O_396,N_8447,N_9935);
nand UO_397 (O_397,N_8323,N_8465);
or UO_398 (O_398,N_8325,N_8113);
nand UO_399 (O_399,N_9561,N_9448);
and UO_400 (O_400,N_9334,N_8284);
or UO_401 (O_401,N_8698,N_8816);
nor UO_402 (O_402,N_8023,N_8295);
nor UO_403 (O_403,N_9184,N_9363);
and UO_404 (O_404,N_8350,N_8826);
nor UO_405 (O_405,N_8742,N_9224);
nand UO_406 (O_406,N_8109,N_9038);
nand UO_407 (O_407,N_9815,N_8376);
xor UO_408 (O_408,N_9582,N_8728);
and UO_409 (O_409,N_9338,N_8043);
nor UO_410 (O_410,N_8842,N_9401);
nand UO_411 (O_411,N_9185,N_9571);
or UO_412 (O_412,N_9233,N_8635);
or UO_413 (O_413,N_9564,N_9965);
and UO_414 (O_414,N_8209,N_9834);
nand UO_415 (O_415,N_9674,N_8461);
and UO_416 (O_416,N_8824,N_8881);
and UO_417 (O_417,N_9518,N_8850);
nand UO_418 (O_418,N_8732,N_9111);
and UO_419 (O_419,N_8180,N_8410);
and UO_420 (O_420,N_8464,N_8813);
nand UO_421 (O_421,N_9226,N_8688);
nand UO_422 (O_422,N_8380,N_8624);
nand UO_423 (O_423,N_8978,N_8954);
nand UO_424 (O_424,N_8831,N_9204);
or UO_425 (O_425,N_9330,N_8176);
and UO_426 (O_426,N_9398,N_9763);
or UO_427 (O_427,N_9329,N_9901);
nand UO_428 (O_428,N_8604,N_9199);
nor UO_429 (O_429,N_8181,N_9115);
nand UO_430 (O_430,N_8250,N_9691);
nor UO_431 (O_431,N_8569,N_9783);
and UO_432 (O_432,N_8333,N_8714);
and UO_433 (O_433,N_9331,N_9195);
nand UO_434 (O_434,N_8489,N_9312);
nand UO_435 (O_435,N_9273,N_9539);
and UO_436 (O_436,N_9430,N_9261);
or UO_437 (O_437,N_9086,N_8123);
and UO_438 (O_438,N_9283,N_8337);
nand UO_439 (O_439,N_9962,N_8298);
nand UO_440 (O_440,N_9738,N_9157);
nand UO_441 (O_441,N_9599,N_9523);
or UO_442 (O_442,N_9903,N_9309);
and UO_443 (O_443,N_9577,N_9254);
or UO_444 (O_444,N_8884,N_9886);
nand UO_445 (O_445,N_9272,N_9421);
nor UO_446 (O_446,N_9460,N_9590);
nand UO_447 (O_447,N_8791,N_8398);
or UO_448 (O_448,N_9646,N_8318);
and UO_449 (O_449,N_8716,N_9890);
or UO_450 (O_450,N_9219,N_8368);
nor UO_451 (O_451,N_8165,N_8494);
or UO_452 (O_452,N_8141,N_9893);
or UO_453 (O_453,N_8687,N_9062);
nor UO_454 (O_454,N_8982,N_9474);
nor UO_455 (O_455,N_8986,N_8454);
or UO_456 (O_456,N_9073,N_8499);
and UO_457 (O_457,N_9900,N_8448);
and UO_458 (O_458,N_9059,N_9007);
and UO_459 (O_459,N_9505,N_8439);
nand UO_460 (O_460,N_8553,N_8923);
or UO_461 (O_461,N_8904,N_9524);
nor UO_462 (O_462,N_8971,N_8773);
or UO_463 (O_463,N_9244,N_8065);
nand UO_464 (O_464,N_9702,N_9091);
and UO_465 (O_465,N_9973,N_8828);
or UO_466 (O_466,N_9688,N_9250);
or UO_467 (O_467,N_8446,N_8482);
and UO_468 (O_468,N_9534,N_9351);
nor UO_469 (O_469,N_9629,N_9380);
and UO_470 (O_470,N_9736,N_8506);
or UO_471 (O_471,N_8501,N_8230);
and UO_472 (O_472,N_9673,N_8255);
or UO_473 (O_473,N_8469,N_8975);
nor UO_474 (O_474,N_9548,N_8741);
or UO_475 (O_475,N_9598,N_9362);
or UO_476 (O_476,N_8679,N_8925);
nor UO_477 (O_477,N_8919,N_8674);
nor UO_478 (O_478,N_8359,N_8424);
nand UO_479 (O_479,N_8866,N_8731);
nand UO_480 (O_480,N_8562,N_9974);
nor UO_481 (O_481,N_8573,N_9498);
nor UO_482 (O_482,N_8477,N_9892);
nor UO_483 (O_483,N_8966,N_8194);
nand UO_484 (O_484,N_9096,N_8832);
or UO_485 (O_485,N_8406,N_9967);
and UO_486 (O_486,N_9269,N_9983);
nand UO_487 (O_487,N_9928,N_9167);
nand UO_488 (O_488,N_9684,N_8264);
nor UO_489 (O_489,N_9681,N_9222);
nand UO_490 (O_490,N_8546,N_8544);
or UO_491 (O_491,N_8921,N_9292);
or UO_492 (O_492,N_8135,N_8937);
or UO_493 (O_493,N_8274,N_8355);
and UO_494 (O_494,N_9126,N_8955);
and UO_495 (O_495,N_9015,N_9004);
or UO_496 (O_496,N_8102,N_9326);
nand UO_497 (O_497,N_8256,N_8152);
and UO_498 (O_498,N_9490,N_8740);
nand UO_499 (O_499,N_9717,N_9208);
nand UO_500 (O_500,N_9034,N_9707);
or UO_501 (O_501,N_9295,N_8985);
nor UO_502 (O_502,N_9779,N_9160);
and UO_503 (O_503,N_8836,N_8331);
and UO_504 (O_504,N_9697,N_9906);
nor UO_505 (O_505,N_9205,N_8042);
nor UO_506 (O_506,N_9857,N_8305);
nor UO_507 (O_507,N_9989,N_8620);
and UO_508 (O_508,N_8691,N_8885);
and UO_509 (O_509,N_9607,N_8435);
xor UO_510 (O_510,N_8508,N_8363);
nand UO_511 (O_511,N_8032,N_8149);
or UO_512 (O_512,N_8000,N_9891);
nor UO_513 (O_513,N_8734,N_9835);
or UO_514 (O_514,N_8664,N_9119);
or UO_515 (O_515,N_9557,N_9041);
or UO_516 (O_516,N_9277,N_9323);
nand UO_517 (O_517,N_9423,N_8536);
nor UO_518 (O_518,N_9223,N_9260);
xor UO_519 (O_519,N_9852,N_9580);
nor UO_520 (O_520,N_9066,N_8348);
nor UO_521 (O_521,N_8909,N_8278);
or UO_522 (O_522,N_8934,N_8496);
or UO_523 (O_523,N_8381,N_8189);
or UO_524 (O_524,N_9141,N_9520);
or UO_525 (O_525,N_9159,N_9844);
nand UO_526 (O_526,N_8663,N_9294);
and UO_527 (O_527,N_8916,N_9961);
or UO_528 (O_528,N_9179,N_9537);
nor UO_529 (O_529,N_9589,N_8229);
nor UO_530 (O_530,N_8632,N_9884);
and UO_531 (O_531,N_8031,N_9418);
or UO_532 (O_532,N_9489,N_9639);
nor UO_533 (O_533,N_9174,N_9770);
or UO_534 (O_534,N_8524,N_8706);
or UO_535 (O_535,N_9992,N_8427);
and UO_536 (O_536,N_8911,N_9843);
nor UO_537 (O_537,N_8631,N_9112);
nor UO_538 (O_538,N_8018,N_9625);
nand UO_539 (O_539,N_8262,N_9169);
and UO_540 (O_540,N_8394,N_8670);
nand UO_541 (O_541,N_9455,N_8805);
or UO_542 (O_542,N_8179,N_9610);
and UO_543 (O_543,N_9289,N_9833);
and UO_544 (O_544,N_8169,N_9247);
and UO_545 (O_545,N_8479,N_9618);
nand UO_546 (O_546,N_8421,N_9819);
and UO_547 (O_547,N_9510,N_8589);
nor UO_548 (O_548,N_9753,N_9026);
and UO_549 (O_549,N_9710,N_9231);
or UO_550 (O_550,N_9016,N_9875);
nor UO_551 (O_551,N_8011,N_8652);
nor UO_552 (O_552,N_8721,N_9726);
nand UO_553 (O_553,N_9651,N_9230);
nor UO_554 (O_554,N_8931,N_8096);
and UO_555 (O_555,N_8992,N_9991);
nor UO_556 (O_556,N_9360,N_8225);
and UO_557 (O_557,N_8107,N_8905);
or UO_558 (O_558,N_9014,N_9859);
nand UO_559 (O_559,N_8581,N_8854);
nand UO_560 (O_560,N_9290,N_9979);
and UO_561 (O_561,N_8078,N_8701);
and UO_562 (O_562,N_8576,N_8879);
nand UO_563 (O_563,N_8600,N_9166);
or UO_564 (O_564,N_9916,N_8126);
xnor UO_565 (O_565,N_9013,N_8840);
nand UO_566 (O_566,N_9267,N_8236);
nand UO_567 (O_567,N_8882,N_8766);
and UO_568 (O_568,N_9516,N_9766);
and UO_569 (O_569,N_8770,N_8798);
nor UO_570 (O_570,N_8800,N_8818);
and UO_571 (O_571,N_8656,N_8384);
or UO_572 (O_572,N_8028,N_9728);
nor UO_573 (O_573,N_9399,N_9070);
or UO_574 (O_574,N_8902,N_9103);
nand UO_575 (O_575,N_8112,N_8248);
nor UO_576 (O_576,N_8170,N_8283);
or UO_577 (O_577,N_8626,N_9145);
or UO_578 (O_578,N_8686,N_8865);
or UO_579 (O_579,N_9856,N_9147);
nand UO_580 (O_580,N_8060,N_9711);
nor UO_581 (O_581,N_9001,N_9742);
or UO_582 (O_582,N_8239,N_8315);
nor UO_583 (O_583,N_8330,N_8222);
nand UO_584 (O_584,N_9148,N_9622);
nor UO_585 (O_585,N_8175,N_8666);
and UO_586 (O_586,N_9671,N_9288);
and UO_587 (O_587,N_8563,N_8361);
or UO_588 (O_588,N_8903,N_9672);
or UO_589 (O_589,N_8775,N_9768);
nor UO_590 (O_590,N_8598,N_9486);
and UO_591 (O_591,N_9407,N_8403);
nand UO_592 (O_592,N_9592,N_9494);
and UO_593 (O_593,N_9031,N_9632);
and UO_594 (O_594,N_8976,N_9842);
nand UO_595 (O_595,N_9895,N_9374);
xnor UO_596 (O_596,N_9718,N_8723);
or UO_597 (O_597,N_9931,N_8118);
or UO_598 (O_598,N_8712,N_9341);
nor UO_599 (O_599,N_9027,N_8334);
xnor UO_600 (O_600,N_8837,N_9619);
nor UO_601 (O_601,N_8395,N_9354);
nand UO_602 (O_602,N_8592,N_9854);
nand UO_603 (O_603,N_9874,N_9102);
nand UO_604 (O_604,N_8374,N_8103);
or UO_605 (O_605,N_8950,N_9099);
and UO_606 (O_606,N_9186,N_9390);
nand UO_607 (O_607,N_8253,N_8896);
nand UO_608 (O_608,N_8864,N_9532);
nor UO_609 (O_609,N_8871,N_8827);
and UO_610 (O_610,N_9125,N_8010);
and UO_611 (O_611,N_8206,N_9550);
nor UO_612 (O_612,N_8609,N_8144);
and UO_613 (O_613,N_9851,N_8156);
nor UO_614 (O_614,N_8124,N_9347);
and UO_615 (O_615,N_9307,N_9270);
and UO_616 (O_616,N_9104,N_9535);
and UO_617 (O_617,N_9719,N_9462);
nand UO_618 (O_618,N_8719,N_9396);
and UO_619 (O_619,N_8806,N_8657);
nor UO_620 (O_620,N_9776,N_9547);
and UO_621 (O_621,N_8796,N_8980);
nand UO_622 (O_622,N_9907,N_9573);
nand UO_623 (O_623,N_8205,N_8335);
nor UO_624 (O_624,N_8539,N_8200);
nand UO_625 (O_625,N_8019,N_9400);
nand UO_626 (O_626,N_8660,N_9274);
nor UO_627 (O_627,N_8155,N_8747);
and UO_628 (O_628,N_8409,N_9264);
nor UO_629 (O_629,N_8640,N_8899);
and UO_630 (O_630,N_9836,N_9882);
or UO_631 (O_631,N_9461,N_9491);
nand UO_632 (O_632,N_8276,N_9470);
or UO_633 (O_633,N_8081,N_9092);
nor UO_634 (O_634,N_9079,N_8226);
and UO_635 (O_635,N_9789,N_9558);
or UO_636 (O_636,N_9203,N_9596);
or UO_637 (O_637,N_8313,N_8538);
and UO_638 (O_638,N_9740,N_9994);
nand UO_639 (O_639,N_9170,N_9065);
or UO_640 (O_640,N_9988,N_9832);
xnor UO_641 (O_641,N_9654,N_9530);
and UO_642 (O_642,N_8700,N_9214);
or UO_643 (O_643,N_8617,N_8044);
xnor UO_644 (O_644,N_8549,N_9243);
nand UO_645 (O_645,N_9355,N_8606);
or UO_646 (O_646,N_8476,N_9465);
and UO_647 (O_647,N_9909,N_8809);
nor UO_648 (O_648,N_8322,N_8697);
or UO_649 (O_649,N_8168,N_8970);
nor UO_650 (O_650,N_9340,N_9504);
nor UO_651 (O_651,N_8420,N_9860);
or UO_652 (O_652,N_9376,N_9085);
xor UO_653 (O_653,N_9335,N_8695);
nor UO_654 (O_654,N_9982,N_8936);
nor UO_655 (O_655,N_9957,N_9082);
nor UO_656 (O_656,N_8070,N_9379);
nor UO_657 (O_657,N_8273,N_8083);
and UO_658 (O_658,N_9737,N_9493);
nand UO_659 (O_659,N_9315,N_8780);
nor UO_660 (O_660,N_9995,N_8694);
nand UO_661 (O_661,N_9908,N_9220);
or UO_662 (O_662,N_8786,N_8952);
or UO_663 (O_663,N_8638,N_9584);
or UO_664 (O_664,N_9482,N_8192);
nor UO_665 (O_665,N_8561,N_8529);
nand UO_666 (O_666,N_9661,N_8441);
and UO_667 (O_667,N_9769,N_9370);
and UO_668 (O_668,N_9899,N_8166);
nor UO_669 (O_669,N_8685,N_8100);
and UO_670 (O_670,N_9521,N_8332);
and UO_671 (O_671,N_8812,N_9266);
or UO_672 (O_672,N_8795,N_8843);
and UO_673 (O_673,N_8901,N_8216);
nor UO_674 (O_674,N_8819,N_8271);
or UO_675 (O_675,N_8558,N_8402);
nor UO_676 (O_676,N_8528,N_8729);
nor UO_677 (O_677,N_8260,N_9787);
nand UO_678 (O_678,N_9551,N_9507);
and UO_679 (O_679,N_8999,N_8279);
or UO_680 (O_680,N_9352,N_9182);
and UO_681 (O_681,N_9636,N_9042);
nor UO_682 (O_682,N_9712,N_8037);
or UO_683 (O_683,N_9431,N_9814);
and UO_684 (O_684,N_8422,N_9784);
and UO_685 (O_685,N_8735,N_8682);
nand UO_686 (O_686,N_8897,N_8516);
nand UO_687 (O_687,N_8847,N_8079);
nand UO_688 (O_688,N_9439,N_8075);
nor UO_689 (O_689,N_9054,N_9183);
nor UO_690 (O_690,N_8839,N_8148);
and UO_691 (O_691,N_8857,N_9310);
nor UO_692 (O_692,N_9129,N_9949);
and UO_693 (O_693,N_8228,N_8048);
or UO_694 (O_694,N_8545,N_8433);
or UO_695 (O_695,N_9215,N_8204);
nand UO_696 (O_696,N_8675,N_9225);
and UO_697 (O_697,N_9705,N_9381);
or UO_698 (O_698,N_9828,N_9955);
and UO_699 (O_699,N_9499,N_9251);
nor UO_700 (O_700,N_8616,N_8932);
and UO_701 (O_701,N_9706,N_9180);
nor UO_702 (O_702,N_8673,N_9793);
or UO_703 (O_703,N_8167,N_8511);
and UO_704 (O_704,N_8396,N_8680);
and UO_705 (O_705,N_9324,N_8303);
or UO_706 (O_706,N_9318,N_9816);
and UO_707 (O_707,N_9271,N_9643);
nand UO_708 (O_708,N_8746,N_8639);
nand UO_709 (O_709,N_8586,N_8214);
and UO_710 (O_710,N_8137,N_8537);
or UO_711 (O_711,N_9917,N_9820);
nor UO_712 (O_712,N_9980,N_9951);
or UO_713 (O_713,N_9475,N_8759);
or UO_714 (O_714,N_8436,N_8389);
nand UO_715 (O_715,N_8878,N_9680);
nor UO_716 (O_716,N_9960,N_9734);
xnor UO_717 (O_717,N_8016,N_8575);
and UO_718 (O_718,N_9841,N_8237);
and UO_719 (O_719,N_9511,N_9853);
and UO_720 (O_720,N_9642,N_8106);
nor UO_721 (O_721,N_9545,N_9193);
or UO_722 (O_722,N_8790,N_9194);
nor UO_723 (O_723,N_8500,N_9950);
nand UO_724 (O_724,N_8371,N_9087);
nand UO_725 (O_725,N_8473,N_9464);
nand UO_726 (O_726,N_8055,N_9513);
or UO_727 (O_727,N_9747,N_8187);
and UO_728 (O_728,N_8211,N_9649);
and UO_729 (O_729,N_8411,N_8503);
nand UO_730 (O_730,N_8292,N_9855);
nand UO_731 (O_731,N_8163,N_8646);
or UO_732 (O_732,N_8689,N_9452);
or UO_733 (O_733,N_8998,N_9663);
nor UO_734 (O_734,N_8162,N_9030);
or UO_735 (O_735,N_9878,N_8808);
nand UO_736 (O_736,N_8767,N_8855);
or UO_737 (O_737,N_8470,N_9450);
and UO_738 (O_738,N_8392,N_8533);
nand UO_739 (O_739,N_9077,N_8071);
nor UO_740 (O_740,N_9682,N_9359);
and UO_741 (O_741,N_9417,N_9790);
and UO_742 (O_742,N_9388,N_8320);
or UO_743 (O_743,N_8705,N_8076);
xor UO_744 (O_744,N_8920,N_9052);
or UO_745 (O_745,N_9613,N_8463);
and UO_746 (O_746,N_9144,N_8369);
nand UO_747 (O_747,N_8880,N_9239);
and UO_748 (O_748,N_9248,N_9813);
nor UO_749 (O_749,N_8707,N_8084);
nand UO_750 (O_750,N_9898,N_9206);
nand UO_751 (O_751,N_9128,N_9803);
or UO_752 (O_752,N_8199,N_9496);
and UO_753 (O_753,N_8772,N_8086);
and UO_754 (O_754,N_9746,N_9094);
nor UO_755 (O_755,N_9010,N_8552);
and UO_756 (O_756,N_9121,N_8956);
nand UO_757 (O_757,N_8505,N_8423);
and UO_758 (O_758,N_8400,N_8711);
and UO_759 (O_759,N_9572,N_8627);
or UO_760 (O_760,N_8122,N_8502);
or UO_761 (O_761,N_9422,N_8257);
or UO_762 (O_762,N_9959,N_8414);
nand UO_763 (O_763,N_9089,N_8930);
or UO_764 (O_764,N_9667,N_9756);
nor UO_765 (O_765,N_8601,N_9721);
or UO_766 (O_766,N_9837,N_8983);
and UO_767 (O_767,N_9689,N_9286);
or UO_768 (O_768,N_8540,N_8357);
nand UO_769 (O_769,N_9946,N_8159);
nand UO_770 (O_770,N_8763,N_9686);
nor UO_771 (O_771,N_9114,N_9581);
nand UO_772 (O_772,N_8231,N_8845);
or UO_773 (O_773,N_9656,N_9164);
nor UO_774 (O_774,N_8684,N_9645);
and UO_775 (O_775,N_8869,N_8997);
nor UO_776 (O_776,N_8035,N_8153);
nand UO_777 (O_777,N_8668,N_8906);
or UO_778 (O_778,N_9845,N_9913);
nand UO_779 (O_779,N_8440,N_9650);
nor UO_780 (O_780,N_8299,N_9727);
and UO_781 (O_781,N_9411,N_8541);
and UO_782 (O_782,N_9522,N_8462);
or UO_783 (O_783,N_8892,N_8848);
and UO_784 (O_784,N_9149,N_9948);
nor UO_785 (O_785,N_9045,N_8690);
nor UO_786 (O_786,N_8282,N_9531);
nor UO_787 (O_787,N_9700,N_9003);
and UO_788 (O_788,N_9268,N_8914);
nor UO_789 (O_789,N_8339,N_9078);
and UO_790 (O_790,N_9755,N_8893);
nand UO_791 (O_791,N_8634,N_8661);
nor UO_792 (O_792,N_8312,N_8651);
and UO_793 (O_793,N_8724,N_9093);
nand UO_794 (O_794,N_8963,N_9538);
or UO_795 (O_795,N_8565,N_9554);
nand UO_796 (O_796,N_8849,N_9709);
or UO_797 (O_797,N_8353,N_8020);
nor UO_798 (O_798,N_8259,N_9929);
or UO_799 (O_799,N_8468,N_8890);
and UO_800 (O_800,N_9611,N_9227);
or UO_801 (O_801,N_8622,N_8061);
nand UO_802 (O_802,N_8390,N_8603);
nand UO_803 (O_803,N_8996,N_9419);
nor UO_804 (O_804,N_9084,N_9151);
and UO_805 (O_805,N_8887,N_8889);
or UO_806 (O_806,N_9301,N_8267);
and UO_807 (O_807,N_9978,N_8116);
nand UO_808 (O_808,N_8993,N_8090);
nor UO_809 (O_809,N_9795,N_9476);
and UO_810 (O_810,N_8415,N_8873);
or UO_811 (O_811,N_8088,N_9123);
or UO_812 (O_812,N_8672,N_9977);
or UO_813 (O_813,N_9546,N_8726);
and UO_814 (O_814,N_8752,N_8057);
nand UO_815 (O_815,N_8870,N_9319);
or UO_816 (O_816,N_8277,N_8781);
or UO_817 (O_817,N_8310,N_9152);
nor UO_818 (O_818,N_9263,N_8861);
or UO_819 (O_819,N_8136,N_9322);
nor UO_820 (O_820,N_8453,N_8608);
nor UO_821 (O_821,N_9676,N_9207);
and UO_822 (O_822,N_9653,N_9438);
and UO_823 (O_823,N_9506,N_8922);
nor UO_824 (O_824,N_9176,N_9748);
nand UO_825 (O_825,N_9210,N_8430);
nand UO_826 (O_826,N_9648,N_8036);
or UO_827 (O_827,N_9046,N_8560);
nand UO_828 (O_828,N_9633,N_9368);
nand UO_829 (O_829,N_8487,N_8807);
or UO_830 (O_830,N_8094,N_9552);
and UO_831 (O_831,N_9759,N_8662);
and UO_832 (O_832,N_8777,N_8343);
and UO_833 (O_833,N_8022,N_8050);
or UO_834 (O_834,N_8426,N_9902);
and UO_835 (O_835,N_9501,N_8405);
nor UO_836 (O_836,N_8649,N_9923);
or UO_837 (O_837,N_9311,N_8517);
and UO_838 (O_838,N_9200,N_8585);
and UO_839 (O_839,N_8519,N_9122);
and UO_840 (O_840,N_8091,N_8188);
or UO_841 (O_841,N_8459,N_9621);
and UO_842 (O_842,N_9911,N_8177);
nand UO_843 (O_843,N_8467,N_8150);
and UO_844 (O_844,N_8142,N_8853);
nor UO_845 (O_845,N_8471,N_9986);
nor UO_846 (O_846,N_9601,N_8294);
nand UO_847 (O_847,N_8444,N_8633);
nor UO_848 (O_848,N_9945,N_9775);
nor UO_849 (O_849,N_8556,N_8875);
nand UO_850 (O_850,N_8951,N_9807);
and UO_851 (O_851,N_8713,N_8481);
and UO_852 (O_852,N_8208,N_8308);
or UO_853 (O_853,N_9257,N_8172);
and UO_854 (O_854,N_8653,N_9767);
nor UO_855 (O_855,N_9420,N_9553);
xor UO_856 (O_856,N_8383,N_8591);
or UO_857 (O_857,N_8981,N_9306);
nand UO_858 (O_858,N_9178,N_8610);
nor UO_859 (O_859,N_9519,N_8991);
nor UO_860 (O_860,N_8571,N_9032);
or UO_861 (O_861,N_9729,N_9120);
nand UO_862 (O_862,N_8736,N_8989);
nor UO_863 (O_863,N_9757,N_9050);
nand UO_864 (O_864,N_8030,N_8041);
nand UO_865 (O_865,N_8940,N_9958);
nor UO_866 (O_866,N_8249,N_8314);
nor UO_867 (O_867,N_9118,N_8949);
or UO_868 (O_868,N_8578,N_8757);
or UO_869 (O_869,N_9871,N_9367);
or UO_870 (O_870,N_9867,N_9500);
and UO_871 (O_871,N_9830,N_8108);
nor UO_872 (O_872,N_8327,N_8202);
nor UO_873 (O_873,N_9829,N_9804);
and UO_874 (O_874,N_9556,N_8316);
or UO_875 (O_875,N_8867,N_9321);
and UO_876 (O_876,N_8221,N_9177);
nor UO_877 (O_877,N_9035,N_9808);
nor UO_878 (O_878,N_8507,N_9593);
nand UO_879 (O_879,N_8472,N_8064);
nand UO_880 (O_880,N_9872,N_8551);
or UO_881 (O_881,N_8615,N_8475);
and UO_882 (O_882,N_9107,N_8730);
or UO_883 (O_883,N_8484,N_9358);
or UO_884 (O_884,N_9336,N_9799);
nand UO_885 (O_885,N_8708,N_8778);
or UO_886 (O_886,N_8297,N_8280);
nand UO_887 (O_887,N_9603,N_8643);
or UO_888 (O_888,N_8737,N_8557);
nand UO_889 (O_889,N_8197,N_8883);
nand UO_890 (O_890,N_9870,N_8815);
nand UO_891 (O_891,N_9060,N_9640);
or UO_892 (O_892,N_8203,N_8784);
and UO_893 (O_893,N_8972,N_9436);
or UO_894 (O_894,N_8580,N_8006);
nand UO_895 (O_895,N_8416,N_9694);
nor UO_896 (O_896,N_9562,N_8891);
or UO_897 (O_897,N_8822,N_9588);
nand UO_898 (O_898,N_9011,N_8480);
and UO_899 (O_899,N_8699,N_8825);
and UO_900 (O_900,N_8625,N_9069);
nand UO_901 (O_901,N_9525,N_8756);
nor UO_902 (O_902,N_9074,N_9773);
or UO_903 (O_903,N_8027,N_8001);
or UO_904 (O_904,N_8373,N_8645);
nor UO_905 (O_905,N_9415,N_9594);
nand UO_906 (O_906,N_8058,N_9585);
nand UO_907 (O_907,N_8296,N_9142);
or UO_908 (O_908,N_8218,N_8935);
nor UO_909 (O_909,N_8868,N_8838);
nor UO_910 (O_910,N_8968,N_9384);
or UO_911 (O_911,N_8510,N_8644);
and UO_912 (O_912,N_8105,N_9865);
nand UO_913 (O_913,N_8754,N_8618);
nand UO_914 (O_914,N_9497,N_9291);
nor UO_915 (O_915,N_8820,N_8630);
and UO_916 (O_916,N_9583,N_9240);
nand UO_917 (O_917,N_9037,N_8196);
nor UO_918 (O_918,N_9075,N_8393);
and UO_919 (O_919,N_9761,N_9302);
nor UO_920 (O_920,N_8201,N_8442);
or UO_921 (O_921,N_9217,N_8092);
or UO_922 (O_922,N_8801,N_8588);
nand UO_923 (O_923,N_9566,N_8344);
and UO_924 (O_924,N_9679,N_8099);
or UO_925 (O_925,N_9357,N_9308);
or UO_926 (O_926,N_9824,N_8595);
or UO_927 (O_927,N_9109,N_8895);
and UO_928 (O_928,N_8974,N_8329);
nor UO_929 (O_929,N_8291,N_9378);
nor UO_930 (O_930,N_9920,N_8863);
nor UO_931 (O_931,N_9345,N_8451);
nor UO_932 (O_932,N_8659,N_9090);
or UO_933 (O_933,N_9432,N_8171);
nor UO_934 (O_934,N_9471,N_9140);
or UO_935 (O_935,N_8797,N_8449);
or UO_936 (O_936,N_9668,N_9049);
nand UO_937 (O_937,N_9941,N_8720);
or UO_938 (O_938,N_8005,N_9293);
or UO_939 (O_939,N_9692,N_9040);
nand UO_940 (O_940,N_9888,N_9876);
and UO_941 (O_941,N_8938,N_9932);
and UO_942 (O_942,N_9527,N_9606);
nor UO_943 (O_943,N_9165,N_8678);
and UO_944 (O_944,N_9213,N_8647);
and UO_945 (O_945,N_8988,N_9009);
nand UO_946 (O_946,N_9634,N_8504);
and UO_947 (O_947,N_8733,N_9402);
nand UO_948 (O_948,N_8455,N_8572);
nor UO_949 (O_949,N_9366,N_8918);
or UO_950 (O_950,N_9924,N_9246);
nor UO_951 (O_951,N_9998,N_8045);
or UO_952 (O_952,N_9927,N_9036);
nand UO_953 (O_953,N_8356,N_8128);
and UO_954 (O_954,N_9887,N_8748);
and UO_955 (O_955,N_8382,N_9785);
nand UO_956 (O_956,N_9459,N_9683);
nor UO_957 (O_957,N_8641,N_8072);
nand UO_958 (O_958,N_8370,N_9492);
nand UO_959 (O_959,N_9265,N_9797);
nor UO_960 (O_960,N_8207,N_8125);
nor UO_961 (O_961,N_9565,N_8810);
and UO_962 (O_962,N_8995,N_8067);
and UO_963 (O_963,N_9956,N_8139);
or UO_964 (O_964,N_9197,N_9098);
or UO_965 (O_965,N_8024,N_8364);
and UO_966 (O_966,N_8117,N_9528);
and UO_967 (O_967,N_8287,N_8860);
and UO_968 (O_968,N_8525,N_9342);
nand UO_969 (O_969,N_9127,N_9880);
nor UO_970 (O_970,N_8434,N_8223);
nand UO_971 (O_971,N_9447,N_9630);
and UO_972 (O_972,N_9337,N_8319);
or UO_973 (O_973,N_9022,N_8942);
or UO_974 (O_974,N_9020,N_8429);
nor UO_975 (O_975,N_8491,N_9454);
nor UO_976 (O_976,N_8093,N_8611);
or UO_977 (O_977,N_9238,N_9730);
or UO_978 (O_978,N_9655,N_9153);
and UO_979 (O_979,N_8568,N_9299);
nand UO_980 (O_980,N_9996,N_8360);
nand UO_981 (O_981,N_8753,N_9617);
nand UO_982 (O_982,N_8445,N_8101);
or UO_983 (O_983,N_9724,N_8408);
or UO_984 (O_984,N_9373,N_9201);
or UO_985 (O_985,N_8365,N_9604);
and UO_986 (O_986,N_9670,N_8910);
or UO_987 (O_987,N_8802,N_9971);
or UO_988 (O_988,N_8243,N_9158);
nand UO_989 (O_989,N_8367,N_8460);
nand UO_990 (O_990,N_8111,N_9896);
and UO_991 (O_991,N_8385,N_9409);
nand UO_992 (O_992,N_9139,N_9333);
or UO_993 (O_993,N_9332,N_9934);
nor UO_994 (O_994,N_8846,N_9017);
and UO_995 (O_995,N_9981,N_8033);
and UO_996 (O_996,N_8834,N_8246);
and UO_997 (O_997,N_9171,N_9990);
and UO_998 (O_998,N_8425,N_8758);
nand UO_999 (O_999,N_8193,N_8593);
and UO_1000 (O_1000,N_8967,N_8268);
or UO_1001 (O_1001,N_8951,N_8760);
nor UO_1002 (O_1002,N_9650,N_9476);
or UO_1003 (O_1003,N_9764,N_8587);
nor UO_1004 (O_1004,N_9041,N_8613);
nand UO_1005 (O_1005,N_8159,N_8747);
or UO_1006 (O_1006,N_9845,N_8459);
or UO_1007 (O_1007,N_9543,N_9287);
and UO_1008 (O_1008,N_8423,N_8524);
or UO_1009 (O_1009,N_8663,N_8000);
nor UO_1010 (O_1010,N_9855,N_8351);
or UO_1011 (O_1011,N_8818,N_9571);
nor UO_1012 (O_1012,N_9202,N_9265);
nor UO_1013 (O_1013,N_8058,N_9604);
or UO_1014 (O_1014,N_8627,N_8582);
nand UO_1015 (O_1015,N_9948,N_9986);
and UO_1016 (O_1016,N_9698,N_8020);
and UO_1017 (O_1017,N_9458,N_8542);
or UO_1018 (O_1018,N_8326,N_8576);
nand UO_1019 (O_1019,N_9571,N_9121);
and UO_1020 (O_1020,N_9812,N_8599);
or UO_1021 (O_1021,N_9997,N_8805);
nand UO_1022 (O_1022,N_8294,N_8228);
nand UO_1023 (O_1023,N_9462,N_9467);
or UO_1024 (O_1024,N_8882,N_8944);
or UO_1025 (O_1025,N_8595,N_8634);
and UO_1026 (O_1026,N_9128,N_8738);
nor UO_1027 (O_1027,N_9858,N_8698);
nand UO_1028 (O_1028,N_8687,N_8224);
or UO_1029 (O_1029,N_8165,N_8536);
xor UO_1030 (O_1030,N_8161,N_8011);
nand UO_1031 (O_1031,N_8873,N_9707);
or UO_1032 (O_1032,N_8578,N_9256);
and UO_1033 (O_1033,N_9681,N_9455);
nand UO_1034 (O_1034,N_8947,N_9977);
nor UO_1035 (O_1035,N_9301,N_8776);
or UO_1036 (O_1036,N_8576,N_9776);
nand UO_1037 (O_1037,N_9610,N_9341);
and UO_1038 (O_1038,N_8432,N_9019);
or UO_1039 (O_1039,N_9711,N_9624);
or UO_1040 (O_1040,N_8644,N_8030);
and UO_1041 (O_1041,N_8815,N_9003);
and UO_1042 (O_1042,N_8303,N_8699);
or UO_1043 (O_1043,N_9172,N_9603);
nor UO_1044 (O_1044,N_9385,N_9992);
and UO_1045 (O_1045,N_8144,N_9054);
or UO_1046 (O_1046,N_8970,N_8669);
nand UO_1047 (O_1047,N_9220,N_8768);
or UO_1048 (O_1048,N_8804,N_8924);
or UO_1049 (O_1049,N_9736,N_9535);
nand UO_1050 (O_1050,N_8633,N_9413);
and UO_1051 (O_1051,N_9291,N_8858);
nand UO_1052 (O_1052,N_8014,N_9126);
nor UO_1053 (O_1053,N_8186,N_9720);
nand UO_1054 (O_1054,N_8019,N_9274);
nor UO_1055 (O_1055,N_9068,N_9294);
and UO_1056 (O_1056,N_9990,N_9698);
and UO_1057 (O_1057,N_9127,N_9830);
nand UO_1058 (O_1058,N_9376,N_9234);
or UO_1059 (O_1059,N_9034,N_9274);
nor UO_1060 (O_1060,N_8391,N_9018);
or UO_1061 (O_1061,N_8436,N_8674);
nand UO_1062 (O_1062,N_8254,N_9990);
nor UO_1063 (O_1063,N_8610,N_8305);
nand UO_1064 (O_1064,N_9468,N_9611);
and UO_1065 (O_1065,N_9326,N_9458);
nand UO_1066 (O_1066,N_8905,N_8672);
nor UO_1067 (O_1067,N_8907,N_9508);
and UO_1068 (O_1068,N_9633,N_8098);
nand UO_1069 (O_1069,N_9061,N_8681);
or UO_1070 (O_1070,N_8692,N_8757);
and UO_1071 (O_1071,N_9166,N_9044);
and UO_1072 (O_1072,N_8959,N_8834);
nand UO_1073 (O_1073,N_9893,N_9123);
and UO_1074 (O_1074,N_8246,N_8002);
or UO_1075 (O_1075,N_9577,N_8689);
nor UO_1076 (O_1076,N_8563,N_8151);
nand UO_1077 (O_1077,N_8586,N_9966);
or UO_1078 (O_1078,N_9220,N_8688);
or UO_1079 (O_1079,N_9588,N_8200);
nor UO_1080 (O_1080,N_9679,N_8275);
nand UO_1081 (O_1081,N_8277,N_8044);
nor UO_1082 (O_1082,N_9041,N_8560);
or UO_1083 (O_1083,N_9965,N_9499);
and UO_1084 (O_1084,N_9176,N_8581);
or UO_1085 (O_1085,N_9679,N_8236);
or UO_1086 (O_1086,N_8326,N_9994);
or UO_1087 (O_1087,N_9326,N_8767);
and UO_1088 (O_1088,N_9989,N_9908);
nand UO_1089 (O_1089,N_8364,N_8225);
or UO_1090 (O_1090,N_8176,N_9410);
nand UO_1091 (O_1091,N_9133,N_9514);
nand UO_1092 (O_1092,N_8096,N_8793);
nand UO_1093 (O_1093,N_8263,N_9086);
nor UO_1094 (O_1094,N_9203,N_8750);
and UO_1095 (O_1095,N_8343,N_9401);
and UO_1096 (O_1096,N_9119,N_9897);
and UO_1097 (O_1097,N_8672,N_9958);
and UO_1098 (O_1098,N_9800,N_8836);
nand UO_1099 (O_1099,N_9728,N_8144);
or UO_1100 (O_1100,N_8207,N_9683);
or UO_1101 (O_1101,N_8636,N_8615);
nor UO_1102 (O_1102,N_9693,N_9123);
or UO_1103 (O_1103,N_9390,N_8782);
nand UO_1104 (O_1104,N_8601,N_9378);
or UO_1105 (O_1105,N_9593,N_9610);
or UO_1106 (O_1106,N_9826,N_9752);
and UO_1107 (O_1107,N_9026,N_9382);
nand UO_1108 (O_1108,N_8920,N_9345);
nor UO_1109 (O_1109,N_9465,N_8212);
nand UO_1110 (O_1110,N_9478,N_9613);
and UO_1111 (O_1111,N_9593,N_8745);
and UO_1112 (O_1112,N_8681,N_8118);
and UO_1113 (O_1113,N_8757,N_9962);
nand UO_1114 (O_1114,N_8820,N_9920);
nand UO_1115 (O_1115,N_8120,N_9027);
and UO_1116 (O_1116,N_8597,N_8685);
or UO_1117 (O_1117,N_8265,N_8698);
or UO_1118 (O_1118,N_8535,N_9320);
xor UO_1119 (O_1119,N_8034,N_9600);
nor UO_1120 (O_1120,N_9889,N_9450);
nor UO_1121 (O_1121,N_8826,N_8193);
nand UO_1122 (O_1122,N_8762,N_9916);
or UO_1123 (O_1123,N_9224,N_8178);
or UO_1124 (O_1124,N_8147,N_9646);
nor UO_1125 (O_1125,N_9395,N_8165);
and UO_1126 (O_1126,N_8767,N_9327);
and UO_1127 (O_1127,N_8399,N_8213);
or UO_1128 (O_1128,N_9406,N_8927);
nand UO_1129 (O_1129,N_9470,N_9958);
nand UO_1130 (O_1130,N_8079,N_9154);
nor UO_1131 (O_1131,N_8189,N_8535);
nor UO_1132 (O_1132,N_8847,N_8754);
nand UO_1133 (O_1133,N_8926,N_8287);
nor UO_1134 (O_1134,N_9777,N_9206);
and UO_1135 (O_1135,N_9433,N_9900);
or UO_1136 (O_1136,N_8443,N_9082);
or UO_1137 (O_1137,N_9086,N_8197);
nand UO_1138 (O_1138,N_9819,N_8813);
and UO_1139 (O_1139,N_9464,N_9348);
and UO_1140 (O_1140,N_8757,N_8748);
nor UO_1141 (O_1141,N_9728,N_9210);
or UO_1142 (O_1142,N_8138,N_9422);
nand UO_1143 (O_1143,N_9942,N_9419);
or UO_1144 (O_1144,N_8499,N_8347);
nand UO_1145 (O_1145,N_9955,N_9324);
and UO_1146 (O_1146,N_8761,N_9040);
or UO_1147 (O_1147,N_9203,N_8192);
nand UO_1148 (O_1148,N_9424,N_8456);
or UO_1149 (O_1149,N_9848,N_8863);
nor UO_1150 (O_1150,N_8326,N_8376);
nor UO_1151 (O_1151,N_8922,N_8443);
or UO_1152 (O_1152,N_8968,N_8956);
nand UO_1153 (O_1153,N_9195,N_9558);
nand UO_1154 (O_1154,N_9305,N_8503);
nand UO_1155 (O_1155,N_9446,N_8432);
nand UO_1156 (O_1156,N_9054,N_9114);
nor UO_1157 (O_1157,N_9018,N_9362);
and UO_1158 (O_1158,N_9548,N_8631);
xor UO_1159 (O_1159,N_9104,N_9180);
nand UO_1160 (O_1160,N_9163,N_8906);
or UO_1161 (O_1161,N_8501,N_8136);
or UO_1162 (O_1162,N_9708,N_9555);
nor UO_1163 (O_1163,N_9919,N_8021);
nor UO_1164 (O_1164,N_8625,N_8981);
nor UO_1165 (O_1165,N_8182,N_9539);
nand UO_1166 (O_1166,N_9305,N_9898);
or UO_1167 (O_1167,N_8313,N_8082);
nor UO_1168 (O_1168,N_9361,N_8221);
nand UO_1169 (O_1169,N_8657,N_9736);
nor UO_1170 (O_1170,N_8046,N_9169);
or UO_1171 (O_1171,N_9703,N_9880);
or UO_1172 (O_1172,N_8156,N_9180);
nand UO_1173 (O_1173,N_8287,N_8983);
or UO_1174 (O_1174,N_9287,N_8861);
and UO_1175 (O_1175,N_8055,N_9846);
and UO_1176 (O_1176,N_9188,N_8575);
nor UO_1177 (O_1177,N_8432,N_8930);
nor UO_1178 (O_1178,N_8114,N_9264);
or UO_1179 (O_1179,N_9764,N_8355);
or UO_1180 (O_1180,N_8470,N_9874);
or UO_1181 (O_1181,N_8234,N_8106);
nor UO_1182 (O_1182,N_8949,N_8537);
nand UO_1183 (O_1183,N_8074,N_8360);
nand UO_1184 (O_1184,N_8306,N_8268);
or UO_1185 (O_1185,N_9962,N_8352);
or UO_1186 (O_1186,N_8317,N_8625);
nor UO_1187 (O_1187,N_8833,N_9193);
nor UO_1188 (O_1188,N_9771,N_9495);
or UO_1189 (O_1189,N_8219,N_9819);
nand UO_1190 (O_1190,N_8958,N_8699);
nand UO_1191 (O_1191,N_8978,N_9794);
nor UO_1192 (O_1192,N_8298,N_8737);
nor UO_1193 (O_1193,N_9587,N_9690);
nand UO_1194 (O_1194,N_9290,N_8650);
and UO_1195 (O_1195,N_9749,N_9259);
nor UO_1196 (O_1196,N_8498,N_9430);
nor UO_1197 (O_1197,N_8359,N_8770);
nand UO_1198 (O_1198,N_8762,N_9968);
or UO_1199 (O_1199,N_8463,N_9377);
or UO_1200 (O_1200,N_9115,N_9490);
and UO_1201 (O_1201,N_9990,N_9139);
and UO_1202 (O_1202,N_9679,N_8653);
and UO_1203 (O_1203,N_9912,N_8615);
nand UO_1204 (O_1204,N_9473,N_8661);
nand UO_1205 (O_1205,N_8026,N_9302);
nor UO_1206 (O_1206,N_9196,N_9965);
or UO_1207 (O_1207,N_8504,N_9618);
nand UO_1208 (O_1208,N_9297,N_8903);
nand UO_1209 (O_1209,N_9295,N_8139);
nand UO_1210 (O_1210,N_8914,N_9356);
nor UO_1211 (O_1211,N_8698,N_9754);
nor UO_1212 (O_1212,N_8782,N_8196);
and UO_1213 (O_1213,N_8256,N_9110);
or UO_1214 (O_1214,N_9536,N_9450);
nor UO_1215 (O_1215,N_9189,N_9592);
and UO_1216 (O_1216,N_8149,N_8757);
and UO_1217 (O_1217,N_8892,N_9887);
nand UO_1218 (O_1218,N_8782,N_8038);
nor UO_1219 (O_1219,N_8910,N_9381);
nor UO_1220 (O_1220,N_8726,N_8190);
or UO_1221 (O_1221,N_9402,N_8570);
and UO_1222 (O_1222,N_9073,N_9346);
nand UO_1223 (O_1223,N_8009,N_9829);
nor UO_1224 (O_1224,N_8876,N_9861);
nand UO_1225 (O_1225,N_9817,N_9397);
nor UO_1226 (O_1226,N_9833,N_8280);
and UO_1227 (O_1227,N_9279,N_9137);
nand UO_1228 (O_1228,N_8604,N_8953);
and UO_1229 (O_1229,N_9509,N_9576);
and UO_1230 (O_1230,N_9873,N_8940);
nand UO_1231 (O_1231,N_8384,N_9344);
nor UO_1232 (O_1232,N_8822,N_9854);
nand UO_1233 (O_1233,N_9805,N_8487);
and UO_1234 (O_1234,N_9544,N_9262);
or UO_1235 (O_1235,N_9829,N_8797);
and UO_1236 (O_1236,N_9024,N_8145);
nor UO_1237 (O_1237,N_8191,N_8428);
or UO_1238 (O_1238,N_9950,N_8652);
or UO_1239 (O_1239,N_9997,N_8860);
nand UO_1240 (O_1240,N_9053,N_8544);
or UO_1241 (O_1241,N_8283,N_8545);
and UO_1242 (O_1242,N_9302,N_9924);
nand UO_1243 (O_1243,N_8449,N_8552);
nor UO_1244 (O_1244,N_8051,N_9552);
nor UO_1245 (O_1245,N_9079,N_9291);
nor UO_1246 (O_1246,N_8762,N_9733);
and UO_1247 (O_1247,N_9088,N_8009);
or UO_1248 (O_1248,N_9019,N_8724);
nor UO_1249 (O_1249,N_9125,N_9002);
xnor UO_1250 (O_1250,N_8972,N_9874);
or UO_1251 (O_1251,N_8490,N_9246);
or UO_1252 (O_1252,N_9457,N_9302);
and UO_1253 (O_1253,N_8150,N_8418);
nand UO_1254 (O_1254,N_9603,N_8047);
xnor UO_1255 (O_1255,N_9001,N_8753);
and UO_1256 (O_1256,N_9272,N_8092);
or UO_1257 (O_1257,N_9603,N_8419);
and UO_1258 (O_1258,N_9464,N_9724);
nand UO_1259 (O_1259,N_8709,N_8217);
and UO_1260 (O_1260,N_9022,N_9612);
or UO_1261 (O_1261,N_8088,N_8092);
nand UO_1262 (O_1262,N_9534,N_9086);
or UO_1263 (O_1263,N_9686,N_8324);
nand UO_1264 (O_1264,N_9185,N_9736);
nand UO_1265 (O_1265,N_8368,N_9269);
and UO_1266 (O_1266,N_9131,N_9580);
or UO_1267 (O_1267,N_9224,N_9237);
nand UO_1268 (O_1268,N_9650,N_8804);
or UO_1269 (O_1269,N_9450,N_9649);
and UO_1270 (O_1270,N_9831,N_9172);
nand UO_1271 (O_1271,N_8963,N_8320);
nor UO_1272 (O_1272,N_8590,N_9354);
or UO_1273 (O_1273,N_9606,N_8798);
and UO_1274 (O_1274,N_8614,N_8015);
or UO_1275 (O_1275,N_8737,N_8607);
nor UO_1276 (O_1276,N_8106,N_9339);
and UO_1277 (O_1277,N_9513,N_8803);
nand UO_1278 (O_1278,N_9146,N_9367);
nor UO_1279 (O_1279,N_8893,N_9535);
and UO_1280 (O_1280,N_8729,N_9700);
or UO_1281 (O_1281,N_9604,N_8993);
nor UO_1282 (O_1282,N_9135,N_9366);
nand UO_1283 (O_1283,N_9085,N_9738);
nor UO_1284 (O_1284,N_8413,N_8457);
xnor UO_1285 (O_1285,N_8247,N_8451);
nor UO_1286 (O_1286,N_9730,N_9635);
and UO_1287 (O_1287,N_8346,N_8531);
and UO_1288 (O_1288,N_9818,N_8808);
and UO_1289 (O_1289,N_9751,N_8063);
or UO_1290 (O_1290,N_8318,N_9323);
nand UO_1291 (O_1291,N_8423,N_8354);
or UO_1292 (O_1292,N_8486,N_9021);
nor UO_1293 (O_1293,N_8885,N_8855);
nor UO_1294 (O_1294,N_8211,N_8834);
and UO_1295 (O_1295,N_8142,N_8323);
or UO_1296 (O_1296,N_9004,N_9048);
or UO_1297 (O_1297,N_8141,N_8066);
nor UO_1298 (O_1298,N_8586,N_8516);
or UO_1299 (O_1299,N_8724,N_8322);
and UO_1300 (O_1300,N_9313,N_9088);
and UO_1301 (O_1301,N_9123,N_9810);
and UO_1302 (O_1302,N_8782,N_9330);
and UO_1303 (O_1303,N_8165,N_8522);
and UO_1304 (O_1304,N_8812,N_9995);
and UO_1305 (O_1305,N_9905,N_8364);
nor UO_1306 (O_1306,N_9886,N_9761);
nor UO_1307 (O_1307,N_9865,N_8084);
and UO_1308 (O_1308,N_8982,N_9282);
nor UO_1309 (O_1309,N_9892,N_9522);
xor UO_1310 (O_1310,N_8381,N_8900);
nor UO_1311 (O_1311,N_8117,N_9884);
or UO_1312 (O_1312,N_9943,N_9798);
or UO_1313 (O_1313,N_9341,N_8958);
and UO_1314 (O_1314,N_8110,N_8960);
and UO_1315 (O_1315,N_8957,N_9304);
nor UO_1316 (O_1316,N_9327,N_8550);
nand UO_1317 (O_1317,N_8567,N_8287);
or UO_1318 (O_1318,N_8824,N_8901);
nor UO_1319 (O_1319,N_8625,N_8044);
nand UO_1320 (O_1320,N_9136,N_9622);
or UO_1321 (O_1321,N_8697,N_9629);
and UO_1322 (O_1322,N_9232,N_9512);
nor UO_1323 (O_1323,N_8553,N_9622);
nor UO_1324 (O_1324,N_8717,N_9472);
and UO_1325 (O_1325,N_9653,N_9910);
and UO_1326 (O_1326,N_8501,N_8861);
and UO_1327 (O_1327,N_9500,N_8871);
nand UO_1328 (O_1328,N_9356,N_8940);
nor UO_1329 (O_1329,N_9173,N_8902);
nor UO_1330 (O_1330,N_8156,N_9268);
and UO_1331 (O_1331,N_8088,N_8422);
and UO_1332 (O_1332,N_8207,N_9694);
and UO_1333 (O_1333,N_8641,N_9691);
and UO_1334 (O_1334,N_8765,N_9793);
nor UO_1335 (O_1335,N_8240,N_8741);
or UO_1336 (O_1336,N_8848,N_9193);
nor UO_1337 (O_1337,N_8638,N_9186);
nor UO_1338 (O_1338,N_8117,N_9039);
nand UO_1339 (O_1339,N_8854,N_9858);
nor UO_1340 (O_1340,N_9810,N_9344);
or UO_1341 (O_1341,N_8667,N_8973);
nand UO_1342 (O_1342,N_8192,N_9879);
or UO_1343 (O_1343,N_8129,N_8097);
nand UO_1344 (O_1344,N_8868,N_9989);
nand UO_1345 (O_1345,N_8229,N_8293);
and UO_1346 (O_1346,N_9000,N_8987);
nand UO_1347 (O_1347,N_9654,N_9257);
xnor UO_1348 (O_1348,N_9198,N_9582);
nor UO_1349 (O_1349,N_9769,N_9617);
nand UO_1350 (O_1350,N_9345,N_9034);
or UO_1351 (O_1351,N_9067,N_9285);
nand UO_1352 (O_1352,N_9626,N_9379);
and UO_1353 (O_1353,N_8962,N_9872);
nor UO_1354 (O_1354,N_9595,N_8178);
nand UO_1355 (O_1355,N_8400,N_9004);
or UO_1356 (O_1356,N_8435,N_8081);
or UO_1357 (O_1357,N_9219,N_8741);
nor UO_1358 (O_1358,N_9099,N_9810);
nor UO_1359 (O_1359,N_8088,N_9625);
and UO_1360 (O_1360,N_9282,N_9956);
or UO_1361 (O_1361,N_9277,N_8315);
nand UO_1362 (O_1362,N_9844,N_9612);
nand UO_1363 (O_1363,N_8712,N_9382);
and UO_1364 (O_1364,N_8042,N_9832);
or UO_1365 (O_1365,N_9763,N_8215);
and UO_1366 (O_1366,N_8677,N_9247);
nand UO_1367 (O_1367,N_8670,N_8654);
nand UO_1368 (O_1368,N_8607,N_8926);
and UO_1369 (O_1369,N_9356,N_9909);
nand UO_1370 (O_1370,N_8397,N_9794);
or UO_1371 (O_1371,N_9889,N_8270);
nand UO_1372 (O_1372,N_8148,N_8034);
or UO_1373 (O_1373,N_8028,N_8843);
nand UO_1374 (O_1374,N_8107,N_8847);
nand UO_1375 (O_1375,N_8136,N_9194);
nand UO_1376 (O_1376,N_9541,N_9210);
nor UO_1377 (O_1377,N_9557,N_8597);
nor UO_1378 (O_1378,N_8701,N_9795);
nand UO_1379 (O_1379,N_8454,N_9155);
and UO_1380 (O_1380,N_9557,N_9359);
and UO_1381 (O_1381,N_9492,N_8114);
and UO_1382 (O_1382,N_8874,N_9856);
or UO_1383 (O_1383,N_8442,N_8194);
or UO_1384 (O_1384,N_8709,N_9545);
nor UO_1385 (O_1385,N_9407,N_9459);
xnor UO_1386 (O_1386,N_9304,N_8574);
and UO_1387 (O_1387,N_9778,N_8530);
or UO_1388 (O_1388,N_8766,N_9675);
nand UO_1389 (O_1389,N_8448,N_9657);
nand UO_1390 (O_1390,N_8595,N_9544);
or UO_1391 (O_1391,N_8694,N_8707);
nor UO_1392 (O_1392,N_9123,N_9784);
nand UO_1393 (O_1393,N_8574,N_8908);
or UO_1394 (O_1394,N_9061,N_8374);
xor UO_1395 (O_1395,N_8905,N_9655);
or UO_1396 (O_1396,N_9007,N_9978);
and UO_1397 (O_1397,N_9223,N_9577);
or UO_1398 (O_1398,N_8574,N_9413);
nor UO_1399 (O_1399,N_8659,N_8448);
nand UO_1400 (O_1400,N_9031,N_9775);
nand UO_1401 (O_1401,N_9659,N_8231);
or UO_1402 (O_1402,N_8174,N_8114);
and UO_1403 (O_1403,N_9992,N_8881);
nand UO_1404 (O_1404,N_8056,N_9940);
xor UO_1405 (O_1405,N_9298,N_8961);
xnor UO_1406 (O_1406,N_8682,N_8163);
nor UO_1407 (O_1407,N_9384,N_8563);
and UO_1408 (O_1408,N_9100,N_8993);
or UO_1409 (O_1409,N_8021,N_9760);
or UO_1410 (O_1410,N_9254,N_8767);
and UO_1411 (O_1411,N_8123,N_8130);
and UO_1412 (O_1412,N_8228,N_9943);
or UO_1413 (O_1413,N_8793,N_9474);
nor UO_1414 (O_1414,N_8475,N_9657);
nand UO_1415 (O_1415,N_9728,N_9206);
or UO_1416 (O_1416,N_9379,N_9168);
nand UO_1417 (O_1417,N_8575,N_8606);
nand UO_1418 (O_1418,N_9269,N_8652);
nand UO_1419 (O_1419,N_9055,N_8214);
nand UO_1420 (O_1420,N_9902,N_8187);
nor UO_1421 (O_1421,N_9867,N_8107);
nand UO_1422 (O_1422,N_8135,N_9726);
and UO_1423 (O_1423,N_9752,N_9864);
or UO_1424 (O_1424,N_9427,N_9642);
and UO_1425 (O_1425,N_8780,N_9721);
or UO_1426 (O_1426,N_8032,N_8748);
nand UO_1427 (O_1427,N_8034,N_8026);
or UO_1428 (O_1428,N_9944,N_8952);
nor UO_1429 (O_1429,N_8756,N_8737);
nand UO_1430 (O_1430,N_8827,N_8291);
and UO_1431 (O_1431,N_9446,N_8888);
and UO_1432 (O_1432,N_9956,N_9973);
or UO_1433 (O_1433,N_8324,N_9690);
nor UO_1434 (O_1434,N_9252,N_9511);
and UO_1435 (O_1435,N_8060,N_9007);
nand UO_1436 (O_1436,N_8423,N_9898);
nand UO_1437 (O_1437,N_8870,N_8379);
and UO_1438 (O_1438,N_9033,N_8136);
and UO_1439 (O_1439,N_8890,N_9416);
and UO_1440 (O_1440,N_8876,N_8884);
nor UO_1441 (O_1441,N_9989,N_8323);
and UO_1442 (O_1442,N_9743,N_8416);
nor UO_1443 (O_1443,N_8232,N_9477);
nand UO_1444 (O_1444,N_9430,N_9812);
and UO_1445 (O_1445,N_9418,N_8933);
nor UO_1446 (O_1446,N_8606,N_8487);
nor UO_1447 (O_1447,N_9859,N_9098);
or UO_1448 (O_1448,N_8614,N_9409);
or UO_1449 (O_1449,N_9278,N_9792);
or UO_1450 (O_1450,N_8447,N_9111);
nor UO_1451 (O_1451,N_8943,N_8309);
nand UO_1452 (O_1452,N_8806,N_8077);
or UO_1453 (O_1453,N_8312,N_9379);
nand UO_1454 (O_1454,N_9087,N_8499);
or UO_1455 (O_1455,N_9426,N_9445);
and UO_1456 (O_1456,N_9817,N_8066);
or UO_1457 (O_1457,N_8190,N_8199);
or UO_1458 (O_1458,N_8990,N_8010);
or UO_1459 (O_1459,N_8678,N_8746);
and UO_1460 (O_1460,N_9897,N_8134);
nand UO_1461 (O_1461,N_9235,N_8502);
nand UO_1462 (O_1462,N_9239,N_8574);
and UO_1463 (O_1463,N_9285,N_9029);
or UO_1464 (O_1464,N_9110,N_9152);
or UO_1465 (O_1465,N_9211,N_8485);
nor UO_1466 (O_1466,N_9992,N_8453);
nor UO_1467 (O_1467,N_9148,N_8093);
nor UO_1468 (O_1468,N_8256,N_9497);
and UO_1469 (O_1469,N_8631,N_9065);
nand UO_1470 (O_1470,N_9175,N_8465);
nand UO_1471 (O_1471,N_9199,N_8058);
and UO_1472 (O_1472,N_8470,N_8302);
and UO_1473 (O_1473,N_8125,N_8269);
nand UO_1474 (O_1474,N_8135,N_8852);
nor UO_1475 (O_1475,N_9427,N_8177);
and UO_1476 (O_1476,N_8319,N_9542);
and UO_1477 (O_1477,N_8088,N_9151);
or UO_1478 (O_1478,N_9371,N_8348);
nand UO_1479 (O_1479,N_8005,N_8733);
nor UO_1480 (O_1480,N_9442,N_8685);
or UO_1481 (O_1481,N_8931,N_9480);
nor UO_1482 (O_1482,N_8436,N_9659);
nand UO_1483 (O_1483,N_8966,N_9737);
nand UO_1484 (O_1484,N_8362,N_9259);
nor UO_1485 (O_1485,N_9999,N_8875);
or UO_1486 (O_1486,N_9012,N_8300);
nand UO_1487 (O_1487,N_8082,N_9541);
or UO_1488 (O_1488,N_8034,N_9999);
nor UO_1489 (O_1489,N_9713,N_9568);
nor UO_1490 (O_1490,N_9384,N_9866);
or UO_1491 (O_1491,N_9737,N_8434);
or UO_1492 (O_1492,N_9594,N_9679);
nor UO_1493 (O_1493,N_8672,N_8530);
nor UO_1494 (O_1494,N_9893,N_9553);
or UO_1495 (O_1495,N_8864,N_8346);
or UO_1496 (O_1496,N_9142,N_8675);
or UO_1497 (O_1497,N_8637,N_8455);
nand UO_1498 (O_1498,N_8233,N_8297);
nor UO_1499 (O_1499,N_9461,N_9186);
endmodule