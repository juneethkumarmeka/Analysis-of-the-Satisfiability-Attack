module basic_1000_10000_1500_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_197,In_819);
nand U1 (N_1,In_17,In_973);
or U2 (N_2,In_807,In_225);
nor U3 (N_3,In_558,In_206);
and U4 (N_4,In_897,In_810);
or U5 (N_5,In_813,In_560);
nor U6 (N_6,In_556,In_536);
nor U7 (N_7,In_296,In_626);
or U8 (N_8,In_471,In_417);
or U9 (N_9,In_55,In_373);
or U10 (N_10,In_306,In_575);
xnor U11 (N_11,In_227,In_261);
and U12 (N_12,In_912,In_426);
and U13 (N_13,In_133,In_984);
nor U14 (N_14,In_634,In_397);
or U15 (N_15,In_765,In_484);
or U16 (N_16,In_169,In_120);
and U17 (N_17,In_616,In_95);
nor U18 (N_18,In_787,In_809);
nor U19 (N_19,In_13,In_563);
and U20 (N_20,In_972,In_326);
xor U21 (N_21,In_140,In_670);
and U22 (N_22,In_685,In_486);
and U23 (N_23,In_806,In_996);
nor U24 (N_24,In_91,In_549);
or U25 (N_25,In_262,In_396);
nand U26 (N_26,In_528,In_938);
nor U27 (N_27,In_249,In_155);
and U28 (N_28,In_950,In_219);
or U29 (N_29,In_242,In_450);
nand U30 (N_30,In_156,In_998);
nor U31 (N_31,In_708,In_791);
and U32 (N_32,In_257,In_435);
nand U33 (N_33,In_707,In_901);
nand U34 (N_34,In_237,In_508);
nor U35 (N_35,In_478,In_105);
xnor U36 (N_36,In_14,In_11);
or U37 (N_37,In_775,In_762);
or U38 (N_38,In_644,In_183);
and U39 (N_39,In_48,In_758);
and U40 (N_40,In_504,In_266);
or U41 (N_41,In_684,In_121);
nor U42 (N_42,In_908,In_401);
nand U43 (N_43,In_128,In_20);
or U44 (N_44,In_94,In_369);
nor U45 (N_45,In_691,In_49);
nor U46 (N_46,In_655,In_36);
nand U47 (N_47,In_904,In_232);
nand U48 (N_48,In_959,In_291);
and U49 (N_49,In_304,In_951);
nand U50 (N_50,In_454,In_805);
or U51 (N_51,In_713,In_365);
and U52 (N_52,In_35,In_717);
nand U53 (N_53,In_190,In_917);
and U54 (N_54,In_970,In_579);
nor U55 (N_55,In_916,In_308);
or U56 (N_56,In_492,In_376);
xnor U57 (N_57,In_537,In_16);
and U58 (N_58,In_940,In_289);
nor U59 (N_59,In_413,In_994);
xor U60 (N_60,In_424,In_759);
nor U61 (N_61,In_876,In_661);
nor U62 (N_62,In_463,In_464);
or U63 (N_63,In_301,In_406);
nor U64 (N_64,In_638,In_542);
and U65 (N_65,In_459,In_148);
and U66 (N_66,In_506,In_989);
or U67 (N_67,In_297,In_774);
or U68 (N_68,In_46,In_112);
and U69 (N_69,In_28,In_754);
and U70 (N_70,In_960,In_336);
or U71 (N_71,In_719,In_602);
nand U72 (N_72,In_766,In_735);
or U73 (N_73,In_161,In_773);
and U74 (N_74,In_519,In_514);
and U75 (N_75,In_677,In_597);
xnor U76 (N_76,In_33,In_134);
nor U77 (N_77,In_172,In_864);
or U78 (N_78,In_390,In_927);
xor U79 (N_79,In_247,In_393);
xnor U80 (N_80,In_381,In_321);
nor U81 (N_81,In_830,In_207);
nor U82 (N_82,In_419,In_932);
nand U83 (N_83,In_353,In_144);
and U84 (N_84,In_117,In_250);
and U85 (N_85,In_694,In_838);
xor U86 (N_86,In_693,In_298);
or U87 (N_87,In_467,In_865);
xor U88 (N_88,In_573,In_106);
xor U89 (N_89,In_841,In_578);
or U90 (N_90,In_84,In_890);
or U91 (N_91,In_267,In_153);
nand U92 (N_92,In_955,In_609);
or U93 (N_93,In_38,In_588);
and U94 (N_94,In_939,In_92);
nand U95 (N_95,In_907,In_361);
and U96 (N_96,In_294,In_354);
and U97 (N_97,In_44,In_629);
nand U98 (N_98,In_898,In_997);
and U99 (N_99,In_166,In_313);
nand U100 (N_100,In_392,In_154);
and U101 (N_101,In_667,In_742);
nor U102 (N_102,In_359,In_391);
xnor U103 (N_103,In_697,In_276);
xor U104 (N_104,In_186,In_10);
or U105 (N_105,In_615,In_711);
nand U106 (N_106,In_213,In_619);
nand U107 (N_107,In_233,In_348);
nand U108 (N_108,In_601,In_62);
xor U109 (N_109,In_650,In_505);
nor U110 (N_110,In_83,In_906);
or U111 (N_111,In_462,In_768);
or U112 (N_112,In_705,In_600);
and U113 (N_113,In_681,In_926);
nor U114 (N_114,In_891,In_198);
xor U115 (N_115,In_309,In_420);
and U116 (N_116,In_503,In_56);
nor U117 (N_117,In_696,In_745);
nor U118 (N_118,In_975,In_531);
nor U119 (N_119,In_256,In_944);
or U120 (N_120,In_200,In_613);
or U121 (N_121,In_310,In_714);
or U122 (N_122,In_223,In_568);
xor U123 (N_123,In_164,In_974);
nand U124 (N_124,In_721,In_914);
xnor U125 (N_125,In_637,In_682);
nand U126 (N_126,In_272,In_577);
xor U127 (N_127,In_239,In_130);
or U128 (N_128,In_982,In_852);
nor U129 (N_129,In_870,In_957);
xnor U130 (N_130,In_849,In_332);
or U131 (N_131,In_138,In_100);
and U132 (N_132,In_31,In_176);
xor U133 (N_133,In_189,In_544);
or U134 (N_134,In_980,In_243);
and U135 (N_135,In_19,In_933);
xor U136 (N_136,In_45,In_781);
and U137 (N_137,In_652,In_518);
nor U138 (N_138,In_442,In_330);
nor U139 (N_139,In_47,In_888);
and U140 (N_140,In_69,In_386);
and U141 (N_141,In_760,In_611);
nand U142 (N_142,In_533,In_541);
xor U143 (N_143,In_590,In_937);
nand U144 (N_144,In_653,In_458);
and U145 (N_145,In_312,In_792);
nor U146 (N_146,In_226,In_152);
nor U147 (N_147,In_210,In_222);
nor U148 (N_148,In_837,In_999);
nand U149 (N_149,In_594,In_827);
or U150 (N_150,In_202,In_779);
xor U151 (N_151,In_18,In_340);
and U152 (N_152,In_674,In_523);
nor U153 (N_153,In_798,In_598);
nand U154 (N_154,In_96,In_546);
and U155 (N_155,In_220,In_561);
nand U156 (N_156,In_911,In_77);
and U157 (N_157,In_345,In_388);
nand U158 (N_158,In_65,In_816);
nor U159 (N_159,In_270,In_292);
nand U160 (N_160,In_80,In_265);
or U161 (N_161,In_969,In_203);
and U162 (N_162,In_315,In_79);
xnor U163 (N_163,In_281,In_803);
xnor U164 (N_164,In_800,In_151);
xnor U165 (N_165,In_868,In_633);
xor U166 (N_166,In_886,In_763);
nor U167 (N_167,In_251,In_165);
nand U168 (N_168,In_127,In_322);
nand U169 (N_169,In_67,In_562);
xnor U170 (N_170,In_498,In_517);
xor U171 (N_171,In_452,In_509);
nor U172 (N_172,In_483,In_961);
xor U173 (N_173,In_286,In_212);
nand U174 (N_174,In_41,In_481);
nand U175 (N_175,In_820,In_358);
nor U176 (N_176,In_608,In_116);
and U177 (N_177,In_490,In_143);
nand U178 (N_178,In_446,In_173);
and U179 (N_179,In_967,In_107);
xor U180 (N_180,In_74,In_698);
and U181 (N_181,In_612,In_636);
and U182 (N_182,In_122,In_734);
nor U183 (N_183,In_377,In_844);
and U184 (N_184,In_229,In_668);
nor U185 (N_185,In_741,In_953);
or U186 (N_186,In_535,In_241);
or U187 (N_187,In_187,In_945);
nand U188 (N_188,In_649,In_25);
nor U189 (N_189,In_701,In_570);
xor U190 (N_190,In_709,In_526);
and U191 (N_191,In_630,In_82);
nand U192 (N_192,In_761,In_753);
nor U193 (N_193,In_769,In_954);
nand U194 (N_194,In_522,In_331);
nand U195 (N_195,In_441,In_167);
xor U196 (N_196,In_995,In_565);
xnor U197 (N_197,In_287,In_293);
or U198 (N_198,In_328,In_473);
or U199 (N_199,In_314,In_727);
or U200 (N_200,In_716,N_51);
nand U201 (N_201,N_189,In_875);
xnor U202 (N_202,In_862,N_1);
nand U203 (N_203,In_40,In_137);
nand U204 (N_204,N_191,In_675);
xor U205 (N_205,In_97,In_706);
nand U206 (N_206,In_60,N_11);
nor U207 (N_207,In_409,In_737);
nor U208 (N_208,In_295,N_163);
nor U209 (N_209,N_88,N_131);
xor U210 (N_210,N_5,In_181);
and U211 (N_211,N_152,In_382);
nand U212 (N_212,In_909,N_4);
or U213 (N_213,N_42,N_80);
or U214 (N_214,In_363,N_43);
xor U215 (N_215,In_543,N_183);
or U216 (N_216,In_510,In_379);
nand U217 (N_217,In_723,In_260);
nor U218 (N_218,In_280,In_125);
and U219 (N_219,In_660,In_855);
or U220 (N_220,In_624,N_181);
nand U221 (N_221,In_924,N_54);
or U222 (N_222,N_56,In_255);
nor U223 (N_223,N_33,In_866);
and U224 (N_224,N_168,In_513);
or U225 (N_225,N_153,N_39);
and U226 (N_226,In_86,In_248);
and U227 (N_227,N_145,N_197);
or U228 (N_228,In_412,N_2);
or U229 (N_229,In_440,In_443);
xnor U230 (N_230,N_85,In_421);
and U231 (N_231,In_288,N_100);
xnor U232 (N_232,In_114,N_63);
nand U233 (N_233,In_700,In_78);
or U234 (N_234,In_163,In_796);
nand U235 (N_235,In_337,In_869);
and U236 (N_236,In_240,In_274);
or U237 (N_237,In_867,In_718);
and U238 (N_238,In_34,N_90);
and U239 (N_239,In_87,N_57);
and U240 (N_240,In_666,In_979);
and U241 (N_241,N_77,N_115);
nand U242 (N_242,N_140,In_99);
nor U243 (N_243,In_593,In_271);
or U244 (N_244,In_715,In_686);
or U245 (N_245,In_739,In_234);
xnor U246 (N_246,In_783,N_93);
nand U247 (N_247,In_177,In_436);
nor U248 (N_248,In_461,N_65);
nand U249 (N_249,N_109,In_736);
nor U250 (N_250,In_930,N_47);
nor U251 (N_251,In_214,In_591);
xor U252 (N_252,In_669,N_172);
xnor U253 (N_253,In_576,In_671);
xor U254 (N_254,In_218,In_437);
or U255 (N_255,N_38,In_339);
nor U256 (N_256,In_992,In_958);
xnor U257 (N_257,In_977,In_456);
or U258 (N_258,N_104,N_134);
or U259 (N_259,In_710,N_147);
nor U260 (N_260,In_521,In_703);
xnor U261 (N_261,In_224,In_731);
nand U262 (N_262,In_102,In_320);
xor U263 (N_263,In_622,In_662);
nor U264 (N_264,N_97,In_264);
nand U265 (N_265,In_746,N_170);
xor U266 (N_266,N_173,N_184);
or U267 (N_267,In_1,N_138);
or U268 (N_268,In_515,In_672);
xnor U269 (N_269,In_191,In_948);
or U270 (N_270,In_673,In_434);
xnor U271 (N_271,In_607,In_351);
xnor U272 (N_272,In_548,In_496);
xnor U273 (N_273,N_108,In_29);
nand U274 (N_274,In_439,N_67);
nor U275 (N_275,In_453,In_427);
or U276 (N_276,In_51,In_174);
xnor U277 (N_277,In_882,In_679);
nand U278 (N_278,In_4,N_185);
nand U279 (N_279,In_688,In_825);
xnor U280 (N_280,In_178,In_894);
xor U281 (N_281,N_17,In_665);
nor U282 (N_282,In_433,In_7);
xor U283 (N_283,In_73,N_154);
and U284 (N_284,N_157,In_21);
nand U285 (N_285,In_495,N_110);
or U286 (N_286,In_569,N_177);
nand U287 (N_287,In_976,In_129);
xor U288 (N_288,N_81,N_141);
nor U289 (N_289,N_64,In_755);
xor U290 (N_290,In_93,In_683);
or U291 (N_291,In_511,In_729);
and U292 (N_292,N_52,In_194);
xor U293 (N_293,N_20,In_552);
xor U294 (N_294,N_139,N_10);
or U295 (N_295,In_325,In_863);
xor U296 (N_296,In_524,In_687);
nand U297 (N_297,In_764,In_851);
nor U298 (N_298,In_702,In_952);
xnor U299 (N_299,N_123,In_853);
xnor U300 (N_300,N_50,In_324);
nand U301 (N_301,In_482,In_804);
nand U302 (N_302,In_278,N_129);
nor U303 (N_303,In_889,In_394);
and U304 (N_304,In_534,N_144);
and U305 (N_305,In_50,In_857);
and U306 (N_306,In_494,In_491);
or U307 (N_307,In_457,In_277);
nand U308 (N_308,In_66,In_68);
nor U309 (N_309,N_92,In_547);
or U310 (N_310,In_192,In_586);
and U311 (N_311,In_162,In_146);
xnor U312 (N_312,In_712,In_928);
or U313 (N_313,In_445,In_258);
nand U314 (N_314,In_822,In_583);
and U315 (N_315,N_142,In_808);
xor U316 (N_316,In_70,In_829);
nand U317 (N_317,N_37,In_53);
nor U318 (N_318,In_170,In_317);
and U319 (N_319,N_136,N_98);
nand U320 (N_320,N_73,In_216);
xnor U321 (N_321,In_404,In_357);
or U322 (N_322,N_6,In_585);
or U323 (N_323,N_117,N_13);
nand U324 (N_324,In_362,In_283);
or U325 (N_325,In_854,In_244);
or U326 (N_326,N_112,In_168);
nor U327 (N_327,N_3,In_338);
or U328 (N_328,In_777,In_299);
nand U329 (N_329,In_582,N_84);
xnor U330 (N_330,In_799,In_329);
nor U331 (N_331,In_346,In_182);
xnor U332 (N_332,In_113,In_370);
xnor U333 (N_333,N_68,In_316);
xor U334 (N_334,In_303,N_195);
xnor U335 (N_335,In_567,In_185);
and U336 (N_336,In_311,In_188);
nand U337 (N_337,N_126,In_126);
and U338 (N_338,N_31,In_57);
nor U339 (N_339,In_39,In_581);
or U340 (N_340,N_35,In_52);
xor U341 (N_341,In_387,In_756);
or U342 (N_342,In_628,In_770);
nand U343 (N_343,In_551,In_968);
and U344 (N_344,In_416,In_899);
and U345 (N_345,In_689,N_27);
nand U346 (N_346,In_195,In_918);
and U347 (N_347,In_26,In_596);
or U348 (N_348,In_343,In_877);
and U349 (N_349,N_187,N_127);
nand U350 (N_350,In_217,N_199);
or U351 (N_351,N_94,In_946);
nand U352 (N_352,In_923,N_78);
and U353 (N_353,N_32,In_589);
and U354 (N_354,In_902,In_411);
or U355 (N_355,In_493,In_54);
and U356 (N_356,In_269,In_385);
and U357 (N_357,In_142,In_858);
nor U358 (N_358,In_395,In_695);
nor U359 (N_359,In_318,In_448);
xnor U360 (N_360,N_96,In_840);
nor U361 (N_361,In_784,In_733);
nor U362 (N_362,In_43,In_801);
nand U363 (N_363,N_107,N_192);
xnor U364 (N_364,In_32,In_103);
or U365 (N_365,N_91,In_610);
or U366 (N_366,In_978,In_432);
or U367 (N_367,In_835,In_451);
and U368 (N_368,In_988,In_566);
and U369 (N_369,In_418,N_16);
xnor U370 (N_370,N_101,In_231);
xor U371 (N_371,In_527,In_360);
nor U372 (N_372,In_159,In_815);
and U373 (N_373,N_158,N_188);
nand U374 (N_374,N_75,In_180);
and U375 (N_375,In_5,In_149);
and U376 (N_376,N_86,In_89);
or U377 (N_377,In_993,In_651);
or U378 (N_378,N_89,N_114);
or U379 (N_379,In_850,In_476);
xor U380 (N_380,In_884,In_344);
nand U381 (N_381,In_380,In_726);
or U382 (N_382,In_678,In_228);
and U383 (N_383,In_500,N_14);
xnor U384 (N_384,In_966,In_640);
xnor U385 (N_385,In_512,In_132);
or U386 (N_386,In_557,In_290);
xor U387 (N_387,In_776,In_211);
nand U388 (N_388,In_620,N_180);
xor U389 (N_389,N_133,In_215);
nor U390 (N_390,In_874,In_399);
or U391 (N_391,In_410,In_872);
nand U392 (N_392,In_895,In_880);
nand U393 (N_393,In_184,In_72);
nand U394 (N_394,In_9,In_635);
nor U395 (N_395,In_883,N_149);
and U396 (N_396,In_525,In_971);
or U397 (N_397,In_141,In_732);
nand U398 (N_398,In_253,N_116);
and U399 (N_399,In_352,N_171);
or U400 (N_400,In_929,N_294);
and U401 (N_401,N_23,In_507);
or U402 (N_402,In_375,N_291);
nor U403 (N_403,N_255,N_210);
nand U404 (N_404,N_318,In_414);
nand U405 (N_405,N_62,N_241);
xnor U406 (N_406,In_477,In_323);
or U407 (N_407,N_128,In_400);
nor U408 (N_408,N_346,N_382);
xor U409 (N_409,N_132,N_275);
xnor U410 (N_410,In_757,N_317);
xnor U411 (N_411,N_366,N_311);
nor U412 (N_412,N_70,In_108);
xnor U413 (N_413,N_253,N_329);
xor U414 (N_414,In_540,In_539);
nor U415 (N_415,In_587,N_214);
nor U416 (N_416,N_356,In_845);
and U417 (N_417,N_113,N_8);
nand U418 (N_418,N_246,In_364);
or U419 (N_419,N_338,N_324);
xnor U420 (N_420,In_423,N_234);
or U421 (N_421,In_722,In_744);
nor U422 (N_422,N_319,In_300);
xnor U423 (N_423,In_209,N_66);
and U424 (N_424,N_146,In_199);
nor U425 (N_425,In_572,N_244);
or U426 (N_426,N_371,N_217);
or U427 (N_427,In_887,N_309);
and U428 (N_428,N_186,In_470);
or U429 (N_429,In_748,In_111);
or U430 (N_430,N_190,In_554);
nor U431 (N_431,In_109,In_663);
nor U432 (N_432,In_124,In_942);
or U433 (N_433,N_335,N_326);
and U434 (N_434,N_207,N_135);
xor U435 (N_435,In_555,N_340);
and U436 (N_436,N_383,N_240);
and U437 (N_437,N_82,In_821);
xor U438 (N_438,In_574,N_299);
nand U439 (N_439,N_386,In_931);
nand U440 (N_440,N_222,N_231);
xnor U441 (N_441,N_350,In_368);
xor U442 (N_442,In_614,N_21);
nor U443 (N_443,N_369,N_229);
nor U444 (N_444,In_750,N_296);
xor U445 (N_445,N_44,N_365);
nor U446 (N_446,N_59,In_502);
nor U447 (N_447,N_102,In_430);
xor U448 (N_448,N_304,N_26);
nand U449 (N_449,N_363,N_205);
or U450 (N_450,In_991,N_200);
nor U451 (N_451,In_811,N_219);
xor U452 (N_452,N_242,N_247);
nor U453 (N_453,In_425,In_963);
or U454 (N_454,In_135,N_36);
or U455 (N_455,N_374,N_119);
and U456 (N_456,In_794,In_468);
nand U457 (N_457,In_472,N_150);
nand U458 (N_458,N_353,N_28);
or U459 (N_459,N_155,In_145);
and U460 (N_460,N_69,In_843);
xnor U461 (N_461,In_802,N_22);
and U462 (N_462,N_159,In_657);
and U463 (N_463,In_341,N_358);
xor U464 (N_464,In_488,In_366);
nor U465 (N_465,In_664,N_357);
nand U466 (N_466,In_529,In_499);
and U467 (N_467,In_355,In_842);
xor U468 (N_468,In_63,N_164);
xor U469 (N_469,N_372,N_233);
and U470 (N_470,N_212,In_371);
and U471 (N_471,In_422,N_121);
and U472 (N_472,In_403,In_915);
nor U473 (N_473,In_384,N_314);
and U474 (N_474,In_981,N_213);
nand U475 (N_475,In_680,In_230);
and U476 (N_476,N_307,N_352);
nand U477 (N_477,In_449,N_194);
or U478 (N_478,In_305,N_72);
nor U479 (N_479,In_647,In_632);
nand U480 (N_480,In_848,N_333);
nor U481 (N_481,N_273,N_364);
nor U482 (N_482,N_316,N_283);
xor U483 (N_483,In_538,In_150);
nand U484 (N_484,N_373,In_618);
or U485 (N_485,In_469,N_169);
and U486 (N_486,In_642,In_790);
and U487 (N_487,In_943,N_193);
nand U488 (N_488,N_156,N_396);
nand U489 (N_489,N_292,In_160);
or U490 (N_490,In_221,N_223);
nand U491 (N_491,N_111,N_249);
nor U492 (N_492,In_778,In_913);
nor U493 (N_493,N_285,N_351);
and U494 (N_494,In_859,N_315);
nand U495 (N_495,In_347,In_625);
nor U496 (N_496,N_201,N_279);
nand U497 (N_497,N_248,N_120);
nand U498 (N_498,N_376,In_627);
and U499 (N_499,In_372,N_293);
and U500 (N_500,N_243,In_98);
nor U501 (N_501,N_397,In_740);
xor U502 (N_502,N_198,In_3);
or U503 (N_503,In_428,In_545);
nor U504 (N_504,N_289,N_160);
xnor U505 (N_505,In_88,In_30);
nand U506 (N_506,In_646,N_263);
and U507 (N_507,N_343,N_348);
nor U508 (N_508,In_592,N_384);
and U509 (N_509,N_337,In_6);
and U510 (N_510,In_720,In_879);
nand U511 (N_511,In_751,N_302);
nand U512 (N_512,N_208,N_272);
or U513 (N_513,In_893,In_648);
nor U514 (N_514,N_40,In_447);
or U515 (N_515,In_692,In_302);
or U516 (N_516,In_90,In_860);
nor U517 (N_517,In_730,In_438);
or U518 (N_518,In_823,In_782);
xor U519 (N_519,In_24,In_839);
xnor U520 (N_520,In_724,In_263);
nand U521 (N_521,In_964,N_182);
nand U522 (N_522,N_381,N_295);
and U523 (N_523,N_345,In_936);
xnor U524 (N_524,N_261,In_772);
or U525 (N_525,In_171,N_395);
and U526 (N_526,In_475,In_606);
or U527 (N_527,In_236,In_747);
xor U528 (N_528,N_71,N_29);
or U529 (N_529,In_641,In_881);
and U530 (N_530,In_817,N_323);
nand U531 (N_531,In_282,N_280);
xnor U532 (N_532,In_76,N_325);
nor U533 (N_533,In_789,In_603);
and U534 (N_534,In_812,N_230);
and U535 (N_535,In_402,In_530);
nand U536 (N_536,In_101,N_0);
or U537 (N_537,In_749,N_380);
and U538 (N_538,In_595,N_377);
or U539 (N_539,N_306,N_360);
nor U540 (N_540,In_407,In_487);
or U541 (N_541,In_175,In_356);
nand U542 (N_542,In_834,N_178);
xor U543 (N_543,In_408,N_130);
nor U544 (N_544,In_64,N_179);
or U545 (N_545,In_949,N_105);
nand U546 (N_546,N_122,In_350);
nand U547 (N_547,In_623,In_268);
and U548 (N_548,In_157,N_103);
nor U549 (N_549,In_983,In_444);
or U550 (N_550,N_174,In_516);
nand U551 (N_551,N_305,In_246);
nand U552 (N_552,N_176,In_905);
and U553 (N_553,N_19,In_205);
or U554 (N_554,N_79,In_824);
nand U555 (N_555,N_9,In_921);
xnor U556 (N_556,In_847,In_245);
nor U557 (N_557,N_46,N_166);
and U558 (N_558,N_48,In_690);
nor U559 (N_559,N_278,In_643);
or U560 (N_560,In_429,N_399);
xor U561 (N_561,N_61,In_571);
nand U562 (N_562,N_308,N_303);
nand U563 (N_563,In_8,In_676);
and U564 (N_564,N_209,In_285);
nor U565 (N_565,N_55,N_288);
nor U566 (N_566,N_298,N_12);
nand U567 (N_567,In_728,N_388);
xnor U568 (N_568,In_460,N_124);
xnor U569 (N_569,N_167,In_910);
nand U570 (N_570,N_252,In_147);
nor U571 (N_571,In_956,In_501);
nand U572 (N_572,N_251,In_335);
xnor U573 (N_573,N_264,N_218);
xnor U574 (N_574,N_60,N_290);
and U575 (N_575,In_238,In_920);
nand U576 (N_576,In_617,In_605);
or U577 (N_577,N_53,In_333);
nand U578 (N_578,In_474,In_743);
or U579 (N_579,In_136,N_257);
nor U580 (N_580,In_639,In_658);
nor U581 (N_581,N_321,In_903);
nand U582 (N_582,N_312,In_179);
or U583 (N_583,N_281,In_832);
and U584 (N_584,N_320,N_270);
nand U585 (N_585,In_235,In_104);
xor U586 (N_586,N_245,N_239);
nor U587 (N_587,N_58,In_59);
nor U588 (N_588,In_725,In_962);
xor U589 (N_589,N_331,N_328);
nor U590 (N_590,N_297,In_23);
nand U591 (N_591,N_225,In_327);
nor U592 (N_592,N_259,In_656);
or U593 (N_593,N_392,In_374);
xnor U594 (N_594,In_654,In_621);
xor U595 (N_595,N_224,N_250);
nor U596 (N_596,In_785,N_389);
and U597 (N_597,N_74,In_61);
or U598 (N_598,In_123,In_389);
xnor U599 (N_599,N_260,N_375);
and U600 (N_600,In_85,In_873);
xnor U601 (N_601,N_524,N_83);
xor U602 (N_602,N_284,N_596);
nand U603 (N_603,In_532,N_416);
nor U604 (N_604,In_405,In_196);
nand U605 (N_605,N_445,N_532);
xor U606 (N_606,N_453,N_393);
xor U607 (N_607,N_349,N_417);
xor U608 (N_608,N_444,N_519);
nand U609 (N_609,N_547,In_2);
and U610 (N_610,In_71,N_162);
xnor U611 (N_611,In_415,N_428);
xor U612 (N_612,In_941,In_631);
and U613 (N_613,N_265,N_443);
and U614 (N_614,N_588,N_587);
nand U615 (N_615,N_221,N_277);
xnor U616 (N_616,In_378,In_900);
xor U617 (N_617,N_282,N_354);
or U618 (N_618,N_555,N_462);
and U619 (N_619,In_780,N_483);
nand U620 (N_620,In_0,N_505);
xnor U621 (N_621,In_252,N_568);
xor U622 (N_622,N_549,In_833);
xor U623 (N_623,N_472,N_347);
xor U624 (N_624,N_495,N_24);
nand U625 (N_625,N_237,In_828);
xor U626 (N_626,N_535,In_986);
and U627 (N_627,In_398,N_466);
xnor U628 (N_628,N_529,N_408);
nor U629 (N_629,N_414,N_514);
nor U630 (N_630,In_580,In_208);
nand U631 (N_631,N_513,N_301);
and U632 (N_632,N_531,N_512);
and U633 (N_633,N_579,N_421);
or U634 (N_634,N_342,N_287);
or U635 (N_635,N_359,N_438);
or U636 (N_636,N_566,N_562);
and U637 (N_637,N_500,In_520);
xor U638 (N_638,N_266,N_477);
and U639 (N_639,N_534,N_409);
xnor U640 (N_640,N_268,N_591);
nor U641 (N_641,N_508,In_793);
and U642 (N_642,N_143,In_831);
nand U643 (N_643,N_576,N_578);
nand U644 (N_644,In_131,In_752);
and U645 (N_645,In_885,In_158);
nand U646 (N_646,N_228,N_523);
nor U647 (N_647,In_81,N_589);
nand U648 (N_648,N_449,N_402);
or U649 (N_649,N_330,N_406);
nor U650 (N_650,N_457,N_378);
xor U651 (N_651,N_528,In_896);
nor U652 (N_652,N_470,In_479);
and U653 (N_653,N_425,In_836);
nor U654 (N_654,N_537,N_30);
nand U655 (N_655,In_115,N_341);
or U656 (N_656,N_25,In_273);
xor U657 (N_657,N_593,N_211);
and U658 (N_658,In_466,N_429);
or U659 (N_659,N_411,In_925);
nand U660 (N_660,N_484,In_27);
xor U661 (N_661,In_110,N_427);
xnor U662 (N_662,N_256,N_434);
or U663 (N_663,N_398,N_262);
nand U664 (N_664,N_583,N_405);
nor U665 (N_665,N_570,N_269);
or U666 (N_666,In_489,N_517);
nand U667 (N_667,N_452,N_95);
nor U668 (N_668,In_818,In_15);
nand U669 (N_669,N_548,In_139);
xor U670 (N_670,In_659,N_594);
and U671 (N_671,In_704,N_271);
nand U672 (N_672,N_538,N_595);
or U673 (N_673,N_454,N_276);
or U674 (N_674,In_383,In_553);
xnor U675 (N_675,N_254,N_530);
nand U676 (N_676,In_279,N_367);
nor U677 (N_677,In_934,N_286);
and U678 (N_678,N_327,N_451);
and U679 (N_679,N_45,N_522);
or U680 (N_680,In_645,N_76);
nand U681 (N_681,N_564,N_571);
or U682 (N_682,In_604,N_99);
or U683 (N_683,N_545,N_161);
nand U684 (N_684,N_412,N_520);
and U685 (N_685,N_361,N_533);
nand U686 (N_686,N_420,N_471);
nor U687 (N_687,N_202,N_336);
or U688 (N_688,N_165,N_226);
nand U689 (N_689,N_459,N_580);
and U690 (N_690,N_274,N_446);
nor U691 (N_691,N_464,N_450);
nand U692 (N_692,N_498,N_322);
xnor U693 (N_693,N_423,In_795);
nand U694 (N_694,N_511,N_232);
or U695 (N_695,N_502,In_797);
xor U696 (N_696,N_41,N_267);
and U697 (N_697,In_254,N_490);
nand U698 (N_698,N_592,N_572);
and U699 (N_699,N_18,N_461);
nor U700 (N_700,N_597,N_488);
and U701 (N_701,N_540,N_518);
xnor U702 (N_702,N_404,N_447);
xnor U703 (N_703,In_342,In_485);
nor U704 (N_704,In_935,N_491);
xor U705 (N_705,N_137,In_947);
and U706 (N_706,In_856,In_892);
nand U707 (N_707,N_506,In_767);
nand U708 (N_708,N_49,In_284);
nor U709 (N_709,N_216,N_458);
nand U710 (N_710,In_990,N_148);
or U711 (N_711,In_985,N_34);
or U712 (N_712,N_493,In_550);
nor U713 (N_713,N_344,N_504);
nand U714 (N_714,N_516,N_440);
nor U715 (N_715,N_487,N_439);
or U716 (N_716,N_332,N_455);
or U717 (N_717,N_536,N_478);
nor U718 (N_718,In_58,N_485);
and U719 (N_719,In_559,In_599);
and U720 (N_720,N_196,N_424);
and U721 (N_721,N_480,N_559);
nor U722 (N_722,N_118,N_460);
and U723 (N_723,N_550,N_565);
nor U724 (N_724,N_563,N_390);
and U725 (N_725,In_334,N_473);
and U726 (N_726,N_476,In_193);
nand U727 (N_727,N_481,N_313);
xnor U728 (N_728,N_574,N_501);
and U729 (N_729,N_391,N_407);
xnor U730 (N_730,N_557,N_539);
xnor U731 (N_731,In_204,In_431);
xnor U732 (N_732,N_551,N_15);
nor U733 (N_733,N_401,N_258);
or U734 (N_734,N_236,N_598);
or U735 (N_735,In_846,N_599);
and U736 (N_736,N_525,N_475);
xor U737 (N_737,N_300,N_560);
or U738 (N_738,N_507,N_499);
nor U739 (N_739,N_552,In_814);
or U740 (N_740,N_486,N_422);
and U741 (N_741,N_482,N_415);
xnor U742 (N_742,In_367,N_400);
or U743 (N_743,In_75,N_432);
and U744 (N_744,N_235,In_119);
and U745 (N_745,N_556,In_42);
or U746 (N_746,N_585,N_220);
and U747 (N_747,N_503,In_987);
nor U748 (N_748,In_22,N_586);
xor U749 (N_749,N_419,N_125);
and U750 (N_750,N_437,N_526);
or U751 (N_751,N_418,In_699);
nor U752 (N_752,N_569,In_771);
and U753 (N_753,N_510,N_515);
nor U754 (N_754,N_543,N_496);
nor U755 (N_755,N_203,N_334);
xor U756 (N_756,N_87,N_410);
nand U757 (N_757,N_238,N_413);
nor U758 (N_758,N_456,N_573);
and U759 (N_759,In_349,N_541);
nor U760 (N_760,In_259,N_441);
xnor U761 (N_761,N_215,In_307);
nand U762 (N_762,N_431,N_435);
and U763 (N_763,In_201,N_465);
xor U764 (N_764,In_319,N_468);
nand U765 (N_765,N_584,N_433);
nor U766 (N_766,N_509,In_275);
and U767 (N_767,N_436,N_567);
or U768 (N_768,N_497,N_542);
xnor U769 (N_769,In_564,In_922);
or U770 (N_770,N_492,In_871);
nand U771 (N_771,In_786,N_394);
nand U772 (N_772,N_442,N_430);
nand U773 (N_773,N_175,N_581);
nor U774 (N_774,N_387,In_738);
xor U775 (N_775,In_584,N_553);
and U776 (N_776,N_467,N_561);
and U777 (N_777,In_919,N_227);
xnor U778 (N_778,N_403,N_474);
and U779 (N_779,N_544,N_521);
or U780 (N_780,N_362,N_355);
and U781 (N_781,In_480,N_379);
nand U782 (N_782,N_479,In_118);
nor U783 (N_783,N_106,N_577);
nand U784 (N_784,N_339,In_861);
nor U785 (N_785,N_558,N_448);
nor U786 (N_786,In_465,N_489);
xor U787 (N_787,In_878,N_310);
nor U788 (N_788,N_546,N_206);
nand U789 (N_789,In_12,N_370);
nand U790 (N_790,In_788,In_965);
nor U791 (N_791,N_385,N_469);
and U792 (N_792,In_497,N_554);
and U793 (N_793,N_7,N_151);
nor U794 (N_794,N_527,N_582);
or U795 (N_795,In_455,In_37);
nand U796 (N_796,N_368,N_590);
nand U797 (N_797,N_426,In_826);
xnor U798 (N_798,N_463,N_494);
nand U799 (N_799,N_575,N_204);
nor U800 (N_800,N_663,N_668);
xnor U801 (N_801,N_722,N_703);
nand U802 (N_802,N_607,N_677);
nand U803 (N_803,N_613,N_636);
nand U804 (N_804,N_610,N_725);
nand U805 (N_805,N_767,N_716);
and U806 (N_806,N_752,N_742);
and U807 (N_807,N_642,N_632);
or U808 (N_808,N_760,N_713);
nor U809 (N_809,N_667,N_705);
xor U810 (N_810,N_675,N_627);
nor U811 (N_811,N_624,N_690);
nor U812 (N_812,N_738,N_774);
xnor U813 (N_813,N_604,N_741);
nor U814 (N_814,N_676,N_683);
nor U815 (N_815,N_631,N_794);
xor U816 (N_816,N_798,N_757);
and U817 (N_817,N_630,N_748);
xor U818 (N_818,N_720,N_765);
nor U819 (N_819,N_626,N_608);
nand U820 (N_820,N_645,N_773);
and U821 (N_821,N_664,N_617);
xnor U822 (N_822,N_777,N_646);
or U823 (N_823,N_669,N_731);
nand U824 (N_824,N_761,N_644);
or U825 (N_825,N_749,N_739);
xnor U826 (N_826,N_605,N_737);
nor U827 (N_827,N_660,N_651);
nor U828 (N_828,N_601,N_784);
xnor U829 (N_829,N_671,N_785);
nand U830 (N_830,N_776,N_696);
nand U831 (N_831,N_790,N_662);
or U832 (N_832,N_754,N_715);
and U833 (N_833,N_609,N_672);
and U834 (N_834,N_674,N_734);
nand U835 (N_835,N_718,N_727);
and U836 (N_836,N_775,N_701);
xnor U837 (N_837,N_770,N_755);
or U838 (N_838,N_666,N_686);
or U839 (N_839,N_768,N_633);
xnor U840 (N_840,N_622,N_733);
and U841 (N_841,N_652,N_657);
nand U842 (N_842,N_614,N_619);
xnor U843 (N_843,N_635,N_693);
nor U844 (N_844,N_641,N_621);
xor U845 (N_845,N_732,N_628);
or U846 (N_846,N_638,N_661);
nor U847 (N_847,N_637,N_769);
nor U848 (N_848,N_712,N_747);
xor U849 (N_849,N_656,N_740);
xor U850 (N_850,N_751,N_788);
nand U851 (N_851,N_684,N_759);
nand U852 (N_852,N_654,N_623);
nand U853 (N_853,N_717,N_762);
or U854 (N_854,N_706,N_698);
and U855 (N_855,N_649,N_781);
nor U856 (N_856,N_797,N_681);
and U857 (N_857,N_707,N_723);
nand U858 (N_858,N_692,N_689);
nand U859 (N_859,N_659,N_772);
nor U860 (N_860,N_764,N_730);
xnor U861 (N_861,N_615,N_606);
nand U862 (N_862,N_600,N_673);
xnor U863 (N_863,N_665,N_780);
nand U864 (N_864,N_799,N_708);
and U865 (N_865,N_700,N_744);
or U866 (N_866,N_688,N_679);
or U867 (N_867,N_753,N_640);
and U868 (N_868,N_766,N_616);
xnor U869 (N_869,N_736,N_699);
or U870 (N_870,N_625,N_603);
nand U871 (N_871,N_795,N_735);
and U872 (N_872,N_729,N_658);
nand U873 (N_873,N_724,N_650);
nand U874 (N_874,N_634,N_728);
nor U875 (N_875,N_710,N_702);
or U876 (N_876,N_745,N_704);
or U877 (N_877,N_648,N_643);
or U878 (N_878,N_639,N_743);
xor U879 (N_879,N_691,N_618);
xor U880 (N_880,N_758,N_779);
nand U881 (N_881,N_771,N_778);
nand U882 (N_882,N_678,N_647);
or U883 (N_883,N_620,N_792);
or U884 (N_884,N_789,N_746);
nand U885 (N_885,N_787,N_685);
or U886 (N_886,N_687,N_793);
xnor U887 (N_887,N_695,N_680);
nand U888 (N_888,N_602,N_655);
and U889 (N_889,N_653,N_612);
nor U890 (N_890,N_786,N_711);
nor U891 (N_891,N_782,N_726);
nand U892 (N_892,N_714,N_783);
and U893 (N_893,N_719,N_721);
or U894 (N_894,N_670,N_629);
nand U895 (N_895,N_697,N_682);
xor U896 (N_896,N_750,N_611);
and U897 (N_897,N_709,N_756);
nand U898 (N_898,N_796,N_763);
xor U899 (N_899,N_791,N_694);
and U900 (N_900,N_607,N_695);
nand U901 (N_901,N_659,N_771);
or U902 (N_902,N_728,N_754);
xnor U903 (N_903,N_652,N_656);
or U904 (N_904,N_626,N_628);
nor U905 (N_905,N_636,N_619);
nand U906 (N_906,N_727,N_741);
and U907 (N_907,N_651,N_798);
nor U908 (N_908,N_747,N_761);
nand U909 (N_909,N_683,N_732);
and U910 (N_910,N_763,N_630);
or U911 (N_911,N_602,N_699);
xnor U912 (N_912,N_603,N_669);
nor U913 (N_913,N_744,N_792);
xor U914 (N_914,N_651,N_781);
or U915 (N_915,N_744,N_781);
nand U916 (N_916,N_677,N_741);
and U917 (N_917,N_708,N_748);
and U918 (N_918,N_650,N_686);
nor U919 (N_919,N_696,N_695);
and U920 (N_920,N_789,N_719);
nor U921 (N_921,N_642,N_702);
or U922 (N_922,N_710,N_749);
xnor U923 (N_923,N_748,N_602);
nor U924 (N_924,N_663,N_733);
or U925 (N_925,N_687,N_704);
xnor U926 (N_926,N_696,N_781);
nand U927 (N_927,N_709,N_641);
nand U928 (N_928,N_692,N_688);
or U929 (N_929,N_697,N_796);
and U930 (N_930,N_782,N_658);
nand U931 (N_931,N_756,N_614);
or U932 (N_932,N_704,N_724);
nand U933 (N_933,N_607,N_783);
and U934 (N_934,N_635,N_697);
or U935 (N_935,N_737,N_651);
nor U936 (N_936,N_735,N_631);
nand U937 (N_937,N_704,N_648);
nand U938 (N_938,N_757,N_604);
nand U939 (N_939,N_739,N_696);
and U940 (N_940,N_724,N_696);
xor U941 (N_941,N_693,N_671);
or U942 (N_942,N_637,N_646);
xor U943 (N_943,N_662,N_694);
nor U944 (N_944,N_616,N_619);
nand U945 (N_945,N_771,N_734);
nor U946 (N_946,N_692,N_640);
or U947 (N_947,N_661,N_719);
nand U948 (N_948,N_639,N_750);
nand U949 (N_949,N_770,N_752);
nand U950 (N_950,N_731,N_792);
nand U951 (N_951,N_706,N_785);
nor U952 (N_952,N_656,N_685);
xnor U953 (N_953,N_680,N_688);
nor U954 (N_954,N_617,N_736);
and U955 (N_955,N_632,N_640);
xnor U956 (N_956,N_726,N_610);
nor U957 (N_957,N_631,N_775);
xnor U958 (N_958,N_767,N_697);
and U959 (N_959,N_741,N_661);
or U960 (N_960,N_671,N_734);
or U961 (N_961,N_641,N_721);
and U962 (N_962,N_699,N_686);
nand U963 (N_963,N_763,N_753);
nand U964 (N_964,N_633,N_739);
or U965 (N_965,N_603,N_697);
nand U966 (N_966,N_613,N_758);
nor U967 (N_967,N_676,N_784);
and U968 (N_968,N_782,N_646);
xor U969 (N_969,N_668,N_673);
or U970 (N_970,N_707,N_698);
nor U971 (N_971,N_674,N_764);
and U972 (N_972,N_630,N_651);
and U973 (N_973,N_629,N_762);
and U974 (N_974,N_765,N_744);
nor U975 (N_975,N_630,N_669);
or U976 (N_976,N_676,N_682);
xor U977 (N_977,N_739,N_768);
or U978 (N_978,N_725,N_604);
xnor U979 (N_979,N_764,N_680);
and U980 (N_980,N_641,N_717);
and U981 (N_981,N_617,N_702);
nor U982 (N_982,N_670,N_681);
nor U983 (N_983,N_714,N_626);
xnor U984 (N_984,N_708,N_730);
or U985 (N_985,N_789,N_664);
and U986 (N_986,N_728,N_646);
xor U987 (N_987,N_699,N_653);
and U988 (N_988,N_771,N_755);
nand U989 (N_989,N_657,N_693);
or U990 (N_990,N_644,N_788);
and U991 (N_991,N_711,N_778);
nand U992 (N_992,N_674,N_714);
and U993 (N_993,N_731,N_637);
nor U994 (N_994,N_726,N_742);
nand U995 (N_995,N_602,N_646);
xor U996 (N_996,N_738,N_704);
xor U997 (N_997,N_749,N_654);
nand U998 (N_998,N_652,N_798);
nand U999 (N_999,N_733,N_728);
nand U1000 (N_1000,N_994,N_946);
or U1001 (N_1001,N_947,N_934);
xnor U1002 (N_1002,N_851,N_948);
or U1003 (N_1003,N_996,N_945);
nor U1004 (N_1004,N_972,N_915);
nor U1005 (N_1005,N_818,N_888);
nand U1006 (N_1006,N_866,N_995);
nand U1007 (N_1007,N_839,N_925);
nor U1008 (N_1008,N_922,N_989);
or U1009 (N_1009,N_809,N_846);
and U1010 (N_1010,N_817,N_858);
nand U1011 (N_1011,N_831,N_992);
or U1012 (N_1012,N_845,N_918);
and U1013 (N_1013,N_813,N_834);
and U1014 (N_1014,N_990,N_808);
and U1015 (N_1015,N_886,N_859);
or U1016 (N_1016,N_953,N_853);
or U1017 (N_1017,N_904,N_971);
and U1018 (N_1018,N_826,N_832);
or U1019 (N_1019,N_816,N_857);
and U1020 (N_1020,N_889,N_968);
xnor U1021 (N_1021,N_824,N_967);
nand U1022 (N_1022,N_890,N_867);
nor U1023 (N_1023,N_969,N_923);
nand U1024 (N_1024,N_898,N_848);
and U1025 (N_1025,N_981,N_927);
or U1026 (N_1026,N_962,N_951);
nor U1027 (N_1027,N_812,N_840);
or U1028 (N_1028,N_957,N_805);
or U1029 (N_1029,N_895,N_985);
nor U1030 (N_1030,N_865,N_965);
nor U1031 (N_1031,N_928,N_833);
or U1032 (N_1032,N_872,N_932);
nor U1033 (N_1033,N_862,N_884);
nor U1034 (N_1034,N_823,N_900);
nor U1035 (N_1035,N_970,N_893);
and U1036 (N_1036,N_949,N_986);
nor U1037 (N_1037,N_885,N_863);
xor U1038 (N_1038,N_919,N_850);
xnor U1039 (N_1039,N_973,N_984);
nand U1040 (N_1040,N_997,N_914);
nand U1041 (N_1041,N_933,N_838);
and U1042 (N_1042,N_881,N_908);
or U1043 (N_1043,N_912,N_894);
nor U1044 (N_1044,N_978,N_950);
xor U1045 (N_1045,N_980,N_938);
xor U1046 (N_1046,N_982,N_899);
or U1047 (N_1047,N_937,N_926);
nand U1048 (N_1048,N_993,N_820);
nor U1049 (N_1049,N_916,N_963);
xor U1050 (N_1050,N_920,N_860);
xnor U1051 (N_1051,N_913,N_902);
and U1052 (N_1052,N_954,N_873);
and U1053 (N_1053,N_880,N_979);
or U1054 (N_1054,N_877,N_905);
or U1055 (N_1055,N_958,N_806);
xnor U1056 (N_1056,N_906,N_959);
and U1057 (N_1057,N_821,N_829);
nor U1058 (N_1058,N_856,N_909);
nor U1059 (N_1059,N_956,N_944);
and U1060 (N_1060,N_861,N_952);
xnor U1061 (N_1061,N_935,N_819);
xor U1062 (N_1062,N_843,N_849);
nor U1063 (N_1063,N_929,N_942);
xor U1064 (N_1064,N_868,N_921);
xor U1065 (N_1065,N_847,N_977);
or U1066 (N_1066,N_910,N_917);
nor U1067 (N_1067,N_842,N_800);
xnor U1068 (N_1068,N_987,N_869);
or U1069 (N_1069,N_966,N_924);
or U1070 (N_1070,N_930,N_961);
and U1071 (N_1071,N_907,N_991);
nand U1072 (N_1072,N_830,N_943);
and U1073 (N_1073,N_998,N_854);
or U1074 (N_1074,N_988,N_941);
nand U1075 (N_1075,N_828,N_803);
and U1076 (N_1076,N_999,N_883);
nand U1077 (N_1077,N_825,N_835);
xnor U1078 (N_1078,N_976,N_960);
nand U1079 (N_1079,N_882,N_837);
nand U1080 (N_1080,N_855,N_807);
nor U1081 (N_1081,N_804,N_964);
nand U1082 (N_1082,N_827,N_844);
and U1083 (N_1083,N_870,N_802);
and U1084 (N_1084,N_911,N_891);
nor U1085 (N_1085,N_975,N_879);
nand U1086 (N_1086,N_852,N_814);
xor U1087 (N_1087,N_822,N_874);
or U1088 (N_1088,N_887,N_801);
and U1089 (N_1089,N_864,N_931);
and U1090 (N_1090,N_815,N_836);
nand U1091 (N_1091,N_811,N_955);
xnor U1092 (N_1092,N_897,N_936);
and U1093 (N_1093,N_878,N_876);
nand U1094 (N_1094,N_892,N_903);
xnor U1095 (N_1095,N_841,N_974);
and U1096 (N_1096,N_939,N_983);
and U1097 (N_1097,N_896,N_810);
xnor U1098 (N_1098,N_875,N_871);
nor U1099 (N_1099,N_901,N_940);
nand U1100 (N_1100,N_908,N_882);
and U1101 (N_1101,N_994,N_890);
and U1102 (N_1102,N_960,N_888);
or U1103 (N_1103,N_931,N_873);
nor U1104 (N_1104,N_973,N_978);
and U1105 (N_1105,N_981,N_807);
nor U1106 (N_1106,N_844,N_974);
xnor U1107 (N_1107,N_905,N_879);
or U1108 (N_1108,N_813,N_911);
nor U1109 (N_1109,N_995,N_992);
xnor U1110 (N_1110,N_976,N_854);
or U1111 (N_1111,N_898,N_869);
or U1112 (N_1112,N_836,N_816);
or U1113 (N_1113,N_984,N_865);
or U1114 (N_1114,N_879,N_809);
xor U1115 (N_1115,N_834,N_944);
xnor U1116 (N_1116,N_828,N_977);
nor U1117 (N_1117,N_893,N_838);
nand U1118 (N_1118,N_918,N_988);
nand U1119 (N_1119,N_880,N_872);
and U1120 (N_1120,N_949,N_840);
xnor U1121 (N_1121,N_991,N_981);
xnor U1122 (N_1122,N_938,N_933);
nand U1123 (N_1123,N_881,N_873);
nor U1124 (N_1124,N_903,N_817);
nand U1125 (N_1125,N_974,N_804);
xnor U1126 (N_1126,N_866,N_965);
and U1127 (N_1127,N_835,N_803);
xnor U1128 (N_1128,N_872,N_924);
or U1129 (N_1129,N_898,N_958);
nand U1130 (N_1130,N_910,N_983);
or U1131 (N_1131,N_855,N_816);
or U1132 (N_1132,N_802,N_998);
xor U1133 (N_1133,N_802,N_949);
nor U1134 (N_1134,N_807,N_991);
nand U1135 (N_1135,N_952,N_980);
and U1136 (N_1136,N_897,N_802);
and U1137 (N_1137,N_826,N_995);
nand U1138 (N_1138,N_927,N_923);
xor U1139 (N_1139,N_812,N_860);
and U1140 (N_1140,N_811,N_936);
and U1141 (N_1141,N_823,N_811);
and U1142 (N_1142,N_974,N_966);
nor U1143 (N_1143,N_999,N_806);
xor U1144 (N_1144,N_847,N_963);
xnor U1145 (N_1145,N_859,N_936);
xor U1146 (N_1146,N_989,N_888);
and U1147 (N_1147,N_831,N_801);
xnor U1148 (N_1148,N_965,N_856);
and U1149 (N_1149,N_985,N_885);
nand U1150 (N_1150,N_844,N_981);
xor U1151 (N_1151,N_894,N_994);
xnor U1152 (N_1152,N_983,N_878);
or U1153 (N_1153,N_909,N_857);
or U1154 (N_1154,N_939,N_826);
or U1155 (N_1155,N_852,N_951);
nand U1156 (N_1156,N_976,N_836);
nor U1157 (N_1157,N_933,N_856);
and U1158 (N_1158,N_811,N_942);
and U1159 (N_1159,N_949,N_960);
or U1160 (N_1160,N_924,N_909);
and U1161 (N_1161,N_905,N_841);
and U1162 (N_1162,N_851,N_935);
and U1163 (N_1163,N_956,N_932);
nand U1164 (N_1164,N_915,N_835);
nor U1165 (N_1165,N_940,N_866);
and U1166 (N_1166,N_936,N_990);
xnor U1167 (N_1167,N_923,N_812);
xor U1168 (N_1168,N_847,N_913);
nor U1169 (N_1169,N_958,N_858);
and U1170 (N_1170,N_805,N_874);
or U1171 (N_1171,N_939,N_842);
nand U1172 (N_1172,N_826,N_809);
nor U1173 (N_1173,N_860,N_872);
nor U1174 (N_1174,N_804,N_897);
nand U1175 (N_1175,N_988,N_814);
or U1176 (N_1176,N_995,N_984);
or U1177 (N_1177,N_992,N_976);
and U1178 (N_1178,N_876,N_885);
xnor U1179 (N_1179,N_963,N_901);
nand U1180 (N_1180,N_801,N_937);
nor U1181 (N_1181,N_975,N_866);
xor U1182 (N_1182,N_948,N_847);
xor U1183 (N_1183,N_960,N_860);
nor U1184 (N_1184,N_838,N_836);
nand U1185 (N_1185,N_845,N_997);
or U1186 (N_1186,N_826,N_964);
xor U1187 (N_1187,N_842,N_941);
and U1188 (N_1188,N_941,N_839);
and U1189 (N_1189,N_919,N_836);
or U1190 (N_1190,N_993,N_910);
nor U1191 (N_1191,N_804,N_891);
nor U1192 (N_1192,N_828,N_931);
nand U1193 (N_1193,N_966,N_875);
xor U1194 (N_1194,N_961,N_842);
nand U1195 (N_1195,N_909,N_992);
nand U1196 (N_1196,N_982,N_990);
or U1197 (N_1197,N_958,N_870);
and U1198 (N_1198,N_803,N_847);
or U1199 (N_1199,N_904,N_960);
nand U1200 (N_1200,N_1095,N_1179);
nor U1201 (N_1201,N_1079,N_1115);
nand U1202 (N_1202,N_1043,N_1122);
and U1203 (N_1203,N_1015,N_1141);
xor U1204 (N_1204,N_1076,N_1157);
nor U1205 (N_1205,N_1128,N_1192);
nand U1206 (N_1206,N_1139,N_1045);
or U1207 (N_1207,N_1172,N_1006);
and U1208 (N_1208,N_1107,N_1037);
and U1209 (N_1209,N_1022,N_1024);
or U1210 (N_1210,N_1193,N_1099);
nor U1211 (N_1211,N_1170,N_1199);
nor U1212 (N_1212,N_1121,N_1031);
nor U1213 (N_1213,N_1020,N_1028);
and U1214 (N_1214,N_1194,N_1191);
nand U1215 (N_1215,N_1035,N_1077);
or U1216 (N_1216,N_1181,N_1018);
or U1217 (N_1217,N_1110,N_1019);
xor U1218 (N_1218,N_1174,N_1142);
xnor U1219 (N_1219,N_1027,N_1114);
nor U1220 (N_1220,N_1113,N_1053);
nand U1221 (N_1221,N_1066,N_1189);
nor U1222 (N_1222,N_1080,N_1117);
nor U1223 (N_1223,N_1176,N_1138);
nor U1224 (N_1224,N_1106,N_1088);
nor U1225 (N_1225,N_1148,N_1153);
nor U1226 (N_1226,N_1162,N_1118);
xnor U1227 (N_1227,N_1154,N_1057);
nor U1228 (N_1228,N_1007,N_1084);
nor U1229 (N_1229,N_1071,N_1186);
or U1230 (N_1230,N_1047,N_1078);
xor U1231 (N_1231,N_1168,N_1145);
or U1232 (N_1232,N_1041,N_1025);
or U1233 (N_1233,N_1184,N_1159);
or U1234 (N_1234,N_1188,N_1091);
nand U1235 (N_1235,N_1119,N_1166);
nand U1236 (N_1236,N_1001,N_1058);
nor U1237 (N_1237,N_1010,N_1152);
nand U1238 (N_1238,N_1120,N_1131);
xor U1239 (N_1239,N_1195,N_1156);
xnor U1240 (N_1240,N_1090,N_1158);
and U1241 (N_1241,N_1144,N_1161);
and U1242 (N_1242,N_1070,N_1183);
and U1243 (N_1243,N_1116,N_1044);
nor U1244 (N_1244,N_1173,N_1180);
xnor U1245 (N_1245,N_1002,N_1125);
xnor U1246 (N_1246,N_1013,N_1177);
xnor U1247 (N_1247,N_1187,N_1032);
and U1248 (N_1248,N_1096,N_1178);
nor U1249 (N_1249,N_1038,N_1104);
nor U1250 (N_1250,N_1069,N_1029);
xor U1251 (N_1251,N_1050,N_1127);
nand U1252 (N_1252,N_1098,N_1101);
and U1253 (N_1253,N_1124,N_1163);
nor U1254 (N_1254,N_1137,N_1075);
nor U1255 (N_1255,N_1169,N_1133);
nor U1256 (N_1256,N_1059,N_1065);
or U1257 (N_1257,N_1112,N_1033);
xnor U1258 (N_1258,N_1060,N_1012);
and U1259 (N_1259,N_1140,N_1083);
nand U1260 (N_1260,N_1042,N_1171);
and U1261 (N_1261,N_1009,N_1100);
xor U1262 (N_1262,N_1052,N_1064);
xor U1263 (N_1263,N_1026,N_1167);
or U1264 (N_1264,N_1061,N_1000);
or U1265 (N_1265,N_1132,N_1040);
or U1266 (N_1266,N_1087,N_1198);
and U1267 (N_1267,N_1067,N_1185);
nand U1268 (N_1268,N_1062,N_1004);
nand U1269 (N_1269,N_1092,N_1164);
or U1270 (N_1270,N_1046,N_1036);
nor U1271 (N_1271,N_1126,N_1103);
or U1272 (N_1272,N_1051,N_1021);
nand U1273 (N_1273,N_1135,N_1094);
nor U1274 (N_1274,N_1182,N_1014);
and U1275 (N_1275,N_1097,N_1034);
nor U1276 (N_1276,N_1196,N_1081);
xor U1277 (N_1277,N_1109,N_1160);
or U1278 (N_1278,N_1049,N_1017);
or U1279 (N_1279,N_1111,N_1011);
or U1280 (N_1280,N_1030,N_1054);
nor U1281 (N_1281,N_1197,N_1149);
or U1282 (N_1282,N_1063,N_1143);
and U1283 (N_1283,N_1102,N_1086);
nand U1284 (N_1284,N_1136,N_1165);
xor U1285 (N_1285,N_1039,N_1008);
nor U1286 (N_1286,N_1175,N_1130);
nor U1287 (N_1287,N_1023,N_1146);
nor U1288 (N_1288,N_1190,N_1072);
or U1289 (N_1289,N_1134,N_1129);
nor U1290 (N_1290,N_1093,N_1147);
nand U1291 (N_1291,N_1155,N_1151);
xnor U1292 (N_1292,N_1150,N_1082);
or U1293 (N_1293,N_1003,N_1016);
xnor U1294 (N_1294,N_1068,N_1055);
nor U1295 (N_1295,N_1089,N_1123);
nor U1296 (N_1296,N_1073,N_1005);
xor U1297 (N_1297,N_1074,N_1105);
xnor U1298 (N_1298,N_1108,N_1085);
nand U1299 (N_1299,N_1048,N_1056);
nand U1300 (N_1300,N_1135,N_1078);
xor U1301 (N_1301,N_1115,N_1178);
nor U1302 (N_1302,N_1161,N_1134);
nor U1303 (N_1303,N_1110,N_1103);
nor U1304 (N_1304,N_1067,N_1146);
and U1305 (N_1305,N_1017,N_1031);
or U1306 (N_1306,N_1130,N_1119);
nand U1307 (N_1307,N_1107,N_1134);
xnor U1308 (N_1308,N_1148,N_1037);
nor U1309 (N_1309,N_1103,N_1081);
or U1310 (N_1310,N_1085,N_1069);
xnor U1311 (N_1311,N_1129,N_1117);
and U1312 (N_1312,N_1172,N_1093);
or U1313 (N_1313,N_1026,N_1127);
xor U1314 (N_1314,N_1104,N_1135);
xnor U1315 (N_1315,N_1026,N_1131);
or U1316 (N_1316,N_1122,N_1077);
or U1317 (N_1317,N_1143,N_1044);
and U1318 (N_1318,N_1103,N_1199);
nor U1319 (N_1319,N_1109,N_1083);
nand U1320 (N_1320,N_1172,N_1199);
xnor U1321 (N_1321,N_1051,N_1112);
nor U1322 (N_1322,N_1195,N_1065);
and U1323 (N_1323,N_1106,N_1125);
xor U1324 (N_1324,N_1011,N_1174);
xnor U1325 (N_1325,N_1034,N_1009);
nand U1326 (N_1326,N_1167,N_1047);
nand U1327 (N_1327,N_1175,N_1033);
xor U1328 (N_1328,N_1091,N_1100);
or U1329 (N_1329,N_1122,N_1066);
nor U1330 (N_1330,N_1110,N_1038);
nor U1331 (N_1331,N_1135,N_1164);
xor U1332 (N_1332,N_1031,N_1020);
nor U1333 (N_1333,N_1170,N_1049);
or U1334 (N_1334,N_1081,N_1111);
nor U1335 (N_1335,N_1124,N_1003);
xor U1336 (N_1336,N_1082,N_1019);
nand U1337 (N_1337,N_1123,N_1090);
xnor U1338 (N_1338,N_1174,N_1090);
or U1339 (N_1339,N_1106,N_1080);
xnor U1340 (N_1340,N_1026,N_1071);
and U1341 (N_1341,N_1029,N_1098);
nand U1342 (N_1342,N_1169,N_1017);
nor U1343 (N_1343,N_1049,N_1048);
nor U1344 (N_1344,N_1170,N_1091);
and U1345 (N_1345,N_1065,N_1187);
xnor U1346 (N_1346,N_1110,N_1055);
xnor U1347 (N_1347,N_1087,N_1052);
xor U1348 (N_1348,N_1149,N_1103);
xor U1349 (N_1349,N_1075,N_1033);
xor U1350 (N_1350,N_1032,N_1028);
and U1351 (N_1351,N_1041,N_1082);
xor U1352 (N_1352,N_1149,N_1157);
nand U1353 (N_1353,N_1152,N_1081);
nand U1354 (N_1354,N_1195,N_1095);
nor U1355 (N_1355,N_1011,N_1082);
xnor U1356 (N_1356,N_1043,N_1198);
or U1357 (N_1357,N_1140,N_1164);
or U1358 (N_1358,N_1051,N_1132);
and U1359 (N_1359,N_1035,N_1110);
and U1360 (N_1360,N_1157,N_1108);
nor U1361 (N_1361,N_1177,N_1109);
xnor U1362 (N_1362,N_1023,N_1194);
and U1363 (N_1363,N_1125,N_1118);
or U1364 (N_1364,N_1132,N_1073);
nor U1365 (N_1365,N_1039,N_1160);
and U1366 (N_1366,N_1061,N_1177);
xnor U1367 (N_1367,N_1182,N_1064);
or U1368 (N_1368,N_1170,N_1142);
or U1369 (N_1369,N_1126,N_1178);
and U1370 (N_1370,N_1166,N_1057);
nand U1371 (N_1371,N_1152,N_1082);
nor U1372 (N_1372,N_1000,N_1047);
nor U1373 (N_1373,N_1143,N_1110);
nand U1374 (N_1374,N_1054,N_1104);
and U1375 (N_1375,N_1070,N_1187);
or U1376 (N_1376,N_1193,N_1129);
xor U1377 (N_1377,N_1108,N_1074);
or U1378 (N_1378,N_1050,N_1051);
nand U1379 (N_1379,N_1056,N_1006);
or U1380 (N_1380,N_1152,N_1061);
xnor U1381 (N_1381,N_1159,N_1143);
and U1382 (N_1382,N_1115,N_1012);
and U1383 (N_1383,N_1097,N_1166);
or U1384 (N_1384,N_1009,N_1072);
nand U1385 (N_1385,N_1048,N_1109);
nor U1386 (N_1386,N_1154,N_1005);
nand U1387 (N_1387,N_1092,N_1045);
and U1388 (N_1388,N_1098,N_1043);
nor U1389 (N_1389,N_1186,N_1121);
nor U1390 (N_1390,N_1065,N_1080);
xor U1391 (N_1391,N_1160,N_1118);
nor U1392 (N_1392,N_1016,N_1127);
nor U1393 (N_1393,N_1175,N_1152);
nand U1394 (N_1394,N_1060,N_1166);
or U1395 (N_1395,N_1081,N_1056);
and U1396 (N_1396,N_1177,N_1028);
nand U1397 (N_1397,N_1183,N_1087);
nand U1398 (N_1398,N_1104,N_1024);
or U1399 (N_1399,N_1038,N_1195);
xor U1400 (N_1400,N_1378,N_1278);
and U1401 (N_1401,N_1321,N_1319);
xor U1402 (N_1402,N_1209,N_1362);
or U1403 (N_1403,N_1316,N_1385);
xor U1404 (N_1404,N_1365,N_1358);
xnor U1405 (N_1405,N_1201,N_1202);
xnor U1406 (N_1406,N_1324,N_1268);
nor U1407 (N_1407,N_1375,N_1264);
and U1408 (N_1408,N_1370,N_1219);
nand U1409 (N_1409,N_1253,N_1303);
nand U1410 (N_1410,N_1223,N_1386);
nand U1411 (N_1411,N_1363,N_1346);
or U1412 (N_1412,N_1329,N_1397);
or U1413 (N_1413,N_1238,N_1298);
or U1414 (N_1414,N_1206,N_1311);
nand U1415 (N_1415,N_1340,N_1344);
nor U1416 (N_1416,N_1350,N_1280);
nor U1417 (N_1417,N_1301,N_1244);
nand U1418 (N_1418,N_1338,N_1247);
nor U1419 (N_1419,N_1282,N_1312);
nor U1420 (N_1420,N_1214,N_1334);
xnor U1421 (N_1421,N_1349,N_1366);
or U1422 (N_1422,N_1302,N_1304);
or U1423 (N_1423,N_1360,N_1377);
and U1424 (N_1424,N_1314,N_1291);
xor U1425 (N_1425,N_1277,N_1379);
nor U1426 (N_1426,N_1242,N_1252);
nand U1427 (N_1427,N_1216,N_1293);
or U1428 (N_1428,N_1212,N_1345);
or U1429 (N_1429,N_1336,N_1269);
xnor U1430 (N_1430,N_1305,N_1315);
nand U1431 (N_1431,N_1390,N_1245);
and U1432 (N_1432,N_1234,N_1309);
and U1433 (N_1433,N_1289,N_1263);
nor U1434 (N_1434,N_1356,N_1207);
xor U1435 (N_1435,N_1287,N_1297);
nor U1436 (N_1436,N_1387,N_1359);
xor U1437 (N_1437,N_1307,N_1352);
xnor U1438 (N_1438,N_1208,N_1230);
xnor U1439 (N_1439,N_1273,N_1200);
nor U1440 (N_1440,N_1239,N_1257);
or U1441 (N_1441,N_1317,N_1267);
nor U1442 (N_1442,N_1355,N_1380);
or U1443 (N_1443,N_1279,N_1292);
or U1444 (N_1444,N_1233,N_1225);
or U1445 (N_1445,N_1384,N_1248);
nor U1446 (N_1446,N_1299,N_1367);
nor U1447 (N_1447,N_1294,N_1353);
nand U1448 (N_1448,N_1393,N_1373);
and U1449 (N_1449,N_1332,N_1271);
nand U1450 (N_1450,N_1284,N_1262);
nand U1451 (N_1451,N_1213,N_1295);
or U1452 (N_1452,N_1374,N_1330);
xor U1453 (N_1453,N_1333,N_1325);
or U1454 (N_1454,N_1327,N_1256);
nand U1455 (N_1455,N_1364,N_1221);
and U1456 (N_1456,N_1335,N_1371);
xnor U1457 (N_1457,N_1396,N_1236);
nand U1458 (N_1458,N_1341,N_1235);
nand U1459 (N_1459,N_1226,N_1288);
and U1460 (N_1460,N_1372,N_1210);
nand U1461 (N_1461,N_1237,N_1222);
nor U1462 (N_1462,N_1231,N_1328);
nand U1463 (N_1463,N_1394,N_1398);
nand U1464 (N_1464,N_1337,N_1211);
xnor U1465 (N_1465,N_1250,N_1205);
xnor U1466 (N_1466,N_1218,N_1272);
nand U1467 (N_1467,N_1283,N_1204);
or U1468 (N_1468,N_1227,N_1246);
or U1469 (N_1469,N_1266,N_1389);
and U1470 (N_1470,N_1251,N_1254);
nand U1471 (N_1471,N_1348,N_1351);
xor U1472 (N_1472,N_1382,N_1376);
nand U1473 (N_1473,N_1260,N_1395);
and U1474 (N_1474,N_1275,N_1391);
or U1475 (N_1475,N_1331,N_1383);
nand U1476 (N_1476,N_1229,N_1215);
xor U1477 (N_1477,N_1381,N_1354);
nand U1478 (N_1478,N_1347,N_1342);
nor U1479 (N_1479,N_1296,N_1399);
and U1480 (N_1480,N_1217,N_1241);
nand U1481 (N_1481,N_1243,N_1249);
nand U1482 (N_1482,N_1228,N_1258);
or U1483 (N_1483,N_1240,N_1300);
or U1484 (N_1484,N_1286,N_1270);
nor U1485 (N_1485,N_1388,N_1310);
xor U1486 (N_1486,N_1224,N_1290);
xor U1487 (N_1487,N_1285,N_1232);
or U1488 (N_1488,N_1274,N_1392);
xor U1489 (N_1489,N_1281,N_1339);
xor U1490 (N_1490,N_1343,N_1306);
and U1491 (N_1491,N_1313,N_1322);
xnor U1492 (N_1492,N_1203,N_1265);
nor U1493 (N_1493,N_1308,N_1369);
xor U1494 (N_1494,N_1255,N_1361);
xor U1495 (N_1495,N_1323,N_1318);
nor U1496 (N_1496,N_1326,N_1320);
or U1497 (N_1497,N_1259,N_1261);
xnor U1498 (N_1498,N_1220,N_1357);
nand U1499 (N_1499,N_1368,N_1276);
xor U1500 (N_1500,N_1372,N_1383);
xor U1501 (N_1501,N_1245,N_1284);
or U1502 (N_1502,N_1212,N_1379);
nor U1503 (N_1503,N_1276,N_1250);
nand U1504 (N_1504,N_1362,N_1278);
nor U1505 (N_1505,N_1396,N_1224);
nor U1506 (N_1506,N_1347,N_1265);
and U1507 (N_1507,N_1262,N_1372);
nor U1508 (N_1508,N_1336,N_1228);
and U1509 (N_1509,N_1336,N_1283);
nor U1510 (N_1510,N_1398,N_1358);
xor U1511 (N_1511,N_1286,N_1376);
xor U1512 (N_1512,N_1292,N_1372);
nand U1513 (N_1513,N_1232,N_1264);
and U1514 (N_1514,N_1321,N_1216);
xnor U1515 (N_1515,N_1241,N_1222);
nand U1516 (N_1516,N_1274,N_1302);
or U1517 (N_1517,N_1334,N_1271);
xnor U1518 (N_1518,N_1233,N_1368);
nor U1519 (N_1519,N_1249,N_1367);
or U1520 (N_1520,N_1270,N_1202);
or U1521 (N_1521,N_1370,N_1293);
xor U1522 (N_1522,N_1210,N_1220);
xnor U1523 (N_1523,N_1386,N_1373);
nand U1524 (N_1524,N_1380,N_1314);
nand U1525 (N_1525,N_1208,N_1385);
or U1526 (N_1526,N_1348,N_1240);
xnor U1527 (N_1527,N_1287,N_1240);
and U1528 (N_1528,N_1237,N_1293);
or U1529 (N_1529,N_1333,N_1266);
nor U1530 (N_1530,N_1359,N_1398);
nand U1531 (N_1531,N_1219,N_1373);
or U1532 (N_1532,N_1245,N_1223);
xor U1533 (N_1533,N_1321,N_1234);
nand U1534 (N_1534,N_1362,N_1374);
and U1535 (N_1535,N_1355,N_1253);
xnor U1536 (N_1536,N_1200,N_1261);
or U1537 (N_1537,N_1306,N_1243);
or U1538 (N_1538,N_1384,N_1308);
xor U1539 (N_1539,N_1339,N_1324);
and U1540 (N_1540,N_1361,N_1395);
or U1541 (N_1541,N_1380,N_1301);
nand U1542 (N_1542,N_1295,N_1238);
nor U1543 (N_1543,N_1384,N_1216);
or U1544 (N_1544,N_1313,N_1301);
nand U1545 (N_1545,N_1322,N_1230);
and U1546 (N_1546,N_1368,N_1330);
nand U1547 (N_1547,N_1259,N_1366);
and U1548 (N_1548,N_1350,N_1243);
xor U1549 (N_1549,N_1213,N_1308);
nor U1550 (N_1550,N_1294,N_1224);
nor U1551 (N_1551,N_1329,N_1265);
nor U1552 (N_1552,N_1274,N_1399);
xnor U1553 (N_1553,N_1382,N_1235);
nand U1554 (N_1554,N_1341,N_1282);
and U1555 (N_1555,N_1239,N_1249);
nand U1556 (N_1556,N_1334,N_1331);
nor U1557 (N_1557,N_1251,N_1207);
xnor U1558 (N_1558,N_1328,N_1327);
xor U1559 (N_1559,N_1223,N_1330);
nor U1560 (N_1560,N_1278,N_1345);
nor U1561 (N_1561,N_1371,N_1364);
xnor U1562 (N_1562,N_1218,N_1298);
nor U1563 (N_1563,N_1242,N_1220);
nor U1564 (N_1564,N_1366,N_1203);
nand U1565 (N_1565,N_1269,N_1204);
xnor U1566 (N_1566,N_1224,N_1281);
nor U1567 (N_1567,N_1300,N_1343);
nand U1568 (N_1568,N_1399,N_1283);
nor U1569 (N_1569,N_1268,N_1354);
and U1570 (N_1570,N_1323,N_1378);
nand U1571 (N_1571,N_1306,N_1395);
or U1572 (N_1572,N_1296,N_1304);
nor U1573 (N_1573,N_1247,N_1379);
nor U1574 (N_1574,N_1349,N_1299);
nand U1575 (N_1575,N_1266,N_1309);
nand U1576 (N_1576,N_1207,N_1220);
xor U1577 (N_1577,N_1256,N_1276);
or U1578 (N_1578,N_1377,N_1370);
nand U1579 (N_1579,N_1261,N_1256);
nand U1580 (N_1580,N_1288,N_1247);
nand U1581 (N_1581,N_1391,N_1352);
or U1582 (N_1582,N_1351,N_1248);
or U1583 (N_1583,N_1270,N_1323);
or U1584 (N_1584,N_1391,N_1343);
xnor U1585 (N_1585,N_1382,N_1367);
xnor U1586 (N_1586,N_1328,N_1398);
xor U1587 (N_1587,N_1273,N_1315);
nor U1588 (N_1588,N_1382,N_1236);
nand U1589 (N_1589,N_1291,N_1323);
nor U1590 (N_1590,N_1358,N_1253);
or U1591 (N_1591,N_1310,N_1379);
nor U1592 (N_1592,N_1365,N_1211);
nand U1593 (N_1593,N_1291,N_1262);
or U1594 (N_1594,N_1349,N_1310);
and U1595 (N_1595,N_1320,N_1256);
and U1596 (N_1596,N_1228,N_1290);
nor U1597 (N_1597,N_1282,N_1253);
xnor U1598 (N_1598,N_1355,N_1393);
nor U1599 (N_1599,N_1325,N_1235);
and U1600 (N_1600,N_1433,N_1582);
nor U1601 (N_1601,N_1503,N_1404);
xnor U1602 (N_1602,N_1578,N_1484);
or U1603 (N_1603,N_1471,N_1499);
nand U1604 (N_1604,N_1485,N_1421);
and U1605 (N_1605,N_1406,N_1436);
xor U1606 (N_1606,N_1464,N_1599);
nor U1607 (N_1607,N_1512,N_1491);
and U1608 (N_1608,N_1497,N_1530);
nor U1609 (N_1609,N_1567,N_1597);
or U1610 (N_1610,N_1462,N_1495);
and U1611 (N_1611,N_1415,N_1532);
nor U1612 (N_1612,N_1470,N_1524);
and U1613 (N_1613,N_1443,N_1453);
or U1614 (N_1614,N_1434,N_1549);
or U1615 (N_1615,N_1487,N_1452);
and U1616 (N_1616,N_1423,N_1427);
or U1617 (N_1617,N_1554,N_1426);
nand U1618 (N_1618,N_1449,N_1456);
xnor U1619 (N_1619,N_1569,N_1528);
and U1620 (N_1620,N_1424,N_1454);
xnor U1621 (N_1621,N_1508,N_1409);
nand U1622 (N_1622,N_1593,N_1498);
or U1623 (N_1623,N_1517,N_1515);
nand U1624 (N_1624,N_1442,N_1475);
and U1625 (N_1625,N_1510,N_1556);
nand U1626 (N_1626,N_1403,N_1466);
and U1627 (N_1627,N_1457,N_1521);
xnor U1628 (N_1628,N_1458,N_1565);
and U1629 (N_1629,N_1420,N_1562);
nand U1630 (N_1630,N_1410,N_1496);
nand U1631 (N_1631,N_1438,N_1579);
nor U1632 (N_1632,N_1505,N_1595);
nor U1633 (N_1633,N_1504,N_1555);
nor U1634 (N_1634,N_1586,N_1590);
or U1635 (N_1635,N_1402,N_1479);
or U1636 (N_1636,N_1523,N_1440);
nand U1637 (N_1637,N_1494,N_1511);
and U1638 (N_1638,N_1489,N_1463);
xnor U1639 (N_1639,N_1431,N_1537);
nand U1640 (N_1640,N_1576,N_1450);
xor U1641 (N_1641,N_1455,N_1577);
nor U1642 (N_1642,N_1566,N_1563);
xnor U1643 (N_1643,N_1430,N_1509);
or U1644 (N_1644,N_1535,N_1570);
xnor U1645 (N_1645,N_1414,N_1598);
xnor U1646 (N_1646,N_1544,N_1437);
xor U1647 (N_1647,N_1529,N_1413);
nor U1648 (N_1648,N_1407,N_1435);
nand U1649 (N_1649,N_1419,N_1575);
nand U1650 (N_1650,N_1416,N_1520);
and U1651 (N_1651,N_1418,N_1518);
or U1652 (N_1652,N_1459,N_1548);
nor U1653 (N_1653,N_1506,N_1501);
nand U1654 (N_1654,N_1559,N_1568);
nor U1655 (N_1655,N_1592,N_1447);
xnor U1656 (N_1656,N_1468,N_1526);
xor U1657 (N_1657,N_1461,N_1588);
xor U1658 (N_1658,N_1561,N_1546);
nand U1659 (N_1659,N_1467,N_1401);
xnor U1660 (N_1660,N_1451,N_1589);
xor U1661 (N_1661,N_1581,N_1533);
nor U1662 (N_1662,N_1465,N_1596);
xor U1663 (N_1663,N_1448,N_1584);
and U1664 (N_1664,N_1490,N_1486);
and U1665 (N_1665,N_1408,N_1591);
xor U1666 (N_1666,N_1432,N_1594);
and U1667 (N_1667,N_1560,N_1516);
and U1668 (N_1668,N_1543,N_1445);
or U1669 (N_1669,N_1514,N_1527);
xor U1670 (N_1670,N_1564,N_1477);
xor U1671 (N_1671,N_1488,N_1476);
or U1672 (N_1672,N_1552,N_1412);
nor U1673 (N_1673,N_1580,N_1478);
nor U1674 (N_1674,N_1553,N_1531);
nand U1675 (N_1675,N_1460,N_1469);
xor U1676 (N_1676,N_1583,N_1541);
or U1677 (N_1677,N_1472,N_1439);
xnor U1678 (N_1678,N_1500,N_1446);
and U1679 (N_1679,N_1539,N_1473);
xnor U1680 (N_1680,N_1441,N_1502);
and U1681 (N_1681,N_1571,N_1558);
nand U1682 (N_1682,N_1405,N_1400);
or U1683 (N_1683,N_1425,N_1481);
xnor U1684 (N_1684,N_1482,N_1429);
and U1685 (N_1685,N_1492,N_1483);
xor U1686 (N_1686,N_1587,N_1540);
nor U1687 (N_1687,N_1574,N_1545);
nand U1688 (N_1688,N_1551,N_1519);
nor U1689 (N_1689,N_1417,N_1538);
and U1690 (N_1690,N_1585,N_1411);
nor U1691 (N_1691,N_1444,N_1557);
xnor U1692 (N_1692,N_1480,N_1474);
nand U1693 (N_1693,N_1536,N_1428);
and U1694 (N_1694,N_1542,N_1573);
xnor U1695 (N_1695,N_1522,N_1550);
nor U1696 (N_1696,N_1493,N_1507);
nand U1697 (N_1697,N_1525,N_1513);
xor U1698 (N_1698,N_1547,N_1534);
or U1699 (N_1699,N_1572,N_1422);
nor U1700 (N_1700,N_1419,N_1574);
or U1701 (N_1701,N_1571,N_1581);
or U1702 (N_1702,N_1599,N_1593);
xnor U1703 (N_1703,N_1554,N_1450);
nor U1704 (N_1704,N_1525,N_1530);
nand U1705 (N_1705,N_1567,N_1547);
xnor U1706 (N_1706,N_1417,N_1500);
and U1707 (N_1707,N_1433,N_1576);
nand U1708 (N_1708,N_1541,N_1489);
or U1709 (N_1709,N_1471,N_1425);
nand U1710 (N_1710,N_1429,N_1521);
or U1711 (N_1711,N_1481,N_1593);
xnor U1712 (N_1712,N_1456,N_1586);
nand U1713 (N_1713,N_1412,N_1544);
nor U1714 (N_1714,N_1502,N_1487);
xnor U1715 (N_1715,N_1571,N_1559);
and U1716 (N_1716,N_1407,N_1538);
xor U1717 (N_1717,N_1425,N_1569);
nor U1718 (N_1718,N_1521,N_1496);
nand U1719 (N_1719,N_1534,N_1539);
nor U1720 (N_1720,N_1526,N_1518);
or U1721 (N_1721,N_1539,N_1584);
and U1722 (N_1722,N_1401,N_1503);
nand U1723 (N_1723,N_1556,N_1483);
nor U1724 (N_1724,N_1578,N_1478);
nand U1725 (N_1725,N_1535,N_1598);
and U1726 (N_1726,N_1547,N_1557);
nand U1727 (N_1727,N_1540,N_1535);
xnor U1728 (N_1728,N_1541,N_1454);
nor U1729 (N_1729,N_1527,N_1422);
nand U1730 (N_1730,N_1501,N_1596);
nand U1731 (N_1731,N_1402,N_1530);
or U1732 (N_1732,N_1484,N_1479);
or U1733 (N_1733,N_1539,N_1564);
nand U1734 (N_1734,N_1465,N_1429);
xnor U1735 (N_1735,N_1434,N_1443);
and U1736 (N_1736,N_1518,N_1520);
nand U1737 (N_1737,N_1510,N_1569);
xor U1738 (N_1738,N_1522,N_1430);
and U1739 (N_1739,N_1454,N_1552);
or U1740 (N_1740,N_1519,N_1579);
nand U1741 (N_1741,N_1571,N_1570);
or U1742 (N_1742,N_1544,N_1563);
and U1743 (N_1743,N_1475,N_1514);
xnor U1744 (N_1744,N_1468,N_1460);
or U1745 (N_1745,N_1438,N_1493);
xnor U1746 (N_1746,N_1535,N_1594);
nor U1747 (N_1747,N_1572,N_1481);
nand U1748 (N_1748,N_1454,N_1588);
and U1749 (N_1749,N_1530,N_1403);
nor U1750 (N_1750,N_1496,N_1488);
nor U1751 (N_1751,N_1433,N_1407);
nor U1752 (N_1752,N_1586,N_1481);
nand U1753 (N_1753,N_1491,N_1470);
nand U1754 (N_1754,N_1533,N_1506);
nor U1755 (N_1755,N_1596,N_1505);
nand U1756 (N_1756,N_1504,N_1458);
nand U1757 (N_1757,N_1489,N_1406);
nand U1758 (N_1758,N_1448,N_1509);
and U1759 (N_1759,N_1456,N_1580);
or U1760 (N_1760,N_1429,N_1419);
nor U1761 (N_1761,N_1420,N_1555);
and U1762 (N_1762,N_1515,N_1427);
nor U1763 (N_1763,N_1527,N_1525);
xnor U1764 (N_1764,N_1432,N_1557);
and U1765 (N_1765,N_1414,N_1445);
nor U1766 (N_1766,N_1424,N_1440);
and U1767 (N_1767,N_1426,N_1436);
or U1768 (N_1768,N_1535,N_1448);
nand U1769 (N_1769,N_1474,N_1516);
or U1770 (N_1770,N_1472,N_1560);
nand U1771 (N_1771,N_1489,N_1520);
or U1772 (N_1772,N_1532,N_1445);
xnor U1773 (N_1773,N_1534,N_1496);
or U1774 (N_1774,N_1579,N_1537);
xor U1775 (N_1775,N_1594,N_1475);
nand U1776 (N_1776,N_1454,N_1429);
nand U1777 (N_1777,N_1535,N_1509);
xnor U1778 (N_1778,N_1444,N_1411);
nand U1779 (N_1779,N_1503,N_1593);
xnor U1780 (N_1780,N_1561,N_1420);
or U1781 (N_1781,N_1510,N_1588);
nor U1782 (N_1782,N_1450,N_1483);
and U1783 (N_1783,N_1584,N_1462);
or U1784 (N_1784,N_1455,N_1535);
and U1785 (N_1785,N_1454,N_1595);
nor U1786 (N_1786,N_1545,N_1407);
xor U1787 (N_1787,N_1534,N_1592);
or U1788 (N_1788,N_1416,N_1454);
or U1789 (N_1789,N_1531,N_1551);
or U1790 (N_1790,N_1555,N_1511);
nor U1791 (N_1791,N_1559,N_1534);
and U1792 (N_1792,N_1528,N_1455);
nand U1793 (N_1793,N_1552,N_1476);
nor U1794 (N_1794,N_1576,N_1571);
nand U1795 (N_1795,N_1509,N_1596);
and U1796 (N_1796,N_1534,N_1562);
nand U1797 (N_1797,N_1507,N_1414);
xnor U1798 (N_1798,N_1418,N_1575);
or U1799 (N_1799,N_1525,N_1449);
nor U1800 (N_1800,N_1643,N_1687);
nand U1801 (N_1801,N_1600,N_1619);
nor U1802 (N_1802,N_1707,N_1751);
xnor U1803 (N_1803,N_1676,N_1659);
nor U1804 (N_1804,N_1628,N_1649);
nand U1805 (N_1805,N_1704,N_1702);
or U1806 (N_1806,N_1775,N_1694);
nand U1807 (N_1807,N_1716,N_1605);
and U1808 (N_1808,N_1798,N_1749);
nand U1809 (N_1809,N_1720,N_1698);
nand U1810 (N_1810,N_1647,N_1757);
nor U1811 (N_1811,N_1708,N_1705);
and U1812 (N_1812,N_1753,N_1756);
nor U1813 (N_1813,N_1731,N_1760);
or U1814 (N_1814,N_1642,N_1604);
or U1815 (N_1815,N_1664,N_1733);
nand U1816 (N_1816,N_1791,N_1685);
or U1817 (N_1817,N_1710,N_1742);
xnor U1818 (N_1818,N_1729,N_1671);
or U1819 (N_1819,N_1774,N_1673);
nor U1820 (N_1820,N_1657,N_1703);
or U1821 (N_1821,N_1741,N_1669);
xnor U1822 (N_1822,N_1624,N_1660);
nor U1823 (N_1823,N_1674,N_1721);
nor U1824 (N_1824,N_1693,N_1736);
or U1825 (N_1825,N_1670,N_1792);
nor U1826 (N_1826,N_1651,N_1725);
and U1827 (N_1827,N_1750,N_1747);
nand U1828 (N_1828,N_1691,N_1712);
nor U1829 (N_1829,N_1767,N_1606);
and U1830 (N_1830,N_1633,N_1745);
and U1831 (N_1831,N_1645,N_1728);
and U1832 (N_1832,N_1677,N_1778);
or U1833 (N_1833,N_1779,N_1615);
nor U1834 (N_1834,N_1630,N_1679);
nand U1835 (N_1835,N_1635,N_1709);
xor U1836 (N_1836,N_1672,N_1734);
and U1837 (N_1837,N_1607,N_1603);
or U1838 (N_1838,N_1795,N_1601);
nor U1839 (N_1839,N_1625,N_1665);
or U1840 (N_1840,N_1621,N_1663);
xor U1841 (N_1841,N_1675,N_1667);
xor U1842 (N_1842,N_1695,N_1688);
xnor U1843 (N_1843,N_1797,N_1771);
nor U1844 (N_1844,N_1654,N_1655);
or U1845 (N_1845,N_1656,N_1782);
nor U1846 (N_1846,N_1781,N_1784);
nor U1847 (N_1847,N_1769,N_1786);
or U1848 (N_1848,N_1648,N_1783);
xor U1849 (N_1849,N_1787,N_1761);
xor U1850 (N_1850,N_1653,N_1641);
and U1851 (N_1851,N_1780,N_1788);
xor U1852 (N_1852,N_1746,N_1732);
nor U1853 (N_1853,N_1699,N_1722);
or U1854 (N_1854,N_1661,N_1613);
or U1855 (N_1855,N_1759,N_1717);
nand U1856 (N_1856,N_1764,N_1730);
nand U1857 (N_1857,N_1611,N_1686);
xnor U1858 (N_1858,N_1714,N_1680);
xor U1859 (N_1859,N_1618,N_1754);
nor U1860 (N_1860,N_1683,N_1636);
xnor U1861 (N_1861,N_1627,N_1715);
nand U1862 (N_1862,N_1622,N_1637);
or U1863 (N_1863,N_1632,N_1638);
xor U1864 (N_1864,N_1737,N_1662);
xnor U1865 (N_1865,N_1614,N_1616);
nand U1866 (N_1866,N_1696,N_1748);
nand U1867 (N_1867,N_1689,N_1706);
or U1868 (N_1868,N_1773,N_1739);
xnor U1869 (N_1869,N_1765,N_1650);
nor U1870 (N_1870,N_1617,N_1793);
nor U1871 (N_1871,N_1701,N_1763);
xor U1872 (N_1872,N_1718,N_1738);
or U1873 (N_1873,N_1666,N_1678);
nor U1874 (N_1874,N_1755,N_1640);
or U1875 (N_1875,N_1724,N_1602);
and U1876 (N_1876,N_1770,N_1713);
or U1877 (N_1877,N_1629,N_1789);
nand U1878 (N_1878,N_1719,N_1668);
xnor U1879 (N_1879,N_1772,N_1639);
nor U1880 (N_1880,N_1612,N_1776);
and U1881 (N_1881,N_1652,N_1610);
and U1882 (N_1882,N_1758,N_1799);
or U1883 (N_1883,N_1684,N_1690);
or U1884 (N_1884,N_1609,N_1777);
or U1885 (N_1885,N_1631,N_1626);
nor U1886 (N_1886,N_1620,N_1796);
nor U1887 (N_1887,N_1681,N_1608);
xnor U1888 (N_1888,N_1723,N_1794);
and U1889 (N_1889,N_1646,N_1644);
xor U1890 (N_1890,N_1790,N_1700);
nand U1891 (N_1891,N_1623,N_1768);
nor U1892 (N_1892,N_1727,N_1711);
nor U1893 (N_1893,N_1634,N_1740);
and U1894 (N_1894,N_1785,N_1735);
nand U1895 (N_1895,N_1726,N_1692);
nor U1896 (N_1896,N_1766,N_1743);
or U1897 (N_1897,N_1752,N_1744);
nor U1898 (N_1898,N_1697,N_1682);
nand U1899 (N_1899,N_1658,N_1762);
and U1900 (N_1900,N_1767,N_1741);
nand U1901 (N_1901,N_1766,N_1798);
nand U1902 (N_1902,N_1777,N_1790);
nand U1903 (N_1903,N_1667,N_1668);
xor U1904 (N_1904,N_1748,N_1727);
and U1905 (N_1905,N_1650,N_1731);
or U1906 (N_1906,N_1610,N_1671);
nand U1907 (N_1907,N_1658,N_1737);
and U1908 (N_1908,N_1654,N_1630);
nor U1909 (N_1909,N_1646,N_1709);
or U1910 (N_1910,N_1773,N_1740);
and U1911 (N_1911,N_1788,N_1711);
xor U1912 (N_1912,N_1684,N_1648);
or U1913 (N_1913,N_1626,N_1668);
nor U1914 (N_1914,N_1677,N_1619);
or U1915 (N_1915,N_1720,N_1733);
nand U1916 (N_1916,N_1691,N_1660);
nand U1917 (N_1917,N_1651,N_1715);
or U1918 (N_1918,N_1631,N_1671);
or U1919 (N_1919,N_1653,N_1645);
and U1920 (N_1920,N_1707,N_1721);
xor U1921 (N_1921,N_1630,N_1644);
xor U1922 (N_1922,N_1777,N_1617);
nor U1923 (N_1923,N_1791,N_1662);
xnor U1924 (N_1924,N_1652,N_1770);
nor U1925 (N_1925,N_1689,N_1756);
and U1926 (N_1926,N_1601,N_1748);
and U1927 (N_1927,N_1772,N_1786);
nor U1928 (N_1928,N_1661,N_1692);
or U1929 (N_1929,N_1741,N_1736);
nand U1930 (N_1930,N_1743,N_1677);
or U1931 (N_1931,N_1678,N_1750);
nor U1932 (N_1932,N_1776,N_1651);
and U1933 (N_1933,N_1613,N_1649);
and U1934 (N_1934,N_1693,N_1661);
nand U1935 (N_1935,N_1692,N_1734);
or U1936 (N_1936,N_1677,N_1635);
nand U1937 (N_1937,N_1671,N_1790);
or U1938 (N_1938,N_1677,N_1672);
nand U1939 (N_1939,N_1767,N_1773);
or U1940 (N_1940,N_1645,N_1708);
and U1941 (N_1941,N_1653,N_1692);
or U1942 (N_1942,N_1617,N_1654);
xnor U1943 (N_1943,N_1604,N_1708);
or U1944 (N_1944,N_1734,N_1689);
and U1945 (N_1945,N_1655,N_1653);
nand U1946 (N_1946,N_1752,N_1653);
nand U1947 (N_1947,N_1618,N_1654);
and U1948 (N_1948,N_1691,N_1643);
nor U1949 (N_1949,N_1746,N_1627);
or U1950 (N_1950,N_1606,N_1724);
nand U1951 (N_1951,N_1653,N_1771);
xnor U1952 (N_1952,N_1757,N_1794);
and U1953 (N_1953,N_1622,N_1710);
nand U1954 (N_1954,N_1700,N_1799);
nand U1955 (N_1955,N_1751,N_1691);
nand U1956 (N_1956,N_1649,N_1687);
nand U1957 (N_1957,N_1662,N_1618);
or U1958 (N_1958,N_1614,N_1607);
and U1959 (N_1959,N_1776,N_1668);
and U1960 (N_1960,N_1757,N_1692);
xor U1961 (N_1961,N_1680,N_1643);
and U1962 (N_1962,N_1669,N_1676);
and U1963 (N_1963,N_1691,N_1656);
nand U1964 (N_1964,N_1681,N_1738);
nor U1965 (N_1965,N_1731,N_1728);
or U1966 (N_1966,N_1631,N_1787);
nor U1967 (N_1967,N_1671,N_1787);
and U1968 (N_1968,N_1777,N_1753);
or U1969 (N_1969,N_1710,N_1660);
or U1970 (N_1970,N_1607,N_1742);
nand U1971 (N_1971,N_1747,N_1763);
nand U1972 (N_1972,N_1628,N_1692);
and U1973 (N_1973,N_1606,N_1656);
xor U1974 (N_1974,N_1798,N_1709);
nand U1975 (N_1975,N_1638,N_1775);
xnor U1976 (N_1976,N_1716,N_1670);
xor U1977 (N_1977,N_1612,N_1685);
nand U1978 (N_1978,N_1678,N_1728);
or U1979 (N_1979,N_1771,N_1675);
and U1980 (N_1980,N_1798,N_1606);
and U1981 (N_1981,N_1611,N_1601);
xor U1982 (N_1982,N_1778,N_1661);
and U1983 (N_1983,N_1717,N_1792);
xor U1984 (N_1984,N_1628,N_1765);
or U1985 (N_1985,N_1757,N_1724);
nor U1986 (N_1986,N_1701,N_1655);
nand U1987 (N_1987,N_1734,N_1788);
and U1988 (N_1988,N_1674,N_1643);
or U1989 (N_1989,N_1773,N_1717);
xnor U1990 (N_1990,N_1658,N_1706);
or U1991 (N_1991,N_1733,N_1783);
and U1992 (N_1992,N_1631,N_1713);
nand U1993 (N_1993,N_1713,N_1671);
or U1994 (N_1994,N_1665,N_1660);
and U1995 (N_1995,N_1626,N_1624);
or U1996 (N_1996,N_1713,N_1775);
nor U1997 (N_1997,N_1740,N_1625);
nand U1998 (N_1998,N_1773,N_1704);
or U1999 (N_1999,N_1762,N_1621);
and U2000 (N_2000,N_1972,N_1940);
nand U2001 (N_2001,N_1961,N_1958);
or U2002 (N_2002,N_1866,N_1831);
nand U2003 (N_2003,N_1906,N_1800);
and U2004 (N_2004,N_1846,N_1809);
xnor U2005 (N_2005,N_1949,N_1818);
nand U2006 (N_2006,N_1914,N_1950);
nand U2007 (N_2007,N_1937,N_1882);
xnor U2008 (N_2008,N_1841,N_1852);
xor U2009 (N_2009,N_1998,N_1879);
nor U2010 (N_2010,N_1811,N_1808);
xnor U2011 (N_2011,N_1933,N_1918);
nor U2012 (N_2012,N_1920,N_1839);
nor U2013 (N_2013,N_1995,N_1911);
or U2014 (N_2014,N_1858,N_1985);
nand U2015 (N_2015,N_1968,N_1883);
and U2016 (N_2016,N_1910,N_1843);
nand U2017 (N_2017,N_1983,N_1942);
nor U2018 (N_2018,N_1824,N_1885);
and U2019 (N_2019,N_1963,N_1916);
nand U2020 (N_2020,N_1993,N_1935);
or U2021 (N_2021,N_1919,N_1817);
nand U2022 (N_2022,N_1897,N_1930);
nor U2023 (N_2023,N_1991,N_1978);
and U2024 (N_2024,N_1863,N_1975);
nand U2025 (N_2025,N_1842,N_1909);
xnor U2026 (N_2026,N_1861,N_1854);
nor U2027 (N_2027,N_1860,N_1871);
nand U2028 (N_2028,N_1822,N_1834);
xor U2029 (N_2029,N_1819,N_1801);
and U2030 (N_2030,N_1867,N_1838);
nor U2031 (N_2031,N_1812,N_1884);
nand U2032 (N_2032,N_1803,N_1954);
or U2033 (N_2033,N_1981,N_1980);
nor U2034 (N_2034,N_1889,N_1925);
nor U2035 (N_2035,N_1806,N_1924);
xor U2036 (N_2036,N_1965,N_1896);
and U2037 (N_2037,N_1805,N_1945);
nor U2038 (N_2038,N_1835,N_1874);
nand U2039 (N_2039,N_1880,N_1984);
or U2040 (N_2040,N_1959,N_1892);
or U2041 (N_2041,N_1922,N_1830);
nand U2042 (N_2042,N_1876,N_1999);
nand U2043 (N_2043,N_1888,N_1931);
nand U2044 (N_2044,N_1948,N_1926);
nand U2045 (N_2045,N_1979,N_1873);
and U2046 (N_2046,N_1836,N_1951);
nor U2047 (N_2047,N_1990,N_1849);
and U2048 (N_2048,N_1987,N_1804);
and U2049 (N_2049,N_1815,N_1820);
and U2050 (N_2050,N_1810,N_1960);
and U2051 (N_2051,N_1966,N_1977);
xnor U2052 (N_2052,N_1970,N_1992);
or U2053 (N_2053,N_1821,N_1816);
nor U2054 (N_2054,N_1907,N_1862);
xnor U2055 (N_2055,N_1807,N_1869);
or U2056 (N_2056,N_1957,N_1917);
and U2057 (N_2057,N_1829,N_1823);
nor U2058 (N_2058,N_1964,N_1886);
xnor U2059 (N_2059,N_1994,N_1974);
or U2060 (N_2060,N_1851,N_1915);
xnor U2061 (N_2061,N_1962,N_1941);
nor U2062 (N_2062,N_1996,N_1814);
nor U2063 (N_2063,N_1890,N_1899);
nor U2064 (N_2064,N_1903,N_1894);
and U2065 (N_2065,N_1900,N_1813);
or U2066 (N_2066,N_1904,N_1929);
nand U2067 (N_2067,N_1947,N_1825);
xnor U2068 (N_2068,N_1932,N_1912);
xnor U2069 (N_2069,N_1943,N_1967);
and U2070 (N_2070,N_1921,N_1895);
nor U2071 (N_2071,N_1857,N_1946);
and U2072 (N_2072,N_1971,N_1982);
nor U2073 (N_2073,N_1870,N_1905);
and U2074 (N_2074,N_1872,N_1848);
or U2075 (N_2075,N_1898,N_1908);
nor U2076 (N_2076,N_1901,N_1875);
nand U2077 (N_2077,N_1855,N_1850);
nor U2078 (N_2078,N_1923,N_1955);
or U2079 (N_2079,N_1826,N_1878);
nand U2080 (N_2080,N_1847,N_1988);
nor U2081 (N_2081,N_1939,N_1827);
nand U2082 (N_2082,N_1927,N_1853);
and U2083 (N_2083,N_1893,N_1856);
xor U2084 (N_2084,N_1868,N_1837);
and U2085 (N_2085,N_1865,N_1956);
nand U2086 (N_2086,N_1997,N_1986);
and U2087 (N_2087,N_1944,N_1840);
or U2088 (N_2088,N_1859,N_1928);
and U2089 (N_2089,N_1845,N_1891);
and U2090 (N_2090,N_1934,N_1989);
nor U2091 (N_2091,N_1832,N_1833);
nor U2092 (N_2092,N_1864,N_1828);
and U2093 (N_2093,N_1881,N_1887);
nand U2094 (N_2094,N_1952,N_1973);
nand U2095 (N_2095,N_1877,N_1976);
nand U2096 (N_2096,N_1902,N_1844);
nand U2097 (N_2097,N_1969,N_1802);
and U2098 (N_2098,N_1936,N_1938);
or U2099 (N_2099,N_1913,N_1953);
xnor U2100 (N_2100,N_1988,N_1955);
or U2101 (N_2101,N_1995,N_1910);
nand U2102 (N_2102,N_1986,N_1829);
nor U2103 (N_2103,N_1861,N_1856);
nand U2104 (N_2104,N_1935,N_1876);
and U2105 (N_2105,N_1919,N_1861);
and U2106 (N_2106,N_1895,N_1928);
xor U2107 (N_2107,N_1916,N_1990);
or U2108 (N_2108,N_1918,N_1959);
or U2109 (N_2109,N_1921,N_1891);
xnor U2110 (N_2110,N_1939,N_1850);
nand U2111 (N_2111,N_1875,N_1992);
or U2112 (N_2112,N_1884,N_1931);
nand U2113 (N_2113,N_1804,N_1949);
or U2114 (N_2114,N_1811,N_1830);
nor U2115 (N_2115,N_1820,N_1954);
xor U2116 (N_2116,N_1894,N_1929);
nand U2117 (N_2117,N_1869,N_1823);
or U2118 (N_2118,N_1879,N_1804);
nand U2119 (N_2119,N_1986,N_1957);
and U2120 (N_2120,N_1902,N_1965);
nor U2121 (N_2121,N_1998,N_1921);
nand U2122 (N_2122,N_1976,N_1852);
nor U2123 (N_2123,N_1837,N_1887);
nor U2124 (N_2124,N_1984,N_1936);
and U2125 (N_2125,N_1899,N_1835);
and U2126 (N_2126,N_1981,N_1817);
and U2127 (N_2127,N_1934,N_1923);
nand U2128 (N_2128,N_1949,N_1817);
and U2129 (N_2129,N_1971,N_1830);
nor U2130 (N_2130,N_1938,N_1863);
xor U2131 (N_2131,N_1940,N_1956);
and U2132 (N_2132,N_1923,N_1914);
and U2133 (N_2133,N_1865,N_1885);
or U2134 (N_2134,N_1843,N_1914);
xnor U2135 (N_2135,N_1862,N_1853);
and U2136 (N_2136,N_1964,N_1962);
xnor U2137 (N_2137,N_1920,N_1990);
nand U2138 (N_2138,N_1857,N_1886);
nand U2139 (N_2139,N_1987,N_1815);
or U2140 (N_2140,N_1949,N_1966);
nor U2141 (N_2141,N_1986,N_1810);
nand U2142 (N_2142,N_1995,N_1883);
and U2143 (N_2143,N_1859,N_1940);
or U2144 (N_2144,N_1911,N_1998);
nand U2145 (N_2145,N_1990,N_1986);
nor U2146 (N_2146,N_1967,N_1908);
xnor U2147 (N_2147,N_1824,N_1946);
nand U2148 (N_2148,N_1893,N_1984);
nand U2149 (N_2149,N_1838,N_1837);
xor U2150 (N_2150,N_1849,N_1912);
and U2151 (N_2151,N_1981,N_1803);
or U2152 (N_2152,N_1865,N_1839);
nand U2153 (N_2153,N_1828,N_1883);
or U2154 (N_2154,N_1919,N_1984);
or U2155 (N_2155,N_1981,N_1813);
xor U2156 (N_2156,N_1974,N_1873);
and U2157 (N_2157,N_1944,N_1921);
xnor U2158 (N_2158,N_1971,N_1859);
or U2159 (N_2159,N_1813,N_1851);
or U2160 (N_2160,N_1954,N_1943);
nor U2161 (N_2161,N_1993,N_1933);
nand U2162 (N_2162,N_1863,N_1867);
xnor U2163 (N_2163,N_1913,N_1881);
and U2164 (N_2164,N_1848,N_1871);
nand U2165 (N_2165,N_1925,N_1896);
or U2166 (N_2166,N_1863,N_1816);
or U2167 (N_2167,N_1890,N_1840);
nand U2168 (N_2168,N_1860,N_1855);
nor U2169 (N_2169,N_1927,N_1888);
and U2170 (N_2170,N_1810,N_1823);
or U2171 (N_2171,N_1846,N_1869);
nor U2172 (N_2172,N_1905,N_1877);
and U2173 (N_2173,N_1812,N_1994);
or U2174 (N_2174,N_1807,N_1993);
nand U2175 (N_2175,N_1931,N_1953);
and U2176 (N_2176,N_1900,N_1884);
nor U2177 (N_2177,N_1926,N_1951);
and U2178 (N_2178,N_1869,N_1885);
xnor U2179 (N_2179,N_1803,N_1946);
nand U2180 (N_2180,N_1922,N_1992);
xor U2181 (N_2181,N_1841,N_1907);
xnor U2182 (N_2182,N_1874,N_1915);
and U2183 (N_2183,N_1853,N_1837);
nor U2184 (N_2184,N_1862,N_1968);
or U2185 (N_2185,N_1913,N_1958);
or U2186 (N_2186,N_1951,N_1906);
and U2187 (N_2187,N_1993,N_1971);
and U2188 (N_2188,N_1926,N_1960);
or U2189 (N_2189,N_1975,N_1808);
nand U2190 (N_2190,N_1947,N_1861);
nand U2191 (N_2191,N_1905,N_1850);
xnor U2192 (N_2192,N_1854,N_1871);
nand U2193 (N_2193,N_1916,N_1993);
nand U2194 (N_2194,N_1805,N_1884);
nor U2195 (N_2195,N_1853,N_1925);
nand U2196 (N_2196,N_1950,N_1844);
or U2197 (N_2197,N_1999,N_1853);
and U2198 (N_2198,N_1997,N_1918);
xnor U2199 (N_2199,N_1955,N_1832);
or U2200 (N_2200,N_2003,N_2116);
nor U2201 (N_2201,N_2112,N_2167);
or U2202 (N_2202,N_2026,N_2121);
or U2203 (N_2203,N_2045,N_2031);
nor U2204 (N_2204,N_2170,N_2155);
and U2205 (N_2205,N_2118,N_2176);
or U2206 (N_2206,N_2127,N_2133);
nor U2207 (N_2207,N_2130,N_2050);
and U2208 (N_2208,N_2110,N_2099);
xnor U2209 (N_2209,N_2069,N_2179);
nand U2210 (N_2210,N_2189,N_2135);
xnor U2211 (N_2211,N_2140,N_2108);
nor U2212 (N_2212,N_2191,N_2005);
nor U2213 (N_2213,N_2035,N_2012);
nor U2214 (N_2214,N_2101,N_2146);
nand U2215 (N_2215,N_2095,N_2122);
and U2216 (N_2216,N_2089,N_2052);
nor U2217 (N_2217,N_2180,N_2072);
xnor U2218 (N_2218,N_2196,N_2156);
nor U2219 (N_2219,N_2047,N_2150);
nor U2220 (N_2220,N_2102,N_2080);
or U2221 (N_2221,N_2165,N_2083);
or U2222 (N_2222,N_2015,N_2096);
nor U2223 (N_2223,N_2126,N_2039);
nand U2224 (N_2224,N_2004,N_2065);
and U2225 (N_2225,N_2190,N_2002);
and U2226 (N_2226,N_2000,N_2001);
nand U2227 (N_2227,N_2142,N_2182);
xnor U2228 (N_2228,N_2062,N_2006);
nand U2229 (N_2229,N_2007,N_2168);
or U2230 (N_2230,N_2107,N_2103);
nor U2231 (N_2231,N_2042,N_2061);
and U2232 (N_2232,N_2158,N_2046);
nand U2233 (N_2233,N_2022,N_2017);
nor U2234 (N_2234,N_2036,N_2100);
and U2235 (N_2235,N_2125,N_2068);
nand U2236 (N_2236,N_2136,N_2067);
or U2237 (N_2237,N_2066,N_2011);
or U2238 (N_2238,N_2051,N_2041);
nand U2239 (N_2239,N_2123,N_2178);
xor U2240 (N_2240,N_2070,N_2161);
or U2241 (N_2241,N_2145,N_2085);
and U2242 (N_2242,N_2131,N_2034);
nand U2243 (N_2243,N_2097,N_2029);
nor U2244 (N_2244,N_2027,N_2019);
xor U2245 (N_2245,N_2059,N_2128);
and U2246 (N_2246,N_2199,N_2049);
nor U2247 (N_2247,N_2166,N_2149);
or U2248 (N_2248,N_2129,N_2162);
and U2249 (N_2249,N_2093,N_2109);
xor U2250 (N_2250,N_2020,N_2030);
nand U2251 (N_2251,N_2028,N_2177);
or U2252 (N_2252,N_2138,N_2181);
and U2253 (N_2253,N_2185,N_2154);
nand U2254 (N_2254,N_2139,N_2195);
nand U2255 (N_2255,N_2198,N_2053);
nor U2256 (N_2256,N_2078,N_2064);
nor U2257 (N_2257,N_2148,N_2119);
xnor U2258 (N_2258,N_2075,N_2106);
xor U2259 (N_2259,N_2111,N_2144);
or U2260 (N_2260,N_2194,N_2160);
xor U2261 (N_2261,N_2120,N_2092);
nor U2262 (N_2262,N_2082,N_2077);
xor U2263 (N_2263,N_2117,N_2063);
and U2264 (N_2264,N_2172,N_2113);
nand U2265 (N_2265,N_2071,N_2021);
and U2266 (N_2266,N_2141,N_2009);
and U2267 (N_2267,N_2151,N_2132);
xnor U2268 (N_2268,N_2073,N_2043);
and U2269 (N_2269,N_2187,N_2137);
and U2270 (N_2270,N_2060,N_2040);
nor U2271 (N_2271,N_2054,N_2184);
and U2272 (N_2272,N_2056,N_2076);
nand U2273 (N_2273,N_2057,N_2183);
or U2274 (N_2274,N_2037,N_2171);
xnor U2275 (N_2275,N_2163,N_2164);
and U2276 (N_2276,N_2174,N_2134);
xnor U2277 (N_2277,N_2084,N_2114);
and U2278 (N_2278,N_2159,N_2008);
nor U2279 (N_2279,N_2013,N_2152);
and U2280 (N_2280,N_2094,N_2044);
nor U2281 (N_2281,N_2088,N_2157);
and U2282 (N_2282,N_2193,N_2153);
and U2283 (N_2283,N_2016,N_2147);
or U2284 (N_2284,N_2169,N_2098);
nand U2285 (N_2285,N_2086,N_2186);
nand U2286 (N_2286,N_2055,N_2115);
nor U2287 (N_2287,N_2105,N_2091);
xnor U2288 (N_2288,N_2192,N_2188);
and U2289 (N_2289,N_2023,N_2081);
or U2290 (N_2290,N_2079,N_2048);
nor U2291 (N_2291,N_2104,N_2010);
or U2292 (N_2292,N_2024,N_2175);
or U2293 (N_2293,N_2018,N_2032);
nand U2294 (N_2294,N_2014,N_2090);
or U2295 (N_2295,N_2143,N_2074);
xor U2296 (N_2296,N_2038,N_2197);
xor U2297 (N_2297,N_2025,N_2124);
nor U2298 (N_2298,N_2058,N_2087);
nor U2299 (N_2299,N_2033,N_2173);
nor U2300 (N_2300,N_2147,N_2100);
or U2301 (N_2301,N_2119,N_2010);
nor U2302 (N_2302,N_2041,N_2062);
xor U2303 (N_2303,N_2006,N_2197);
or U2304 (N_2304,N_2023,N_2044);
and U2305 (N_2305,N_2099,N_2123);
xnor U2306 (N_2306,N_2050,N_2057);
or U2307 (N_2307,N_2144,N_2185);
or U2308 (N_2308,N_2025,N_2047);
and U2309 (N_2309,N_2160,N_2193);
xnor U2310 (N_2310,N_2069,N_2143);
and U2311 (N_2311,N_2060,N_2129);
nand U2312 (N_2312,N_2131,N_2111);
nand U2313 (N_2313,N_2154,N_2065);
xor U2314 (N_2314,N_2100,N_2119);
or U2315 (N_2315,N_2155,N_2180);
and U2316 (N_2316,N_2096,N_2039);
and U2317 (N_2317,N_2059,N_2171);
nand U2318 (N_2318,N_2166,N_2187);
xnor U2319 (N_2319,N_2097,N_2108);
and U2320 (N_2320,N_2105,N_2103);
and U2321 (N_2321,N_2172,N_2019);
nand U2322 (N_2322,N_2109,N_2102);
xnor U2323 (N_2323,N_2084,N_2071);
and U2324 (N_2324,N_2181,N_2110);
or U2325 (N_2325,N_2151,N_2173);
nand U2326 (N_2326,N_2157,N_2133);
nand U2327 (N_2327,N_2149,N_2168);
nor U2328 (N_2328,N_2151,N_2139);
xnor U2329 (N_2329,N_2018,N_2157);
nand U2330 (N_2330,N_2122,N_2041);
nand U2331 (N_2331,N_2114,N_2182);
nand U2332 (N_2332,N_2111,N_2123);
xor U2333 (N_2333,N_2163,N_2158);
nor U2334 (N_2334,N_2045,N_2151);
and U2335 (N_2335,N_2069,N_2136);
nand U2336 (N_2336,N_2105,N_2016);
xnor U2337 (N_2337,N_2052,N_2167);
nor U2338 (N_2338,N_2045,N_2170);
nand U2339 (N_2339,N_2080,N_2078);
and U2340 (N_2340,N_2167,N_2069);
nand U2341 (N_2341,N_2057,N_2185);
nor U2342 (N_2342,N_2131,N_2132);
xnor U2343 (N_2343,N_2186,N_2005);
or U2344 (N_2344,N_2109,N_2070);
or U2345 (N_2345,N_2104,N_2100);
xor U2346 (N_2346,N_2096,N_2058);
nor U2347 (N_2347,N_2198,N_2159);
nand U2348 (N_2348,N_2082,N_2054);
and U2349 (N_2349,N_2011,N_2039);
xor U2350 (N_2350,N_2169,N_2087);
and U2351 (N_2351,N_2115,N_2032);
xor U2352 (N_2352,N_2105,N_2050);
or U2353 (N_2353,N_2153,N_2198);
xnor U2354 (N_2354,N_2057,N_2170);
or U2355 (N_2355,N_2115,N_2009);
or U2356 (N_2356,N_2097,N_2171);
nor U2357 (N_2357,N_2032,N_2041);
and U2358 (N_2358,N_2101,N_2108);
or U2359 (N_2359,N_2130,N_2192);
and U2360 (N_2360,N_2118,N_2004);
nor U2361 (N_2361,N_2088,N_2166);
xnor U2362 (N_2362,N_2082,N_2015);
nand U2363 (N_2363,N_2010,N_2001);
and U2364 (N_2364,N_2166,N_2195);
nor U2365 (N_2365,N_2003,N_2034);
and U2366 (N_2366,N_2031,N_2073);
nor U2367 (N_2367,N_2156,N_2005);
or U2368 (N_2368,N_2162,N_2107);
or U2369 (N_2369,N_2187,N_2087);
nor U2370 (N_2370,N_2148,N_2087);
nor U2371 (N_2371,N_2103,N_2106);
nand U2372 (N_2372,N_2131,N_2044);
nor U2373 (N_2373,N_2070,N_2000);
nand U2374 (N_2374,N_2076,N_2154);
nand U2375 (N_2375,N_2165,N_2078);
xor U2376 (N_2376,N_2085,N_2065);
xnor U2377 (N_2377,N_2022,N_2065);
nor U2378 (N_2378,N_2006,N_2183);
or U2379 (N_2379,N_2021,N_2171);
nand U2380 (N_2380,N_2090,N_2102);
nor U2381 (N_2381,N_2163,N_2049);
xor U2382 (N_2382,N_2122,N_2079);
xnor U2383 (N_2383,N_2077,N_2179);
nor U2384 (N_2384,N_2033,N_2132);
or U2385 (N_2385,N_2077,N_2038);
and U2386 (N_2386,N_2112,N_2026);
or U2387 (N_2387,N_2173,N_2163);
xnor U2388 (N_2388,N_2045,N_2122);
nor U2389 (N_2389,N_2048,N_2121);
xor U2390 (N_2390,N_2127,N_2098);
nor U2391 (N_2391,N_2042,N_2101);
and U2392 (N_2392,N_2006,N_2159);
nand U2393 (N_2393,N_2150,N_2112);
or U2394 (N_2394,N_2119,N_2174);
xnor U2395 (N_2395,N_2102,N_2196);
nor U2396 (N_2396,N_2005,N_2010);
nor U2397 (N_2397,N_2180,N_2039);
nand U2398 (N_2398,N_2185,N_2052);
and U2399 (N_2399,N_2104,N_2143);
and U2400 (N_2400,N_2325,N_2290);
nand U2401 (N_2401,N_2339,N_2269);
or U2402 (N_2402,N_2265,N_2329);
nor U2403 (N_2403,N_2291,N_2307);
nand U2404 (N_2404,N_2374,N_2341);
or U2405 (N_2405,N_2360,N_2318);
and U2406 (N_2406,N_2382,N_2228);
nor U2407 (N_2407,N_2347,N_2385);
nor U2408 (N_2408,N_2392,N_2369);
and U2409 (N_2409,N_2217,N_2313);
or U2410 (N_2410,N_2299,N_2232);
xor U2411 (N_2411,N_2306,N_2398);
nor U2412 (N_2412,N_2214,N_2233);
and U2413 (N_2413,N_2344,N_2253);
xnor U2414 (N_2414,N_2321,N_2315);
nor U2415 (N_2415,N_2272,N_2387);
nor U2416 (N_2416,N_2366,N_2292);
nand U2417 (N_2417,N_2216,N_2316);
and U2418 (N_2418,N_2367,N_2317);
xor U2419 (N_2419,N_2297,N_2305);
and U2420 (N_2420,N_2311,N_2322);
or U2421 (N_2421,N_2331,N_2391);
nor U2422 (N_2422,N_2319,N_2300);
nand U2423 (N_2423,N_2260,N_2261);
xnor U2424 (N_2424,N_2239,N_2224);
xor U2425 (N_2425,N_2264,N_2220);
and U2426 (N_2426,N_2204,N_2310);
nor U2427 (N_2427,N_2377,N_2352);
nor U2428 (N_2428,N_2263,N_2309);
and U2429 (N_2429,N_2363,N_2215);
xor U2430 (N_2430,N_2373,N_2244);
and U2431 (N_2431,N_2207,N_2255);
xnor U2432 (N_2432,N_2247,N_2288);
or U2433 (N_2433,N_2355,N_2298);
and U2434 (N_2434,N_2379,N_2296);
nor U2435 (N_2435,N_2289,N_2268);
xnor U2436 (N_2436,N_2205,N_2277);
xor U2437 (N_2437,N_2389,N_2267);
or U2438 (N_2438,N_2303,N_2249);
and U2439 (N_2439,N_2350,N_2386);
nor U2440 (N_2440,N_2237,N_2332);
and U2441 (N_2441,N_2286,N_2200);
or U2442 (N_2442,N_2294,N_2270);
nor U2443 (N_2443,N_2383,N_2257);
nand U2444 (N_2444,N_2203,N_2262);
nand U2445 (N_2445,N_2308,N_2221);
xnor U2446 (N_2446,N_2312,N_2356);
xor U2447 (N_2447,N_2376,N_2370);
nor U2448 (N_2448,N_2326,N_2304);
xnor U2449 (N_2449,N_2229,N_2397);
and U2450 (N_2450,N_2256,N_2324);
nand U2451 (N_2451,N_2372,N_2380);
nand U2452 (N_2452,N_2337,N_2285);
or U2453 (N_2453,N_2258,N_2284);
nor U2454 (N_2454,N_2276,N_2219);
or U2455 (N_2455,N_2279,N_2302);
and U2456 (N_2456,N_2314,N_2342);
nor U2457 (N_2457,N_2245,N_2371);
xnor U2458 (N_2458,N_2378,N_2362);
nand U2459 (N_2459,N_2251,N_2301);
xnor U2460 (N_2460,N_2334,N_2348);
nor U2461 (N_2461,N_2273,N_2236);
or U2462 (N_2462,N_2252,N_2240);
or U2463 (N_2463,N_2282,N_2283);
nor U2464 (N_2464,N_2340,N_2231);
nand U2465 (N_2465,N_2323,N_2234);
xnor U2466 (N_2466,N_2368,N_2343);
or U2467 (N_2467,N_2351,N_2235);
and U2468 (N_2468,N_2333,N_2238);
nand U2469 (N_2469,N_2230,N_2280);
or U2470 (N_2470,N_2211,N_2212);
and U2471 (N_2471,N_2327,N_2226);
nor U2472 (N_2472,N_2209,N_2357);
or U2473 (N_2473,N_2375,N_2393);
nor U2474 (N_2474,N_2250,N_2248);
nand U2475 (N_2475,N_2223,N_2281);
and U2476 (N_2476,N_2210,N_2243);
nor U2477 (N_2477,N_2225,N_2330);
or U2478 (N_2478,N_2274,N_2346);
xnor U2479 (N_2479,N_2395,N_2202);
xor U2480 (N_2480,N_2359,N_2328);
nor U2481 (N_2481,N_2394,N_2361);
nor U2482 (N_2482,N_2278,N_2335);
and U2483 (N_2483,N_2208,N_2388);
nand U2484 (N_2484,N_2206,N_2384);
or U2485 (N_2485,N_2242,N_2399);
or U2486 (N_2486,N_2271,N_2320);
or U2487 (N_2487,N_2390,N_2287);
or U2488 (N_2488,N_2354,N_2365);
nand U2489 (N_2489,N_2259,N_2254);
nand U2490 (N_2490,N_2381,N_2345);
or U2491 (N_2491,N_2218,N_2349);
or U2492 (N_2492,N_2293,N_2295);
or U2493 (N_2493,N_2246,N_2396);
or U2494 (N_2494,N_2241,N_2213);
or U2495 (N_2495,N_2201,N_2353);
nand U2496 (N_2496,N_2338,N_2364);
nor U2497 (N_2497,N_2336,N_2358);
or U2498 (N_2498,N_2227,N_2275);
nor U2499 (N_2499,N_2222,N_2266);
nand U2500 (N_2500,N_2360,N_2377);
and U2501 (N_2501,N_2302,N_2398);
and U2502 (N_2502,N_2211,N_2223);
and U2503 (N_2503,N_2368,N_2297);
xnor U2504 (N_2504,N_2335,N_2214);
nand U2505 (N_2505,N_2332,N_2352);
and U2506 (N_2506,N_2249,N_2277);
nor U2507 (N_2507,N_2311,N_2393);
or U2508 (N_2508,N_2273,N_2262);
and U2509 (N_2509,N_2307,N_2378);
and U2510 (N_2510,N_2229,N_2220);
nand U2511 (N_2511,N_2309,N_2380);
nor U2512 (N_2512,N_2242,N_2386);
or U2513 (N_2513,N_2281,N_2224);
nor U2514 (N_2514,N_2201,N_2348);
and U2515 (N_2515,N_2360,N_2293);
and U2516 (N_2516,N_2394,N_2297);
and U2517 (N_2517,N_2263,N_2271);
nand U2518 (N_2518,N_2379,N_2244);
xnor U2519 (N_2519,N_2298,N_2317);
nand U2520 (N_2520,N_2380,N_2331);
nand U2521 (N_2521,N_2298,N_2352);
nor U2522 (N_2522,N_2256,N_2353);
nand U2523 (N_2523,N_2343,N_2293);
xnor U2524 (N_2524,N_2328,N_2268);
and U2525 (N_2525,N_2205,N_2256);
nand U2526 (N_2526,N_2261,N_2311);
and U2527 (N_2527,N_2365,N_2244);
or U2528 (N_2528,N_2224,N_2253);
or U2529 (N_2529,N_2272,N_2230);
and U2530 (N_2530,N_2351,N_2231);
or U2531 (N_2531,N_2261,N_2319);
nand U2532 (N_2532,N_2393,N_2297);
nand U2533 (N_2533,N_2273,N_2353);
nor U2534 (N_2534,N_2212,N_2285);
and U2535 (N_2535,N_2310,N_2351);
nor U2536 (N_2536,N_2336,N_2272);
xor U2537 (N_2537,N_2365,N_2376);
nor U2538 (N_2538,N_2230,N_2321);
nand U2539 (N_2539,N_2213,N_2242);
nor U2540 (N_2540,N_2373,N_2380);
and U2541 (N_2541,N_2248,N_2210);
nor U2542 (N_2542,N_2227,N_2228);
and U2543 (N_2543,N_2262,N_2317);
xor U2544 (N_2544,N_2274,N_2341);
nand U2545 (N_2545,N_2244,N_2207);
nand U2546 (N_2546,N_2375,N_2250);
or U2547 (N_2547,N_2311,N_2375);
or U2548 (N_2548,N_2306,N_2356);
nand U2549 (N_2549,N_2335,N_2242);
and U2550 (N_2550,N_2348,N_2374);
nor U2551 (N_2551,N_2271,N_2211);
nor U2552 (N_2552,N_2286,N_2381);
xnor U2553 (N_2553,N_2211,N_2333);
or U2554 (N_2554,N_2318,N_2341);
nor U2555 (N_2555,N_2292,N_2328);
nand U2556 (N_2556,N_2233,N_2329);
or U2557 (N_2557,N_2205,N_2323);
and U2558 (N_2558,N_2206,N_2390);
nand U2559 (N_2559,N_2336,N_2399);
nor U2560 (N_2560,N_2362,N_2251);
nand U2561 (N_2561,N_2243,N_2305);
nand U2562 (N_2562,N_2348,N_2261);
nor U2563 (N_2563,N_2383,N_2295);
xnor U2564 (N_2564,N_2265,N_2253);
and U2565 (N_2565,N_2392,N_2275);
and U2566 (N_2566,N_2230,N_2316);
xor U2567 (N_2567,N_2306,N_2322);
or U2568 (N_2568,N_2207,N_2232);
nand U2569 (N_2569,N_2216,N_2350);
and U2570 (N_2570,N_2294,N_2318);
and U2571 (N_2571,N_2335,N_2259);
nand U2572 (N_2572,N_2277,N_2347);
nand U2573 (N_2573,N_2387,N_2268);
nor U2574 (N_2574,N_2229,N_2389);
or U2575 (N_2575,N_2239,N_2262);
and U2576 (N_2576,N_2255,N_2235);
nand U2577 (N_2577,N_2391,N_2299);
nor U2578 (N_2578,N_2290,N_2397);
nand U2579 (N_2579,N_2272,N_2249);
nor U2580 (N_2580,N_2224,N_2307);
nor U2581 (N_2581,N_2259,N_2251);
nor U2582 (N_2582,N_2269,N_2279);
and U2583 (N_2583,N_2346,N_2302);
nand U2584 (N_2584,N_2310,N_2292);
xor U2585 (N_2585,N_2361,N_2261);
nand U2586 (N_2586,N_2315,N_2309);
or U2587 (N_2587,N_2254,N_2396);
or U2588 (N_2588,N_2286,N_2256);
and U2589 (N_2589,N_2302,N_2305);
and U2590 (N_2590,N_2230,N_2244);
or U2591 (N_2591,N_2310,N_2215);
nand U2592 (N_2592,N_2398,N_2375);
nor U2593 (N_2593,N_2233,N_2247);
nor U2594 (N_2594,N_2358,N_2284);
or U2595 (N_2595,N_2242,N_2229);
nand U2596 (N_2596,N_2374,N_2257);
xor U2597 (N_2597,N_2234,N_2239);
nand U2598 (N_2598,N_2206,N_2236);
nand U2599 (N_2599,N_2228,N_2293);
xor U2600 (N_2600,N_2496,N_2443);
nor U2601 (N_2601,N_2599,N_2513);
and U2602 (N_2602,N_2427,N_2435);
and U2603 (N_2603,N_2503,N_2429);
xor U2604 (N_2604,N_2425,N_2400);
or U2605 (N_2605,N_2577,N_2421);
nor U2606 (N_2606,N_2420,N_2520);
and U2607 (N_2607,N_2511,N_2477);
and U2608 (N_2608,N_2542,N_2475);
nor U2609 (N_2609,N_2414,N_2498);
nand U2610 (N_2610,N_2521,N_2406);
or U2611 (N_2611,N_2438,N_2573);
nor U2612 (N_2612,N_2556,N_2537);
or U2613 (N_2613,N_2489,N_2452);
nor U2614 (N_2614,N_2541,N_2555);
xor U2615 (N_2615,N_2418,N_2433);
and U2616 (N_2616,N_2422,N_2572);
nor U2617 (N_2617,N_2579,N_2562);
or U2618 (N_2618,N_2479,N_2592);
nand U2619 (N_2619,N_2545,N_2580);
or U2620 (N_2620,N_2597,N_2461);
nand U2621 (N_2621,N_2410,N_2539);
or U2622 (N_2622,N_2527,N_2500);
nor U2623 (N_2623,N_2446,N_2561);
or U2624 (N_2624,N_2459,N_2423);
nand U2625 (N_2625,N_2499,N_2486);
or U2626 (N_2626,N_2581,N_2462);
nor U2627 (N_2627,N_2440,N_2432);
xnor U2628 (N_2628,N_2550,N_2492);
or U2629 (N_2629,N_2405,N_2557);
nor U2630 (N_2630,N_2518,N_2549);
nand U2631 (N_2631,N_2442,N_2566);
nor U2632 (N_2632,N_2578,N_2588);
xnor U2633 (N_2633,N_2428,N_2554);
xnor U2634 (N_2634,N_2403,N_2582);
and U2635 (N_2635,N_2487,N_2531);
nor U2636 (N_2636,N_2546,N_2424);
or U2637 (N_2637,N_2510,N_2548);
nor U2638 (N_2638,N_2483,N_2449);
nand U2639 (N_2639,N_2434,N_2552);
or U2640 (N_2640,N_2468,N_2538);
xor U2641 (N_2641,N_2476,N_2463);
and U2642 (N_2642,N_2575,N_2493);
xor U2643 (N_2643,N_2466,N_2517);
xor U2644 (N_2644,N_2570,N_2441);
nand U2645 (N_2645,N_2519,N_2530);
or U2646 (N_2646,N_2535,N_2485);
or U2647 (N_2647,N_2504,N_2586);
and U2648 (N_2648,N_2506,N_2482);
or U2649 (N_2649,N_2437,N_2471);
or U2650 (N_2650,N_2591,N_2419);
nor U2651 (N_2651,N_2457,N_2563);
xor U2652 (N_2652,N_2407,N_2553);
and U2653 (N_2653,N_2560,N_2516);
and U2654 (N_2654,N_2491,N_2514);
or U2655 (N_2655,N_2484,N_2447);
nand U2656 (N_2656,N_2544,N_2455);
nand U2657 (N_2657,N_2559,N_2430);
nor U2658 (N_2658,N_2533,N_2590);
xor U2659 (N_2659,N_2456,N_2416);
nor U2660 (N_2660,N_2401,N_2569);
xnor U2661 (N_2661,N_2558,N_2509);
nand U2662 (N_2662,N_2480,N_2412);
xor U2663 (N_2663,N_2565,N_2417);
nor U2664 (N_2664,N_2502,N_2547);
xor U2665 (N_2665,N_2584,N_2598);
and U2666 (N_2666,N_2488,N_2522);
and U2667 (N_2667,N_2505,N_2585);
or U2668 (N_2668,N_2472,N_2583);
nor U2669 (N_2669,N_2564,N_2478);
xor U2670 (N_2670,N_2495,N_2543);
nand U2671 (N_2671,N_2460,N_2523);
and U2672 (N_2672,N_2574,N_2587);
xnor U2673 (N_2673,N_2413,N_2551);
xor U2674 (N_2674,N_2453,N_2567);
and U2675 (N_2675,N_2431,N_2451);
nor U2676 (N_2676,N_2409,N_2494);
nand U2677 (N_2677,N_2444,N_2529);
nand U2678 (N_2678,N_2571,N_2404);
and U2679 (N_2679,N_2445,N_2454);
or U2680 (N_2680,N_2540,N_2426);
or U2681 (N_2681,N_2402,N_2525);
or U2682 (N_2682,N_2458,N_2526);
or U2683 (N_2683,N_2595,N_2464);
or U2684 (N_2684,N_2497,N_2436);
xor U2685 (N_2685,N_2450,N_2439);
xnor U2686 (N_2686,N_2524,N_2490);
nor U2687 (N_2687,N_2532,N_2415);
nand U2688 (N_2688,N_2528,N_2508);
xor U2689 (N_2689,N_2512,N_2473);
and U2690 (N_2690,N_2474,N_2589);
nand U2691 (N_2691,N_2408,N_2515);
nor U2692 (N_2692,N_2536,N_2470);
or U2693 (N_2693,N_2467,N_2596);
or U2694 (N_2694,N_2534,N_2469);
or U2695 (N_2695,N_2576,N_2448);
nor U2696 (N_2696,N_2507,N_2593);
nand U2697 (N_2697,N_2568,N_2481);
or U2698 (N_2698,N_2411,N_2465);
and U2699 (N_2699,N_2594,N_2501);
or U2700 (N_2700,N_2435,N_2470);
nand U2701 (N_2701,N_2437,N_2562);
nand U2702 (N_2702,N_2505,N_2438);
xor U2703 (N_2703,N_2597,N_2435);
nand U2704 (N_2704,N_2448,N_2525);
or U2705 (N_2705,N_2403,N_2446);
nor U2706 (N_2706,N_2458,N_2475);
nor U2707 (N_2707,N_2434,N_2562);
nand U2708 (N_2708,N_2462,N_2571);
nand U2709 (N_2709,N_2442,N_2501);
and U2710 (N_2710,N_2410,N_2438);
or U2711 (N_2711,N_2402,N_2562);
and U2712 (N_2712,N_2441,N_2505);
xnor U2713 (N_2713,N_2481,N_2551);
xor U2714 (N_2714,N_2554,N_2537);
and U2715 (N_2715,N_2520,N_2507);
nor U2716 (N_2716,N_2546,N_2410);
and U2717 (N_2717,N_2462,N_2533);
xor U2718 (N_2718,N_2451,N_2488);
and U2719 (N_2719,N_2404,N_2523);
nand U2720 (N_2720,N_2452,N_2439);
or U2721 (N_2721,N_2596,N_2468);
xnor U2722 (N_2722,N_2526,N_2478);
and U2723 (N_2723,N_2544,N_2498);
and U2724 (N_2724,N_2405,N_2506);
and U2725 (N_2725,N_2496,N_2504);
xnor U2726 (N_2726,N_2511,N_2510);
and U2727 (N_2727,N_2438,N_2491);
and U2728 (N_2728,N_2406,N_2430);
and U2729 (N_2729,N_2423,N_2584);
nand U2730 (N_2730,N_2454,N_2582);
xnor U2731 (N_2731,N_2484,N_2439);
nand U2732 (N_2732,N_2441,N_2410);
or U2733 (N_2733,N_2505,N_2448);
or U2734 (N_2734,N_2522,N_2489);
and U2735 (N_2735,N_2578,N_2430);
nand U2736 (N_2736,N_2406,N_2490);
or U2737 (N_2737,N_2551,N_2425);
xor U2738 (N_2738,N_2564,N_2475);
xor U2739 (N_2739,N_2443,N_2426);
or U2740 (N_2740,N_2433,N_2406);
nand U2741 (N_2741,N_2461,N_2514);
and U2742 (N_2742,N_2459,N_2446);
nor U2743 (N_2743,N_2517,N_2599);
nor U2744 (N_2744,N_2545,N_2558);
or U2745 (N_2745,N_2593,N_2453);
and U2746 (N_2746,N_2468,N_2561);
xor U2747 (N_2747,N_2510,N_2525);
nand U2748 (N_2748,N_2518,N_2532);
nor U2749 (N_2749,N_2468,N_2545);
nand U2750 (N_2750,N_2551,N_2538);
and U2751 (N_2751,N_2442,N_2429);
xor U2752 (N_2752,N_2557,N_2453);
xnor U2753 (N_2753,N_2529,N_2518);
nor U2754 (N_2754,N_2414,N_2547);
xor U2755 (N_2755,N_2515,N_2434);
or U2756 (N_2756,N_2588,N_2429);
and U2757 (N_2757,N_2529,N_2509);
xnor U2758 (N_2758,N_2437,N_2519);
and U2759 (N_2759,N_2417,N_2534);
and U2760 (N_2760,N_2416,N_2525);
or U2761 (N_2761,N_2543,N_2535);
xor U2762 (N_2762,N_2440,N_2580);
nor U2763 (N_2763,N_2586,N_2479);
and U2764 (N_2764,N_2518,N_2531);
nor U2765 (N_2765,N_2523,N_2585);
nor U2766 (N_2766,N_2481,N_2537);
or U2767 (N_2767,N_2418,N_2456);
and U2768 (N_2768,N_2559,N_2533);
and U2769 (N_2769,N_2559,N_2588);
xor U2770 (N_2770,N_2513,N_2497);
or U2771 (N_2771,N_2444,N_2478);
and U2772 (N_2772,N_2480,N_2576);
nand U2773 (N_2773,N_2466,N_2492);
or U2774 (N_2774,N_2515,N_2524);
and U2775 (N_2775,N_2535,N_2462);
and U2776 (N_2776,N_2424,N_2574);
xor U2777 (N_2777,N_2521,N_2522);
or U2778 (N_2778,N_2557,N_2460);
and U2779 (N_2779,N_2515,N_2441);
or U2780 (N_2780,N_2520,N_2436);
xnor U2781 (N_2781,N_2401,N_2426);
xor U2782 (N_2782,N_2500,N_2588);
xnor U2783 (N_2783,N_2462,N_2402);
and U2784 (N_2784,N_2521,N_2421);
and U2785 (N_2785,N_2494,N_2448);
or U2786 (N_2786,N_2598,N_2443);
and U2787 (N_2787,N_2599,N_2582);
xor U2788 (N_2788,N_2502,N_2540);
or U2789 (N_2789,N_2434,N_2430);
xnor U2790 (N_2790,N_2483,N_2528);
nor U2791 (N_2791,N_2554,N_2524);
nor U2792 (N_2792,N_2437,N_2402);
xor U2793 (N_2793,N_2476,N_2581);
nand U2794 (N_2794,N_2583,N_2491);
nand U2795 (N_2795,N_2558,N_2506);
xnor U2796 (N_2796,N_2596,N_2510);
or U2797 (N_2797,N_2529,N_2590);
and U2798 (N_2798,N_2551,N_2455);
nand U2799 (N_2799,N_2419,N_2402);
or U2800 (N_2800,N_2698,N_2780);
nand U2801 (N_2801,N_2776,N_2653);
nor U2802 (N_2802,N_2729,N_2759);
nand U2803 (N_2803,N_2721,N_2710);
nor U2804 (N_2804,N_2766,N_2662);
xor U2805 (N_2805,N_2643,N_2799);
and U2806 (N_2806,N_2788,N_2702);
or U2807 (N_2807,N_2727,N_2618);
nand U2808 (N_2808,N_2623,N_2775);
or U2809 (N_2809,N_2751,N_2650);
nor U2810 (N_2810,N_2703,N_2708);
and U2811 (N_2811,N_2683,N_2648);
xor U2812 (N_2812,N_2691,N_2634);
nor U2813 (N_2813,N_2645,N_2677);
and U2814 (N_2814,N_2616,N_2668);
xor U2815 (N_2815,N_2633,N_2709);
and U2816 (N_2816,N_2654,N_2744);
and U2817 (N_2817,N_2635,N_2608);
xnor U2818 (N_2818,N_2606,N_2646);
nor U2819 (N_2819,N_2605,N_2636);
nand U2820 (N_2820,N_2725,N_2738);
nor U2821 (N_2821,N_2764,N_2601);
nand U2822 (N_2822,N_2724,N_2617);
xor U2823 (N_2823,N_2745,N_2620);
xor U2824 (N_2824,N_2789,N_2656);
nand U2825 (N_2825,N_2626,N_2660);
and U2826 (N_2826,N_2768,N_2701);
xnor U2827 (N_2827,N_2673,N_2795);
and U2828 (N_2828,N_2659,N_2749);
and U2829 (N_2829,N_2640,N_2675);
or U2830 (N_2830,N_2637,N_2732);
xnor U2831 (N_2831,N_2603,N_2609);
xor U2832 (N_2832,N_2647,N_2624);
or U2833 (N_2833,N_2705,N_2733);
or U2834 (N_2834,N_2782,N_2737);
nand U2835 (N_2835,N_2771,N_2706);
xnor U2836 (N_2836,N_2684,N_2607);
nor U2837 (N_2837,N_2792,N_2719);
and U2838 (N_2838,N_2786,N_2754);
or U2839 (N_2839,N_2629,N_2704);
xnor U2840 (N_2840,N_2652,N_2611);
xor U2841 (N_2841,N_2685,N_2730);
xor U2842 (N_2842,N_2707,N_2641);
nor U2843 (N_2843,N_2723,N_2682);
xor U2844 (N_2844,N_2794,N_2734);
nor U2845 (N_2845,N_2664,N_2755);
nand U2846 (N_2846,N_2665,N_2696);
nor U2847 (N_2847,N_2763,N_2644);
nor U2848 (N_2848,N_2663,N_2791);
or U2849 (N_2849,N_2674,N_2772);
nor U2850 (N_2850,N_2672,N_2686);
and U2851 (N_2851,N_2630,N_2785);
and U2852 (N_2852,N_2639,N_2642);
or U2853 (N_2853,N_2657,N_2742);
or U2854 (N_2854,N_2739,N_2761);
or U2855 (N_2855,N_2676,N_2767);
or U2856 (N_2856,N_2613,N_2666);
nor U2857 (N_2857,N_2602,N_2714);
xnor U2858 (N_2858,N_2681,N_2715);
and U2859 (N_2859,N_2712,N_2697);
and U2860 (N_2860,N_2790,N_2756);
or U2861 (N_2861,N_2655,N_2713);
or U2862 (N_2862,N_2753,N_2781);
nor U2863 (N_2863,N_2778,N_2765);
xor U2864 (N_2864,N_2787,N_2651);
xnor U2865 (N_2865,N_2774,N_2770);
or U2866 (N_2866,N_2622,N_2614);
or U2867 (N_2867,N_2793,N_2746);
xnor U2868 (N_2868,N_2671,N_2798);
nand U2869 (N_2869,N_2638,N_2680);
xnor U2870 (N_2870,N_2649,N_2760);
nor U2871 (N_2871,N_2699,N_2688);
and U2872 (N_2872,N_2718,N_2726);
and U2873 (N_2873,N_2783,N_2621);
xor U2874 (N_2874,N_2731,N_2690);
xnor U2875 (N_2875,N_2695,N_2700);
and U2876 (N_2876,N_2604,N_2658);
xor U2877 (N_2877,N_2625,N_2758);
and U2878 (N_2878,N_2741,N_2736);
xnor U2879 (N_2879,N_2716,N_2612);
and U2880 (N_2880,N_2693,N_2735);
nor U2881 (N_2881,N_2757,N_2694);
or U2882 (N_2882,N_2687,N_2762);
or U2883 (N_2883,N_2670,N_2669);
xor U2884 (N_2884,N_2720,N_2769);
or U2885 (N_2885,N_2619,N_2747);
or U2886 (N_2886,N_2740,N_2784);
nor U2887 (N_2887,N_2711,N_2692);
or U2888 (N_2888,N_2717,N_2627);
and U2889 (N_2889,N_2632,N_2631);
nand U2890 (N_2890,N_2678,N_2667);
nand U2891 (N_2891,N_2779,N_2752);
or U2892 (N_2892,N_2743,N_2628);
or U2893 (N_2893,N_2722,N_2748);
or U2894 (N_2894,N_2679,N_2796);
nand U2895 (N_2895,N_2610,N_2773);
nand U2896 (N_2896,N_2777,N_2750);
xor U2897 (N_2897,N_2600,N_2728);
xor U2898 (N_2898,N_2797,N_2661);
and U2899 (N_2899,N_2615,N_2689);
xor U2900 (N_2900,N_2743,N_2660);
xor U2901 (N_2901,N_2735,N_2780);
nand U2902 (N_2902,N_2773,N_2752);
xnor U2903 (N_2903,N_2732,N_2769);
or U2904 (N_2904,N_2700,N_2649);
and U2905 (N_2905,N_2767,N_2710);
xnor U2906 (N_2906,N_2625,N_2709);
nand U2907 (N_2907,N_2675,N_2652);
xnor U2908 (N_2908,N_2664,N_2645);
or U2909 (N_2909,N_2750,N_2633);
nor U2910 (N_2910,N_2720,N_2652);
nor U2911 (N_2911,N_2700,N_2709);
and U2912 (N_2912,N_2744,N_2643);
xor U2913 (N_2913,N_2777,N_2604);
xor U2914 (N_2914,N_2716,N_2721);
or U2915 (N_2915,N_2604,N_2687);
or U2916 (N_2916,N_2752,N_2665);
nand U2917 (N_2917,N_2792,N_2687);
nand U2918 (N_2918,N_2616,N_2676);
and U2919 (N_2919,N_2646,N_2635);
or U2920 (N_2920,N_2737,N_2755);
nor U2921 (N_2921,N_2687,N_2667);
nand U2922 (N_2922,N_2753,N_2682);
and U2923 (N_2923,N_2729,N_2685);
nor U2924 (N_2924,N_2702,N_2620);
nand U2925 (N_2925,N_2653,N_2684);
and U2926 (N_2926,N_2692,N_2715);
nor U2927 (N_2927,N_2616,N_2639);
xor U2928 (N_2928,N_2754,N_2725);
or U2929 (N_2929,N_2763,N_2679);
or U2930 (N_2930,N_2656,N_2710);
and U2931 (N_2931,N_2738,N_2636);
xnor U2932 (N_2932,N_2756,N_2784);
nand U2933 (N_2933,N_2781,N_2709);
nand U2934 (N_2934,N_2715,N_2745);
nor U2935 (N_2935,N_2727,N_2689);
nand U2936 (N_2936,N_2745,N_2796);
or U2937 (N_2937,N_2625,N_2686);
and U2938 (N_2938,N_2725,N_2632);
xnor U2939 (N_2939,N_2656,N_2750);
or U2940 (N_2940,N_2683,N_2741);
and U2941 (N_2941,N_2732,N_2602);
nand U2942 (N_2942,N_2736,N_2785);
nor U2943 (N_2943,N_2753,N_2617);
xor U2944 (N_2944,N_2798,N_2794);
xor U2945 (N_2945,N_2744,N_2659);
nor U2946 (N_2946,N_2655,N_2721);
nand U2947 (N_2947,N_2653,N_2702);
xor U2948 (N_2948,N_2684,N_2783);
nor U2949 (N_2949,N_2630,N_2699);
or U2950 (N_2950,N_2761,N_2622);
and U2951 (N_2951,N_2779,N_2754);
or U2952 (N_2952,N_2783,N_2711);
or U2953 (N_2953,N_2654,N_2632);
or U2954 (N_2954,N_2726,N_2772);
nand U2955 (N_2955,N_2704,N_2651);
xor U2956 (N_2956,N_2664,N_2765);
and U2957 (N_2957,N_2763,N_2738);
and U2958 (N_2958,N_2793,N_2622);
nand U2959 (N_2959,N_2636,N_2633);
nand U2960 (N_2960,N_2734,N_2609);
and U2961 (N_2961,N_2686,N_2726);
or U2962 (N_2962,N_2693,N_2663);
and U2963 (N_2963,N_2776,N_2711);
xnor U2964 (N_2964,N_2697,N_2784);
or U2965 (N_2965,N_2651,N_2682);
or U2966 (N_2966,N_2758,N_2744);
nand U2967 (N_2967,N_2789,N_2711);
and U2968 (N_2968,N_2702,N_2731);
or U2969 (N_2969,N_2712,N_2726);
or U2970 (N_2970,N_2690,N_2644);
nor U2971 (N_2971,N_2676,N_2780);
and U2972 (N_2972,N_2687,N_2705);
nand U2973 (N_2973,N_2680,N_2688);
nor U2974 (N_2974,N_2718,N_2723);
or U2975 (N_2975,N_2700,N_2606);
xnor U2976 (N_2976,N_2619,N_2679);
and U2977 (N_2977,N_2624,N_2728);
or U2978 (N_2978,N_2787,N_2786);
xor U2979 (N_2979,N_2668,N_2643);
and U2980 (N_2980,N_2691,N_2666);
xor U2981 (N_2981,N_2744,N_2756);
and U2982 (N_2982,N_2668,N_2628);
or U2983 (N_2983,N_2786,N_2772);
nor U2984 (N_2984,N_2646,N_2695);
nand U2985 (N_2985,N_2719,N_2698);
and U2986 (N_2986,N_2633,N_2645);
and U2987 (N_2987,N_2645,N_2669);
and U2988 (N_2988,N_2745,N_2691);
nand U2989 (N_2989,N_2667,N_2750);
xnor U2990 (N_2990,N_2622,N_2768);
and U2991 (N_2991,N_2788,N_2715);
xor U2992 (N_2992,N_2763,N_2689);
nor U2993 (N_2993,N_2670,N_2724);
xnor U2994 (N_2994,N_2744,N_2764);
or U2995 (N_2995,N_2632,N_2739);
or U2996 (N_2996,N_2732,N_2748);
nor U2997 (N_2997,N_2760,N_2646);
nand U2998 (N_2998,N_2760,N_2609);
xor U2999 (N_2999,N_2602,N_2797);
and U3000 (N_3000,N_2984,N_2904);
and U3001 (N_3001,N_2851,N_2919);
and U3002 (N_3002,N_2835,N_2921);
or U3003 (N_3003,N_2867,N_2970);
nand U3004 (N_3004,N_2979,N_2838);
nand U3005 (N_3005,N_2840,N_2988);
xor U3006 (N_3006,N_2866,N_2998);
nor U3007 (N_3007,N_2828,N_2910);
nor U3008 (N_3008,N_2994,N_2961);
xnor U3009 (N_3009,N_2923,N_2848);
xnor U3010 (N_3010,N_2981,N_2876);
or U3011 (N_3011,N_2859,N_2858);
xnor U3012 (N_3012,N_2800,N_2845);
xnor U3013 (N_3013,N_2999,N_2992);
nand U3014 (N_3014,N_2829,N_2985);
or U3015 (N_3015,N_2802,N_2882);
nor U3016 (N_3016,N_2817,N_2836);
nand U3017 (N_3017,N_2839,N_2930);
nand U3018 (N_3018,N_2831,N_2844);
nand U3019 (N_3019,N_2947,N_2865);
nand U3020 (N_3020,N_2819,N_2911);
nor U3021 (N_3021,N_2812,N_2937);
nand U3022 (N_3022,N_2815,N_2962);
nor U3023 (N_3023,N_2888,N_2933);
nor U3024 (N_3024,N_2920,N_2833);
xor U3025 (N_3025,N_2901,N_2890);
or U3026 (N_3026,N_2931,N_2906);
or U3027 (N_3027,N_2908,N_2941);
or U3028 (N_3028,N_2944,N_2991);
nand U3029 (N_3029,N_2913,N_2987);
nor U3030 (N_3030,N_2965,N_2932);
xor U3031 (N_3031,N_2915,N_2873);
or U3032 (N_3032,N_2943,N_2814);
or U3033 (N_3033,N_2874,N_2816);
and U3034 (N_3034,N_2942,N_2973);
nand U3035 (N_3035,N_2898,N_2824);
or U3036 (N_3036,N_2891,N_2966);
or U3037 (N_3037,N_2989,N_2903);
and U3038 (N_3038,N_2870,N_2804);
or U3039 (N_3039,N_2995,N_2878);
xnor U3040 (N_3040,N_2809,N_2905);
and U3041 (N_3041,N_2823,N_2886);
nand U3042 (N_3042,N_2821,N_2883);
nor U3043 (N_3043,N_2830,N_2952);
or U3044 (N_3044,N_2955,N_2801);
xnor U3045 (N_3045,N_2875,N_2841);
nand U3046 (N_3046,N_2860,N_2949);
and U3047 (N_3047,N_2916,N_2813);
and U3048 (N_3048,N_2900,N_2959);
nor U3049 (N_3049,N_2997,N_2894);
nor U3050 (N_3050,N_2971,N_2986);
and U3051 (N_3051,N_2934,N_2917);
or U3052 (N_3052,N_2884,N_2951);
nor U3053 (N_3053,N_2918,N_2850);
nand U3054 (N_3054,N_2837,N_2803);
and U3055 (N_3055,N_2869,N_2857);
nor U3056 (N_3056,N_2826,N_2963);
xnor U3057 (N_3057,N_2902,N_2895);
xnor U3058 (N_3058,N_2983,N_2909);
nor U3059 (N_3059,N_2864,N_2974);
nor U3060 (N_3060,N_2810,N_2877);
and U3061 (N_3061,N_2927,N_2928);
nor U3062 (N_3062,N_2868,N_2855);
or U3063 (N_3063,N_2982,N_2948);
or U3064 (N_3064,N_2842,N_2935);
and U3065 (N_3065,N_2912,N_2972);
and U3066 (N_3066,N_2968,N_2940);
nor U3067 (N_3067,N_2957,N_2827);
or U3068 (N_3068,N_2976,N_2846);
and U3069 (N_3069,N_2945,N_2881);
xor U3070 (N_3070,N_2825,N_2978);
xor U3071 (N_3071,N_2980,N_2853);
or U3072 (N_3072,N_2924,N_2849);
nor U3073 (N_3073,N_2922,N_2892);
and U3074 (N_3074,N_2852,N_2960);
and U3075 (N_3075,N_2863,N_2862);
and U3076 (N_3076,N_2897,N_2977);
nor U3077 (N_3077,N_2808,N_2899);
and U3078 (N_3078,N_2954,N_2969);
nand U3079 (N_3079,N_2996,N_2811);
xnor U3080 (N_3080,N_2914,N_2889);
nor U3081 (N_3081,N_2893,N_2926);
xnor U3082 (N_3082,N_2990,N_2818);
nor U3083 (N_3083,N_2807,N_2929);
or U3084 (N_3084,N_2856,N_2975);
nor U3085 (N_3085,N_2847,N_2925);
nor U3086 (N_3086,N_2871,N_2967);
xor U3087 (N_3087,N_2854,N_2956);
nand U3088 (N_3088,N_2806,N_2885);
or U3089 (N_3089,N_2939,N_2936);
xnor U3090 (N_3090,N_2832,N_2953);
nand U3091 (N_3091,N_2820,N_2861);
and U3092 (N_3092,N_2938,N_2907);
nor U3093 (N_3093,N_2887,N_2993);
xor U3094 (N_3094,N_2950,N_2958);
nor U3095 (N_3095,N_2880,N_2896);
nand U3096 (N_3096,N_2879,N_2872);
or U3097 (N_3097,N_2843,N_2946);
or U3098 (N_3098,N_2964,N_2805);
and U3099 (N_3099,N_2834,N_2822);
xor U3100 (N_3100,N_2832,N_2959);
nor U3101 (N_3101,N_2859,N_2907);
xor U3102 (N_3102,N_2856,N_2916);
xnor U3103 (N_3103,N_2954,N_2940);
and U3104 (N_3104,N_2930,N_2829);
nor U3105 (N_3105,N_2909,N_2968);
or U3106 (N_3106,N_2859,N_2886);
and U3107 (N_3107,N_2949,N_2974);
xor U3108 (N_3108,N_2830,N_2888);
and U3109 (N_3109,N_2840,N_2995);
nor U3110 (N_3110,N_2856,N_2927);
xor U3111 (N_3111,N_2981,N_2810);
and U3112 (N_3112,N_2850,N_2879);
nand U3113 (N_3113,N_2813,N_2883);
or U3114 (N_3114,N_2868,N_2979);
nand U3115 (N_3115,N_2869,N_2811);
xnor U3116 (N_3116,N_2950,N_2979);
nand U3117 (N_3117,N_2820,N_2980);
nor U3118 (N_3118,N_2930,N_2981);
or U3119 (N_3119,N_2860,N_2982);
nor U3120 (N_3120,N_2916,N_2846);
nor U3121 (N_3121,N_2960,N_2972);
nor U3122 (N_3122,N_2921,N_2977);
and U3123 (N_3123,N_2880,N_2835);
nor U3124 (N_3124,N_2891,N_2962);
nor U3125 (N_3125,N_2881,N_2853);
xnor U3126 (N_3126,N_2977,N_2944);
nor U3127 (N_3127,N_2952,N_2938);
and U3128 (N_3128,N_2868,N_2898);
and U3129 (N_3129,N_2838,N_2816);
and U3130 (N_3130,N_2928,N_2979);
nor U3131 (N_3131,N_2993,N_2975);
nor U3132 (N_3132,N_2813,N_2885);
xnor U3133 (N_3133,N_2866,N_2950);
nand U3134 (N_3134,N_2968,N_2848);
or U3135 (N_3135,N_2985,N_2941);
xor U3136 (N_3136,N_2883,N_2805);
xnor U3137 (N_3137,N_2954,N_2955);
nand U3138 (N_3138,N_2896,N_2898);
nor U3139 (N_3139,N_2810,N_2813);
nand U3140 (N_3140,N_2883,N_2824);
xnor U3141 (N_3141,N_2999,N_2897);
xor U3142 (N_3142,N_2800,N_2906);
nor U3143 (N_3143,N_2884,N_2838);
xor U3144 (N_3144,N_2957,N_2869);
nor U3145 (N_3145,N_2990,N_2941);
nand U3146 (N_3146,N_2936,N_2965);
xor U3147 (N_3147,N_2980,N_2817);
nor U3148 (N_3148,N_2870,N_2957);
nor U3149 (N_3149,N_2916,N_2885);
nand U3150 (N_3150,N_2875,N_2923);
nand U3151 (N_3151,N_2809,N_2983);
xnor U3152 (N_3152,N_2921,N_2975);
or U3153 (N_3153,N_2809,N_2964);
xor U3154 (N_3154,N_2813,N_2889);
and U3155 (N_3155,N_2819,N_2979);
and U3156 (N_3156,N_2899,N_2914);
nand U3157 (N_3157,N_2989,N_2847);
xnor U3158 (N_3158,N_2937,N_2953);
xnor U3159 (N_3159,N_2836,N_2826);
nand U3160 (N_3160,N_2809,N_2837);
nor U3161 (N_3161,N_2967,N_2912);
nand U3162 (N_3162,N_2860,N_2820);
and U3163 (N_3163,N_2891,N_2827);
nand U3164 (N_3164,N_2829,N_2986);
or U3165 (N_3165,N_2849,N_2936);
or U3166 (N_3166,N_2935,N_2912);
nor U3167 (N_3167,N_2894,N_2926);
xnor U3168 (N_3168,N_2898,N_2880);
xor U3169 (N_3169,N_2920,N_2868);
nand U3170 (N_3170,N_2872,N_2920);
or U3171 (N_3171,N_2962,N_2884);
xnor U3172 (N_3172,N_2843,N_2881);
nand U3173 (N_3173,N_2908,N_2925);
xnor U3174 (N_3174,N_2820,N_2910);
or U3175 (N_3175,N_2920,N_2847);
and U3176 (N_3176,N_2941,N_2923);
xnor U3177 (N_3177,N_2815,N_2960);
nand U3178 (N_3178,N_2984,N_2934);
and U3179 (N_3179,N_2835,N_2883);
nand U3180 (N_3180,N_2812,N_2899);
nor U3181 (N_3181,N_2858,N_2973);
or U3182 (N_3182,N_2805,N_2979);
nor U3183 (N_3183,N_2863,N_2811);
nor U3184 (N_3184,N_2807,N_2874);
nand U3185 (N_3185,N_2879,N_2807);
and U3186 (N_3186,N_2988,N_2998);
or U3187 (N_3187,N_2960,N_2929);
and U3188 (N_3188,N_2978,N_2913);
nand U3189 (N_3189,N_2939,N_2965);
xor U3190 (N_3190,N_2848,N_2810);
and U3191 (N_3191,N_2859,N_2956);
xor U3192 (N_3192,N_2880,N_2839);
nand U3193 (N_3193,N_2909,N_2894);
nand U3194 (N_3194,N_2974,N_2963);
and U3195 (N_3195,N_2861,N_2977);
xor U3196 (N_3196,N_2855,N_2916);
nor U3197 (N_3197,N_2962,N_2812);
nand U3198 (N_3198,N_2845,N_2935);
xor U3199 (N_3199,N_2863,N_2870);
and U3200 (N_3200,N_3034,N_3145);
nor U3201 (N_3201,N_3055,N_3048);
nor U3202 (N_3202,N_3190,N_3119);
and U3203 (N_3203,N_3180,N_3162);
nor U3204 (N_3204,N_3142,N_3179);
xor U3205 (N_3205,N_3030,N_3023);
and U3206 (N_3206,N_3136,N_3068);
and U3207 (N_3207,N_3133,N_3026);
xnor U3208 (N_3208,N_3138,N_3005);
or U3209 (N_3209,N_3065,N_3058);
nand U3210 (N_3210,N_3094,N_3092);
nor U3211 (N_3211,N_3012,N_3175);
nor U3212 (N_3212,N_3010,N_3037);
xnor U3213 (N_3213,N_3118,N_3062);
or U3214 (N_3214,N_3041,N_3036);
nor U3215 (N_3215,N_3021,N_3165);
nor U3216 (N_3216,N_3115,N_3053);
and U3217 (N_3217,N_3131,N_3150);
nor U3218 (N_3218,N_3097,N_3069);
and U3219 (N_3219,N_3017,N_3122);
and U3220 (N_3220,N_3160,N_3124);
and U3221 (N_3221,N_3089,N_3176);
and U3222 (N_3222,N_3170,N_3045);
or U3223 (N_3223,N_3066,N_3099);
nand U3224 (N_3224,N_3128,N_3006);
nand U3225 (N_3225,N_3171,N_3156);
nand U3226 (N_3226,N_3052,N_3117);
xor U3227 (N_3227,N_3166,N_3109);
nor U3228 (N_3228,N_3191,N_3051);
or U3229 (N_3229,N_3095,N_3152);
and U3230 (N_3230,N_3046,N_3087);
or U3231 (N_3231,N_3147,N_3125);
nor U3232 (N_3232,N_3072,N_3009);
xor U3233 (N_3233,N_3135,N_3003);
or U3234 (N_3234,N_3144,N_3085);
and U3235 (N_3235,N_3088,N_3093);
nor U3236 (N_3236,N_3137,N_3130);
and U3237 (N_3237,N_3127,N_3015);
nor U3238 (N_3238,N_3004,N_3000);
xnor U3239 (N_3239,N_3129,N_3140);
and U3240 (N_3240,N_3159,N_3107);
nand U3241 (N_3241,N_3164,N_3047);
xnor U3242 (N_3242,N_3103,N_3054);
or U3243 (N_3243,N_3100,N_3035);
xnor U3244 (N_3244,N_3077,N_3024);
xnor U3245 (N_3245,N_3078,N_3187);
xor U3246 (N_3246,N_3032,N_3161);
xor U3247 (N_3247,N_3007,N_3090);
nor U3248 (N_3248,N_3141,N_3192);
nand U3249 (N_3249,N_3033,N_3020);
and U3250 (N_3250,N_3168,N_3173);
and U3251 (N_3251,N_3148,N_3183);
nand U3252 (N_3252,N_3126,N_3178);
xor U3253 (N_3253,N_3157,N_3081);
nand U3254 (N_3254,N_3027,N_3114);
and U3255 (N_3255,N_3070,N_3080);
or U3256 (N_3256,N_3182,N_3086);
nand U3257 (N_3257,N_3177,N_3057);
nand U3258 (N_3258,N_3013,N_3056);
and U3259 (N_3259,N_3043,N_3050);
nor U3260 (N_3260,N_3042,N_3084);
xor U3261 (N_3261,N_3174,N_3016);
or U3262 (N_3262,N_3181,N_3172);
nand U3263 (N_3263,N_3038,N_3031);
nand U3264 (N_3264,N_3146,N_3059);
nor U3265 (N_3265,N_3132,N_3195);
and U3266 (N_3266,N_3101,N_3002);
xor U3267 (N_3267,N_3096,N_3075);
nor U3268 (N_3268,N_3102,N_3083);
or U3269 (N_3269,N_3149,N_3098);
nand U3270 (N_3270,N_3163,N_3108);
or U3271 (N_3271,N_3064,N_3196);
or U3272 (N_3272,N_3061,N_3199);
nor U3273 (N_3273,N_3197,N_3113);
nand U3274 (N_3274,N_3029,N_3067);
or U3275 (N_3275,N_3001,N_3008);
and U3276 (N_3276,N_3193,N_3076);
xor U3277 (N_3277,N_3151,N_3022);
nand U3278 (N_3278,N_3186,N_3049);
nor U3279 (N_3279,N_3019,N_3106);
nor U3280 (N_3280,N_3185,N_3079);
and U3281 (N_3281,N_3073,N_3014);
nand U3282 (N_3282,N_3104,N_3091);
nand U3283 (N_3283,N_3071,N_3121);
nand U3284 (N_3284,N_3120,N_3154);
or U3285 (N_3285,N_3167,N_3110);
nor U3286 (N_3286,N_3028,N_3082);
or U3287 (N_3287,N_3112,N_3188);
and U3288 (N_3288,N_3189,N_3040);
nand U3289 (N_3289,N_3060,N_3158);
nor U3290 (N_3290,N_3169,N_3044);
or U3291 (N_3291,N_3198,N_3063);
or U3292 (N_3292,N_3194,N_3184);
and U3293 (N_3293,N_3153,N_3123);
nand U3294 (N_3294,N_3018,N_3105);
or U3295 (N_3295,N_3134,N_3116);
or U3296 (N_3296,N_3074,N_3155);
xnor U3297 (N_3297,N_3111,N_3039);
xor U3298 (N_3298,N_3025,N_3011);
or U3299 (N_3299,N_3143,N_3139);
or U3300 (N_3300,N_3167,N_3078);
xor U3301 (N_3301,N_3187,N_3027);
and U3302 (N_3302,N_3107,N_3151);
nand U3303 (N_3303,N_3195,N_3116);
xnor U3304 (N_3304,N_3007,N_3120);
nand U3305 (N_3305,N_3000,N_3185);
xor U3306 (N_3306,N_3051,N_3178);
and U3307 (N_3307,N_3086,N_3105);
or U3308 (N_3308,N_3082,N_3083);
xor U3309 (N_3309,N_3057,N_3155);
and U3310 (N_3310,N_3144,N_3024);
and U3311 (N_3311,N_3083,N_3131);
or U3312 (N_3312,N_3140,N_3138);
nor U3313 (N_3313,N_3176,N_3120);
nand U3314 (N_3314,N_3159,N_3037);
nand U3315 (N_3315,N_3073,N_3085);
or U3316 (N_3316,N_3133,N_3064);
xor U3317 (N_3317,N_3103,N_3179);
nand U3318 (N_3318,N_3022,N_3053);
nor U3319 (N_3319,N_3120,N_3169);
xnor U3320 (N_3320,N_3155,N_3148);
and U3321 (N_3321,N_3064,N_3125);
or U3322 (N_3322,N_3020,N_3105);
and U3323 (N_3323,N_3025,N_3021);
or U3324 (N_3324,N_3027,N_3105);
nand U3325 (N_3325,N_3004,N_3153);
nor U3326 (N_3326,N_3139,N_3085);
and U3327 (N_3327,N_3002,N_3067);
xor U3328 (N_3328,N_3009,N_3180);
nor U3329 (N_3329,N_3092,N_3026);
nor U3330 (N_3330,N_3067,N_3006);
xor U3331 (N_3331,N_3136,N_3078);
and U3332 (N_3332,N_3023,N_3183);
nor U3333 (N_3333,N_3086,N_3139);
nand U3334 (N_3334,N_3186,N_3009);
nand U3335 (N_3335,N_3113,N_3130);
and U3336 (N_3336,N_3128,N_3072);
nor U3337 (N_3337,N_3071,N_3018);
and U3338 (N_3338,N_3078,N_3084);
nand U3339 (N_3339,N_3036,N_3003);
nor U3340 (N_3340,N_3180,N_3151);
nand U3341 (N_3341,N_3003,N_3012);
nand U3342 (N_3342,N_3198,N_3193);
nor U3343 (N_3343,N_3124,N_3191);
or U3344 (N_3344,N_3197,N_3130);
or U3345 (N_3345,N_3160,N_3142);
and U3346 (N_3346,N_3141,N_3098);
and U3347 (N_3347,N_3179,N_3092);
nor U3348 (N_3348,N_3085,N_3005);
nand U3349 (N_3349,N_3178,N_3074);
nand U3350 (N_3350,N_3116,N_3174);
and U3351 (N_3351,N_3015,N_3061);
and U3352 (N_3352,N_3064,N_3198);
or U3353 (N_3353,N_3093,N_3136);
and U3354 (N_3354,N_3003,N_3185);
nor U3355 (N_3355,N_3075,N_3093);
or U3356 (N_3356,N_3020,N_3021);
or U3357 (N_3357,N_3128,N_3013);
or U3358 (N_3358,N_3087,N_3025);
xor U3359 (N_3359,N_3035,N_3054);
or U3360 (N_3360,N_3154,N_3123);
nand U3361 (N_3361,N_3142,N_3109);
or U3362 (N_3362,N_3033,N_3165);
or U3363 (N_3363,N_3126,N_3084);
and U3364 (N_3364,N_3133,N_3088);
xnor U3365 (N_3365,N_3019,N_3094);
and U3366 (N_3366,N_3177,N_3192);
and U3367 (N_3367,N_3143,N_3092);
nor U3368 (N_3368,N_3089,N_3049);
and U3369 (N_3369,N_3142,N_3058);
xor U3370 (N_3370,N_3024,N_3173);
or U3371 (N_3371,N_3152,N_3081);
or U3372 (N_3372,N_3108,N_3157);
nor U3373 (N_3373,N_3064,N_3021);
nor U3374 (N_3374,N_3152,N_3147);
or U3375 (N_3375,N_3174,N_3196);
and U3376 (N_3376,N_3025,N_3036);
nor U3377 (N_3377,N_3136,N_3170);
nor U3378 (N_3378,N_3193,N_3123);
xor U3379 (N_3379,N_3014,N_3085);
or U3380 (N_3380,N_3013,N_3137);
or U3381 (N_3381,N_3063,N_3022);
and U3382 (N_3382,N_3096,N_3044);
or U3383 (N_3383,N_3199,N_3056);
and U3384 (N_3384,N_3000,N_3148);
xor U3385 (N_3385,N_3185,N_3179);
nor U3386 (N_3386,N_3036,N_3047);
nand U3387 (N_3387,N_3068,N_3191);
xor U3388 (N_3388,N_3175,N_3099);
nor U3389 (N_3389,N_3162,N_3167);
nand U3390 (N_3390,N_3051,N_3141);
and U3391 (N_3391,N_3159,N_3177);
nor U3392 (N_3392,N_3150,N_3166);
nor U3393 (N_3393,N_3044,N_3053);
and U3394 (N_3394,N_3137,N_3093);
or U3395 (N_3395,N_3023,N_3126);
or U3396 (N_3396,N_3193,N_3173);
or U3397 (N_3397,N_3016,N_3142);
or U3398 (N_3398,N_3095,N_3080);
nor U3399 (N_3399,N_3084,N_3157);
xor U3400 (N_3400,N_3200,N_3305);
and U3401 (N_3401,N_3205,N_3394);
or U3402 (N_3402,N_3201,N_3358);
and U3403 (N_3403,N_3218,N_3342);
nor U3404 (N_3404,N_3360,N_3254);
or U3405 (N_3405,N_3301,N_3211);
and U3406 (N_3406,N_3294,N_3379);
or U3407 (N_3407,N_3202,N_3264);
xnor U3408 (N_3408,N_3380,N_3232);
nand U3409 (N_3409,N_3224,N_3214);
or U3410 (N_3410,N_3398,N_3287);
xnor U3411 (N_3411,N_3251,N_3312);
nand U3412 (N_3412,N_3340,N_3243);
xor U3413 (N_3413,N_3392,N_3395);
nor U3414 (N_3414,N_3275,N_3223);
nand U3415 (N_3415,N_3249,N_3337);
nand U3416 (N_3416,N_3366,N_3383);
or U3417 (N_3417,N_3262,N_3245);
xnor U3418 (N_3418,N_3210,N_3276);
and U3419 (N_3419,N_3246,N_3391);
and U3420 (N_3420,N_3336,N_3300);
xor U3421 (N_3421,N_3384,N_3373);
nand U3422 (N_3422,N_3348,N_3216);
and U3423 (N_3423,N_3284,N_3319);
nor U3424 (N_3424,N_3356,N_3330);
nand U3425 (N_3425,N_3368,N_3256);
nor U3426 (N_3426,N_3209,N_3268);
or U3427 (N_3427,N_3274,N_3215);
and U3428 (N_3428,N_3381,N_3248);
xor U3429 (N_3429,N_3213,N_3206);
nand U3430 (N_3430,N_3230,N_3282);
and U3431 (N_3431,N_3203,N_3372);
nand U3432 (N_3432,N_3280,N_3322);
and U3433 (N_3433,N_3204,N_3387);
or U3434 (N_3434,N_3389,N_3285);
xnor U3435 (N_3435,N_3378,N_3364);
xor U3436 (N_3436,N_3354,N_3258);
and U3437 (N_3437,N_3252,N_3344);
nor U3438 (N_3438,N_3307,N_3244);
and U3439 (N_3439,N_3236,N_3396);
or U3440 (N_3440,N_3329,N_3388);
nand U3441 (N_3441,N_3212,N_3234);
or U3442 (N_3442,N_3318,N_3334);
and U3443 (N_3443,N_3314,N_3221);
xnor U3444 (N_3444,N_3365,N_3207);
and U3445 (N_3445,N_3390,N_3367);
nor U3446 (N_3446,N_3238,N_3313);
and U3447 (N_3447,N_3260,N_3267);
nand U3448 (N_3448,N_3283,N_3240);
xor U3449 (N_3449,N_3349,N_3227);
and U3450 (N_3450,N_3361,N_3304);
xor U3451 (N_3451,N_3363,N_3325);
xor U3452 (N_3452,N_3352,N_3316);
xnor U3453 (N_3453,N_3257,N_3362);
xnor U3454 (N_3454,N_3225,N_3270);
nor U3455 (N_3455,N_3253,N_3332);
xnor U3456 (N_3456,N_3228,N_3317);
nand U3457 (N_3457,N_3350,N_3311);
xnor U3458 (N_3458,N_3242,N_3231);
nor U3459 (N_3459,N_3296,N_3297);
nor U3460 (N_3460,N_3339,N_3382);
and U3461 (N_3461,N_3347,N_3278);
xnor U3462 (N_3462,N_3385,N_3235);
nor U3463 (N_3463,N_3255,N_3226);
nand U3464 (N_3464,N_3217,N_3273);
or U3465 (N_3465,N_3341,N_3265);
or U3466 (N_3466,N_3393,N_3370);
xor U3467 (N_3467,N_3298,N_3292);
and U3468 (N_3468,N_3247,N_3327);
and U3469 (N_3469,N_3371,N_3353);
or U3470 (N_3470,N_3386,N_3374);
or U3471 (N_3471,N_3323,N_3291);
nand U3472 (N_3472,N_3399,N_3293);
and U3473 (N_3473,N_3355,N_3376);
nor U3474 (N_3474,N_3328,N_3208);
xor U3475 (N_3475,N_3281,N_3220);
and U3476 (N_3476,N_3306,N_3277);
or U3477 (N_3477,N_3315,N_3266);
nor U3478 (N_3478,N_3331,N_3303);
and U3479 (N_3479,N_3343,N_3357);
or U3480 (N_3480,N_3279,N_3271);
nand U3481 (N_3481,N_3239,N_3286);
and U3482 (N_3482,N_3259,N_3222);
or U3483 (N_3483,N_3359,N_3263);
xnor U3484 (N_3484,N_3333,N_3369);
nand U3485 (N_3485,N_3345,N_3321);
xor U3486 (N_3486,N_3320,N_3290);
nand U3487 (N_3487,N_3261,N_3237);
and U3488 (N_3488,N_3397,N_3241);
nor U3489 (N_3489,N_3351,N_3302);
and U3490 (N_3490,N_3335,N_3219);
or U3491 (N_3491,N_3377,N_3299);
nand U3492 (N_3492,N_3295,N_3250);
or U3493 (N_3493,N_3324,N_3338);
xnor U3494 (N_3494,N_3233,N_3310);
nand U3495 (N_3495,N_3272,N_3308);
nand U3496 (N_3496,N_3289,N_3288);
nor U3497 (N_3497,N_3229,N_3309);
xor U3498 (N_3498,N_3326,N_3346);
and U3499 (N_3499,N_3269,N_3375);
nand U3500 (N_3500,N_3361,N_3385);
or U3501 (N_3501,N_3378,N_3363);
or U3502 (N_3502,N_3260,N_3233);
nand U3503 (N_3503,N_3217,N_3281);
and U3504 (N_3504,N_3239,N_3347);
and U3505 (N_3505,N_3344,N_3308);
nand U3506 (N_3506,N_3269,N_3384);
nor U3507 (N_3507,N_3334,N_3394);
xor U3508 (N_3508,N_3362,N_3317);
and U3509 (N_3509,N_3265,N_3347);
nor U3510 (N_3510,N_3355,N_3242);
and U3511 (N_3511,N_3276,N_3213);
or U3512 (N_3512,N_3367,N_3345);
xor U3513 (N_3513,N_3289,N_3298);
or U3514 (N_3514,N_3380,N_3306);
or U3515 (N_3515,N_3333,N_3245);
or U3516 (N_3516,N_3301,N_3346);
or U3517 (N_3517,N_3323,N_3370);
xnor U3518 (N_3518,N_3343,N_3397);
xnor U3519 (N_3519,N_3271,N_3273);
or U3520 (N_3520,N_3281,N_3202);
nor U3521 (N_3521,N_3379,N_3267);
nor U3522 (N_3522,N_3342,N_3381);
nor U3523 (N_3523,N_3221,N_3227);
nor U3524 (N_3524,N_3251,N_3328);
nand U3525 (N_3525,N_3327,N_3266);
and U3526 (N_3526,N_3353,N_3229);
xor U3527 (N_3527,N_3202,N_3379);
and U3528 (N_3528,N_3323,N_3278);
xnor U3529 (N_3529,N_3265,N_3232);
nor U3530 (N_3530,N_3342,N_3324);
and U3531 (N_3531,N_3304,N_3367);
or U3532 (N_3532,N_3306,N_3371);
and U3533 (N_3533,N_3268,N_3222);
xor U3534 (N_3534,N_3280,N_3326);
xor U3535 (N_3535,N_3241,N_3373);
nand U3536 (N_3536,N_3349,N_3280);
nand U3537 (N_3537,N_3314,N_3331);
xnor U3538 (N_3538,N_3302,N_3300);
nand U3539 (N_3539,N_3355,N_3236);
nand U3540 (N_3540,N_3365,N_3211);
xnor U3541 (N_3541,N_3325,N_3313);
xnor U3542 (N_3542,N_3354,N_3257);
xor U3543 (N_3543,N_3280,N_3361);
and U3544 (N_3544,N_3342,N_3302);
or U3545 (N_3545,N_3260,N_3258);
nand U3546 (N_3546,N_3349,N_3358);
and U3547 (N_3547,N_3260,N_3327);
xor U3548 (N_3548,N_3277,N_3385);
nor U3549 (N_3549,N_3206,N_3258);
or U3550 (N_3550,N_3343,N_3398);
or U3551 (N_3551,N_3262,N_3231);
or U3552 (N_3552,N_3227,N_3218);
xor U3553 (N_3553,N_3328,N_3321);
nand U3554 (N_3554,N_3244,N_3225);
nand U3555 (N_3555,N_3273,N_3278);
nor U3556 (N_3556,N_3300,N_3246);
nand U3557 (N_3557,N_3342,N_3397);
nor U3558 (N_3558,N_3229,N_3318);
or U3559 (N_3559,N_3368,N_3339);
nand U3560 (N_3560,N_3382,N_3303);
xnor U3561 (N_3561,N_3303,N_3260);
nor U3562 (N_3562,N_3366,N_3215);
xor U3563 (N_3563,N_3269,N_3311);
or U3564 (N_3564,N_3203,N_3264);
or U3565 (N_3565,N_3264,N_3258);
and U3566 (N_3566,N_3254,N_3274);
nand U3567 (N_3567,N_3216,N_3280);
or U3568 (N_3568,N_3237,N_3349);
nor U3569 (N_3569,N_3214,N_3234);
or U3570 (N_3570,N_3347,N_3247);
xnor U3571 (N_3571,N_3312,N_3273);
nand U3572 (N_3572,N_3348,N_3311);
nand U3573 (N_3573,N_3250,N_3360);
nand U3574 (N_3574,N_3302,N_3279);
nor U3575 (N_3575,N_3224,N_3365);
and U3576 (N_3576,N_3258,N_3313);
xor U3577 (N_3577,N_3334,N_3274);
and U3578 (N_3578,N_3207,N_3318);
nor U3579 (N_3579,N_3312,N_3264);
and U3580 (N_3580,N_3278,N_3226);
or U3581 (N_3581,N_3367,N_3298);
and U3582 (N_3582,N_3223,N_3383);
nor U3583 (N_3583,N_3348,N_3282);
and U3584 (N_3584,N_3221,N_3217);
nor U3585 (N_3585,N_3293,N_3251);
nand U3586 (N_3586,N_3291,N_3310);
nand U3587 (N_3587,N_3313,N_3394);
nor U3588 (N_3588,N_3393,N_3231);
and U3589 (N_3589,N_3236,N_3260);
nand U3590 (N_3590,N_3394,N_3342);
or U3591 (N_3591,N_3213,N_3384);
and U3592 (N_3592,N_3239,N_3288);
nor U3593 (N_3593,N_3214,N_3238);
or U3594 (N_3594,N_3211,N_3317);
nand U3595 (N_3595,N_3200,N_3218);
or U3596 (N_3596,N_3350,N_3328);
nand U3597 (N_3597,N_3369,N_3309);
or U3598 (N_3598,N_3221,N_3269);
xnor U3599 (N_3599,N_3342,N_3375);
xnor U3600 (N_3600,N_3468,N_3433);
or U3601 (N_3601,N_3464,N_3547);
nor U3602 (N_3602,N_3504,N_3535);
nor U3603 (N_3603,N_3518,N_3491);
nand U3604 (N_3604,N_3505,N_3563);
nand U3605 (N_3605,N_3465,N_3417);
nand U3606 (N_3606,N_3447,N_3531);
nor U3607 (N_3607,N_3428,N_3446);
nor U3608 (N_3608,N_3499,N_3544);
and U3609 (N_3609,N_3474,N_3415);
xor U3610 (N_3610,N_3508,N_3423);
xor U3611 (N_3611,N_3469,N_3488);
nand U3612 (N_3612,N_3419,N_3459);
or U3613 (N_3613,N_3557,N_3455);
nor U3614 (N_3614,N_3462,N_3536);
or U3615 (N_3615,N_3525,N_3421);
xor U3616 (N_3616,N_3451,N_3479);
or U3617 (N_3617,N_3414,N_3411);
nand U3618 (N_3618,N_3556,N_3425);
nor U3619 (N_3619,N_3475,N_3591);
nor U3620 (N_3620,N_3486,N_3485);
and U3621 (N_3621,N_3438,N_3461);
nor U3622 (N_3622,N_3506,N_3522);
and U3623 (N_3623,N_3532,N_3590);
nor U3624 (N_3624,N_3408,N_3534);
and U3625 (N_3625,N_3496,N_3574);
and U3626 (N_3626,N_3489,N_3598);
nand U3627 (N_3627,N_3568,N_3422);
and U3628 (N_3628,N_3510,N_3529);
nand U3629 (N_3629,N_3429,N_3467);
or U3630 (N_3630,N_3418,N_3426);
and U3631 (N_3631,N_3424,N_3542);
nor U3632 (N_3632,N_3502,N_3517);
nor U3633 (N_3633,N_3523,N_3498);
nand U3634 (N_3634,N_3443,N_3587);
nand U3635 (N_3635,N_3595,N_3541);
nand U3636 (N_3636,N_3445,N_3472);
or U3637 (N_3637,N_3543,N_3588);
nand U3638 (N_3638,N_3530,N_3483);
nand U3639 (N_3639,N_3580,N_3401);
xnor U3640 (N_3640,N_3537,N_3512);
and U3641 (N_3641,N_3520,N_3495);
nor U3642 (N_3642,N_3589,N_3549);
nand U3643 (N_3643,N_3457,N_3561);
and U3644 (N_3644,N_3404,N_3403);
nor U3645 (N_3645,N_3473,N_3487);
or U3646 (N_3646,N_3454,N_3503);
or U3647 (N_3647,N_3493,N_3481);
nand U3648 (N_3648,N_3400,N_3584);
nand U3649 (N_3649,N_3416,N_3579);
nand U3650 (N_3650,N_3482,N_3507);
nor U3651 (N_3651,N_3463,N_3578);
xor U3652 (N_3652,N_3453,N_3514);
nand U3653 (N_3653,N_3492,N_3406);
and U3654 (N_3654,N_3560,N_3427);
and U3655 (N_3655,N_3405,N_3448);
nor U3656 (N_3656,N_3494,N_3439);
and U3657 (N_3657,N_3511,N_3430);
or U3658 (N_3658,N_3476,N_3555);
or U3659 (N_3659,N_3599,N_3435);
nor U3660 (N_3660,N_3596,N_3449);
nor U3661 (N_3661,N_3594,N_3456);
xor U3662 (N_3662,N_3500,N_3582);
nor U3663 (N_3663,N_3524,N_3509);
and U3664 (N_3664,N_3466,N_3539);
nand U3665 (N_3665,N_3553,N_3413);
and U3666 (N_3666,N_3478,N_3576);
nand U3667 (N_3667,N_3527,N_3558);
nor U3668 (N_3668,N_3597,N_3420);
and U3669 (N_3669,N_3444,N_3480);
nand U3670 (N_3670,N_3432,N_3565);
nand U3671 (N_3671,N_3572,N_3501);
and U3672 (N_3672,N_3442,N_3450);
or U3673 (N_3673,N_3583,N_3460);
and U3674 (N_3674,N_3564,N_3516);
nor U3675 (N_3675,N_3410,N_3548);
and U3676 (N_3676,N_3551,N_3592);
nor U3677 (N_3677,N_3533,N_3571);
xor U3678 (N_3678,N_3559,N_3581);
nor U3679 (N_3679,N_3513,N_3437);
or U3680 (N_3680,N_3528,N_3562);
and U3681 (N_3681,N_3402,N_3471);
nand U3682 (N_3682,N_3573,N_3497);
xor U3683 (N_3683,N_3409,N_3526);
or U3684 (N_3684,N_3577,N_3585);
or U3685 (N_3685,N_3452,N_3434);
and U3686 (N_3686,N_3575,N_3593);
nor U3687 (N_3687,N_3436,N_3458);
nand U3688 (N_3688,N_3570,N_3554);
nand U3689 (N_3689,N_3552,N_3519);
nor U3690 (N_3690,N_3586,N_3470);
or U3691 (N_3691,N_3521,N_3545);
nand U3692 (N_3692,N_3407,N_3440);
xnor U3693 (N_3693,N_3569,N_3550);
or U3694 (N_3694,N_3431,N_3441);
nand U3695 (N_3695,N_3490,N_3412);
nor U3696 (N_3696,N_3538,N_3566);
nor U3697 (N_3697,N_3540,N_3515);
nor U3698 (N_3698,N_3546,N_3477);
nand U3699 (N_3699,N_3567,N_3484);
and U3700 (N_3700,N_3586,N_3425);
or U3701 (N_3701,N_3562,N_3522);
or U3702 (N_3702,N_3526,N_3517);
nor U3703 (N_3703,N_3514,N_3451);
xnor U3704 (N_3704,N_3455,N_3523);
or U3705 (N_3705,N_3499,N_3445);
nor U3706 (N_3706,N_3478,N_3512);
nand U3707 (N_3707,N_3557,N_3588);
xor U3708 (N_3708,N_3526,N_3521);
and U3709 (N_3709,N_3512,N_3595);
xor U3710 (N_3710,N_3493,N_3542);
and U3711 (N_3711,N_3487,N_3495);
xnor U3712 (N_3712,N_3553,N_3465);
xnor U3713 (N_3713,N_3496,N_3441);
nor U3714 (N_3714,N_3536,N_3599);
nor U3715 (N_3715,N_3598,N_3490);
nand U3716 (N_3716,N_3467,N_3595);
nand U3717 (N_3717,N_3581,N_3583);
nand U3718 (N_3718,N_3404,N_3503);
nand U3719 (N_3719,N_3479,N_3402);
or U3720 (N_3720,N_3444,N_3557);
nor U3721 (N_3721,N_3412,N_3447);
and U3722 (N_3722,N_3563,N_3487);
and U3723 (N_3723,N_3490,N_3406);
and U3724 (N_3724,N_3465,N_3567);
or U3725 (N_3725,N_3588,N_3534);
or U3726 (N_3726,N_3543,N_3571);
or U3727 (N_3727,N_3511,N_3550);
nor U3728 (N_3728,N_3512,N_3502);
or U3729 (N_3729,N_3548,N_3428);
or U3730 (N_3730,N_3587,N_3545);
nand U3731 (N_3731,N_3488,N_3519);
and U3732 (N_3732,N_3423,N_3506);
nor U3733 (N_3733,N_3463,N_3492);
nand U3734 (N_3734,N_3476,N_3489);
or U3735 (N_3735,N_3509,N_3437);
nor U3736 (N_3736,N_3591,N_3543);
xor U3737 (N_3737,N_3455,N_3422);
xnor U3738 (N_3738,N_3523,N_3426);
xor U3739 (N_3739,N_3478,N_3477);
and U3740 (N_3740,N_3401,N_3421);
nand U3741 (N_3741,N_3599,N_3456);
nand U3742 (N_3742,N_3481,N_3486);
and U3743 (N_3743,N_3510,N_3484);
and U3744 (N_3744,N_3547,N_3524);
nor U3745 (N_3745,N_3530,N_3566);
nand U3746 (N_3746,N_3423,N_3507);
or U3747 (N_3747,N_3462,N_3522);
and U3748 (N_3748,N_3575,N_3524);
or U3749 (N_3749,N_3565,N_3506);
nor U3750 (N_3750,N_3588,N_3559);
nand U3751 (N_3751,N_3568,N_3571);
xor U3752 (N_3752,N_3451,N_3481);
nand U3753 (N_3753,N_3466,N_3533);
xnor U3754 (N_3754,N_3573,N_3461);
or U3755 (N_3755,N_3426,N_3423);
nand U3756 (N_3756,N_3483,N_3510);
xor U3757 (N_3757,N_3415,N_3441);
or U3758 (N_3758,N_3407,N_3447);
nand U3759 (N_3759,N_3562,N_3545);
or U3760 (N_3760,N_3493,N_3567);
xnor U3761 (N_3761,N_3546,N_3442);
nor U3762 (N_3762,N_3425,N_3569);
nand U3763 (N_3763,N_3483,N_3467);
or U3764 (N_3764,N_3598,N_3436);
nor U3765 (N_3765,N_3439,N_3421);
nor U3766 (N_3766,N_3416,N_3587);
nand U3767 (N_3767,N_3583,N_3417);
xor U3768 (N_3768,N_3424,N_3518);
nor U3769 (N_3769,N_3579,N_3442);
xnor U3770 (N_3770,N_3568,N_3468);
or U3771 (N_3771,N_3512,N_3461);
nor U3772 (N_3772,N_3500,N_3518);
xnor U3773 (N_3773,N_3491,N_3587);
nor U3774 (N_3774,N_3577,N_3545);
nand U3775 (N_3775,N_3595,N_3582);
nand U3776 (N_3776,N_3445,N_3422);
and U3777 (N_3777,N_3578,N_3427);
xnor U3778 (N_3778,N_3456,N_3431);
xnor U3779 (N_3779,N_3441,N_3452);
nor U3780 (N_3780,N_3585,N_3555);
and U3781 (N_3781,N_3402,N_3409);
or U3782 (N_3782,N_3577,N_3479);
xnor U3783 (N_3783,N_3417,N_3438);
nor U3784 (N_3784,N_3436,N_3566);
nor U3785 (N_3785,N_3441,N_3449);
and U3786 (N_3786,N_3558,N_3533);
xor U3787 (N_3787,N_3402,N_3458);
xnor U3788 (N_3788,N_3589,N_3551);
and U3789 (N_3789,N_3440,N_3591);
or U3790 (N_3790,N_3595,N_3453);
xor U3791 (N_3791,N_3419,N_3503);
or U3792 (N_3792,N_3510,N_3573);
nor U3793 (N_3793,N_3453,N_3455);
nor U3794 (N_3794,N_3499,N_3401);
or U3795 (N_3795,N_3476,N_3446);
xor U3796 (N_3796,N_3543,N_3436);
and U3797 (N_3797,N_3575,N_3448);
xnor U3798 (N_3798,N_3545,N_3544);
and U3799 (N_3799,N_3580,N_3512);
xnor U3800 (N_3800,N_3667,N_3753);
xor U3801 (N_3801,N_3682,N_3605);
nand U3802 (N_3802,N_3771,N_3660);
nor U3803 (N_3803,N_3649,N_3726);
nor U3804 (N_3804,N_3714,N_3701);
nor U3805 (N_3805,N_3683,N_3748);
nor U3806 (N_3806,N_3708,N_3722);
xnor U3807 (N_3807,N_3624,N_3739);
nor U3808 (N_3808,N_3681,N_3703);
nor U3809 (N_3809,N_3740,N_3719);
and U3810 (N_3810,N_3652,N_3710);
or U3811 (N_3811,N_3784,N_3777);
nand U3812 (N_3812,N_3775,N_3735);
nand U3813 (N_3813,N_3713,N_3687);
xnor U3814 (N_3814,N_3761,N_3688);
nor U3815 (N_3815,N_3659,N_3680);
and U3816 (N_3816,N_3643,N_3693);
or U3817 (N_3817,N_3615,N_3795);
and U3818 (N_3818,N_3706,N_3621);
nand U3819 (N_3819,N_3647,N_3782);
nor U3820 (N_3820,N_3675,N_3712);
nor U3821 (N_3821,N_3611,N_3689);
and U3822 (N_3822,N_3750,N_3655);
nor U3823 (N_3823,N_3796,N_3639);
and U3824 (N_3824,N_3634,N_3670);
or U3825 (N_3825,N_3696,N_3603);
and U3826 (N_3826,N_3769,N_3671);
nor U3827 (N_3827,N_3785,N_3786);
nor U3828 (N_3828,N_3653,N_3763);
nand U3829 (N_3829,N_3674,N_3736);
xor U3830 (N_3830,N_3664,N_3705);
and U3831 (N_3831,N_3610,N_3730);
xnor U3832 (N_3832,N_3749,N_3656);
nand U3833 (N_3833,N_3773,N_3791);
nand U3834 (N_3834,N_3768,N_3690);
xor U3835 (N_3835,N_3640,N_3751);
nand U3836 (N_3836,N_3737,N_3756);
and U3837 (N_3837,N_3702,N_3633);
nor U3838 (N_3838,N_3704,N_3684);
nand U3839 (N_3839,N_3745,N_3755);
or U3840 (N_3840,N_3698,N_3743);
nor U3841 (N_3841,N_3758,N_3757);
nand U3842 (N_3842,N_3691,N_3759);
and U3843 (N_3843,N_3678,N_3685);
xnor U3844 (N_3844,N_3789,N_3642);
xor U3845 (N_3845,N_3723,N_3629);
xor U3846 (N_3846,N_3613,N_3648);
xor U3847 (N_3847,N_3651,N_3631);
and U3848 (N_3848,N_3774,N_3793);
and U3849 (N_3849,N_3742,N_3665);
nor U3850 (N_3850,N_3733,N_3673);
or U3851 (N_3851,N_3646,N_3746);
and U3852 (N_3852,N_3731,N_3715);
xnor U3853 (N_3853,N_3609,N_3741);
nor U3854 (N_3854,N_3754,N_3669);
nand U3855 (N_3855,N_3744,N_3732);
nand U3856 (N_3856,N_3620,N_3707);
and U3857 (N_3857,N_3636,N_3630);
xnor U3858 (N_3858,N_3632,N_3614);
and U3859 (N_3859,N_3650,N_3627);
and U3860 (N_3860,N_3622,N_3792);
nor U3861 (N_3861,N_3637,N_3764);
nor U3862 (N_3862,N_3720,N_3602);
and U3863 (N_3863,N_3607,N_3677);
or U3864 (N_3864,N_3770,N_3716);
nand U3865 (N_3865,N_3697,N_3781);
nor U3866 (N_3866,N_3663,N_3676);
nand U3867 (N_3867,N_3625,N_3619);
and U3868 (N_3868,N_3600,N_3725);
or U3869 (N_3869,N_3699,N_3641);
nand U3870 (N_3870,N_3721,N_3612);
xor U3871 (N_3871,N_3779,N_3700);
nand U3872 (N_3872,N_3794,N_3658);
xor U3873 (N_3873,N_3606,N_3662);
nor U3874 (N_3874,N_3727,N_3601);
xnor U3875 (N_3875,N_3760,N_3790);
xnor U3876 (N_3876,N_3762,N_3724);
or U3877 (N_3877,N_3772,N_3797);
nor U3878 (N_3878,N_3766,N_3668);
nor U3879 (N_3879,N_3711,N_3752);
xnor U3880 (N_3880,N_3626,N_3628);
nand U3881 (N_3881,N_3788,N_3776);
or U3882 (N_3882,N_3717,N_3686);
nand U3883 (N_3883,N_3635,N_3780);
or U3884 (N_3884,N_3787,N_3617);
nor U3885 (N_3885,N_3666,N_3604);
xor U3886 (N_3886,N_3644,N_3661);
or U3887 (N_3887,N_3694,N_3734);
xnor U3888 (N_3888,N_3709,N_3654);
or U3889 (N_3889,N_3672,N_3623);
and U3890 (N_3890,N_3608,N_3778);
nor U3891 (N_3891,N_3738,N_3747);
or U3892 (N_3892,N_3657,N_3638);
and U3893 (N_3893,N_3692,N_3645);
xor U3894 (N_3894,N_3729,N_3618);
nor U3895 (N_3895,N_3765,N_3616);
nand U3896 (N_3896,N_3783,N_3767);
or U3897 (N_3897,N_3695,N_3718);
and U3898 (N_3898,N_3798,N_3679);
xor U3899 (N_3899,N_3799,N_3728);
xnor U3900 (N_3900,N_3614,N_3687);
xor U3901 (N_3901,N_3625,N_3678);
nor U3902 (N_3902,N_3789,N_3611);
and U3903 (N_3903,N_3680,N_3676);
xnor U3904 (N_3904,N_3763,N_3600);
and U3905 (N_3905,N_3701,N_3798);
nor U3906 (N_3906,N_3634,N_3672);
xnor U3907 (N_3907,N_3620,N_3792);
or U3908 (N_3908,N_3742,N_3686);
nand U3909 (N_3909,N_3732,N_3724);
nand U3910 (N_3910,N_3755,N_3748);
nand U3911 (N_3911,N_3713,N_3714);
and U3912 (N_3912,N_3755,N_3656);
nand U3913 (N_3913,N_3695,N_3611);
and U3914 (N_3914,N_3675,N_3605);
nor U3915 (N_3915,N_3650,N_3641);
xor U3916 (N_3916,N_3705,N_3771);
or U3917 (N_3917,N_3703,N_3759);
nand U3918 (N_3918,N_3796,N_3769);
xor U3919 (N_3919,N_3604,N_3799);
xnor U3920 (N_3920,N_3612,N_3605);
nor U3921 (N_3921,N_3662,N_3723);
or U3922 (N_3922,N_3643,N_3629);
and U3923 (N_3923,N_3709,N_3740);
nor U3924 (N_3924,N_3646,N_3787);
xor U3925 (N_3925,N_3786,N_3684);
or U3926 (N_3926,N_3727,N_3672);
nor U3927 (N_3927,N_3628,N_3676);
or U3928 (N_3928,N_3654,N_3795);
and U3929 (N_3929,N_3608,N_3764);
nor U3930 (N_3930,N_3752,N_3764);
xor U3931 (N_3931,N_3720,N_3744);
nand U3932 (N_3932,N_3798,N_3614);
nand U3933 (N_3933,N_3747,N_3653);
or U3934 (N_3934,N_3793,N_3621);
nand U3935 (N_3935,N_3631,N_3713);
xnor U3936 (N_3936,N_3685,N_3650);
and U3937 (N_3937,N_3744,N_3678);
or U3938 (N_3938,N_3688,N_3737);
nand U3939 (N_3939,N_3752,N_3616);
nor U3940 (N_3940,N_3751,N_3646);
nand U3941 (N_3941,N_3644,N_3781);
xor U3942 (N_3942,N_3771,N_3619);
or U3943 (N_3943,N_3628,N_3648);
nor U3944 (N_3944,N_3760,N_3650);
and U3945 (N_3945,N_3623,N_3732);
xor U3946 (N_3946,N_3745,N_3680);
or U3947 (N_3947,N_3618,N_3645);
nand U3948 (N_3948,N_3745,N_3763);
xnor U3949 (N_3949,N_3762,N_3798);
nor U3950 (N_3950,N_3754,N_3667);
nor U3951 (N_3951,N_3661,N_3601);
nand U3952 (N_3952,N_3735,N_3649);
and U3953 (N_3953,N_3782,N_3708);
nor U3954 (N_3954,N_3719,N_3730);
nand U3955 (N_3955,N_3658,N_3732);
or U3956 (N_3956,N_3621,N_3636);
and U3957 (N_3957,N_3760,N_3789);
or U3958 (N_3958,N_3699,N_3766);
nand U3959 (N_3959,N_3759,N_3655);
and U3960 (N_3960,N_3603,N_3604);
nor U3961 (N_3961,N_3632,N_3664);
or U3962 (N_3962,N_3761,N_3792);
or U3963 (N_3963,N_3723,N_3708);
xnor U3964 (N_3964,N_3650,N_3649);
and U3965 (N_3965,N_3745,N_3770);
nor U3966 (N_3966,N_3718,N_3771);
xnor U3967 (N_3967,N_3737,N_3720);
or U3968 (N_3968,N_3651,N_3725);
or U3969 (N_3969,N_3652,N_3603);
and U3970 (N_3970,N_3725,N_3787);
nor U3971 (N_3971,N_3782,N_3729);
or U3972 (N_3972,N_3683,N_3764);
or U3973 (N_3973,N_3782,N_3654);
nand U3974 (N_3974,N_3627,N_3628);
nor U3975 (N_3975,N_3667,N_3771);
or U3976 (N_3976,N_3785,N_3670);
nand U3977 (N_3977,N_3718,N_3773);
nand U3978 (N_3978,N_3681,N_3619);
nor U3979 (N_3979,N_3751,N_3652);
or U3980 (N_3980,N_3617,N_3688);
xnor U3981 (N_3981,N_3615,N_3704);
or U3982 (N_3982,N_3739,N_3688);
nor U3983 (N_3983,N_3751,N_3644);
nand U3984 (N_3984,N_3644,N_3663);
xnor U3985 (N_3985,N_3730,N_3688);
or U3986 (N_3986,N_3676,N_3693);
xnor U3987 (N_3987,N_3747,N_3610);
nand U3988 (N_3988,N_3746,N_3652);
xor U3989 (N_3989,N_3606,N_3687);
nand U3990 (N_3990,N_3615,N_3683);
and U3991 (N_3991,N_3606,N_3774);
nand U3992 (N_3992,N_3635,N_3742);
xor U3993 (N_3993,N_3703,N_3669);
nor U3994 (N_3994,N_3712,N_3661);
nand U3995 (N_3995,N_3779,N_3703);
and U3996 (N_3996,N_3639,N_3750);
xor U3997 (N_3997,N_3735,N_3777);
or U3998 (N_3998,N_3638,N_3619);
nand U3999 (N_3999,N_3682,N_3668);
nor U4000 (N_4000,N_3977,N_3855);
xor U4001 (N_4001,N_3821,N_3847);
nor U4002 (N_4002,N_3919,N_3917);
and U4003 (N_4003,N_3932,N_3955);
nor U4004 (N_4004,N_3882,N_3818);
or U4005 (N_4005,N_3935,N_3870);
or U4006 (N_4006,N_3999,N_3952);
or U4007 (N_4007,N_3968,N_3939);
or U4008 (N_4008,N_3898,N_3918);
nand U4009 (N_4009,N_3865,N_3947);
nor U4010 (N_4010,N_3989,N_3943);
or U4011 (N_4011,N_3931,N_3853);
and U4012 (N_4012,N_3892,N_3885);
xnor U4013 (N_4013,N_3881,N_3899);
xor U4014 (N_4014,N_3913,N_3831);
nand U4015 (N_4015,N_3975,N_3927);
nor U4016 (N_4016,N_3872,N_3914);
nand U4017 (N_4017,N_3996,N_3871);
and U4018 (N_4018,N_3967,N_3969);
or U4019 (N_4019,N_3922,N_3905);
xor U4020 (N_4020,N_3906,N_3866);
xor U4021 (N_4021,N_3985,N_3805);
nor U4022 (N_4022,N_3976,N_3860);
nor U4023 (N_4023,N_3819,N_3948);
or U4024 (N_4024,N_3813,N_3994);
nand U4025 (N_4025,N_3848,N_3876);
nor U4026 (N_4026,N_3957,N_3891);
xor U4027 (N_4027,N_3960,N_3873);
and U4028 (N_4028,N_3824,N_3949);
nand U4029 (N_4029,N_3861,N_3953);
and U4030 (N_4030,N_3904,N_3907);
nand U4031 (N_4031,N_3897,N_3941);
and U4032 (N_4032,N_3950,N_3979);
nor U4033 (N_4033,N_3852,N_3808);
xnor U4034 (N_4034,N_3962,N_3921);
and U4035 (N_4035,N_3961,N_3856);
nor U4036 (N_4036,N_3886,N_3820);
xor U4037 (N_4037,N_3851,N_3844);
or U4038 (N_4038,N_3846,N_3997);
or U4039 (N_4039,N_3837,N_3988);
nand U4040 (N_4040,N_3990,N_3814);
nand U4041 (N_4041,N_3938,N_3909);
or U4042 (N_4042,N_3836,N_3830);
or U4043 (N_4043,N_3812,N_3958);
nand U4044 (N_4044,N_3835,N_3911);
nand U4045 (N_4045,N_3964,N_3959);
xor U4046 (N_4046,N_3845,N_3995);
nor U4047 (N_4047,N_3804,N_3936);
nand U4048 (N_4048,N_3928,N_3840);
or U4049 (N_4049,N_3912,N_3889);
and U4050 (N_4050,N_3972,N_3884);
or U4051 (N_4051,N_3890,N_3838);
nand U4052 (N_4052,N_3803,N_3992);
nand U4053 (N_4053,N_3822,N_3887);
nor U4054 (N_4054,N_3900,N_3862);
nor U4055 (N_4055,N_3933,N_3903);
nor U4056 (N_4056,N_3893,N_3987);
nand U4057 (N_4057,N_3827,N_3825);
nand U4058 (N_4058,N_3924,N_3880);
or U4059 (N_4059,N_3809,N_3920);
or U4060 (N_4060,N_3815,N_3857);
xnor U4061 (N_4061,N_3910,N_3956);
nor U4062 (N_4062,N_3894,N_3883);
and U4063 (N_4063,N_3951,N_3946);
xnor U4064 (N_4064,N_3858,N_3937);
nand U4065 (N_4065,N_3929,N_3841);
and U4066 (N_4066,N_3930,N_3954);
and U4067 (N_4067,N_3925,N_3877);
and U4068 (N_4068,N_3971,N_3826);
nor U4069 (N_4069,N_3980,N_3878);
nand U4070 (N_4070,N_3801,N_3916);
or U4071 (N_4071,N_3864,N_3902);
nor U4072 (N_4072,N_3966,N_3807);
or U4073 (N_4073,N_3998,N_3895);
nor U4074 (N_4074,N_3986,N_3973);
or U4075 (N_4075,N_3832,N_3970);
and U4076 (N_4076,N_3854,N_3923);
or U4077 (N_4077,N_3879,N_3810);
xnor U4078 (N_4078,N_3817,N_3940);
and U4079 (N_4079,N_3843,N_3974);
nor U4080 (N_4080,N_3828,N_3816);
xor U4081 (N_4081,N_3850,N_3875);
or U4082 (N_4082,N_3867,N_3863);
nand U4083 (N_4083,N_3896,N_3978);
nor U4084 (N_4084,N_3983,N_3839);
nor U4085 (N_4085,N_3944,N_3926);
xor U4086 (N_4086,N_3842,N_3806);
nand U4087 (N_4087,N_3945,N_3874);
nor U4088 (N_4088,N_3982,N_3800);
or U4089 (N_4089,N_3888,N_3823);
nand U4090 (N_4090,N_3834,N_3942);
xnor U4091 (N_4091,N_3869,N_3915);
xor U4092 (N_4092,N_3802,N_3963);
or U4093 (N_4093,N_3829,N_3908);
nand U4094 (N_4094,N_3984,N_3991);
xnor U4095 (N_4095,N_3849,N_3934);
nand U4096 (N_4096,N_3833,N_3868);
nor U4097 (N_4097,N_3981,N_3965);
nand U4098 (N_4098,N_3859,N_3993);
and U4099 (N_4099,N_3811,N_3901);
nand U4100 (N_4100,N_3843,N_3932);
nor U4101 (N_4101,N_3888,N_3856);
and U4102 (N_4102,N_3856,N_3863);
nand U4103 (N_4103,N_3990,N_3860);
and U4104 (N_4104,N_3838,N_3843);
or U4105 (N_4105,N_3890,N_3986);
xnor U4106 (N_4106,N_3870,N_3846);
nor U4107 (N_4107,N_3925,N_3931);
and U4108 (N_4108,N_3944,N_3955);
and U4109 (N_4109,N_3949,N_3839);
and U4110 (N_4110,N_3998,N_3831);
nand U4111 (N_4111,N_3971,N_3890);
nor U4112 (N_4112,N_3862,N_3898);
and U4113 (N_4113,N_3950,N_3982);
xnor U4114 (N_4114,N_3958,N_3893);
or U4115 (N_4115,N_3984,N_3850);
or U4116 (N_4116,N_3827,N_3901);
nand U4117 (N_4117,N_3808,N_3886);
xor U4118 (N_4118,N_3987,N_3957);
nand U4119 (N_4119,N_3930,N_3882);
and U4120 (N_4120,N_3960,N_3860);
and U4121 (N_4121,N_3879,N_3906);
nor U4122 (N_4122,N_3932,N_3824);
or U4123 (N_4123,N_3932,N_3921);
or U4124 (N_4124,N_3956,N_3953);
and U4125 (N_4125,N_3933,N_3859);
nor U4126 (N_4126,N_3827,N_3938);
nand U4127 (N_4127,N_3869,N_3847);
and U4128 (N_4128,N_3868,N_3969);
or U4129 (N_4129,N_3843,N_3984);
or U4130 (N_4130,N_3813,N_3895);
nor U4131 (N_4131,N_3808,N_3912);
nor U4132 (N_4132,N_3981,N_3898);
and U4133 (N_4133,N_3819,N_3829);
nor U4134 (N_4134,N_3940,N_3831);
nor U4135 (N_4135,N_3929,N_3991);
nor U4136 (N_4136,N_3918,N_3830);
nand U4137 (N_4137,N_3967,N_3986);
and U4138 (N_4138,N_3937,N_3919);
nor U4139 (N_4139,N_3916,N_3980);
nor U4140 (N_4140,N_3927,N_3939);
nor U4141 (N_4141,N_3968,N_3970);
nand U4142 (N_4142,N_3879,N_3953);
nand U4143 (N_4143,N_3822,N_3884);
and U4144 (N_4144,N_3876,N_3967);
xor U4145 (N_4145,N_3823,N_3863);
nand U4146 (N_4146,N_3881,N_3901);
xnor U4147 (N_4147,N_3992,N_3813);
nand U4148 (N_4148,N_3965,N_3980);
and U4149 (N_4149,N_3855,N_3840);
nand U4150 (N_4150,N_3817,N_3904);
xnor U4151 (N_4151,N_3835,N_3945);
and U4152 (N_4152,N_3907,N_3917);
nand U4153 (N_4153,N_3974,N_3813);
nor U4154 (N_4154,N_3954,N_3848);
nand U4155 (N_4155,N_3917,N_3890);
or U4156 (N_4156,N_3844,N_3805);
and U4157 (N_4157,N_3864,N_3863);
or U4158 (N_4158,N_3942,N_3935);
nand U4159 (N_4159,N_3893,N_3812);
nor U4160 (N_4160,N_3887,N_3943);
and U4161 (N_4161,N_3885,N_3911);
xnor U4162 (N_4162,N_3852,N_3933);
or U4163 (N_4163,N_3996,N_3907);
nand U4164 (N_4164,N_3975,N_3834);
xnor U4165 (N_4165,N_3980,N_3877);
nor U4166 (N_4166,N_3970,N_3821);
or U4167 (N_4167,N_3900,N_3999);
xnor U4168 (N_4168,N_3899,N_3898);
xor U4169 (N_4169,N_3851,N_3873);
xor U4170 (N_4170,N_3941,N_3853);
and U4171 (N_4171,N_3843,N_3989);
nand U4172 (N_4172,N_3955,N_3827);
nor U4173 (N_4173,N_3991,N_3922);
and U4174 (N_4174,N_3998,N_3897);
nor U4175 (N_4175,N_3832,N_3839);
nand U4176 (N_4176,N_3906,N_3986);
and U4177 (N_4177,N_3821,N_3956);
or U4178 (N_4178,N_3921,N_3938);
nand U4179 (N_4179,N_3830,N_3928);
nor U4180 (N_4180,N_3937,N_3970);
xnor U4181 (N_4181,N_3944,N_3843);
nand U4182 (N_4182,N_3966,N_3927);
nand U4183 (N_4183,N_3885,N_3877);
and U4184 (N_4184,N_3874,N_3835);
and U4185 (N_4185,N_3983,N_3940);
xor U4186 (N_4186,N_3831,N_3876);
xor U4187 (N_4187,N_3940,N_3908);
nor U4188 (N_4188,N_3897,N_3840);
nand U4189 (N_4189,N_3854,N_3850);
nor U4190 (N_4190,N_3904,N_3964);
nand U4191 (N_4191,N_3829,N_3926);
nand U4192 (N_4192,N_3864,N_3841);
nor U4193 (N_4193,N_3922,N_3863);
xnor U4194 (N_4194,N_3918,N_3955);
nand U4195 (N_4195,N_3921,N_3945);
nor U4196 (N_4196,N_3960,N_3986);
and U4197 (N_4197,N_3895,N_3908);
and U4198 (N_4198,N_3866,N_3991);
or U4199 (N_4199,N_3826,N_3931);
and U4200 (N_4200,N_4063,N_4163);
xnor U4201 (N_4201,N_4155,N_4026);
and U4202 (N_4202,N_4179,N_4191);
or U4203 (N_4203,N_4118,N_4029);
nand U4204 (N_4204,N_4126,N_4106);
nor U4205 (N_4205,N_4059,N_4197);
xor U4206 (N_4206,N_4123,N_4154);
nor U4207 (N_4207,N_4164,N_4115);
and U4208 (N_4208,N_4032,N_4168);
nand U4209 (N_4209,N_4028,N_4084);
and U4210 (N_4210,N_4109,N_4045);
and U4211 (N_4211,N_4050,N_4167);
nor U4212 (N_4212,N_4113,N_4087);
xor U4213 (N_4213,N_4127,N_4170);
and U4214 (N_4214,N_4122,N_4002);
nor U4215 (N_4215,N_4158,N_4035);
and U4216 (N_4216,N_4007,N_4120);
and U4217 (N_4217,N_4053,N_4047);
nand U4218 (N_4218,N_4147,N_4131);
nor U4219 (N_4219,N_4042,N_4077);
and U4220 (N_4220,N_4114,N_4015);
nand U4221 (N_4221,N_4186,N_4088);
xnor U4222 (N_4222,N_4130,N_4143);
xor U4223 (N_4223,N_4112,N_4004);
nand U4224 (N_4224,N_4055,N_4136);
or U4225 (N_4225,N_4001,N_4038);
nor U4226 (N_4226,N_4018,N_4082);
xnor U4227 (N_4227,N_4171,N_4150);
or U4228 (N_4228,N_4085,N_4091);
nand U4229 (N_4229,N_4036,N_4068);
nand U4230 (N_4230,N_4030,N_4116);
nor U4231 (N_4231,N_4098,N_4173);
or U4232 (N_4232,N_4041,N_4064);
nand U4233 (N_4233,N_4110,N_4194);
and U4234 (N_4234,N_4095,N_4067);
and U4235 (N_4235,N_4017,N_4121);
xnor U4236 (N_4236,N_4025,N_4149);
nand U4237 (N_4237,N_4195,N_4180);
nor U4238 (N_4238,N_4153,N_4099);
nor U4239 (N_4239,N_4052,N_4156);
nor U4240 (N_4240,N_4071,N_4006);
xnor U4241 (N_4241,N_4145,N_4048);
nor U4242 (N_4242,N_4097,N_4016);
nor U4243 (N_4243,N_4184,N_4056);
and U4244 (N_4244,N_4160,N_4135);
and U4245 (N_4245,N_4005,N_4040);
or U4246 (N_4246,N_4037,N_4092);
xnor U4247 (N_4247,N_4176,N_4117);
xor U4248 (N_4248,N_4061,N_4076);
and U4249 (N_4249,N_4043,N_4196);
nand U4250 (N_4250,N_4054,N_4020);
or U4251 (N_4251,N_4192,N_4079);
nand U4252 (N_4252,N_4003,N_4125);
nand U4253 (N_4253,N_4011,N_4057);
xnor U4254 (N_4254,N_4174,N_4014);
and U4255 (N_4255,N_4102,N_4103);
nand U4256 (N_4256,N_4137,N_4146);
nor U4257 (N_4257,N_4090,N_4175);
xor U4258 (N_4258,N_4101,N_4024);
nor U4259 (N_4259,N_4012,N_4138);
and U4260 (N_4260,N_4044,N_4078);
xor U4261 (N_4261,N_4039,N_4083);
and U4262 (N_4262,N_4144,N_4013);
or U4263 (N_4263,N_4129,N_4198);
nand U4264 (N_4264,N_4193,N_4065);
xnor U4265 (N_4265,N_4075,N_4148);
and U4266 (N_4266,N_4069,N_4060);
and U4267 (N_4267,N_4027,N_4031);
or U4268 (N_4268,N_4051,N_4151);
and U4269 (N_4269,N_4072,N_4188);
or U4270 (N_4270,N_4134,N_4178);
xnor U4271 (N_4271,N_4166,N_4073);
xor U4272 (N_4272,N_4157,N_4133);
nor U4273 (N_4273,N_4119,N_4187);
nor U4274 (N_4274,N_4066,N_4034);
nand U4275 (N_4275,N_4089,N_4107);
or U4276 (N_4276,N_4033,N_4189);
nor U4277 (N_4277,N_4141,N_4019);
nand U4278 (N_4278,N_4165,N_4049);
nor U4279 (N_4279,N_4086,N_4021);
nor U4280 (N_4280,N_4111,N_4142);
or U4281 (N_4281,N_4093,N_4161);
or U4282 (N_4282,N_4022,N_4162);
xnor U4283 (N_4283,N_4183,N_4074);
and U4284 (N_4284,N_4182,N_4159);
or U4285 (N_4285,N_4094,N_4190);
xnor U4286 (N_4286,N_4100,N_4199);
nand U4287 (N_4287,N_4062,N_4140);
nor U4288 (N_4288,N_4081,N_4181);
or U4289 (N_4289,N_4124,N_4105);
nand U4290 (N_4290,N_4046,N_4023);
or U4291 (N_4291,N_4108,N_4008);
xnor U4292 (N_4292,N_4096,N_4128);
nand U4293 (N_4293,N_4080,N_4169);
xnor U4294 (N_4294,N_4139,N_4152);
and U4295 (N_4295,N_4058,N_4177);
xnor U4296 (N_4296,N_4185,N_4172);
nand U4297 (N_4297,N_4010,N_4070);
nor U4298 (N_4298,N_4104,N_4000);
xor U4299 (N_4299,N_4132,N_4009);
nor U4300 (N_4300,N_4132,N_4062);
xor U4301 (N_4301,N_4088,N_4080);
and U4302 (N_4302,N_4026,N_4195);
xnor U4303 (N_4303,N_4186,N_4174);
or U4304 (N_4304,N_4046,N_4122);
nand U4305 (N_4305,N_4199,N_4073);
nor U4306 (N_4306,N_4106,N_4066);
nand U4307 (N_4307,N_4038,N_4037);
xor U4308 (N_4308,N_4176,N_4118);
nand U4309 (N_4309,N_4084,N_4185);
nor U4310 (N_4310,N_4177,N_4123);
xor U4311 (N_4311,N_4104,N_4121);
and U4312 (N_4312,N_4022,N_4114);
and U4313 (N_4313,N_4101,N_4076);
or U4314 (N_4314,N_4088,N_4178);
nor U4315 (N_4315,N_4199,N_4125);
nand U4316 (N_4316,N_4004,N_4138);
or U4317 (N_4317,N_4198,N_4004);
nand U4318 (N_4318,N_4196,N_4063);
nor U4319 (N_4319,N_4148,N_4087);
and U4320 (N_4320,N_4150,N_4024);
or U4321 (N_4321,N_4139,N_4040);
nor U4322 (N_4322,N_4064,N_4147);
nor U4323 (N_4323,N_4066,N_4078);
xnor U4324 (N_4324,N_4042,N_4120);
xor U4325 (N_4325,N_4056,N_4097);
nor U4326 (N_4326,N_4050,N_4072);
nor U4327 (N_4327,N_4093,N_4114);
xor U4328 (N_4328,N_4127,N_4189);
nor U4329 (N_4329,N_4025,N_4117);
nand U4330 (N_4330,N_4040,N_4076);
and U4331 (N_4331,N_4032,N_4053);
and U4332 (N_4332,N_4073,N_4009);
nor U4333 (N_4333,N_4111,N_4141);
xor U4334 (N_4334,N_4195,N_4077);
nor U4335 (N_4335,N_4133,N_4093);
and U4336 (N_4336,N_4047,N_4042);
xnor U4337 (N_4337,N_4114,N_4179);
nor U4338 (N_4338,N_4024,N_4165);
nand U4339 (N_4339,N_4149,N_4158);
nand U4340 (N_4340,N_4165,N_4061);
or U4341 (N_4341,N_4104,N_4183);
nand U4342 (N_4342,N_4021,N_4059);
xor U4343 (N_4343,N_4118,N_4124);
nand U4344 (N_4344,N_4105,N_4174);
nand U4345 (N_4345,N_4106,N_4162);
or U4346 (N_4346,N_4095,N_4085);
nor U4347 (N_4347,N_4008,N_4189);
nand U4348 (N_4348,N_4120,N_4034);
nor U4349 (N_4349,N_4048,N_4173);
or U4350 (N_4350,N_4031,N_4028);
and U4351 (N_4351,N_4072,N_4134);
nand U4352 (N_4352,N_4166,N_4117);
xnor U4353 (N_4353,N_4169,N_4121);
or U4354 (N_4354,N_4030,N_4067);
and U4355 (N_4355,N_4177,N_4171);
nand U4356 (N_4356,N_4196,N_4122);
or U4357 (N_4357,N_4184,N_4011);
nand U4358 (N_4358,N_4184,N_4159);
nand U4359 (N_4359,N_4150,N_4094);
and U4360 (N_4360,N_4124,N_4087);
and U4361 (N_4361,N_4093,N_4113);
nor U4362 (N_4362,N_4019,N_4046);
xor U4363 (N_4363,N_4083,N_4137);
nor U4364 (N_4364,N_4118,N_4017);
nor U4365 (N_4365,N_4064,N_4016);
nor U4366 (N_4366,N_4085,N_4169);
nand U4367 (N_4367,N_4003,N_4132);
nand U4368 (N_4368,N_4058,N_4025);
xnor U4369 (N_4369,N_4183,N_4169);
nand U4370 (N_4370,N_4166,N_4099);
and U4371 (N_4371,N_4101,N_4000);
xor U4372 (N_4372,N_4110,N_4085);
xor U4373 (N_4373,N_4167,N_4035);
or U4374 (N_4374,N_4066,N_4116);
nand U4375 (N_4375,N_4134,N_4121);
and U4376 (N_4376,N_4153,N_4180);
nor U4377 (N_4377,N_4160,N_4063);
nand U4378 (N_4378,N_4013,N_4150);
and U4379 (N_4379,N_4072,N_4026);
nor U4380 (N_4380,N_4040,N_4011);
and U4381 (N_4381,N_4028,N_4179);
or U4382 (N_4382,N_4026,N_4145);
xnor U4383 (N_4383,N_4158,N_4155);
or U4384 (N_4384,N_4184,N_4179);
nor U4385 (N_4385,N_4021,N_4157);
xnor U4386 (N_4386,N_4094,N_4002);
xor U4387 (N_4387,N_4196,N_4125);
xnor U4388 (N_4388,N_4189,N_4060);
or U4389 (N_4389,N_4123,N_4116);
nand U4390 (N_4390,N_4161,N_4086);
nand U4391 (N_4391,N_4142,N_4141);
xnor U4392 (N_4392,N_4144,N_4050);
xnor U4393 (N_4393,N_4100,N_4087);
or U4394 (N_4394,N_4131,N_4070);
and U4395 (N_4395,N_4163,N_4180);
and U4396 (N_4396,N_4170,N_4082);
xor U4397 (N_4397,N_4160,N_4007);
xor U4398 (N_4398,N_4037,N_4187);
xnor U4399 (N_4399,N_4049,N_4010);
and U4400 (N_4400,N_4300,N_4257);
nor U4401 (N_4401,N_4293,N_4276);
or U4402 (N_4402,N_4275,N_4322);
or U4403 (N_4403,N_4218,N_4347);
and U4404 (N_4404,N_4312,N_4336);
nand U4405 (N_4405,N_4205,N_4213);
and U4406 (N_4406,N_4390,N_4295);
xor U4407 (N_4407,N_4305,N_4221);
nor U4408 (N_4408,N_4376,N_4314);
or U4409 (N_4409,N_4219,N_4252);
nand U4410 (N_4410,N_4385,N_4208);
and U4411 (N_4411,N_4259,N_4272);
or U4412 (N_4412,N_4309,N_4350);
and U4413 (N_4413,N_4352,N_4268);
and U4414 (N_4414,N_4212,N_4225);
and U4415 (N_4415,N_4393,N_4311);
and U4416 (N_4416,N_4229,N_4345);
or U4417 (N_4417,N_4273,N_4254);
xor U4418 (N_4418,N_4342,N_4294);
nand U4419 (N_4419,N_4262,N_4230);
nor U4420 (N_4420,N_4223,N_4333);
nand U4421 (N_4421,N_4299,N_4348);
nor U4422 (N_4422,N_4356,N_4337);
and U4423 (N_4423,N_4249,N_4354);
nor U4424 (N_4424,N_4396,N_4383);
xnor U4425 (N_4425,N_4291,N_4387);
and U4426 (N_4426,N_4282,N_4242);
xnor U4427 (N_4427,N_4371,N_4368);
nand U4428 (N_4428,N_4395,N_4277);
xor U4429 (N_4429,N_4329,N_4255);
or U4430 (N_4430,N_4256,N_4214);
and U4431 (N_4431,N_4251,N_4279);
nor U4432 (N_4432,N_4362,N_4215);
and U4433 (N_4433,N_4226,N_4364);
or U4434 (N_4434,N_4304,N_4344);
nor U4435 (N_4435,N_4391,N_4326);
or U4436 (N_4436,N_4301,N_4360);
nand U4437 (N_4437,N_4324,N_4378);
nor U4438 (N_4438,N_4211,N_4222);
or U4439 (N_4439,N_4216,N_4308);
or U4440 (N_4440,N_4233,N_4339);
or U4441 (N_4441,N_4201,N_4346);
nor U4442 (N_4442,N_4238,N_4203);
nand U4443 (N_4443,N_4239,N_4264);
nand U4444 (N_4444,N_4260,N_4319);
and U4445 (N_4445,N_4320,N_4292);
xor U4446 (N_4446,N_4361,N_4297);
nor U4447 (N_4447,N_4397,N_4274);
and U4448 (N_4448,N_4290,N_4349);
and U4449 (N_4449,N_4281,N_4303);
or U4450 (N_4450,N_4232,N_4380);
nand U4451 (N_4451,N_4247,N_4394);
nor U4452 (N_4452,N_4379,N_4278);
and U4453 (N_4453,N_4220,N_4241);
nor U4454 (N_4454,N_4258,N_4366);
xnor U4455 (N_4455,N_4224,N_4302);
or U4456 (N_4456,N_4202,N_4204);
nand U4457 (N_4457,N_4285,N_4321);
nor U4458 (N_4458,N_4351,N_4325);
nor U4459 (N_4459,N_4270,N_4307);
xor U4460 (N_4460,N_4266,N_4353);
nand U4461 (N_4461,N_4341,N_4372);
and U4462 (N_4462,N_4332,N_4398);
or U4463 (N_4463,N_4389,N_4200);
xor U4464 (N_4464,N_4355,N_4289);
xnor U4465 (N_4465,N_4210,N_4373);
nand U4466 (N_4466,N_4263,N_4323);
or U4467 (N_4467,N_4231,N_4374);
and U4468 (N_4468,N_4237,N_4283);
nor U4469 (N_4469,N_4338,N_4228);
nand U4470 (N_4470,N_4253,N_4234);
nand U4471 (N_4471,N_4310,N_4359);
xor U4472 (N_4472,N_4315,N_4358);
and U4473 (N_4473,N_4335,N_4365);
nand U4474 (N_4474,N_4284,N_4209);
or U4475 (N_4475,N_4330,N_4271);
or U4476 (N_4476,N_4392,N_4357);
or U4477 (N_4477,N_4384,N_4261);
nor U4478 (N_4478,N_4206,N_4269);
xnor U4479 (N_4479,N_4250,N_4381);
nand U4480 (N_4480,N_4246,N_4388);
nand U4481 (N_4481,N_4367,N_4377);
nand U4482 (N_4482,N_4331,N_4369);
nor U4483 (N_4483,N_4363,N_4265);
nand U4484 (N_4484,N_4240,N_4227);
nor U4485 (N_4485,N_4298,N_4296);
or U4486 (N_4486,N_4334,N_4343);
nor U4487 (N_4487,N_4306,N_4375);
nor U4488 (N_4488,N_4382,N_4318);
and U4489 (N_4489,N_4286,N_4248);
xnor U4490 (N_4490,N_4288,N_4244);
nand U4491 (N_4491,N_4207,N_4287);
and U4492 (N_4492,N_4217,N_4235);
or U4493 (N_4493,N_4243,N_4327);
or U4494 (N_4494,N_4280,N_4316);
xnor U4495 (N_4495,N_4328,N_4340);
nand U4496 (N_4496,N_4370,N_4317);
xor U4497 (N_4497,N_4386,N_4313);
xor U4498 (N_4498,N_4267,N_4399);
and U4499 (N_4499,N_4236,N_4245);
nand U4500 (N_4500,N_4394,N_4341);
xnor U4501 (N_4501,N_4257,N_4256);
xor U4502 (N_4502,N_4241,N_4292);
or U4503 (N_4503,N_4213,N_4328);
or U4504 (N_4504,N_4329,N_4294);
nor U4505 (N_4505,N_4347,N_4269);
or U4506 (N_4506,N_4210,N_4244);
and U4507 (N_4507,N_4246,N_4241);
xnor U4508 (N_4508,N_4239,N_4355);
and U4509 (N_4509,N_4355,N_4206);
xnor U4510 (N_4510,N_4244,N_4281);
and U4511 (N_4511,N_4290,N_4323);
nor U4512 (N_4512,N_4218,N_4315);
xnor U4513 (N_4513,N_4361,N_4291);
nor U4514 (N_4514,N_4280,N_4248);
nand U4515 (N_4515,N_4261,N_4263);
and U4516 (N_4516,N_4277,N_4266);
and U4517 (N_4517,N_4376,N_4318);
and U4518 (N_4518,N_4361,N_4221);
nand U4519 (N_4519,N_4386,N_4295);
xor U4520 (N_4520,N_4231,N_4268);
or U4521 (N_4521,N_4355,N_4244);
nand U4522 (N_4522,N_4215,N_4261);
or U4523 (N_4523,N_4358,N_4208);
and U4524 (N_4524,N_4373,N_4312);
nor U4525 (N_4525,N_4203,N_4375);
nand U4526 (N_4526,N_4299,N_4290);
or U4527 (N_4527,N_4313,N_4237);
or U4528 (N_4528,N_4250,N_4353);
and U4529 (N_4529,N_4257,N_4231);
xor U4530 (N_4530,N_4399,N_4329);
nor U4531 (N_4531,N_4236,N_4311);
or U4532 (N_4532,N_4205,N_4233);
xnor U4533 (N_4533,N_4295,N_4374);
and U4534 (N_4534,N_4292,N_4389);
or U4535 (N_4535,N_4252,N_4290);
xnor U4536 (N_4536,N_4205,N_4281);
or U4537 (N_4537,N_4312,N_4219);
and U4538 (N_4538,N_4311,N_4318);
xor U4539 (N_4539,N_4383,N_4321);
nand U4540 (N_4540,N_4335,N_4375);
xnor U4541 (N_4541,N_4351,N_4389);
nor U4542 (N_4542,N_4293,N_4234);
xnor U4543 (N_4543,N_4325,N_4244);
nor U4544 (N_4544,N_4208,N_4235);
or U4545 (N_4545,N_4216,N_4318);
nor U4546 (N_4546,N_4215,N_4219);
or U4547 (N_4547,N_4383,N_4309);
xor U4548 (N_4548,N_4375,N_4269);
nand U4549 (N_4549,N_4315,N_4312);
xor U4550 (N_4550,N_4220,N_4250);
nor U4551 (N_4551,N_4293,N_4257);
and U4552 (N_4552,N_4288,N_4266);
nand U4553 (N_4553,N_4240,N_4290);
or U4554 (N_4554,N_4260,N_4326);
xor U4555 (N_4555,N_4261,N_4237);
and U4556 (N_4556,N_4252,N_4328);
or U4557 (N_4557,N_4351,N_4361);
or U4558 (N_4558,N_4331,N_4334);
or U4559 (N_4559,N_4243,N_4366);
nand U4560 (N_4560,N_4247,N_4314);
nand U4561 (N_4561,N_4283,N_4311);
xnor U4562 (N_4562,N_4252,N_4347);
or U4563 (N_4563,N_4247,N_4266);
nor U4564 (N_4564,N_4312,N_4284);
xnor U4565 (N_4565,N_4336,N_4377);
xnor U4566 (N_4566,N_4359,N_4358);
or U4567 (N_4567,N_4230,N_4239);
nand U4568 (N_4568,N_4364,N_4233);
and U4569 (N_4569,N_4398,N_4211);
nor U4570 (N_4570,N_4277,N_4200);
and U4571 (N_4571,N_4336,N_4233);
and U4572 (N_4572,N_4318,N_4260);
and U4573 (N_4573,N_4386,N_4263);
nor U4574 (N_4574,N_4201,N_4336);
xnor U4575 (N_4575,N_4259,N_4333);
xnor U4576 (N_4576,N_4348,N_4380);
and U4577 (N_4577,N_4354,N_4210);
and U4578 (N_4578,N_4277,N_4235);
nor U4579 (N_4579,N_4247,N_4281);
nand U4580 (N_4580,N_4397,N_4293);
nand U4581 (N_4581,N_4311,N_4394);
nor U4582 (N_4582,N_4261,N_4227);
xnor U4583 (N_4583,N_4393,N_4388);
xor U4584 (N_4584,N_4211,N_4282);
nor U4585 (N_4585,N_4243,N_4279);
and U4586 (N_4586,N_4215,N_4396);
and U4587 (N_4587,N_4309,N_4279);
or U4588 (N_4588,N_4396,N_4210);
nor U4589 (N_4589,N_4328,N_4215);
or U4590 (N_4590,N_4231,N_4334);
nand U4591 (N_4591,N_4397,N_4309);
nor U4592 (N_4592,N_4228,N_4336);
xor U4593 (N_4593,N_4260,N_4249);
xnor U4594 (N_4594,N_4211,N_4371);
nor U4595 (N_4595,N_4279,N_4304);
nor U4596 (N_4596,N_4373,N_4252);
or U4597 (N_4597,N_4252,N_4379);
xnor U4598 (N_4598,N_4343,N_4324);
xor U4599 (N_4599,N_4222,N_4385);
xor U4600 (N_4600,N_4539,N_4578);
and U4601 (N_4601,N_4452,N_4460);
nor U4602 (N_4602,N_4484,N_4479);
and U4603 (N_4603,N_4419,N_4449);
nor U4604 (N_4604,N_4402,N_4561);
or U4605 (N_4605,N_4410,N_4577);
xnor U4606 (N_4606,N_4424,N_4517);
nor U4607 (N_4607,N_4412,N_4499);
nand U4608 (N_4608,N_4508,N_4477);
and U4609 (N_4609,N_4551,N_4450);
and U4610 (N_4610,N_4458,N_4557);
or U4611 (N_4611,N_4533,N_4514);
nand U4612 (N_4612,N_4409,N_4573);
nand U4613 (N_4613,N_4475,N_4437);
nand U4614 (N_4614,N_4520,N_4465);
or U4615 (N_4615,N_4583,N_4505);
or U4616 (N_4616,N_4472,N_4589);
xor U4617 (N_4617,N_4441,N_4525);
or U4618 (N_4618,N_4459,N_4552);
and U4619 (N_4619,N_4495,N_4462);
or U4620 (N_4620,N_4540,N_4426);
and U4621 (N_4621,N_4554,N_4575);
nor U4622 (N_4622,N_4509,N_4443);
nand U4623 (N_4623,N_4457,N_4558);
nor U4624 (N_4624,N_4580,N_4444);
and U4625 (N_4625,N_4598,N_4474);
nand U4626 (N_4626,N_4469,N_4478);
nand U4627 (N_4627,N_4454,N_4564);
and U4628 (N_4628,N_4542,N_4581);
xnor U4629 (N_4629,N_4430,N_4545);
xor U4630 (N_4630,N_4556,N_4538);
nor U4631 (N_4631,N_4497,N_4596);
and U4632 (N_4632,N_4595,N_4588);
and U4633 (N_4633,N_4547,N_4515);
xnor U4634 (N_4634,N_4486,N_4492);
and U4635 (N_4635,N_4476,N_4512);
and U4636 (N_4636,N_4500,N_4587);
nand U4637 (N_4637,N_4593,N_4591);
nor U4638 (N_4638,N_4467,N_4543);
xnor U4639 (N_4639,N_4516,N_4507);
and U4640 (N_4640,N_4511,N_4524);
nand U4641 (N_4641,N_4544,N_4546);
nor U4642 (N_4642,N_4572,N_4416);
and U4643 (N_4643,N_4471,N_4521);
nor U4644 (N_4644,N_4565,N_4406);
nor U4645 (N_4645,N_4548,N_4498);
or U4646 (N_4646,N_4429,N_4481);
nor U4647 (N_4647,N_4405,N_4582);
and U4648 (N_4648,N_4493,N_4563);
nand U4649 (N_4649,N_4504,N_4531);
nand U4650 (N_4650,N_4599,N_4448);
nand U4651 (N_4651,N_4488,N_4569);
or U4652 (N_4652,N_4442,N_4527);
nand U4653 (N_4653,N_4529,N_4526);
nand U4654 (N_4654,N_4464,N_4480);
nor U4655 (N_4655,N_4560,N_4528);
or U4656 (N_4656,N_4550,N_4483);
or U4657 (N_4657,N_4435,N_4559);
nand U4658 (N_4658,N_4463,N_4453);
and U4659 (N_4659,N_4473,N_4534);
nor U4660 (N_4660,N_4414,N_4567);
or U4661 (N_4661,N_4418,N_4536);
nand U4662 (N_4662,N_4468,N_4502);
or U4663 (N_4663,N_4438,N_4420);
nor U4664 (N_4664,N_4425,N_4553);
nor U4665 (N_4665,N_4549,N_4571);
and U4666 (N_4666,N_4407,N_4446);
and U4667 (N_4667,N_4482,N_4413);
nand U4668 (N_4668,N_4506,N_4592);
or U4669 (N_4669,N_4594,N_4456);
nand U4670 (N_4670,N_4421,N_4586);
and U4671 (N_4671,N_4401,N_4439);
xnor U4672 (N_4672,N_4494,N_4487);
nor U4673 (N_4673,N_4496,N_4518);
xor U4674 (N_4674,N_4451,N_4510);
xor U4675 (N_4675,N_4503,N_4447);
and U4676 (N_4676,N_4574,N_4562);
nor U4677 (N_4677,N_4436,N_4585);
or U4678 (N_4678,N_4568,N_4555);
and U4679 (N_4679,N_4522,N_4440);
and U4680 (N_4680,N_4490,N_4432);
and U4681 (N_4681,N_4422,N_4434);
or U4682 (N_4682,N_4489,N_4427);
and U4683 (N_4683,N_4535,N_4576);
nor U4684 (N_4684,N_4433,N_4423);
nand U4685 (N_4685,N_4579,N_4530);
xnor U4686 (N_4686,N_4411,N_4570);
and U4687 (N_4687,N_4597,N_4455);
and U4688 (N_4688,N_4400,N_4403);
nand U4689 (N_4689,N_4584,N_4417);
nor U4690 (N_4690,N_4537,N_4501);
nor U4691 (N_4691,N_4415,N_4513);
and U4692 (N_4692,N_4404,N_4523);
and U4693 (N_4693,N_4590,N_4541);
xor U4694 (N_4694,N_4466,N_4566);
or U4695 (N_4695,N_4461,N_4431);
and U4696 (N_4696,N_4428,N_4470);
nand U4697 (N_4697,N_4491,N_4408);
or U4698 (N_4698,N_4532,N_4445);
or U4699 (N_4699,N_4485,N_4519);
nand U4700 (N_4700,N_4570,N_4443);
or U4701 (N_4701,N_4518,N_4443);
or U4702 (N_4702,N_4453,N_4544);
nand U4703 (N_4703,N_4574,N_4534);
and U4704 (N_4704,N_4570,N_4506);
and U4705 (N_4705,N_4456,N_4472);
and U4706 (N_4706,N_4414,N_4560);
and U4707 (N_4707,N_4565,N_4461);
nand U4708 (N_4708,N_4574,N_4419);
or U4709 (N_4709,N_4488,N_4571);
nand U4710 (N_4710,N_4451,N_4421);
or U4711 (N_4711,N_4448,N_4456);
xnor U4712 (N_4712,N_4460,N_4412);
or U4713 (N_4713,N_4589,N_4467);
and U4714 (N_4714,N_4482,N_4523);
or U4715 (N_4715,N_4400,N_4462);
nand U4716 (N_4716,N_4486,N_4498);
nor U4717 (N_4717,N_4480,N_4425);
and U4718 (N_4718,N_4445,N_4442);
nor U4719 (N_4719,N_4591,N_4509);
and U4720 (N_4720,N_4595,N_4483);
or U4721 (N_4721,N_4479,N_4522);
nand U4722 (N_4722,N_4549,N_4538);
and U4723 (N_4723,N_4558,N_4404);
nand U4724 (N_4724,N_4404,N_4557);
or U4725 (N_4725,N_4471,N_4535);
or U4726 (N_4726,N_4547,N_4516);
or U4727 (N_4727,N_4501,N_4444);
and U4728 (N_4728,N_4485,N_4504);
nor U4729 (N_4729,N_4448,N_4547);
xor U4730 (N_4730,N_4449,N_4479);
or U4731 (N_4731,N_4596,N_4404);
nand U4732 (N_4732,N_4451,N_4580);
nor U4733 (N_4733,N_4420,N_4593);
nor U4734 (N_4734,N_4424,N_4479);
xor U4735 (N_4735,N_4563,N_4467);
or U4736 (N_4736,N_4547,N_4592);
nor U4737 (N_4737,N_4575,N_4556);
nand U4738 (N_4738,N_4460,N_4583);
nor U4739 (N_4739,N_4477,N_4566);
xnor U4740 (N_4740,N_4573,N_4484);
nand U4741 (N_4741,N_4416,N_4598);
nor U4742 (N_4742,N_4571,N_4598);
nand U4743 (N_4743,N_4425,N_4507);
xnor U4744 (N_4744,N_4414,N_4472);
nor U4745 (N_4745,N_4500,N_4564);
and U4746 (N_4746,N_4474,N_4576);
nor U4747 (N_4747,N_4428,N_4579);
nand U4748 (N_4748,N_4562,N_4592);
or U4749 (N_4749,N_4579,N_4438);
xor U4750 (N_4750,N_4587,N_4401);
nand U4751 (N_4751,N_4508,N_4478);
and U4752 (N_4752,N_4555,N_4472);
xor U4753 (N_4753,N_4453,N_4547);
and U4754 (N_4754,N_4580,N_4516);
nor U4755 (N_4755,N_4453,N_4534);
nor U4756 (N_4756,N_4463,N_4588);
and U4757 (N_4757,N_4594,N_4423);
or U4758 (N_4758,N_4504,N_4570);
nand U4759 (N_4759,N_4504,N_4559);
xnor U4760 (N_4760,N_4465,N_4524);
or U4761 (N_4761,N_4566,N_4514);
nand U4762 (N_4762,N_4445,N_4418);
nand U4763 (N_4763,N_4424,N_4549);
xor U4764 (N_4764,N_4544,N_4408);
and U4765 (N_4765,N_4524,N_4546);
nand U4766 (N_4766,N_4431,N_4506);
nand U4767 (N_4767,N_4562,N_4561);
and U4768 (N_4768,N_4458,N_4570);
xnor U4769 (N_4769,N_4501,N_4569);
and U4770 (N_4770,N_4577,N_4412);
nor U4771 (N_4771,N_4520,N_4400);
xnor U4772 (N_4772,N_4517,N_4415);
xor U4773 (N_4773,N_4475,N_4561);
nor U4774 (N_4774,N_4470,N_4496);
xnor U4775 (N_4775,N_4442,N_4578);
or U4776 (N_4776,N_4400,N_4574);
or U4777 (N_4777,N_4498,N_4578);
xnor U4778 (N_4778,N_4500,N_4451);
xnor U4779 (N_4779,N_4460,N_4547);
nand U4780 (N_4780,N_4541,N_4574);
and U4781 (N_4781,N_4542,N_4576);
and U4782 (N_4782,N_4405,N_4453);
and U4783 (N_4783,N_4568,N_4561);
nor U4784 (N_4784,N_4588,N_4445);
and U4785 (N_4785,N_4502,N_4427);
nor U4786 (N_4786,N_4475,N_4598);
xor U4787 (N_4787,N_4417,N_4459);
nor U4788 (N_4788,N_4527,N_4499);
xor U4789 (N_4789,N_4447,N_4508);
and U4790 (N_4790,N_4491,N_4401);
and U4791 (N_4791,N_4501,N_4475);
or U4792 (N_4792,N_4432,N_4473);
nor U4793 (N_4793,N_4545,N_4443);
nand U4794 (N_4794,N_4440,N_4463);
nor U4795 (N_4795,N_4497,N_4403);
and U4796 (N_4796,N_4470,N_4408);
xnor U4797 (N_4797,N_4553,N_4449);
nand U4798 (N_4798,N_4588,N_4407);
or U4799 (N_4799,N_4549,N_4409);
nand U4800 (N_4800,N_4774,N_4621);
nand U4801 (N_4801,N_4703,N_4605);
and U4802 (N_4802,N_4637,N_4799);
and U4803 (N_4803,N_4602,N_4796);
or U4804 (N_4804,N_4770,N_4677);
nor U4805 (N_4805,N_4624,N_4603);
nand U4806 (N_4806,N_4751,N_4639);
xnor U4807 (N_4807,N_4693,N_4660);
nand U4808 (N_4808,N_4626,N_4788);
nand U4809 (N_4809,N_4680,N_4606);
nand U4810 (N_4810,N_4627,N_4675);
nand U4811 (N_4811,N_4750,N_4792);
and U4812 (N_4812,N_4689,N_4729);
or U4813 (N_4813,N_4704,N_4659);
xor U4814 (N_4814,N_4688,N_4607);
or U4815 (N_4815,N_4611,N_4628);
and U4816 (N_4816,N_4712,N_4658);
nand U4817 (N_4817,N_4647,N_4775);
nand U4818 (N_4818,N_4779,N_4697);
xnor U4819 (N_4819,N_4715,N_4630);
xnor U4820 (N_4820,N_4650,N_4694);
xnor U4821 (N_4821,N_4633,N_4777);
or U4822 (N_4822,N_4778,N_4634);
nand U4823 (N_4823,N_4696,N_4731);
nand U4824 (N_4824,N_4684,N_4641);
or U4825 (N_4825,N_4601,N_4657);
nor U4826 (N_4826,N_4743,N_4656);
xor U4827 (N_4827,N_4764,N_4625);
and U4828 (N_4828,N_4719,N_4752);
xor U4829 (N_4829,N_4683,N_4669);
nand U4830 (N_4830,N_4717,N_4789);
nor U4831 (N_4831,N_4762,N_4672);
or U4832 (N_4832,N_4766,N_4609);
nand U4833 (N_4833,N_4741,N_4784);
and U4834 (N_4834,N_4685,N_4645);
nand U4835 (N_4835,N_4758,N_4738);
xnor U4836 (N_4836,N_4765,N_4782);
or U4837 (N_4837,N_4727,N_4620);
xor U4838 (N_4838,N_4691,N_4600);
nor U4839 (N_4839,N_4733,N_4768);
or U4840 (N_4840,N_4740,N_4746);
xnor U4841 (N_4841,N_4776,N_4797);
xnor U4842 (N_4842,N_4739,N_4794);
xor U4843 (N_4843,N_4686,N_4726);
xnor U4844 (N_4844,N_4711,N_4612);
nand U4845 (N_4845,N_4749,N_4618);
or U4846 (N_4846,N_4616,N_4720);
nor U4847 (N_4847,N_4674,N_4610);
xor U4848 (N_4848,N_4747,N_4723);
and U4849 (N_4849,N_4663,N_4702);
nand U4850 (N_4850,N_4773,N_4724);
nand U4851 (N_4851,N_4635,N_4756);
nand U4852 (N_4852,N_4662,N_4783);
or U4853 (N_4853,N_4757,N_4709);
xnor U4854 (N_4854,N_4640,N_4692);
and U4855 (N_4855,N_4732,N_4654);
nor U4856 (N_4856,N_4786,N_4771);
xnor U4857 (N_4857,N_4655,N_4695);
and U4858 (N_4858,N_4636,N_4714);
nor U4859 (N_4859,N_4622,N_4613);
xnor U4860 (N_4860,N_4676,N_4793);
nand U4861 (N_4861,N_4632,N_4795);
and U4862 (N_4862,N_4615,N_4679);
xnor U4863 (N_4863,N_4748,N_4608);
or U4864 (N_4864,N_4707,N_4665);
nor U4865 (N_4865,N_4755,N_4742);
nand U4866 (N_4866,N_4699,N_4767);
or U4867 (N_4867,N_4706,N_4629);
and U4868 (N_4868,N_4798,N_4698);
and U4869 (N_4869,N_4721,N_4614);
nand U4870 (N_4870,N_4631,N_4744);
nand U4871 (N_4871,N_4780,N_4648);
nor U4872 (N_4872,N_4646,N_4690);
xnor U4873 (N_4873,N_4763,N_4666);
and U4874 (N_4874,N_4772,N_4759);
xor U4875 (N_4875,N_4644,N_4701);
and U4876 (N_4876,N_4678,N_4673);
nor U4877 (N_4877,N_4754,N_4725);
or U4878 (N_4878,N_4781,N_4664);
and U4879 (N_4879,N_4745,N_4728);
nand U4880 (N_4880,N_4787,N_4713);
and U4881 (N_4881,N_4652,N_4785);
nand U4882 (N_4882,N_4643,N_4604);
nor U4883 (N_4883,N_4661,N_4653);
xor U4884 (N_4884,N_4700,N_4722);
or U4885 (N_4885,N_4737,N_4667);
or U4886 (N_4886,N_4791,N_4790);
nor U4887 (N_4887,N_4769,N_4671);
and U4888 (N_4888,N_4670,N_4735);
nand U4889 (N_4889,N_4705,N_4760);
or U4890 (N_4890,N_4710,N_4619);
and U4891 (N_4891,N_4716,N_4753);
nor U4892 (N_4892,N_4734,N_4681);
or U4893 (N_4893,N_4708,N_4623);
xnor U4894 (N_4894,N_4736,N_4682);
and U4895 (N_4895,N_4617,N_4687);
nand U4896 (N_4896,N_4638,N_4718);
xor U4897 (N_4897,N_4642,N_4730);
nand U4898 (N_4898,N_4761,N_4651);
nor U4899 (N_4899,N_4649,N_4668);
and U4900 (N_4900,N_4615,N_4632);
nor U4901 (N_4901,N_4793,N_4758);
or U4902 (N_4902,N_4707,N_4661);
and U4903 (N_4903,N_4792,N_4654);
and U4904 (N_4904,N_4635,N_4709);
and U4905 (N_4905,N_4695,N_4747);
or U4906 (N_4906,N_4637,N_4708);
or U4907 (N_4907,N_4768,N_4782);
nor U4908 (N_4908,N_4752,N_4683);
or U4909 (N_4909,N_4763,N_4778);
and U4910 (N_4910,N_4723,N_4602);
or U4911 (N_4911,N_4670,N_4745);
nor U4912 (N_4912,N_4792,N_4610);
nor U4913 (N_4913,N_4648,N_4727);
nor U4914 (N_4914,N_4697,N_4626);
or U4915 (N_4915,N_4723,N_4621);
and U4916 (N_4916,N_4734,N_4662);
or U4917 (N_4917,N_4707,N_4708);
xnor U4918 (N_4918,N_4738,N_4636);
or U4919 (N_4919,N_4767,N_4682);
or U4920 (N_4920,N_4627,N_4760);
and U4921 (N_4921,N_4714,N_4606);
xnor U4922 (N_4922,N_4765,N_4604);
nand U4923 (N_4923,N_4684,N_4701);
xnor U4924 (N_4924,N_4696,N_4797);
nor U4925 (N_4925,N_4737,N_4678);
nor U4926 (N_4926,N_4742,N_4791);
and U4927 (N_4927,N_4660,N_4732);
or U4928 (N_4928,N_4727,N_4659);
nor U4929 (N_4929,N_4682,N_4664);
and U4930 (N_4930,N_4696,N_4637);
and U4931 (N_4931,N_4610,N_4669);
xor U4932 (N_4932,N_4648,N_4775);
nand U4933 (N_4933,N_4793,N_4786);
xor U4934 (N_4934,N_4792,N_4788);
and U4935 (N_4935,N_4681,N_4697);
nand U4936 (N_4936,N_4782,N_4761);
and U4937 (N_4937,N_4687,N_4698);
and U4938 (N_4938,N_4685,N_4646);
nor U4939 (N_4939,N_4649,N_4688);
xor U4940 (N_4940,N_4718,N_4627);
xnor U4941 (N_4941,N_4769,N_4787);
nor U4942 (N_4942,N_4694,N_4604);
nand U4943 (N_4943,N_4719,N_4644);
and U4944 (N_4944,N_4708,N_4618);
xnor U4945 (N_4945,N_4626,N_4724);
and U4946 (N_4946,N_4791,N_4797);
or U4947 (N_4947,N_4616,N_4614);
nor U4948 (N_4948,N_4630,N_4605);
nor U4949 (N_4949,N_4749,N_4714);
and U4950 (N_4950,N_4747,N_4749);
or U4951 (N_4951,N_4671,N_4720);
nand U4952 (N_4952,N_4655,N_4633);
nor U4953 (N_4953,N_4737,N_4766);
nand U4954 (N_4954,N_4741,N_4690);
or U4955 (N_4955,N_4690,N_4751);
xor U4956 (N_4956,N_4687,N_4674);
and U4957 (N_4957,N_4729,N_4686);
nand U4958 (N_4958,N_4772,N_4680);
or U4959 (N_4959,N_4626,N_4702);
nor U4960 (N_4960,N_4787,N_4705);
nor U4961 (N_4961,N_4718,N_4760);
nand U4962 (N_4962,N_4629,N_4707);
nor U4963 (N_4963,N_4601,N_4755);
nor U4964 (N_4964,N_4717,N_4659);
and U4965 (N_4965,N_4660,N_4755);
nor U4966 (N_4966,N_4679,N_4692);
or U4967 (N_4967,N_4673,N_4799);
nand U4968 (N_4968,N_4761,N_4747);
nor U4969 (N_4969,N_4630,N_4672);
xor U4970 (N_4970,N_4621,N_4620);
and U4971 (N_4971,N_4779,N_4787);
or U4972 (N_4972,N_4644,N_4794);
nor U4973 (N_4973,N_4726,N_4774);
xor U4974 (N_4974,N_4646,N_4718);
xnor U4975 (N_4975,N_4799,N_4755);
nor U4976 (N_4976,N_4710,N_4653);
or U4977 (N_4977,N_4601,N_4772);
nor U4978 (N_4978,N_4770,N_4737);
xor U4979 (N_4979,N_4673,N_4631);
nand U4980 (N_4980,N_4767,N_4670);
nand U4981 (N_4981,N_4764,N_4776);
nand U4982 (N_4982,N_4762,N_4665);
and U4983 (N_4983,N_4679,N_4639);
or U4984 (N_4984,N_4669,N_4714);
nand U4985 (N_4985,N_4768,N_4629);
xor U4986 (N_4986,N_4709,N_4784);
nor U4987 (N_4987,N_4754,N_4649);
and U4988 (N_4988,N_4669,N_4787);
nand U4989 (N_4989,N_4719,N_4794);
or U4990 (N_4990,N_4609,N_4664);
xnor U4991 (N_4991,N_4769,N_4651);
nor U4992 (N_4992,N_4602,N_4662);
or U4993 (N_4993,N_4752,N_4727);
nand U4994 (N_4994,N_4748,N_4695);
xnor U4995 (N_4995,N_4738,N_4788);
or U4996 (N_4996,N_4628,N_4758);
or U4997 (N_4997,N_4634,N_4738);
nand U4998 (N_4998,N_4627,N_4683);
nand U4999 (N_4999,N_4692,N_4682);
or U5000 (N_5000,N_4970,N_4911);
and U5001 (N_5001,N_4804,N_4841);
nor U5002 (N_5002,N_4820,N_4950);
nand U5003 (N_5003,N_4846,N_4964);
or U5004 (N_5004,N_4868,N_4811);
and U5005 (N_5005,N_4853,N_4848);
and U5006 (N_5006,N_4844,N_4893);
nand U5007 (N_5007,N_4997,N_4818);
or U5008 (N_5008,N_4819,N_4895);
nor U5009 (N_5009,N_4887,N_4927);
nor U5010 (N_5010,N_4917,N_4965);
nand U5011 (N_5011,N_4978,N_4913);
nor U5012 (N_5012,N_4945,N_4828);
nand U5013 (N_5013,N_4956,N_4886);
or U5014 (N_5014,N_4881,N_4892);
and U5015 (N_5015,N_4930,N_4986);
and U5016 (N_5016,N_4949,N_4875);
or U5017 (N_5017,N_4829,N_4941);
xnor U5018 (N_5018,N_4972,N_4873);
and U5019 (N_5019,N_4865,N_4852);
nor U5020 (N_5020,N_4864,N_4889);
and U5021 (N_5021,N_4810,N_4981);
or U5022 (N_5022,N_4826,N_4954);
nor U5023 (N_5023,N_4832,N_4980);
xor U5024 (N_5024,N_4938,N_4903);
nand U5025 (N_5025,N_4993,N_4976);
xnor U5026 (N_5026,N_4837,N_4948);
or U5027 (N_5027,N_4975,N_4859);
or U5028 (N_5028,N_4883,N_4998);
xnor U5029 (N_5029,N_4932,N_4985);
and U5030 (N_5030,N_4928,N_4940);
or U5031 (N_5031,N_4803,N_4925);
or U5032 (N_5032,N_4802,N_4900);
nand U5033 (N_5033,N_4880,N_4856);
nor U5034 (N_5034,N_4860,N_4821);
or U5035 (N_5035,N_4806,N_4935);
nor U5036 (N_5036,N_4874,N_4984);
or U5037 (N_5037,N_4918,N_4952);
and U5038 (N_5038,N_4987,N_4813);
and U5039 (N_5039,N_4834,N_4857);
and U5040 (N_5040,N_4946,N_4891);
nand U5041 (N_5041,N_4801,N_4990);
or U5042 (N_5042,N_4825,N_4924);
xor U5043 (N_5043,N_4808,N_4833);
and U5044 (N_5044,N_4850,N_4899);
xnor U5045 (N_5045,N_4914,N_4877);
nor U5046 (N_5046,N_4912,N_4831);
xnor U5047 (N_5047,N_4835,N_4994);
nor U5048 (N_5048,N_4977,N_4896);
or U5049 (N_5049,N_4839,N_4996);
and U5050 (N_5050,N_4906,N_4840);
or U5051 (N_5051,N_4955,N_4888);
nor U5052 (N_5052,N_4807,N_4960);
nand U5053 (N_5053,N_4910,N_4897);
or U5054 (N_5054,N_4805,N_4992);
nand U5055 (N_5055,N_4885,N_4999);
nand U5056 (N_5056,N_4929,N_4947);
xor U5057 (N_5057,N_4971,N_4816);
nor U5058 (N_5058,N_4974,N_4812);
and U5059 (N_5059,N_4869,N_4942);
nand U5060 (N_5060,N_4923,N_4824);
or U5061 (N_5061,N_4894,N_4855);
and U5062 (N_5062,N_4890,N_4908);
nor U5063 (N_5063,N_4863,N_4836);
or U5064 (N_5064,N_4934,N_4926);
or U5065 (N_5065,N_4962,N_4838);
nand U5066 (N_5066,N_4961,N_4915);
nor U5067 (N_5067,N_4901,N_4866);
nor U5068 (N_5068,N_4827,N_4854);
nor U5069 (N_5069,N_4872,N_4876);
and U5070 (N_5070,N_4862,N_4989);
nand U5071 (N_5071,N_4870,N_4867);
or U5072 (N_5072,N_4815,N_4861);
nand U5073 (N_5073,N_4902,N_4943);
nor U5074 (N_5074,N_4982,N_4898);
xnor U5075 (N_5075,N_4830,N_4937);
nor U5076 (N_5076,N_4871,N_4951);
nor U5077 (N_5077,N_4973,N_4845);
or U5078 (N_5078,N_4967,N_4843);
nand U5079 (N_5079,N_4847,N_4968);
nor U5080 (N_5080,N_4969,N_4966);
nor U5081 (N_5081,N_4983,N_4988);
xnor U5082 (N_5082,N_4878,N_4822);
xor U5083 (N_5083,N_4979,N_4842);
nand U5084 (N_5084,N_4959,N_4922);
xor U5085 (N_5085,N_4944,N_4907);
or U5086 (N_5086,N_4817,N_4936);
nor U5087 (N_5087,N_4931,N_4958);
nand U5088 (N_5088,N_4916,N_4920);
and U5089 (N_5089,N_4823,N_4995);
nand U5090 (N_5090,N_4882,N_4905);
xor U5091 (N_5091,N_4939,N_4858);
or U5092 (N_5092,N_4909,N_4814);
and U5093 (N_5093,N_4921,N_4991);
nand U5094 (N_5094,N_4851,N_4809);
xnor U5095 (N_5095,N_4904,N_4957);
and U5096 (N_5096,N_4849,N_4884);
nand U5097 (N_5097,N_4879,N_4933);
or U5098 (N_5098,N_4953,N_4800);
or U5099 (N_5099,N_4963,N_4919);
nand U5100 (N_5100,N_4843,N_4808);
xor U5101 (N_5101,N_4870,N_4853);
nand U5102 (N_5102,N_4958,N_4946);
nor U5103 (N_5103,N_4980,N_4892);
or U5104 (N_5104,N_4889,N_4871);
nand U5105 (N_5105,N_4995,N_4905);
and U5106 (N_5106,N_4832,N_4875);
and U5107 (N_5107,N_4800,N_4884);
nor U5108 (N_5108,N_4932,N_4831);
or U5109 (N_5109,N_4979,N_4971);
and U5110 (N_5110,N_4983,N_4884);
or U5111 (N_5111,N_4836,N_4811);
xor U5112 (N_5112,N_4963,N_4844);
nor U5113 (N_5113,N_4944,N_4975);
nand U5114 (N_5114,N_4909,N_4940);
nor U5115 (N_5115,N_4843,N_4991);
nor U5116 (N_5116,N_4828,N_4868);
nand U5117 (N_5117,N_4894,N_4901);
nand U5118 (N_5118,N_4997,N_4865);
and U5119 (N_5119,N_4957,N_4959);
nor U5120 (N_5120,N_4892,N_4857);
nor U5121 (N_5121,N_4803,N_4996);
or U5122 (N_5122,N_4952,N_4832);
and U5123 (N_5123,N_4933,N_4857);
and U5124 (N_5124,N_4987,N_4873);
or U5125 (N_5125,N_4912,N_4913);
and U5126 (N_5126,N_4978,N_4962);
or U5127 (N_5127,N_4916,N_4840);
nand U5128 (N_5128,N_4902,N_4946);
and U5129 (N_5129,N_4995,N_4893);
and U5130 (N_5130,N_4853,N_4810);
nand U5131 (N_5131,N_4801,N_4821);
and U5132 (N_5132,N_4853,N_4872);
nand U5133 (N_5133,N_4909,N_4934);
and U5134 (N_5134,N_4879,N_4839);
nand U5135 (N_5135,N_4846,N_4946);
nor U5136 (N_5136,N_4979,N_4858);
xnor U5137 (N_5137,N_4994,N_4898);
and U5138 (N_5138,N_4907,N_4845);
xor U5139 (N_5139,N_4820,N_4934);
xnor U5140 (N_5140,N_4858,N_4963);
nand U5141 (N_5141,N_4935,N_4858);
nor U5142 (N_5142,N_4998,N_4873);
and U5143 (N_5143,N_4823,N_4805);
and U5144 (N_5144,N_4922,N_4936);
nand U5145 (N_5145,N_4943,N_4885);
xor U5146 (N_5146,N_4947,N_4925);
xnor U5147 (N_5147,N_4939,N_4815);
nand U5148 (N_5148,N_4885,N_4883);
and U5149 (N_5149,N_4910,N_4873);
and U5150 (N_5150,N_4905,N_4979);
nand U5151 (N_5151,N_4825,N_4827);
xor U5152 (N_5152,N_4965,N_4940);
and U5153 (N_5153,N_4940,N_4835);
nor U5154 (N_5154,N_4903,N_4955);
nor U5155 (N_5155,N_4910,N_4855);
or U5156 (N_5156,N_4922,N_4862);
and U5157 (N_5157,N_4923,N_4870);
xor U5158 (N_5158,N_4990,N_4803);
nor U5159 (N_5159,N_4850,N_4821);
nor U5160 (N_5160,N_4907,N_4889);
or U5161 (N_5161,N_4925,N_4863);
and U5162 (N_5162,N_4916,N_4972);
nor U5163 (N_5163,N_4958,N_4922);
and U5164 (N_5164,N_4907,N_4859);
or U5165 (N_5165,N_4932,N_4881);
nand U5166 (N_5166,N_4970,N_4931);
or U5167 (N_5167,N_4861,N_4982);
or U5168 (N_5168,N_4976,N_4972);
or U5169 (N_5169,N_4915,N_4960);
nand U5170 (N_5170,N_4931,N_4946);
xor U5171 (N_5171,N_4944,N_4955);
and U5172 (N_5172,N_4979,N_4952);
or U5173 (N_5173,N_4855,N_4992);
nand U5174 (N_5174,N_4905,N_4841);
xor U5175 (N_5175,N_4996,N_4967);
xnor U5176 (N_5176,N_4863,N_4870);
and U5177 (N_5177,N_4877,N_4841);
xnor U5178 (N_5178,N_4895,N_4980);
nor U5179 (N_5179,N_4890,N_4872);
or U5180 (N_5180,N_4978,N_4938);
nor U5181 (N_5181,N_4952,N_4803);
or U5182 (N_5182,N_4915,N_4863);
xor U5183 (N_5183,N_4941,N_4821);
and U5184 (N_5184,N_4876,N_4900);
or U5185 (N_5185,N_4874,N_4869);
and U5186 (N_5186,N_4870,N_4902);
nand U5187 (N_5187,N_4888,N_4997);
or U5188 (N_5188,N_4989,N_4973);
nor U5189 (N_5189,N_4991,N_4917);
nor U5190 (N_5190,N_4998,N_4982);
nor U5191 (N_5191,N_4977,N_4866);
or U5192 (N_5192,N_4968,N_4841);
xnor U5193 (N_5193,N_4845,N_4867);
xor U5194 (N_5194,N_4861,N_4869);
nor U5195 (N_5195,N_4963,N_4961);
xnor U5196 (N_5196,N_4826,N_4837);
xor U5197 (N_5197,N_4943,N_4870);
or U5198 (N_5198,N_4818,N_4901);
xnor U5199 (N_5199,N_4860,N_4913);
and U5200 (N_5200,N_5014,N_5093);
nand U5201 (N_5201,N_5095,N_5030);
nor U5202 (N_5202,N_5061,N_5059);
nor U5203 (N_5203,N_5158,N_5003);
or U5204 (N_5204,N_5146,N_5064);
xor U5205 (N_5205,N_5124,N_5173);
and U5206 (N_5206,N_5111,N_5006);
or U5207 (N_5207,N_5034,N_5120);
xor U5208 (N_5208,N_5119,N_5132);
or U5209 (N_5209,N_5052,N_5103);
and U5210 (N_5210,N_5101,N_5066);
xnor U5211 (N_5211,N_5191,N_5040);
xor U5212 (N_5212,N_5032,N_5089);
and U5213 (N_5213,N_5099,N_5174);
nand U5214 (N_5214,N_5039,N_5025);
or U5215 (N_5215,N_5046,N_5041);
or U5216 (N_5216,N_5126,N_5058);
or U5217 (N_5217,N_5017,N_5016);
or U5218 (N_5218,N_5086,N_5028);
nand U5219 (N_5219,N_5113,N_5198);
nor U5220 (N_5220,N_5148,N_5050);
and U5221 (N_5221,N_5183,N_5021);
nand U5222 (N_5222,N_5091,N_5133);
and U5223 (N_5223,N_5096,N_5194);
nor U5224 (N_5224,N_5171,N_5170);
xor U5225 (N_5225,N_5131,N_5189);
nor U5226 (N_5226,N_5060,N_5062);
and U5227 (N_5227,N_5184,N_5165);
nand U5228 (N_5228,N_5180,N_5082);
or U5229 (N_5229,N_5164,N_5038);
or U5230 (N_5230,N_5051,N_5011);
and U5231 (N_5231,N_5172,N_5186);
nor U5232 (N_5232,N_5122,N_5185);
or U5233 (N_5233,N_5110,N_5007);
xor U5234 (N_5234,N_5027,N_5013);
nor U5235 (N_5235,N_5199,N_5105);
or U5236 (N_5236,N_5100,N_5085);
xnor U5237 (N_5237,N_5197,N_5090);
nand U5238 (N_5238,N_5143,N_5104);
and U5239 (N_5239,N_5080,N_5115);
nor U5240 (N_5240,N_5192,N_5123);
and U5241 (N_5241,N_5175,N_5002);
nand U5242 (N_5242,N_5035,N_5010);
nor U5243 (N_5243,N_5151,N_5130);
xor U5244 (N_5244,N_5162,N_5138);
or U5245 (N_5245,N_5083,N_5142);
nand U5246 (N_5246,N_5020,N_5154);
nor U5247 (N_5247,N_5106,N_5125);
xnor U5248 (N_5248,N_5055,N_5094);
nand U5249 (N_5249,N_5166,N_5156);
nand U5250 (N_5250,N_5152,N_5134);
and U5251 (N_5251,N_5144,N_5077);
nor U5252 (N_5252,N_5056,N_5098);
and U5253 (N_5253,N_5141,N_5190);
nand U5254 (N_5254,N_5179,N_5063);
or U5255 (N_5255,N_5159,N_5157);
and U5256 (N_5256,N_5069,N_5187);
xor U5257 (N_5257,N_5147,N_5068);
nor U5258 (N_5258,N_5000,N_5121);
and U5259 (N_5259,N_5114,N_5137);
nor U5260 (N_5260,N_5107,N_5178);
nor U5261 (N_5261,N_5065,N_5042);
or U5262 (N_5262,N_5048,N_5181);
or U5263 (N_5263,N_5015,N_5070);
nor U5264 (N_5264,N_5153,N_5193);
nor U5265 (N_5265,N_5116,N_5117);
xor U5266 (N_5266,N_5005,N_5024);
nand U5267 (N_5267,N_5088,N_5112);
or U5268 (N_5268,N_5075,N_5169);
nor U5269 (N_5269,N_5195,N_5087);
nand U5270 (N_5270,N_5031,N_5053);
xnor U5271 (N_5271,N_5135,N_5071);
xor U5272 (N_5272,N_5150,N_5092);
and U5273 (N_5273,N_5196,N_5047);
nor U5274 (N_5274,N_5177,N_5129);
or U5275 (N_5275,N_5074,N_5081);
nor U5276 (N_5276,N_5168,N_5076);
xnor U5277 (N_5277,N_5097,N_5176);
or U5278 (N_5278,N_5012,N_5043);
and U5279 (N_5279,N_5026,N_5022);
or U5280 (N_5280,N_5118,N_5023);
and U5281 (N_5281,N_5054,N_5033);
xnor U5282 (N_5282,N_5160,N_5009);
or U5283 (N_5283,N_5102,N_5149);
nor U5284 (N_5284,N_5004,N_5188);
xnor U5285 (N_5285,N_5161,N_5001);
nand U5286 (N_5286,N_5163,N_5084);
or U5287 (N_5287,N_5018,N_5139);
xnor U5288 (N_5288,N_5072,N_5079);
xor U5289 (N_5289,N_5128,N_5127);
nor U5290 (N_5290,N_5029,N_5108);
or U5291 (N_5291,N_5167,N_5057);
and U5292 (N_5292,N_5036,N_5019);
nor U5293 (N_5293,N_5008,N_5044);
nor U5294 (N_5294,N_5049,N_5145);
or U5295 (N_5295,N_5037,N_5155);
and U5296 (N_5296,N_5136,N_5045);
or U5297 (N_5297,N_5078,N_5109);
nand U5298 (N_5298,N_5073,N_5067);
nand U5299 (N_5299,N_5182,N_5140);
and U5300 (N_5300,N_5142,N_5096);
xor U5301 (N_5301,N_5062,N_5159);
or U5302 (N_5302,N_5102,N_5116);
and U5303 (N_5303,N_5108,N_5110);
xor U5304 (N_5304,N_5160,N_5193);
and U5305 (N_5305,N_5114,N_5125);
nor U5306 (N_5306,N_5179,N_5153);
or U5307 (N_5307,N_5146,N_5124);
nor U5308 (N_5308,N_5081,N_5011);
xnor U5309 (N_5309,N_5172,N_5042);
or U5310 (N_5310,N_5112,N_5018);
nor U5311 (N_5311,N_5005,N_5029);
nand U5312 (N_5312,N_5131,N_5162);
and U5313 (N_5313,N_5040,N_5106);
nor U5314 (N_5314,N_5054,N_5047);
nand U5315 (N_5315,N_5065,N_5002);
nor U5316 (N_5316,N_5036,N_5082);
and U5317 (N_5317,N_5087,N_5160);
or U5318 (N_5318,N_5146,N_5030);
nor U5319 (N_5319,N_5030,N_5101);
nor U5320 (N_5320,N_5134,N_5094);
xnor U5321 (N_5321,N_5033,N_5178);
and U5322 (N_5322,N_5004,N_5052);
and U5323 (N_5323,N_5070,N_5088);
nor U5324 (N_5324,N_5193,N_5152);
or U5325 (N_5325,N_5155,N_5190);
or U5326 (N_5326,N_5164,N_5167);
or U5327 (N_5327,N_5122,N_5147);
nor U5328 (N_5328,N_5032,N_5148);
and U5329 (N_5329,N_5070,N_5101);
nand U5330 (N_5330,N_5133,N_5054);
nor U5331 (N_5331,N_5009,N_5197);
nor U5332 (N_5332,N_5087,N_5003);
nand U5333 (N_5333,N_5089,N_5116);
or U5334 (N_5334,N_5022,N_5113);
xnor U5335 (N_5335,N_5165,N_5164);
or U5336 (N_5336,N_5071,N_5063);
and U5337 (N_5337,N_5078,N_5050);
xor U5338 (N_5338,N_5012,N_5161);
nand U5339 (N_5339,N_5058,N_5031);
xnor U5340 (N_5340,N_5120,N_5197);
and U5341 (N_5341,N_5159,N_5105);
nand U5342 (N_5342,N_5086,N_5163);
and U5343 (N_5343,N_5057,N_5107);
or U5344 (N_5344,N_5128,N_5065);
xor U5345 (N_5345,N_5081,N_5035);
nand U5346 (N_5346,N_5026,N_5111);
nand U5347 (N_5347,N_5161,N_5089);
nand U5348 (N_5348,N_5179,N_5177);
nor U5349 (N_5349,N_5031,N_5161);
and U5350 (N_5350,N_5033,N_5053);
nand U5351 (N_5351,N_5014,N_5049);
nand U5352 (N_5352,N_5020,N_5115);
or U5353 (N_5353,N_5158,N_5196);
nor U5354 (N_5354,N_5018,N_5020);
or U5355 (N_5355,N_5021,N_5160);
and U5356 (N_5356,N_5046,N_5177);
nor U5357 (N_5357,N_5078,N_5018);
and U5358 (N_5358,N_5041,N_5114);
or U5359 (N_5359,N_5145,N_5066);
nand U5360 (N_5360,N_5102,N_5070);
and U5361 (N_5361,N_5088,N_5173);
or U5362 (N_5362,N_5008,N_5002);
and U5363 (N_5363,N_5050,N_5068);
and U5364 (N_5364,N_5058,N_5077);
or U5365 (N_5365,N_5077,N_5002);
xor U5366 (N_5366,N_5036,N_5163);
nand U5367 (N_5367,N_5102,N_5092);
or U5368 (N_5368,N_5012,N_5136);
nor U5369 (N_5369,N_5125,N_5008);
and U5370 (N_5370,N_5156,N_5128);
or U5371 (N_5371,N_5036,N_5094);
xnor U5372 (N_5372,N_5051,N_5016);
and U5373 (N_5373,N_5080,N_5169);
or U5374 (N_5374,N_5045,N_5053);
nand U5375 (N_5375,N_5119,N_5033);
or U5376 (N_5376,N_5006,N_5132);
nor U5377 (N_5377,N_5082,N_5153);
nor U5378 (N_5378,N_5041,N_5076);
nor U5379 (N_5379,N_5099,N_5121);
nor U5380 (N_5380,N_5123,N_5095);
xnor U5381 (N_5381,N_5109,N_5000);
nand U5382 (N_5382,N_5151,N_5036);
nor U5383 (N_5383,N_5154,N_5184);
and U5384 (N_5384,N_5143,N_5033);
nand U5385 (N_5385,N_5021,N_5015);
xnor U5386 (N_5386,N_5185,N_5198);
and U5387 (N_5387,N_5190,N_5031);
nor U5388 (N_5388,N_5118,N_5133);
xnor U5389 (N_5389,N_5029,N_5196);
nand U5390 (N_5390,N_5087,N_5140);
nor U5391 (N_5391,N_5107,N_5129);
nand U5392 (N_5392,N_5009,N_5191);
and U5393 (N_5393,N_5016,N_5166);
nor U5394 (N_5394,N_5126,N_5060);
nand U5395 (N_5395,N_5138,N_5093);
or U5396 (N_5396,N_5193,N_5106);
xnor U5397 (N_5397,N_5036,N_5103);
xor U5398 (N_5398,N_5017,N_5161);
nand U5399 (N_5399,N_5052,N_5044);
xor U5400 (N_5400,N_5378,N_5202);
nand U5401 (N_5401,N_5311,N_5365);
xor U5402 (N_5402,N_5310,N_5295);
xor U5403 (N_5403,N_5376,N_5286);
and U5404 (N_5404,N_5366,N_5335);
nand U5405 (N_5405,N_5301,N_5364);
or U5406 (N_5406,N_5354,N_5352);
nor U5407 (N_5407,N_5343,N_5231);
and U5408 (N_5408,N_5339,N_5261);
or U5409 (N_5409,N_5347,N_5203);
or U5410 (N_5410,N_5332,N_5341);
nor U5411 (N_5411,N_5383,N_5307);
nor U5412 (N_5412,N_5234,N_5221);
or U5413 (N_5413,N_5395,N_5204);
nor U5414 (N_5414,N_5269,N_5390);
and U5415 (N_5415,N_5326,N_5399);
nor U5416 (N_5416,N_5283,N_5226);
or U5417 (N_5417,N_5353,N_5329);
xnor U5418 (N_5418,N_5370,N_5220);
or U5419 (N_5419,N_5244,N_5218);
nor U5420 (N_5420,N_5211,N_5206);
xor U5421 (N_5421,N_5267,N_5287);
or U5422 (N_5422,N_5299,N_5268);
and U5423 (N_5423,N_5227,N_5340);
and U5424 (N_5424,N_5358,N_5213);
nand U5425 (N_5425,N_5371,N_5263);
or U5426 (N_5426,N_5298,N_5276);
xnor U5427 (N_5427,N_5316,N_5271);
xnor U5428 (N_5428,N_5259,N_5273);
or U5429 (N_5429,N_5387,N_5249);
and U5430 (N_5430,N_5323,N_5243);
or U5431 (N_5431,N_5264,N_5318);
or U5432 (N_5432,N_5388,N_5367);
nor U5433 (N_5433,N_5360,N_5246);
xnor U5434 (N_5434,N_5214,N_5230);
nand U5435 (N_5435,N_5377,N_5241);
xor U5436 (N_5436,N_5331,N_5205);
nand U5437 (N_5437,N_5348,N_5351);
nor U5438 (N_5438,N_5284,N_5215);
nor U5439 (N_5439,N_5277,N_5285);
nor U5440 (N_5440,N_5305,N_5201);
or U5441 (N_5441,N_5274,N_5229);
xnor U5442 (N_5442,N_5328,N_5278);
xnor U5443 (N_5443,N_5294,N_5210);
or U5444 (N_5444,N_5398,N_5223);
and U5445 (N_5445,N_5315,N_5336);
nand U5446 (N_5446,N_5345,N_5260);
nand U5447 (N_5447,N_5280,N_5355);
and U5448 (N_5448,N_5225,N_5281);
or U5449 (N_5449,N_5372,N_5303);
nor U5450 (N_5450,N_5302,N_5306);
and U5451 (N_5451,N_5275,N_5250);
nor U5452 (N_5452,N_5209,N_5382);
xor U5453 (N_5453,N_5253,N_5312);
nor U5454 (N_5454,N_5346,N_5368);
and U5455 (N_5455,N_5247,N_5232);
and U5456 (N_5456,N_5394,N_5289);
nor U5457 (N_5457,N_5252,N_5397);
xor U5458 (N_5458,N_5321,N_5389);
nand U5459 (N_5459,N_5380,N_5219);
nand U5460 (N_5460,N_5379,N_5291);
or U5461 (N_5461,N_5308,N_5359);
and U5462 (N_5462,N_5304,N_5393);
and U5463 (N_5463,N_5237,N_5208);
and U5464 (N_5464,N_5207,N_5338);
or U5465 (N_5465,N_5248,N_5314);
nor U5466 (N_5466,N_5242,N_5319);
nor U5467 (N_5467,N_5236,N_5235);
or U5468 (N_5468,N_5320,N_5245);
or U5469 (N_5469,N_5391,N_5369);
or U5470 (N_5470,N_5309,N_5279);
and U5471 (N_5471,N_5349,N_5333);
or U5472 (N_5472,N_5266,N_5292);
or U5473 (N_5473,N_5216,N_5255);
nand U5474 (N_5474,N_5384,N_5363);
or U5475 (N_5475,N_5344,N_5375);
nor U5476 (N_5476,N_5381,N_5386);
xnor U5477 (N_5477,N_5288,N_5240);
nand U5478 (N_5478,N_5293,N_5313);
and U5479 (N_5479,N_5300,N_5222);
xnor U5480 (N_5480,N_5337,N_5282);
nand U5481 (N_5481,N_5373,N_5330);
or U5482 (N_5482,N_5356,N_5385);
nand U5483 (N_5483,N_5256,N_5396);
and U5484 (N_5484,N_5257,N_5224);
nand U5485 (N_5485,N_5357,N_5392);
nand U5486 (N_5486,N_5317,N_5350);
nor U5487 (N_5487,N_5296,N_5334);
nor U5488 (N_5488,N_5239,N_5265);
nor U5489 (N_5489,N_5322,N_5290);
nor U5490 (N_5490,N_5217,N_5362);
and U5491 (N_5491,N_5327,N_5325);
xnor U5492 (N_5492,N_5200,N_5251);
nand U5493 (N_5493,N_5258,N_5238);
and U5494 (N_5494,N_5297,N_5212);
and U5495 (N_5495,N_5342,N_5228);
nor U5496 (N_5496,N_5233,N_5272);
and U5497 (N_5497,N_5324,N_5361);
and U5498 (N_5498,N_5254,N_5374);
or U5499 (N_5499,N_5270,N_5262);
and U5500 (N_5500,N_5363,N_5336);
nor U5501 (N_5501,N_5380,N_5342);
or U5502 (N_5502,N_5263,N_5231);
or U5503 (N_5503,N_5378,N_5356);
or U5504 (N_5504,N_5332,N_5372);
nor U5505 (N_5505,N_5388,N_5371);
and U5506 (N_5506,N_5251,N_5383);
and U5507 (N_5507,N_5249,N_5238);
nand U5508 (N_5508,N_5330,N_5282);
or U5509 (N_5509,N_5291,N_5373);
nor U5510 (N_5510,N_5258,N_5216);
nand U5511 (N_5511,N_5399,N_5383);
nand U5512 (N_5512,N_5393,N_5253);
and U5513 (N_5513,N_5377,N_5334);
nand U5514 (N_5514,N_5245,N_5344);
nor U5515 (N_5515,N_5394,N_5256);
and U5516 (N_5516,N_5357,N_5204);
nor U5517 (N_5517,N_5258,N_5250);
and U5518 (N_5518,N_5365,N_5201);
and U5519 (N_5519,N_5328,N_5324);
nand U5520 (N_5520,N_5273,N_5276);
nand U5521 (N_5521,N_5292,N_5302);
nand U5522 (N_5522,N_5330,N_5331);
nand U5523 (N_5523,N_5220,N_5253);
nand U5524 (N_5524,N_5309,N_5371);
nand U5525 (N_5525,N_5270,N_5342);
nor U5526 (N_5526,N_5286,N_5363);
nand U5527 (N_5527,N_5361,N_5282);
and U5528 (N_5528,N_5236,N_5202);
or U5529 (N_5529,N_5262,N_5211);
nand U5530 (N_5530,N_5225,N_5270);
xnor U5531 (N_5531,N_5353,N_5324);
and U5532 (N_5532,N_5394,N_5249);
nor U5533 (N_5533,N_5277,N_5334);
xnor U5534 (N_5534,N_5324,N_5359);
and U5535 (N_5535,N_5280,N_5360);
or U5536 (N_5536,N_5253,N_5309);
nor U5537 (N_5537,N_5334,N_5275);
xnor U5538 (N_5538,N_5262,N_5251);
nor U5539 (N_5539,N_5217,N_5344);
or U5540 (N_5540,N_5254,N_5290);
nand U5541 (N_5541,N_5213,N_5322);
or U5542 (N_5542,N_5352,N_5362);
nor U5543 (N_5543,N_5334,N_5213);
and U5544 (N_5544,N_5346,N_5373);
or U5545 (N_5545,N_5345,N_5237);
and U5546 (N_5546,N_5211,N_5316);
nand U5547 (N_5547,N_5262,N_5280);
xor U5548 (N_5548,N_5347,N_5362);
and U5549 (N_5549,N_5280,N_5358);
nor U5550 (N_5550,N_5345,N_5236);
nor U5551 (N_5551,N_5289,N_5340);
or U5552 (N_5552,N_5348,N_5225);
xnor U5553 (N_5553,N_5266,N_5229);
and U5554 (N_5554,N_5372,N_5358);
nor U5555 (N_5555,N_5301,N_5370);
xor U5556 (N_5556,N_5205,N_5359);
nor U5557 (N_5557,N_5348,N_5316);
and U5558 (N_5558,N_5209,N_5271);
nor U5559 (N_5559,N_5218,N_5307);
or U5560 (N_5560,N_5260,N_5275);
xnor U5561 (N_5561,N_5316,N_5309);
or U5562 (N_5562,N_5324,N_5265);
and U5563 (N_5563,N_5305,N_5267);
and U5564 (N_5564,N_5206,N_5281);
nor U5565 (N_5565,N_5348,N_5312);
or U5566 (N_5566,N_5275,N_5304);
nor U5567 (N_5567,N_5333,N_5207);
and U5568 (N_5568,N_5245,N_5340);
xnor U5569 (N_5569,N_5339,N_5380);
and U5570 (N_5570,N_5222,N_5340);
or U5571 (N_5571,N_5267,N_5227);
nor U5572 (N_5572,N_5369,N_5298);
or U5573 (N_5573,N_5284,N_5232);
nand U5574 (N_5574,N_5351,N_5297);
and U5575 (N_5575,N_5375,N_5255);
xnor U5576 (N_5576,N_5285,N_5321);
and U5577 (N_5577,N_5344,N_5349);
xnor U5578 (N_5578,N_5308,N_5314);
xor U5579 (N_5579,N_5361,N_5275);
nor U5580 (N_5580,N_5321,N_5221);
xor U5581 (N_5581,N_5316,N_5270);
nor U5582 (N_5582,N_5334,N_5241);
or U5583 (N_5583,N_5218,N_5321);
and U5584 (N_5584,N_5342,N_5361);
nand U5585 (N_5585,N_5291,N_5363);
nand U5586 (N_5586,N_5326,N_5372);
xnor U5587 (N_5587,N_5374,N_5337);
nor U5588 (N_5588,N_5317,N_5306);
and U5589 (N_5589,N_5279,N_5397);
xor U5590 (N_5590,N_5389,N_5381);
xor U5591 (N_5591,N_5395,N_5351);
xnor U5592 (N_5592,N_5370,N_5346);
or U5593 (N_5593,N_5326,N_5302);
nor U5594 (N_5594,N_5299,N_5308);
xor U5595 (N_5595,N_5244,N_5209);
and U5596 (N_5596,N_5229,N_5321);
and U5597 (N_5597,N_5320,N_5242);
and U5598 (N_5598,N_5275,N_5378);
and U5599 (N_5599,N_5217,N_5297);
xor U5600 (N_5600,N_5560,N_5510);
nand U5601 (N_5601,N_5473,N_5407);
and U5602 (N_5602,N_5515,N_5493);
nor U5603 (N_5603,N_5518,N_5503);
and U5604 (N_5604,N_5438,N_5543);
and U5605 (N_5605,N_5440,N_5486);
nand U5606 (N_5606,N_5405,N_5457);
nor U5607 (N_5607,N_5437,N_5491);
or U5608 (N_5608,N_5451,N_5542);
xnor U5609 (N_5609,N_5428,N_5441);
nor U5610 (N_5610,N_5481,N_5466);
nor U5611 (N_5611,N_5580,N_5410);
and U5612 (N_5612,N_5596,N_5423);
and U5613 (N_5613,N_5482,N_5448);
nor U5614 (N_5614,N_5462,N_5562);
or U5615 (N_5615,N_5402,N_5586);
xor U5616 (N_5616,N_5498,N_5544);
or U5617 (N_5617,N_5570,N_5413);
nand U5618 (N_5618,N_5599,N_5558);
nand U5619 (N_5619,N_5431,N_5537);
xor U5620 (N_5620,N_5576,N_5519);
or U5621 (N_5621,N_5589,N_5533);
nor U5622 (N_5622,N_5495,N_5546);
and U5623 (N_5623,N_5531,N_5517);
or U5624 (N_5624,N_5587,N_5508);
nand U5625 (N_5625,N_5568,N_5447);
xor U5626 (N_5626,N_5427,N_5574);
or U5627 (N_5627,N_5496,N_5461);
or U5628 (N_5628,N_5528,N_5480);
xor U5629 (N_5629,N_5585,N_5455);
and U5630 (N_5630,N_5475,N_5442);
and U5631 (N_5631,N_5549,N_5488);
nand U5632 (N_5632,N_5532,N_5535);
or U5633 (N_5633,N_5408,N_5563);
or U5634 (N_5634,N_5581,N_5584);
and U5635 (N_5635,N_5567,N_5575);
nor U5636 (N_5636,N_5534,N_5504);
nor U5637 (N_5637,N_5404,N_5520);
xnor U5638 (N_5638,N_5500,N_5446);
nand U5639 (N_5639,N_5460,N_5470);
and U5640 (N_5640,N_5434,N_5595);
xor U5641 (N_5641,N_5468,N_5529);
nor U5642 (N_5642,N_5497,N_5458);
xnor U5643 (N_5643,N_5536,N_5483);
or U5644 (N_5644,N_5416,N_5444);
nand U5645 (N_5645,N_5527,N_5573);
or U5646 (N_5646,N_5465,N_5569);
and U5647 (N_5647,N_5530,N_5545);
xor U5648 (N_5648,N_5400,N_5538);
nand U5649 (N_5649,N_5594,N_5523);
and U5650 (N_5650,N_5422,N_5474);
or U5651 (N_5651,N_5578,N_5555);
xor U5652 (N_5652,N_5456,N_5565);
xnor U5653 (N_5653,N_5540,N_5501);
and U5654 (N_5654,N_5541,N_5472);
nor U5655 (N_5655,N_5450,N_5430);
nor U5656 (N_5656,N_5424,N_5453);
xnor U5657 (N_5657,N_5494,N_5526);
and U5658 (N_5658,N_5484,N_5499);
xnor U5659 (N_5659,N_5443,N_5445);
or U5660 (N_5660,N_5554,N_5598);
nand U5661 (N_5661,N_5582,N_5566);
and U5662 (N_5662,N_5487,N_5583);
xor U5663 (N_5663,N_5525,N_5425);
nor U5664 (N_5664,N_5561,N_5509);
nor U5665 (N_5665,N_5521,N_5469);
nor U5666 (N_5666,N_5556,N_5577);
xor U5667 (N_5667,N_5511,N_5421);
and U5668 (N_5668,N_5571,N_5432);
nor U5669 (N_5669,N_5479,N_5507);
xor U5670 (N_5670,N_5471,N_5435);
nor U5671 (N_5671,N_5512,N_5513);
nor U5672 (N_5672,N_5489,N_5579);
xor U5673 (N_5673,N_5492,N_5426);
nor U5674 (N_5674,N_5552,N_5464);
nand U5675 (N_5675,N_5415,N_5477);
nor U5676 (N_5676,N_5502,N_5505);
and U5677 (N_5677,N_5406,N_5522);
and U5678 (N_5678,N_5597,N_5412);
and U5679 (N_5679,N_5524,N_5417);
or U5680 (N_5680,N_5449,N_5551);
or U5681 (N_5681,N_5452,N_5419);
and U5682 (N_5682,N_5553,N_5514);
or U5683 (N_5683,N_5559,N_5459);
nor U5684 (N_5684,N_5564,N_5409);
and U5685 (N_5685,N_5433,N_5485);
nand U5686 (N_5686,N_5429,N_5516);
or U5687 (N_5687,N_5490,N_5548);
or U5688 (N_5688,N_5550,N_5590);
xnor U5689 (N_5689,N_5403,N_5420);
xnor U5690 (N_5690,N_5463,N_5467);
and U5691 (N_5691,N_5478,N_5439);
or U5692 (N_5692,N_5557,N_5414);
nor U5693 (N_5693,N_5591,N_5401);
nand U5694 (N_5694,N_5454,N_5506);
xnor U5695 (N_5695,N_5411,N_5593);
and U5696 (N_5696,N_5539,N_5547);
xor U5697 (N_5697,N_5418,N_5588);
or U5698 (N_5698,N_5572,N_5436);
nor U5699 (N_5699,N_5476,N_5592);
or U5700 (N_5700,N_5419,N_5496);
or U5701 (N_5701,N_5427,N_5591);
nand U5702 (N_5702,N_5591,N_5459);
or U5703 (N_5703,N_5508,N_5455);
and U5704 (N_5704,N_5467,N_5414);
and U5705 (N_5705,N_5426,N_5441);
or U5706 (N_5706,N_5478,N_5512);
or U5707 (N_5707,N_5489,N_5596);
nor U5708 (N_5708,N_5510,N_5471);
nor U5709 (N_5709,N_5547,N_5559);
nor U5710 (N_5710,N_5538,N_5543);
and U5711 (N_5711,N_5443,N_5534);
nand U5712 (N_5712,N_5490,N_5594);
nor U5713 (N_5713,N_5576,N_5425);
nand U5714 (N_5714,N_5548,N_5542);
nand U5715 (N_5715,N_5414,N_5453);
and U5716 (N_5716,N_5425,N_5501);
xor U5717 (N_5717,N_5422,N_5574);
nand U5718 (N_5718,N_5597,N_5567);
or U5719 (N_5719,N_5521,N_5457);
nor U5720 (N_5720,N_5549,N_5554);
nand U5721 (N_5721,N_5554,N_5497);
or U5722 (N_5722,N_5434,N_5427);
xnor U5723 (N_5723,N_5516,N_5446);
nand U5724 (N_5724,N_5598,N_5520);
or U5725 (N_5725,N_5512,N_5505);
and U5726 (N_5726,N_5431,N_5533);
or U5727 (N_5727,N_5430,N_5556);
xnor U5728 (N_5728,N_5599,N_5539);
nor U5729 (N_5729,N_5499,N_5589);
and U5730 (N_5730,N_5568,N_5478);
nor U5731 (N_5731,N_5403,N_5557);
and U5732 (N_5732,N_5479,N_5445);
nand U5733 (N_5733,N_5514,N_5536);
xor U5734 (N_5734,N_5466,N_5534);
xnor U5735 (N_5735,N_5462,N_5571);
or U5736 (N_5736,N_5471,N_5532);
or U5737 (N_5737,N_5528,N_5491);
xor U5738 (N_5738,N_5496,N_5475);
nor U5739 (N_5739,N_5452,N_5515);
xor U5740 (N_5740,N_5506,N_5437);
or U5741 (N_5741,N_5550,N_5459);
nor U5742 (N_5742,N_5400,N_5541);
nor U5743 (N_5743,N_5455,N_5526);
nor U5744 (N_5744,N_5499,N_5447);
xor U5745 (N_5745,N_5419,N_5501);
and U5746 (N_5746,N_5559,N_5585);
nand U5747 (N_5747,N_5478,N_5593);
and U5748 (N_5748,N_5532,N_5545);
and U5749 (N_5749,N_5542,N_5558);
xor U5750 (N_5750,N_5514,N_5492);
or U5751 (N_5751,N_5554,N_5531);
nand U5752 (N_5752,N_5586,N_5418);
nand U5753 (N_5753,N_5576,N_5478);
xnor U5754 (N_5754,N_5593,N_5449);
or U5755 (N_5755,N_5513,N_5428);
nor U5756 (N_5756,N_5435,N_5550);
or U5757 (N_5757,N_5521,N_5594);
nand U5758 (N_5758,N_5531,N_5494);
and U5759 (N_5759,N_5445,N_5414);
or U5760 (N_5760,N_5475,N_5407);
and U5761 (N_5761,N_5570,N_5523);
and U5762 (N_5762,N_5432,N_5417);
or U5763 (N_5763,N_5493,N_5421);
nor U5764 (N_5764,N_5478,N_5557);
or U5765 (N_5765,N_5571,N_5450);
nor U5766 (N_5766,N_5518,N_5523);
nand U5767 (N_5767,N_5439,N_5503);
nand U5768 (N_5768,N_5566,N_5508);
nor U5769 (N_5769,N_5587,N_5547);
xnor U5770 (N_5770,N_5439,N_5583);
nand U5771 (N_5771,N_5557,N_5408);
or U5772 (N_5772,N_5406,N_5453);
nor U5773 (N_5773,N_5557,N_5428);
xor U5774 (N_5774,N_5434,N_5536);
or U5775 (N_5775,N_5559,N_5412);
or U5776 (N_5776,N_5536,N_5521);
xor U5777 (N_5777,N_5416,N_5432);
nor U5778 (N_5778,N_5505,N_5448);
or U5779 (N_5779,N_5405,N_5430);
nand U5780 (N_5780,N_5570,N_5507);
nor U5781 (N_5781,N_5404,N_5400);
xnor U5782 (N_5782,N_5558,N_5512);
or U5783 (N_5783,N_5531,N_5461);
nand U5784 (N_5784,N_5525,N_5592);
and U5785 (N_5785,N_5489,N_5404);
or U5786 (N_5786,N_5536,N_5437);
or U5787 (N_5787,N_5494,N_5453);
nand U5788 (N_5788,N_5435,N_5517);
and U5789 (N_5789,N_5564,N_5407);
xnor U5790 (N_5790,N_5527,N_5412);
nor U5791 (N_5791,N_5567,N_5588);
xnor U5792 (N_5792,N_5455,N_5555);
nand U5793 (N_5793,N_5513,N_5530);
nand U5794 (N_5794,N_5507,N_5431);
xor U5795 (N_5795,N_5482,N_5420);
xor U5796 (N_5796,N_5418,N_5446);
and U5797 (N_5797,N_5472,N_5426);
and U5798 (N_5798,N_5451,N_5593);
or U5799 (N_5799,N_5432,N_5514);
and U5800 (N_5800,N_5751,N_5602);
or U5801 (N_5801,N_5639,N_5611);
nor U5802 (N_5802,N_5755,N_5708);
and U5803 (N_5803,N_5651,N_5649);
nand U5804 (N_5804,N_5785,N_5773);
nand U5805 (N_5805,N_5682,N_5605);
nand U5806 (N_5806,N_5713,N_5673);
or U5807 (N_5807,N_5608,N_5614);
xor U5808 (N_5808,N_5739,N_5712);
and U5809 (N_5809,N_5670,N_5694);
and U5810 (N_5810,N_5724,N_5618);
and U5811 (N_5811,N_5658,N_5625);
nand U5812 (N_5812,N_5722,N_5632);
or U5813 (N_5813,N_5696,N_5648);
or U5814 (N_5814,N_5681,N_5669);
xnor U5815 (N_5815,N_5684,N_5686);
and U5816 (N_5816,N_5750,N_5638);
xnor U5817 (N_5817,N_5645,N_5788);
and U5818 (N_5818,N_5716,N_5742);
and U5819 (N_5819,N_5757,N_5704);
xnor U5820 (N_5820,N_5607,N_5626);
nor U5821 (N_5821,N_5616,N_5775);
nand U5822 (N_5822,N_5679,N_5737);
nand U5823 (N_5823,N_5705,N_5703);
and U5824 (N_5824,N_5759,N_5663);
or U5825 (N_5825,N_5765,N_5784);
xnor U5826 (N_5826,N_5695,N_5767);
or U5827 (N_5827,N_5671,N_5760);
or U5828 (N_5828,N_5702,N_5701);
or U5829 (N_5829,N_5640,N_5735);
xor U5830 (N_5830,N_5680,N_5762);
or U5831 (N_5831,N_5698,N_5706);
nor U5832 (N_5832,N_5672,N_5627);
or U5833 (N_5833,N_5661,N_5783);
and U5834 (N_5834,N_5769,N_5726);
xor U5835 (N_5835,N_5718,N_5675);
nor U5836 (N_5836,N_5655,N_5752);
xnor U5837 (N_5837,N_5652,N_5609);
or U5838 (N_5838,N_5644,N_5728);
nand U5839 (N_5839,N_5710,N_5600);
xnor U5840 (N_5840,N_5711,N_5794);
or U5841 (N_5841,N_5657,N_5761);
nand U5842 (N_5842,N_5787,N_5641);
or U5843 (N_5843,N_5779,N_5789);
nor U5844 (N_5844,N_5612,N_5615);
and U5845 (N_5845,N_5601,N_5631);
and U5846 (N_5846,N_5633,N_5778);
and U5847 (N_5847,N_5690,N_5668);
or U5848 (N_5848,N_5731,N_5709);
or U5849 (N_5849,N_5624,N_5717);
and U5850 (N_5850,N_5629,N_5674);
xnor U5851 (N_5851,N_5666,N_5730);
and U5852 (N_5852,N_5781,N_5768);
or U5853 (N_5853,N_5683,N_5746);
nand U5854 (N_5854,N_5797,N_5749);
or U5855 (N_5855,N_5720,N_5772);
xnor U5856 (N_5856,N_5656,N_5707);
nand U5857 (N_5857,N_5798,N_5620);
nand U5858 (N_5858,N_5741,N_5721);
nor U5859 (N_5859,N_5736,N_5604);
and U5860 (N_5860,N_5770,N_5771);
nand U5861 (N_5861,N_5685,N_5693);
nor U5862 (N_5862,N_5753,N_5660);
and U5863 (N_5863,N_5723,N_5740);
nor U5864 (N_5864,N_5756,N_5795);
and U5865 (N_5865,N_5744,N_5699);
nand U5866 (N_5866,N_5617,N_5630);
nand U5867 (N_5867,N_5745,N_5662);
nand U5868 (N_5868,N_5733,N_5636);
or U5869 (N_5869,N_5623,N_5621);
or U5870 (N_5870,N_5606,N_5790);
and U5871 (N_5871,N_5635,N_5764);
xor U5872 (N_5872,N_5793,N_5637);
xor U5873 (N_5873,N_5650,N_5715);
xor U5874 (N_5874,N_5763,N_5747);
and U5875 (N_5875,N_5697,N_5610);
and U5876 (N_5876,N_5729,N_5667);
or U5877 (N_5877,N_5748,N_5774);
xnor U5878 (N_5878,N_5603,N_5688);
xor U5879 (N_5879,N_5725,N_5678);
nand U5880 (N_5880,N_5734,N_5792);
nand U5881 (N_5881,N_5692,N_5714);
nand U5882 (N_5882,N_5727,N_5796);
nand U5883 (N_5883,N_5738,N_5776);
or U5884 (N_5884,N_5647,N_5689);
and U5885 (N_5885,N_5619,N_5613);
nor U5886 (N_5886,N_5622,N_5766);
xnor U5887 (N_5887,N_5719,N_5628);
or U5888 (N_5888,N_5642,N_5732);
or U5889 (N_5889,N_5687,N_5791);
or U5890 (N_5890,N_5646,N_5780);
nand U5891 (N_5891,N_5758,N_5665);
and U5892 (N_5892,N_5799,N_5659);
and U5893 (N_5893,N_5782,N_5786);
nor U5894 (N_5894,N_5777,N_5691);
xnor U5895 (N_5895,N_5654,N_5653);
and U5896 (N_5896,N_5664,N_5634);
nor U5897 (N_5897,N_5676,N_5643);
and U5898 (N_5898,N_5700,N_5743);
nand U5899 (N_5899,N_5754,N_5677);
nor U5900 (N_5900,N_5743,N_5689);
or U5901 (N_5901,N_5648,N_5619);
xnor U5902 (N_5902,N_5649,N_5776);
and U5903 (N_5903,N_5698,N_5732);
nand U5904 (N_5904,N_5762,N_5730);
and U5905 (N_5905,N_5674,N_5705);
and U5906 (N_5906,N_5776,N_5616);
nand U5907 (N_5907,N_5756,N_5713);
and U5908 (N_5908,N_5765,N_5720);
or U5909 (N_5909,N_5754,N_5786);
nand U5910 (N_5910,N_5602,N_5722);
nand U5911 (N_5911,N_5661,N_5755);
nor U5912 (N_5912,N_5704,N_5618);
xor U5913 (N_5913,N_5613,N_5649);
or U5914 (N_5914,N_5647,N_5620);
nor U5915 (N_5915,N_5647,N_5673);
and U5916 (N_5916,N_5794,N_5749);
xor U5917 (N_5917,N_5664,N_5605);
nand U5918 (N_5918,N_5661,N_5718);
xnor U5919 (N_5919,N_5797,N_5653);
nand U5920 (N_5920,N_5693,N_5648);
nor U5921 (N_5921,N_5683,N_5744);
nand U5922 (N_5922,N_5715,N_5654);
or U5923 (N_5923,N_5632,N_5739);
nor U5924 (N_5924,N_5690,N_5674);
and U5925 (N_5925,N_5668,N_5693);
xor U5926 (N_5926,N_5625,N_5603);
nor U5927 (N_5927,N_5641,N_5746);
and U5928 (N_5928,N_5615,N_5702);
nand U5929 (N_5929,N_5768,N_5767);
nor U5930 (N_5930,N_5714,N_5734);
or U5931 (N_5931,N_5778,N_5732);
or U5932 (N_5932,N_5769,N_5667);
and U5933 (N_5933,N_5673,N_5674);
or U5934 (N_5934,N_5683,N_5620);
or U5935 (N_5935,N_5674,N_5683);
or U5936 (N_5936,N_5677,N_5749);
xor U5937 (N_5937,N_5686,N_5732);
nand U5938 (N_5938,N_5688,N_5739);
and U5939 (N_5939,N_5713,N_5608);
nor U5940 (N_5940,N_5649,N_5791);
xnor U5941 (N_5941,N_5688,N_5613);
or U5942 (N_5942,N_5612,N_5737);
nand U5943 (N_5943,N_5799,N_5703);
nand U5944 (N_5944,N_5635,N_5723);
nand U5945 (N_5945,N_5639,N_5756);
nor U5946 (N_5946,N_5681,N_5680);
xnor U5947 (N_5947,N_5642,N_5753);
and U5948 (N_5948,N_5772,N_5731);
nand U5949 (N_5949,N_5787,N_5637);
xnor U5950 (N_5950,N_5636,N_5777);
nor U5951 (N_5951,N_5755,N_5689);
nand U5952 (N_5952,N_5670,N_5612);
and U5953 (N_5953,N_5727,N_5615);
nor U5954 (N_5954,N_5767,N_5798);
nand U5955 (N_5955,N_5622,N_5665);
or U5956 (N_5956,N_5626,N_5628);
nor U5957 (N_5957,N_5676,N_5636);
nor U5958 (N_5958,N_5633,N_5654);
nand U5959 (N_5959,N_5788,N_5701);
nor U5960 (N_5960,N_5685,N_5747);
xnor U5961 (N_5961,N_5733,N_5618);
or U5962 (N_5962,N_5667,N_5631);
and U5963 (N_5963,N_5779,N_5741);
or U5964 (N_5964,N_5794,N_5632);
xnor U5965 (N_5965,N_5733,N_5781);
nor U5966 (N_5966,N_5685,N_5655);
or U5967 (N_5967,N_5756,N_5679);
xor U5968 (N_5968,N_5635,N_5744);
nor U5969 (N_5969,N_5666,N_5684);
or U5970 (N_5970,N_5700,N_5731);
or U5971 (N_5971,N_5763,N_5618);
and U5972 (N_5972,N_5758,N_5638);
nand U5973 (N_5973,N_5644,N_5709);
nor U5974 (N_5974,N_5712,N_5781);
or U5975 (N_5975,N_5665,N_5712);
nand U5976 (N_5976,N_5683,N_5648);
nor U5977 (N_5977,N_5670,N_5642);
nand U5978 (N_5978,N_5660,N_5698);
nand U5979 (N_5979,N_5762,N_5783);
and U5980 (N_5980,N_5681,N_5738);
nand U5981 (N_5981,N_5696,N_5603);
nand U5982 (N_5982,N_5726,N_5655);
nor U5983 (N_5983,N_5709,N_5602);
xor U5984 (N_5984,N_5744,N_5743);
xor U5985 (N_5985,N_5600,N_5784);
and U5986 (N_5986,N_5763,N_5681);
nor U5987 (N_5987,N_5684,N_5631);
or U5988 (N_5988,N_5620,N_5637);
nand U5989 (N_5989,N_5615,N_5724);
or U5990 (N_5990,N_5692,N_5717);
nand U5991 (N_5991,N_5749,N_5640);
nor U5992 (N_5992,N_5779,N_5735);
xnor U5993 (N_5993,N_5750,N_5740);
nand U5994 (N_5994,N_5790,N_5693);
nand U5995 (N_5995,N_5752,N_5611);
or U5996 (N_5996,N_5698,N_5731);
nor U5997 (N_5997,N_5758,N_5607);
or U5998 (N_5998,N_5770,N_5676);
nor U5999 (N_5999,N_5667,N_5606);
or U6000 (N_6000,N_5801,N_5942);
nand U6001 (N_6001,N_5851,N_5911);
and U6002 (N_6002,N_5953,N_5803);
nor U6003 (N_6003,N_5881,N_5980);
and U6004 (N_6004,N_5805,N_5869);
or U6005 (N_6005,N_5894,N_5884);
nand U6006 (N_6006,N_5877,N_5843);
xor U6007 (N_6007,N_5943,N_5825);
nand U6008 (N_6008,N_5863,N_5833);
nor U6009 (N_6009,N_5928,N_5835);
nand U6010 (N_6010,N_5907,N_5978);
xor U6011 (N_6011,N_5821,N_5817);
or U6012 (N_6012,N_5872,N_5968);
nand U6013 (N_6013,N_5908,N_5929);
nand U6014 (N_6014,N_5822,N_5946);
xnor U6015 (N_6015,N_5889,N_5897);
or U6016 (N_6016,N_5847,N_5922);
xnor U6017 (N_6017,N_5974,N_5827);
xnor U6018 (N_6018,N_5807,N_5837);
xnor U6019 (N_6019,N_5850,N_5971);
and U6020 (N_6020,N_5853,N_5988);
and U6021 (N_6021,N_5886,N_5948);
nand U6022 (N_6022,N_5918,N_5826);
nor U6023 (N_6023,N_5998,N_5984);
or U6024 (N_6024,N_5997,N_5800);
or U6025 (N_6025,N_5986,N_5887);
or U6026 (N_6026,N_5861,N_5926);
nand U6027 (N_6027,N_5808,N_5999);
nand U6028 (N_6028,N_5823,N_5959);
nand U6029 (N_6029,N_5882,N_5979);
or U6030 (N_6030,N_5901,N_5873);
nor U6031 (N_6031,N_5956,N_5931);
and U6032 (N_6032,N_5944,N_5875);
nand U6033 (N_6033,N_5809,N_5913);
and U6034 (N_6034,N_5891,N_5836);
or U6035 (N_6035,N_5903,N_5914);
nand U6036 (N_6036,N_5860,N_5934);
nand U6037 (N_6037,N_5831,N_5976);
nand U6038 (N_6038,N_5975,N_5815);
or U6039 (N_6039,N_5846,N_5862);
or U6040 (N_6040,N_5938,N_5947);
xnor U6041 (N_6041,N_5924,N_5952);
nor U6042 (N_6042,N_5910,N_5965);
or U6043 (N_6043,N_5856,N_5842);
nand U6044 (N_6044,N_5993,N_5954);
and U6045 (N_6045,N_5937,N_5985);
and U6046 (N_6046,N_5950,N_5879);
nor U6047 (N_6047,N_5804,N_5994);
nand U6048 (N_6048,N_5973,N_5857);
nor U6049 (N_6049,N_5810,N_5900);
or U6050 (N_6050,N_5841,N_5878);
nor U6051 (N_6051,N_5870,N_5838);
nor U6052 (N_6052,N_5859,N_5936);
nor U6053 (N_6053,N_5819,N_5813);
or U6054 (N_6054,N_5923,N_5935);
nor U6055 (N_6055,N_5921,N_5949);
nor U6056 (N_6056,N_5987,N_5834);
or U6057 (N_6057,N_5962,N_5854);
nor U6058 (N_6058,N_5883,N_5874);
xnor U6059 (N_6059,N_5888,N_5902);
nor U6060 (N_6060,N_5876,N_5945);
nand U6061 (N_6061,N_5989,N_5905);
nor U6062 (N_6062,N_5868,N_5927);
xor U6063 (N_6063,N_5848,N_5829);
or U6064 (N_6064,N_5852,N_5940);
xnor U6065 (N_6065,N_5867,N_5820);
or U6066 (N_6066,N_5933,N_5816);
nor U6067 (N_6067,N_5812,N_5916);
and U6068 (N_6068,N_5951,N_5865);
nand U6069 (N_6069,N_5991,N_5866);
xor U6070 (N_6070,N_5871,N_5832);
xnor U6071 (N_6071,N_5920,N_5828);
nand U6072 (N_6072,N_5895,N_5972);
and U6073 (N_6073,N_5930,N_5830);
nor U6074 (N_6074,N_5939,N_5845);
nand U6075 (N_6075,N_5824,N_5983);
xor U6076 (N_6076,N_5840,N_5996);
nand U6077 (N_6077,N_5858,N_5802);
or U6078 (N_6078,N_5919,N_5969);
nor U6079 (N_6079,N_5982,N_5932);
xnor U6080 (N_6080,N_5915,N_5961);
nand U6081 (N_6081,N_5880,N_5909);
or U6082 (N_6082,N_5963,N_5818);
nor U6083 (N_6083,N_5912,N_5925);
and U6084 (N_6084,N_5849,N_5906);
and U6085 (N_6085,N_5995,N_5896);
and U6086 (N_6086,N_5864,N_5977);
nor U6087 (N_6087,N_5855,N_5904);
nand U6088 (N_6088,N_5899,N_5964);
or U6089 (N_6089,N_5992,N_5844);
or U6090 (N_6090,N_5892,N_5814);
or U6091 (N_6091,N_5957,N_5885);
or U6092 (N_6092,N_5811,N_5839);
or U6093 (N_6093,N_5960,N_5981);
nor U6094 (N_6094,N_5970,N_5893);
and U6095 (N_6095,N_5941,N_5958);
xor U6096 (N_6096,N_5917,N_5967);
xnor U6097 (N_6097,N_5898,N_5966);
nor U6098 (N_6098,N_5990,N_5890);
nor U6099 (N_6099,N_5806,N_5955);
nor U6100 (N_6100,N_5992,N_5800);
xor U6101 (N_6101,N_5950,N_5842);
nor U6102 (N_6102,N_5859,N_5939);
and U6103 (N_6103,N_5888,N_5972);
nor U6104 (N_6104,N_5805,N_5815);
xnor U6105 (N_6105,N_5966,N_5971);
and U6106 (N_6106,N_5985,N_5871);
nor U6107 (N_6107,N_5806,N_5962);
or U6108 (N_6108,N_5863,N_5901);
nand U6109 (N_6109,N_5879,N_5883);
or U6110 (N_6110,N_5842,N_5919);
nor U6111 (N_6111,N_5814,N_5869);
nor U6112 (N_6112,N_5978,N_5865);
and U6113 (N_6113,N_5858,N_5850);
or U6114 (N_6114,N_5994,N_5952);
and U6115 (N_6115,N_5965,N_5966);
and U6116 (N_6116,N_5946,N_5938);
or U6117 (N_6117,N_5951,N_5975);
nand U6118 (N_6118,N_5882,N_5823);
or U6119 (N_6119,N_5804,N_5858);
nand U6120 (N_6120,N_5971,N_5898);
xor U6121 (N_6121,N_5888,N_5808);
xnor U6122 (N_6122,N_5947,N_5830);
nand U6123 (N_6123,N_5805,N_5833);
xnor U6124 (N_6124,N_5885,N_5892);
nand U6125 (N_6125,N_5836,N_5958);
and U6126 (N_6126,N_5889,N_5904);
and U6127 (N_6127,N_5915,N_5840);
nand U6128 (N_6128,N_5901,N_5958);
or U6129 (N_6129,N_5937,N_5856);
nand U6130 (N_6130,N_5919,N_5998);
or U6131 (N_6131,N_5924,N_5848);
and U6132 (N_6132,N_5884,N_5991);
nand U6133 (N_6133,N_5875,N_5868);
nand U6134 (N_6134,N_5993,N_5947);
nor U6135 (N_6135,N_5839,N_5942);
xnor U6136 (N_6136,N_5849,N_5945);
nor U6137 (N_6137,N_5877,N_5845);
nand U6138 (N_6138,N_5929,N_5941);
and U6139 (N_6139,N_5892,N_5818);
xnor U6140 (N_6140,N_5932,N_5878);
xnor U6141 (N_6141,N_5968,N_5898);
or U6142 (N_6142,N_5879,N_5949);
and U6143 (N_6143,N_5808,N_5985);
and U6144 (N_6144,N_5873,N_5982);
nand U6145 (N_6145,N_5837,N_5833);
nor U6146 (N_6146,N_5946,N_5819);
nor U6147 (N_6147,N_5901,N_5858);
xnor U6148 (N_6148,N_5963,N_5898);
or U6149 (N_6149,N_5959,N_5994);
or U6150 (N_6150,N_5921,N_5903);
nor U6151 (N_6151,N_5958,N_5921);
or U6152 (N_6152,N_5917,N_5890);
or U6153 (N_6153,N_5811,N_5991);
nor U6154 (N_6154,N_5899,N_5986);
or U6155 (N_6155,N_5812,N_5987);
xor U6156 (N_6156,N_5952,N_5982);
nor U6157 (N_6157,N_5966,N_5964);
and U6158 (N_6158,N_5956,N_5891);
xnor U6159 (N_6159,N_5843,N_5973);
or U6160 (N_6160,N_5933,N_5930);
nand U6161 (N_6161,N_5905,N_5853);
or U6162 (N_6162,N_5874,N_5938);
and U6163 (N_6163,N_5981,N_5802);
nand U6164 (N_6164,N_5863,N_5945);
nor U6165 (N_6165,N_5997,N_5817);
or U6166 (N_6166,N_5912,N_5994);
or U6167 (N_6167,N_5827,N_5824);
xnor U6168 (N_6168,N_5917,N_5831);
and U6169 (N_6169,N_5831,N_5835);
nand U6170 (N_6170,N_5983,N_5919);
nor U6171 (N_6171,N_5927,N_5992);
xor U6172 (N_6172,N_5868,N_5924);
or U6173 (N_6173,N_5901,N_5903);
nand U6174 (N_6174,N_5859,N_5870);
xor U6175 (N_6175,N_5983,N_5857);
and U6176 (N_6176,N_5855,N_5841);
nor U6177 (N_6177,N_5912,N_5866);
and U6178 (N_6178,N_5985,N_5823);
nand U6179 (N_6179,N_5830,N_5978);
and U6180 (N_6180,N_5975,N_5916);
xor U6181 (N_6181,N_5956,N_5998);
nor U6182 (N_6182,N_5967,N_5912);
or U6183 (N_6183,N_5932,N_5968);
nand U6184 (N_6184,N_5904,N_5842);
nor U6185 (N_6185,N_5980,N_5855);
and U6186 (N_6186,N_5936,N_5966);
xnor U6187 (N_6187,N_5970,N_5870);
nand U6188 (N_6188,N_5971,N_5951);
or U6189 (N_6189,N_5924,N_5916);
xor U6190 (N_6190,N_5945,N_5913);
nor U6191 (N_6191,N_5846,N_5947);
xor U6192 (N_6192,N_5924,N_5802);
or U6193 (N_6193,N_5949,N_5937);
nand U6194 (N_6194,N_5880,N_5823);
xor U6195 (N_6195,N_5984,N_5840);
and U6196 (N_6196,N_5877,N_5923);
nand U6197 (N_6197,N_5925,N_5920);
nor U6198 (N_6198,N_5974,N_5925);
nand U6199 (N_6199,N_5858,N_5834);
xnor U6200 (N_6200,N_6048,N_6061);
and U6201 (N_6201,N_6001,N_6090);
nand U6202 (N_6202,N_6062,N_6144);
nand U6203 (N_6203,N_6009,N_6112);
or U6204 (N_6204,N_6071,N_6084);
nor U6205 (N_6205,N_6191,N_6136);
or U6206 (N_6206,N_6147,N_6010);
or U6207 (N_6207,N_6189,N_6047);
or U6208 (N_6208,N_6079,N_6058);
xnor U6209 (N_6209,N_6183,N_6069);
and U6210 (N_6210,N_6187,N_6169);
xnor U6211 (N_6211,N_6148,N_6007);
xor U6212 (N_6212,N_6190,N_6070);
xor U6213 (N_6213,N_6102,N_6173);
nor U6214 (N_6214,N_6133,N_6128);
or U6215 (N_6215,N_6160,N_6121);
or U6216 (N_6216,N_6197,N_6114);
nand U6217 (N_6217,N_6124,N_6171);
nor U6218 (N_6218,N_6170,N_6129);
nand U6219 (N_6219,N_6164,N_6181);
and U6220 (N_6220,N_6095,N_6146);
or U6221 (N_6221,N_6158,N_6065);
nand U6222 (N_6222,N_6060,N_6076);
or U6223 (N_6223,N_6175,N_6097);
nand U6224 (N_6224,N_6043,N_6142);
or U6225 (N_6225,N_6134,N_6059);
or U6226 (N_6226,N_6052,N_6176);
xnor U6227 (N_6227,N_6022,N_6089);
nor U6228 (N_6228,N_6081,N_6074);
nor U6229 (N_6229,N_6032,N_6083);
or U6230 (N_6230,N_6143,N_6162);
xnor U6231 (N_6231,N_6100,N_6174);
nand U6232 (N_6232,N_6101,N_6019);
xnor U6233 (N_6233,N_6149,N_6028);
or U6234 (N_6234,N_6077,N_6157);
or U6235 (N_6235,N_6178,N_6163);
nand U6236 (N_6236,N_6110,N_6150);
nor U6237 (N_6237,N_6046,N_6137);
xor U6238 (N_6238,N_6020,N_6055);
nor U6239 (N_6239,N_6013,N_6036);
xnor U6240 (N_6240,N_6122,N_6063);
nor U6241 (N_6241,N_6056,N_6027);
nor U6242 (N_6242,N_6082,N_6024);
or U6243 (N_6243,N_6011,N_6154);
nor U6244 (N_6244,N_6140,N_6194);
xor U6245 (N_6245,N_6172,N_6080);
nand U6246 (N_6246,N_6044,N_6002);
or U6247 (N_6247,N_6096,N_6057);
and U6248 (N_6248,N_6088,N_6188);
or U6249 (N_6249,N_6186,N_6015);
nor U6250 (N_6250,N_6039,N_6123);
and U6251 (N_6251,N_6118,N_6117);
or U6252 (N_6252,N_6033,N_6093);
xor U6253 (N_6253,N_6092,N_6042);
xnor U6254 (N_6254,N_6165,N_6131);
xnor U6255 (N_6255,N_6086,N_6116);
and U6256 (N_6256,N_6198,N_6021);
xnor U6257 (N_6257,N_6153,N_6066);
xor U6258 (N_6258,N_6008,N_6041);
or U6259 (N_6259,N_6072,N_6105);
or U6260 (N_6260,N_6054,N_6195);
or U6261 (N_6261,N_6155,N_6091);
and U6262 (N_6262,N_6156,N_6199);
or U6263 (N_6263,N_6000,N_6006);
xnor U6264 (N_6264,N_6045,N_6053);
and U6265 (N_6265,N_6180,N_6168);
xor U6266 (N_6266,N_6068,N_6005);
or U6267 (N_6267,N_6139,N_6037);
or U6268 (N_6268,N_6064,N_6023);
nor U6269 (N_6269,N_6111,N_6040);
and U6270 (N_6270,N_6184,N_6145);
nand U6271 (N_6271,N_6161,N_6004);
and U6272 (N_6272,N_6026,N_6135);
nor U6273 (N_6273,N_6109,N_6051);
xnor U6274 (N_6274,N_6003,N_6106);
xor U6275 (N_6275,N_6138,N_6182);
nor U6276 (N_6276,N_6029,N_6141);
xnor U6277 (N_6277,N_6099,N_6038);
nand U6278 (N_6278,N_6192,N_6196);
xnor U6279 (N_6279,N_6151,N_6034);
and U6280 (N_6280,N_6098,N_6067);
or U6281 (N_6281,N_6120,N_6193);
nand U6282 (N_6282,N_6030,N_6087);
nor U6283 (N_6283,N_6017,N_6012);
nor U6284 (N_6284,N_6094,N_6159);
nand U6285 (N_6285,N_6130,N_6103);
nand U6286 (N_6286,N_6119,N_6115);
or U6287 (N_6287,N_6126,N_6113);
xnor U6288 (N_6288,N_6085,N_6127);
xnor U6289 (N_6289,N_6035,N_6179);
and U6290 (N_6290,N_6185,N_6078);
nand U6291 (N_6291,N_6104,N_6031);
xor U6292 (N_6292,N_6016,N_6107);
and U6293 (N_6293,N_6152,N_6166);
xnor U6294 (N_6294,N_6073,N_6050);
xor U6295 (N_6295,N_6075,N_6049);
and U6296 (N_6296,N_6025,N_6014);
xnor U6297 (N_6297,N_6177,N_6108);
and U6298 (N_6298,N_6018,N_6125);
and U6299 (N_6299,N_6167,N_6132);
nor U6300 (N_6300,N_6017,N_6111);
xor U6301 (N_6301,N_6195,N_6066);
nand U6302 (N_6302,N_6142,N_6024);
or U6303 (N_6303,N_6038,N_6036);
or U6304 (N_6304,N_6187,N_6141);
nand U6305 (N_6305,N_6039,N_6007);
nor U6306 (N_6306,N_6145,N_6199);
and U6307 (N_6307,N_6106,N_6092);
xnor U6308 (N_6308,N_6068,N_6039);
xnor U6309 (N_6309,N_6192,N_6038);
nor U6310 (N_6310,N_6021,N_6078);
or U6311 (N_6311,N_6154,N_6144);
and U6312 (N_6312,N_6199,N_6049);
xor U6313 (N_6313,N_6040,N_6182);
xnor U6314 (N_6314,N_6057,N_6160);
and U6315 (N_6315,N_6134,N_6103);
xor U6316 (N_6316,N_6063,N_6092);
or U6317 (N_6317,N_6197,N_6155);
xnor U6318 (N_6318,N_6119,N_6038);
and U6319 (N_6319,N_6151,N_6063);
nor U6320 (N_6320,N_6189,N_6117);
xnor U6321 (N_6321,N_6190,N_6010);
nor U6322 (N_6322,N_6000,N_6122);
and U6323 (N_6323,N_6113,N_6045);
nand U6324 (N_6324,N_6179,N_6184);
xor U6325 (N_6325,N_6085,N_6158);
xnor U6326 (N_6326,N_6071,N_6064);
nor U6327 (N_6327,N_6130,N_6136);
xor U6328 (N_6328,N_6028,N_6102);
nand U6329 (N_6329,N_6190,N_6076);
nand U6330 (N_6330,N_6040,N_6133);
or U6331 (N_6331,N_6150,N_6059);
nor U6332 (N_6332,N_6040,N_6154);
xor U6333 (N_6333,N_6186,N_6196);
nor U6334 (N_6334,N_6034,N_6028);
and U6335 (N_6335,N_6130,N_6097);
nor U6336 (N_6336,N_6092,N_6154);
nand U6337 (N_6337,N_6035,N_6150);
nand U6338 (N_6338,N_6172,N_6120);
or U6339 (N_6339,N_6177,N_6009);
xor U6340 (N_6340,N_6147,N_6197);
or U6341 (N_6341,N_6043,N_6055);
nand U6342 (N_6342,N_6054,N_6137);
xor U6343 (N_6343,N_6043,N_6169);
nand U6344 (N_6344,N_6024,N_6177);
xnor U6345 (N_6345,N_6016,N_6124);
nor U6346 (N_6346,N_6121,N_6125);
nor U6347 (N_6347,N_6032,N_6113);
nand U6348 (N_6348,N_6085,N_6047);
nor U6349 (N_6349,N_6088,N_6093);
nor U6350 (N_6350,N_6031,N_6106);
nand U6351 (N_6351,N_6182,N_6061);
nor U6352 (N_6352,N_6006,N_6097);
nand U6353 (N_6353,N_6071,N_6029);
nor U6354 (N_6354,N_6132,N_6012);
nand U6355 (N_6355,N_6177,N_6011);
xor U6356 (N_6356,N_6133,N_6037);
or U6357 (N_6357,N_6162,N_6070);
or U6358 (N_6358,N_6035,N_6187);
nor U6359 (N_6359,N_6049,N_6140);
or U6360 (N_6360,N_6119,N_6012);
or U6361 (N_6361,N_6099,N_6048);
xnor U6362 (N_6362,N_6083,N_6177);
or U6363 (N_6363,N_6115,N_6013);
and U6364 (N_6364,N_6104,N_6181);
xnor U6365 (N_6365,N_6132,N_6029);
nand U6366 (N_6366,N_6137,N_6083);
and U6367 (N_6367,N_6040,N_6109);
nor U6368 (N_6368,N_6144,N_6050);
xnor U6369 (N_6369,N_6168,N_6003);
or U6370 (N_6370,N_6132,N_6051);
or U6371 (N_6371,N_6040,N_6020);
and U6372 (N_6372,N_6022,N_6111);
or U6373 (N_6373,N_6169,N_6120);
or U6374 (N_6374,N_6052,N_6166);
xor U6375 (N_6375,N_6063,N_6040);
xnor U6376 (N_6376,N_6186,N_6184);
and U6377 (N_6377,N_6135,N_6023);
or U6378 (N_6378,N_6183,N_6196);
nand U6379 (N_6379,N_6094,N_6029);
xnor U6380 (N_6380,N_6197,N_6050);
nand U6381 (N_6381,N_6148,N_6026);
xor U6382 (N_6382,N_6026,N_6109);
nand U6383 (N_6383,N_6090,N_6129);
and U6384 (N_6384,N_6057,N_6125);
nand U6385 (N_6385,N_6188,N_6080);
or U6386 (N_6386,N_6058,N_6049);
or U6387 (N_6387,N_6103,N_6083);
xnor U6388 (N_6388,N_6072,N_6066);
nand U6389 (N_6389,N_6127,N_6163);
xor U6390 (N_6390,N_6116,N_6143);
or U6391 (N_6391,N_6102,N_6086);
xor U6392 (N_6392,N_6061,N_6006);
nand U6393 (N_6393,N_6089,N_6097);
nor U6394 (N_6394,N_6069,N_6059);
or U6395 (N_6395,N_6134,N_6071);
or U6396 (N_6396,N_6076,N_6186);
nor U6397 (N_6397,N_6087,N_6011);
nor U6398 (N_6398,N_6015,N_6081);
and U6399 (N_6399,N_6002,N_6094);
nand U6400 (N_6400,N_6267,N_6291);
nand U6401 (N_6401,N_6353,N_6298);
or U6402 (N_6402,N_6302,N_6367);
nand U6403 (N_6403,N_6396,N_6274);
nand U6404 (N_6404,N_6352,N_6280);
or U6405 (N_6405,N_6384,N_6212);
or U6406 (N_6406,N_6284,N_6290);
and U6407 (N_6407,N_6234,N_6215);
nor U6408 (N_6408,N_6216,N_6255);
nor U6409 (N_6409,N_6305,N_6257);
and U6410 (N_6410,N_6209,N_6232);
xnor U6411 (N_6411,N_6286,N_6323);
nor U6412 (N_6412,N_6268,N_6242);
nor U6413 (N_6413,N_6301,N_6293);
and U6414 (N_6414,N_6303,N_6230);
xor U6415 (N_6415,N_6326,N_6392);
and U6416 (N_6416,N_6347,N_6233);
nor U6417 (N_6417,N_6208,N_6204);
xnor U6418 (N_6418,N_6377,N_6225);
nand U6419 (N_6419,N_6245,N_6357);
or U6420 (N_6420,N_6213,N_6235);
nor U6421 (N_6421,N_6358,N_6260);
or U6422 (N_6422,N_6254,N_6276);
or U6423 (N_6423,N_6288,N_6202);
nor U6424 (N_6424,N_6211,N_6334);
or U6425 (N_6425,N_6243,N_6217);
nand U6426 (N_6426,N_6341,N_6295);
nand U6427 (N_6427,N_6324,N_6318);
and U6428 (N_6428,N_6278,N_6256);
xor U6429 (N_6429,N_6389,N_6344);
xnor U6430 (N_6430,N_6348,N_6270);
and U6431 (N_6431,N_6244,N_6259);
nor U6432 (N_6432,N_6361,N_6360);
or U6433 (N_6433,N_6201,N_6397);
nor U6434 (N_6434,N_6369,N_6387);
xnor U6435 (N_6435,N_6264,N_6335);
nand U6436 (N_6436,N_6240,N_6206);
xnor U6437 (N_6437,N_6218,N_6246);
or U6438 (N_6438,N_6277,N_6214);
nand U6439 (N_6439,N_6336,N_6252);
or U6440 (N_6440,N_6329,N_6289);
xor U6441 (N_6441,N_6351,N_6356);
and U6442 (N_6442,N_6381,N_6363);
nor U6443 (N_6443,N_6285,N_6330);
and U6444 (N_6444,N_6247,N_6379);
nand U6445 (N_6445,N_6287,N_6383);
or U6446 (N_6446,N_6390,N_6297);
nand U6447 (N_6447,N_6258,N_6299);
or U6448 (N_6448,N_6273,N_6313);
nor U6449 (N_6449,N_6393,N_6269);
and U6450 (N_6450,N_6311,N_6370);
and U6451 (N_6451,N_6325,N_6333);
or U6452 (N_6452,N_6223,N_6316);
or U6453 (N_6453,N_6275,N_6261);
nand U6454 (N_6454,N_6307,N_6385);
and U6455 (N_6455,N_6251,N_6283);
xor U6456 (N_6456,N_6321,N_6391);
nor U6457 (N_6457,N_6374,N_6364);
nand U6458 (N_6458,N_6312,N_6343);
nor U6459 (N_6459,N_6355,N_6395);
xor U6460 (N_6460,N_6386,N_6376);
nor U6461 (N_6461,N_6362,N_6237);
xnor U6462 (N_6462,N_6310,N_6203);
xnor U6463 (N_6463,N_6372,N_6339);
xor U6464 (N_6464,N_6226,N_6296);
or U6465 (N_6465,N_6236,N_6375);
and U6466 (N_6466,N_6373,N_6319);
xnor U6467 (N_6467,N_6342,N_6365);
nor U6468 (N_6468,N_6345,N_6294);
or U6469 (N_6469,N_6262,N_6281);
or U6470 (N_6470,N_6368,N_6228);
nor U6471 (N_6471,N_6327,N_6309);
nand U6472 (N_6472,N_6322,N_6315);
nor U6473 (N_6473,N_6388,N_6219);
nand U6474 (N_6474,N_6338,N_6227);
and U6475 (N_6475,N_6354,N_6231);
xnor U6476 (N_6476,N_6253,N_6317);
or U6477 (N_6477,N_6249,N_6399);
or U6478 (N_6478,N_6207,N_6200);
xor U6479 (N_6479,N_6263,N_6220);
nor U6480 (N_6480,N_6265,N_6314);
nand U6481 (N_6481,N_6282,N_6349);
xnor U6482 (N_6482,N_6359,N_6378);
or U6483 (N_6483,N_6350,N_6320);
xor U6484 (N_6484,N_6221,N_6346);
and U6485 (N_6485,N_6308,N_6300);
xor U6486 (N_6486,N_6304,N_6328);
nand U6487 (N_6487,N_6229,N_6394);
xor U6488 (N_6488,N_6272,N_6248);
nor U6489 (N_6489,N_6340,N_6279);
nor U6490 (N_6490,N_6250,N_6366);
nand U6491 (N_6491,N_6332,N_6238);
or U6492 (N_6492,N_6210,N_6224);
nor U6493 (N_6493,N_6382,N_6292);
xnor U6494 (N_6494,N_6222,N_6271);
or U6495 (N_6495,N_6266,N_6306);
nand U6496 (N_6496,N_6239,N_6241);
or U6497 (N_6497,N_6371,N_6380);
and U6498 (N_6498,N_6337,N_6398);
and U6499 (N_6499,N_6205,N_6331);
xnor U6500 (N_6500,N_6279,N_6241);
and U6501 (N_6501,N_6278,N_6398);
and U6502 (N_6502,N_6330,N_6291);
nor U6503 (N_6503,N_6255,N_6262);
nand U6504 (N_6504,N_6391,N_6277);
and U6505 (N_6505,N_6240,N_6291);
or U6506 (N_6506,N_6270,N_6260);
xnor U6507 (N_6507,N_6225,N_6315);
nand U6508 (N_6508,N_6209,N_6300);
or U6509 (N_6509,N_6310,N_6275);
and U6510 (N_6510,N_6284,N_6202);
nor U6511 (N_6511,N_6331,N_6337);
nor U6512 (N_6512,N_6263,N_6222);
or U6513 (N_6513,N_6329,N_6321);
xnor U6514 (N_6514,N_6288,N_6270);
nand U6515 (N_6515,N_6300,N_6205);
nand U6516 (N_6516,N_6264,N_6289);
and U6517 (N_6517,N_6354,N_6259);
or U6518 (N_6518,N_6245,N_6202);
xor U6519 (N_6519,N_6252,N_6236);
or U6520 (N_6520,N_6330,N_6287);
or U6521 (N_6521,N_6227,N_6350);
nor U6522 (N_6522,N_6322,N_6368);
nor U6523 (N_6523,N_6338,N_6384);
nor U6524 (N_6524,N_6296,N_6232);
or U6525 (N_6525,N_6284,N_6294);
nor U6526 (N_6526,N_6224,N_6323);
nand U6527 (N_6527,N_6325,N_6245);
nand U6528 (N_6528,N_6385,N_6245);
nor U6529 (N_6529,N_6326,N_6217);
or U6530 (N_6530,N_6368,N_6220);
nand U6531 (N_6531,N_6397,N_6303);
xnor U6532 (N_6532,N_6207,N_6361);
or U6533 (N_6533,N_6205,N_6364);
or U6534 (N_6534,N_6347,N_6340);
nand U6535 (N_6535,N_6215,N_6261);
nor U6536 (N_6536,N_6373,N_6363);
and U6537 (N_6537,N_6292,N_6229);
nor U6538 (N_6538,N_6241,N_6322);
nand U6539 (N_6539,N_6280,N_6360);
and U6540 (N_6540,N_6311,N_6249);
nor U6541 (N_6541,N_6385,N_6386);
or U6542 (N_6542,N_6305,N_6347);
or U6543 (N_6543,N_6257,N_6252);
nand U6544 (N_6544,N_6338,N_6253);
xor U6545 (N_6545,N_6341,N_6200);
xnor U6546 (N_6546,N_6253,N_6320);
xor U6547 (N_6547,N_6349,N_6389);
xor U6548 (N_6548,N_6280,N_6241);
or U6549 (N_6549,N_6368,N_6309);
xnor U6550 (N_6550,N_6330,N_6325);
nor U6551 (N_6551,N_6331,N_6288);
nand U6552 (N_6552,N_6207,N_6334);
nor U6553 (N_6553,N_6307,N_6260);
or U6554 (N_6554,N_6286,N_6218);
and U6555 (N_6555,N_6330,N_6388);
or U6556 (N_6556,N_6348,N_6255);
nand U6557 (N_6557,N_6393,N_6216);
and U6558 (N_6558,N_6325,N_6315);
and U6559 (N_6559,N_6311,N_6373);
or U6560 (N_6560,N_6227,N_6270);
nor U6561 (N_6561,N_6242,N_6292);
nand U6562 (N_6562,N_6291,N_6263);
or U6563 (N_6563,N_6368,N_6205);
xnor U6564 (N_6564,N_6244,N_6378);
nand U6565 (N_6565,N_6355,N_6296);
nand U6566 (N_6566,N_6300,N_6258);
or U6567 (N_6567,N_6261,N_6217);
or U6568 (N_6568,N_6291,N_6351);
nor U6569 (N_6569,N_6200,N_6283);
xnor U6570 (N_6570,N_6240,N_6390);
nor U6571 (N_6571,N_6207,N_6218);
nor U6572 (N_6572,N_6254,N_6389);
nand U6573 (N_6573,N_6264,N_6240);
nor U6574 (N_6574,N_6234,N_6283);
and U6575 (N_6575,N_6259,N_6276);
xor U6576 (N_6576,N_6234,N_6322);
xor U6577 (N_6577,N_6228,N_6379);
xor U6578 (N_6578,N_6259,N_6315);
xor U6579 (N_6579,N_6201,N_6243);
nand U6580 (N_6580,N_6393,N_6204);
xor U6581 (N_6581,N_6337,N_6234);
nand U6582 (N_6582,N_6352,N_6330);
or U6583 (N_6583,N_6332,N_6266);
and U6584 (N_6584,N_6362,N_6250);
nand U6585 (N_6585,N_6380,N_6319);
nand U6586 (N_6586,N_6237,N_6270);
xnor U6587 (N_6587,N_6392,N_6370);
xor U6588 (N_6588,N_6366,N_6277);
nor U6589 (N_6589,N_6231,N_6369);
nor U6590 (N_6590,N_6211,N_6394);
and U6591 (N_6591,N_6281,N_6321);
xor U6592 (N_6592,N_6342,N_6348);
nor U6593 (N_6593,N_6203,N_6314);
and U6594 (N_6594,N_6321,N_6358);
nand U6595 (N_6595,N_6269,N_6338);
nand U6596 (N_6596,N_6304,N_6380);
xor U6597 (N_6597,N_6327,N_6364);
and U6598 (N_6598,N_6253,N_6354);
and U6599 (N_6599,N_6244,N_6368);
nand U6600 (N_6600,N_6499,N_6598);
nor U6601 (N_6601,N_6472,N_6426);
nor U6602 (N_6602,N_6455,N_6527);
or U6603 (N_6603,N_6479,N_6456);
xnor U6604 (N_6604,N_6594,N_6484);
xor U6605 (N_6605,N_6563,N_6558);
or U6606 (N_6606,N_6464,N_6517);
xnor U6607 (N_6607,N_6581,N_6588);
and U6608 (N_6608,N_6593,N_6437);
nor U6609 (N_6609,N_6431,N_6512);
and U6610 (N_6610,N_6539,N_6515);
nor U6611 (N_6611,N_6599,N_6532);
xor U6612 (N_6612,N_6438,N_6490);
nor U6613 (N_6613,N_6414,N_6468);
and U6614 (N_6614,N_6425,N_6434);
xnor U6615 (N_6615,N_6502,N_6582);
nand U6616 (N_6616,N_6510,N_6530);
or U6617 (N_6617,N_6554,N_6422);
or U6618 (N_6618,N_6404,N_6578);
nor U6619 (N_6619,N_6571,N_6442);
or U6620 (N_6620,N_6560,N_6500);
nor U6621 (N_6621,N_6580,N_6548);
or U6622 (N_6622,N_6595,N_6450);
and U6623 (N_6623,N_6522,N_6482);
and U6624 (N_6624,N_6400,N_6430);
nand U6625 (N_6625,N_6424,N_6494);
and U6626 (N_6626,N_6576,N_6407);
and U6627 (N_6627,N_6474,N_6497);
or U6628 (N_6628,N_6546,N_6496);
nand U6629 (N_6629,N_6592,N_6421);
nand U6630 (N_6630,N_6433,N_6428);
nand U6631 (N_6631,N_6403,N_6534);
and U6632 (N_6632,N_6507,N_6480);
or U6633 (N_6633,N_6445,N_6493);
nand U6634 (N_6634,N_6524,N_6568);
xor U6635 (N_6635,N_6420,N_6491);
or U6636 (N_6636,N_6516,N_6543);
nor U6637 (N_6637,N_6467,N_6526);
nand U6638 (N_6638,N_6409,N_6401);
nor U6639 (N_6639,N_6521,N_6441);
xnor U6640 (N_6640,N_6531,N_6410);
and U6641 (N_6641,N_6478,N_6448);
nor U6642 (N_6642,N_6462,N_6565);
xor U6643 (N_6643,N_6569,N_6589);
or U6644 (N_6644,N_6460,N_6453);
xnor U6645 (N_6645,N_6585,N_6423);
nand U6646 (N_6646,N_6485,N_6454);
nand U6647 (N_6647,N_6457,N_6488);
or U6648 (N_6648,N_6519,N_6486);
nor U6649 (N_6649,N_6575,N_6473);
and U6650 (N_6650,N_6597,N_6552);
and U6651 (N_6651,N_6528,N_6529);
xnor U6652 (N_6652,N_6447,N_6550);
and U6653 (N_6653,N_6412,N_6446);
and U6654 (N_6654,N_6536,N_6542);
and U6655 (N_6655,N_6570,N_6574);
or U6656 (N_6656,N_6406,N_6476);
or U6657 (N_6657,N_6465,N_6587);
and U6658 (N_6658,N_6544,N_6583);
or U6659 (N_6659,N_6561,N_6432);
or U6660 (N_6660,N_6564,N_6440);
nand U6661 (N_6661,N_6419,N_6596);
xnor U6662 (N_6662,N_6525,N_6584);
xnor U6663 (N_6663,N_6503,N_6509);
and U6664 (N_6664,N_6439,N_6572);
nor U6665 (N_6665,N_6586,N_6402);
and U6666 (N_6666,N_6540,N_6506);
nor U6667 (N_6667,N_6449,N_6477);
xnor U6668 (N_6668,N_6466,N_6579);
or U6669 (N_6669,N_6487,N_6508);
nand U6670 (N_6670,N_6523,N_6538);
or U6671 (N_6671,N_6418,N_6498);
nand U6672 (N_6672,N_6555,N_6417);
nand U6673 (N_6673,N_6567,N_6415);
or U6674 (N_6674,N_6411,N_6444);
nand U6675 (N_6675,N_6470,N_6501);
or U6676 (N_6676,N_6562,N_6459);
and U6677 (N_6677,N_6429,N_6443);
nor U6678 (N_6678,N_6551,N_6408);
nor U6679 (N_6679,N_6591,N_6435);
nor U6680 (N_6680,N_6436,N_6495);
or U6681 (N_6681,N_6452,N_6545);
and U6682 (N_6682,N_6413,N_6577);
nor U6683 (N_6683,N_6556,N_6547);
or U6684 (N_6684,N_6475,N_6590);
nand U6685 (N_6685,N_6513,N_6427);
nor U6686 (N_6686,N_6416,N_6471);
nor U6687 (N_6687,N_6505,N_6518);
nand U6688 (N_6688,N_6557,N_6520);
nor U6689 (N_6689,N_6405,N_6537);
xnor U6690 (N_6690,N_6533,N_6514);
and U6691 (N_6691,N_6535,N_6481);
or U6692 (N_6692,N_6469,N_6451);
and U6693 (N_6693,N_6483,N_6461);
and U6694 (N_6694,N_6573,N_6553);
and U6695 (N_6695,N_6489,N_6549);
and U6696 (N_6696,N_6463,N_6559);
and U6697 (N_6697,N_6504,N_6458);
xor U6698 (N_6698,N_6566,N_6541);
xor U6699 (N_6699,N_6511,N_6492);
xor U6700 (N_6700,N_6510,N_6518);
nor U6701 (N_6701,N_6428,N_6425);
and U6702 (N_6702,N_6455,N_6495);
or U6703 (N_6703,N_6544,N_6464);
and U6704 (N_6704,N_6580,N_6449);
and U6705 (N_6705,N_6570,N_6465);
and U6706 (N_6706,N_6569,N_6499);
nor U6707 (N_6707,N_6435,N_6574);
xor U6708 (N_6708,N_6582,N_6528);
nand U6709 (N_6709,N_6522,N_6544);
xnor U6710 (N_6710,N_6500,N_6447);
nor U6711 (N_6711,N_6508,N_6489);
xnor U6712 (N_6712,N_6597,N_6442);
and U6713 (N_6713,N_6453,N_6572);
xor U6714 (N_6714,N_6475,N_6508);
xor U6715 (N_6715,N_6440,N_6403);
and U6716 (N_6716,N_6404,N_6552);
nand U6717 (N_6717,N_6534,N_6553);
and U6718 (N_6718,N_6513,N_6415);
and U6719 (N_6719,N_6587,N_6411);
nand U6720 (N_6720,N_6452,N_6471);
nand U6721 (N_6721,N_6534,N_6463);
xnor U6722 (N_6722,N_6459,N_6494);
nor U6723 (N_6723,N_6486,N_6523);
or U6724 (N_6724,N_6551,N_6466);
nor U6725 (N_6725,N_6502,N_6538);
or U6726 (N_6726,N_6470,N_6588);
xnor U6727 (N_6727,N_6504,N_6428);
xnor U6728 (N_6728,N_6429,N_6570);
nor U6729 (N_6729,N_6475,N_6458);
nand U6730 (N_6730,N_6546,N_6423);
or U6731 (N_6731,N_6580,N_6559);
nor U6732 (N_6732,N_6592,N_6560);
and U6733 (N_6733,N_6420,N_6402);
nor U6734 (N_6734,N_6429,N_6584);
xor U6735 (N_6735,N_6571,N_6579);
or U6736 (N_6736,N_6592,N_6413);
nor U6737 (N_6737,N_6583,N_6587);
and U6738 (N_6738,N_6496,N_6513);
xor U6739 (N_6739,N_6554,N_6519);
xor U6740 (N_6740,N_6474,N_6418);
or U6741 (N_6741,N_6506,N_6570);
nand U6742 (N_6742,N_6446,N_6528);
or U6743 (N_6743,N_6593,N_6498);
nand U6744 (N_6744,N_6437,N_6575);
and U6745 (N_6745,N_6533,N_6493);
and U6746 (N_6746,N_6568,N_6532);
nand U6747 (N_6747,N_6558,N_6529);
xor U6748 (N_6748,N_6583,N_6463);
nand U6749 (N_6749,N_6462,N_6579);
xor U6750 (N_6750,N_6401,N_6506);
or U6751 (N_6751,N_6597,N_6521);
or U6752 (N_6752,N_6482,N_6538);
nand U6753 (N_6753,N_6572,N_6480);
and U6754 (N_6754,N_6584,N_6406);
nand U6755 (N_6755,N_6482,N_6514);
nor U6756 (N_6756,N_6406,N_6588);
or U6757 (N_6757,N_6576,N_6433);
nor U6758 (N_6758,N_6586,N_6478);
and U6759 (N_6759,N_6508,N_6484);
nor U6760 (N_6760,N_6585,N_6513);
nor U6761 (N_6761,N_6426,N_6474);
xnor U6762 (N_6762,N_6445,N_6523);
nor U6763 (N_6763,N_6574,N_6525);
nor U6764 (N_6764,N_6518,N_6454);
xnor U6765 (N_6765,N_6426,N_6596);
xnor U6766 (N_6766,N_6409,N_6547);
or U6767 (N_6767,N_6574,N_6575);
xor U6768 (N_6768,N_6555,N_6408);
nor U6769 (N_6769,N_6529,N_6542);
nor U6770 (N_6770,N_6517,N_6577);
nand U6771 (N_6771,N_6432,N_6522);
nor U6772 (N_6772,N_6444,N_6532);
or U6773 (N_6773,N_6538,N_6412);
or U6774 (N_6774,N_6584,N_6593);
xor U6775 (N_6775,N_6574,N_6486);
xnor U6776 (N_6776,N_6544,N_6454);
xnor U6777 (N_6777,N_6427,N_6554);
and U6778 (N_6778,N_6540,N_6590);
xnor U6779 (N_6779,N_6466,N_6442);
nor U6780 (N_6780,N_6583,N_6540);
nand U6781 (N_6781,N_6587,N_6452);
or U6782 (N_6782,N_6464,N_6574);
xor U6783 (N_6783,N_6406,N_6554);
nor U6784 (N_6784,N_6566,N_6472);
xnor U6785 (N_6785,N_6416,N_6467);
xor U6786 (N_6786,N_6599,N_6421);
or U6787 (N_6787,N_6423,N_6557);
nor U6788 (N_6788,N_6428,N_6429);
nor U6789 (N_6789,N_6563,N_6459);
and U6790 (N_6790,N_6449,N_6424);
and U6791 (N_6791,N_6409,N_6561);
or U6792 (N_6792,N_6448,N_6503);
and U6793 (N_6793,N_6419,N_6462);
xnor U6794 (N_6794,N_6574,N_6577);
xnor U6795 (N_6795,N_6513,N_6468);
xor U6796 (N_6796,N_6457,N_6404);
or U6797 (N_6797,N_6439,N_6512);
nand U6798 (N_6798,N_6561,N_6476);
and U6799 (N_6799,N_6415,N_6429);
and U6800 (N_6800,N_6730,N_6651);
xor U6801 (N_6801,N_6676,N_6609);
nand U6802 (N_6802,N_6661,N_6718);
xnor U6803 (N_6803,N_6741,N_6755);
nand U6804 (N_6804,N_6637,N_6633);
nand U6805 (N_6805,N_6725,N_6796);
xor U6806 (N_6806,N_6789,N_6762);
or U6807 (N_6807,N_6715,N_6620);
and U6808 (N_6808,N_6728,N_6736);
nor U6809 (N_6809,N_6785,N_6663);
and U6810 (N_6810,N_6703,N_6775);
nor U6811 (N_6811,N_6691,N_6710);
or U6812 (N_6812,N_6756,N_6722);
nand U6813 (N_6813,N_6662,N_6638);
or U6814 (N_6814,N_6717,N_6660);
nor U6815 (N_6815,N_6742,N_6679);
nor U6816 (N_6816,N_6708,N_6761);
nand U6817 (N_6817,N_6772,N_6634);
nand U6818 (N_6818,N_6681,N_6607);
nand U6819 (N_6819,N_6626,N_6774);
or U6820 (N_6820,N_6746,N_6733);
xor U6821 (N_6821,N_6677,N_6627);
nand U6822 (N_6822,N_6606,N_6683);
or U6823 (N_6823,N_6667,N_6668);
or U6824 (N_6824,N_6738,N_6793);
xor U6825 (N_6825,N_6672,N_6768);
nor U6826 (N_6826,N_6619,N_6754);
xnor U6827 (N_6827,N_6763,N_6674);
or U6828 (N_6828,N_6686,N_6706);
nor U6829 (N_6829,N_6630,N_6740);
or U6830 (N_6830,N_6723,N_6605);
xnor U6831 (N_6831,N_6788,N_6751);
or U6832 (N_6832,N_6747,N_6799);
or U6833 (N_6833,N_6743,N_6732);
or U6834 (N_6834,N_6666,N_6680);
nand U6835 (N_6835,N_6776,N_6645);
and U6836 (N_6836,N_6658,N_6659);
nor U6837 (N_6837,N_6695,N_6713);
nor U6838 (N_6838,N_6734,N_6781);
and U6839 (N_6839,N_6798,N_6650);
and U6840 (N_6840,N_6783,N_6694);
or U6841 (N_6841,N_6735,N_6737);
and U6842 (N_6842,N_6636,N_6639);
nand U6843 (N_6843,N_6702,N_6784);
or U6844 (N_6844,N_6608,N_6601);
xnor U6845 (N_6845,N_6682,N_6787);
nor U6846 (N_6846,N_6640,N_6709);
and U6847 (N_6847,N_6675,N_6777);
xnor U6848 (N_6848,N_6687,N_6729);
nor U6849 (N_6849,N_6611,N_6773);
nor U6850 (N_6850,N_6724,N_6669);
xnor U6851 (N_6851,N_6649,N_6684);
or U6852 (N_6852,N_6720,N_6794);
nand U6853 (N_6853,N_6604,N_6616);
xnor U6854 (N_6854,N_6644,N_6707);
and U6855 (N_6855,N_6642,N_6771);
nor U6856 (N_6856,N_6646,N_6665);
or U6857 (N_6857,N_6652,N_6778);
xor U6858 (N_6858,N_6750,N_6690);
or U6859 (N_6859,N_6745,N_6765);
xnor U6860 (N_6860,N_6780,N_6602);
xnor U6861 (N_6861,N_6716,N_6657);
nor U6862 (N_6862,N_6625,N_6739);
or U6863 (N_6863,N_6617,N_6635);
nand U6864 (N_6864,N_6757,N_6603);
xnor U6865 (N_6865,N_6767,N_6622);
and U6866 (N_6866,N_6779,N_6610);
xnor U6867 (N_6867,N_6795,N_6760);
nor U6868 (N_6868,N_6701,N_6647);
nand U6869 (N_6869,N_6719,N_6643);
nand U6870 (N_6870,N_6670,N_6654);
xor U6871 (N_6871,N_6698,N_6731);
and U6872 (N_6872,N_6697,N_6671);
nand U6873 (N_6873,N_6759,N_6700);
nor U6874 (N_6874,N_6621,N_6692);
nor U6875 (N_6875,N_6749,N_6678);
nor U6876 (N_6876,N_6614,N_6753);
xor U6877 (N_6877,N_6766,N_6615);
and U6878 (N_6878,N_6726,N_6699);
and U6879 (N_6879,N_6688,N_6712);
nor U6880 (N_6880,N_6653,N_6748);
nand U6881 (N_6881,N_6790,N_6769);
nor U6882 (N_6882,N_6689,N_6721);
nor U6883 (N_6883,N_6632,N_6624);
nand U6884 (N_6884,N_6628,N_6656);
nand U6885 (N_6885,N_6782,N_6696);
xnor U6886 (N_6886,N_6764,N_6631);
xor U6887 (N_6887,N_6613,N_6704);
xnor U6888 (N_6888,N_6711,N_6623);
and U6889 (N_6889,N_6752,N_6664);
or U6890 (N_6890,N_6786,N_6648);
nor U6891 (N_6891,N_6693,N_6673);
nor U6892 (N_6892,N_6612,N_6727);
xor U6893 (N_6893,N_6600,N_6797);
xnor U6894 (N_6894,N_6770,N_6791);
nor U6895 (N_6895,N_6792,N_6629);
xnor U6896 (N_6896,N_6705,N_6744);
nand U6897 (N_6897,N_6758,N_6655);
nand U6898 (N_6898,N_6714,N_6685);
nor U6899 (N_6899,N_6641,N_6618);
nand U6900 (N_6900,N_6733,N_6750);
nand U6901 (N_6901,N_6746,N_6730);
nand U6902 (N_6902,N_6646,N_6678);
or U6903 (N_6903,N_6722,N_6625);
or U6904 (N_6904,N_6715,N_6749);
or U6905 (N_6905,N_6797,N_6786);
xor U6906 (N_6906,N_6781,N_6682);
nand U6907 (N_6907,N_6635,N_6681);
nor U6908 (N_6908,N_6764,N_6660);
xor U6909 (N_6909,N_6627,N_6745);
nor U6910 (N_6910,N_6634,N_6612);
nand U6911 (N_6911,N_6687,N_6706);
nor U6912 (N_6912,N_6729,N_6694);
and U6913 (N_6913,N_6741,N_6697);
or U6914 (N_6914,N_6760,N_6718);
nor U6915 (N_6915,N_6673,N_6709);
nand U6916 (N_6916,N_6687,N_6786);
xnor U6917 (N_6917,N_6762,N_6616);
nand U6918 (N_6918,N_6646,N_6739);
and U6919 (N_6919,N_6797,N_6692);
nand U6920 (N_6920,N_6716,N_6754);
or U6921 (N_6921,N_6612,N_6619);
or U6922 (N_6922,N_6647,N_6792);
nor U6923 (N_6923,N_6675,N_6680);
nor U6924 (N_6924,N_6736,N_6797);
or U6925 (N_6925,N_6705,N_6684);
or U6926 (N_6926,N_6739,N_6768);
nand U6927 (N_6927,N_6707,N_6629);
or U6928 (N_6928,N_6725,N_6664);
nor U6929 (N_6929,N_6613,N_6689);
nor U6930 (N_6930,N_6740,N_6704);
xor U6931 (N_6931,N_6710,N_6712);
or U6932 (N_6932,N_6788,N_6748);
nand U6933 (N_6933,N_6799,N_6734);
xor U6934 (N_6934,N_6767,N_6759);
or U6935 (N_6935,N_6716,N_6717);
or U6936 (N_6936,N_6739,N_6602);
nor U6937 (N_6937,N_6769,N_6761);
xnor U6938 (N_6938,N_6661,N_6644);
nor U6939 (N_6939,N_6787,N_6616);
xor U6940 (N_6940,N_6755,N_6680);
xor U6941 (N_6941,N_6624,N_6681);
xnor U6942 (N_6942,N_6612,N_6663);
nand U6943 (N_6943,N_6623,N_6729);
xor U6944 (N_6944,N_6738,N_6619);
or U6945 (N_6945,N_6603,N_6685);
xnor U6946 (N_6946,N_6632,N_6780);
and U6947 (N_6947,N_6702,N_6727);
nor U6948 (N_6948,N_6671,N_6764);
or U6949 (N_6949,N_6669,N_6723);
xnor U6950 (N_6950,N_6781,N_6608);
nand U6951 (N_6951,N_6695,N_6614);
nand U6952 (N_6952,N_6631,N_6797);
nor U6953 (N_6953,N_6743,N_6615);
or U6954 (N_6954,N_6798,N_6712);
xor U6955 (N_6955,N_6657,N_6690);
or U6956 (N_6956,N_6663,N_6718);
and U6957 (N_6957,N_6714,N_6667);
or U6958 (N_6958,N_6638,N_6719);
and U6959 (N_6959,N_6722,N_6637);
nand U6960 (N_6960,N_6652,N_6718);
and U6961 (N_6961,N_6613,N_6630);
xnor U6962 (N_6962,N_6695,N_6736);
nor U6963 (N_6963,N_6609,N_6718);
and U6964 (N_6964,N_6603,N_6700);
xnor U6965 (N_6965,N_6682,N_6603);
xnor U6966 (N_6966,N_6695,N_6717);
and U6967 (N_6967,N_6625,N_6659);
and U6968 (N_6968,N_6638,N_6798);
or U6969 (N_6969,N_6789,N_6701);
xnor U6970 (N_6970,N_6667,N_6736);
xnor U6971 (N_6971,N_6760,N_6623);
nand U6972 (N_6972,N_6682,N_6777);
and U6973 (N_6973,N_6738,N_6794);
xor U6974 (N_6974,N_6716,N_6712);
or U6975 (N_6975,N_6603,N_6779);
and U6976 (N_6976,N_6618,N_6672);
nor U6977 (N_6977,N_6624,N_6676);
or U6978 (N_6978,N_6795,N_6672);
or U6979 (N_6979,N_6798,N_6721);
xnor U6980 (N_6980,N_6613,N_6719);
xnor U6981 (N_6981,N_6637,N_6769);
nor U6982 (N_6982,N_6787,N_6799);
xor U6983 (N_6983,N_6704,N_6743);
nand U6984 (N_6984,N_6679,N_6784);
and U6985 (N_6985,N_6724,N_6682);
xor U6986 (N_6986,N_6676,N_6684);
xor U6987 (N_6987,N_6781,N_6787);
and U6988 (N_6988,N_6743,N_6783);
xnor U6989 (N_6989,N_6799,N_6644);
nand U6990 (N_6990,N_6763,N_6776);
xor U6991 (N_6991,N_6634,N_6739);
xnor U6992 (N_6992,N_6648,N_6617);
nand U6993 (N_6993,N_6724,N_6717);
nor U6994 (N_6994,N_6647,N_6668);
xor U6995 (N_6995,N_6623,N_6744);
nor U6996 (N_6996,N_6667,N_6719);
nor U6997 (N_6997,N_6626,N_6752);
and U6998 (N_6998,N_6771,N_6669);
nor U6999 (N_6999,N_6697,N_6666);
and U7000 (N_7000,N_6871,N_6807);
xor U7001 (N_7001,N_6835,N_6929);
and U7002 (N_7002,N_6952,N_6914);
xor U7003 (N_7003,N_6859,N_6974);
xor U7004 (N_7004,N_6831,N_6959);
or U7005 (N_7005,N_6842,N_6918);
and U7006 (N_7006,N_6978,N_6957);
or U7007 (N_7007,N_6970,N_6839);
and U7008 (N_7008,N_6927,N_6928);
xnor U7009 (N_7009,N_6853,N_6900);
xnor U7010 (N_7010,N_6815,N_6947);
nand U7011 (N_7011,N_6820,N_6850);
xnor U7012 (N_7012,N_6823,N_6824);
nand U7013 (N_7013,N_6896,N_6955);
nand U7014 (N_7014,N_6817,N_6979);
xnor U7015 (N_7015,N_6805,N_6991);
xnor U7016 (N_7016,N_6884,N_6951);
or U7017 (N_7017,N_6844,N_6862);
nand U7018 (N_7018,N_6975,N_6892);
or U7019 (N_7019,N_6837,N_6933);
xnor U7020 (N_7020,N_6990,N_6827);
nand U7021 (N_7021,N_6903,N_6941);
xnor U7022 (N_7022,N_6905,N_6940);
nand U7023 (N_7023,N_6982,N_6867);
nor U7024 (N_7024,N_6911,N_6986);
nand U7025 (N_7025,N_6998,N_6804);
nor U7026 (N_7026,N_6973,N_6812);
nor U7027 (N_7027,N_6818,N_6863);
xor U7028 (N_7028,N_6856,N_6981);
or U7029 (N_7029,N_6907,N_6870);
xor U7030 (N_7030,N_6932,N_6864);
or U7031 (N_7031,N_6891,N_6868);
xor U7032 (N_7032,N_6936,N_6874);
xor U7033 (N_7033,N_6972,N_6888);
nand U7034 (N_7034,N_6886,N_6917);
and U7035 (N_7035,N_6883,N_6920);
xor U7036 (N_7036,N_6816,N_6866);
and U7037 (N_7037,N_6819,N_6953);
nor U7038 (N_7038,N_6915,N_6993);
or U7039 (N_7039,N_6985,N_6930);
and U7040 (N_7040,N_6901,N_6832);
or U7041 (N_7041,N_6987,N_6875);
or U7042 (N_7042,N_6880,N_6814);
xor U7043 (N_7043,N_6865,N_6902);
nor U7044 (N_7044,N_6899,N_6904);
or U7045 (N_7045,N_6833,N_6912);
or U7046 (N_7046,N_6822,N_6997);
nor U7047 (N_7047,N_6942,N_6977);
nand U7048 (N_7048,N_6906,N_6924);
nor U7049 (N_7049,N_6836,N_6908);
nand U7050 (N_7050,N_6829,N_6960);
xnor U7051 (N_7051,N_6992,N_6821);
nand U7052 (N_7052,N_6950,N_6931);
nand U7053 (N_7053,N_6848,N_6855);
or U7054 (N_7054,N_6857,N_6858);
nor U7055 (N_7055,N_6995,N_6845);
and U7056 (N_7056,N_6935,N_6851);
xor U7057 (N_7057,N_6889,N_6852);
nor U7058 (N_7058,N_6800,N_6963);
nand U7059 (N_7059,N_6898,N_6872);
and U7060 (N_7060,N_6954,N_6873);
nand U7061 (N_7061,N_6847,N_6809);
and U7062 (N_7062,N_6802,N_6897);
nor U7063 (N_7063,N_6937,N_6962);
nand U7064 (N_7064,N_6830,N_6885);
nand U7065 (N_7065,N_6968,N_6948);
or U7066 (N_7066,N_6909,N_6934);
xor U7067 (N_7067,N_6910,N_6984);
and U7068 (N_7068,N_6840,N_6943);
nand U7069 (N_7069,N_6980,N_6877);
nand U7070 (N_7070,N_6861,N_6989);
nor U7071 (N_7071,N_6834,N_6882);
or U7072 (N_7072,N_6921,N_6879);
xnor U7073 (N_7073,N_6876,N_6976);
nand U7074 (N_7074,N_6838,N_6826);
xor U7075 (N_7075,N_6843,N_6841);
xnor U7076 (N_7076,N_6916,N_6988);
or U7077 (N_7077,N_6849,N_6944);
xnor U7078 (N_7078,N_6971,N_6945);
nor U7079 (N_7079,N_6894,N_6887);
nor U7080 (N_7080,N_6808,N_6811);
and U7081 (N_7081,N_6994,N_6922);
nand U7082 (N_7082,N_6893,N_6828);
or U7083 (N_7083,N_6961,N_6913);
or U7084 (N_7084,N_6938,N_6996);
nor U7085 (N_7085,N_6881,N_6810);
nand U7086 (N_7086,N_6869,N_6969);
nand U7087 (N_7087,N_6983,N_6967);
xor U7088 (N_7088,N_6806,N_6958);
xor U7089 (N_7089,N_6946,N_6965);
nor U7090 (N_7090,N_6966,N_6925);
xnor U7091 (N_7091,N_6964,N_6926);
nor U7092 (N_7092,N_6890,N_6854);
nand U7093 (N_7093,N_6999,N_6895);
nand U7094 (N_7094,N_6878,N_6803);
or U7095 (N_7095,N_6939,N_6813);
and U7096 (N_7096,N_6919,N_6801);
or U7097 (N_7097,N_6956,N_6825);
or U7098 (N_7098,N_6949,N_6846);
xor U7099 (N_7099,N_6860,N_6923);
xor U7100 (N_7100,N_6917,N_6943);
nand U7101 (N_7101,N_6851,N_6889);
and U7102 (N_7102,N_6920,N_6995);
and U7103 (N_7103,N_6891,N_6999);
xnor U7104 (N_7104,N_6915,N_6860);
and U7105 (N_7105,N_6978,N_6835);
or U7106 (N_7106,N_6999,N_6844);
nand U7107 (N_7107,N_6919,N_6835);
nor U7108 (N_7108,N_6992,N_6924);
nor U7109 (N_7109,N_6818,N_6807);
xnor U7110 (N_7110,N_6927,N_6903);
nand U7111 (N_7111,N_6931,N_6823);
nor U7112 (N_7112,N_6849,N_6977);
xnor U7113 (N_7113,N_6873,N_6883);
nand U7114 (N_7114,N_6888,N_6846);
and U7115 (N_7115,N_6833,N_6828);
nand U7116 (N_7116,N_6843,N_6860);
xor U7117 (N_7117,N_6852,N_6805);
nor U7118 (N_7118,N_6845,N_6800);
nor U7119 (N_7119,N_6820,N_6818);
nand U7120 (N_7120,N_6919,N_6819);
and U7121 (N_7121,N_6920,N_6909);
xnor U7122 (N_7122,N_6905,N_6817);
or U7123 (N_7123,N_6917,N_6930);
nand U7124 (N_7124,N_6822,N_6835);
xor U7125 (N_7125,N_6821,N_6916);
nand U7126 (N_7126,N_6851,N_6932);
or U7127 (N_7127,N_6923,N_6904);
nor U7128 (N_7128,N_6864,N_6969);
and U7129 (N_7129,N_6836,N_6853);
and U7130 (N_7130,N_6958,N_6870);
and U7131 (N_7131,N_6820,N_6898);
nor U7132 (N_7132,N_6918,N_6930);
nor U7133 (N_7133,N_6942,N_6868);
and U7134 (N_7134,N_6854,N_6899);
nor U7135 (N_7135,N_6945,N_6894);
xnor U7136 (N_7136,N_6915,N_6851);
or U7137 (N_7137,N_6934,N_6810);
nor U7138 (N_7138,N_6898,N_6936);
and U7139 (N_7139,N_6916,N_6819);
or U7140 (N_7140,N_6899,N_6867);
and U7141 (N_7141,N_6865,N_6995);
nand U7142 (N_7142,N_6979,N_6834);
xor U7143 (N_7143,N_6986,N_6924);
xor U7144 (N_7144,N_6858,N_6826);
and U7145 (N_7145,N_6848,N_6966);
nor U7146 (N_7146,N_6990,N_6811);
nor U7147 (N_7147,N_6952,N_6881);
or U7148 (N_7148,N_6911,N_6898);
or U7149 (N_7149,N_6942,N_6844);
nand U7150 (N_7150,N_6849,N_6808);
nand U7151 (N_7151,N_6814,N_6823);
and U7152 (N_7152,N_6923,N_6852);
and U7153 (N_7153,N_6907,N_6800);
and U7154 (N_7154,N_6890,N_6904);
nand U7155 (N_7155,N_6931,N_6989);
or U7156 (N_7156,N_6999,N_6942);
and U7157 (N_7157,N_6963,N_6818);
nor U7158 (N_7158,N_6969,N_6998);
nor U7159 (N_7159,N_6924,N_6817);
or U7160 (N_7160,N_6845,N_6851);
or U7161 (N_7161,N_6974,N_6942);
xnor U7162 (N_7162,N_6958,N_6834);
and U7163 (N_7163,N_6871,N_6918);
nor U7164 (N_7164,N_6934,N_6809);
nor U7165 (N_7165,N_6861,N_6830);
or U7166 (N_7166,N_6896,N_6970);
xnor U7167 (N_7167,N_6831,N_6991);
or U7168 (N_7168,N_6986,N_6965);
xnor U7169 (N_7169,N_6937,N_6920);
nor U7170 (N_7170,N_6930,N_6861);
and U7171 (N_7171,N_6915,N_6954);
nor U7172 (N_7172,N_6904,N_6913);
or U7173 (N_7173,N_6915,N_6974);
and U7174 (N_7174,N_6942,N_6896);
or U7175 (N_7175,N_6980,N_6938);
or U7176 (N_7176,N_6839,N_6954);
and U7177 (N_7177,N_6885,N_6848);
or U7178 (N_7178,N_6836,N_6861);
and U7179 (N_7179,N_6879,N_6932);
and U7180 (N_7180,N_6887,N_6966);
nor U7181 (N_7181,N_6991,N_6844);
or U7182 (N_7182,N_6933,N_6944);
or U7183 (N_7183,N_6815,N_6810);
and U7184 (N_7184,N_6876,N_6858);
or U7185 (N_7185,N_6959,N_6867);
xnor U7186 (N_7186,N_6945,N_6905);
xnor U7187 (N_7187,N_6986,N_6829);
or U7188 (N_7188,N_6874,N_6840);
nor U7189 (N_7189,N_6921,N_6857);
and U7190 (N_7190,N_6898,N_6847);
and U7191 (N_7191,N_6952,N_6969);
nand U7192 (N_7192,N_6967,N_6885);
nand U7193 (N_7193,N_6885,N_6897);
or U7194 (N_7194,N_6888,N_6841);
nor U7195 (N_7195,N_6857,N_6914);
or U7196 (N_7196,N_6973,N_6835);
or U7197 (N_7197,N_6928,N_6814);
and U7198 (N_7198,N_6819,N_6932);
nor U7199 (N_7199,N_6957,N_6851);
nand U7200 (N_7200,N_7038,N_7099);
xnor U7201 (N_7201,N_7134,N_7132);
xor U7202 (N_7202,N_7000,N_7156);
nand U7203 (N_7203,N_7009,N_7042);
or U7204 (N_7204,N_7128,N_7158);
xor U7205 (N_7205,N_7104,N_7024);
and U7206 (N_7206,N_7111,N_7192);
nand U7207 (N_7207,N_7143,N_7157);
xor U7208 (N_7208,N_7007,N_7141);
and U7209 (N_7209,N_7089,N_7135);
or U7210 (N_7210,N_7129,N_7116);
and U7211 (N_7211,N_7119,N_7100);
and U7212 (N_7212,N_7062,N_7076);
xnor U7213 (N_7213,N_7010,N_7101);
nor U7214 (N_7214,N_7117,N_7155);
and U7215 (N_7215,N_7088,N_7166);
xnor U7216 (N_7216,N_7035,N_7096);
nor U7217 (N_7217,N_7081,N_7118);
xnor U7218 (N_7218,N_7018,N_7026);
or U7219 (N_7219,N_7110,N_7025);
and U7220 (N_7220,N_7053,N_7122);
nand U7221 (N_7221,N_7151,N_7040);
nor U7222 (N_7222,N_7072,N_7093);
and U7223 (N_7223,N_7033,N_7073);
or U7224 (N_7224,N_7184,N_7123);
nand U7225 (N_7225,N_7080,N_7049);
and U7226 (N_7226,N_7127,N_7070);
nor U7227 (N_7227,N_7142,N_7091);
xor U7228 (N_7228,N_7055,N_7161);
nor U7229 (N_7229,N_7021,N_7162);
nor U7230 (N_7230,N_7092,N_7068);
or U7231 (N_7231,N_7121,N_7163);
nor U7232 (N_7232,N_7060,N_7150);
nor U7233 (N_7233,N_7034,N_7175);
or U7234 (N_7234,N_7145,N_7082);
xor U7235 (N_7235,N_7047,N_7176);
and U7236 (N_7236,N_7011,N_7057);
or U7237 (N_7237,N_7044,N_7144);
nor U7238 (N_7238,N_7027,N_7036);
and U7239 (N_7239,N_7168,N_7196);
and U7240 (N_7240,N_7147,N_7125);
xnor U7241 (N_7241,N_7001,N_7051);
nand U7242 (N_7242,N_7113,N_7194);
and U7243 (N_7243,N_7006,N_7002);
and U7244 (N_7244,N_7066,N_7191);
xnor U7245 (N_7245,N_7065,N_7085);
or U7246 (N_7246,N_7005,N_7064);
or U7247 (N_7247,N_7102,N_7003);
nand U7248 (N_7248,N_7138,N_7094);
and U7249 (N_7249,N_7059,N_7029);
or U7250 (N_7250,N_7074,N_7189);
or U7251 (N_7251,N_7130,N_7137);
nor U7252 (N_7252,N_7139,N_7187);
nand U7253 (N_7253,N_7045,N_7146);
nor U7254 (N_7254,N_7061,N_7133);
nor U7255 (N_7255,N_7182,N_7058);
or U7256 (N_7256,N_7171,N_7179);
xor U7257 (N_7257,N_7183,N_7030);
xor U7258 (N_7258,N_7106,N_7077);
and U7259 (N_7259,N_7014,N_7109);
and U7260 (N_7260,N_7165,N_7012);
and U7261 (N_7261,N_7195,N_7015);
nand U7262 (N_7262,N_7004,N_7185);
and U7263 (N_7263,N_7050,N_7079);
nand U7264 (N_7264,N_7198,N_7039);
and U7265 (N_7265,N_7098,N_7063);
or U7266 (N_7266,N_7032,N_7178);
xnor U7267 (N_7267,N_7078,N_7105);
nor U7268 (N_7268,N_7186,N_7197);
nand U7269 (N_7269,N_7052,N_7019);
and U7270 (N_7270,N_7124,N_7028);
nand U7271 (N_7271,N_7152,N_7086);
xnor U7272 (N_7272,N_7154,N_7188);
nand U7273 (N_7273,N_7159,N_7108);
and U7274 (N_7274,N_7084,N_7020);
xnor U7275 (N_7275,N_7016,N_7090);
nand U7276 (N_7276,N_7172,N_7041);
xor U7277 (N_7277,N_7180,N_7170);
and U7278 (N_7278,N_7103,N_7031);
or U7279 (N_7279,N_7114,N_7131);
and U7280 (N_7280,N_7174,N_7173);
and U7281 (N_7281,N_7097,N_7177);
and U7282 (N_7282,N_7013,N_7056);
and U7283 (N_7283,N_7022,N_7160);
nand U7284 (N_7284,N_7140,N_7164);
xor U7285 (N_7285,N_7069,N_7136);
or U7286 (N_7286,N_7120,N_7148);
and U7287 (N_7287,N_7199,N_7153);
xor U7288 (N_7288,N_7046,N_7037);
xor U7289 (N_7289,N_7054,N_7043);
nor U7290 (N_7290,N_7112,N_7087);
nand U7291 (N_7291,N_7017,N_7167);
and U7292 (N_7292,N_7071,N_7126);
and U7293 (N_7293,N_7107,N_7008);
or U7294 (N_7294,N_7067,N_7095);
or U7295 (N_7295,N_7181,N_7115);
nand U7296 (N_7296,N_7149,N_7169);
and U7297 (N_7297,N_7190,N_7083);
and U7298 (N_7298,N_7193,N_7075);
and U7299 (N_7299,N_7048,N_7023);
nand U7300 (N_7300,N_7034,N_7141);
nor U7301 (N_7301,N_7062,N_7140);
and U7302 (N_7302,N_7098,N_7009);
nand U7303 (N_7303,N_7186,N_7092);
nor U7304 (N_7304,N_7184,N_7034);
nor U7305 (N_7305,N_7175,N_7182);
nor U7306 (N_7306,N_7056,N_7026);
nand U7307 (N_7307,N_7044,N_7001);
xor U7308 (N_7308,N_7053,N_7003);
and U7309 (N_7309,N_7101,N_7025);
xnor U7310 (N_7310,N_7100,N_7037);
or U7311 (N_7311,N_7056,N_7060);
xnor U7312 (N_7312,N_7166,N_7123);
nand U7313 (N_7313,N_7106,N_7165);
nand U7314 (N_7314,N_7187,N_7055);
or U7315 (N_7315,N_7135,N_7199);
xnor U7316 (N_7316,N_7138,N_7122);
and U7317 (N_7317,N_7110,N_7018);
nand U7318 (N_7318,N_7150,N_7052);
and U7319 (N_7319,N_7169,N_7171);
nor U7320 (N_7320,N_7154,N_7064);
nand U7321 (N_7321,N_7095,N_7169);
xor U7322 (N_7322,N_7184,N_7145);
nor U7323 (N_7323,N_7109,N_7053);
nor U7324 (N_7324,N_7087,N_7007);
or U7325 (N_7325,N_7019,N_7154);
nor U7326 (N_7326,N_7168,N_7144);
xnor U7327 (N_7327,N_7145,N_7152);
and U7328 (N_7328,N_7106,N_7047);
xor U7329 (N_7329,N_7186,N_7072);
nand U7330 (N_7330,N_7037,N_7143);
or U7331 (N_7331,N_7158,N_7104);
and U7332 (N_7332,N_7053,N_7001);
nand U7333 (N_7333,N_7180,N_7126);
nand U7334 (N_7334,N_7005,N_7053);
nand U7335 (N_7335,N_7165,N_7008);
or U7336 (N_7336,N_7029,N_7045);
xnor U7337 (N_7337,N_7147,N_7046);
xor U7338 (N_7338,N_7004,N_7107);
nor U7339 (N_7339,N_7053,N_7004);
nor U7340 (N_7340,N_7123,N_7189);
xor U7341 (N_7341,N_7046,N_7103);
or U7342 (N_7342,N_7081,N_7106);
and U7343 (N_7343,N_7046,N_7067);
nand U7344 (N_7344,N_7184,N_7106);
xnor U7345 (N_7345,N_7184,N_7156);
nor U7346 (N_7346,N_7181,N_7127);
nand U7347 (N_7347,N_7076,N_7092);
nor U7348 (N_7348,N_7061,N_7096);
and U7349 (N_7349,N_7056,N_7190);
xnor U7350 (N_7350,N_7197,N_7046);
and U7351 (N_7351,N_7000,N_7138);
nand U7352 (N_7352,N_7008,N_7004);
and U7353 (N_7353,N_7002,N_7169);
nand U7354 (N_7354,N_7175,N_7067);
or U7355 (N_7355,N_7198,N_7038);
or U7356 (N_7356,N_7129,N_7135);
xnor U7357 (N_7357,N_7030,N_7186);
nand U7358 (N_7358,N_7136,N_7194);
nand U7359 (N_7359,N_7150,N_7030);
nand U7360 (N_7360,N_7154,N_7010);
nand U7361 (N_7361,N_7145,N_7179);
or U7362 (N_7362,N_7111,N_7185);
nor U7363 (N_7363,N_7073,N_7109);
nand U7364 (N_7364,N_7168,N_7042);
or U7365 (N_7365,N_7132,N_7136);
or U7366 (N_7366,N_7199,N_7059);
and U7367 (N_7367,N_7002,N_7148);
nand U7368 (N_7368,N_7104,N_7108);
and U7369 (N_7369,N_7045,N_7122);
nand U7370 (N_7370,N_7095,N_7073);
or U7371 (N_7371,N_7196,N_7052);
nor U7372 (N_7372,N_7099,N_7152);
and U7373 (N_7373,N_7176,N_7190);
xnor U7374 (N_7374,N_7030,N_7064);
nor U7375 (N_7375,N_7032,N_7153);
nand U7376 (N_7376,N_7060,N_7091);
xor U7377 (N_7377,N_7089,N_7005);
and U7378 (N_7378,N_7034,N_7100);
xor U7379 (N_7379,N_7131,N_7127);
and U7380 (N_7380,N_7188,N_7177);
nor U7381 (N_7381,N_7143,N_7119);
or U7382 (N_7382,N_7107,N_7047);
nand U7383 (N_7383,N_7042,N_7119);
nor U7384 (N_7384,N_7008,N_7122);
xnor U7385 (N_7385,N_7023,N_7192);
and U7386 (N_7386,N_7085,N_7196);
nor U7387 (N_7387,N_7188,N_7004);
nand U7388 (N_7388,N_7076,N_7153);
nor U7389 (N_7389,N_7161,N_7162);
and U7390 (N_7390,N_7089,N_7083);
xor U7391 (N_7391,N_7151,N_7028);
or U7392 (N_7392,N_7051,N_7072);
nand U7393 (N_7393,N_7086,N_7005);
nand U7394 (N_7394,N_7040,N_7140);
xor U7395 (N_7395,N_7197,N_7110);
nor U7396 (N_7396,N_7125,N_7155);
or U7397 (N_7397,N_7064,N_7070);
or U7398 (N_7398,N_7190,N_7039);
nor U7399 (N_7399,N_7032,N_7071);
xnor U7400 (N_7400,N_7326,N_7250);
nor U7401 (N_7401,N_7206,N_7272);
xor U7402 (N_7402,N_7372,N_7279);
and U7403 (N_7403,N_7374,N_7258);
or U7404 (N_7404,N_7382,N_7362);
xnor U7405 (N_7405,N_7331,N_7240);
nand U7406 (N_7406,N_7268,N_7229);
or U7407 (N_7407,N_7398,N_7364);
and U7408 (N_7408,N_7275,N_7211);
nor U7409 (N_7409,N_7249,N_7218);
xor U7410 (N_7410,N_7308,N_7378);
nor U7411 (N_7411,N_7292,N_7337);
nor U7412 (N_7412,N_7306,N_7304);
and U7413 (N_7413,N_7271,N_7365);
and U7414 (N_7414,N_7359,N_7289);
or U7415 (N_7415,N_7269,N_7393);
nor U7416 (N_7416,N_7366,N_7300);
and U7417 (N_7417,N_7252,N_7223);
xor U7418 (N_7418,N_7373,N_7236);
xnor U7419 (N_7419,N_7287,N_7233);
nand U7420 (N_7420,N_7286,N_7376);
xor U7421 (N_7421,N_7384,N_7387);
nand U7422 (N_7422,N_7343,N_7358);
nor U7423 (N_7423,N_7309,N_7338);
and U7424 (N_7424,N_7330,N_7302);
and U7425 (N_7425,N_7231,N_7251);
nor U7426 (N_7426,N_7277,N_7392);
nand U7427 (N_7427,N_7363,N_7237);
nor U7428 (N_7428,N_7307,N_7242);
and U7429 (N_7429,N_7342,N_7361);
nand U7430 (N_7430,N_7284,N_7349);
and U7431 (N_7431,N_7369,N_7347);
nor U7432 (N_7432,N_7296,N_7243);
nor U7433 (N_7433,N_7260,N_7219);
nor U7434 (N_7434,N_7346,N_7340);
or U7435 (N_7435,N_7247,N_7210);
xor U7436 (N_7436,N_7221,N_7238);
nor U7437 (N_7437,N_7323,N_7344);
xnor U7438 (N_7438,N_7246,N_7266);
or U7439 (N_7439,N_7394,N_7334);
or U7440 (N_7440,N_7263,N_7336);
nor U7441 (N_7441,N_7214,N_7375);
nand U7442 (N_7442,N_7341,N_7348);
and U7443 (N_7443,N_7322,N_7383);
or U7444 (N_7444,N_7248,N_7391);
and U7445 (N_7445,N_7314,N_7215);
xnor U7446 (N_7446,N_7311,N_7312);
xnor U7447 (N_7447,N_7294,N_7316);
nand U7448 (N_7448,N_7253,N_7385);
xor U7449 (N_7449,N_7230,N_7379);
nand U7450 (N_7450,N_7293,N_7232);
or U7451 (N_7451,N_7209,N_7282);
or U7452 (N_7452,N_7389,N_7318);
nor U7453 (N_7453,N_7224,N_7390);
and U7454 (N_7454,N_7357,N_7396);
or U7455 (N_7455,N_7368,N_7327);
and U7456 (N_7456,N_7239,N_7261);
and U7457 (N_7457,N_7299,N_7255);
xor U7458 (N_7458,N_7280,N_7370);
xnor U7459 (N_7459,N_7297,N_7328);
or U7460 (N_7460,N_7360,N_7320);
or U7461 (N_7461,N_7332,N_7371);
or U7462 (N_7462,N_7202,N_7386);
or U7463 (N_7463,N_7291,N_7228);
nand U7464 (N_7464,N_7213,N_7352);
xnor U7465 (N_7465,N_7208,N_7325);
xnor U7466 (N_7466,N_7305,N_7257);
xnor U7467 (N_7467,N_7259,N_7333);
and U7468 (N_7468,N_7301,N_7273);
nand U7469 (N_7469,N_7354,N_7205);
or U7470 (N_7470,N_7399,N_7234);
nand U7471 (N_7471,N_7350,N_7329);
xor U7472 (N_7472,N_7324,N_7315);
xnor U7473 (N_7473,N_7212,N_7339);
and U7474 (N_7474,N_7226,N_7265);
and U7475 (N_7475,N_7283,N_7235);
or U7476 (N_7476,N_7380,N_7298);
nor U7477 (N_7477,N_7245,N_7256);
or U7478 (N_7478,N_7270,N_7225);
or U7479 (N_7479,N_7274,N_7303);
and U7480 (N_7480,N_7313,N_7317);
and U7481 (N_7481,N_7222,N_7321);
and U7482 (N_7482,N_7345,N_7377);
nand U7483 (N_7483,N_7281,N_7288);
xor U7484 (N_7484,N_7355,N_7220);
xnor U7485 (N_7485,N_7356,N_7278);
nor U7486 (N_7486,N_7227,N_7267);
nor U7487 (N_7487,N_7241,N_7264);
nor U7488 (N_7488,N_7388,N_7254);
nand U7489 (N_7489,N_7262,N_7203);
nor U7490 (N_7490,N_7353,N_7319);
nand U7491 (N_7491,N_7276,N_7381);
nor U7492 (N_7492,N_7207,N_7351);
and U7493 (N_7493,N_7204,N_7285);
nand U7494 (N_7494,N_7244,N_7216);
nor U7495 (N_7495,N_7201,N_7335);
nand U7496 (N_7496,N_7290,N_7295);
or U7497 (N_7497,N_7217,N_7310);
xor U7498 (N_7498,N_7200,N_7367);
or U7499 (N_7499,N_7395,N_7397);
nand U7500 (N_7500,N_7257,N_7217);
or U7501 (N_7501,N_7398,N_7215);
nand U7502 (N_7502,N_7305,N_7229);
nand U7503 (N_7503,N_7315,N_7339);
nor U7504 (N_7504,N_7275,N_7373);
and U7505 (N_7505,N_7375,N_7251);
nor U7506 (N_7506,N_7248,N_7219);
nor U7507 (N_7507,N_7315,N_7383);
nor U7508 (N_7508,N_7321,N_7383);
nor U7509 (N_7509,N_7220,N_7324);
nand U7510 (N_7510,N_7376,N_7387);
xor U7511 (N_7511,N_7275,N_7397);
nand U7512 (N_7512,N_7300,N_7269);
nand U7513 (N_7513,N_7297,N_7291);
and U7514 (N_7514,N_7339,N_7205);
and U7515 (N_7515,N_7368,N_7296);
nor U7516 (N_7516,N_7343,N_7366);
or U7517 (N_7517,N_7354,N_7207);
xnor U7518 (N_7518,N_7301,N_7362);
nand U7519 (N_7519,N_7210,N_7252);
nor U7520 (N_7520,N_7239,N_7281);
and U7521 (N_7521,N_7377,N_7327);
or U7522 (N_7522,N_7334,N_7281);
nor U7523 (N_7523,N_7235,N_7248);
or U7524 (N_7524,N_7351,N_7249);
xor U7525 (N_7525,N_7311,N_7230);
nand U7526 (N_7526,N_7321,N_7231);
nor U7527 (N_7527,N_7397,N_7369);
xor U7528 (N_7528,N_7313,N_7247);
or U7529 (N_7529,N_7376,N_7205);
nand U7530 (N_7530,N_7301,N_7244);
nand U7531 (N_7531,N_7277,N_7357);
nand U7532 (N_7532,N_7233,N_7308);
and U7533 (N_7533,N_7344,N_7263);
xnor U7534 (N_7534,N_7348,N_7312);
xor U7535 (N_7535,N_7287,N_7217);
or U7536 (N_7536,N_7210,N_7309);
and U7537 (N_7537,N_7361,N_7264);
nand U7538 (N_7538,N_7311,N_7385);
xor U7539 (N_7539,N_7225,N_7375);
nand U7540 (N_7540,N_7310,N_7342);
nand U7541 (N_7541,N_7373,N_7330);
or U7542 (N_7542,N_7275,N_7276);
nor U7543 (N_7543,N_7360,N_7273);
nor U7544 (N_7544,N_7284,N_7321);
xnor U7545 (N_7545,N_7207,N_7230);
nor U7546 (N_7546,N_7329,N_7304);
or U7547 (N_7547,N_7295,N_7396);
and U7548 (N_7548,N_7275,N_7225);
or U7549 (N_7549,N_7237,N_7342);
or U7550 (N_7550,N_7247,N_7357);
xnor U7551 (N_7551,N_7320,N_7210);
nand U7552 (N_7552,N_7238,N_7287);
or U7553 (N_7553,N_7260,N_7379);
nor U7554 (N_7554,N_7215,N_7328);
or U7555 (N_7555,N_7346,N_7260);
and U7556 (N_7556,N_7362,N_7280);
nand U7557 (N_7557,N_7242,N_7391);
xor U7558 (N_7558,N_7213,N_7301);
nand U7559 (N_7559,N_7397,N_7206);
xor U7560 (N_7560,N_7242,N_7283);
nor U7561 (N_7561,N_7223,N_7326);
nand U7562 (N_7562,N_7261,N_7325);
and U7563 (N_7563,N_7389,N_7225);
nor U7564 (N_7564,N_7269,N_7383);
xor U7565 (N_7565,N_7290,N_7388);
or U7566 (N_7566,N_7389,N_7321);
nor U7567 (N_7567,N_7250,N_7205);
nor U7568 (N_7568,N_7234,N_7357);
or U7569 (N_7569,N_7341,N_7367);
and U7570 (N_7570,N_7271,N_7358);
or U7571 (N_7571,N_7227,N_7259);
or U7572 (N_7572,N_7388,N_7280);
and U7573 (N_7573,N_7260,N_7256);
or U7574 (N_7574,N_7221,N_7317);
xor U7575 (N_7575,N_7314,N_7312);
nand U7576 (N_7576,N_7288,N_7373);
and U7577 (N_7577,N_7301,N_7393);
nand U7578 (N_7578,N_7283,N_7267);
or U7579 (N_7579,N_7201,N_7279);
or U7580 (N_7580,N_7247,N_7320);
and U7581 (N_7581,N_7255,N_7249);
or U7582 (N_7582,N_7229,N_7228);
nand U7583 (N_7583,N_7304,N_7315);
nor U7584 (N_7584,N_7241,N_7343);
nand U7585 (N_7585,N_7212,N_7352);
and U7586 (N_7586,N_7338,N_7251);
nor U7587 (N_7587,N_7220,N_7363);
xnor U7588 (N_7588,N_7258,N_7245);
xnor U7589 (N_7589,N_7352,N_7344);
nor U7590 (N_7590,N_7203,N_7215);
nor U7591 (N_7591,N_7382,N_7302);
nor U7592 (N_7592,N_7283,N_7389);
nand U7593 (N_7593,N_7354,N_7211);
nor U7594 (N_7594,N_7210,N_7363);
nor U7595 (N_7595,N_7297,N_7390);
xor U7596 (N_7596,N_7399,N_7385);
xor U7597 (N_7597,N_7317,N_7304);
nand U7598 (N_7598,N_7339,N_7372);
or U7599 (N_7599,N_7287,N_7262);
nor U7600 (N_7600,N_7564,N_7551);
nand U7601 (N_7601,N_7405,N_7486);
nand U7602 (N_7602,N_7423,N_7567);
xor U7603 (N_7603,N_7541,N_7442);
or U7604 (N_7604,N_7538,N_7488);
or U7605 (N_7605,N_7414,N_7419);
xnor U7606 (N_7606,N_7556,N_7415);
nand U7607 (N_7607,N_7444,N_7484);
nor U7608 (N_7608,N_7420,N_7437);
xor U7609 (N_7609,N_7540,N_7451);
nor U7610 (N_7610,N_7453,N_7510);
or U7611 (N_7611,N_7557,N_7574);
or U7612 (N_7612,N_7578,N_7464);
xnor U7613 (N_7613,N_7555,N_7589);
nand U7614 (N_7614,N_7591,N_7468);
or U7615 (N_7615,N_7482,N_7568);
nor U7616 (N_7616,N_7470,N_7410);
nor U7617 (N_7617,N_7594,N_7586);
nand U7618 (N_7618,N_7448,N_7479);
nand U7619 (N_7619,N_7549,N_7471);
and U7620 (N_7620,N_7490,N_7435);
and U7621 (N_7621,N_7411,N_7558);
and U7622 (N_7622,N_7472,N_7565);
xnor U7623 (N_7623,N_7450,N_7544);
xor U7624 (N_7624,N_7581,N_7501);
or U7625 (N_7625,N_7449,N_7548);
or U7626 (N_7626,N_7559,N_7563);
and U7627 (N_7627,N_7452,N_7493);
xor U7628 (N_7628,N_7598,N_7439);
and U7629 (N_7629,N_7462,N_7480);
and U7630 (N_7630,N_7447,N_7489);
or U7631 (N_7631,N_7536,N_7456);
nand U7632 (N_7632,N_7432,N_7426);
nand U7633 (N_7633,N_7441,N_7575);
nand U7634 (N_7634,N_7593,N_7529);
and U7635 (N_7635,N_7408,N_7505);
nor U7636 (N_7636,N_7511,N_7531);
xnor U7637 (N_7637,N_7539,N_7545);
nand U7638 (N_7638,N_7503,N_7403);
or U7639 (N_7639,N_7569,N_7552);
or U7640 (N_7640,N_7517,N_7576);
nor U7641 (N_7641,N_7431,N_7495);
nand U7642 (N_7642,N_7504,N_7446);
nor U7643 (N_7643,N_7436,N_7553);
and U7644 (N_7644,N_7583,N_7460);
or U7645 (N_7645,N_7445,N_7554);
or U7646 (N_7646,N_7580,N_7412);
or U7647 (N_7647,N_7418,N_7469);
and U7648 (N_7648,N_7582,N_7595);
nor U7649 (N_7649,N_7430,N_7509);
xor U7650 (N_7650,N_7428,N_7465);
or U7651 (N_7651,N_7535,N_7526);
and U7652 (N_7652,N_7476,N_7457);
nand U7653 (N_7653,N_7562,N_7425);
or U7654 (N_7654,N_7587,N_7400);
and U7655 (N_7655,N_7443,N_7494);
xor U7656 (N_7656,N_7566,N_7487);
or U7657 (N_7657,N_7596,N_7475);
xnor U7658 (N_7658,N_7514,N_7550);
nand U7659 (N_7659,N_7599,N_7427);
nand U7660 (N_7660,N_7516,N_7491);
nor U7661 (N_7661,N_7467,N_7592);
nand U7662 (N_7662,N_7584,N_7473);
nor U7663 (N_7663,N_7597,N_7530);
nor U7664 (N_7664,N_7571,N_7496);
or U7665 (N_7665,N_7527,N_7458);
and U7666 (N_7666,N_7542,N_7506);
and U7667 (N_7667,N_7406,N_7533);
and U7668 (N_7668,N_7474,N_7513);
or U7669 (N_7669,N_7417,N_7477);
and U7670 (N_7670,N_7466,N_7485);
and U7671 (N_7671,N_7577,N_7507);
and U7672 (N_7672,N_7537,N_7404);
or U7673 (N_7673,N_7519,N_7573);
nand U7674 (N_7674,N_7433,N_7434);
xnor U7675 (N_7675,N_7528,N_7534);
xor U7676 (N_7676,N_7520,N_7518);
nor U7677 (N_7677,N_7498,N_7463);
and U7678 (N_7678,N_7572,N_7407);
xnor U7679 (N_7679,N_7522,N_7585);
nand U7680 (N_7680,N_7579,N_7461);
xnor U7681 (N_7681,N_7515,N_7416);
nand U7682 (N_7682,N_7547,N_7523);
and U7683 (N_7683,N_7512,N_7402);
nor U7684 (N_7684,N_7401,N_7409);
and U7685 (N_7685,N_7459,N_7543);
nor U7686 (N_7686,N_7588,N_7413);
or U7687 (N_7687,N_7478,N_7422);
and U7688 (N_7688,N_7546,N_7561);
xor U7689 (N_7689,N_7590,N_7454);
xnor U7690 (N_7690,N_7532,N_7525);
xor U7691 (N_7691,N_7502,N_7492);
nand U7692 (N_7692,N_7570,N_7421);
xor U7693 (N_7693,N_7424,N_7481);
and U7694 (N_7694,N_7560,N_7497);
nor U7695 (N_7695,N_7440,N_7521);
nor U7696 (N_7696,N_7455,N_7500);
or U7697 (N_7697,N_7499,N_7438);
nor U7698 (N_7698,N_7508,N_7483);
nor U7699 (N_7699,N_7429,N_7524);
and U7700 (N_7700,N_7443,N_7463);
and U7701 (N_7701,N_7537,N_7512);
and U7702 (N_7702,N_7575,N_7496);
nand U7703 (N_7703,N_7451,N_7479);
nand U7704 (N_7704,N_7462,N_7538);
nor U7705 (N_7705,N_7438,N_7464);
xor U7706 (N_7706,N_7492,N_7488);
xor U7707 (N_7707,N_7542,N_7492);
nand U7708 (N_7708,N_7577,N_7573);
xor U7709 (N_7709,N_7458,N_7426);
xor U7710 (N_7710,N_7435,N_7479);
and U7711 (N_7711,N_7495,N_7521);
nor U7712 (N_7712,N_7418,N_7571);
or U7713 (N_7713,N_7405,N_7573);
xnor U7714 (N_7714,N_7405,N_7460);
and U7715 (N_7715,N_7515,N_7546);
nand U7716 (N_7716,N_7500,N_7496);
xnor U7717 (N_7717,N_7535,N_7471);
nand U7718 (N_7718,N_7589,N_7505);
nand U7719 (N_7719,N_7573,N_7522);
nor U7720 (N_7720,N_7555,N_7590);
and U7721 (N_7721,N_7463,N_7436);
nand U7722 (N_7722,N_7560,N_7593);
and U7723 (N_7723,N_7467,N_7452);
or U7724 (N_7724,N_7463,N_7496);
or U7725 (N_7725,N_7429,N_7550);
and U7726 (N_7726,N_7563,N_7412);
xnor U7727 (N_7727,N_7411,N_7592);
nor U7728 (N_7728,N_7487,N_7423);
xor U7729 (N_7729,N_7438,N_7542);
nor U7730 (N_7730,N_7416,N_7485);
nand U7731 (N_7731,N_7510,N_7598);
and U7732 (N_7732,N_7595,N_7519);
nand U7733 (N_7733,N_7578,N_7456);
nand U7734 (N_7734,N_7584,N_7452);
xnor U7735 (N_7735,N_7508,N_7520);
xnor U7736 (N_7736,N_7445,N_7579);
or U7737 (N_7737,N_7458,N_7555);
nand U7738 (N_7738,N_7545,N_7585);
xnor U7739 (N_7739,N_7445,N_7525);
nand U7740 (N_7740,N_7421,N_7459);
and U7741 (N_7741,N_7496,N_7486);
nand U7742 (N_7742,N_7513,N_7429);
nor U7743 (N_7743,N_7499,N_7437);
nand U7744 (N_7744,N_7581,N_7465);
or U7745 (N_7745,N_7598,N_7442);
nor U7746 (N_7746,N_7574,N_7445);
nand U7747 (N_7747,N_7529,N_7422);
xnor U7748 (N_7748,N_7510,N_7526);
xor U7749 (N_7749,N_7439,N_7419);
nor U7750 (N_7750,N_7439,N_7567);
xor U7751 (N_7751,N_7438,N_7424);
or U7752 (N_7752,N_7477,N_7438);
and U7753 (N_7753,N_7563,N_7523);
nor U7754 (N_7754,N_7579,N_7549);
xor U7755 (N_7755,N_7539,N_7489);
nand U7756 (N_7756,N_7408,N_7403);
xnor U7757 (N_7757,N_7564,N_7483);
nor U7758 (N_7758,N_7417,N_7499);
or U7759 (N_7759,N_7486,N_7538);
and U7760 (N_7760,N_7433,N_7559);
nor U7761 (N_7761,N_7466,N_7578);
nor U7762 (N_7762,N_7593,N_7464);
nand U7763 (N_7763,N_7505,N_7460);
xor U7764 (N_7764,N_7450,N_7440);
and U7765 (N_7765,N_7574,N_7469);
nor U7766 (N_7766,N_7470,N_7527);
or U7767 (N_7767,N_7544,N_7461);
or U7768 (N_7768,N_7529,N_7453);
and U7769 (N_7769,N_7441,N_7422);
or U7770 (N_7770,N_7489,N_7418);
nand U7771 (N_7771,N_7577,N_7440);
nor U7772 (N_7772,N_7413,N_7430);
nor U7773 (N_7773,N_7449,N_7490);
and U7774 (N_7774,N_7491,N_7457);
and U7775 (N_7775,N_7470,N_7406);
and U7776 (N_7776,N_7575,N_7541);
nand U7777 (N_7777,N_7472,N_7542);
nor U7778 (N_7778,N_7471,N_7488);
xnor U7779 (N_7779,N_7464,N_7400);
and U7780 (N_7780,N_7560,N_7402);
and U7781 (N_7781,N_7525,N_7517);
nand U7782 (N_7782,N_7542,N_7574);
xnor U7783 (N_7783,N_7557,N_7414);
xor U7784 (N_7784,N_7558,N_7476);
nor U7785 (N_7785,N_7483,N_7514);
nand U7786 (N_7786,N_7507,N_7469);
and U7787 (N_7787,N_7486,N_7462);
nand U7788 (N_7788,N_7522,N_7434);
nand U7789 (N_7789,N_7502,N_7558);
nor U7790 (N_7790,N_7496,N_7483);
nor U7791 (N_7791,N_7539,N_7479);
xnor U7792 (N_7792,N_7599,N_7487);
nor U7793 (N_7793,N_7535,N_7512);
or U7794 (N_7794,N_7430,N_7585);
xnor U7795 (N_7795,N_7419,N_7598);
xor U7796 (N_7796,N_7545,N_7575);
and U7797 (N_7797,N_7402,N_7510);
nand U7798 (N_7798,N_7578,N_7482);
nand U7799 (N_7799,N_7470,N_7493);
nand U7800 (N_7800,N_7664,N_7763);
nand U7801 (N_7801,N_7651,N_7733);
or U7802 (N_7802,N_7615,N_7633);
or U7803 (N_7803,N_7775,N_7748);
xor U7804 (N_7804,N_7739,N_7690);
or U7805 (N_7805,N_7602,N_7776);
or U7806 (N_7806,N_7650,N_7732);
and U7807 (N_7807,N_7754,N_7620);
nand U7808 (N_7808,N_7736,N_7625);
or U7809 (N_7809,N_7706,N_7710);
or U7810 (N_7810,N_7790,N_7792);
xnor U7811 (N_7811,N_7670,N_7671);
nor U7812 (N_7812,N_7668,N_7685);
xnor U7813 (N_7813,N_7719,N_7647);
and U7814 (N_7814,N_7663,N_7661);
nand U7815 (N_7815,N_7683,N_7774);
nand U7816 (N_7816,N_7642,N_7798);
nand U7817 (N_7817,N_7780,N_7743);
or U7818 (N_7818,N_7606,N_7695);
and U7819 (N_7819,N_7722,N_7746);
or U7820 (N_7820,N_7692,N_7762);
and U7821 (N_7821,N_7702,N_7645);
nor U7822 (N_7822,N_7600,N_7669);
nand U7823 (N_7823,N_7751,N_7704);
xor U7824 (N_7824,N_7644,N_7788);
nand U7825 (N_7825,N_7745,N_7629);
nor U7826 (N_7826,N_7636,N_7787);
or U7827 (N_7827,N_7614,N_7797);
nor U7828 (N_7828,N_7727,N_7653);
xnor U7829 (N_7829,N_7618,N_7741);
nand U7830 (N_7830,N_7665,N_7613);
or U7831 (N_7831,N_7691,N_7696);
or U7832 (N_7832,N_7711,N_7771);
nor U7833 (N_7833,N_7603,N_7682);
xnor U7834 (N_7834,N_7742,N_7799);
and U7835 (N_7835,N_7648,N_7631);
nand U7836 (N_7836,N_7667,N_7655);
and U7837 (N_7837,N_7765,N_7693);
nand U7838 (N_7838,N_7649,N_7755);
or U7839 (N_7839,N_7720,N_7604);
xnor U7840 (N_7840,N_7680,N_7725);
nor U7841 (N_7841,N_7652,N_7697);
nand U7842 (N_7842,N_7657,N_7635);
xnor U7843 (N_7843,N_7786,N_7601);
nor U7844 (N_7844,N_7791,N_7674);
xnor U7845 (N_7845,N_7617,N_7772);
nor U7846 (N_7846,N_7658,N_7611);
nor U7847 (N_7847,N_7634,N_7714);
nand U7848 (N_7848,N_7750,N_7782);
or U7849 (N_7849,N_7639,N_7698);
and U7850 (N_7850,N_7777,N_7764);
nand U7851 (N_7851,N_7627,N_7752);
nand U7852 (N_7852,N_7605,N_7723);
nor U7853 (N_7853,N_7724,N_7638);
and U7854 (N_7854,N_7785,N_7770);
and U7855 (N_7855,N_7758,N_7796);
and U7856 (N_7856,N_7630,N_7646);
xnor U7857 (N_7857,N_7623,N_7659);
xnor U7858 (N_7858,N_7678,N_7660);
and U7859 (N_7859,N_7621,N_7713);
nand U7860 (N_7860,N_7795,N_7749);
xor U7861 (N_7861,N_7728,N_7740);
nor U7862 (N_7862,N_7793,N_7734);
nor U7863 (N_7863,N_7759,N_7640);
or U7864 (N_7864,N_7688,N_7619);
nor U7865 (N_7865,N_7712,N_7654);
xor U7866 (N_7866,N_7672,N_7753);
and U7867 (N_7867,N_7738,N_7773);
and U7868 (N_7868,N_7689,N_7705);
and U7869 (N_7869,N_7694,N_7632);
nor U7870 (N_7870,N_7616,N_7781);
nand U7871 (N_7871,N_7610,N_7700);
nand U7872 (N_7872,N_7612,N_7676);
nor U7873 (N_7873,N_7784,N_7721);
xor U7874 (N_7874,N_7608,N_7756);
nor U7875 (N_7875,N_7744,N_7794);
nand U7876 (N_7876,N_7747,N_7673);
and U7877 (N_7877,N_7628,N_7679);
or U7878 (N_7878,N_7609,N_7662);
or U7879 (N_7879,N_7760,N_7624);
nor U7880 (N_7880,N_7731,N_7715);
xnor U7881 (N_7881,N_7607,N_7737);
and U7882 (N_7882,N_7643,N_7708);
and U7883 (N_7883,N_7709,N_7666);
and U7884 (N_7884,N_7735,N_7789);
nand U7885 (N_7885,N_7717,N_7684);
nand U7886 (N_7886,N_7716,N_7707);
and U7887 (N_7887,N_7637,N_7768);
and U7888 (N_7888,N_7699,N_7718);
nand U7889 (N_7889,N_7703,N_7687);
nand U7890 (N_7890,N_7729,N_7757);
xor U7891 (N_7891,N_7626,N_7778);
nand U7892 (N_7892,N_7766,N_7769);
nor U7893 (N_7893,N_7779,N_7726);
nor U7894 (N_7894,N_7622,N_7681);
xor U7895 (N_7895,N_7783,N_7761);
nor U7896 (N_7896,N_7686,N_7677);
nand U7897 (N_7897,N_7656,N_7701);
xnor U7898 (N_7898,N_7730,N_7767);
nor U7899 (N_7899,N_7641,N_7675);
or U7900 (N_7900,N_7608,N_7778);
nand U7901 (N_7901,N_7756,N_7691);
nor U7902 (N_7902,N_7704,N_7706);
xor U7903 (N_7903,N_7740,N_7630);
nand U7904 (N_7904,N_7608,N_7796);
or U7905 (N_7905,N_7744,N_7644);
or U7906 (N_7906,N_7726,N_7795);
nor U7907 (N_7907,N_7718,N_7705);
nand U7908 (N_7908,N_7748,N_7731);
xor U7909 (N_7909,N_7691,N_7757);
or U7910 (N_7910,N_7634,N_7770);
and U7911 (N_7911,N_7602,N_7704);
nand U7912 (N_7912,N_7662,N_7788);
and U7913 (N_7913,N_7780,N_7673);
nand U7914 (N_7914,N_7775,N_7664);
xor U7915 (N_7915,N_7719,N_7699);
xnor U7916 (N_7916,N_7605,N_7642);
nand U7917 (N_7917,N_7613,N_7692);
nand U7918 (N_7918,N_7722,N_7747);
nor U7919 (N_7919,N_7783,N_7601);
xnor U7920 (N_7920,N_7723,N_7672);
nand U7921 (N_7921,N_7773,N_7612);
and U7922 (N_7922,N_7697,N_7743);
nor U7923 (N_7923,N_7660,N_7622);
xnor U7924 (N_7924,N_7788,N_7753);
or U7925 (N_7925,N_7690,N_7710);
nand U7926 (N_7926,N_7672,N_7724);
xor U7927 (N_7927,N_7742,N_7757);
nor U7928 (N_7928,N_7711,N_7751);
nor U7929 (N_7929,N_7685,N_7617);
or U7930 (N_7930,N_7611,N_7647);
nor U7931 (N_7931,N_7648,N_7679);
xor U7932 (N_7932,N_7729,N_7785);
nor U7933 (N_7933,N_7678,N_7721);
or U7934 (N_7934,N_7701,N_7718);
and U7935 (N_7935,N_7706,N_7754);
and U7936 (N_7936,N_7683,N_7611);
nor U7937 (N_7937,N_7789,N_7632);
xnor U7938 (N_7938,N_7694,N_7790);
and U7939 (N_7939,N_7749,N_7779);
and U7940 (N_7940,N_7712,N_7706);
nand U7941 (N_7941,N_7717,N_7798);
nor U7942 (N_7942,N_7724,N_7651);
xnor U7943 (N_7943,N_7688,N_7609);
or U7944 (N_7944,N_7674,N_7666);
xnor U7945 (N_7945,N_7658,N_7750);
or U7946 (N_7946,N_7764,N_7690);
and U7947 (N_7947,N_7705,N_7737);
and U7948 (N_7948,N_7660,N_7669);
xnor U7949 (N_7949,N_7758,N_7743);
xor U7950 (N_7950,N_7798,N_7638);
nor U7951 (N_7951,N_7679,N_7761);
nor U7952 (N_7952,N_7659,N_7633);
nor U7953 (N_7953,N_7713,N_7640);
or U7954 (N_7954,N_7614,N_7604);
and U7955 (N_7955,N_7693,N_7636);
and U7956 (N_7956,N_7742,N_7729);
nor U7957 (N_7957,N_7609,N_7698);
nand U7958 (N_7958,N_7726,N_7642);
or U7959 (N_7959,N_7772,N_7653);
xnor U7960 (N_7960,N_7734,N_7783);
or U7961 (N_7961,N_7749,N_7792);
nand U7962 (N_7962,N_7738,N_7748);
xor U7963 (N_7963,N_7740,N_7798);
and U7964 (N_7964,N_7654,N_7798);
xor U7965 (N_7965,N_7631,N_7704);
and U7966 (N_7966,N_7691,N_7649);
or U7967 (N_7967,N_7639,N_7742);
nor U7968 (N_7968,N_7603,N_7640);
nand U7969 (N_7969,N_7772,N_7616);
or U7970 (N_7970,N_7648,N_7700);
nor U7971 (N_7971,N_7794,N_7600);
nand U7972 (N_7972,N_7776,N_7798);
or U7973 (N_7973,N_7607,N_7683);
xnor U7974 (N_7974,N_7770,N_7717);
or U7975 (N_7975,N_7760,N_7709);
nor U7976 (N_7976,N_7702,N_7699);
or U7977 (N_7977,N_7674,N_7622);
nand U7978 (N_7978,N_7751,N_7694);
nor U7979 (N_7979,N_7694,N_7687);
xnor U7980 (N_7980,N_7704,N_7715);
and U7981 (N_7981,N_7688,N_7713);
nand U7982 (N_7982,N_7672,N_7742);
and U7983 (N_7983,N_7676,N_7692);
or U7984 (N_7984,N_7710,N_7773);
nor U7985 (N_7985,N_7676,N_7642);
nor U7986 (N_7986,N_7628,N_7764);
or U7987 (N_7987,N_7790,N_7637);
xnor U7988 (N_7988,N_7609,N_7677);
nand U7989 (N_7989,N_7690,N_7726);
and U7990 (N_7990,N_7753,N_7782);
or U7991 (N_7991,N_7713,N_7606);
nand U7992 (N_7992,N_7612,N_7664);
nand U7993 (N_7993,N_7685,N_7608);
or U7994 (N_7994,N_7705,N_7796);
or U7995 (N_7995,N_7703,N_7650);
xnor U7996 (N_7996,N_7649,N_7762);
and U7997 (N_7997,N_7710,N_7713);
or U7998 (N_7998,N_7793,N_7637);
and U7999 (N_7999,N_7752,N_7707);
xnor U8000 (N_8000,N_7974,N_7899);
and U8001 (N_8001,N_7991,N_7937);
nand U8002 (N_8002,N_7979,N_7823);
nand U8003 (N_8003,N_7866,N_7980);
nor U8004 (N_8004,N_7958,N_7912);
or U8005 (N_8005,N_7850,N_7869);
and U8006 (N_8006,N_7857,N_7889);
or U8007 (N_8007,N_7978,N_7872);
xor U8008 (N_8008,N_7911,N_7812);
nor U8009 (N_8009,N_7841,N_7842);
xnor U8010 (N_8010,N_7882,N_7894);
and U8011 (N_8011,N_7952,N_7854);
nand U8012 (N_8012,N_7888,N_7830);
nand U8013 (N_8013,N_7898,N_7943);
and U8014 (N_8014,N_7802,N_7834);
and U8015 (N_8015,N_7901,N_7821);
nand U8016 (N_8016,N_7907,N_7950);
and U8017 (N_8017,N_7849,N_7805);
nand U8018 (N_8018,N_7997,N_7946);
nand U8019 (N_8019,N_7864,N_7836);
or U8020 (N_8020,N_7846,N_7862);
xor U8021 (N_8021,N_7935,N_7878);
nand U8022 (N_8022,N_7856,N_7963);
nor U8023 (N_8023,N_7909,N_7871);
or U8024 (N_8024,N_7884,N_7896);
nand U8025 (N_8025,N_7861,N_7829);
xnor U8026 (N_8026,N_7905,N_7967);
nand U8027 (N_8027,N_7904,N_7918);
nand U8028 (N_8028,N_7895,N_7916);
nand U8029 (N_8029,N_7927,N_7932);
nor U8030 (N_8030,N_7993,N_7951);
or U8031 (N_8031,N_7810,N_7945);
nand U8032 (N_8032,N_7835,N_7971);
nand U8033 (N_8033,N_7964,N_7915);
nand U8034 (N_8034,N_7908,N_7987);
nand U8035 (N_8035,N_7928,N_7936);
xnor U8036 (N_8036,N_7879,N_7989);
nor U8037 (N_8037,N_7920,N_7970);
and U8038 (N_8038,N_7931,N_7972);
xor U8039 (N_8039,N_7876,N_7825);
xor U8040 (N_8040,N_7944,N_7953);
nor U8041 (N_8041,N_7968,N_7806);
and U8042 (N_8042,N_7839,N_7921);
xnor U8043 (N_8043,N_7845,N_7977);
and U8044 (N_8044,N_7995,N_7893);
xnor U8045 (N_8045,N_7949,N_7832);
nor U8046 (N_8046,N_7969,N_7965);
xor U8047 (N_8047,N_7811,N_7847);
nor U8048 (N_8048,N_7962,N_7807);
nand U8049 (N_8049,N_7831,N_7828);
or U8050 (N_8050,N_7827,N_7902);
xor U8051 (N_8051,N_7957,N_7852);
or U8052 (N_8052,N_7887,N_7880);
nor U8053 (N_8053,N_7985,N_7929);
nand U8054 (N_8054,N_7955,N_7804);
xor U8055 (N_8055,N_7900,N_7881);
xnor U8056 (N_8056,N_7800,N_7926);
nand U8057 (N_8057,N_7860,N_7853);
xor U8058 (N_8058,N_7976,N_7919);
or U8059 (N_8059,N_7984,N_7981);
xnor U8060 (N_8060,N_7824,N_7877);
xnor U8061 (N_8061,N_7817,N_7865);
and U8062 (N_8062,N_7875,N_7966);
or U8063 (N_8063,N_7973,N_7886);
and U8064 (N_8064,N_7990,N_7867);
and U8065 (N_8065,N_7992,N_7982);
xor U8066 (N_8066,N_7814,N_7988);
and U8067 (N_8067,N_7922,N_7942);
xnor U8068 (N_8068,N_7975,N_7947);
nor U8069 (N_8069,N_7816,N_7983);
nand U8070 (N_8070,N_7959,N_7820);
nor U8071 (N_8071,N_7848,N_7885);
nor U8072 (N_8072,N_7890,N_7933);
and U8073 (N_8073,N_7851,N_7940);
or U8074 (N_8074,N_7859,N_7868);
and U8075 (N_8075,N_7994,N_7874);
nor U8076 (N_8076,N_7934,N_7954);
nand U8077 (N_8077,N_7941,N_7913);
nand U8078 (N_8078,N_7910,N_7996);
xor U8079 (N_8079,N_7923,N_7998);
nor U8080 (N_8080,N_7999,N_7956);
nand U8081 (N_8081,N_7960,N_7801);
nand U8082 (N_8082,N_7891,N_7858);
nor U8083 (N_8083,N_7925,N_7924);
or U8084 (N_8084,N_7897,N_7855);
or U8085 (N_8085,N_7870,N_7903);
and U8086 (N_8086,N_7948,N_7822);
nor U8087 (N_8087,N_7803,N_7843);
nand U8088 (N_8088,N_7838,N_7892);
nand U8089 (N_8089,N_7930,N_7863);
or U8090 (N_8090,N_7833,N_7939);
nand U8091 (N_8091,N_7809,N_7914);
nor U8092 (N_8092,N_7826,N_7837);
nor U8093 (N_8093,N_7819,N_7808);
nand U8094 (N_8094,N_7818,N_7986);
xnor U8095 (N_8095,N_7883,N_7813);
xnor U8096 (N_8096,N_7815,N_7844);
and U8097 (N_8097,N_7873,N_7917);
and U8098 (N_8098,N_7961,N_7938);
nor U8099 (N_8099,N_7906,N_7840);
nor U8100 (N_8100,N_7868,N_7825);
nand U8101 (N_8101,N_7918,N_7970);
or U8102 (N_8102,N_7919,N_7860);
or U8103 (N_8103,N_7881,N_7884);
and U8104 (N_8104,N_7912,N_7935);
xor U8105 (N_8105,N_7800,N_7831);
xnor U8106 (N_8106,N_7858,N_7994);
or U8107 (N_8107,N_7974,N_7934);
nor U8108 (N_8108,N_7973,N_7900);
xnor U8109 (N_8109,N_7832,N_7834);
nand U8110 (N_8110,N_7867,N_7960);
and U8111 (N_8111,N_7892,N_7976);
nor U8112 (N_8112,N_7837,N_7975);
xnor U8113 (N_8113,N_7874,N_7821);
and U8114 (N_8114,N_7967,N_7961);
xor U8115 (N_8115,N_7970,N_7821);
or U8116 (N_8116,N_7951,N_7913);
nand U8117 (N_8117,N_7894,N_7975);
nor U8118 (N_8118,N_7930,N_7939);
and U8119 (N_8119,N_7802,N_7986);
or U8120 (N_8120,N_7803,N_7914);
or U8121 (N_8121,N_7891,N_7879);
xor U8122 (N_8122,N_7954,N_7821);
nand U8123 (N_8123,N_7828,N_7876);
and U8124 (N_8124,N_7829,N_7957);
nor U8125 (N_8125,N_7859,N_7907);
nor U8126 (N_8126,N_7833,N_7855);
or U8127 (N_8127,N_7934,N_7999);
xnor U8128 (N_8128,N_7986,N_7806);
xor U8129 (N_8129,N_7935,N_7819);
nand U8130 (N_8130,N_7852,N_7918);
and U8131 (N_8131,N_7901,N_7972);
and U8132 (N_8132,N_7822,N_7919);
xor U8133 (N_8133,N_7802,N_7914);
nand U8134 (N_8134,N_7981,N_7943);
nand U8135 (N_8135,N_7954,N_7923);
nor U8136 (N_8136,N_7984,N_7866);
or U8137 (N_8137,N_7971,N_7941);
nor U8138 (N_8138,N_7918,N_7994);
and U8139 (N_8139,N_7911,N_7982);
or U8140 (N_8140,N_7939,N_7875);
or U8141 (N_8141,N_7859,N_7863);
nand U8142 (N_8142,N_7974,N_7883);
nor U8143 (N_8143,N_7950,N_7838);
nor U8144 (N_8144,N_7940,N_7919);
nand U8145 (N_8145,N_7897,N_7929);
nand U8146 (N_8146,N_7969,N_7982);
nor U8147 (N_8147,N_7832,N_7854);
nor U8148 (N_8148,N_7807,N_7958);
nand U8149 (N_8149,N_7831,N_7852);
and U8150 (N_8150,N_7925,N_7832);
and U8151 (N_8151,N_7960,N_7870);
nor U8152 (N_8152,N_7979,N_7962);
xnor U8153 (N_8153,N_7903,N_7964);
or U8154 (N_8154,N_7827,N_7986);
xnor U8155 (N_8155,N_7853,N_7822);
and U8156 (N_8156,N_7980,N_7815);
nor U8157 (N_8157,N_7806,N_7969);
nor U8158 (N_8158,N_7915,N_7953);
xor U8159 (N_8159,N_7819,N_7924);
or U8160 (N_8160,N_7810,N_7901);
nor U8161 (N_8161,N_7952,N_7824);
or U8162 (N_8162,N_7988,N_7961);
xnor U8163 (N_8163,N_7870,N_7872);
xor U8164 (N_8164,N_7841,N_7816);
and U8165 (N_8165,N_7836,N_7802);
xor U8166 (N_8166,N_7831,N_7814);
nand U8167 (N_8167,N_7915,N_7994);
nor U8168 (N_8168,N_7982,N_7966);
or U8169 (N_8169,N_7855,N_7974);
or U8170 (N_8170,N_7899,N_7987);
xnor U8171 (N_8171,N_7958,N_7935);
nand U8172 (N_8172,N_7977,N_7919);
xor U8173 (N_8173,N_7834,N_7883);
nand U8174 (N_8174,N_7831,N_7857);
or U8175 (N_8175,N_7981,N_7861);
nand U8176 (N_8176,N_7848,N_7986);
nor U8177 (N_8177,N_7950,N_7998);
or U8178 (N_8178,N_7806,N_7808);
and U8179 (N_8179,N_7852,N_7811);
and U8180 (N_8180,N_7956,N_7915);
or U8181 (N_8181,N_7817,N_7824);
nor U8182 (N_8182,N_7861,N_7864);
and U8183 (N_8183,N_7948,N_7971);
or U8184 (N_8184,N_7994,N_7992);
nand U8185 (N_8185,N_7889,N_7861);
nand U8186 (N_8186,N_7987,N_7874);
and U8187 (N_8187,N_7809,N_7860);
nor U8188 (N_8188,N_7910,N_7806);
nand U8189 (N_8189,N_7813,N_7925);
xnor U8190 (N_8190,N_7977,N_7819);
or U8191 (N_8191,N_7887,N_7973);
nor U8192 (N_8192,N_7958,N_7981);
nor U8193 (N_8193,N_7933,N_7935);
nor U8194 (N_8194,N_7983,N_7887);
nand U8195 (N_8195,N_7972,N_7936);
and U8196 (N_8196,N_7871,N_7918);
nand U8197 (N_8197,N_7867,N_7821);
nand U8198 (N_8198,N_7928,N_7837);
nand U8199 (N_8199,N_7878,N_7874);
nand U8200 (N_8200,N_8002,N_8140);
xor U8201 (N_8201,N_8141,N_8186);
nand U8202 (N_8202,N_8136,N_8039);
nand U8203 (N_8203,N_8035,N_8001);
xor U8204 (N_8204,N_8183,N_8057);
xor U8205 (N_8205,N_8011,N_8025);
nand U8206 (N_8206,N_8132,N_8086);
nor U8207 (N_8207,N_8172,N_8037);
and U8208 (N_8208,N_8061,N_8159);
nand U8209 (N_8209,N_8152,N_8189);
xor U8210 (N_8210,N_8103,N_8041);
xor U8211 (N_8211,N_8145,N_8082);
and U8212 (N_8212,N_8195,N_8164);
or U8213 (N_8213,N_8079,N_8015);
nand U8214 (N_8214,N_8122,N_8089);
or U8215 (N_8215,N_8078,N_8150);
and U8216 (N_8216,N_8180,N_8157);
xor U8217 (N_8217,N_8014,N_8131);
or U8218 (N_8218,N_8040,N_8034);
nor U8219 (N_8219,N_8052,N_8104);
nor U8220 (N_8220,N_8064,N_8139);
and U8221 (N_8221,N_8044,N_8087);
xor U8222 (N_8222,N_8051,N_8065);
nand U8223 (N_8223,N_8028,N_8162);
xor U8224 (N_8224,N_8017,N_8054);
xnor U8225 (N_8225,N_8097,N_8032);
and U8226 (N_8226,N_8042,N_8059);
nand U8227 (N_8227,N_8080,N_8009);
or U8228 (N_8228,N_8096,N_8113);
nand U8229 (N_8229,N_8175,N_8111);
nand U8230 (N_8230,N_8194,N_8135);
and U8231 (N_8231,N_8003,N_8105);
and U8232 (N_8232,N_8013,N_8010);
or U8233 (N_8233,N_8036,N_8119);
nor U8234 (N_8234,N_8165,N_8134);
and U8235 (N_8235,N_8112,N_8045);
or U8236 (N_8236,N_8053,N_8121);
and U8237 (N_8237,N_8169,N_8149);
xor U8238 (N_8238,N_8107,N_8153);
or U8239 (N_8239,N_8008,N_8148);
nor U8240 (N_8240,N_8127,N_8088);
or U8241 (N_8241,N_8171,N_8117);
nor U8242 (N_8242,N_8048,N_8160);
and U8243 (N_8243,N_8047,N_8043);
and U8244 (N_8244,N_8144,N_8049);
or U8245 (N_8245,N_8055,N_8120);
xnor U8246 (N_8246,N_8137,N_8075);
or U8247 (N_8247,N_8093,N_8038);
xnor U8248 (N_8248,N_8099,N_8147);
nor U8249 (N_8249,N_8109,N_8155);
xnor U8250 (N_8250,N_8068,N_8181);
xor U8251 (N_8251,N_8158,N_8197);
and U8252 (N_8252,N_8161,N_8006);
nor U8253 (N_8253,N_8170,N_8138);
or U8254 (N_8254,N_8023,N_8072);
or U8255 (N_8255,N_8187,N_8090);
nand U8256 (N_8256,N_8179,N_8026);
nand U8257 (N_8257,N_8128,N_8033);
nor U8258 (N_8258,N_8108,N_8130);
nand U8259 (N_8259,N_8046,N_8004);
and U8260 (N_8260,N_8074,N_8178);
nand U8261 (N_8261,N_8116,N_8110);
nand U8262 (N_8262,N_8174,N_8166);
and U8263 (N_8263,N_8063,N_8142);
or U8264 (N_8264,N_8073,N_8083);
or U8265 (N_8265,N_8076,N_8114);
and U8266 (N_8266,N_8071,N_8177);
nand U8267 (N_8267,N_8118,N_8196);
nand U8268 (N_8268,N_8007,N_8115);
xor U8269 (N_8269,N_8021,N_8173);
xor U8270 (N_8270,N_8094,N_8184);
and U8271 (N_8271,N_8192,N_8066);
and U8272 (N_8272,N_8106,N_8024);
nor U8273 (N_8273,N_8019,N_8124);
nor U8274 (N_8274,N_8081,N_8022);
xor U8275 (N_8275,N_8069,N_8000);
and U8276 (N_8276,N_8091,N_8016);
and U8277 (N_8277,N_8198,N_8129);
xor U8278 (N_8278,N_8146,N_8005);
nand U8279 (N_8279,N_8070,N_8077);
and U8280 (N_8280,N_8182,N_8067);
nand U8281 (N_8281,N_8056,N_8143);
nand U8282 (N_8282,N_8050,N_8154);
or U8283 (N_8283,N_8133,N_8084);
and U8284 (N_8284,N_8100,N_8092);
nand U8285 (N_8285,N_8102,N_8190);
and U8286 (N_8286,N_8191,N_8012);
xor U8287 (N_8287,N_8176,N_8185);
nand U8288 (N_8288,N_8123,N_8101);
nor U8289 (N_8289,N_8060,N_8167);
xor U8290 (N_8290,N_8095,N_8085);
nand U8291 (N_8291,N_8151,N_8098);
or U8292 (N_8292,N_8126,N_8193);
and U8293 (N_8293,N_8168,N_8018);
nand U8294 (N_8294,N_8163,N_8058);
nand U8295 (N_8295,N_8027,N_8199);
nand U8296 (N_8296,N_8031,N_8030);
nor U8297 (N_8297,N_8062,N_8020);
xor U8298 (N_8298,N_8029,N_8188);
or U8299 (N_8299,N_8125,N_8156);
or U8300 (N_8300,N_8126,N_8006);
nand U8301 (N_8301,N_8098,N_8095);
nor U8302 (N_8302,N_8036,N_8003);
xor U8303 (N_8303,N_8110,N_8184);
xor U8304 (N_8304,N_8050,N_8026);
nand U8305 (N_8305,N_8141,N_8027);
or U8306 (N_8306,N_8087,N_8006);
and U8307 (N_8307,N_8094,N_8163);
xnor U8308 (N_8308,N_8198,N_8158);
nor U8309 (N_8309,N_8079,N_8166);
xnor U8310 (N_8310,N_8148,N_8138);
nor U8311 (N_8311,N_8118,N_8103);
and U8312 (N_8312,N_8048,N_8056);
nand U8313 (N_8313,N_8185,N_8190);
nand U8314 (N_8314,N_8032,N_8153);
nand U8315 (N_8315,N_8115,N_8093);
nor U8316 (N_8316,N_8082,N_8125);
and U8317 (N_8317,N_8039,N_8182);
nor U8318 (N_8318,N_8009,N_8073);
and U8319 (N_8319,N_8042,N_8144);
xnor U8320 (N_8320,N_8047,N_8111);
nor U8321 (N_8321,N_8027,N_8167);
nor U8322 (N_8322,N_8066,N_8063);
nor U8323 (N_8323,N_8168,N_8062);
and U8324 (N_8324,N_8152,N_8030);
or U8325 (N_8325,N_8117,N_8087);
or U8326 (N_8326,N_8045,N_8188);
nor U8327 (N_8327,N_8083,N_8126);
nor U8328 (N_8328,N_8062,N_8111);
nor U8329 (N_8329,N_8013,N_8130);
nand U8330 (N_8330,N_8104,N_8063);
nand U8331 (N_8331,N_8041,N_8018);
or U8332 (N_8332,N_8066,N_8176);
nand U8333 (N_8333,N_8085,N_8198);
or U8334 (N_8334,N_8186,N_8060);
xnor U8335 (N_8335,N_8015,N_8007);
nand U8336 (N_8336,N_8189,N_8062);
and U8337 (N_8337,N_8074,N_8155);
xor U8338 (N_8338,N_8052,N_8102);
nor U8339 (N_8339,N_8145,N_8110);
or U8340 (N_8340,N_8074,N_8141);
nand U8341 (N_8341,N_8192,N_8100);
or U8342 (N_8342,N_8116,N_8043);
or U8343 (N_8343,N_8022,N_8000);
or U8344 (N_8344,N_8190,N_8091);
and U8345 (N_8345,N_8176,N_8069);
nand U8346 (N_8346,N_8056,N_8053);
nand U8347 (N_8347,N_8090,N_8171);
nand U8348 (N_8348,N_8014,N_8183);
nand U8349 (N_8349,N_8194,N_8197);
nand U8350 (N_8350,N_8014,N_8040);
nor U8351 (N_8351,N_8155,N_8057);
nand U8352 (N_8352,N_8029,N_8192);
xor U8353 (N_8353,N_8029,N_8038);
or U8354 (N_8354,N_8188,N_8081);
or U8355 (N_8355,N_8162,N_8097);
nand U8356 (N_8356,N_8184,N_8148);
or U8357 (N_8357,N_8194,N_8063);
xor U8358 (N_8358,N_8180,N_8123);
nand U8359 (N_8359,N_8121,N_8197);
or U8360 (N_8360,N_8141,N_8018);
or U8361 (N_8361,N_8179,N_8075);
and U8362 (N_8362,N_8010,N_8105);
and U8363 (N_8363,N_8008,N_8132);
nor U8364 (N_8364,N_8088,N_8074);
nor U8365 (N_8365,N_8081,N_8054);
and U8366 (N_8366,N_8036,N_8090);
nand U8367 (N_8367,N_8073,N_8186);
nor U8368 (N_8368,N_8198,N_8092);
nand U8369 (N_8369,N_8156,N_8003);
nor U8370 (N_8370,N_8068,N_8008);
xnor U8371 (N_8371,N_8074,N_8186);
nor U8372 (N_8372,N_8110,N_8094);
xor U8373 (N_8373,N_8038,N_8070);
nor U8374 (N_8374,N_8089,N_8147);
or U8375 (N_8375,N_8042,N_8099);
nand U8376 (N_8376,N_8114,N_8077);
nor U8377 (N_8377,N_8187,N_8178);
xnor U8378 (N_8378,N_8116,N_8170);
nand U8379 (N_8379,N_8189,N_8188);
nor U8380 (N_8380,N_8130,N_8159);
xnor U8381 (N_8381,N_8089,N_8018);
nor U8382 (N_8382,N_8099,N_8017);
nor U8383 (N_8383,N_8028,N_8159);
and U8384 (N_8384,N_8050,N_8176);
xor U8385 (N_8385,N_8085,N_8112);
or U8386 (N_8386,N_8091,N_8057);
or U8387 (N_8387,N_8170,N_8007);
and U8388 (N_8388,N_8130,N_8165);
or U8389 (N_8389,N_8182,N_8031);
or U8390 (N_8390,N_8001,N_8060);
xnor U8391 (N_8391,N_8160,N_8158);
nor U8392 (N_8392,N_8174,N_8183);
or U8393 (N_8393,N_8170,N_8133);
nor U8394 (N_8394,N_8145,N_8111);
nor U8395 (N_8395,N_8104,N_8161);
xnor U8396 (N_8396,N_8187,N_8108);
or U8397 (N_8397,N_8087,N_8041);
or U8398 (N_8398,N_8114,N_8159);
or U8399 (N_8399,N_8027,N_8056);
xnor U8400 (N_8400,N_8311,N_8226);
and U8401 (N_8401,N_8396,N_8343);
nor U8402 (N_8402,N_8379,N_8253);
and U8403 (N_8403,N_8377,N_8242);
xor U8404 (N_8404,N_8262,N_8299);
and U8405 (N_8405,N_8326,N_8254);
nand U8406 (N_8406,N_8295,N_8392);
xnor U8407 (N_8407,N_8364,N_8237);
xnor U8408 (N_8408,N_8363,N_8244);
nor U8409 (N_8409,N_8276,N_8283);
or U8410 (N_8410,N_8315,N_8266);
nor U8411 (N_8411,N_8212,N_8227);
and U8412 (N_8412,N_8230,N_8210);
and U8413 (N_8413,N_8308,N_8313);
xor U8414 (N_8414,N_8232,N_8294);
or U8415 (N_8415,N_8215,N_8289);
and U8416 (N_8416,N_8307,N_8332);
nand U8417 (N_8417,N_8274,N_8290);
nor U8418 (N_8418,N_8269,N_8324);
and U8419 (N_8419,N_8345,N_8355);
nor U8420 (N_8420,N_8206,N_8383);
and U8421 (N_8421,N_8257,N_8261);
xnor U8422 (N_8422,N_8204,N_8318);
nand U8423 (N_8423,N_8368,N_8342);
nor U8424 (N_8424,N_8258,N_8301);
and U8425 (N_8425,N_8293,N_8325);
and U8426 (N_8426,N_8217,N_8229);
nor U8427 (N_8427,N_8251,N_8200);
and U8428 (N_8428,N_8391,N_8234);
nand U8429 (N_8429,N_8225,N_8341);
xnor U8430 (N_8430,N_8216,N_8384);
or U8431 (N_8431,N_8298,N_8213);
nor U8432 (N_8432,N_8334,N_8281);
nor U8433 (N_8433,N_8287,N_8279);
or U8434 (N_8434,N_8390,N_8310);
xor U8435 (N_8435,N_8350,N_8381);
xnor U8436 (N_8436,N_8271,N_8248);
nand U8437 (N_8437,N_8344,N_8359);
or U8438 (N_8438,N_8238,N_8235);
xor U8439 (N_8439,N_8354,N_8277);
or U8440 (N_8440,N_8399,N_8208);
nand U8441 (N_8441,N_8314,N_8241);
xor U8442 (N_8442,N_8265,N_8239);
nor U8443 (N_8443,N_8221,N_8317);
nand U8444 (N_8444,N_8339,N_8353);
nand U8445 (N_8445,N_8367,N_8246);
or U8446 (N_8446,N_8340,N_8349);
or U8447 (N_8447,N_8267,N_8275);
and U8448 (N_8448,N_8333,N_8236);
nand U8449 (N_8449,N_8320,N_8321);
nor U8450 (N_8450,N_8338,N_8323);
or U8451 (N_8451,N_8375,N_8231);
nor U8452 (N_8452,N_8336,N_8385);
and U8453 (N_8453,N_8365,N_8335);
xor U8454 (N_8454,N_8280,N_8263);
xor U8455 (N_8455,N_8366,N_8376);
nand U8456 (N_8456,N_8252,N_8233);
and U8457 (N_8457,N_8331,N_8347);
nand U8458 (N_8458,N_8218,N_8352);
nor U8459 (N_8459,N_8291,N_8249);
and U8460 (N_8460,N_8296,N_8305);
nand U8461 (N_8461,N_8322,N_8360);
or U8462 (N_8462,N_8386,N_8316);
or U8463 (N_8463,N_8374,N_8205);
or U8464 (N_8464,N_8378,N_8203);
nor U8465 (N_8465,N_8398,N_8348);
nor U8466 (N_8466,N_8369,N_8223);
xnor U8467 (N_8467,N_8397,N_8211);
or U8468 (N_8468,N_8201,N_8243);
or U8469 (N_8469,N_8288,N_8255);
and U8470 (N_8470,N_8319,N_8260);
xor U8471 (N_8471,N_8395,N_8282);
nor U8472 (N_8472,N_8330,N_8380);
xor U8473 (N_8473,N_8264,N_8222);
nand U8474 (N_8474,N_8302,N_8224);
nand U8475 (N_8475,N_8207,N_8303);
nor U8476 (N_8476,N_8270,N_8245);
or U8477 (N_8477,N_8328,N_8358);
nor U8478 (N_8478,N_8373,N_8361);
nand U8479 (N_8479,N_8284,N_8312);
or U8480 (N_8480,N_8300,N_8393);
or U8481 (N_8481,N_8346,N_8268);
nand U8482 (N_8482,N_8259,N_8309);
xnor U8483 (N_8483,N_8329,N_8273);
or U8484 (N_8484,N_8256,N_8388);
nand U8485 (N_8485,N_8228,N_8219);
xor U8486 (N_8486,N_8327,N_8247);
xor U8487 (N_8487,N_8214,N_8371);
nor U8488 (N_8488,N_8357,N_8278);
or U8489 (N_8489,N_8286,N_8372);
or U8490 (N_8490,N_8202,N_8337);
xnor U8491 (N_8491,N_8250,N_8389);
or U8492 (N_8492,N_8394,N_8292);
nor U8493 (N_8493,N_8220,N_8285);
nor U8494 (N_8494,N_8272,N_8304);
and U8495 (N_8495,N_8209,N_8362);
or U8496 (N_8496,N_8356,N_8306);
nor U8497 (N_8497,N_8370,N_8351);
xor U8498 (N_8498,N_8297,N_8240);
xor U8499 (N_8499,N_8382,N_8387);
nor U8500 (N_8500,N_8203,N_8236);
xor U8501 (N_8501,N_8358,N_8324);
and U8502 (N_8502,N_8325,N_8273);
or U8503 (N_8503,N_8245,N_8341);
nand U8504 (N_8504,N_8347,N_8222);
xnor U8505 (N_8505,N_8343,N_8260);
or U8506 (N_8506,N_8318,N_8233);
xor U8507 (N_8507,N_8297,N_8235);
or U8508 (N_8508,N_8387,N_8302);
and U8509 (N_8509,N_8321,N_8353);
nand U8510 (N_8510,N_8220,N_8294);
nor U8511 (N_8511,N_8315,N_8208);
xnor U8512 (N_8512,N_8282,N_8290);
or U8513 (N_8513,N_8349,N_8374);
xnor U8514 (N_8514,N_8320,N_8217);
nand U8515 (N_8515,N_8323,N_8213);
or U8516 (N_8516,N_8280,N_8226);
and U8517 (N_8517,N_8213,N_8273);
nand U8518 (N_8518,N_8257,N_8392);
xnor U8519 (N_8519,N_8251,N_8243);
xor U8520 (N_8520,N_8227,N_8294);
nand U8521 (N_8521,N_8201,N_8396);
and U8522 (N_8522,N_8340,N_8263);
nand U8523 (N_8523,N_8224,N_8222);
nand U8524 (N_8524,N_8250,N_8355);
and U8525 (N_8525,N_8336,N_8350);
nand U8526 (N_8526,N_8303,N_8202);
xnor U8527 (N_8527,N_8378,N_8228);
nor U8528 (N_8528,N_8216,N_8228);
nor U8529 (N_8529,N_8326,N_8284);
or U8530 (N_8530,N_8225,N_8243);
xnor U8531 (N_8531,N_8339,N_8306);
and U8532 (N_8532,N_8387,N_8365);
xnor U8533 (N_8533,N_8280,N_8393);
and U8534 (N_8534,N_8258,N_8352);
and U8535 (N_8535,N_8326,N_8317);
and U8536 (N_8536,N_8297,N_8289);
and U8537 (N_8537,N_8366,N_8309);
nand U8538 (N_8538,N_8212,N_8284);
xor U8539 (N_8539,N_8236,N_8220);
xor U8540 (N_8540,N_8356,N_8340);
nor U8541 (N_8541,N_8259,N_8393);
nor U8542 (N_8542,N_8373,N_8308);
or U8543 (N_8543,N_8350,N_8379);
nor U8544 (N_8544,N_8238,N_8294);
xnor U8545 (N_8545,N_8260,N_8308);
nor U8546 (N_8546,N_8245,N_8212);
xor U8547 (N_8547,N_8302,N_8297);
nor U8548 (N_8548,N_8228,N_8304);
xnor U8549 (N_8549,N_8202,N_8220);
nor U8550 (N_8550,N_8317,N_8268);
nand U8551 (N_8551,N_8200,N_8238);
xnor U8552 (N_8552,N_8311,N_8253);
nor U8553 (N_8553,N_8358,N_8332);
nand U8554 (N_8554,N_8201,N_8297);
and U8555 (N_8555,N_8356,N_8300);
and U8556 (N_8556,N_8271,N_8272);
or U8557 (N_8557,N_8266,N_8371);
nand U8558 (N_8558,N_8350,N_8241);
and U8559 (N_8559,N_8245,N_8379);
nor U8560 (N_8560,N_8319,N_8386);
or U8561 (N_8561,N_8271,N_8393);
nand U8562 (N_8562,N_8286,N_8274);
xor U8563 (N_8563,N_8252,N_8310);
and U8564 (N_8564,N_8225,N_8397);
or U8565 (N_8565,N_8378,N_8273);
xnor U8566 (N_8566,N_8265,N_8388);
and U8567 (N_8567,N_8386,N_8212);
nor U8568 (N_8568,N_8303,N_8225);
nand U8569 (N_8569,N_8317,N_8312);
xor U8570 (N_8570,N_8255,N_8289);
nor U8571 (N_8571,N_8353,N_8300);
and U8572 (N_8572,N_8256,N_8345);
or U8573 (N_8573,N_8298,N_8273);
and U8574 (N_8574,N_8252,N_8204);
xor U8575 (N_8575,N_8379,N_8331);
or U8576 (N_8576,N_8292,N_8228);
or U8577 (N_8577,N_8385,N_8352);
and U8578 (N_8578,N_8206,N_8303);
xor U8579 (N_8579,N_8298,N_8208);
xnor U8580 (N_8580,N_8219,N_8223);
xnor U8581 (N_8581,N_8338,N_8361);
xor U8582 (N_8582,N_8250,N_8330);
and U8583 (N_8583,N_8234,N_8283);
xor U8584 (N_8584,N_8305,N_8209);
nor U8585 (N_8585,N_8250,N_8270);
xor U8586 (N_8586,N_8375,N_8235);
xnor U8587 (N_8587,N_8377,N_8298);
nand U8588 (N_8588,N_8387,N_8353);
xnor U8589 (N_8589,N_8384,N_8256);
nand U8590 (N_8590,N_8251,N_8261);
or U8591 (N_8591,N_8208,N_8274);
and U8592 (N_8592,N_8345,N_8259);
nor U8593 (N_8593,N_8365,N_8263);
or U8594 (N_8594,N_8258,N_8306);
and U8595 (N_8595,N_8323,N_8307);
and U8596 (N_8596,N_8205,N_8204);
or U8597 (N_8597,N_8215,N_8210);
and U8598 (N_8598,N_8274,N_8387);
nand U8599 (N_8599,N_8223,N_8251);
nand U8600 (N_8600,N_8518,N_8533);
or U8601 (N_8601,N_8467,N_8411);
and U8602 (N_8602,N_8549,N_8548);
nor U8603 (N_8603,N_8406,N_8568);
nor U8604 (N_8604,N_8538,N_8443);
or U8605 (N_8605,N_8501,N_8546);
nand U8606 (N_8606,N_8488,N_8410);
nor U8607 (N_8607,N_8516,N_8480);
or U8608 (N_8608,N_8553,N_8560);
and U8609 (N_8609,N_8595,N_8508);
and U8610 (N_8610,N_8441,N_8456);
nand U8611 (N_8611,N_8412,N_8517);
nor U8612 (N_8612,N_8558,N_8529);
and U8613 (N_8613,N_8557,N_8421);
nor U8614 (N_8614,N_8453,N_8449);
xnor U8615 (N_8615,N_8567,N_8524);
nor U8616 (N_8616,N_8485,N_8445);
xor U8617 (N_8617,N_8500,N_8520);
nor U8618 (N_8618,N_8574,N_8489);
or U8619 (N_8619,N_8572,N_8483);
nor U8620 (N_8620,N_8461,N_8432);
nand U8621 (N_8621,N_8505,N_8593);
nand U8622 (N_8622,N_8576,N_8434);
nor U8623 (N_8623,N_8436,N_8504);
xnor U8624 (N_8624,N_8550,N_8519);
or U8625 (N_8625,N_8458,N_8440);
or U8626 (N_8626,N_8506,N_8400);
xor U8627 (N_8627,N_8472,N_8465);
nand U8628 (N_8628,N_8405,N_8507);
nor U8629 (N_8629,N_8455,N_8495);
xnor U8630 (N_8630,N_8589,N_8464);
nor U8631 (N_8631,N_8466,N_8578);
nor U8632 (N_8632,N_8566,N_8498);
and U8633 (N_8633,N_8547,N_8424);
or U8634 (N_8634,N_8484,N_8562);
and U8635 (N_8635,N_8428,N_8515);
or U8636 (N_8636,N_8552,N_8462);
or U8637 (N_8637,N_8563,N_8570);
nand U8638 (N_8638,N_8571,N_8527);
nand U8639 (N_8639,N_8435,N_8426);
xnor U8640 (N_8640,N_8569,N_8477);
or U8641 (N_8641,N_8416,N_8418);
nand U8642 (N_8642,N_8404,N_8536);
nor U8643 (N_8643,N_8584,N_8540);
nor U8644 (N_8644,N_8448,N_8414);
xnor U8645 (N_8645,N_8523,N_8587);
or U8646 (N_8646,N_8486,N_8582);
xnor U8647 (N_8647,N_8544,N_8564);
and U8648 (N_8648,N_8588,N_8542);
or U8649 (N_8649,N_8473,N_8402);
and U8650 (N_8650,N_8471,N_8452);
nor U8651 (N_8651,N_8450,N_8497);
xnor U8652 (N_8652,N_8415,N_8522);
nand U8653 (N_8653,N_8460,N_8541);
or U8654 (N_8654,N_8511,N_8451);
nand U8655 (N_8655,N_8401,N_8429);
nand U8656 (N_8656,N_8512,N_8407);
and U8657 (N_8657,N_8598,N_8559);
nand U8658 (N_8658,N_8446,N_8437);
xor U8659 (N_8659,N_8534,N_8439);
or U8660 (N_8660,N_8463,N_8438);
and U8661 (N_8661,N_8459,N_8554);
or U8662 (N_8662,N_8444,N_8430);
or U8663 (N_8663,N_8528,N_8478);
nand U8664 (N_8664,N_8509,N_8590);
and U8665 (N_8665,N_8510,N_8491);
and U8666 (N_8666,N_8532,N_8475);
nand U8667 (N_8667,N_8565,N_8530);
nand U8668 (N_8668,N_8585,N_8499);
nand U8669 (N_8669,N_8513,N_8575);
or U8670 (N_8670,N_8420,N_8427);
or U8671 (N_8671,N_8413,N_8408);
and U8672 (N_8672,N_8470,N_8599);
or U8673 (N_8673,N_8417,N_8592);
and U8674 (N_8674,N_8537,N_8469);
nor U8675 (N_8675,N_8403,N_8577);
xnor U8676 (N_8676,N_8531,N_8454);
xor U8677 (N_8677,N_8580,N_8545);
nor U8678 (N_8678,N_8457,N_8502);
or U8679 (N_8679,N_8481,N_8526);
or U8680 (N_8680,N_8597,N_8479);
xor U8681 (N_8681,N_8423,N_8442);
nor U8682 (N_8682,N_8419,N_8521);
and U8683 (N_8683,N_8583,N_8543);
or U8684 (N_8684,N_8490,N_8492);
nand U8685 (N_8685,N_8433,N_8596);
nand U8686 (N_8686,N_8482,N_8573);
or U8687 (N_8687,N_8539,N_8535);
nand U8688 (N_8688,N_8586,N_8409);
and U8689 (N_8689,N_8561,N_8487);
or U8690 (N_8690,N_8431,N_8591);
and U8691 (N_8691,N_8555,N_8476);
and U8692 (N_8692,N_8581,N_8556);
and U8693 (N_8693,N_8594,N_8422);
and U8694 (N_8694,N_8425,N_8496);
and U8695 (N_8695,N_8494,N_8493);
nor U8696 (N_8696,N_8579,N_8503);
nor U8697 (N_8697,N_8525,N_8551);
and U8698 (N_8698,N_8474,N_8447);
xnor U8699 (N_8699,N_8468,N_8514);
nor U8700 (N_8700,N_8490,N_8515);
and U8701 (N_8701,N_8417,N_8525);
nand U8702 (N_8702,N_8571,N_8472);
or U8703 (N_8703,N_8454,N_8414);
and U8704 (N_8704,N_8446,N_8417);
nor U8705 (N_8705,N_8510,N_8422);
nor U8706 (N_8706,N_8496,N_8581);
or U8707 (N_8707,N_8532,N_8578);
and U8708 (N_8708,N_8536,N_8576);
nand U8709 (N_8709,N_8544,N_8455);
and U8710 (N_8710,N_8501,N_8582);
nor U8711 (N_8711,N_8437,N_8506);
nor U8712 (N_8712,N_8567,N_8465);
nor U8713 (N_8713,N_8552,N_8543);
and U8714 (N_8714,N_8580,N_8499);
nand U8715 (N_8715,N_8509,N_8586);
nor U8716 (N_8716,N_8448,N_8458);
or U8717 (N_8717,N_8538,N_8445);
xnor U8718 (N_8718,N_8507,N_8463);
or U8719 (N_8719,N_8409,N_8582);
nor U8720 (N_8720,N_8501,N_8453);
nor U8721 (N_8721,N_8453,N_8423);
xor U8722 (N_8722,N_8443,N_8550);
nand U8723 (N_8723,N_8412,N_8592);
nand U8724 (N_8724,N_8499,N_8537);
or U8725 (N_8725,N_8481,N_8584);
or U8726 (N_8726,N_8560,N_8423);
and U8727 (N_8727,N_8426,N_8555);
and U8728 (N_8728,N_8563,N_8463);
and U8729 (N_8729,N_8581,N_8456);
nor U8730 (N_8730,N_8464,N_8569);
and U8731 (N_8731,N_8572,N_8433);
and U8732 (N_8732,N_8575,N_8534);
and U8733 (N_8733,N_8575,N_8493);
xnor U8734 (N_8734,N_8576,N_8586);
nand U8735 (N_8735,N_8460,N_8463);
xnor U8736 (N_8736,N_8450,N_8561);
nor U8737 (N_8737,N_8554,N_8476);
nor U8738 (N_8738,N_8575,N_8570);
nand U8739 (N_8739,N_8424,N_8418);
or U8740 (N_8740,N_8442,N_8519);
nor U8741 (N_8741,N_8410,N_8562);
and U8742 (N_8742,N_8511,N_8518);
and U8743 (N_8743,N_8503,N_8568);
and U8744 (N_8744,N_8560,N_8426);
nor U8745 (N_8745,N_8525,N_8557);
and U8746 (N_8746,N_8598,N_8431);
nand U8747 (N_8747,N_8485,N_8407);
nor U8748 (N_8748,N_8422,N_8477);
and U8749 (N_8749,N_8457,N_8415);
nor U8750 (N_8750,N_8423,N_8526);
and U8751 (N_8751,N_8547,N_8452);
xnor U8752 (N_8752,N_8582,N_8412);
nand U8753 (N_8753,N_8571,N_8500);
nor U8754 (N_8754,N_8457,N_8528);
and U8755 (N_8755,N_8548,N_8477);
xor U8756 (N_8756,N_8441,N_8401);
or U8757 (N_8757,N_8468,N_8589);
or U8758 (N_8758,N_8400,N_8413);
nand U8759 (N_8759,N_8513,N_8549);
xor U8760 (N_8760,N_8560,N_8531);
or U8761 (N_8761,N_8584,N_8559);
or U8762 (N_8762,N_8516,N_8477);
or U8763 (N_8763,N_8590,N_8517);
nor U8764 (N_8764,N_8534,N_8495);
nand U8765 (N_8765,N_8565,N_8545);
or U8766 (N_8766,N_8495,N_8506);
nand U8767 (N_8767,N_8400,N_8554);
and U8768 (N_8768,N_8451,N_8513);
nand U8769 (N_8769,N_8433,N_8496);
and U8770 (N_8770,N_8412,N_8404);
xor U8771 (N_8771,N_8594,N_8576);
nor U8772 (N_8772,N_8448,N_8553);
nor U8773 (N_8773,N_8475,N_8474);
nor U8774 (N_8774,N_8588,N_8412);
and U8775 (N_8775,N_8453,N_8570);
nor U8776 (N_8776,N_8508,N_8598);
nor U8777 (N_8777,N_8553,N_8525);
and U8778 (N_8778,N_8499,N_8474);
xnor U8779 (N_8779,N_8580,N_8495);
nor U8780 (N_8780,N_8492,N_8530);
xnor U8781 (N_8781,N_8517,N_8534);
nand U8782 (N_8782,N_8521,N_8568);
nand U8783 (N_8783,N_8547,N_8463);
or U8784 (N_8784,N_8408,N_8449);
or U8785 (N_8785,N_8592,N_8527);
nor U8786 (N_8786,N_8560,N_8424);
xnor U8787 (N_8787,N_8555,N_8533);
xnor U8788 (N_8788,N_8598,N_8558);
or U8789 (N_8789,N_8437,N_8447);
nor U8790 (N_8790,N_8568,N_8545);
or U8791 (N_8791,N_8500,N_8417);
or U8792 (N_8792,N_8435,N_8434);
nor U8793 (N_8793,N_8405,N_8481);
nand U8794 (N_8794,N_8526,N_8471);
and U8795 (N_8795,N_8570,N_8541);
or U8796 (N_8796,N_8414,N_8553);
or U8797 (N_8797,N_8417,N_8458);
nand U8798 (N_8798,N_8505,N_8499);
nand U8799 (N_8799,N_8467,N_8529);
and U8800 (N_8800,N_8757,N_8645);
and U8801 (N_8801,N_8661,N_8706);
nand U8802 (N_8802,N_8654,N_8644);
or U8803 (N_8803,N_8603,N_8610);
or U8804 (N_8804,N_8673,N_8617);
xor U8805 (N_8805,N_8724,N_8682);
nor U8806 (N_8806,N_8620,N_8747);
nor U8807 (N_8807,N_8798,N_8771);
nand U8808 (N_8808,N_8625,N_8745);
nor U8809 (N_8809,N_8780,N_8729);
nor U8810 (N_8810,N_8611,N_8762);
nand U8811 (N_8811,N_8672,N_8664);
or U8812 (N_8812,N_8693,N_8643);
nor U8813 (N_8813,N_8632,N_8769);
and U8814 (N_8814,N_8731,N_8739);
nand U8815 (N_8815,N_8680,N_8770);
nand U8816 (N_8816,N_8707,N_8733);
and U8817 (N_8817,N_8789,N_8716);
or U8818 (N_8818,N_8709,N_8776);
xnor U8819 (N_8819,N_8640,N_8656);
and U8820 (N_8820,N_8718,N_8691);
or U8821 (N_8821,N_8658,N_8665);
xor U8822 (N_8822,N_8626,N_8607);
or U8823 (N_8823,N_8649,N_8767);
nand U8824 (N_8824,N_8773,N_8705);
nand U8825 (N_8825,N_8622,N_8734);
and U8826 (N_8826,N_8676,N_8655);
xor U8827 (N_8827,N_8786,N_8624);
nand U8828 (N_8828,N_8646,N_8638);
nor U8829 (N_8829,N_8618,N_8712);
nand U8830 (N_8830,N_8764,N_8717);
nand U8831 (N_8831,N_8668,N_8787);
nor U8832 (N_8832,N_8799,N_8621);
xor U8833 (N_8833,N_8779,N_8660);
nand U8834 (N_8834,N_8698,N_8736);
nor U8835 (N_8835,N_8600,N_8659);
xor U8836 (N_8836,N_8781,N_8761);
xnor U8837 (N_8837,N_8637,N_8768);
or U8838 (N_8838,N_8641,N_8687);
or U8839 (N_8839,N_8627,N_8679);
and U8840 (N_8840,N_8633,N_8681);
nand U8841 (N_8841,N_8666,N_8636);
nor U8842 (N_8842,N_8721,N_8732);
nand U8843 (N_8843,N_8752,N_8735);
nor U8844 (N_8844,N_8606,N_8697);
and U8845 (N_8845,N_8675,N_8642);
nand U8846 (N_8846,N_8604,N_8631);
or U8847 (N_8847,N_8727,N_8674);
nor U8848 (N_8848,N_8628,N_8728);
xnor U8849 (N_8849,N_8737,N_8652);
nand U8850 (N_8850,N_8684,N_8790);
xor U8851 (N_8851,N_8692,N_8630);
nand U8852 (N_8852,N_8651,N_8722);
nand U8853 (N_8853,N_8602,N_8743);
and U8854 (N_8854,N_8695,N_8702);
or U8855 (N_8855,N_8609,N_8700);
nor U8856 (N_8856,N_8726,N_8748);
nor U8857 (N_8857,N_8758,N_8775);
xor U8858 (N_8858,N_8614,N_8797);
and U8859 (N_8859,N_8784,N_8714);
or U8860 (N_8860,N_8696,N_8763);
nor U8861 (N_8861,N_8785,N_8608);
and U8862 (N_8862,N_8663,N_8788);
and U8863 (N_8863,N_8635,N_8662);
nand U8864 (N_8864,N_8791,N_8647);
and U8865 (N_8865,N_8694,N_8751);
nand U8866 (N_8866,N_8794,N_8754);
and U8867 (N_8867,N_8669,N_8738);
xnor U8868 (N_8868,N_8605,N_8629);
nand U8869 (N_8869,N_8750,N_8760);
or U8870 (N_8870,N_8612,N_8653);
or U8871 (N_8871,N_8723,N_8701);
or U8872 (N_8872,N_8708,N_8753);
xnor U8873 (N_8873,N_8657,N_8783);
nor U8874 (N_8874,N_8616,N_8686);
nor U8875 (N_8875,N_8678,N_8782);
nor U8876 (N_8876,N_8746,N_8766);
and U8877 (N_8877,N_8650,N_8710);
xnor U8878 (N_8878,N_8615,N_8756);
and U8879 (N_8879,N_8699,N_8740);
nor U8880 (N_8880,N_8741,N_8703);
and U8881 (N_8881,N_8759,N_8793);
nor U8882 (N_8882,N_8619,N_8765);
nand U8883 (N_8883,N_8755,N_8796);
nor U8884 (N_8884,N_8742,N_8670);
xnor U8885 (N_8885,N_8725,N_8667);
and U8886 (N_8886,N_8720,N_8685);
nand U8887 (N_8887,N_8730,N_8774);
nand U8888 (N_8888,N_8648,N_8795);
nor U8889 (N_8889,N_8690,N_8683);
nor U8890 (N_8890,N_8677,N_8792);
xor U8891 (N_8891,N_8778,N_8719);
nor U8892 (N_8892,N_8711,N_8671);
and U8893 (N_8893,N_8601,N_8623);
xor U8894 (N_8894,N_8772,N_8688);
and U8895 (N_8895,N_8613,N_8713);
nor U8896 (N_8896,N_8715,N_8749);
xor U8897 (N_8897,N_8777,N_8689);
and U8898 (N_8898,N_8639,N_8634);
nand U8899 (N_8899,N_8704,N_8744);
xor U8900 (N_8900,N_8711,N_8798);
xnor U8901 (N_8901,N_8649,N_8772);
or U8902 (N_8902,N_8600,N_8654);
nor U8903 (N_8903,N_8752,N_8794);
or U8904 (N_8904,N_8676,N_8656);
xnor U8905 (N_8905,N_8669,N_8656);
nor U8906 (N_8906,N_8652,N_8635);
nor U8907 (N_8907,N_8792,N_8619);
and U8908 (N_8908,N_8754,N_8763);
and U8909 (N_8909,N_8737,N_8789);
nor U8910 (N_8910,N_8650,N_8784);
nor U8911 (N_8911,N_8785,N_8736);
nand U8912 (N_8912,N_8669,N_8692);
or U8913 (N_8913,N_8612,N_8724);
nand U8914 (N_8914,N_8701,N_8630);
or U8915 (N_8915,N_8797,N_8777);
or U8916 (N_8916,N_8680,N_8753);
nor U8917 (N_8917,N_8711,N_8612);
or U8918 (N_8918,N_8609,N_8772);
and U8919 (N_8919,N_8735,N_8672);
or U8920 (N_8920,N_8728,N_8725);
xor U8921 (N_8921,N_8724,N_8699);
and U8922 (N_8922,N_8733,N_8784);
or U8923 (N_8923,N_8770,N_8774);
nor U8924 (N_8924,N_8750,N_8650);
nand U8925 (N_8925,N_8774,N_8657);
and U8926 (N_8926,N_8636,N_8762);
xor U8927 (N_8927,N_8742,N_8724);
or U8928 (N_8928,N_8612,N_8652);
xor U8929 (N_8929,N_8726,N_8794);
xor U8930 (N_8930,N_8658,N_8691);
xnor U8931 (N_8931,N_8768,N_8757);
or U8932 (N_8932,N_8697,N_8779);
or U8933 (N_8933,N_8669,N_8649);
nand U8934 (N_8934,N_8751,N_8799);
or U8935 (N_8935,N_8698,N_8678);
nand U8936 (N_8936,N_8670,N_8603);
nor U8937 (N_8937,N_8710,N_8660);
nand U8938 (N_8938,N_8741,N_8701);
nor U8939 (N_8939,N_8743,N_8797);
xnor U8940 (N_8940,N_8725,N_8726);
and U8941 (N_8941,N_8763,N_8790);
and U8942 (N_8942,N_8792,N_8612);
xor U8943 (N_8943,N_8680,N_8701);
nand U8944 (N_8944,N_8674,N_8790);
or U8945 (N_8945,N_8631,N_8619);
xnor U8946 (N_8946,N_8632,N_8609);
xor U8947 (N_8947,N_8698,N_8654);
and U8948 (N_8948,N_8679,N_8621);
or U8949 (N_8949,N_8622,N_8736);
xnor U8950 (N_8950,N_8727,N_8672);
xor U8951 (N_8951,N_8711,N_8610);
nand U8952 (N_8952,N_8647,N_8744);
or U8953 (N_8953,N_8773,N_8739);
or U8954 (N_8954,N_8617,N_8631);
xor U8955 (N_8955,N_8786,N_8784);
nor U8956 (N_8956,N_8670,N_8717);
and U8957 (N_8957,N_8647,N_8600);
and U8958 (N_8958,N_8626,N_8649);
nor U8959 (N_8959,N_8756,N_8698);
nor U8960 (N_8960,N_8704,N_8601);
or U8961 (N_8961,N_8785,N_8796);
or U8962 (N_8962,N_8618,N_8700);
nand U8963 (N_8963,N_8721,N_8779);
nand U8964 (N_8964,N_8658,N_8707);
nand U8965 (N_8965,N_8605,N_8712);
nor U8966 (N_8966,N_8739,N_8716);
and U8967 (N_8967,N_8677,N_8662);
xnor U8968 (N_8968,N_8607,N_8692);
xor U8969 (N_8969,N_8671,N_8646);
or U8970 (N_8970,N_8616,N_8689);
and U8971 (N_8971,N_8758,N_8760);
or U8972 (N_8972,N_8615,N_8682);
and U8973 (N_8973,N_8765,N_8731);
nor U8974 (N_8974,N_8783,N_8684);
and U8975 (N_8975,N_8753,N_8764);
and U8976 (N_8976,N_8629,N_8700);
and U8977 (N_8977,N_8626,N_8666);
nand U8978 (N_8978,N_8764,N_8693);
xor U8979 (N_8979,N_8613,N_8690);
or U8980 (N_8980,N_8628,N_8691);
nand U8981 (N_8981,N_8795,N_8638);
and U8982 (N_8982,N_8685,N_8648);
nand U8983 (N_8983,N_8735,N_8760);
and U8984 (N_8984,N_8648,N_8742);
and U8985 (N_8985,N_8725,N_8781);
nor U8986 (N_8986,N_8618,N_8703);
nand U8987 (N_8987,N_8664,N_8687);
and U8988 (N_8988,N_8607,N_8735);
or U8989 (N_8989,N_8700,N_8706);
and U8990 (N_8990,N_8786,N_8799);
xnor U8991 (N_8991,N_8677,N_8779);
xor U8992 (N_8992,N_8702,N_8690);
xor U8993 (N_8993,N_8616,N_8743);
nor U8994 (N_8994,N_8744,N_8669);
or U8995 (N_8995,N_8732,N_8656);
or U8996 (N_8996,N_8636,N_8601);
nor U8997 (N_8997,N_8610,N_8691);
nor U8998 (N_8998,N_8727,N_8635);
and U8999 (N_8999,N_8649,N_8740);
and U9000 (N_9000,N_8930,N_8870);
nand U9001 (N_9001,N_8827,N_8951);
nand U9002 (N_9002,N_8859,N_8865);
nor U9003 (N_9003,N_8809,N_8824);
xor U9004 (N_9004,N_8835,N_8920);
or U9005 (N_9005,N_8862,N_8852);
or U9006 (N_9006,N_8869,N_8937);
xnor U9007 (N_9007,N_8975,N_8887);
nor U9008 (N_9008,N_8810,N_8800);
or U9009 (N_9009,N_8844,N_8886);
and U9010 (N_9010,N_8861,N_8998);
or U9011 (N_9011,N_8933,N_8897);
nand U9012 (N_9012,N_8899,N_8855);
nand U9013 (N_9013,N_8927,N_8866);
xnor U9014 (N_9014,N_8907,N_8985);
xor U9015 (N_9015,N_8893,N_8945);
nor U9016 (N_9016,N_8939,N_8989);
or U9017 (N_9017,N_8812,N_8890);
xnor U9018 (N_9018,N_8978,N_8884);
and U9019 (N_9019,N_8938,N_8815);
or U9020 (N_9020,N_8949,N_8857);
nor U9021 (N_9021,N_8842,N_8901);
nor U9022 (N_9022,N_8839,N_8950);
nor U9023 (N_9023,N_8993,N_8928);
or U9024 (N_9024,N_8954,N_8801);
xor U9025 (N_9025,N_8996,N_8984);
or U9026 (N_9026,N_8836,N_8878);
xor U9027 (N_9027,N_8995,N_8941);
and U9028 (N_9028,N_8999,N_8896);
nand U9029 (N_9029,N_8988,N_8846);
nor U9030 (N_9030,N_8822,N_8858);
or U9031 (N_9031,N_8931,N_8957);
and U9032 (N_9032,N_8948,N_8850);
nor U9033 (N_9033,N_8911,N_8841);
xor U9034 (N_9034,N_8943,N_8871);
xnor U9035 (N_9035,N_8912,N_8952);
and U9036 (N_9036,N_8924,N_8921);
or U9037 (N_9037,N_8905,N_8906);
nor U9038 (N_9038,N_8838,N_8986);
and U9039 (N_9039,N_8867,N_8940);
xnor U9040 (N_9040,N_8994,N_8923);
or U9041 (N_9041,N_8803,N_8991);
nand U9042 (N_9042,N_8823,N_8942);
and U9043 (N_9043,N_8902,N_8900);
nor U9044 (N_9044,N_8965,N_8864);
and U9045 (N_9045,N_8854,N_8898);
and U9046 (N_9046,N_8992,N_8926);
and U9047 (N_9047,N_8904,N_8817);
or U9048 (N_9048,N_8826,N_8953);
or U9049 (N_9049,N_8935,N_8974);
nor U9050 (N_9050,N_8845,N_8970);
xnor U9051 (N_9051,N_8947,N_8847);
nor U9052 (N_9052,N_8875,N_8971);
or U9053 (N_9053,N_8881,N_8922);
xnor U9054 (N_9054,N_8895,N_8874);
and U9055 (N_9055,N_8888,N_8892);
xor U9056 (N_9056,N_8982,N_8963);
nor U9057 (N_9057,N_8832,N_8972);
nor U9058 (N_9058,N_8833,N_8894);
and U9059 (N_9059,N_8969,N_8880);
or U9060 (N_9060,N_8977,N_8914);
or U9061 (N_9061,N_8849,N_8962);
or U9062 (N_9062,N_8917,N_8932);
nand U9063 (N_9063,N_8925,N_8818);
nor U9064 (N_9064,N_8946,N_8981);
or U9065 (N_9065,N_8851,N_8837);
and U9066 (N_9066,N_8955,N_8910);
xor U9067 (N_9067,N_8856,N_8967);
or U9068 (N_9068,N_8959,N_8879);
nand U9069 (N_9069,N_8909,N_8820);
and U9070 (N_9070,N_8825,N_8868);
xnor U9071 (N_9071,N_8983,N_8811);
nor U9072 (N_9072,N_8819,N_8903);
xnor U9073 (N_9073,N_8990,N_8882);
nor U9074 (N_9074,N_8830,N_8973);
and U9075 (N_9075,N_8891,N_8831);
and U9076 (N_9076,N_8929,N_8936);
or U9077 (N_9077,N_8966,N_8889);
nor U9078 (N_9078,N_8853,N_8872);
nand U9079 (N_9079,N_8848,N_8997);
xor U9080 (N_9080,N_8960,N_8860);
and U9081 (N_9081,N_8873,N_8813);
xnor U9082 (N_9082,N_8968,N_8956);
and U9083 (N_9083,N_8806,N_8961);
nor U9084 (N_9084,N_8915,N_8816);
and U9085 (N_9085,N_8805,N_8828);
and U9086 (N_9086,N_8918,N_8834);
or U9087 (N_9087,N_8821,N_8934);
and U9088 (N_9088,N_8876,N_8807);
nor U9089 (N_9089,N_8843,N_8883);
xnor U9090 (N_9090,N_8808,N_8919);
or U9091 (N_9091,N_8885,N_8829);
nand U9092 (N_9092,N_8958,N_8814);
nor U9093 (N_9093,N_8804,N_8976);
nand U9094 (N_9094,N_8916,N_8802);
nor U9095 (N_9095,N_8944,N_8987);
or U9096 (N_9096,N_8877,N_8908);
nor U9097 (N_9097,N_8964,N_8979);
nor U9098 (N_9098,N_8913,N_8840);
nand U9099 (N_9099,N_8980,N_8863);
and U9100 (N_9100,N_8854,N_8911);
xor U9101 (N_9101,N_8871,N_8925);
and U9102 (N_9102,N_8857,N_8910);
nor U9103 (N_9103,N_8968,N_8907);
xor U9104 (N_9104,N_8908,N_8949);
xnor U9105 (N_9105,N_8995,N_8942);
nor U9106 (N_9106,N_8802,N_8946);
nor U9107 (N_9107,N_8946,N_8970);
xor U9108 (N_9108,N_8911,N_8955);
nand U9109 (N_9109,N_8932,N_8984);
nand U9110 (N_9110,N_8953,N_8801);
and U9111 (N_9111,N_8963,N_8837);
and U9112 (N_9112,N_8996,N_8826);
nand U9113 (N_9113,N_8975,N_8902);
or U9114 (N_9114,N_8872,N_8810);
and U9115 (N_9115,N_8847,N_8823);
and U9116 (N_9116,N_8833,N_8942);
or U9117 (N_9117,N_8895,N_8989);
or U9118 (N_9118,N_8816,N_8985);
and U9119 (N_9119,N_8804,N_8816);
xnor U9120 (N_9120,N_8923,N_8997);
nand U9121 (N_9121,N_8895,N_8976);
and U9122 (N_9122,N_8908,N_8808);
nand U9123 (N_9123,N_8856,N_8992);
or U9124 (N_9124,N_8985,N_8983);
or U9125 (N_9125,N_8964,N_8945);
and U9126 (N_9126,N_8884,N_8898);
and U9127 (N_9127,N_8804,N_8975);
nor U9128 (N_9128,N_8980,N_8978);
xor U9129 (N_9129,N_8931,N_8801);
nor U9130 (N_9130,N_8988,N_8950);
xor U9131 (N_9131,N_8927,N_8935);
or U9132 (N_9132,N_8983,N_8822);
nand U9133 (N_9133,N_8942,N_8864);
nor U9134 (N_9134,N_8873,N_8836);
xnor U9135 (N_9135,N_8827,N_8885);
xor U9136 (N_9136,N_8966,N_8801);
xor U9137 (N_9137,N_8846,N_8975);
nand U9138 (N_9138,N_8919,N_8874);
xor U9139 (N_9139,N_8873,N_8839);
xnor U9140 (N_9140,N_8915,N_8922);
xor U9141 (N_9141,N_8897,N_8805);
nand U9142 (N_9142,N_8989,N_8995);
or U9143 (N_9143,N_8865,N_8995);
and U9144 (N_9144,N_8853,N_8835);
and U9145 (N_9145,N_8992,N_8970);
nand U9146 (N_9146,N_8837,N_8981);
or U9147 (N_9147,N_8981,N_8958);
and U9148 (N_9148,N_8810,N_8894);
and U9149 (N_9149,N_8858,N_8975);
nand U9150 (N_9150,N_8916,N_8957);
nand U9151 (N_9151,N_8803,N_8914);
nand U9152 (N_9152,N_8962,N_8880);
nor U9153 (N_9153,N_8854,N_8909);
nor U9154 (N_9154,N_8807,N_8865);
xnor U9155 (N_9155,N_8953,N_8901);
and U9156 (N_9156,N_8991,N_8859);
and U9157 (N_9157,N_8872,N_8859);
and U9158 (N_9158,N_8861,N_8860);
nor U9159 (N_9159,N_8934,N_8880);
and U9160 (N_9160,N_8862,N_8920);
and U9161 (N_9161,N_8927,N_8832);
xor U9162 (N_9162,N_8874,N_8872);
nand U9163 (N_9163,N_8852,N_8878);
xor U9164 (N_9164,N_8807,N_8874);
and U9165 (N_9165,N_8971,N_8855);
or U9166 (N_9166,N_8809,N_8960);
or U9167 (N_9167,N_8872,N_8961);
nand U9168 (N_9168,N_8944,N_8839);
or U9169 (N_9169,N_8803,N_8998);
nor U9170 (N_9170,N_8933,N_8856);
or U9171 (N_9171,N_8961,N_8852);
xor U9172 (N_9172,N_8890,N_8914);
and U9173 (N_9173,N_8936,N_8874);
nand U9174 (N_9174,N_8952,N_8943);
nor U9175 (N_9175,N_8981,N_8913);
or U9176 (N_9176,N_8879,N_8923);
xor U9177 (N_9177,N_8855,N_8834);
nor U9178 (N_9178,N_8960,N_8987);
and U9179 (N_9179,N_8877,N_8981);
or U9180 (N_9180,N_8896,N_8914);
or U9181 (N_9181,N_8832,N_8910);
nor U9182 (N_9182,N_8942,N_8978);
xnor U9183 (N_9183,N_8952,N_8951);
or U9184 (N_9184,N_8950,N_8896);
and U9185 (N_9185,N_8976,N_8886);
xnor U9186 (N_9186,N_8991,N_8989);
and U9187 (N_9187,N_8860,N_8986);
or U9188 (N_9188,N_8919,N_8884);
or U9189 (N_9189,N_8861,N_8985);
xnor U9190 (N_9190,N_8986,N_8815);
nand U9191 (N_9191,N_8862,N_8992);
nand U9192 (N_9192,N_8804,N_8981);
and U9193 (N_9193,N_8887,N_8993);
nand U9194 (N_9194,N_8951,N_8980);
nor U9195 (N_9195,N_8968,N_8871);
nor U9196 (N_9196,N_8948,N_8999);
xnor U9197 (N_9197,N_8867,N_8999);
nor U9198 (N_9198,N_8803,N_8844);
nand U9199 (N_9199,N_8858,N_8819);
or U9200 (N_9200,N_9094,N_9135);
or U9201 (N_9201,N_9052,N_9139);
xor U9202 (N_9202,N_9018,N_9141);
xnor U9203 (N_9203,N_9132,N_9169);
nor U9204 (N_9204,N_9030,N_9190);
and U9205 (N_9205,N_9066,N_9105);
nor U9206 (N_9206,N_9024,N_9186);
or U9207 (N_9207,N_9173,N_9022);
and U9208 (N_9208,N_9187,N_9163);
nor U9209 (N_9209,N_9008,N_9060);
nand U9210 (N_9210,N_9082,N_9128);
nand U9211 (N_9211,N_9111,N_9110);
xnor U9212 (N_9212,N_9087,N_9177);
nand U9213 (N_9213,N_9154,N_9062);
nand U9214 (N_9214,N_9080,N_9119);
nand U9215 (N_9215,N_9003,N_9100);
and U9216 (N_9216,N_9027,N_9140);
or U9217 (N_9217,N_9101,N_9007);
or U9218 (N_9218,N_9120,N_9109);
xnor U9219 (N_9219,N_9172,N_9099);
xnor U9220 (N_9220,N_9175,N_9193);
nand U9221 (N_9221,N_9155,N_9189);
or U9222 (N_9222,N_9164,N_9199);
nand U9223 (N_9223,N_9181,N_9061);
nor U9224 (N_9224,N_9002,N_9151);
nand U9225 (N_9225,N_9038,N_9084);
nor U9226 (N_9226,N_9058,N_9176);
or U9227 (N_9227,N_9166,N_9083);
nor U9228 (N_9228,N_9108,N_9106);
xor U9229 (N_9229,N_9170,N_9016);
or U9230 (N_9230,N_9095,N_9075);
nor U9231 (N_9231,N_9138,N_9197);
nand U9232 (N_9232,N_9015,N_9157);
xnor U9233 (N_9233,N_9019,N_9188);
nor U9234 (N_9234,N_9085,N_9160);
and U9235 (N_9235,N_9045,N_9179);
or U9236 (N_9236,N_9073,N_9171);
nand U9237 (N_9237,N_9035,N_9156);
nor U9238 (N_9238,N_9009,N_9092);
xor U9239 (N_9239,N_9043,N_9020);
nor U9240 (N_9240,N_9049,N_9134);
nor U9241 (N_9241,N_9097,N_9098);
nand U9242 (N_9242,N_9126,N_9137);
nand U9243 (N_9243,N_9127,N_9077);
nand U9244 (N_9244,N_9129,N_9053);
and U9245 (N_9245,N_9167,N_9112);
xnor U9246 (N_9246,N_9054,N_9124);
or U9247 (N_9247,N_9150,N_9072);
nor U9248 (N_9248,N_9182,N_9042);
or U9249 (N_9249,N_9068,N_9192);
and U9250 (N_9250,N_9034,N_9162);
nor U9251 (N_9251,N_9076,N_9089);
and U9252 (N_9252,N_9194,N_9051);
xnor U9253 (N_9253,N_9044,N_9021);
and U9254 (N_9254,N_9004,N_9136);
nor U9255 (N_9255,N_9057,N_9103);
nand U9256 (N_9256,N_9158,N_9130);
and U9257 (N_9257,N_9116,N_9107);
and U9258 (N_9258,N_9168,N_9183);
and U9259 (N_9259,N_9064,N_9050);
and U9260 (N_9260,N_9113,N_9196);
nor U9261 (N_9261,N_9055,N_9131);
nor U9262 (N_9262,N_9104,N_9037);
xnor U9263 (N_9263,N_9153,N_9174);
xor U9264 (N_9264,N_9031,N_9025);
and U9265 (N_9265,N_9148,N_9033);
or U9266 (N_9266,N_9198,N_9102);
nand U9267 (N_9267,N_9001,N_9056);
xnor U9268 (N_9268,N_9178,N_9159);
and U9269 (N_9269,N_9152,N_9133);
xnor U9270 (N_9270,N_9046,N_9145);
nor U9271 (N_9271,N_9059,N_9115);
or U9272 (N_9272,N_9028,N_9040);
or U9273 (N_9273,N_9091,N_9195);
or U9274 (N_9274,N_9191,N_9142);
nand U9275 (N_9275,N_9041,N_9017);
nand U9276 (N_9276,N_9000,N_9088);
and U9277 (N_9277,N_9123,N_9165);
xor U9278 (N_9278,N_9014,N_9065);
nor U9279 (N_9279,N_9185,N_9122);
nand U9280 (N_9280,N_9023,N_9074);
and U9281 (N_9281,N_9070,N_9117);
xor U9282 (N_9282,N_9063,N_9032);
nor U9283 (N_9283,N_9149,N_9144);
and U9284 (N_9284,N_9005,N_9026);
nand U9285 (N_9285,N_9093,N_9039);
xor U9286 (N_9286,N_9114,N_9180);
nand U9287 (N_9287,N_9096,N_9121);
nor U9288 (N_9288,N_9013,N_9047);
and U9289 (N_9289,N_9079,N_9036);
and U9290 (N_9290,N_9078,N_9086);
xnor U9291 (N_9291,N_9081,N_9006);
nor U9292 (N_9292,N_9069,N_9029);
nor U9293 (N_9293,N_9067,N_9161);
or U9294 (N_9294,N_9011,N_9146);
xor U9295 (N_9295,N_9147,N_9012);
and U9296 (N_9296,N_9125,N_9143);
nor U9297 (N_9297,N_9048,N_9071);
or U9298 (N_9298,N_9118,N_9090);
nor U9299 (N_9299,N_9010,N_9184);
nand U9300 (N_9300,N_9107,N_9097);
or U9301 (N_9301,N_9082,N_9148);
xnor U9302 (N_9302,N_9085,N_9002);
and U9303 (N_9303,N_9182,N_9004);
nor U9304 (N_9304,N_9073,N_9122);
and U9305 (N_9305,N_9191,N_9140);
nor U9306 (N_9306,N_9084,N_9149);
nor U9307 (N_9307,N_9167,N_9129);
nand U9308 (N_9308,N_9184,N_9112);
or U9309 (N_9309,N_9176,N_9191);
or U9310 (N_9310,N_9118,N_9146);
xor U9311 (N_9311,N_9091,N_9197);
xnor U9312 (N_9312,N_9069,N_9197);
nor U9313 (N_9313,N_9111,N_9180);
or U9314 (N_9314,N_9109,N_9052);
and U9315 (N_9315,N_9033,N_9121);
or U9316 (N_9316,N_9108,N_9144);
xnor U9317 (N_9317,N_9163,N_9045);
nor U9318 (N_9318,N_9132,N_9063);
and U9319 (N_9319,N_9069,N_9118);
nor U9320 (N_9320,N_9091,N_9043);
nand U9321 (N_9321,N_9195,N_9128);
nand U9322 (N_9322,N_9111,N_9160);
nand U9323 (N_9323,N_9143,N_9190);
xnor U9324 (N_9324,N_9172,N_9006);
or U9325 (N_9325,N_9158,N_9161);
nor U9326 (N_9326,N_9128,N_9126);
xnor U9327 (N_9327,N_9054,N_9008);
xor U9328 (N_9328,N_9073,N_9160);
and U9329 (N_9329,N_9029,N_9003);
nand U9330 (N_9330,N_9145,N_9156);
xnor U9331 (N_9331,N_9029,N_9022);
nand U9332 (N_9332,N_9159,N_9057);
nand U9333 (N_9333,N_9044,N_9150);
or U9334 (N_9334,N_9194,N_9047);
xor U9335 (N_9335,N_9180,N_9177);
nand U9336 (N_9336,N_9195,N_9160);
and U9337 (N_9337,N_9157,N_9072);
or U9338 (N_9338,N_9089,N_9126);
xnor U9339 (N_9339,N_9195,N_9130);
nor U9340 (N_9340,N_9065,N_9019);
nand U9341 (N_9341,N_9161,N_9185);
nor U9342 (N_9342,N_9040,N_9162);
nand U9343 (N_9343,N_9187,N_9169);
or U9344 (N_9344,N_9111,N_9127);
nand U9345 (N_9345,N_9177,N_9101);
and U9346 (N_9346,N_9027,N_9122);
nor U9347 (N_9347,N_9087,N_9019);
xor U9348 (N_9348,N_9150,N_9028);
and U9349 (N_9349,N_9096,N_9117);
nand U9350 (N_9350,N_9011,N_9139);
and U9351 (N_9351,N_9118,N_9107);
nand U9352 (N_9352,N_9070,N_9041);
or U9353 (N_9353,N_9116,N_9022);
or U9354 (N_9354,N_9041,N_9046);
or U9355 (N_9355,N_9039,N_9136);
or U9356 (N_9356,N_9075,N_9053);
nor U9357 (N_9357,N_9108,N_9093);
and U9358 (N_9358,N_9023,N_9142);
nand U9359 (N_9359,N_9124,N_9078);
and U9360 (N_9360,N_9067,N_9125);
or U9361 (N_9361,N_9095,N_9166);
nor U9362 (N_9362,N_9100,N_9035);
and U9363 (N_9363,N_9026,N_9190);
nand U9364 (N_9364,N_9039,N_9160);
or U9365 (N_9365,N_9071,N_9062);
nor U9366 (N_9366,N_9088,N_9180);
and U9367 (N_9367,N_9080,N_9034);
nor U9368 (N_9368,N_9132,N_9059);
nor U9369 (N_9369,N_9000,N_9179);
nor U9370 (N_9370,N_9170,N_9103);
nor U9371 (N_9371,N_9052,N_9189);
nand U9372 (N_9372,N_9109,N_9150);
nand U9373 (N_9373,N_9175,N_9083);
xnor U9374 (N_9374,N_9059,N_9190);
nand U9375 (N_9375,N_9176,N_9121);
or U9376 (N_9376,N_9152,N_9173);
or U9377 (N_9377,N_9130,N_9155);
and U9378 (N_9378,N_9137,N_9164);
nor U9379 (N_9379,N_9193,N_9027);
or U9380 (N_9380,N_9085,N_9080);
and U9381 (N_9381,N_9018,N_9098);
or U9382 (N_9382,N_9185,N_9112);
or U9383 (N_9383,N_9043,N_9108);
and U9384 (N_9384,N_9174,N_9166);
nor U9385 (N_9385,N_9114,N_9089);
nand U9386 (N_9386,N_9199,N_9065);
and U9387 (N_9387,N_9019,N_9086);
or U9388 (N_9388,N_9194,N_9164);
or U9389 (N_9389,N_9001,N_9089);
xnor U9390 (N_9390,N_9176,N_9104);
nand U9391 (N_9391,N_9082,N_9109);
xnor U9392 (N_9392,N_9011,N_9088);
or U9393 (N_9393,N_9105,N_9182);
or U9394 (N_9394,N_9084,N_9144);
xnor U9395 (N_9395,N_9030,N_9147);
or U9396 (N_9396,N_9185,N_9128);
xor U9397 (N_9397,N_9051,N_9193);
nor U9398 (N_9398,N_9113,N_9002);
and U9399 (N_9399,N_9177,N_9110);
or U9400 (N_9400,N_9243,N_9315);
or U9401 (N_9401,N_9391,N_9353);
nand U9402 (N_9402,N_9258,N_9218);
xnor U9403 (N_9403,N_9381,N_9282);
nand U9404 (N_9404,N_9328,N_9200);
xnor U9405 (N_9405,N_9370,N_9375);
nor U9406 (N_9406,N_9257,N_9244);
nand U9407 (N_9407,N_9389,N_9277);
xnor U9408 (N_9408,N_9351,N_9354);
xor U9409 (N_9409,N_9209,N_9227);
and U9410 (N_9410,N_9260,N_9206);
and U9411 (N_9411,N_9372,N_9398);
nand U9412 (N_9412,N_9291,N_9284);
and U9413 (N_9413,N_9306,N_9292);
nand U9414 (N_9414,N_9390,N_9300);
nand U9415 (N_9415,N_9376,N_9274);
nand U9416 (N_9416,N_9270,N_9216);
nor U9417 (N_9417,N_9271,N_9297);
xor U9418 (N_9418,N_9397,N_9288);
xnor U9419 (N_9419,N_9302,N_9343);
xnor U9420 (N_9420,N_9323,N_9210);
nor U9421 (N_9421,N_9326,N_9380);
nand U9422 (N_9422,N_9252,N_9399);
and U9423 (N_9423,N_9336,N_9232);
and U9424 (N_9424,N_9221,N_9369);
xnor U9425 (N_9425,N_9382,N_9269);
xnor U9426 (N_9426,N_9267,N_9395);
nor U9427 (N_9427,N_9347,N_9251);
and U9428 (N_9428,N_9374,N_9239);
nor U9429 (N_9429,N_9219,N_9309);
nand U9430 (N_9430,N_9314,N_9246);
xor U9431 (N_9431,N_9341,N_9366);
and U9432 (N_9432,N_9394,N_9331);
nand U9433 (N_9433,N_9261,N_9237);
nor U9434 (N_9434,N_9259,N_9342);
xnor U9435 (N_9435,N_9281,N_9253);
and U9436 (N_9436,N_9355,N_9283);
xor U9437 (N_9437,N_9208,N_9329);
nand U9438 (N_9438,N_9396,N_9339);
nor U9439 (N_9439,N_9305,N_9363);
or U9440 (N_9440,N_9320,N_9255);
xor U9441 (N_9441,N_9350,N_9346);
and U9442 (N_9442,N_9308,N_9265);
nand U9443 (N_9443,N_9304,N_9276);
and U9444 (N_9444,N_9358,N_9280);
xnor U9445 (N_9445,N_9290,N_9201);
nand U9446 (N_9446,N_9325,N_9334);
xor U9447 (N_9447,N_9245,N_9362);
nor U9448 (N_9448,N_9316,N_9324);
nor U9449 (N_9449,N_9371,N_9225);
xor U9450 (N_9450,N_9337,N_9321);
xnor U9451 (N_9451,N_9333,N_9330);
xnor U9452 (N_9452,N_9234,N_9286);
nand U9453 (N_9453,N_9217,N_9377);
and U9454 (N_9454,N_9357,N_9263);
and U9455 (N_9455,N_9213,N_9240);
xnor U9456 (N_9456,N_9338,N_9272);
and U9457 (N_9457,N_9236,N_9360);
nand U9458 (N_9458,N_9349,N_9344);
or U9459 (N_9459,N_9295,N_9298);
nand U9460 (N_9460,N_9311,N_9268);
nand U9461 (N_9461,N_9310,N_9254);
nand U9462 (N_9462,N_9299,N_9289);
nor U9463 (N_9463,N_9278,N_9285);
or U9464 (N_9464,N_9296,N_9242);
nand U9465 (N_9465,N_9204,N_9365);
nand U9466 (N_9466,N_9359,N_9238);
nor U9467 (N_9467,N_9250,N_9224);
or U9468 (N_9468,N_9207,N_9279);
nand U9469 (N_9469,N_9256,N_9222);
nor U9470 (N_9470,N_9312,N_9262);
nand U9471 (N_9471,N_9214,N_9220);
nor U9472 (N_9472,N_9388,N_9229);
nand U9473 (N_9473,N_9340,N_9223);
xnor U9474 (N_9474,N_9383,N_9335);
or U9475 (N_9475,N_9228,N_9212);
nand U9476 (N_9476,N_9384,N_9235);
nor U9477 (N_9477,N_9327,N_9273);
and U9478 (N_9478,N_9367,N_9303);
and U9479 (N_9479,N_9313,N_9202);
xnor U9480 (N_9480,N_9247,N_9352);
and U9481 (N_9481,N_9248,N_9231);
and U9482 (N_9482,N_9249,N_9364);
nor U9483 (N_9483,N_9294,N_9215);
or U9484 (N_9484,N_9266,N_9307);
nor U9485 (N_9485,N_9287,N_9203);
xor U9486 (N_9486,N_9322,N_9368);
xor U9487 (N_9487,N_9378,N_9345);
xnor U9488 (N_9488,N_9319,N_9387);
xnor U9489 (N_9489,N_9293,N_9356);
or U9490 (N_9490,N_9241,N_9385);
or U9491 (N_9491,N_9275,N_9386);
and U9492 (N_9492,N_9230,N_9205);
nand U9493 (N_9493,N_9361,N_9393);
and U9494 (N_9494,N_9392,N_9301);
and U9495 (N_9495,N_9379,N_9211);
nand U9496 (N_9496,N_9317,N_9373);
and U9497 (N_9497,N_9332,N_9264);
nor U9498 (N_9498,N_9318,N_9226);
or U9499 (N_9499,N_9348,N_9233);
and U9500 (N_9500,N_9203,N_9204);
or U9501 (N_9501,N_9269,N_9229);
xor U9502 (N_9502,N_9300,N_9291);
nor U9503 (N_9503,N_9211,N_9371);
xnor U9504 (N_9504,N_9343,N_9206);
nor U9505 (N_9505,N_9368,N_9251);
and U9506 (N_9506,N_9359,N_9232);
or U9507 (N_9507,N_9381,N_9389);
and U9508 (N_9508,N_9378,N_9363);
nor U9509 (N_9509,N_9324,N_9273);
and U9510 (N_9510,N_9291,N_9311);
or U9511 (N_9511,N_9320,N_9326);
xor U9512 (N_9512,N_9351,N_9287);
xor U9513 (N_9513,N_9395,N_9215);
nor U9514 (N_9514,N_9214,N_9327);
nand U9515 (N_9515,N_9321,N_9368);
xnor U9516 (N_9516,N_9239,N_9264);
nor U9517 (N_9517,N_9240,N_9261);
xnor U9518 (N_9518,N_9385,N_9380);
or U9519 (N_9519,N_9279,N_9264);
or U9520 (N_9520,N_9228,N_9287);
and U9521 (N_9521,N_9206,N_9374);
nor U9522 (N_9522,N_9257,N_9317);
nor U9523 (N_9523,N_9285,N_9258);
xor U9524 (N_9524,N_9224,N_9253);
or U9525 (N_9525,N_9302,N_9336);
nor U9526 (N_9526,N_9271,N_9368);
nand U9527 (N_9527,N_9270,N_9294);
and U9528 (N_9528,N_9364,N_9350);
nor U9529 (N_9529,N_9283,N_9319);
and U9530 (N_9530,N_9388,N_9321);
xnor U9531 (N_9531,N_9261,N_9337);
nand U9532 (N_9532,N_9235,N_9380);
nand U9533 (N_9533,N_9253,N_9284);
nand U9534 (N_9534,N_9397,N_9205);
nand U9535 (N_9535,N_9298,N_9312);
or U9536 (N_9536,N_9286,N_9316);
and U9537 (N_9537,N_9200,N_9355);
nor U9538 (N_9538,N_9290,N_9316);
nand U9539 (N_9539,N_9332,N_9288);
and U9540 (N_9540,N_9317,N_9300);
nand U9541 (N_9541,N_9277,N_9366);
and U9542 (N_9542,N_9360,N_9359);
and U9543 (N_9543,N_9207,N_9209);
nand U9544 (N_9544,N_9383,N_9390);
or U9545 (N_9545,N_9380,N_9310);
nand U9546 (N_9546,N_9312,N_9359);
or U9547 (N_9547,N_9322,N_9397);
xnor U9548 (N_9548,N_9224,N_9258);
nor U9549 (N_9549,N_9369,N_9350);
nand U9550 (N_9550,N_9346,N_9223);
nand U9551 (N_9551,N_9235,N_9285);
nand U9552 (N_9552,N_9273,N_9336);
or U9553 (N_9553,N_9257,N_9276);
and U9554 (N_9554,N_9361,N_9275);
nor U9555 (N_9555,N_9258,N_9335);
nand U9556 (N_9556,N_9273,N_9267);
xnor U9557 (N_9557,N_9206,N_9266);
or U9558 (N_9558,N_9314,N_9287);
xnor U9559 (N_9559,N_9383,N_9317);
and U9560 (N_9560,N_9228,N_9396);
xnor U9561 (N_9561,N_9328,N_9209);
nor U9562 (N_9562,N_9232,N_9287);
or U9563 (N_9563,N_9324,N_9315);
or U9564 (N_9564,N_9279,N_9249);
xnor U9565 (N_9565,N_9279,N_9353);
and U9566 (N_9566,N_9349,N_9351);
xor U9567 (N_9567,N_9354,N_9213);
nand U9568 (N_9568,N_9290,N_9247);
and U9569 (N_9569,N_9378,N_9303);
nand U9570 (N_9570,N_9338,N_9286);
and U9571 (N_9571,N_9259,N_9200);
xor U9572 (N_9572,N_9237,N_9343);
nand U9573 (N_9573,N_9301,N_9321);
nor U9574 (N_9574,N_9209,N_9346);
nand U9575 (N_9575,N_9322,N_9330);
xor U9576 (N_9576,N_9392,N_9399);
nand U9577 (N_9577,N_9336,N_9247);
nand U9578 (N_9578,N_9398,N_9229);
nor U9579 (N_9579,N_9383,N_9204);
xnor U9580 (N_9580,N_9296,N_9229);
xor U9581 (N_9581,N_9227,N_9239);
xnor U9582 (N_9582,N_9249,N_9354);
nand U9583 (N_9583,N_9235,N_9334);
nand U9584 (N_9584,N_9211,N_9320);
and U9585 (N_9585,N_9330,N_9203);
and U9586 (N_9586,N_9226,N_9240);
nand U9587 (N_9587,N_9282,N_9380);
or U9588 (N_9588,N_9281,N_9303);
and U9589 (N_9589,N_9327,N_9267);
or U9590 (N_9590,N_9376,N_9371);
nor U9591 (N_9591,N_9381,N_9336);
and U9592 (N_9592,N_9328,N_9246);
nand U9593 (N_9593,N_9321,N_9328);
or U9594 (N_9594,N_9395,N_9270);
nand U9595 (N_9595,N_9343,N_9321);
or U9596 (N_9596,N_9363,N_9371);
nand U9597 (N_9597,N_9383,N_9309);
nor U9598 (N_9598,N_9211,N_9324);
nor U9599 (N_9599,N_9237,N_9361);
nor U9600 (N_9600,N_9540,N_9521);
nand U9601 (N_9601,N_9506,N_9586);
xor U9602 (N_9602,N_9446,N_9522);
nor U9603 (N_9603,N_9460,N_9411);
nor U9604 (N_9604,N_9577,N_9588);
xnor U9605 (N_9605,N_9517,N_9556);
xnor U9606 (N_9606,N_9579,N_9409);
and U9607 (N_9607,N_9596,N_9476);
and U9608 (N_9608,N_9524,N_9499);
nor U9609 (N_9609,N_9491,N_9430);
and U9610 (N_9610,N_9481,N_9544);
nor U9611 (N_9611,N_9508,N_9494);
or U9612 (N_9612,N_9450,N_9572);
xor U9613 (N_9613,N_9578,N_9501);
nor U9614 (N_9614,N_9543,N_9449);
nand U9615 (N_9615,N_9583,N_9441);
nor U9616 (N_9616,N_9545,N_9551);
nor U9617 (N_9617,N_9502,N_9598);
and U9618 (N_9618,N_9439,N_9538);
xor U9619 (N_9619,N_9483,N_9550);
and U9620 (N_9620,N_9554,N_9564);
xor U9621 (N_9621,N_9454,N_9589);
and U9622 (N_9622,N_9492,N_9420);
nor U9623 (N_9623,N_9519,N_9487);
and U9624 (N_9624,N_9473,N_9537);
or U9625 (N_9625,N_9470,N_9448);
xnor U9626 (N_9626,N_9489,N_9552);
nand U9627 (N_9627,N_9488,N_9436);
nor U9628 (N_9628,N_9423,N_9528);
nor U9629 (N_9629,N_9595,N_9558);
xor U9630 (N_9630,N_9445,N_9584);
nor U9631 (N_9631,N_9591,N_9523);
nor U9632 (N_9632,N_9412,N_9443);
nand U9633 (N_9633,N_9425,N_9469);
nor U9634 (N_9634,N_9472,N_9404);
and U9635 (N_9635,N_9510,N_9582);
nand U9636 (N_9636,N_9533,N_9576);
or U9637 (N_9637,N_9566,N_9464);
or U9638 (N_9638,N_9474,N_9532);
nand U9639 (N_9639,N_9453,N_9580);
nand U9640 (N_9640,N_9590,N_9416);
nor U9641 (N_9641,N_9490,N_9403);
and U9642 (N_9642,N_9479,N_9475);
or U9643 (N_9643,N_9563,N_9512);
or U9644 (N_9644,N_9536,N_9561);
xor U9645 (N_9645,N_9539,N_9568);
nor U9646 (N_9646,N_9400,N_9426);
nor U9647 (N_9647,N_9465,N_9593);
and U9648 (N_9648,N_9547,N_9431);
nand U9649 (N_9649,N_9432,N_9405);
nor U9650 (N_9650,N_9562,N_9452);
and U9651 (N_9651,N_9503,N_9511);
or U9652 (N_9652,N_9505,N_9569);
xnor U9653 (N_9653,N_9567,N_9429);
or U9654 (N_9654,N_9406,N_9557);
and U9655 (N_9655,N_9407,N_9520);
nand U9656 (N_9656,N_9574,N_9451);
or U9657 (N_9657,N_9534,N_9471);
and U9658 (N_9658,N_9509,N_9486);
or U9659 (N_9659,N_9535,N_9581);
nand U9660 (N_9660,N_9437,N_9427);
xor U9661 (N_9661,N_9455,N_9599);
nand U9662 (N_9662,N_9456,N_9419);
or U9663 (N_9663,N_9447,N_9482);
or U9664 (N_9664,N_9594,N_9413);
nand U9665 (N_9665,N_9442,N_9478);
xnor U9666 (N_9666,N_9500,N_9434);
nor U9667 (N_9667,N_9458,N_9485);
xor U9668 (N_9668,N_9457,N_9548);
or U9669 (N_9669,N_9559,N_9560);
or U9670 (N_9670,N_9422,N_9497);
xor U9671 (N_9671,N_9440,N_9504);
nor U9672 (N_9672,N_9575,N_9592);
or U9673 (N_9673,N_9438,N_9462);
nor U9674 (N_9674,N_9415,N_9461);
nor U9675 (N_9675,N_9480,N_9424);
nand U9676 (N_9676,N_9421,N_9477);
xor U9677 (N_9677,N_9514,N_9515);
and U9678 (N_9678,N_9467,N_9546);
nor U9679 (N_9679,N_9565,N_9418);
or U9680 (N_9680,N_9433,N_9529);
xor U9681 (N_9681,N_9507,N_9527);
or U9682 (N_9682,N_9541,N_9402);
or U9683 (N_9683,N_9463,N_9498);
and U9684 (N_9684,N_9444,N_9526);
nor U9685 (N_9685,N_9597,N_9496);
or U9686 (N_9686,N_9401,N_9531);
nor U9687 (N_9687,N_9518,N_9571);
and U9688 (N_9688,N_9435,N_9459);
xnor U9689 (N_9689,N_9408,N_9428);
or U9690 (N_9690,N_9468,N_9553);
nand U9691 (N_9691,N_9525,N_9410);
or U9692 (N_9692,N_9484,N_9542);
and U9693 (N_9693,N_9549,N_9466);
nor U9694 (N_9694,N_9495,N_9530);
nand U9695 (N_9695,N_9513,N_9555);
xor U9696 (N_9696,N_9587,N_9414);
and U9697 (N_9697,N_9573,N_9570);
xor U9698 (N_9698,N_9493,N_9417);
nand U9699 (N_9699,N_9585,N_9516);
or U9700 (N_9700,N_9473,N_9453);
nand U9701 (N_9701,N_9404,N_9403);
xor U9702 (N_9702,N_9408,N_9575);
and U9703 (N_9703,N_9518,N_9489);
nor U9704 (N_9704,N_9453,N_9461);
or U9705 (N_9705,N_9439,N_9506);
xor U9706 (N_9706,N_9467,N_9570);
and U9707 (N_9707,N_9474,N_9455);
and U9708 (N_9708,N_9572,N_9467);
and U9709 (N_9709,N_9475,N_9543);
xor U9710 (N_9710,N_9472,N_9597);
or U9711 (N_9711,N_9594,N_9459);
xor U9712 (N_9712,N_9582,N_9515);
nor U9713 (N_9713,N_9478,N_9435);
or U9714 (N_9714,N_9460,N_9512);
nand U9715 (N_9715,N_9401,N_9446);
and U9716 (N_9716,N_9461,N_9480);
nor U9717 (N_9717,N_9568,N_9557);
nand U9718 (N_9718,N_9442,N_9537);
nor U9719 (N_9719,N_9401,N_9530);
xor U9720 (N_9720,N_9428,N_9543);
or U9721 (N_9721,N_9540,N_9494);
nor U9722 (N_9722,N_9469,N_9458);
nor U9723 (N_9723,N_9424,N_9596);
nor U9724 (N_9724,N_9480,N_9486);
or U9725 (N_9725,N_9533,N_9588);
nand U9726 (N_9726,N_9524,N_9577);
or U9727 (N_9727,N_9597,N_9566);
nand U9728 (N_9728,N_9593,N_9597);
nor U9729 (N_9729,N_9471,N_9521);
and U9730 (N_9730,N_9456,N_9572);
and U9731 (N_9731,N_9548,N_9402);
nor U9732 (N_9732,N_9439,N_9541);
xnor U9733 (N_9733,N_9543,N_9546);
and U9734 (N_9734,N_9413,N_9515);
or U9735 (N_9735,N_9453,N_9412);
nor U9736 (N_9736,N_9431,N_9553);
and U9737 (N_9737,N_9535,N_9571);
nand U9738 (N_9738,N_9555,N_9435);
nor U9739 (N_9739,N_9424,N_9529);
or U9740 (N_9740,N_9555,N_9451);
and U9741 (N_9741,N_9526,N_9558);
xor U9742 (N_9742,N_9428,N_9597);
and U9743 (N_9743,N_9559,N_9434);
xnor U9744 (N_9744,N_9589,N_9565);
nand U9745 (N_9745,N_9460,N_9456);
nand U9746 (N_9746,N_9589,N_9528);
nor U9747 (N_9747,N_9559,N_9413);
or U9748 (N_9748,N_9567,N_9444);
or U9749 (N_9749,N_9421,N_9554);
nor U9750 (N_9750,N_9518,N_9525);
or U9751 (N_9751,N_9451,N_9507);
nor U9752 (N_9752,N_9469,N_9416);
nor U9753 (N_9753,N_9528,N_9512);
or U9754 (N_9754,N_9414,N_9446);
nor U9755 (N_9755,N_9451,N_9580);
or U9756 (N_9756,N_9405,N_9426);
nor U9757 (N_9757,N_9475,N_9566);
and U9758 (N_9758,N_9401,N_9454);
and U9759 (N_9759,N_9468,N_9409);
and U9760 (N_9760,N_9508,N_9409);
xor U9761 (N_9761,N_9440,N_9487);
or U9762 (N_9762,N_9564,N_9531);
nand U9763 (N_9763,N_9417,N_9418);
and U9764 (N_9764,N_9597,N_9583);
xor U9765 (N_9765,N_9584,N_9506);
nand U9766 (N_9766,N_9441,N_9505);
and U9767 (N_9767,N_9575,N_9423);
and U9768 (N_9768,N_9584,N_9552);
xor U9769 (N_9769,N_9400,N_9527);
and U9770 (N_9770,N_9531,N_9581);
xor U9771 (N_9771,N_9552,N_9441);
nand U9772 (N_9772,N_9465,N_9537);
xor U9773 (N_9773,N_9541,N_9566);
nand U9774 (N_9774,N_9416,N_9404);
nor U9775 (N_9775,N_9523,N_9518);
nand U9776 (N_9776,N_9467,N_9523);
and U9777 (N_9777,N_9453,N_9584);
nor U9778 (N_9778,N_9418,N_9534);
nand U9779 (N_9779,N_9456,N_9488);
xor U9780 (N_9780,N_9401,N_9475);
and U9781 (N_9781,N_9537,N_9514);
xnor U9782 (N_9782,N_9573,N_9417);
xor U9783 (N_9783,N_9508,N_9418);
nor U9784 (N_9784,N_9447,N_9401);
or U9785 (N_9785,N_9596,N_9505);
xnor U9786 (N_9786,N_9476,N_9530);
nor U9787 (N_9787,N_9501,N_9421);
xor U9788 (N_9788,N_9430,N_9417);
nor U9789 (N_9789,N_9566,N_9418);
nor U9790 (N_9790,N_9461,N_9499);
nand U9791 (N_9791,N_9568,N_9460);
xnor U9792 (N_9792,N_9411,N_9579);
xnor U9793 (N_9793,N_9565,N_9555);
or U9794 (N_9794,N_9456,N_9489);
or U9795 (N_9795,N_9423,N_9480);
or U9796 (N_9796,N_9449,N_9595);
or U9797 (N_9797,N_9472,N_9483);
or U9798 (N_9798,N_9445,N_9554);
and U9799 (N_9799,N_9424,N_9525);
or U9800 (N_9800,N_9760,N_9692);
xor U9801 (N_9801,N_9689,N_9677);
xnor U9802 (N_9802,N_9673,N_9682);
and U9803 (N_9803,N_9762,N_9748);
nand U9804 (N_9804,N_9759,N_9742);
nand U9805 (N_9805,N_9603,N_9707);
and U9806 (N_9806,N_9764,N_9691);
and U9807 (N_9807,N_9661,N_9662);
nor U9808 (N_9808,N_9758,N_9785);
nor U9809 (N_9809,N_9700,N_9616);
and U9810 (N_9810,N_9714,N_9668);
nor U9811 (N_9811,N_9670,N_9724);
xor U9812 (N_9812,N_9791,N_9610);
nor U9813 (N_9813,N_9629,N_9732);
nor U9814 (N_9814,N_9617,N_9765);
and U9815 (N_9815,N_9619,N_9751);
or U9816 (N_9816,N_9740,N_9600);
and U9817 (N_9817,N_9693,N_9623);
nand U9818 (N_9818,N_9776,N_9667);
or U9819 (N_9819,N_9731,N_9716);
xnor U9820 (N_9820,N_9701,N_9757);
xnor U9821 (N_9821,N_9719,N_9672);
and U9822 (N_9822,N_9796,N_9747);
xnor U9823 (N_9823,N_9695,N_9710);
nor U9824 (N_9824,N_9763,N_9637);
nand U9825 (N_9825,N_9643,N_9660);
or U9826 (N_9826,N_9717,N_9745);
nor U9827 (N_9827,N_9620,N_9681);
xor U9828 (N_9828,N_9606,N_9605);
nor U9829 (N_9829,N_9743,N_9738);
nor U9830 (N_9830,N_9683,N_9646);
nand U9831 (N_9831,N_9651,N_9644);
or U9832 (N_9832,N_9795,N_9753);
nor U9833 (N_9833,N_9633,N_9602);
or U9834 (N_9834,N_9655,N_9712);
nand U9835 (N_9835,N_9685,N_9618);
xnor U9836 (N_9836,N_9675,N_9627);
and U9837 (N_9837,N_9657,N_9630);
or U9838 (N_9838,N_9611,N_9642);
and U9839 (N_9839,N_9601,N_9687);
or U9840 (N_9840,N_9767,N_9640);
nand U9841 (N_9841,N_9797,N_9654);
nand U9842 (N_9842,N_9798,N_9628);
and U9843 (N_9843,N_9653,N_9713);
xnor U9844 (N_9844,N_9604,N_9645);
and U9845 (N_9845,N_9631,N_9770);
or U9846 (N_9846,N_9794,N_9784);
xor U9847 (N_9847,N_9786,N_9705);
nor U9848 (N_9848,N_9664,N_9715);
and U9849 (N_9849,N_9621,N_9744);
and U9850 (N_9850,N_9690,N_9725);
nand U9851 (N_9851,N_9639,N_9609);
nand U9852 (N_9852,N_9746,N_9615);
nor U9853 (N_9853,N_9727,N_9789);
nor U9854 (N_9854,N_9775,N_9718);
nand U9855 (N_9855,N_9669,N_9674);
xor U9856 (N_9856,N_9665,N_9638);
nor U9857 (N_9857,N_9787,N_9768);
nor U9858 (N_9858,N_9696,N_9656);
and U9859 (N_9859,N_9635,N_9688);
nand U9860 (N_9860,N_9741,N_9733);
or U9861 (N_9861,N_9790,N_9769);
xnor U9862 (N_9862,N_9608,N_9686);
xor U9863 (N_9863,N_9666,N_9613);
or U9864 (N_9864,N_9739,N_9709);
xor U9865 (N_9865,N_9663,N_9771);
nor U9866 (N_9866,N_9708,N_9774);
nor U9867 (N_9867,N_9703,N_9680);
xnor U9868 (N_9868,N_9699,N_9720);
xnor U9869 (N_9869,N_9799,N_9641);
or U9870 (N_9870,N_9728,N_9788);
or U9871 (N_9871,N_9648,N_9756);
nor U9872 (N_9872,N_9658,N_9752);
nor U9873 (N_9873,N_9734,N_9736);
nor U9874 (N_9874,N_9676,N_9783);
nand U9875 (N_9875,N_9671,N_9698);
xor U9876 (N_9876,N_9702,N_9679);
or U9877 (N_9877,N_9625,N_9754);
nand U9878 (N_9878,N_9761,N_9659);
or U9879 (N_9879,N_9706,N_9647);
nand U9880 (N_9880,N_9792,N_9778);
nand U9881 (N_9881,N_9650,N_9722);
and U9882 (N_9882,N_9622,N_9766);
nand U9883 (N_9883,N_9777,N_9626);
and U9884 (N_9884,N_9678,N_9697);
xor U9885 (N_9885,N_9652,N_9721);
xnor U9886 (N_9886,N_9723,N_9749);
nand U9887 (N_9887,N_9735,N_9750);
nor U9888 (N_9888,N_9781,N_9694);
or U9889 (N_9889,N_9634,N_9624);
xnor U9890 (N_9890,N_9636,N_9755);
and U9891 (N_9891,N_9782,N_9772);
nand U9892 (N_9892,N_9711,N_9726);
xor U9893 (N_9893,N_9780,N_9773);
nand U9894 (N_9894,N_9684,N_9779);
nand U9895 (N_9895,N_9704,N_9737);
and U9896 (N_9896,N_9607,N_9730);
nor U9897 (N_9897,N_9632,N_9793);
xnor U9898 (N_9898,N_9614,N_9612);
or U9899 (N_9899,N_9649,N_9729);
nor U9900 (N_9900,N_9615,N_9697);
nor U9901 (N_9901,N_9768,N_9702);
or U9902 (N_9902,N_9684,N_9737);
nor U9903 (N_9903,N_9752,N_9720);
and U9904 (N_9904,N_9622,N_9730);
or U9905 (N_9905,N_9654,N_9741);
nor U9906 (N_9906,N_9779,N_9653);
and U9907 (N_9907,N_9796,N_9699);
nand U9908 (N_9908,N_9745,N_9761);
nand U9909 (N_9909,N_9639,N_9633);
or U9910 (N_9910,N_9611,N_9627);
or U9911 (N_9911,N_9775,N_9740);
or U9912 (N_9912,N_9693,N_9612);
nand U9913 (N_9913,N_9766,N_9747);
nand U9914 (N_9914,N_9644,N_9719);
or U9915 (N_9915,N_9746,N_9649);
or U9916 (N_9916,N_9664,N_9790);
xnor U9917 (N_9917,N_9678,N_9629);
nor U9918 (N_9918,N_9700,N_9797);
or U9919 (N_9919,N_9606,N_9735);
and U9920 (N_9920,N_9722,N_9655);
nand U9921 (N_9921,N_9762,N_9697);
or U9922 (N_9922,N_9645,N_9785);
nor U9923 (N_9923,N_9647,N_9675);
and U9924 (N_9924,N_9765,N_9745);
xor U9925 (N_9925,N_9675,N_9781);
nand U9926 (N_9926,N_9790,N_9659);
nor U9927 (N_9927,N_9785,N_9600);
and U9928 (N_9928,N_9637,N_9757);
xor U9929 (N_9929,N_9662,N_9678);
xnor U9930 (N_9930,N_9732,N_9702);
nor U9931 (N_9931,N_9768,N_9610);
and U9932 (N_9932,N_9755,N_9702);
nor U9933 (N_9933,N_9615,N_9678);
and U9934 (N_9934,N_9728,N_9738);
and U9935 (N_9935,N_9684,N_9772);
or U9936 (N_9936,N_9682,N_9769);
nand U9937 (N_9937,N_9750,N_9675);
nand U9938 (N_9938,N_9610,N_9721);
nor U9939 (N_9939,N_9707,N_9638);
or U9940 (N_9940,N_9768,N_9609);
xor U9941 (N_9941,N_9794,N_9714);
or U9942 (N_9942,N_9677,N_9660);
and U9943 (N_9943,N_9657,N_9692);
xor U9944 (N_9944,N_9614,N_9738);
or U9945 (N_9945,N_9780,N_9698);
xnor U9946 (N_9946,N_9708,N_9697);
nor U9947 (N_9947,N_9642,N_9632);
and U9948 (N_9948,N_9790,N_9683);
nand U9949 (N_9949,N_9700,N_9704);
nand U9950 (N_9950,N_9730,N_9778);
or U9951 (N_9951,N_9651,N_9785);
nor U9952 (N_9952,N_9771,N_9639);
xor U9953 (N_9953,N_9632,N_9750);
nor U9954 (N_9954,N_9721,N_9732);
nand U9955 (N_9955,N_9765,N_9638);
nor U9956 (N_9956,N_9797,N_9640);
and U9957 (N_9957,N_9631,N_9686);
xor U9958 (N_9958,N_9785,N_9648);
and U9959 (N_9959,N_9732,N_9667);
nand U9960 (N_9960,N_9613,N_9629);
nor U9961 (N_9961,N_9652,N_9606);
xor U9962 (N_9962,N_9620,N_9714);
xnor U9963 (N_9963,N_9694,N_9633);
nor U9964 (N_9964,N_9652,N_9663);
nor U9965 (N_9965,N_9653,N_9673);
nor U9966 (N_9966,N_9612,N_9736);
nor U9967 (N_9967,N_9669,N_9755);
nand U9968 (N_9968,N_9725,N_9676);
or U9969 (N_9969,N_9775,N_9631);
or U9970 (N_9970,N_9611,N_9726);
xor U9971 (N_9971,N_9782,N_9675);
or U9972 (N_9972,N_9617,N_9674);
or U9973 (N_9973,N_9618,N_9765);
nor U9974 (N_9974,N_9629,N_9769);
xnor U9975 (N_9975,N_9788,N_9611);
nand U9976 (N_9976,N_9745,N_9654);
and U9977 (N_9977,N_9790,N_9699);
xnor U9978 (N_9978,N_9625,N_9775);
or U9979 (N_9979,N_9714,N_9768);
and U9980 (N_9980,N_9780,N_9791);
nand U9981 (N_9981,N_9765,N_9643);
xor U9982 (N_9982,N_9784,N_9718);
and U9983 (N_9983,N_9700,N_9742);
and U9984 (N_9984,N_9619,N_9687);
and U9985 (N_9985,N_9776,N_9643);
or U9986 (N_9986,N_9765,N_9740);
xnor U9987 (N_9987,N_9787,N_9685);
or U9988 (N_9988,N_9664,N_9798);
and U9989 (N_9989,N_9624,N_9723);
or U9990 (N_9990,N_9716,N_9730);
nor U9991 (N_9991,N_9684,N_9730);
nor U9992 (N_9992,N_9611,N_9683);
nor U9993 (N_9993,N_9781,N_9727);
or U9994 (N_9994,N_9646,N_9671);
and U9995 (N_9995,N_9768,N_9699);
nand U9996 (N_9996,N_9773,N_9642);
or U9997 (N_9997,N_9665,N_9676);
nor U9998 (N_9998,N_9629,N_9640);
nand U9999 (N_9999,N_9779,N_9734);
nor UO_0 (O_0,N_9940,N_9805);
nor UO_1 (O_1,N_9999,N_9995);
xnor UO_2 (O_2,N_9920,N_9934);
xor UO_3 (O_3,N_9837,N_9935);
and UO_4 (O_4,N_9840,N_9833);
or UO_5 (O_5,N_9976,N_9858);
or UO_6 (O_6,N_9907,N_9811);
and UO_7 (O_7,N_9830,N_9926);
nor UO_8 (O_8,N_9952,N_9975);
or UO_9 (O_9,N_9890,N_9897);
xor UO_10 (O_10,N_9984,N_9855);
and UO_11 (O_11,N_9803,N_9870);
nor UO_12 (O_12,N_9889,N_9950);
nand UO_13 (O_13,N_9836,N_9945);
nor UO_14 (O_14,N_9941,N_9816);
nor UO_15 (O_15,N_9997,N_9987);
xor UO_16 (O_16,N_9958,N_9972);
xnor UO_17 (O_17,N_9949,N_9887);
nor UO_18 (O_18,N_9882,N_9823);
and UO_19 (O_19,N_9939,N_9861);
nand UO_20 (O_20,N_9872,N_9894);
and UO_21 (O_21,N_9996,N_9961);
nor UO_22 (O_22,N_9905,N_9914);
nor UO_23 (O_23,N_9839,N_9919);
or UO_24 (O_24,N_9970,N_9865);
nand UO_25 (O_25,N_9822,N_9866);
xnor UO_26 (O_26,N_9802,N_9883);
nand UO_27 (O_27,N_9832,N_9899);
nand UO_28 (O_28,N_9967,N_9843);
nand UO_29 (O_29,N_9925,N_9814);
and UO_30 (O_30,N_9885,N_9928);
nor UO_31 (O_31,N_9978,N_9847);
or UO_32 (O_32,N_9924,N_9902);
or UO_33 (O_33,N_9810,N_9977);
xnor UO_34 (O_34,N_9871,N_9842);
and UO_35 (O_35,N_9827,N_9844);
xnor UO_36 (O_36,N_9900,N_9821);
xnor UO_37 (O_37,N_9981,N_9955);
and UO_38 (O_38,N_9850,N_9909);
nand UO_39 (O_39,N_9876,N_9906);
nor UO_40 (O_40,N_9912,N_9910);
nor UO_41 (O_41,N_9852,N_9911);
and UO_42 (O_42,N_9988,N_9942);
nand UO_43 (O_43,N_9971,N_9983);
xnor UO_44 (O_44,N_9886,N_9953);
xnor UO_45 (O_45,N_9916,N_9834);
and UO_46 (O_46,N_9820,N_9923);
xnor UO_47 (O_47,N_9835,N_9956);
nand UO_48 (O_48,N_9884,N_9938);
nor UO_49 (O_49,N_9895,N_9980);
nor UO_50 (O_50,N_9807,N_9809);
and UO_51 (O_51,N_9918,N_9812);
and UO_52 (O_52,N_9829,N_9892);
nand UO_53 (O_53,N_9936,N_9873);
nand UO_54 (O_54,N_9990,N_9888);
and UO_55 (O_55,N_9854,N_9903);
or UO_56 (O_56,N_9891,N_9915);
or UO_57 (O_57,N_9825,N_9921);
xor UO_58 (O_58,N_9960,N_9878);
or UO_59 (O_59,N_9845,N_9946);
and UO_60 (O_60,N_9853,N_9904);
and UO_61 (O_61,N_9931,N_9813);
or UO_62 (O_62,N_9879,N_9804);
nand UO_63 (O_63,N_9989,N_9932);
nand UO_64 (O_64,N_9992,N_9859);
xnor UO_65 (O_65,N_9957,N_9969);
xnor UO_66 (O_66,N_9922,N_9857);
and UO_67 (O_67,N_9913,N_9838);
and UO_68 (O_68,N_9896,N_9930);
nand UO_69 (O_69,N_9868,N_9944);
or UO_70 (O_70,N_9929,N_9991);
or UO_71 (O_71,N_9968,N_9801);
or UO_72 (O_72,N_9826,N_9874);
nor UO_73 (O_73,N_9828,N_9943);
and UO_74 (O_74,N_9849,N_9948);
nand UO_75 (O_75,N_9806,N_9862);
nand UO_76 (O_76,N_9841,N_9817);
nand UO_77 (O_77,N_9993,N_9860);
and UO_78 (O_78,N_9962,N_9927);
and UO_79 (O_79,N_9815,N_9964);
xnor UO_80 (O_80,N_9898,N_9937);
and UO_81 (O_81,N_9863,N_9951);
xnor UO_82 (O_82,N_9875,N_9994);
or UO_83 (O_83,N_9985,N_9848);
nand UO_84 (O_84,N_9881,N_9893);
or UO_85 (O_85,N_9986,N_9908);
nand UO_86 (O_86,N_9954,N_9851);
nand UO_87 (O_87,N_9864,N_9959);
nand UO_88 (O_88,N_9947,N_9856);
or UO_89 (O_89,N_9819,N_9880);
and UO_90 (O_90,N_9998,N_9818);
and UO_91 (O_91,N_9869,N_9831);
and UO_92 (O_92,N_9966,N_9867);
nor UO_93 (O_93,N_9877,N_9917);
and UO_94 (O_94,N_9973,N_9963);
or UO_95 (O_95,N_9901,N_9933);
and UO_96 (O_96,N_9808,N_9982);
nand UO_97 (O_97,N_9846,N_9800);
nor UO_98 (O_98,N_9974,N_9979);
nand UO_99 (O_99,N_9965,N_9824);
nor UO_100 (O_100,N_9882,N_9825);
nor UO_101 (O_101,N_9889,N_9891);
nor UO_102 (O_102,N_9810,N_9829);
xor UO_103 (O_103,N_9977,N_9818);
nand UO_104 (O_104,N_9842,N_9883);
xnor UO_105 (O_105,N_9967,N_9958);
nor UO_106 (O_106,N_9892,N_9862);
nor UO_107 (O_107,N_9847,N_9892);
nor UO_108 (O_108,N_9954,N_9910);
or UO_109 (O_109,N_9999,N_9824);
xor UO_110 (O_110,N_9860,N_9819);
nand UO_111 (O_111,N_9834,N_9889);
nand UO_112 (O_112,N_9887,N_9869);
nand UO_113 (O_113,N_9803,N_9844);
nand UO_114 (O_114,N_9882,N_9868);
nand UO_115 (O_115,N_9886,N_9908);
or UO_116 (O_116,N_9989,N_9892);
xor UO_117 (O_117,N_9883,N_9979);
xor UO_118 (O_118,N_9821,N_9944);
xor UO_119 (O_119,N_9873,N_9882);
or UO_120 (O_120,N_9923,N_9917);
xnor UO_121 (O_121,N_9833,N_9849);
or UO_122 (O_122,N_9983,N_9801);
xor UO_123 (O_123,N_9999,N_9955);
nand UO_124 (O_124,N_9926,N_9848);
nor UO_125 (O_125,N_9933,N_9966);
or UO_126 (O_126,N_9829,N_9927);
and UO_127 (O_127,N_9974,N_9864);
nor UO_128 (O_128,N_9991,N_9899);
xor UO_129 (O_129,N_9888,N_9847);
or UO_130 (O_130,N_9957,N_9984);
xnor UO_131 (O_131,N_9906,N_9844);
or UO_132 (O_132,N_9818,N_9813);
and UO_133 (O_133,N_9801,N_9902);
xnor UO_134 (O_134,N_9822,N_9842);
nor UO_135 (O_135,N_9849,N_9963);
xnor UO_136 (O_136,N_9959,N_9822);
xor UO_137 (O_137,N_9844,N_9915);
nor UO_138 (O_138,N_9894,N_9957);
xnor UO_139 (O_139,N_9906,N_9804);
xor UO_140 (O_140,N_9999,N_9975);
or UO_141 (O_141,N_9837,N_9985);
and UO_142 (O_142,N_9934,N_9820);
nor UO_143 (O_143,N_9834,N_9870);
and UO_144 (O_144,N_9840,N_9963);
xnor UO_145 (O_145,N_9908,N_9838);
or UO_146 (O_146,N_9823,N_9895);
nor UO_147 (O_147,N_9992,N_9963);
and UO_148 (O_148,N_9998,N_9878);
nor UO_149 (O_149,N_9982,N_9839);
nand UO_150 (O_150,N_9833,N_9875);
and UO_151 (O_151,N_9815,N_9970);
or UO_152 (O_152,N_9883,N_9975);
xor UO_153 (O_153,N_9904,N_9859);
nor UO_154 (O_154,N_9963,N_9877);
or UO_155 (O_155,N_9902,N_9828);
nor UO_156 (O_156,N_9874,N_9891);
or UO_157 (O_157,N_9853,N_9881);
nand UO_158 (O_158,N_9803,N_9986);
xor UO_159 (O_159,N_9866,N_9970);
and UO_160 (O_160,N_9843,N_9875);
xnor UO_161 (O_161,N_9902,N_9872);
xor UO_162 (O_162,N_9980,N_9965);
or UO_163 (O_163,N_9828,N_9909);
or UO_164 (O_164,N_9997,N_9954);
and UO_165 (O_165,N_9972,N_9909);
nand UO_166 (O_166,N_9894,N_9812);
and UO_167 (O_167,N_9923,N_9880);
nand UO_168 (O_168,N_9864,N_9842);
nor UO_169 (O_169,N_9894,N_9913);
nand UO_170 (O_170,N_9910,N_9941);
nand UO_171 (O_171,N_9975,N_9953);
xnor UO_172 (O_172,N_9881,N_9999);
nor UO_173 (O_173,N_9945,N_9946);
or UO_174 (O_174,N_9865,N_9890);
or UO_175 (O_175,N_9982,N_9948);
xnor UO_176 (O_176,N_9812,N_9992);
nor UO_177 (O_177,N_9849,N_9914);
or UO_178 (O_178,N_9840,N_9814);
and UO_179 (O_179,N_9995,N_9809);
xnor UO_180 (O_180,N_9820,N_9814);
xnor UO_181 (O_181,N_9917,N_9808);
nor UO_182 (O_182,N_9859,N_9879);
nand UO_183 (O_183,N_9873,N_9983);
or UO_184 (O_184,N_9932,N_9852);
nand UO_185 (O_185,N_9889,N_9916);
and UO_186 (O_186,N_9811,N_9865);
nand UO_187 (O_187,N_9913,N_9890);
nor UO_188 (O_188,N_9806,N_9859);
nand UO_189 (O_189,N_9872,N_9877);
or UO_190 (O_190,N_9819,N_9879);
or UO_191 (O_191,N_9863,N_9927);
nor UO_192 (O_192,N_9912,N_9849);
nor UO_193 (O_193,N_9887,N_9993);
xnor UO_194 (O_194,N_9812,N_9978);
xnor UO_195 (O_195,N_9903,N_9869);
and UO_196 (O_196,N_9998,N_9838);
xor UO_197 (O_197,N_9979,N_9961);
and UO_198 (O_198,N_9825,N_9806);
nor UO_199 (O_199,N_9826,N_9818);
or UO_200 (O_200,N_9990,N_9898);
or UO_201 (O_201,N_9843,N_9857);
or UO_202 (O_202,N_9852,N_9962);
xnor UO_203 (O_203,N_9858,N_9951);
xnor UO_204 (O_204,N_9842,N_9974);
xor UO_205 (O_205,N_9874,N_9932);
or UO_206 (O_206,N_9849,N_9871);
or UO_207 (O_207,N_9803,N_9928);
nand UO_208 (O_208,N_9846,N_9866);
or UO_209 (O_209,N_9835,N_9981);
xor UO_210 (O_210,N_9848,N_9927);
xnor UO_211 (O_211,N_9999,N_9914);
nand UO_212 (O_212,N_9931,N_9869);
xor UO_213 (O_213,N_9997,N_9837);
xnor UO_214 (O_214,N_9923,N_9833);
or UO_215 (O_215,N_9935,N_9803);
xor UO_216 (O_216,N_9962,N_9837);
nor UO_217 (O_217,N_9956,N_9906);
and UO_218 (O_218,N_9939,N_9974);
nand UO_219 (O_219,N_9939,N_9847);
nand UO_220 (O_220,N_9854,N_9998);
and UO_221 (O_221,N_9937,N_9911);
nand UO_222 (O_222,N_9938,N_9987);
nor UO_223 (O_223,N_9976,N_9825);
nor UO_224 (O_224,N_9810,N_9804);
and UO_225 (O_225,N_9832,N_9913);
nand UO_226 (O_226,N_9996,N_9845);
or UO_227 (O_227,N_9817,N_9936);
xor UO_228 (O_228,N_9983,N_9949);
xor UO_229 (O_229,N_9930,N_9924);
nor UO_230 (O_230,N_9820,N_9829);
nor UO_231 (O_231,N_9871,N_9964);
nor UO_232 (O_232,N_9817,N_9880);
or UO_233 (O_233,N_9846,N_9986);
and UO_234 (O_234,N_9854,N_9946);
and UO_235 (O_235,N_9973,N_9884);
and UO_236 (O_236,N_9927,N_9832);
and UO_237 (O_237,N_9901,N_9987);
xor UO_238 (O_238,N_9802,N_9890);
or UO_239 (O_239,N_9989,N_9827);
nand UO_240 (O_240,N_9997,N_9862);
or UO_241 (O_241,N_9932,N_9935);
nand UO_242 (O_242,N_9808,N_9945);
or UO_243 (O_243,N_9838,N_9801);
or UO_244 (O_244,N_9973,N_9805);
nand UO_245 (O_245,N_9930,N_9969);
xnor UO_246 (O_246,N_9957,N_9926);
xnor UO_247 (O_247,N_9934,N_9878);
or UO_248 (O_248,N_9956,N_9879);
and UO_249 (O_249,N_9873,N_9853);
or UO_250 (O_250,N_9961,N_9804);
xnor UO_251 (O_251,N_9840,N_9990);
or UO_252 (O_252,N_9804,N_9898);
nor UO_253 (O_253,N_9963,N_9936);
or UO_254 (O_254,N_9865,N_9896);
or UO_255 (O_255,N_9911,N_9957);
xnor UO_256 (O_256,N_9964,N_9811);
or UO_257 (O_257,N_9817,N_9992);
or UO_258 (O_258,N_9802,N_9824);
nand UO_259 (O_259,N_9878,N_9830);
and UO_260 (O_260,N_9835,N_9858);
and UO_261 (O_261,N_9953,N_9898);
nor UO_262 (O_262,N_9843,N_9988);
nand UO_263 (O_263,N_9986,N_9848);
nor UO_264 (O_264,N_9973,N_9888);
and UO_265 (O_265,N_9904,N_9918);
nor UO_266 (O_266,N_9957,N_9815);
and UO_267 (O_267,N_9870,N_9990);
or UO_268 (O_268,N_9891,N_9917);
or UO_269 (O_269,N_9969,N_9864);
or UO_270 (O_270,N_9963,N_9919);
nor UO_271 (O_271,N_9808,N_9847);
and UO_272 (O_272,N_9862,N_9876);
and UO_273 (O_273,N_9853,N_9924);
nor UO_274 (O_274,N_9953,N_9885);
or UO_275 (O_275,N_9937,N_9981);
nand UO_276 (O_276,N_9823,N_9896);
xor UO_277 (O_277,N_9906,N_9967);
xnor UO_278 (O_278,N_9864,N_9898);
and UO_279 (O_279,N_9916,N_9864);
or UO_280 (O_280,N_9824,N_9807);
nand UO_281 (O_281,N_9936,N_9824);
or UO_282 (O_282,N_9823,N_9825);
nand UO_283 (O_283,N_9848,N_9950);
xor UO_284 (O_284,N_9843,N_9990);
xnor UO_285 (O_285,N_9812,N_9823);
nor UO_286 (O_286,N_9822,N_9809);
and UO_287 (O_287,N_9868,N_9815);
or UO_288 (O_288,N_9811,N_9807);
nor UO_289 (O_289,N_9960,N_9906);
or UO_290 (O_290,N_9827,N_9953);
nor UO_291 (O_291,N_9892,N_9932);
nor UO_292 (O_292,N_9880,N_9859);
or UO_293 (O_293,N_9914,N_9935);
nor UO_294 (O_294,N_9922,N_9987);
nor UO_295 (O_295,N_9816,N_9905);
and UO_296 (O_296,N_9856,N_9822);
xnor UO_297 (O_297,N_9858,N_9916);
xor UO_298 (O_298,N_9858,N_9853);
nor UO_299 (O_299,N_9993,N_9911);
or UO_300 (O_300,N_9860,N_9838);
nand UO_301 (O_301,N_9821,N_9986);
and UO_302 (O_302,N_9849,N_9907);
nand UO_303 (O_303,N_9991,N_9835);
or UO_304 (O_304,N_9966,N_9833);
nand UO_305 (O_305,N_9944,N_9974);
nand UO_306 (O_306,N_9906,N_9959);
nand UO_307 (O_307,N_9824,N_9990);
and UO_308 (O_308,N_9936,N_9803);
nand UO_309 (O_309,N_9862,N_9801);
nand UO_310 (O_310,N_9855,N_9836);
or UO_311 (O_311,N_9971,N_9928);
or UO_312 (O_312,N_9885,N_9834);
nor UO_313 (O_313,N_9883,N_9804);
and UO_314 (O_314,N_9862,N_9846);
and UO_315 (O_315,N_9935,N_9807);
and UO_316 (O_316,N_9834,N_9981);
xnor UO_317 (O_317,N_9923,N_9852);
or UO_318 (O_318,N_9887,N_9809);
and UO_319 (O_319,N_9827,N_9969);
nand UO_320 (O_320,N_9842,N_9934);
nor UO_321 (O_321,N_9854,N_9933);
or UO_322 (O_322,N_9947,N_9839);
nand UO_323 (O_323,N_9935,N_9921);
nand UO_324 (O_324,N_9962,N_9838);
nor UO_325 (O_325,N_9841,N_9866);
or UO_326 (O_326,N_9894,N_9928);
nor UO_327 (O_327,N_9862,N_9830);
and UO_328 (O_328,N_9825,N_9848);
or UO_329 (O_329,N_9979,N_9834);
and UO_330 (O_330,N_9900,N_9980);
and UO_331 (O_331,N_9837,N_9803);
xnor UO_332 (O_332,N_9906,N_9932);
nand UO_333 (O_333,N_9802,N_9934);
xor UO_334 (O_334,N_9952,N_9833);
or UO_335 (O_335,N_9886,N_9844);
nand UO_336 (O_336,N_9906,N_9922);
or UO_337 (O_337,N_9837,N_9845);
and UO_338 (O_338,N_9919,N_9905);
nor UO_339 (O_339,N_9952,N_9941);
or UO_340 (O_340,N_9889,N_9930);
and UO_341 (O_341,N_9861,N_9865);
or UO_342 (O_342,N_9958,N_9869);
and UO_343 (O_343,N_9961,N_9903);
xor UO_344 (O_344,N_9883,N_9996);
nor UO_345 (O_345,N_9849,N_9961);
and UO_346 (O_346,N_9803,N_9974);
xnor UO_347 (O_347,N_9865,N_9853);
nand UO_348 (O_348,N_9871,N_9983);
nor UO_349 (O_349,N_9911,N_9874);
or UO_350 (O_350,N_9906,N_9832);
and UO_351 (O_351,N_9956,N_9864);
and UO_352 (O_352,N_9892,N_9887);
xnor UO_353 (O_353,N_9986,N_9931);
nand UO_354 (O_354,N_9979,N_9982);
and UO_355 (O_355,N_9969,N_9805);
and UO_356 (O_356,N_9918,N_9858);
or UO_357 (O_357,N_9828,N_9838);
and UO_358 (O_358,N_9810,N_9923);
nor UO_359 (O_359,N_9976,N_9855);
or UO_360 (O_360,N_9979,N_9995);
or UO_361 (O_361,N_9804,N_9871);
nand UO_362 (O_362,N_9840,N_9953);
nand UO_363 (O_363,N_9969,N_9962);
and UO_364 (O_364,N_9845,N_9872);
and UO_365 (O_365,N_9859,N_9945);
nand UO_366 (O_366,N_9846,N_9854);
nand UO_367 (O_367,N_9856,N_9929);
nor UO_368 (O_368,N_9946,N_9860);
or UO_369 (O_369,N_9945,N_9876);
and UO_370 (O_370,N_9909,N_9819);
or UO_371 (O_371,N_9883,N_9902);
or UO_372 (O_372,N_9959,N_9946);
or UO_373 (O_373,N_9872,N_9926);
and UO_374 (O_374,N_9983,N_9977);
nand UO_375 (O_375,N_9891,N_9852);
or UO_376 (O_376,N_9976,N_9953);
or UO_377 (O_377,N_9974,N_9872);
nor UO_378 (O_378,N_9853,N_9972);
or UO_379 (O_379,N_9941,N_9875);
nor UO_380 (O_380,N_9987,N_9960);
or UO_381 (O_381,N_9928,N_9934);
and UO_382 (O_382,N_9819,N_9854);
and UO_383 (O_383,N_9904,N_9978);
nand UO_384 (O_384,N_9824,N_9878);
or UO_385 (O_385,N_9878,N_9827);
nand UO_386 (O_386,N_9860,N_9981);
and UO_387 (O_387,N_9868,N_9860);
xnor UO_388 (O_388,N_9950,N_9959);
xnor UO_389 (O_389,N_9883,N_9877);
nor UO_390 (O_390,N_9867,N_9855);
xor UO_391 (O_391,N_9893,N_9820);
and UO_392 (O_392,N_9871,N_9854);
or UO_393 (O_393,N_9902,N_9900);
and UO_394 (O_394,N_9847,N_9976);
and UO_395 (O_395,N_9952,N_9926);
xor UO_396 (O_396,N_9850,N_9837);
xnor UO_397 (O_397,N_9944,N_9890);
and UO_398 (O_398,N_9836,N_9944);
nor UO_399 (O_399,N_9822,N_9890);
nor UO_400 (O_400,N_9871,N_9944);
and UO_401 (O_401,N_9995,N_9825);
xor UO_402 (O_402,N_9973,N_9959);
nand UO_403 (O_403,N_9840,N_9914);
or UO_404 (O_404,N_9948,N_9824);
or UO_405 (O_405,N_9822,N_9906);
nand UO_406 (O_406,N_9928,N_9895);
or UO_407 (O_407,N_9886,N_9881);
or UO_408 (O_408,N_9814,N_9897);
nand UO_409 (O_409,N_9819,N_9938);
xnor UO_410 (O_410,N_9921,N_9999);
xnor UO_411 (O_411,N_9917,N_9931);
nand UO_412 (O_412,N_9804,N_9849);
and UO_413 (O_413,N_9993,N_9877);
nor UO_414 (O_414,N_9923,N_9905);
xor UO_415 (O_415,N_9815,N_9840);
and UO_416 (O_416,N_9840,N_9987);
xnor UO_417 (O_417,N_9952,N_9959);
xnor UO_418 (O_418,N_9895,N_9910);
xnor UO_419 (O_419,N_9865,N_9893);
nor UO_420 (O_420,N_9866,N_9967);
nand UO_421 (O_421,N_9928,N_9876);
xnor UO_422 (O_422,N_9994,N_9906);
and UO_423 (O_423,N_9819,N_9883);
xor UO_424 (O_424,N_9868,N_9921);
nor UO_425 (O_425,N_9907,N_9988);
xor UO_426 (O_426,N_9853,N_9991);
xor UO_427 (O_427,N_9804,N_9850);
nand UO_428 (O_428,N_9970,N_9857);
nand UO_429 (O_429,N_9990,N_9957);
xnor UO_430 (O_430,N_9876,N_9925);
nand UO_431 (O_431,N_9924,N_9859);
and UO_432 (O_432,N_9990,N_9907);
nor UO_433 (O_433,N_9942,N_9958);
and UO_434 (O_434,N_9854,N_9805);
nand UO_435 (O_435,N_9843,N_9835);
nand UO_436 (O_436,N_9934,N_9891);
xor UO_437 (O_437,N_9805,N_9868);
and UO_438 (O_438,N_9911,N_9848);
or UO_439 (O_439,N_9876,N_9844);
or UO_440 (O_440,N_9970,N_9861);
or UO_441 (O_441,N_9879,N_9897);
nor UO_442 (O_442,N_9827,N_9850);
or UO_443 (O_443,N_9827,N_9924);
and UO_444 (O_444,N_9829,N_9841);
nor UO_445 (O_445,N_9869,N_9857);
nor UO_446 (O_446,N_9800,N_9904);
nand UO_447 (O_447,N_9967,N_9805);
xor UO_448 (O_448,N_9960,N_9823);
xor UO_449 (O_449,N_9885,N_9871);
or UO_450 (O_450,N_9926,N_9979);
nor UO_451 (O_451,N_9980,N_9921);
xnor UO_452 (O_452,N_9890,N_9851);
and UO_453 (O_453,N_9961,N_9875);
and UO_454 (O_454,N_9937,N_9840);
and UO_455 (O_455,N_9951,N_9882);
xnor UO_456 (O_456,N_9908,N_9964);
nand UO_457 (O_457,N_9820,N_9921);
xor UO_458 (O_458,N_9894,N_9847);
and UO_459 (O_459,N_9831,N_9834);
and UO_460 (O_460,N_9882,N_9803);
xnor UO_461 (O_461,N_9889,N_9880);
nand UO_462 (O_462,N_9861,N_9873);
xnor UO_463 (O_463,N_9996,N_9807);
or UO_464 (O_464,N_9859,N_9824);
nor UO_465 (O_465,N_9977,N_9872);
nand UO_466 (O_466,N_9960,N_9851);
and UO_467 (O_467,N_9997,N_9847);
xnor UO_468 (O_468,N_9932,N_9825);
nand UO_469 (O_469,N_9849,N_9881);
and UO_470 (O_470,N_9998,N_9831);
nor UO_471 (O_471,N_9946,N_9902);
xnor UO_472 (O_472,N_9858,N_9995);
or UO_473 (O_473,N_9806,N_9967);
nor UO_474 (O_474,N_9932,N_9836);
and UO_475 (O_475,N_9961,N_9928);
and UO_476 (O_476,N_9998,N_9853);
or UO_477 (O_477,N_9875,N_9891);
and UO_478 (O_478,N_9942,N_9870);
and UO_479 (O_479,N_9882,N_9906);
and UO_480 (O_480,N_9908,N_9910);
nor UO_481 (O_481,N_9929,N_9973);
or UO_482 (O_482,N_9818,N_9872);
nand UO_483 (O_483,N_9911,N_9814);
xnor UO_484 (O_484,N_9955,N_9950);
nand UO_485 (O_485,N_9918,N_9881);
xor UO_486 (O_486,N_9820,N_9830);
and UO_487 (O_487,N_9817,N_9866);
nor UO_488 (O_488,N_9980,N_9954);
nand UO_489 (O_489,N_9819,N_9885);
or UO_490 (O_490,N_9903,N_9824);
and UO_491 (O_491,N_9842,N_9893);
or UO_492 (O_492,N_9945,N_9848);
nor UO_493 (O_493,N_9920,N_9831);
and UO_494 (O_494,N_9905,N_9836);
nor UO_495 (O_495,N_9851,N_9850);
or UO_496 (O_496,N_9950,N_9985);
nor UO_497 (O_497,N_9866,N_9906);
nor UO_498 (O_498,N_9876,N_9835);
and UO_499 (O_499,N_9839,N_9828);
nor UO_500 (O_500,N_9933,N_9932);
nand UO_501 (O_501,N_9960,N_9991);
or UO_502 (O_502,N_9815,N_9894);
nor UO_503 (O_503,N_9958,N_9856);
nor UO_504 (O_504,N_9996,N_9970);
nand UO_505 (O_505,N_9907,N_9941);
nand UO_506 (O_506,N_9953,N_9818);
nor UO_507 (O_507,N_9807,N_9865);
nor UO_508 (O_508,N_9942,N_9984);
xor UO_509 (O_509,N_9887,N_9866);
nand UO_510 (O_510,N_9843,N_9934);
and UO_511 (O_511,N_9891,N_9976);
and UO_512 (O_512,N_9911,N_9970);
nand UO_513 (O_513,N_9838,N_9857);
and UO_514 (O_514,N_9896,N_9949);
xor UO_515 (O_515,N_9925,N_9828);
or UO_516 (O_516,N_9968,N_9943);
or UO_517 (O_517,N_9897,N_9982);
nand UO_518 (O_518,N_9903,N_9990);
nand UO_519 (O_519,N_9951,N_9967);
or UO_520 (O_520,N_9995,N_9813);
and UO_521 (O_521,N_9846,N_9974);
nor UO_522 (O_522,N_9953,N_9906);
and UO_523 (O_523,N_9943,N_9878);
xor UO_524 (O_524,N_9897,N_9828);
xor UO_525 (O_525,N_9873,N_9978);
and UO_526 (O_526,N_9892,N_9992);
or UO_527 (O_527,N_9893,N_9831);
or UO_528 (O_528,N_9878,N_9917);
or UO_529 (O_529,N_9884,N_9854);
xor UO_530 (O_530,N_9998,N_9939);
or UO_531 (O_531,N_9965,N_9921);
and UO_532 (O_532,N_9996,N_9984);
nor UO_533 (O_533,N_9915,N_9960);
nor UO_534 (O_534,N_9924,N_9879);
nor UO_535 (O_535,N_9839,N_9962);
and UO_536 (O_536,N_9804,N_9921);
nand UO_537 (O_537,N_9926,N_9942);
or UO_538 (O_538,N_9812,N_9953);
or UO_539 (O_539,N_9826,N_9938);
and UO_540 (O_540,N_9948,N_9838);
nor UO_541 (O_541,N_9992,N_9996);
and UO_542 (O_542,N_9997,N_9833);
and UO_543 (O_543,N_9882,N_9946);
nor UO_544 (O_544,N_9813,N_9823);
and UO_545 (O_545,N_9948,N_9818);
nand UO_546 (O_546,N_9945,N_9816);
xnor UO_547 (O_547,N_9814,N_9940);
or UO_548 (O_548,N_9854,N_9994);
and UO_549 (O_549,N_9850,N_9920);
xnor UO_550 (O_550,N_9804,N_9874);
and UO_551 (O_551,N_9917,N_9832);
nand UO_552 (O_552,N_9851,N_9974);
nor UO_553 (O_553,N_9948,N_9813);
xor UO_554 (O_554,N_9865,N_9903);
nand UO_555 (O_555,N_9958,N_9895);
or UO_556 (O_556,N_9954,N_9926);
nor UO_557 (O_557,N_9952,N_9905);
nand UO_558 (O_558,N_9864,N_9878);
nor UO_559 (O_559,N_9930,N_9954);
nor UO_560 (O_560,N_9946,N_9813);
nor UO_561 (O_561,N_9993,N_9822);
and UO_562 (O_562,N_9951,N_9920);
or UO_563 (O_563,N_9975,N_9962);
and UO_564 (O_564,N_9830,N_9902);
or UO_565 (O_565,N_9938,N_9873);
nor UO_566 (O_566,N_9842,N_9910);
or UO_567 (O_567,N_9865,N_9900);
xnor UO_568 (O_568,N_9974,N_9919);
xnor UO_569 (O_569,N_9872,N_9820);
xnor UO_570 (O_570,N_9813,N_9844);
nand UO_571 (O_571,N_9862,N_9805);
and UO_572 (O_572,N_9809,N_9870);
or UO_573 (O_573,N_9967,N_9908);
nand UO_574 (O_574,N_9934,N_9962);
nand UO_575 (O_575,N_9941,N_9815);
xnor UO_576 (O_576,N_9829,N_9885);
and UO_577 (O_577,N_9995,N_9856);
nor UO_578 (O_578,N_9958,N_9943);
or UO_579 (O_579,N_9981,N_9917);
xnor UO_580 (O_580,N_9821,N_9888);
xor UO_581 (O_581,N_9805,N_9803);
nand UO_582 (O_582,N_9802,N_9973);
nand UO_583 (O_583,N_9950,N_9856);
and UO_584 (O_584,N_9877,N_9965);
nand UO_585 (O_585,N_9979,N_9893);
or UO_586 (O_586,N_9989,N_9990);
nor UO_587 (O_587,N_9948,N_9805);
and UO_588 (O_588,N_9842,N_9905);
or UO_589 (O_589,N_9994,N_9874);
and UO_590 (O_590,N_9893,N_9889);
and UO_591 (O_591,N_9818,N_9947);
nand UO_592 (O_592,N_9970,N_9811);
or UO_593 (O_593,N_9813,N_9912);
or UO_594 (O_594,N_9868,N_9963);
or UO_595 (O_595,N_9966,N_9918);
and UO_596 (O_596,N_9985,N_9922);
or UO_597 (O_597,N_9839,N_9897);
nor UO_598 (O_598,N_9991,N_9921);
nor UO_599 (O_599,N_9901,N_9857);
or UO_600 (O_600,N_9994,N_9859);
or UO_601 (O_601,N_9886,N_9948);
or UO_602 (O_602,N_9912,N_9956);
xnor UO_603 (O_603,N_9869,N_9962);
xnor UO_604 (O_604,N_9961,N_9847);
nand UO_605 (O_605,N_9804,N_9950);
nand UO_606 (O_606,N_9859,N_9889);
nand UO_607 (O_607,N_9876,N_9880);
xor UO_608 (O_608,N_9805,N_9987);
xnor UO_609 (O_609,N_9860,N_9927);
and UO_610 (O_610,N_9911,N_9827);
nor UO_611 (O_611,N_9928,N_9897);
xor UO_612 (O_612,N_9858,N_9857);
xnor UO_613 (O_613,N_9899,N_9913);
or UO_614 (O_614,N_9819,N_9817);
xnor UO_615 (O_615,N_9822,N_9836);
nor UO_616 (O_616,N_9940,N_9929);
and UO_617 (O_617,N_9867,N_9805);
and UO_618 (O_618,N_9895,N_9808);
nor UO_619 (O_619,N_9971,N_9838);
and UO_620 (O_620,N_9872,N_9893);
or UO_621 (O_621,N_9872,N_9858);
or UO_622 (O_622,N_9931,N_9969);
xnor UO_623 (O_623,N_9844,N_9849);
nor UO_624 (O_624,N_9835,N_9969);
or UO_625 (O_625,N_9826,N_9955);
xnor UO_626 (O_626,N_9816,N_9843);
or UO_627 (O_627,N_9992,N_9995);
and UO_628 (O_628,N_9900,N_9926);
nand UO_629 (O_629,N_9904,N_9986);
and UO_630 (O_630,N_9838,N_9869);
or UO_631 (O_631,N_9952,N_9940);
or UO_632 (O_632,N_9890,N_9967);
nor UO_633 (O_633,N_9987,N_9858);
xnor UO_634 (O_634,N_9938,N_9876);
xor UO_635 (O_635,N_9877,N_9884);
xnor UO_636 (O_636,N_9800,N_9919);
or UO_637 (O_637,N_9809,N_9974);
and UO_638 (O_638,N_9958,N_9890);
nor UO_639 (O_639,N_9998,N_9999);
and UO_640 (O_640,N_9809,N_9872);
nor UO_641 (O_641,N_9840,N_9887);
xnor UO_642 (O_642,N_9902,N_9974);
or UO_643 (O_643,N_9911,N_9879);
and UO_644 (O_644,N_9818,N_9808);
and UO_645 (O_645,N_9937,N_9814);
nor UO_646 (O_646,N_9935,N_9836);
and UO_647 (O_647,N_9956,N_9880);
and UO_648 (O_648,N_9888,N_9893);
nor UO_649 (O_649,N_9813,N_9871);
nand UO_650 (O_650,N_9927,N_9819);
nand UO_651 (O_651,N_9802,N_9940);
nand UO_652 (O_652,N_9875,N_9885);
or UO_653 (O_653,N_9816,N_9856);
nand UO_654 (O_654,N_9810,N_9987);
nand UO_655 (O_655,N_9996,N_9978);
or UO_656 (O_656,N_9967,N_9802);
xor UO_657 (O_657,N_9914,N_9845);
nand UO_658 (O_658,N_9976,N_9875);
xnor UO_659 (O_659,N_9963,N_9886);
xnor UO_660 (O_660,N_9852,N_9902);
xnor UO_661 (O_661,N_9886,N_9841);
and UO_662 (O_662,N_9939,N_9943);
xor UO_663 (O_663,N_9920,N_9898);
and UO_664 (O_664,N_9980,N_9844);
nor UO_665 (O_665,N_9816,N_9933);
nand UO_666 (O_666,N_9849,N_9814);
xnor UO_667 (O_667,N_9940,N_9821);
nor UO_668 (O_668,N_9847,N_9994);
nand UO_669 (O_669,N_9829,N_9943);
and UO_670 (O_670,N_9953,N_9990);
or UO_671 (O_671,N_9973,N_9872);
and UO_672 (O_672,N_9802,N_9994);
xnor UO_673 (O_673,N_9928,N_9888);
and UO_674 (O_674,N_9851,N_9800);
and UO_675 (O_675,N_9831,N_9960);
nand UO_676 (O_676,N_9936,N_9913);
or UO_677 (O_677,N_9845,N_9990);
nand UO_678 (O_678,N_9946,N_9934);
nand UO_679 (O_679,N_9837,N_9973);
nand UO_680 (O_680,N_9945,N_9994);
and UO_681 (O_681,N_9805,N_9935);
nand UO_682 (O_682,N_9810,N_9903);
and UO_683 (O_683,N_9803,N_9815);
and UO_684 (O_684,N_9995,N_9915);
and UO_685 (O_685,N_9894,N_9992);
or UO_686 (O_686,N_9807,N_9808);
nand UO_687 (O_687,N_9858,N_9948);
xor UO_688 (O_688,N_9855,N_9964);
and UO_689 (O_689,N_9809,N_9908);
nand UO_690 (O_690,N_9950,N_9826);
nor UO_691 (O_691,N_9963,N_9946);
or UO_692 (O_692,N_9889,N_9894);
and UO_693 (O_693,N_9902,N_9885);
nand UO_694 (O_694,N_9963,N_9967);
nor UO_695 (O_695,N_9949,N_9989);
or UO_696 (O_696,N_9962,N_9954);
nand UO_697 (O_697,N_9918,N_9970);
nand UO_698 (O_698,N_9863,N_9800);
xnor UO_699 (O_699,N_9874,N_9888);
and UO_700 (O_700,N_9866,N_9833);
or UO_701 (O_701,N_9889,N_9820);
nand UO_702 (O_702,N_9955,N_9898);
xor UO_703 (O_703,N_9902,N_9973);
and UO_704 (O_704,N_9918,N_9846);
xor UO_705 (O_705,N_9988,N_9842);
and UO_706 (O_706,N_9809,N_9966);
and UO_707 (O_707,N_9958,N_9983);
nand UO_708 (O_708,N_9985,N_9993);
and UO_709 (O_709,N_9949,N_9965);
xnor UO_710 (O_710,N_9970,N_9838);
nor UO_711 (O_711,N_9931,N_9852);
or UO_712 (O_712,N_9946,N_9987);
xor UO_713 (O_713,N_9854,N_9962);
xnor UO_714 (O_714,N_9810,N_9967);
nand UO_715 (O_715,N_9879,N_9932);
nand UO_716 (O_716,N_9969,N_9912);
nand UO_717 (O_717,N_9823,N_9966);
nand UO_718 (O_718,N_9821,N_9819);
xnor UO_719 (O_719,N_9861,N_9928);
nand UO_720 (O_720,N_9926,N_9908);
and UO_721 (O_721,N_9830,N_9807);
xor UO_722 (O_722,N_9823,N_9974);
nor UO_723 (O_723,N_9878,N_9915);
nor UO_724 (O_724,N_9816,N_9893);
nor UO_725 (O_725,N_9949,N_9908);
nor UO_726 (O_726,N_9972,N_9879);
or UO_727 (O_727,N_9968,N_9918);
xor UO_728 (O_728,N_9851,N_9827);
or UO_729 (O_729,N_9935,N_9880);
and UO_730 (O_730,N_9803,N_9982);
xnor UO_731 (O_731,N_9974,N_9891);
and UO_732 (O_732,N_9995,N_9852);
nor UO_733 (O_733,N_9937,N_9908);
nor UO_734 (O_734,N_9815,N_9912);
nor UO_735 (O_735,N_9890,N_9886);
nor UO_736 (O_736,N_9864,N_9982);
nor UO_737 (O_737,N_9949,N_9855);
nand UO_738 (O_738,N_9959,N_9926);
and UO_739 (O_739,N_9998,N_9943);
and UO_740 (O_740,N_9937,N_9881);
xnor UO_741 (O_741,N_9868,N_9945);
nor UO_742 (O_742,N_9883,N_9974);
xor UO_743 (O_743,N_9826,N_9912);
nand UO_744 (O_744,N_9852,N_9918);
nand UO_745 (O_745,N_9961,N_9916);
and UO_746 (O_746,N_9983,N_9816);
nor UO_747 (O_747,N_9960,N_9821);
or UO_748 (O_748,N_9885,N_9825);
and UO_749 (O_749,N_9943,N_9840);
nand UO_750 (O_750,N_9831,N_9921);
xnor UO_751 (O_751,N_9962,N_9921);
and UO_752 (O_752,N_9966,N_9850);
nand UO_753 (O_753,N_9823,N_9910);
xnor UO_754 (O_754,N_9855,N_9844);
and UO_755 (O_755,N_9882,N_9909);
nand UO_756 (O_756,N_9874,N_9914);
xnor UO_757 (O_757,N_9979,N_9887);
or UO_758 (O_758,N_9892,N_9924);
or UO_759 (O_759,N_9946,N_9894);
nand UO_760 (O_760,N_9987,N_9843);
nand UO_761 (O_761,N_9959,N_9969);
and UO_762 (O_762,N_9825,N_9805);
nand UO_763 (O_763,N_9955,N_9919);
and UO_764 (O_764,N_9919,N_9809);
nand UO_765 (O_765,N_9912,N_9844);
nor UO_766 (O_766,N_9960,N_9896);
nand UO_767 (O_767,N_9812,N_9803);
and UO_768 (O_768,N_9806,N_9872);
nand UO_769 (O_769,N_9980,N_9808);
and UO_770 (O_770,N_9970,N_9933);
nor UO_771 (O_771,N_9985,N_9915);
and UO_772 (O_772,N_9973,N_9932);
nand UO_773 (O_773,N_9817,N_9829);
or UO_774 (O_774,N_9827,N_9921);
nor UO_775 (O_775,N_9857,N_9948);
nand UO_776 (O_776,N_9889,N_9872);
nand UO_777 (O_777,N_9960,N_9908);
nor UO_778 (O_778,N_9944,N_9829);
and UO_779 (O_779,N_9954,N_9827);
and UO_780 (O_780,N_9819,N_9981);
xnor UO_781 (O_781,N_9836,N_9805);
nand UO_782 (O_782,N_9835,N_9919);
xor UO_783 (O_783,N_9818,N_9927);
nand UO_784 (O_784,N_9839,N_9860);
nor UO_785 (O_785,N_9976,N_9885);
nor UO_786 (O_786,N_9932,N_9980);
nor UO_787 (O_787,N_9801,N_9982);
xnor UO_788 (O_788,N_9840,N_9979);
nor UO_789 (O_789,N_9879,N_9880);
or UO_790 (O_790,N_9917,N_9914);
nor UO_791 (O_791,N_9995,N_9860);
xnor UO_792 (O_792,N_9935,N_9902);
or UO_793 (O_793,N_9972,N_9821);
xor UO_794 (O_794,N_9845,N_9897);
or UO_795 (O_795,N_9922,N_9989);
nor UO_796 (O_796,N_9842,N_9836);
and UO_797 (O_797,N_9826,N_9957);
nand UO_798 (O_798,N_9940,N_9853);
and UO_799 (O_799,N_9948,N_9963);
nand UO_800 (O_800,N_9830,N_9838);
and UO_801 (O_801,N_9943,N_9937);
nand UO_802 (O_802,N_9835,N_9861);
or UO_803 (O_803,N_9863,N_9914);
or UO_804 (O_804,N_9982,N_9989);
nand UO_805 (O_805,N_9851,N_9820);
xnor UO_806 (O_806,N_9933,N_9962);
and UO_807 (O_807,N_9880,N_9858);
and UO_808 (O_808,N_9960,N_9962);
or UO_809 (O_809,N_9989,N_9917);
nor UO_810 (O_810,N_9873,N_9947);
nor UO_811 (O_811,N_9969,N_9856);
xnor UO_812 (O_812,N_9937,N_9985);
nor UO_813 (O_813,N_9833,N_9964);
or UO_814 (O_814,N_9822,N_9805);
or UO_815 (O_815,N_9866,N_9871);
xor UO_816 (O_816,N_9874,N_9926);
and UO_817 (O_817,N_9904,N_9843);
nor UO_818 (O_818,N_9804,N_9984);
and UO_819 (O_819,N_9980,N_9960);
xor UO_820 (O_820,N_9920,N_9945);
nor UO_821 (O_821,N_9851,N_9841);
nor UO_822 (O_822,N_9968,N_9969);
or UO_823 (O_823,N_9983,N_9904);
and UO_824 (O_824,N_9890,N_9991);
nor UO_825 (O_825,N_9999,N_9948);
nor UO_826 (O_826,N_9889,N_9983);
or UO_827 (O_827,N_9849,N_9895);
nor UO_828 (O_828,N_9844,N_9902);
or UO_829 (O_829,N_9884,N_9879);
or UO_830 (O_830,N_9973,N_9925);
nor UO_831 (O_831,N_9831,N_9897);
nor UO_832 (O_832,N_9828,N_9975);
nor UO_833 (O_833,N_9871,N_9827);
and UO_834 (O_834,N_9958,N_9981);
nor UO_835 (O_835,N_9855,N_9843);
or UO_836 (O_836,N_9935,N_9839);
xor UO_837 (O_837,N_9852,N_9890);
nor UO_838 (O_838,N_9818,N_9982);
nand UO_839 (O_839,N_9865,N_9915);
xor UO_840 (O_840,N_9921,N_9850);
xor UO_841 (O_841,N_9842,N_9951);
nor UO_842 (O_842,N_9897,N_9924);
nor UO_843 (O_843,N_9854,N_9874);
nor UO_844 (O_844,N_9869,N_9822);
nand UO_845 (O_845,N_9967,N_9953);
or UO_846 (O_846,N_9882,N_9847);
nor UO_847 (O_847,N_9977,N_9923);
xnor UO_848 (O_848,N_9953,N_9970);
or UO_849 (O_849,N_9870,N_9858);
nand UO_850 (O_850,N_9817,N_9922);
xor UO_851 (O_851,N_9808,N_9926);
and UO_852 (O_852,N_9831,N_9844);
nor UO_853 (O_853,N_9969,N_9853);
and UO_854 (O_854,N_9857,N_9850);
nand UO_855 (O_855,N_9801,N_9802);
and UO_856 (O_856,N_9913,N_9846);
xnor UO_857 (O_857,N_9905,N_9805);
and UO_858 (O_858,N_9973,N_9994);
and UO_859 (O_859,N_9881,N_9915);
and UO_860 (O_860,N_9895,N_9832);
nor UO_861 (O_861,N_9812,N_9818);
nor UO_862 (O_862,N_9948,N_9807);
nand UO_863 (O_863,N_9878,N_9995);
or UO_864 (O_864,N_9916,N_9845);
nor UO_865 (O_865,N_9959,N_9860);
and UO_866 (O_866,N_9808,N_9986);
and UO_867 (O_867,N_9918,N_9861);
nand UO_868 (O_868,N_9935,N_9924);
and UO_869 (O_869,N_9851,N_9962);
and UO_870 (O_870,N_9908,N_9901);
nand UO_871 (O_871,N_9887,N_9913);
and UO_872 (O_872,N_9825,N_9883);
nand UO_873 (O_873,N_9849,N_9922);
or UO_874 (O_874,N_9916,N_9836);
xor UO_875 (O_875,N_9907,N_9918);
xor UO_876 (O_876,N_9895,N_9867);
nand UO_877 (O_877,N_9879,N_9802);
xnor UO_878 (O_878,N_9877,N_9866);
xnor UO_879 (O_879,N_9841,N_9920);
nor UO_880 (O_880,N_9868,N_9940);
or UO_881 (O_881,N_9898,N_9939);
xor UO_882 (O_882,N_9835,N_9809);
nand UO_883 (O_883,N_9820,N_9949);
or UO_884 (O_884,N_9971,N_9906);
or UO_885 (O_885,N_9856,N_9870);
nor UO_886 (O_886,N_9985,N_9972);
nor UO_887 (O_887,N_9887,N_9816);
and UO_888 (O_888,N_9950,N_9845);
and UO_889 (O_889,N_9945,N_9886);
or UO_890 (O_890,N_9882,N_9832);
or UO_891 (O_891,N_9952,N_9868);
nand UO_892 (O_892,N_9889,N_9982);
and UO_893 (O_893,N_9979,N_9984);
or UO_894 (O_894,N_9801,N_9991);
or UO_895 (O_895,N_9976,N_9807);
xnor UO_896 (O_896,N_9915,N_9856);
xnor UO_897 (O_897,N_9958,N_9813);
nor UO_898 (O_898,N_9921,N_9833);
nand UO_899 (O_899,N_9803,N_9969);
xor UO_900 (O_900,N_9938,N_9932);
xor UO_901 (O_901,N_9898,N_9835);
and UO_902 (O_902,N_9963,N_9955);
nand UO_903 (O_903,N_9932,N_9978);
or UO_904 (O_904,N_9976,N_9815);
xor UO_905 (O_905,N_9844,N_9880);
xor UO_906 (O_906,N_9882,N_9952);
xor UO_907 (O_907,N_9956,N_9961);
and UO_908 (O_908,N_9883,N_9887);
xor UO_909 (O_909,N_9947,N_9912);
nand UO_910 (O_910,N_9927,N_9912);
xnor UO_911 (O_911,N_9972,N_9991);
or UO_912 (O_912,N_9956,N_9953);
xnor UO_913 (O_913,N_9963,N_9921);
or UO_914 (O_914,N_9862,N_9834);
nor UO_915 (O_915,N_9891,N_9926);
nor UO_916 (O_916,N_9931,N_9834);
and UO_917 (O_917,N_9950,N_9854);
xor UO_918 (O_918,N_9961,N_9854);
nor UO_919 (O_919,N_9863,N_9806);
or UO_920 (O_920,N_9944,N_9968);
xor UO_921 (O_921,N_9831,N_9840);
and UO_922 (O_922,N_9981,N_9915);
nor UO_923 (O_923,N_9884,N_9924);
or UO_924 (O_924,N_9935,N_9926);
and UO_925 (O_925,N_9921,N_9940);
nor UO_926 (O_926,N_9809,N_9873);
nor UO_927 (O_927,N_9968,N_9899);
xor UO_928 (O_928,N_9928,N_9856);
xor UO_929 (O_929,N_9866,N_9824);
or UO_930 (O_930,N_9995,N_9936);
xnor UO_931 (O_931,N_9899,N_9925);
nand UO_932 (O_932,N_9899,N_9815);
xnor UO_933 (O_933,N_9877,N_9938);
nand UO_934 (O_934,N_9926,N_9829);
nor UO_935 (O_935,N_9854,N_9898);
or UO_936 (O_936,N_9889,N_9908);
nor UO_937 (O_937,N_9900,N_9931);
nor UO_938 (O_938,N_9802,N_9918);
or UO_939 (O_939,N_9805,N_9804);
or UO_940 (O_940,N_9853,N_9856);
nand UO_941 (O_941,N_9992,N_9846);
nand UO_942 (O_942,N_9838,N_9839);
nor UO_943 (O_943,N_9933,N_9885);
nor UO_944 (O_944,N_9903,N_9883);
nor UO_945 (O_945,N_9981,N_9984);
nor UO_946 (O_946,N_9922,N_9957);
nor UO_947 (O_947,N_9892,N_9873);
and UO_948 (O_948,N_9830,N_9822);
and UO_949 (O_949,N_9801,N_9851);
xnor UO_950 (O_950,N_9834,N_9843);
nor UO_951 (O_951,N_9907,N_9812);
nand UO_952 (O_952,N_9858,N_9843);
and UO_953 (O_953,N_9972,N_9947);
nor UO_954 (O_954,N_9982,N_9933);
and UO_955 (O_955,N_9991,N_9996);
and UO_956 (O_956,N_9894,N_9936);
or UO_957 (O_957,N_9992,N_9931);
and UO_958 (O_958,N_9826,N_9810);
nand UO_959 (O_959,N_9842,N_9821);
and UO_960 (O_960,N_9889,N_9913);
nand UO_961 (O_961,N_9823,N_9912);
xor UO_962 (O_962,N_9824,N_9846);
or UO_963 (O_963,N_9919,N_9958);
nor UO_964 (O_964,N_9969,N_9925);
or UO_965 (O_965,N_9811,N_9878);
nand UO_966 (O_966,N_9926,N_9989);
nor UO_967 (O_967,N_9865,N_9960);
and UO_968 (O_968,N_9862,N_9969);
nor UO_969 (O_969,N_9879,N_9807);
and UO_970 (O_970,N_9963,N_9838);
nor UO_971 (O_971,N_9923,N_9849);
xor UO_972 (O_972,N_9929,N_9955);
xnor UO_973 (O_973,N_9843,N_9903);
nor UO_974 (O_974,N_9916,N_9868);
xnor UO_975 (O_975,N_9977,N_9837);
nor UO_976 (O_976,N_9975,N_9972);
xor UO_977 (O_977,N_9956,N_9865);
nor UO_978 (O_978,N_9852,N_9926);
or UO_979 (O_979,N_9860,N_9947);
and UO_980 (O_980,N_9919,N_9859);
and UO_981 (O_981,N_9888,N_9808);
and UO_982 (O_982,N_9946,N_9898);
nor UO_983 (O_983,N_9938,N_9883);
nor UO_984 (O_984,N_9812,N_9955);
nor UO_985 (O_985,N_9933,N_9814);
xor UO_986 (O_986,N_9977,N_9911);
and UO_987 (O_987,N_9808,N_9872);
and UO_988 (O_988,N_9843,N_9871);
nor UO_989 (O_989,N_9879,N_9907);
nor UO_990 (O_990,N_9860,N_9805);
or UO_991 (O_991,N_9838,N_9898);
xor UO_992 (O_992,N_9893,N_9963);
xnor UO_993 (O_993,N_9870,N_9952);
and UO_994 (O_994,N_9983,N_9928);
and UO_995 (O_995,N_9814,N_9951);
or UO_996 (O_996,N_9803,N_9811);
nand UO_997 (O_997,N_9876,N_9948);
or UO_998 (O_998,N_9917,N_9857);
nand UO_999 (O_999,N_9893,N_9847);
and UO_1000 (O_1000,N_9881,N_9926);
nor UO_1001 (O_1001,N_9879,N_9912);
or UO_1002 (O_1002,N_9922,N_9870);
nand UO_1003 (O_1003,N_9919,N_9976);
and UO_1004 (O_1004,N_9983,N_9886);
nor UO_1005 (O_1005,N_9974,N_9811);
nor UO_1006 (O_1006,N_9820,N_9995);
xnor UO_1007 (O_1007,N_9885,N_9991);
xor UO_1008 (O_1008,N_9987,N_9857);
and UO_1009 (O_1009,N_9895,N_9934);
and UO_1010 (O_1010,N_9931,N_9920);
or UO_1011 (O_1011,N_9837,N_9922);
nand UO_1012 (O_1012,N_9961,N_9811);
xor UO_1013 (O_1013,N_9962,N_9915);
nand UO_1014 (O_1014,N_9957,N_9965);
xor UO_1015 (O_1015,N_9879,N_9980);
xor UO_1016 (O_1016,N_9929,N_9865);
and UO_1017 (O_1017,N_9853,N_9923);
and UO_1018 (O_1018,N_9817,N_9894);
nand UO_1019 (O_1019,N_9812,N_9835);
or UO_1020 (O_1020,N_9951,N_9820);
nand UO_1021 (O_1021,N_9914,N_9911);
nand UO_1022 (O_1022,N_9915,N_9964);
or UO_1023 (O_1023,N_9913,N_9961);
and UO_1024 (O_1024,N_9920,N_9833);
xnor UO_1025 (O_1025,N_9875,N_9859);
nand UO_1026 (O_1026,N_9909,N_9881);
and UO_1027 (O_1027,N_9831,N_9830);
xnor UO_1028 (O_1028,N_9803,N_9874);
xnor UO_1029 (O_1029,N_9842,N_9950);
or UO_1030 (O_1030,N_9863,N_9897);
xnor UO_1031 (O_1031,N_9826,N_9817);
nor UO_1032 (O_1032,N_9924,N_9861);
xnor UO_1033 (O_1033,N_9900,N_9885);
or UO_1034 (O_1034,N_9984,N_9887);
nand UO_1035 (O_1035,N_9815,N_9821);
and UO_1036 (O_1036,N_9978,N_9972);
xor UO_1037 (O_1037,N_9928,N_9905);
nand UO_1038 (O_1038,N_9854,N_9978);
nand UO_1039 (O_1039,N_9955,N_9806);
xnor UO_1040 (O_1040,N_9891,N_9896);
and UO_1041 (O_1041,N_9849,N_9896);
nor UO_1042 (O_1042,N_9864,N_9871);
nor UO_1043 (O_1043,N_9998,N_9957);
and UO_1044 (O_1044,N_9948,N_9835);
nor UO_1045 (O_1045,N_9929,N_9895);
nor UO_1046 (O_1046,N_9895,N_9933);
xor UO_1047 (O_1047,N_9976,N_9995);
and UO_1048 (O_1048,N_9897,N_9805);
nand UO_1049 (O_1049,N_9810,N_9801);
and UO_1050 (O_1050,N_9823,N_9860);
or UO_1051 (O_1051,N_9995,N_9965);
nor UO_1052 (O_1052,N_9918,N_9832);
nand UO_1053 (O_1053,N_9822,N_9907);
or UO_1054 (O_1054,N_9975,N_9910);
nor UO_1055 (O_1055,N_9877,N_9922);
nor UO_1056 (O_1056,N_9805,N_9845);
and UO_1057 (O_1057,N_9877,N_9827);
nor UO_1058 (O_1058,N_9910,N_9963);
and UO_1059 (O_1059,N_9927,N_9897);
nor UO_1060 (O_1060,N_9819,N_9841);
or UO_1061 (O_1061,N_9814,N_9913);
xnor UO_1062 (O_1062,N_9945,N_9985);
or UO_1063 (O_1063,N_9912,N_9899);
and UO_1064 (O_1064,N_9848,N_9800);
nor UO_1065 (O_1065,N_9985,N_9997);
and UO_1066 (O_1066,N_9865,N_9977);
or UO_1067 (O_1067,N_9884,N_9833);
or UO_1068 (O_1068,N_9891,N_9906);
and UO_1069 (O_1069,N_9931,N_9853);
nand UO_1070 (O_1070,N_9838,N_9807);
and UO_1071 (O_1071,N_9927,N_9831);
xnor UO_1072 (O_1072,N_9815,N_9811);
or UO_1073 (O_1073,N_9807,N_9990);
or UO_1074 (O_1074,N_9837,N_9821);
xor UO_1075 (O_1075,N_9911,N_9996);
xor UO_1076 (O_1076,N_9861,N_9985);
nand UO_1077 (O_1077,N_9854,N_9972);
and UO_1078 (O_1078,N_9860,N_9986);
and UO_1079 (O_1079,N_9965,N_9851);
and UO_1080 (O_1080,N_9924,N_9839);
nor UO_1081 (O_1081,N_9854,N_9800);
and UO_1082 (O_1082,N_9993,N_9855);
nand UO_1083 (O_1083,N_9871,N_9874);
nand UO_1084 (O_1084,N_9916,N_9919);
nor UO_1085 (O_1085,N_9906,N_9989);
nand UO_1086 (O_1086,N_9867,N_9807);
xnor UO_1087 (O_1087,N_9914,N_9924);
xnor UO_1088 (O_1088,N_9839,N_9918);
nor UO_1089 (O_1089,N_9962,N_9977);
nor UO_1090 (O_1090,N_9853,N_9864);
and UO_1091 (O_1091,N_9826,N_9900);
nor UO_1092 (O_1092,N_9910,N_9829);
and UO_1093 (O_1093,N_9859,N_9942);
and UO_1094 (O_1094,N_9838,N_9822);
and UO_1095 (O_1095,N_9997,N_9934);
nor UO_1096 (O_1096,N_9891,N_9860);
nor UO_1097 (O_1097,N_9866,N_9987);
nor UO_1098 (O_1098,N_9954,N_9895);
nor UO_1099 (O_1099,N_9901,N_9979);
nor UO_1100 (O_1100,N_9938,N_9942);
nor UO_1101 (O_1101,N_9986,N_9910);
nor UO_1102 (O_1102,N_9945,N_9866);
nand UO_1103 (O_1103,N_9939,N_9976);
and UO_1104 (O_1104,N_9888,N_9810);
xnor UO_1105 (O_1105,N_9901,N_9961);
xnor UO_1106 (O_1106,N_9985,N_9847);
or UO_1107 (O_1107,N_9897,N_9933);
and UO_1108 (O_1108,N_9889,N_9976);
or UO_1109 (O_1109,N_9906,N_9941);
or UO_1110 (O_1110,N_9840,N_9958);
xor UO_1111 (O_1111,N_9858,N_9975);
and UO_1112 (O_1112,N_9813,N_9919);
and UO_1113 (O_1113,N_9935,N_9841);
nand UO_1114 (O_1114,N_9896,N_9827);
and UO_1115 (O_1115,N_9877,N_9939);
and UO_1116 (O_1116,N_9815,N_9916);
nor UO_1117 (O_1117,N_9948,N_9989);
or UO_1118 (O_1118,N_9854,N_9897);
xnor UO_1119 (O_1119,N_9974,N_9871);
nor UO_1120 (O_1120,N_9899,N_9964);
or UO_1121 (O_1121,N_9862,N_9850);
or UO_1122 (O_1122,N_9992,N_9811);
nand UO_1123 (O_1123,N_9940,N_9900);
nand UO_1124 (O_1124,N_9972,N_9858);
nand UO_1125 (O_1125,N_9943,N_9936);
nand UO_1126 (O_1126,N_9923,N_9875);
nand UO_1127 (O_1127,N_9889,N_9875);
or UO_1128 (O_1128,N_9876,N_9827);
nand UO_1129 (O_1129,N_9835,N_9982);
nand UO_1130 (O_1130,N_9982,N_9928);
nor UO_1131 (O_1131,N_9918,N_9961);
xnor UO_1132 (O_1132,N_9923,N_9983);
nor UO_1133 (O_1133,N_9850,N_9894);
or UO_1134 (O_1134,N_9975,N_9811);
nor UO_1135 (O_1135,N_9923,N_9893);
xor UO_1136 (O_1136,N_9965,N_9838);
or UO_1137 (O_1137,N_9984,N_9844);
or UO_1138 (O_1138,N_9930,N_9996);
nand UO_1139 (O_1139,N_9839,N_9869);
nand UO_1140 (O_1140,N_9955,N_9849);
or UO_1141 (O_1141,N_9969,N_9825);
and UO_1142 (O_1142,N_9856,N_9829);
nand UO_1143 (O_1143,N_9829,N_9989);
and UO_1144 (O_1144,N_9985,N_9827);
or UO_1145 (O_1145,N_9933,N_9838);
nor UO_1146 (O_1146,N_9828,N_9855);
and UO_1147 (O_1147,N_9979,N_9864);
nand UO_1148 (O_1148,N_9902,N_9864);
or UO_1149 (O_1149,N_9921,N_9816);
nand UO_1150 (O_1150,N_9835,N_9996);
nand UO_1151 (O_1151,N_9949,N_9915);
or UO_1152 (O_1152,N_9810,N_9983);
and UO_1153 (O_1153,N_9971,N_9888);
and UO_1154 (O_1154,N_9896,N_9906);
xnor UO_1155 (O_1155,N_9922,N_9941);
nor UO_1156 (O_1156,N_9833,N_9906);
xor UO_1157 (O_1157,N_9990,N_9806);
and UO_1158 (O_1158,N_9865,N_9985);
and UO_1159 (O_1159,N_9840,N_9808);
nand UO_1160 (O_1160,N_9832,N_9959);
and UO_1161 (O_1161,N_9916,N_9929);
and UO_1162 (O_1162,N_9960,N_9977);
or UO_1163 (O_1163,N_9983,N_9946);
xor UO_1164 (O_1164,N_9985,N_9921);
nor UO_1165 (O_1165,N_9960,N_9961);
nor UO_1166 (O_1166,N_9994,N_9989);
xor UO_1167 (O_1167,N_9929,N_9808);
and UO_1168 (O_1168,N_9959,N_9977);
and UO_1169 (O_1169,N_9894,N_9919);
xor UO_1170 (O_1170,N_9863,N_9852);
or UO_1171 (O_1171,N_9929,N_9961);
xor UO_1172 (O_1172,N_9817,N_9835);
or UO_1173 (O_1173,N_9926,N_9993);
xor UO_1174 (O_1174,N_9942,N_9941);
or UO_1175 (O_1175,N_9901,N_9830);
nand UO_1176 (O_1176,N_9861,N_9811);
or UO_1177 (O_1177,N_9945,N_9898);
or UO_1178 (O_1178,N_9816,N_9928);
xor UO_1179 (O_1179,N_9890,N_9973);
nand UO_1180 (O_1180,N_9847,N_9914);
nand UO_1181 (O_1181,N_9811,N_9840);
nand UO_1182 (O_1182,N_9862,N_9975);
and UO_1183 (O_1183,N_9845,N_9976);
nor UO_1184 (O_1184,N_9891,N_9872);
and UO_1185 (O_1185,N_9804,N_9844);
and UO_1186 (O_1186,N_9851,N_9942);
nor UO_1187 (O_1187,N_9913,N_9803);
nand UO_1188 (O_1188,N_9865,N_9948);
and UO_1189 (O_1189,N_9952,N_9849);
xnor UO_1190 (O_1190,N_9891,N_9936);
nand UO_1191 (O_1191,N_9830,N_9979);
xnor UO_1192 (O_1192,N_9923,N_9901);
nor UO_1193 (O_1193,N_9839,N_9892);
or UO_1194 (O_1194,N_9986,N_9942);
xnor UO_1195 (O_1195,N_9946,N_9933);
nand UO_1196 (O_1196,N_9889,N_9890);
or UO_1197 (O_1197,N_9938,N_9891);
nand UO_1198 (O_1198,N_9991,N_9863);
nor UO_1199 (O_1199,N_9927,N_9802);
or UO_1200 (O_1200,N_9944,N_9860);
and UO_1201 (O_1201,N_9805,N_9890);
nand UO_1202 (O_1202,N_9815,N_9958);
xor UO_1203 (O_1203,N_9853,N_9802);
nor UO_1204 (O_1204,N_9861,N_9900);
xor UO_1205 (O_1205,N_9933,N_9815);
or UO_1206 (O_1206,N_9835,N_9880);
xor UO_1207 (O_1207,N_9837,N_9931);
and UO_1208 (O_1208,N_9904,N_9997);
and UO_1209 (O_1209,N_9993,N_9982);
nor UO_1210 (O_1210,N_9996,N_9851);
nor UO_1211 (O_1211,N_9977,N_9856);
nand UO_1212 (O_1212,N_9832,N_9940);
xnor UO_1213 (O_1213,N_9903,N_9858);
nand UO_1214 (O_1214,N_9971,N_9954);
xor UO_1215 (O_1215,N_9915,N_9909);
or UO_1216 (O_1216,N_9876,N_9834);
and UO_1217 (O_1217,N_9840,N_9982);
nand UO_1218 (O_1218,N_9900,N_9906);
nor UO_1219 (O_1219,N_9829,N_9984);
and UO_1220 (O_1220,N_9832,N_9809);
nand UO_1221 (O_1221,N_9936,N_9928);
nand UO_1222 (O_1222,N_9809,N_9801);
or UO_1223 (O_1223,N_9825,N_9872);
and UO_1224 (O_1224,N_9968,N_9896);
nor UO_1225 (O_1225,N_9850,N_9965);
or UO_1226 (O_1226,N_9808,N_9869);
nor UO_1227 (O_1227,N_9930,N_9837);
xor UO_1228 (O_1228,N_9976,N_9887);
xnor UO_1229 (O_1229,N_9849,N_9898);
xnor UO_1230 (O_1230,N_9887,N_9893);
and UO_1231 (O_1231,N_9874,N_9936);
xnor UO_1232 (O_1232,N_9806,N_9971);
and UO_1233 (O_1233,N_9812,N_9895);
and UO_1234 (O_1234,N_9918,N_9867);
xor UO_1235 (O_1235,N_9857,N_9865);
nor UO_1236 (O_1236,N_9983,N_9826);
and UO_1237 (O_1237,N_9962,N_9819);
nor UO_1238 (O_1238,N_9951,N_9911);
and UO_1239 (O_1239,N_9885,N_9918);
and UO_1240 (O_1240,N_9987,N_9863);
and UO_1241 (O_1241,N_9803,N_9832);
nand UO_1242 (O_1242,N_9989,N_9956);
nand UO_1243 (O_1243,N_9853,N_9982);
nand UO_1244 (O_1244,N_9809,N_9889);
or UO_1245 (O_1245,N_9954,N_9979);
nor UO_1246 (O_1246,N_9837,N_9948);
and UO_1247 (O_1247,N_9960,N_9840);
xnor UO_1248 (O_1248,N_9925,N_9935);
nand UO_1249 (O_1249,N_9820,N_9868);
nand UO_1250 (O_1250,N_9947,N_9831);
and UO_1251 (O_1251,N_9942,N_9910);
xor UO_1252 (O_1252,N_9804,N_9999);
or UO_1253 (O_1253,N_9875,N_9943);
nor UO_1254 (O_1254,N_9895,N_9991);
xor UO_1255 (O_1255,N_9876,N_9924);
and UO_1256 (O_1256,N_9818,N_9837);
xor UO_1257 (O_1257,N_9954,N_9830);
or UO_1258 (O_1258,N_9824,N_9913);
xor UO_1259 (O_1259,N_9803,N_9861);
or UO_1260 (O_1260,N_9813,N_9881);
nand UO_1261 (O_1261,N_9968,N_9854);
or UO_1262 (O_1262,N_9881,N_9819);
nor UO_1263 (O_1263,N_9815,N_9817);
or UO_1264 (O_1264,N_9947,N_9805);
xor UO_1265 (O_1265,N_9973,N_9956);
xor UO_1266 (O_1266,N_9809,N_9961);
nor UO_1267 (O_1267,N_9943,N_9871);
nor UO_1268 (O_1268,N_9860,N_9852);
and UO_1269 (O_1269,N_9865,N_9883);
nand UO_1270 (O_1270,N_9890,N_9954);
and UO_1271 (O_1271,N_9832,N_9902);
and UO_1272 (O_1272,N_9817,N_9839);
and UO_1273 (O_1273,N_9989,N_9803);
and UO_1274 (O_1274,N_9888,N_9930);
and UO_1275 (O_1275,N_9936,N_9890);
nand UO_1276 (O_1276,N_9963,N_9972);
xnor UO_1277 (O_1277,N_9994,N_9905);
nand UO_1278 (O_1278,N_9907,N_9842);
and UO_1279 (O_1279,N_9881,N_9873);
xnor UO_1280 (O_1280,N_9831,N_9810);
nand UO_1281 (O_1281,N_9947,N_9826);
and UO_1282 (O_1282,N_9941,N_9961);
nand UO_1283 (O_1283,N_9857,N_9977);
or UO_1284 (O_1284,N_9814,N_9968);
nand UO_1285 (O_1285,N_9976,N_9827);
and UO_1286 (O_1286,N_9860,N_9965);
nand UO_1287 (O_1287,N_9942,N_9950);
nor UO_1288 (O_1288,N_9829,N_9870);
xor UO_1289 (O_1289,N_9890,N_9825);
or UO_1290 (O_1290,N_9976,N_9819);
or UO_1291 (O_1291,N_9884,N_9808);
nor UO_1292 (O_1292,N_9899,N_9860);
nor UO_1293 (O_1293,N_9804,N_9947);
nand UO_1294 (O_1294,N_9852,N_9901);
nor UO_1295 (O_1295,N_9881,N_9875);
and UO_1296 (O_1296,N_9830,N_9882);
nor UO_1297 (O_1297,N_9924,N_9811);
nand UO_1298 (O_1298,N_9875,N_9949);
xor UO_1299 (O_1299,N_9869,N_9937);
xor UO_1300 (O_1300,N_9926,N_9972);
nor UO_1301 (O_1301,N_9983,N_9820);
and UO_1302 (O_1302,N_9989,N_9872);
nor UO_1303 (O_1303,N_9985,N_9823);
or UO_1304 (O_1304,N_9965,N_9912);
and UO_1305 (O_1305,N_9999,N_9933);
xnor UO_1306 (O_1306,N_9878,N_9941);
xor UO_1307 (O_1307,N_9910,N_9856);
and UO_1308 (O_1308,N_9813,N_9978);
xnor UO_1309 (O_1309,N_9953,N_9884);
xnor UO_1310 (O_1310,N_9917,N_9807);
or UO_1311 (O_1311,N_9913,N_9839);
xor UO_1312 (O_1312,N_9970,N_9978);
xnor UO_1313 (O_1313,N_9973,N_9816);
nor UO_1314 (O_1314,N_9867,N_9824);
nand UO_1315 (O_1315,N_9918,N_9828);
xnor UO_1316 (O_1316,N_9854,N_9940);
and UO_1317 (O_1317,N_9928,N_9956);
nand UO_1318 (O_1318,N_9862,N_9882);
and UO_1319 (O_1319,N_9878,N_9822);
or UO_1320 (O_1320,N_9865,N_9806);
or UO_1321 (O_1321,N_9855,N_9873);
and UO_1322 (O_1322,N_9869,N_9854);
xnor UO_1323 (O_1323,N_9896,N_9946);
xnor UO_1324 (O_1324,N_9880,N_9997);
xor UO_1325 (O_1325,N_9925,N_9932);
and UO_1326 (O_1326,N_9978,N_9865);
nand UO_1327 (O_1327,N_9849,N_9861);
nand UO_1328 (O_1328,N_9862,N_9967);
and UO_1329 (O_1329,N_9864,N_9823);
xnor UO_1330 (O_1330,N_9948,N_9888);
xor UO_1331 (O_1331,N_9987,N_9817);
nor UO_1332 (O_1332,N_9872,N_9999);
xnor UO_1333 (O_1333,N_9809,N_9842);
xor UO_1334 (O_1334,N_9860,N_9851);
xor UO_1335 (O_1335,N_9804,N_9865);
and UO_1336 (O_1336,N_9895,N_9972);
and UO_1337 (O_1337,N_9880,N_9910);
nand UO_1338 (O_1338,N_9934,N_9976);
or UO_1339 (O_1339,N_9827,N_9858);
and UO_1340 (O_1340,N_9850,N_9821);
nand UO_1341 (O_1341,N_9868,N_9920);
nor UO_1342 (O_1342,N_9993,N_9962);
or UO_1343 (O_1343,N_9895,N_9913);
or UO_1344 (O_1344,N_9806,N_9864);
or UO_1345 (O_1345,N_9804,N_9953);
nor UO_1346 (O_1346,N_9945,N_9853);
nor UO_1347 (O_1347,N_9994,N_9982);
nand UO_1348 (O_1348,N_9992,N_9858);
and UO_1349 (O_1349,N_9901,N_9982);
nand UO_1350 (O_1350,N_9836,N_9819);
and UO_1351 (O_1351,N_9969,N_9800);
xor UO_1352 (O_1352,N_9920,N_9914);
xor UO_1353 (O_1353,N_9815,N_9968);
nor UO_1354 (O_1354,N_9853,N_9811);
nor UO_1355 (O_1355,N_9908,N_9980);
nand UO_1356 (O_1356,N_9855,N_9827);
xor UO_1357 (O_1357,N_9912,N_9839);
and UO_1358 (O_1358,N_9888,N_9961);
nor UO_1359 (O_1359,N_9869,N_9884);
or UO_1360 (O_1360,N_9841,N_9897);
nand UO_1361 (O_1361,N_9918,N_9879);
and UO_1362 (O_1362,N_9906,N_9936);
or UO_1363 (O_1363,N_9838,N_9813);
and UO_1364 (O_1364,N_9874,N_9924);
and UO_1365 (O_1365,N_9827,N_9915);
nand UO_1366 (O_1366,N_9943,N_9990);
nand UO_1367 (O_1367,N_9996,N_9875);
nor UO_1368 (O_1368,N_9921,N_9915);
nand UO_1369 (O_1369,N_9929,N_9998);
nand UO_1370 (O_1370,N_9878,N_9946);
or UO_1371 (O_1371,N_9827,N_9862);
nand UO_1372 (O_1372,N_9945,N_9958);
or UO_1373 (O_1373,N_9836,N_9807);
nand UO_1374 (O_1374,N_9931,N_9848);
nand UO_1375 (O_1375,N_9846,N_9987);
nand UO_1376 (O_1376,N_9880,N_9807);
nor UO_1377 (O_1377,N_9897,N_9921);
nor UO_1378 (O_1378,N_9831,N_9971);
xnor UO_1379 (O_1379,N_9827,N_9887);
nor UO_1380 (O_1380,N_9994,N_9968);
nor UO_1381 (O_1381,N_9842,N_9858);
xnor UO_1382 (O_1382,N_9880,N_9843);
or UO_1383 (O_1383,N_9949,N_9909);
and UO_1384 (O_1384,N_9837,N_9925);
and UO_1385 (O_1385,N_9856,N_9844);
and UO_1386 (O_1386,N_9859,N_9956);
or UO_1387 (O_1387,N_9826,N_9937);
or UO_1388 (O_1388,N_9948,N_9844);
or UO_1389 (O_1389,N_9899,N_9812);
nor UO_1390 (O_1390,N_9817,N_9842);
and UO_1391 (O_1391,N_9840,N_9842);
xor UO_1392 (O_1392,N_9820,N_9809);
nor UO_1393 (O_1393,N_9851,N_9926);
nand UO_1394 (O_1394,N_9822,N_9983);
xor UO_1395 (O_1395,N_9901,N_9859);
and UO_1396 (O_1396,N_9813,N_9831);
nand UO_1397 (O_1397,N_9871,N_9828);
or UO_1398 (O_1398,N_9881,N_9856);
nor UO_1399 (O_1399,N_9961,N_9860);
and UO_1400 (O_1400,N_9975,N_9994);
nor UO_1401 (O_1401,N_9964,N_9992);
or UO_1402 (O_1402,N_9899,N_9976);
nor UO_1403 (O_1403,N_9899,N_9926);
xor UO_1404 (O_1404,N_9879,N_9938);
nor UO_1405 (O_1405,N_9864,N_9962);
or UO_1406 (O_1406,N_9889,N_9801);
xor UO_1407 (O_1407,N_9989,N_9968);
nand UO_1408 (O_1408,N_9976,N_9812);
nor UO_1409 (O_1409,N_9944,N_9924);
nor UO_1410 (O_1410,N_9846,N_9891);
nand UO_1411 (O_1411,N_9877,N_9975);
and UO_1412 (O_1412,N_9997,N_9943);
nand UO_1413 (O_1413,N_9950,N_9849);
nand UO_1414 (O_1414,N_9935,N_9832);
and UO_1415 (O_1415,N_9918,N_9949);
and UO_1416 (O_1416,N_9844,N_9881);
nor UO_1417 (O_1417,N_9947,N_9911);
nor UO_1418 (O_1418,N_9882,N_9908);
nand UO_1419 (O_1419,N_9915,N_9855);
xnor UO_1420 (O_1420,N_9921,N_9972);
xor UO_1421 (O_1421,N_9936,N_9857);
xnor UO_1422 (O_1422,N_9804,N_9854);
nand UO_1423 (O_1423,N_9875,N_9902);
or UO_1424 (O_1424,N_9900,N_9929);
nor UO_1425 (O_1425,N_9922,N_9868);
and UO_1426 (O_1426,N_9954,N_9959);
and UO_1427 (O_1427,N_9855,N_9874);
nand UO_1428 (O_1428,N_9868,N_9918);
nand UO_1429 (O_1429,N_9963,N_9872);
nand UO_1430 (O_1430,N_9986,N_9960);
and UO_1431 (O_1431,N_9845,N_9846);
nand UO_1432 (O_1432,N_9976,N_9838);
nor UO_1433 (O_1433,N_9821,N_9810);
nand UO_1434 (O_1434,N_9930,N_9816);
or UO_1435 (O_1435,N_9808,N_9815);
or UO_1436 (O_1436,N_9872,N_9898);
xor UO_1437 (O_1437,N_9929,N_9878);
nand UO_1438 (O_1438,N_9871,N_9814);
and UO_1439 (O_1439,N_9943,N_9897);
nand UO_1440 (O_1440,N_9880,N_9964);
xnor UO_1441 (O_1441,N_9820,N_9833);
and UO_1442 (O_1442,N_9933,N_9919);
and UO_1443 (O_1443,N_9969,N_9949);
xnor UO_1444 (O_1444,N_9932,N_9800);
xor UO_1445 (O_1445,N_9801,N_9942);
nand UO_1446 (O_1446,N_9991,N_9924);
nor UO_1447 (O_1447,N_9878,N_9817);
nor UO_1448 (O_1448,N_9834,N_9898);
and UO_1449 (O_1449,N_9967,N_9987);
nand UO_1450 (O_1450,N_9857,N_9943);
nand UO_1451 (O_1451,N_9971,N_9809);
or UO_1452 (O_1452,N_9934,N_9816);
or UO_1453 (O_1453,N_9873,N_9834);
nand UO_1454 (O_1454,N_9815,N_9896);
or UO_1455 (O_1455,N_9988,N_9975);
and UO_1456 (O_1456,N_9903,N_9835);
nor UO_1457 (O_1457,N_9920,N_9990);
and UO_1458 (O_1458,N_9994,N_9876);
nand UO_1459 (O_1459,N_9892,N_9821);
or UO_1460 (O_1460,N_9815,N_9830);
or UO_1461 (O_1461,N_9893,N_9857);
or UO_1462 (O_1462,N_9905,N_9855);
nor UO_1463 (O_1463,N_9972,N_9933);
and UO_1464 (O_1464,N_9987,N_9964);
nand UO_1465 (O_1465,N_9929,N_9834);
xnor UO_1466 (O_1466,N_9902,N_9907);
xor UO_1467 (O_1467,N_9943,N_9891);
and UO_1468 (O_1468,N_9922,N_9884);
xnor UO_1469 (O_1469,N_9896,N_9873);
xor UO_1470 (O_1470,N_9849,N_9962);
nand UO_1471 (O_1471,N_9967,N_9840);
or UO_1472 (O_1472,N_9982,N_9879);
and UO_1473 (O_1473,N_9880,N_9947);
and UO_1474 (O_1474,N_9986,N_9801);
or UO_1475 (O_1475,N_9944,N_9819);
nor UO_1476 (O_1476,N_9849,N_9846);
or UO_1477 (O_1477,N_9807,N_9863);
and UO_1478 (O_1478,N_9963,N_9816);
or UO_1479 (O_1479,N_9938,N_9917);
nand UO_1480 (O_1480,N_9875,N_9846);
and UO_1481 (O_1481,N_9936,N_9927);
or UO_1482 (O_1482,N_9823,N_9815);
nor UO_1483 (O_1483,N_9866,N_9838);
xnor UO_1484 (O_1484,N_9910,N_9943);
nand UO_1485 (O_1485,N_9839,N_9819);
xnor UO_1486 (O_1486,N_9927,N_9856);
xnor UO_1487 (O_1487,N_9952,N_9887);
nand UO_1488 (O_1488,N_9858,N_9878);
nand UO_1489 (O_1489,N_9854,N_9829);
nand UO_1490 (O_1490,N_9957,N_9912);
nand UO_1491 (O_1491,N_9882,N_9931);
nor UO_1492 (O_1492,N_9832,N_9999);
and UO_1493 (O_1493,N_9991,N_9873);
xor UO_1494 (O_1494,N_9926,N_9951);
xor UO_1495 (O_1495,N_9827,N_9904);
nor UO_1496 (O_1496,N_9867,N_9904);
xnor UO_1497 (O_1497,N_9837,N_9891);
nor UO_1498 (O_1498,N_9854,N_9827);
xnor UO_1499 (O_1499,N_9931,N_9970);
endmodule