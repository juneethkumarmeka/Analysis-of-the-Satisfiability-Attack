module basic_500_3000_500_5_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_147,In_453);
and U1 (N_1,In_298,In_3);
nand U2 (N_2,In_431,In_376);
and U3 (N_3,In_167,In_483);
and U4 (N_4,In_477,In_427);
nor U5 (N_5,In_449,In_425);
nor U6 (N_6,In_29,In_98);
or U7 (N_7,In_469,In_417);
and U8 (N_8,In_239,In_462);
nor U9 (N_9,In_6,In_319);
or U10 (N_10,In_74,In_198);
nand U11 (N_11,In_341,In_475);
nor U12 (N_12,In_36,In_303);
and U13 (N_13,In_480,In_384);
and U14 (N_14,In_33,In_150);
or U15 (N_15,In_85,In_117);
or U16 (N_16,In_240,In_163);
and U17 (N_17,In_368,In_402);
and U18 (N_18,In_44,In_329);
nand U19 (N_19,In_166,In_424);
or U20 (N_20,In_474,In_231);
and U21 (N_21,In_331,In_126);
or U22 (N_22,In_356,In_302);
xnor U23 (N_23,In_178,In_419);
nor U24 (N_24,In_103,In_313);
or U25 (N_25,In_165,In_411);
or U26 (N_26,In_172,In_413);
nand U27 (N_27,In_288,In_53);
nand U28 (N_28,In_437,In_268);
or U29 (N_29,In_225,In_87);
and U30 (N_30,In_242,In_311);
nor U31 (N_31,In_333,In_304);
and U32 (N_32,In_12,In_9);
nand U33 (N_33,In_406,In_70);
nor U34 (N_34,In_233,In_359);
and U35 (N_35,In_305,In_111);
nand U36 (N_36,In_461,In_248);
nor U37 (N_37,In_39,In_364);
nand U38 (N_38,In_256,In_317);
nand U39 (N_39,In_57,In_50);
nand U40 (N_40,In_360,In_199);
or U41 (N_41,In_306,In_129);
and U42 (N_42,In_105,In_79);
or U43 (N_43,In_136,In_328);
nand U44 (N_44,In_69,In_255);
or U45 (N_45,In_18,In_389);
nor U46 (N_46,In_102,In_206);
nor U47 (N_47,In_337,In_4);
and U48 (N_48,In_435,In_373);
nand U49 (N_49,In_326,In_75);
nand U50 (N_50,In_68,In_309);
nor U51 (N_51,In_452,In_492);
or U52 (N_52,In_34,In_446);
and U53 (N_53,In_344,In_214);
nand U54 (N_54,In_334,In_161);
nand U55 (N_55,In_442,In_276);
and U56 (N_56,In_350,In_149);
and U57 (N_57,In_390,In_301);
nand U58 (N_58,In_321,In_310);
and U59 (N_59,In_164,In_473);
and U60 (N_60,In_491,In_124);
nand U61 (N_61,In_349,In_260);
and U62 (N_62,In_316,In_108);
and U63 (N_63,In_335,In_134);
and U64 (N_64,In_488,In_84);
nand U65 (N_65,In_155,In_495);
nor U66 (N_66,In_455,In_81);
nor U67 (N_67,In_434,In_210);
nand U68 (N_68,In_386,In_369);
xor U69 (N_69,In_433,In_485);
nor U70 (N_70,In_238,In_408);
nor U71 (N_71,In_300,In_380);
or U72 (N_72,In_374,In_202);
and U73 (N_73,In_467,In_92);
nand U74 (N_74,In_464,In_418);
or U75 (N_75,In_459,In_466);
or U76 (N_76,In_141,In_25);
or U77 (N_77,In_381,In_215);
nand U78 (N_78,In_254,In_354);
xnor U79 (N_79,In_139,In_51);
and U80 (N_80,In_5,In_95);
and U81 (N_81,In_426,In_89);
and U82 (N_82,In_403,In_274);
and U83 (N_83,In_100,In_358);
nand U84 (N_84,In_365,In_460);
and U85 (N_85,In_383,In_441);
nor U86 (N_86,In_97,In_193);
or U87 (N_87,In_192,In_204);
nand U88 (N_88,In_497,In_8);
and U89 (N_89,In_11,In_387);
xor U90 (N_90,In_211,In_338);
nand U91 (N_91,In_52,In_289);
and U92 (N_92,In_325,In_38);
or U93 (N_93,In_294,In_388);
and U94 (N_94,In_340,In_203);
nand U95 (N_95,In_451,In_315);
and U96 (N_96,In_363,In_138);
and U97 (N_97,In_130,In_470);
or U98 (N_98,In_284,In_379);
and U99 (N_99,In_96,In_246);
nand U100 (N_100,In_185,In_42);
nor U101 (N_101,In_1,In_207);
and U102 (N_102,In_20,In_237);
or U103 (N_103,In_24,In_16);
or U104 (N_104,In_73,In_481);
nand U105 (N_105,In_83,In_266);
nor U106 (N_106,In_220,In_106);
nor U107 (N_107,In_72,In_450);
nand U108 (N_108,In_375,In_279);
nor U109 (N_109,In_421,In_489);
and U110 (N_110,In_296,In_120);
nor U111 (N_111,In_448,In_235);
nand U112 (N_112,In_241,In_482);
and U113 (N_113,In_41,In_184);
nor U114 (N_114,In_320,In_159);
nand U115 (N_115,In_152,In_228);
xnor U116 (N_116,In_262,In_345);
nor U117 (N_117,In_196,In_158);
and U118 (N_118,In_393,In_420);
and U119 (N_119,In_394,In_348);
nand U120 (N_120,In_324,In_292);
and U121 (N_121,In_456,In_314);
nor U122 (N_122,In_49,In_176);
nor U123 (N_123,In_430,In_145);
or U124 (N_124,In_143,In_447);
and U125 (N_125,In_107,In_55);
nand U126 (N_126,In_367,In_253);
and U127 (N_127,In_259,In_342);
and U128 (N_128,In_61,In_281);
xor U129 (N_129,In_62,In_195);
or U130 (N_130,In_217,In_128);
nand U131 (N_131,In_398,In_131);
and U132 (N_132,In_308,In_287);
and U133 (N_133,In_127,In_30);
nand U134 (N_134,In_370,In_436);
nor U135 (N_135,In_490,In_249);
or U136 (N_136,In_409,In_372);
or U137 (N_137,In_88,In_397);
or U138 (N_138,In_137,In_362);
nor U139 (N_139,In_60,In_201);
or U140 (N_140,In_361,In_188);
or U141 (N_141,In_168,In_382);
or U142 (N_142,In_343,In_10);
nor U143 (N_143,In_54,In_280);
or U144 (N_144,In_91,In_132);
nand U145 (N_145,In_357,In_438);
and U146 (N_146,In_114,In_77);
and U147 (N_147,In_125,In_479);
nor U148 (N_148,In_19,In_58);
nor U149 (N_149,In_400,In_80);
or U150 (N_150,In_282,In_135);
nor U151 (N_151,In_189,In_458);
and U152 (N_152,In_258,In_251);
nand U153 (N_153,In_347,In_429);
nand U154 (N_154,In_187,In_140);
nand U155 (N_155,In_46,In_322);
nor U156 (N_156,In_269,In_67);
nor U157 (N_157,In_121,In_378);
nor U158 (N_158,In_227,In_267);
nor U159 (N_159,In_86,In_21);
and U160 (N_160,In_224,In_116);
nor U161 (N_161,In_415,In_190);
and U162 (N_162,In_133,In_410);
and U163 (N_163,In_56,In_414);
nand U164 (N_164,In_277,In_498);
nand U165 (N_165,In_428,In_396);
or U166 (N_166,In_48,In_0);
or U167 (N_167,In_43,In_177);
and U168 (N_168,In_35,In_407);
or U169 (N_169,In_422,In_232);
or U170 (N_170,In_318,In_154);
nor U171 (N_171,In_17,In_297);
or U172 (N_172,In_160,In_229);
or U173 (N_173,In_47,In_353);
and U174 (N_174,In_40,In_494);
and U175 (N_175,In_183,In_440);
or U176 (N_176,In_271,In_2);
and U177 (N_177,In_366,In_23);
xnor U178 (N_178,In_291,In_286);
and U179 (N_179,In_186,In_493);
nand U180 (N_180,In_323,In_499);
nor U181 (N_181,In_275,In_327);
or U182 (N_182,In_299,In_162);
nand U183 (N_183,In_222,In_226);
and U184 (N_184,In_486,In_454);
nor U185 (N_185,In_463,In_257);
or U186 (N_186,In_157,In_351);
or U187 (N_187,In_295,In_261);
nand U188 (N_188,In_330,In_307);
nand U189 (N_189,In_15,In_148);
nand U190 (N_190,In_173,In_346);
or U191 (N_191,In_37,In_405);
nand U192 (N_192,In_151,In_423);
or U193 (N_193,In_399,In_401);
and U194 (N_194,In_170,In_182);
and U195 (N_195,In_278,In_243);
nor U196 (N_196,In_213,In_478);
nor U197 (N_197,In_416,In_156);
or U198 (N_198,In_13,In_153);
or U199 (N_199,In_412,In_283);
nand U200 (N_200,In_285,In_94);
nand U201 (N_201,In_395,In_28);
nand U202 (N_202,In_31,In_45);
or U203 (N_203,In_212,In_312);
nor U204 (N_204,In_216,In_22);
nand U205 (N_205,In_219,In_336);
nand U206 (N_206,In_122,In_355);
and U207 (N_207,In_487,In_208);
nand U208 (N_208,In_109,In_468);
nand U209 (N_209,In_465,In_90);
and U210 (N_210,In_247,In_123);
or U211 (N_211,In_339,In_293);
nand U212 (N_212,In_146,In_444);
or U213 (N_213,In_223,In_179);
nand U214 (N_214,In_236,In_265);
nand U215 (N_215,In_244,In_273);
nor U216 (N_216,In_119,In_270);
and U217 (N_217,In_26,In_7);
nor U218 (N_218,In_64,In_332);
and U219 (N_219,In_230,In_218);
and U220 (N_220,In_371,In_252);
nor U221 (N_221,In_404,In_352);
nor U222 (N_222,In_144,In_197);
nor U223 (N_223,In_191,In_180);
and U224 (N_224,In_221,In_264);
or U225 (N_225,In_110,In_457);
or U226 (N_226,In_209,In_377);
nor U227 (N_227,In_171,In_194);
nand U228 (N_228,In_476,In_115);
nor U229 (N_229,In_290,In_118);
or U230 (N_230,In_112,In_78);
and U231 (N_231,In_263,In_432);
and U232 (N_232,In_445,In_113);
nand U233 (N_233,In_66,In_471);
and U234 (N_234,In_272,In_63);
nand U235 (N_235,In_93,In_169);
nand U236 (N_236,In_472,In_245);
or U237 (N_237,In_71,In_391);
nor U238 (N_238,In_27,In_175);
or U239 (N_239,In_76,In_250);
or U240 (N_240,In_99,In_439);
or U241 (N_241,In_234,In_82);
or U242 (N_242,In_65,In_14);
nor U243 (N_243,In_443,In_385);
or U244 (N_244,In_205,In_104);
xor U245 (N_245,In_496,In_484);
or U246 (N_246,In_174,In_181);
nor U247 (N_247,In_101,In_59);
and U248 (N_248,In_392,In_142);
nand U249 (N_249,In_32,In_200);
and U250 (N_250,In_69,In_28);
xor U251 (N_251,In_461,In_247);
nand U252 (N_252,In_419,In_415);
nand U253 (N_253,In_137,In_309);
and U254 (N_254,In_13,In_151);
and U255 (N_255,In_411,In_324);
nand U256 (N_256,In_453,In_476);
and U257 (N_257,In_367,In_176);
nand U258 (N_258,In_194,In_379);
and U259 (N_259,In_317,In_476);
nand U260 (N_260,In_401,In_389);
and U261 (N_261,In_294,In_166);
nand U262 (N_262,In_79,In_88);
or U263 (N_263,In_259,In_224);
nor U264 (N_264,In_402,In_289);
or U265 (N_265,In_267,In_445);
or U266 (N_266,In_462,In_102);
and U267 (N_267,In_237,In_457);
or U268 (N_268,In_139,In_188);
nor U269 (N_269,In_8,In_0);
nor U270 (N_270,In_470,In_86);
and U271 (N_271,In_346,In_28);
and U272 (N_272,In_376,In_378);
and U273 (N_273,In_93,In_10);
nand U274 (N_274,In_285,In_458);
and U275 (N_275,In_231,In_36);
or U276 (N_276,In_182,In_390);
or U277 (N_277,In_215,In_34);
or U278 (N_278,In_424,In_387);
and U279 (N_279,In_21,In_198);
nand U280 (N_280,In_405,In_427);
nor U281 (N_281,In_283,In_434);
and U282 (N_282,In_295,In_409);
nand U283 (N_283,In_439,In_203);
nor U284 (N_284,In_232,In_7);
and U285 (N_285,In_266,In_350);
or U286 (N_286,In_96,In_83);
nor U287 (N_287,In_327,In_75);
nand U288 (N_288,In_465,In_305);
nor U289 (N_289,In_322,In_460);
nand U290 (N_290,In_356,In_12);
nor U291 (N_291,In_211,In_278);
nand U292 (N_292,In_350,In_403);
nand U293 (N_293,In_431,In_261);
nor U294 (N_294,In_9,In_281);
nand U295 (N_295,In_435,In_293);
or U296 (N_296,In_472,In_323);
nor U297 (N_297,In_267,In_334);
nor U298 (N_298,In_390,In_392);
and U299 (N_299,In_415,In_336);
and U300 (N_300,In_394,In_52);
and U301 (N_301,In_10,In_250);
nor U302 (N_302,In_308,In_488);
and U303 (N_303,In_393,In_158);
nand U304 (N_304,In_15,In_422);
or U305 (N_305,In_306,In_284);
or U306 (N_306,In_170,In_493);
nor U307 (N_307,In_303,In_77);
nor U308 (N_308,In_382,In_377);
and U309 (N_309,In_116,In_315);
and U310 (N_310,In_6,In_149);
or U311 (N_311,In_203,In_49);
and U312 (N_312,In_438,In_214);
nand U313 (N_313,In_396,In_51);
nand U314 (N_314,In_1,In_28);
and U315 (N_315,In_204,In_265);
or U316 (N_316,In_22,In_447);
and U317 (N_317,In_159,In_90);
nand U318 (N_318,In_415,In_6);
nor U319 (N_319,In_128,In_373);
or U320 (N_320,In_252,In_117);
nand U321 (N_321,In_315,In_275);
and U322 (N_322,In_197,In_427);
and U323 (N_323,In_123,In_4);
nor U324 (N_324,In_52,In_489);
nand U325 (N_325,In_311,In_33);
nor U326 (N_326,In_25,In_46);
nor U327 (N_327,In_499,In_465);
or U328 (N_328,In_188,In_122);
and U329 (N_329,In_315,In_138);
nand U330 (N_330,In_181,In_436);
or U331 (N_331,In_82,In_30);
or U332 (N_332,In_450,In_351);
xnor U333 (N_333,In_248,In_191);
or U334 (N_334,In_268,In_318);
and U335 (N_335,In_246,In_219);
or U336 (N_336,In_138,In_415);
nor U337 (N_337,In_227,In_420);
nand U338 (N_338,In_76,In_278);
nor U339 (N_339,In_342,In_365);
or U340 (N_340,In_384,In_240);
nor U341 (N_341,In_116,In_462);
nand U342 (N_342,In_165,In_79);
and U343 (N_343,In_207,In_445);
and U344 (N_344,In_130,In_17);
or U345 (N_345,In_168,In_162);
or U346 (N_346,In_174,In_483);
nand U347 (N_347,In_60,In_189);
nor U348 (N_348,In_368,In_67);
nand U349 (N_349,In_481,In_485);
nand U350 (N_350,In_424,In_180);
or U351 (N_351,In_23,In_88);
nor U352 (N_352,In_177,In_358);
and U353 (N_353,In_449,In_1);
or U354 (N_354,In_433,In_76);
nand U355 (N_355,In_218,In_331);
and U356 (N_356,In_433,In_355);
or U357 (N_357,In_335,In_436);
or U358 (N_358,In_455,In_166);
nand U359 (N_359,In_48,In_174);
and U360 (N_360,In_71,In_298);
and U361 (N_361,In_316,In_257);
nor U362 (N_362,In_299,In_138);
nand U363 (N_363,In_310,In_385);
nand U364 (N_364,In_205,In_79);
xnor U365 (N_365,In_456,In_290);
or U366 (N_366,In_48,In_76);
nand U367 (N_367,In_109,In_279);
nor U368 (N_368,In_123,In_38);
nand U369 (N_369,In_241,In_20);
and U370 (N_370,In_359,In_134);
nor U371 (N_371,In_495,In_399);
nand U372 (N_372,In_45,In_389);
nand U373 (N_373,In_268,In_232);
nand U374 (N_374,In_331,In_459);
nand U375 (N_375,In_330,In_381);
nor U376 (N_376,In_374,In_182);
or U377 (N_377,In_465,In_128);
xor U378 (N_378,In_422,In_296);
nand U379 (N_379,In_414,In_268);
nand U380 (N_380,In_304,In_156);
nor U381 (N_381,In_214,In_145);
and U382 (N_382,In_327,In_287);
and U383 (N_383,In_275,In_378);
or U384 (N_384,In_19,In_401);
nand U385 (N_385,In_240,In_338);
nand U386 (N_386,In_212,In_242);
nand U387 (N_387,In_99,In_82);
and U388 (N_388,In_137,In_315);
or U389 (N_389,In_198,In_104);
nand U390 (N_390,In_331,In_349);
or U391 (N_391,In_372,In_195);
nand U392 (N_392,In_137,In_421);
and U393 (N_393,In_427,In_33);
or U394 (N_394,In_319,In_401);
or U395 (N_395,In_195,In_220);
or U396 (N_396,In_309,In_266);
or U397 (N_397,In_369,In_192);
nor U398 (N_398,In_176,In_226);
nand U399 (N_399,In_183,In_411);
xnor U400 (N_400,In_308,In_45);
nor U401 (N_401,In_278,In_358);
or U402 (N_402,In_330,In_39);
nand U403 (N_403,In_111,In_317);
or U404 (N_404,In_104,In_193);
nand U405 (N_405,In_23,In_39);
nor U406 (N_406,In_324,In_128);
nand U407 (N_407,In_125,In_289);
or U408 (N_408,In_254,In_440);
or U409 (N_409,In_290,In_100);
nor U410 (N_410,In_484,In_440);
and U411 (N_411,In_397,In_274);
and U412 (N_412,In_413,In_264);
nor U413 (N_413,In_10,In_390);
or U414 (N_414,In_271,In_100);
or U415 (N_415,In_33,In_330);
or U416 (N_416,In_464,In_23);
nor U417 (N_417,In_289,In_489);
nand U418 (N_418,In_316,In_222);
and U419 (N_419,In_488,In_23);
nor U420 (N_420,In_473,In_215);
nand U421 (N_421,In_496,In_142);
and U422 (N_422,In_129,In_494);
nand U423 (N_423,In_56,In_131);
or U424 (N_424,In_78,In_16);
and U425 (N_425,In_284,In_167);
nand U426 (N_426,In_36,In_208);
or U427 (N_427,In_123,In_30);
and U428 (N_428,In_444,In_83);
nand U429 (N_429,In_366,In_153);
and U430 (N_430,In_22,In_372);
or U431 (N_431,In_62,In_29);
or U432 (N_432,In_201,In_99);
nor U433 (N_433,In_60,In_146);
nor U434 (N_434,In_315,In_58);
and U435 (N_435,In_486,In_304);
or U436 (N_436,In_88,In_47);
or U437 (N_437,In_260,In_128);
and U438 (N_438,In_109,In_11);
and U439 (N_439,In_390,In_166);
nor U440 (N_440,In_100,In_431);
nand U441 (N_441,In_199,In_189);
nand U442 (N_442,In_117,In_187);
and U443 (N_443,In_94,In_353);
and U444 (N_444,In_139,In_137);
or U445 (N_445,In_358,In_181);
and U446 (N_446,In_323,In_411);
and U447 (N_447,In_103,In_356);
or U448 (N_448,In_58,In_361);
or U449 (N_449,In_100,In_194);
xnor U450 (N_450,In_93,In_219);
nor U451 (N_451,In_343,In_105);
nand U452 (N_452,In_263,In_359);
nor U453 (N_453,In_211,In_397);
and U454 (N_454,In_303,In_372);
nand U455 (N_455,In_381,In_100);
and U456 (N_456,In_67,In_233);
nand U457 (N_457,In_424,In_441);
nor U458 (N_458,In_348,In_471);
nand U459 (N_459,In_192,In_345);
and U460 (N_460,In_59,In_4);
nor U461 (N_461,In_385,In_164);
and U462 (N_462,In_62,In_464);
nand U463 (N_463,In_365,In_88);
and U464 (N_464,In_82,In_284);
nor U465 (N_465,In_188,In_460);
nand U466 (N_466,In_61,In_190);
nor U467 (N_467,In_26,In_438);
or U468 (N_468,In_352,In_283);
nor U469 (N_469,In_468,In_168);
nor U470 (N_470,In_213,In_275);
and U471 (N_471,In_311,In_268);
or U472 (N_472,In_128,In_329);
nor U473 (N_473,In_389,In_409);
or U474 (N_474,In_59,In_197);
or U475 (N_475,In_438,In_125);
nand U476 (N_476,In_197,In_363);
and U477 (N_477,In_233,In_0);
or U478 (N_478,In_420,In_406);
nor U479 (N_479,In_144,In_446);
and U480 (N_480,In_389,In_289);
nand U481 (N_481,In_137,In_135);
or U482 (N_482,In_341,In_296);
and U483 (N_483,In_354,In_403);
and U484 (N_484,In_220,In_281);
nor U485 (N_485,In_280,In_377);
nand U486 (N_486,In_151,In_386);
nand U487 (N_487,In_183,In_28);
and U488 (N_488,In_421,In_184);
or U489 (N_489,In_297,In_486);
and U490 (N_490,In_10,In_245);
nand U491 (N_491,In_227,In_19);
xor U492 (N_492,In_64,In_290);
nand U493 (N_493,In_41,In_347);
nor U494 (N_494,In_200,In_355);
nand U495 (N_495,In_202,In_352);
or U496 (N_496,In_147,In_318);
or U497 (N_497,In_65,In_471);
and U498 (N_498,In_273,In_33);
nor U499 (N_499,In_102,In_482);
or U500 (N_500,In_233,In_270);
xnor U501 (N_501,In_378,In_499);
or U502 (N_502,In_362,In_96);
nor U503 (N_503,In_305,In_174);
or U504 (N_504,In_10,In_316);
and U505 (N_505,In_61,In_264);
nor U506 (N_506,In_66,In_382);
nand U507 (N_507,In_288,In_490);
nand U508 (N_508,In_445,In_409);
and U509 (N_509,In_498,In_415);
and U510 (N_510,In_119,In_129);
or U511 (N_511,In_106,In_332);
xnor U512 (N_512,In_96,In_81);
or U513 (N_513,In_48,In_449);
nand U514 (N_514,In_246,In_401);
and U515 (N_515,In_362,In_477);
xnor U516 (N_516,In_197,In_131);
nor U517 (N_517,In_216,In_403);
nor U518 (N_518,In_490,In_90);
and U519 (N_519,In_25,In_121);
nand U520 (N_520,In_492,In_249);
and U521 (N_521,In_416,In_18);
and U522 (N_522,In_200,In_297);
nor U523 (N_523,In_102,In_77);
and U524 (N_524,In_481,In_100);
nand U525 (N_525,In_337,In_421);
or U526 (N_526,In_22,In_36);
or U527 (N_527,In_72,In_394);
nor U528 (N_528,In_312,In_197);
or U529 (N_529,In_250,In_326);
nand U530 (N_530,In_134,In_453);
and U531 (N_531,In_163,In_412);
and U532 (N_532,In_490,In_474);
or U533 (N_533,In_174,In_67);
xnor U534 (N_534,In_202,In_491);
xor U535 (N_535,In_247,In_362);
and U536 (N_536,In_284,In_459);
and U537 (N_537,In_276,In_151);
and U538 (N_538,In_119,In_67);
nor U539 (N_539,In_132,In_427);
nor U540 (N_540,In_74,In_415);
nand U541 (N_541,In_368,In_83);
and U542 (N_542,In_495,In_444);
or U543 (N_543,In_167,In_482);
or U544 (N_544,In_271,In_74);
nand U545 (N_545,In_406,In_219);
or U546 (N_546,In_162,In_122);
nor U547 (N_547,In_157,In_120);
and U548 (N_548,In_318,In_123);
nand U549 (N_549,In_72,In_282);
and U550 (N_550,In_410,In_229);
or U551 (N_551,In_133,In_495);
nand U552 (N_552,In_82,In_173);
or U553 (N_553,In_105,In_386);
and U554 (N_554,In_173,In_401);
nand U555 (N_555,In_346,In_481);
nor U556 (N_556,In_140,In_176);
nand U557 (N_557,In_447,In_315);
xnor U558 (N_558,In_443,In_3);
nand U559 (N_559,In_124,In_270);
nand U560 (N_560,In_163,In_397);
and U561 (N_561,In_400,In_297);
nor U562 (N_562,In_482,In_351);
or U563 (N_563,In_249,In_23);
nand U564 (N_564,In_16,In_353);
or U565 (N_565,In_132,In_108);
or U566 (N_566,In_158,In_95);
and U567 (N_567,In_300,In_320);
and U568 (N_568,In_364,In_193);
nand U569 (N_569,In_213,In_259);
nor U570 (N_570,In_245,In_302);
or U571 (N_571,In_171,In_420);
and U572 (N_572,In_337,In_76);
nor U573 (N_573,In_96,In_187);
nand U574 (N_574,In_195,In_442);
or U575 (N_575,In_418,In_301);
or U576 (N_576,In_275,In_32);
or U577 (N_577,In_309,In_397);
or U578 (N_578,In_179,In_252);
or U579 (N_579,In_277,In_29);
nor U580 (N_580,In_213,In_100);
or U581 (N_581,In_319,In_313);
nand U582 (N_582,In_187,In_192);
and U583 (N_583,In_56,In_340);
and U584 (N_584,In_488,In_206);
nor U585 (N_585,In_367,In_335);
nand U586 (N_586,In_92,In_286);
nor U587 (N_587,In_347,In_49);
or U588 (N_588,In_472,In_498);
nand U589 (N_589,In_260,In_79);
xor U590 (N_590,In_364,In_343);
and U591 (N_591,In_451,In_190);
nor U592 (N_592,In_214,In_147);
or U593 (N_593,In_114,In_329);
and U594 (N_594,In_323,In_162);
and U595 (N_595,In_210,In_346);
or U596 (N_596,In_122,In_3);
nor U597 (N_597,In_486,In_257);
nor U598 (N_598,In_454,In_21);
and U599 (N_599,In_12,In_6);
nand U600 (N_600,N_411,N_311);
xnor U601 (N_601,N_442,N_578);
nand U602 (N_602,N_223,N_574);
xnor U603 (N_603,N_191,N_53);
nor U604 (N_604,N_28,N_527);
nand U605 (N_605,N_207,N_392);
nor U606 (N_606,N_219,N_340);
and U607 (N_607,N_593,N_319);
xor U608 (N_608,N_427,N_267);
nor U609 (N_609,N_398,N_355);
or U610 (N_610,N_43,N_93);
nand U611 (N_611,N_499,N_563);
nand U612 (N_612,N_431,N_380);
and U613 (N_613,N_270,N_17);
nor U614 (N_614,N_254,N_146);
and U615 (N_615,N_502,N_14);
and U616 (N_616,N_416,N_540);
nand U617 (N_617,N_297,N_205);
nor U618 (N_618,N_284,N_530);
or U619 (N_619,N_598,N_167);
nor U620 (N_620,N_570,N_389);
xor U621 (N_621,N_538,N_144);
nand U622 (N_622,N_374,N_344);
and U623 (N_623,N_520,N_326);
or U624 (N_624,N_541,N_588);
nor U625 (N_625,N_282,N_20);
nor U626 (N_626,N_34,N_334);
nand U627 (N_627,N_90,N_195);
and U628 (N_628,N_173,N_583);
and U629 (N_629,N_321,N_35);
nand U630 (N_630,N_543,N_368);
and U631 (N_631,N_109,N_187);
nand U632 (N_632,N_57,N_513);
nand U633 (N_633,N_151,N_318);
nand U634 (N_634,N_25,N_115);
nand U635 (N_635,N_573,N_585);
and U636 (N_636,N_479,N_89);
or U637 (N_637,N_100,N_348);
nand U638 (N_638,N_258,N_322);
and U639 (N_639,N_106,N_60);
and U640 (N_640,N_558,N_343);
nor U641 (N_641,N_59,N_303);
nor U642 (N_642,N_256,N_522);
and U643 (N_643,N_568,N_492);
nor U644 (N_644,N_63,N_32);
nor U645 (N_645,N_142,N_189);
xnor U646 (N_646,N_23,N_356);
or U647 (N_647,N_420,N_417);
or U648 (N_648,N_159,N_206);
or U649 (N_649,N_227,N_290);
nand U650 (N_650,N_30,N_208);
nor U651 (N_651,N_122,N_358);
nand U652 (N_652,N_363,N_46);
nor U653 (N_653,N_298,N_504);
and U654 (N_654,N_473,N_87);
nor U655 (N_655,N_529,N_467);
nor U656 (N_656,N_209,N_18);
nand U657 (N_657,N_359,N_266);
nor U658 (N_658,N_350,N_264);
or U659 (N_659,N_535,N_235);
nand U660 (N_660,N_149,N_382);
nand U661 (N_661,N_510,N_413);
nand U662 (N_662,N_73,N_402);
or U663 (N_663,N_460,N_452);
or U664 (N_664,N_346,N_72);
nand U665 (N_665,N_242,N_414);
and U666 (N_666,N_337,N_468);
and U667 (N_667,N_304,N_130);
nand U668 (N_668,N_31,N_472);
nor U669 (N_669,N_58,N_33);
and U670 (N_670,N_203,N_65);
and U671 (N_671,N_103,N_79);
nand U672 (N_672,N_329,N_102);
nand U673 (N_673,N_291,N_86);
and U674 (N_674,N_108,N_199);
xor U675 (N_675,N_105,N_560);
nand U676 (N_676,N_82,N_148);
nand U677 (N_677,N_24,N_566);
and U678 (N_678,N_555,N_4);
and U679 (N_679,N_222,N_596);
or U680 (N_680,N_182,N_478);
and U681 (N_681,N_404,N_474);
and U682 (N_682,N_525,N_327);
or U683 (N_683,N_150,N_331);
or U684 (N_684,N_307,N_325);
or U685 (N_685,N_561,N_459);
and U686 (N_686,N_511,N_597);
nand U687 (N_687,N_455,N_309);
and U688 (N_688,N_381,N_183);
nor U689 (N_689,N_496,N_546);
and U690 (N_690,N_549,N_406);
nand U691 (N_691,N_580,N_260);
or U692 (N_692,N_458,N_456);
or U693 (N_693,N_299,N_582);
and U694 (N_694,N_428,N_202);
nor U695 (N_695,N_412,N_2);
and U696 (N_696,N_579,N_439);
or U697 (N_697,N_247,N_482);
or U698 (N_698,N_237,N_362);
nor U699 (N_699,N_410,N_572);
or U700 (N_700,N_539,N_444);
nor U701 (N_701,N_421,N_295);
nand U702 (N_702,N_367,N_305);
or U703 (N_703,N_172,N_590);
nand U704 (N_704,N_445,N_243);
or U705 (N_705,N_210,N_251);
or U706 (N_706,N_67,N_559);
nand U707 (N_707,N_481,N_567);
and U708 (N_708,N_285,N_551);
or U709 (N_709,N_476,N_391);
and U710 (N_710,N_153,N_193);
or U711 (N_711,N_123,N_438);
and U712 (N_712,N_376,N_75);
nor U713 (N_713,N_261,N_107);
nand U714 (N_714,N_180,N_81);
or U715 (N_715,N_13,N_324);
nand U716 (N_716,N_379,N_516);
nor U717 (N_717,N_451,N_292);
or U718 (N_718,N_250,N_453);
and U719 (N_719,N_253,N_577);
and U720 (N_720,N_232,N_110);
nand U721 (N_721,N_407,N_283);
nand U722 (N_722,N_184,N_587);
and U723 (N_723,N_197,N_211);
nand U724 (N_724,N_276,N_449);
or U725 (N_725,N_220,N_263);
or U726 (N_726,N_228,N_386);
nand U727 (N_727,N_405,N_330);
or U728 (N_728,N_120,N_39);
nand U729 (N_729,N_429,N_308);
nand U730 (N_730,N_104,N_74);
and U731 (N_731,N_19,N_557);
nand U732 (N_732,N_152,N_26);
nand U733 (N_733,N_48,N_171);
or U734 (N_734,N_426,N_338);
nor U735 (N_735,N_8,N_301);
nand U736 (N_736,N_116,N_523);
or U737 (N_737,N_524,N_238);
or U738 (N_738,N_234,N_52);
or U739 (N_739,N_518,N_186);
or U740 (N_740,N_564,N_0);
xnor U741 (N_741,N_378,N_370);
nor U742 (N_742,N_40,N_519);
nand U743 (N_743,N_415,N_514);
and U744 (N_744,N_441,N_395);
and U745 (N_745,N_315,N_138);
or U746 (N_746,N_328,N_181);
and U747 (N_747,N_96,N_506);
or U748 (N_748,N_69,N_169);
and U749 (N_749,N_548,N_259);
or U750 (N_750,N_255,N_168);
and U751 (N_751,N_491,N_517);
and U752 (N_752,N_373,N_268);
and U753 (N_753,N_155,N_36);
or U754 (N_754,N_581,N_88);
or U755 (N_755,N_121,N_469);
nand U756 (N_756,N_157,N_361);
or U757 (N_757,N_226,N_269);
nor U758 (N_758,N_385,N_369);
or U759 (N_759,N_521,N_401);
and U760 (N_760,N_509,N_179);
or U761 (N_761,N_230,N_147);
and U762 (N_762,N_132,N_425);
nor U763 (N_763,N_95,N_281);
nand U764 (N_764,N_38,N_339);
or U765 (N_765,N_351,N_61);
and U766 (N_766,N_317,N_536);
nand U767 (N_767,N_461,N_158);
or U768 (N_768,N_51,N_85);
nor U769 (N_769,N_443,N_200);
and U770 (N_770,N_565,N_400);
and U771 (N_771,N_477,N_508);
nor U772 (N_772,N_434,N_161);
nor U773 (N_773,N_371,N_56);
or U774 (N_774,N_84,N_101);
nand U775 (N_775,N_249,N_165);
and U776 (N_776,N_185,N_77);
and U777 (N_777,N_160,N_9);
or U778 (N_778,N_113,N_224);
nor U779 (N_779,N_133,N_488);
or U780 (N_780,N_7,N_342);
nand U781 (N_781,N_240,N_194);
and U782 (N_782,N_347,N_236);
nor U783 (N_783,N_216,N_277);
or U784 (N_784,N_44,N_125);
and U785 (N_785,N_196,N_366);
nor U786 (N_786,N_534,N_495);
and U787 (N_787,N_372,N_497);
xor U788 (N_788,N_274,N_175);
or U789 (N_789,N_436,N_471);
and U790 (N_790,N_424,N_483);
nor U791 (N_791,N_312,N_225);
nand U792 (N_792,N_248,N_62);
xnor U793 (N_793,N_287,N_569);
nor U794 (N_794,N_515,N_135);
or U795 (N_795,N_537,N_229);
nor U796 (N_796,N_15,N_591);
and U797 (N_797,N_54,N_310);
xnor U798 (N_798,N_599,N_265);
and U799 (N_799,N_71,N_97);
and U800 (N_800,N_198,N_437);
nand U801 (N_801,N_302,N_49);
nand U802 (N_802,N_353,N_545);
or U803 (N_803,N_357,N_447);
or U804 (N_804,N_78,N_393);
nor U805 (N_805,N_475,N_252);
nor U806 (N_806,N_164,N_201);
or U807 (N_807,N_6,N_271);
nor U808 (N_808,N_163,N_141);
nand U809 (N_809,N_76,N_464);
and U810 (N_810,N_112,N_1);
nor U811 (N_811,N_512,N_466);
and U812 (N_812,N_176,N_571);
and U813 (N_813,N_16,N_594);
xnor U814 (N_814,N_245,N_349);
nand U815 (N_815,N_177,N_136);
or U816 (N_816,N_162,N_364);
nor U817 (N_817,N_487,N_231);
nor U818 (N_818,N_531,N_333);
and U819 (N_819,N_463,N_403);
nor U820 (N_820,N_128,N_178);
or U821 (N_821,N_544,N_480);
and U822 (N_822,N_498,N_279);
nor U823 (N_823,N_204,N_239);
nand U824 (N_824,N_306,N_50);
and U825 (N_825,N_589,N_192);
or U826 (N_826,N_432,N_218);
nor U827 (N_827,N_154,N_3);
nor U828 (N_828,N_140,N_12);
and U829 (N_829,N_399,N_505);
and U830 (N_830,N_66,N_91);
or U831 (N_831,N_166,N_503);
and U832 (N_832,N_446,N_99);
or U833 (N_833,N_409,N_419);
nand U834 (N_834,N_134,N_554);
nand U835 (N_835,N_532,N_365);
or U836 (N_836,N_550,N_465);
nor U837 (N_837,N_143,N_280);
nor U838 (N_838,N_332,N_575);
or U839 (N_839,N_22,N_47);
nand U840 (N_840,N_360,N_156);
nor U841 (N_841,N_336,N_42);
or U842 (N_842,N_394,N_390);
xor U843 (N_843,N_119,N_70);
nand U844 (N_844,N_354,N_190);
nor U845 (N_845,N_27,N_5);
nand U846 (N_846,N_387,N_127);
nor U847 (N_847,N_83,N_493);
nand U848 (N_848,N_286,N_526);
nand U849 (N_849,N_556,N_547);
and U850 (N_850,N_430,N_80);
nor U851 (N_851,N_595,N_489);
or U852 (N_852,N_117,N_375);
or U853 (N_853,N_397,N_562);
nand U854 (N_854,N_500,N_507);
nand U855 (N_855,N_462,N_296);
xor U856 (N_856,N_118,N_214);
and U857 (N_857,N_212,N_37);
xnor U858 (N_858,N_422,N_388);
and U859 (N_859,N_542,N_246);
xor U860 (N_860,N_552,N_352);
or U861 (N_861,N_221,N_383);
and U862 (N_862,N_316,N_278);
and U863 (N_863,N_21,N_553);
nand U864 (N_864,N_528,N_289);
and U865 (N_865,N_300,N_94);
nor U866 (N_866,N_418,N_129);
and U867 (N_867,N_188,N_433);
nand U868 (N_868,N_586,N_215);
nand U869 (N_869,N_131,N_244);
nor U870 (N_870,N_275,N_457);
nand U871 (N_871,N_440,N_320);
xor U872 (N_872,N_345,N_533);
nor U873 (N_873,N_11,N_288);
nand U874 (N_874,N_454,N_313);
or U875 (N_875,N_323,N_92);
and U876 (N_876,N_124,N_592);
and U877 (N_877,N_217,N_341);
or U878 (N_878,N_145,N_41);
or U879 (N_879,N_114,N_423);
nand U880 (N_880,N_213,N_448);
nor U881 (N_881,N_314,N_435);
or U882 (N_882,N_29,N_273);
or U883 (N_883,N_584,N_10);
xor U884 (N_884,N_174,N_486);
nand U885 (N_885,N_126,N_257);
or U886 (N_886,N_293,N_470);
nor U887 (N_887,N_45,N_335);
or U888 (N_888,N_377,N_294);
nor U889 (N_889,N_408,N_98);
and U890 (N_890,N_262,N_501);
or U891 (N_891,N_272,N_233);
nand U892 (N_892,N_139,N_111);
or U893 (N_893,N_396,N_484);
nand U894 (N_894,N_576,N_170);
nand U895 (N_895,N_55,N_490);
and U896 (N_896,N_137,N_384);
nor U897 (N_897,N_241,N_494);
or U898 (N_898,N_68,N_485);
nor U899 (N_899,N_450,N_64);
or U900 (N_900,N_133,N_400);
and U901 (N_901,N_555,N_586);
and U902 (N_902,N_259,N_433);
nand U903 (N_903,N_345,N_473);
nand U904 (N_904,N_274,N_270);
xor U905 (N_905,N_450,N_496);
and U906 (N_906,N_151,N_155);
and U907 (N_907,N_334,N_154);
or U908 (N_908,N_509,N_397);
nand U909 (N_909,N_276,N_145);
or U910 (N_910,N_231,N_291);
nand U911 (N_911,N_570,N_559);
nand U912 (N_912,N_351,N_461);
or U913 (N_913,N_105,N_57);
nor U914 (N_914,N_3,N_198);
and U915 (N_915,N_579,N_19);
nor U916 (N_916,N_188,N_314);
xnor U917 (N_917,N_322,N_309);
or U918 (N_918,N_139,N_16);
and U919 (N_919,N_511,N_323);
and U920 (N_920,N_481,N_297);
nand U921 (N_921,N_209,N_34);
nand U922 (N_922,N_179,N_571);
nor U923 (N_923,N_443,N_89);
nor U924 (N_924,N_362,N_235);
xor U925 (N_925,N_417,N_290);
nor U926 (N_926,N_169,N_408);
nand U927 (N_927,N_262,N_447);
nor U928 (N_928,N_301,N_560);
nor U929 (N_929,N_237,N_236);
nand U930 (N_930,N_290,N_62);
nor U931 (N_931,N_226,N_438);
nand U932 (N_932,N_323,N_407);
nand U933 (N_933,N_96,N_138);
and U934 (N_934,N_460,N_537);
nand U935 (N_935,N_233,N_35);
nand U936 (N_936,N_298,N_293);
or U937 (N_937,N_555,N_10);
and U938 (N_938,N_541,N_213);
and U939 (N_939,N_312,N_308);
or U940 (N_940,N_87,N_251);
nor U941 (N_941,N_39,N_93);
nand U942 (N_942,N_267,N_224);
nor U943 (N_943,N_35,N_464);
or U944 (N_944,N_520,N_430);
xor U945 (N_945,N_101,N_249);
nand U946 (N_946,N_101,N_355);
nor U947 (N_947,N_225,N_166);
nor U948 (N_948,N_371,N_180);
nand U949 (N_949,N_488,N_220);
nor U950 (N_950,N_67,N_554);
and U951 (N_951,N_283,N_185);
nand U952 (N_952,N_4,N_9);
or U953 (N_953,N_56,N_316);
and U954 (N_954,N_277,N_103);
nand U955 (N_955,N_97,N_364);
nor U956 (N_956,N_496,N_538);
or U957 (N_957,N_365,N_20);
xor U958 (N_958,N_511,N_214);
and U959 (N_959,N_288,N_9);
or U960 (N_960,N_367,N_560);
or U961 (N_961,N_252,N_314);
or U962 (N_962,N_20,N_138);
or U963 (N_963,N_432,N_119);
nand U964 (N_964,N_32,N_415);
or U965 (N_965,N_117,N_194);
xor U966 (N_966,N_517,N_358);
or U967 (N_967,N_28,N_289);
and U968 (N_968,N_364,N_77);
nor U969 (N_969,N_558,N_181);
nand U970 (N_970,N_3,N_394);
or U971 (N_971,N_261,N_118);
xor U972 (N_972,N_434,N_103);
xor U973 (N_973,N_23,N_290);
nand U974 (N_974,N_530,N_225);
and U975 (N_975,N_84,N_570);
and U976 (N_976,N_580,N_207);
nor U977 (N_977,N_387,N_6);
xnor U978 (N_978,N_95,N_147);
or U979 (N_979,N_524,N_30);
nand U980 (N_980,N_560,N_165);
nand U981 (N_981,N_291,N_394);
and U982 (N_982,N_251,N_160);
nand U983 (N_983,N_20,N_326);
and U984 (N_984,N_559,N_158);
nor U985 (N_985,N_245,N_206);
nand U986 (N_986,N_217,N_561);
and U987 (N_987,N_295,N_405);
nand U988 (N_988,N_373,N_576);
and U989 (N_989,N_94,N_239);
or U990 (N_990,N_59,N_274);
nand U991 (N_991,N_278,N_146);
nor U992 (N_992,N_315,N_142);
and U993 (N_993,N_315,N_13);
nand U994 (N_994,N_16,N_95);
nand U995 (N_995,N_399,N_6);
nor U996 (N_996,N_219,N_575);
or U997 (N_997,N_189,N_514);
nor U998 (N_998,N_579,N_138);
and U999 (N_999,N_471,N_70);
nand U1000 (N_1000,N_0,N_69);
and U1001 (N_1001,N_27,N_236);
nand U1002 (N_1002,N_112,N_190);
xnor U1003 (N_1003,N_433,N_100);
and U1004 (N_1004,N_36,N_349);
and U1005 (N_1005,N_131,N_376);
nand U1006 (N_1006,N_369,N_170);
nand U1007 (N_1007,N_36,N_414);
and U1008 (N_1008,N_465,N_599);
nand U1009 (N_1009,N_528,N_424);
and U1010 (N_1010,N_354,N_60);
and U1011 (N_1011,N_388,N_409);
and U1012 (N_1012,N_184,N_144);
nor U1013 (N_1013,N_185,N_253);
and U1014 (N_1014,N_8,N_1);
and U1015 (N_1015,N_322,N_570);
and U1016 (N_1016,N_246,N_61);
and U1017 (N_1017,N_140,N_150);
or U1018 (N_1018,N_226,N_100);
nor U1019 (N_1019,N_404,N_134);
or U1020 (N_1020,N_81,N_74);
and U1021 (N_1021,N_167,N_596);
or U1022 (N_1022,N_14,N_583);
or U1023 (N_1023,N_35,N_107);
nand U1024 (N_1024,N_196,N_288);
nor U1025 (N_1025,N_377,N_263);
nor U1026 (N_1026,N_375,N_156);
and U1027 (N_1027,N_466,N_505);
or U1028 (N_1028,N_269,N_331);
nand U1029 (N_1029,N_154,N_132);
nor U1030 (N_1030,N_225,N_487);
nand U1031 (N_1031,N_260,N_420);
or U1032 (N_1032,N_141,N_92);
or U1033 (N_1033,N_299,N_557);
nor U1034 (N_1034,N_198,N_540);
and U1035 (N_1035,N_439,N_271);
nand U1036 (N_1036,N_122,N_494);
nand U1037 (N_1037,N_20,N_471);
and U1038 (N_1038,N_124,N_296);
or U1039 (N_1039,N_428,N_51);
xor U1040 (N_1040,N_481,N_214);
nor U1041 (N_1041,N_31,N_174);
and U1042 (N_1042,N_219,N_27);
nor U1043 (N_1043,N_224,N_346);
and U1044 (N_1044,N_492,N_110);
nor U1045 (N_1045,N_445,N_54);
nand U1046 (N_1046,N_504,N_592);
nand U1047 (N_1047,N_298,N_101);
nor U1048 (N_1048,N_10,N_504);
or U1049 (N_1049,N_238,N_561);
nor U1050 (N_1050,N_468,N_593);
nand U1051 (N_1051,N_188,N_431);
or U1052 (N_1052,N_226,N_566);
nand U1053 (N_1053,N_580,N_291);
and U1054 (N_1054,N_348,N_130);
nand U1055 (N_1055,N_123,N_450);
and U1056 (N_1056,N_232,N_218);
nor U1057 (N_1057,N_232,N_44);
or U1058 (N_1058,N_311,N_571);
and U1059 (N_1059,N_157,N_432);
nor U1060 (N_1060,N_51,N_142);
or U1061 (N_1061,N_308,N_244);
nand U1062 (N_1062,N_253,N_159);
or U1063 (N_1063,N_355,N_121);
nor U1064 (N_1064,N_323,N_113);
nor U1065 (N_1065,N_148,N_250);
nor U1066 (N_1066,N_328,N_82);
and U1067 (N_1067,N_352,N_583);
and U1068 (N_1068,N_177,N_502);
or U1069 (N_1069,N_131,N_31);
or U1070 (N_1070,N_231,N_436);
nor U1071 (N_1071,N_386,N_153);
and U1072 (N_1072,N_11,N_306);
and U1073 (N_1073,N_270,N_29);
nand U1074 (N_1074,N_242,N_90);
nor U1075 (N_1075,N_82,N_39);
or U1076 (N_1076,N_165,N_467);
and U1077 (N_1077,N_111,N_60);
or U1078 (N_1078,N_401,N_378);
xnor U1079 (N_1079,N_92,N_367);
nor U1080 (N_1080,N_293,N_114);
nand U1081 (N_1081,N_67,N_233);
or U1082 (N_1082,N_415,N_452);
or U1083 (N_1083,N_31,N_233);
nor U1084 (N_1084,N_159,N_315);
nand U1085 (N_1085,N_204,N_97);
or U1086 (N_1086,N_380,N_186);
or U1087 (N_1087,N_564,N_117);
or U1088 (N_1088,N_445,N_281);
nor U1089 (N_1089,N_145,N_157);
and U1090 (N_1090,N_346,N_512);
nand U1091 (N_1091,N_119,N_329);
xnor U1092 (N_1092,N_57,N_219);
or U1093 (N_1093,N_343,N_485);
and U1094 (N_1094,N_395,N_329);
or U1095 (N_1095,N_288,N_348);
nor U1096 (N_1096,N_379,N_107);
and U1097 (N_1097,N_118,N_520);
nand U1098 (N_1098,N_426,N_347);
and U1099 (N_1099,N_508,N_229);
or U1100 (N_1100,N_253,N_512);
and U1101 (N_1101,N_409,N_321);
or U1102 (N_1102,N_432,N_15);
nor U1103 (N_1103,N_504,N_482);
or U1104 (N_1104,N_437,N_257);
or U1105 (N_1105,N_174,N_497);
nor U1106 (N_1106,N_415,N_547);
nor U1107 (N_1107,N_288,N_239);
and U1108 (N_1108,N_320,N_463);
and U1109 (N_1109,N_449,N_357);
or U1110 (N_1110,N_314,N_78);
nor U1111 (N_1111,N_367,N_242);
xor U1112 (N_1112,N_406,N_111);
or U1113 (N_1113,N_269,N_56);
nor U1114 (N_1114,N_489,N_200);
nor U1115 (N_1115,N_388,N_17);
nor U1116 (N_1116,N_566,N_292);
nor U1117 (N_1117,N_39,N_490);
or U1118 (N_1118,N_593,N_288);
nand U1119 (N_1119,N_363,N_594);
nor U1120 (N_1120,N_385,N_300);
and U1121 (N_1121,N_469,N_560);
nand U1122 (N_1122,N_544,N_493);
or U1123 (N_1123,N_401,N_318);
or U1124 (N_1124,N_61,N_251);
and U1125 (N_1125,N_176,N_301);
and U1126 (N_1126,N_513,N_531);
nor U1127 (N_1127,N_171,N_249);
nor U1128 (N_1128,N_418,N_495);
xnor U1129 (N_1129,N_405,N_39);
nor U1130 (N_1130,N_437,N_295);
or U1131 (N_1131,N_42,N_571);
nand U1132 (N_1132,N_105,N_437);
nor U1133 (N_1133,N_511,N_1);
nor U1134 (N_1134,N_77,N_177);
nor U1135 (N_1135,N_211,N_254);
or U1136 (N_1136,N_63,N_13);
nand U1137 (N_1137,N_394,N_169);
and U1138 (N_1138,N_137,N_298);
and U1139 (N_1139,N_268,N_549);
or U1140 (N_1140,N_413,N_203);
or U1141 (N_1141,N_3,N_266);
nand U1142 (N_1142,N_577,N_121);
and U1143 (N_1143,N_117,N_545);
nand U1144 (N_1144,N_332,N_513);
nand U1145 (N_1145,N_47,N_189);
or U1146 (N_1146,N_76,N_339);
or U1147 (N_1147,N_326,N_583);
and U1148 (N_1148,N_33,N_375);
nand U1149 (N_1149,N_145,N_385);
and U1150 (N_1150,N_244,N_20);
nor U1151 (N_1151,N_339,N_457);
nand U1152 (N_1152,N_585,N_269);
nand U1153 (N_1153,N_227,N_164);
nand U1154 (N_1154,N_94,N_231);
or U1155 (N_1155,N_311,N_466);
nand U1156 (N_1156,N_481,N_310);
or U1157 (N_1157,N_338,N_459);
and U1158 (N_1158,N_331,N_491);
nor U1159 (N_1159,N_515,N_458);
or U1160 (N_1160,N_23,N_530);
nand U1161 (N_1161,N_315,N_340);
nand U1162 (N_1162,N_414,N_251);
and U1163 (N_1163,N_262,N_222);
nand U1164 (N_1164,N_98,N_281);
or U1165 (N_1165,N_379,N_87);
and U1166 (N_1166,N_364,N_583);
and U1167 (N_1167,N_557,N_449);
nand U1168 (N_1168,N_410,N_439);
nor U1169 (N_1169,N_112,N_30);
or U1170 (N_1170,N_354,N_529);
nand U1171 (N_1171,N_556,N_116);
or U1172 (N_1172,N_379,N_464);
or U1173 (N_1173,N_490,N_264);
nand U1174 (N_1174,N_150,N_96);
nor U1175 (N_1175,N_348,N_303);
nor U1176 (N_1176,N_129,N_33);
and U1177 (N_1177,N_354,N_212);
or U1178 (N_1178,N_140,N_442);
nor U1179 (N_1179,N_255,N_582);
and U1180 (N_1180,N_444,N_170);
nor U1181 (N_1181,N_411,N_503);
or U1182 (N_1182,N_144,N_522);
or U1183 (N_1183,N_284,N_565);
and U1184 (N_1184,N_195,N_25);
nand U1185 (N_1185,N_131,N_503);
or U1186 (N_1186,N_5,N_15);
nor U1187 (N_1187,N_249,N_585);
nand U1188 (N_1188,N_544,N_449);
nor U1189 (N_1189,N_591,N_232);
nand U1190 (N_1190,N_582,N_90);
nand U1191 (N_1191,N_318,N_305);
nor U1192 (N_1192,N_507,N_209);
and U1193 (N_1193,N_353,N_4);
nor U1194 (N_1194,N_512,N_151);
nor U1195 (N_1195,N_115,N_44);
nor U1196 (N_1196,N_561,N_118);
or U1197 (N_1197,N_306,N_103);
or U1198 (N_1198,N_430,N_147);
nor U1199 (N_1199,N_259,N_415);
or U1200 (N_1200,N_981,N_694);
nor U1201 (N_1201,N_1080,N_991);
or U1202 (N_1202,N_706,N_768);
nor U1203 (N_1203,N_814,N_720);
or U1204 (N_1204,N_1147,N_773);
nand U1205 (N_1205,N_968,N_942);
nand U1206 (N_1206,N_616,N_961);
nor U1207 (N_1207,N_716,N_827);
nor U1208 (N_1208,N_904,N_841);
nor U1209 (N_1209,N_856,N_691);
nor U1210 (N_1210,N_1008,N_850);
or U1211 (N_1211,N_909,N_703);
xnor U1212 (N_1212,N_869,N_983);
or U1213 (N_1213,N_1104,N_1142);
or U1214 (N_1214,N_969,N_1103);
or U1215 (N_1215,N_656,N_642);
and U1216 (N_1216,N_982,N_1053);
nand U1217 (N_1217,N_820,N_1022);
or U1218 (N_1218,N_821,N_628);
nor U1219 (N_1219,N_1133,N_853);
and U1220 (N_1220,N_1111,N_842);
or U1221 (N_1221,N_621,N_877);
and U1222 (N_1222,N_1191,N_852);
nand U1223 (N_1223,N_1052,N_715);
nand U1224 (N_1224,N_1014,N_844);
nor U1225 (N_1225,N_871,N_947);
nor U1226 (N_1226,N_845,N_746);
nor U1227 (N_1227,N_1000,N_730);
and U1228 (N_1228,N_1027,N_798);
nor U1229 (N_1229,N_708,N_1017);
nor U1230 (N_1230,N_678,N_1062);
nand U1231 (N_1231,N_606,N_625);
nor U1232 (N_1232,N_737,N_879);
or U1233 (N_1233,N_977,N_920);
nand U1234 (N_1234,N_913,N_620);
nor U1235 (N_1235,N_807,N_724);
xor U1236 (N_1236,N_684,N_1106);
and U1237 (N_1237,N_741,N_1109);
nand U1238 (N_1238,N_739,N_902);
and U1239 (N_1239,N_1061,N_1160);
and U1240 (N_1240,N_1116,N_749);
nor U1241 (N_1241,N_808,N_669);
nor U1242 (N_1242,N_661,N_632);
nor U1243 (N_1243,N_1156,N_914);
and U1244 (N_1244,N_915,N_663);
nor U1245 (N_1245,N_613,N_1041);
xnor U1246 (N_1246,N_1150,N_1090);
nand U1247 (N_1247,N_721,N_1197);
xor U1248 (N_1248,N_950,N_674);
nand U1249 (N_1249,N_619,N_1067);
and U1250 (N_1250,N_713,N_908);
and U1251 (N_1251,N_1179,N_757);
or U1252 (N_1252,N_971,N_707);
or U1253 (N_1253,N_1078,N_876);
nand U1254 (N_1254,N_846,N_897);
or U1255 (N_1255,N_782,N_868);
and U1256 (N_1256,N_617,N_847);
nand U1257 (N_1257,N_994,N_1036);
and U1258 (N_1258,N_1066,N_1009);
nand U1259 (N_1259,N_1162,N_1110);
or U1260 (N_1260,N_635,N_819);
nand U1261 (N_1261,N_1007,N_952);
nand U1262 (N_1262,N_733,N_735);
nor U1263 (N_1263,N_818,N_1101);
or U1264 (N_1264,N_673,N_666);
or U1265 (N_1265,N_1087,N_995);
or U1266 (N_1266,N_751,N_1096);
nand U1267 (N_1267,N_833,N_830);
xor U1268 (N_1268,N_917,N_655);
and U1269 (N_1269,N_780,N_788);
xor U1270 (N_1270,N_859,N_1174);
nand U1271 (N_1271,N_797,N_1131);
nor U1272 (N_1272,N_775,N_719);
nor U1273 (N_1273,N_653,N_651);
or U1274 (N_1274,N_1035,N_900);
nor U1275 (N_1275,N_926,N_839);
and U1276 (N_1276,N_989,N_930);
and U1277 (N_1277,N_1178,N_1123);
or U1278 (N_1278,N_1072,N_1049);
nor U1279 (N_1279,N_888,N_993);
and U1280 (N_1280,N_714,N_1166);
nand U1281 (N_1281,N_1070,N_956);
or U1282 (N_1282,N_786,N_829);
nor U1283 (N_1283,N_832,N_1005);
or U1284 (N_1284,N_676,N_1189);
nor U1285 (N_1285,N_1186,N_837);
and U1286 (N_1286,N_857,N_1033);
and U1287 (N_1287,N_664,N_958);
nor U1288 (N_1288,N_967,N_825);
and U1289 (N_1289,N_1056,N_815);
and U1290 (N_1290,N_940,N_802);
or U1291 (N_1291,N_890,N_754);
nand U1292 (N_1292,N_1086,N_903);
nand U1293 (N_1293,N_872,N_1047);
and U1294 (N_1294,N_687,N_864);
nand U1295 (N_1295,N_816,N_1013);
and U1296 (N_1296,N_1089,N_683);
or U1297 (N_1297,N_1012,N_752);
nand U1298 (N_1298,N_791,N_1085);
nor U1299 (N_1299,N_622,N_1184);
and U1300 (N_1300,N_614,N_1190);
nand U1301 (N_1301,N_934,N_863);
and U1302 (N_1302,N_1065,N_1135);
nor U1303 (N_1303,N_1029,N_1032);
and U1304 (N_1304,N_610,N_893);
and U1305 (N_1305,N_718,N_933);
nand U1306 (N_1306,N_1064,N_793);
and U1307 (N_1307,N_759,N_659);
nand U1308 (N_1308,N_1148,N_1141);
nor U1309 (N_1309,N_648,N_1043);
nand U1310 (N_1310,N_608,N_690);
nand U1311 (N_1311,N_1128,N_843);
nand U1312 (N_1312,N_717,N_685);
and U1313 (N_1313,N_1199,N_848);
nor U1314 (N_1314,N_1161,N_826);
nand U1315 (N_1315,N_1016,N_885);
nand U1316 (N_1316,N_725,N_660);
nand U1317 (N_1317,N_1046,N_1112);
and U1318 (N_1318,N_1094,N_889);
or U1319 (N_1319,N_618,N_1028);
nor U1320 (N_1320,N_910,N_729);
and U1321 (N_1321,N_873,N_753);
and U1322 (N_1322,N_1050,N_626);
nor U1323 (N_1323,N_604,N_946);
nand U1324 (N_1324,N_849,N_1076);
nand U1325 (N_1325,N_1113,N_696);
nor U1326 (N_1326,N_1167,N_1175);
and U1327 (N_1327,N_766,N_1192);
nor U1328 (N_1328,N_955,N_627);
nand U1329 (N_1329,N_1138,N_640);
and U1330 (N_1330,N_963,N_1082);
nor U1331 (N_1331,N_1188,N_1118);
nor U1332 (N_1332,N_970,N_763);
nor U1333 (N_1333,N_750,N_945);
or U1334 (N_1334,N_675,N_1127);
or U1335 (N_1335,N_966,N_1193);
or U1336 (N_1336,N_951,N_1074);
nor U1337 (N_1337,N_671,N_810);
and U1338 (N_1338,N_828,N_1018);
nand U1339 (N_1339,N_925,N_886);
nor U1340 (N_1340,N_1020,N_809);
nor U1341 (N_1341,N_1002,N_932);
and U1342 (N_1342,N_665,N_1054);
nor U1343 (N_1343,N_949,N_745);
and U1344 (N_1344,N_1006,N_1187);
nor U1345 (N_1345,N_1095,N_992);
nand U1346 (N_1346,N_1151,N_670);
and U1347 (N_1347,N_633,N_603);
and U1348 (N_1348,N_636,N_1058);
or U1349 (N_1349,N_677,N_974);
or U1350 (N_1350,N_901,N_1099);
and U1351 (N_1351,N_1075,N_1092);
nor U1352 (N_1352,N_858,N_634);
nand U1353 (N_1353,N_1069,N_771);
nor U1354 (N_1354,N_647,N_1137);
and U1355 (N_1355,N_811,N_1119);
nor U1356 (N_1356,N_787,N_1155);
xnor U1357 (N_1357,N_785,N_1145);
nand U1358 (N_1358,N_767,N_672);
nor U1359 (N_1359,N_631,N_605);
nor U1360 (N_1360,N_1068,N_895);
nor U1361 (N_1361,N_1024,N_662);
and U1362 (N_1362,N_1038,N_1117);
nor U1363 (N_1363,N_960,N_792);
or U1364 (N_1364,N_892,N_693);
nor U1365 (N_1365,N_916,N_1158);
nor U1366 (N_1366,N_711,N_1045);
nand U1367 (N_1367,N_1040,N_1180);
or U1368 (N_1368,N_972,N_997);
nand U1369 (N_1369,N_1107,N_806);
or U1370 (N_1370,N_789,N_919);
nand U1371 (N_1371,N_639,N_1176);
and U1372 (N_1372,N_996,N_726);
nor U1373 (N_1373,N_1115,N_629);
nor U1374 (N_1374,N_705,N_1153);
nor U1375 (N_1375,N_747,N_1130);
or U1376 (N_1376,N_1097,N_638);
and U1377 (N_1377,N_681,N_911);
nand U1378 (N_1378,N_883,N_882);
nor U1379 (N_1379,N_1171,N_602);
nand U1380 (N_1380,N_938,N_1026);
nor U1381 (N_1381,N_738,N_1146);
and U1382 (N_1382,N_1181,N_650);
or U1383 (N_1383,N_851,N_1093);
nor U1384 (N_1384,N_1001,N_865);
nand U1385 (N_1385,N_643,N_1154);
or U1386 (N_1386,N_887,N_698);
or U1387 (N_1387,N_1015,N_772);
and U1388 (N_1388,N_1077,N_1037);
nand U1389 (N_1389,N_1168,N_679);
nor U1390 (N_1390,N_601,N_935);
and U1391 (N_1391,N_1102,N_795);
nand U1392 (N_1392,N_990,N_959);
nand U1393 (N_1393,N_1139,N_1083);
nand U1394 (N_1394,N_646,N_1125);
nor U1395 (N_1395,N_762,N_1088);
nor U1396 (N_1396,N_1170,N_878);
and U1397 (N_1397,N_965,N_784);
or U1398 (N_1398,N_800,N_781);
nand U1399 (N_1399,N_701,N_939);
nor U1400 (N_1400,N_998,N_957);
nand U1401 (N_1401,N_831,N_927);
nor U1402 (N_1402,N_861,N_905);
nor U1403 (N_1403,N_898,N_769);
nand U1404 (N_1404,N_697,N_1152);
nor U1405 (N_1405,N_682,N_680);
nand U1406 (N_1406,N_734,N_630);
and U1407 (N_1407,N_838,N_805);
nor U1408 (N_1408,N_931,N_712);
or U1409 (N_1409,N_835,N_756);
or U1410 (N_1410,N_954,N_1149);
xor U1411 (N_1411,N_1194,N_1023);
nand U1412 (N_1412,N_740,N_1132);
nand U1413 (N_1413,N_985,N_723);
nor U1414 (N_1414,N_1122,N_1031);
and U1415 (N_1415,N_645,N_722);
xor U1416 (N_1416,N_1144,N_817);
nand U1417 (N_1417,N_667,N_976);
nand U1418 (N_1418,N_964,N_918);
nor U1419 (N_1419,N_700,N_744);
or U1420 (N_1420,N_803,N_836);
or U1421 (N_1421,N_988,N_1165);
or U1422 (N_1422,N_1048,N_765);
and U1423 (N_1423,N_710,N_922);
and U1424 (N_1424,N_936,N_658);
nand U1425 (N_1425,N_943,N_1060);
nand U1426 (N_1426,N_1120,N_801);
nor U1427 (N_1427,N_906,N_702);
nand U1428 (N_1428,N_728,N_884);
or U1429 (N_1429,N_1195,N_764);
nor U1430 (N_1430,N_1163,N_1055);
or U1431 (N_1431,N_984,N_923);
nand U1432 (N_1432,N_973,N_979);
nor U1433 (N_1433,N_907,N_1051);
nand U1434 (N_1434,N_924,N_777);
or U1435 (N_1435,N_709,N_742);
nand U1436 (N_1436,N_899,N_731);
nor U1437 (N_1437,N_727,N_1091);
xor U1438 (N_1438,N_1098,N_1126);
or U1439 (N_1439,N_774,N_929);
nor U1440 (N_1440,N_1108,N_624);
and U1441 (N_1441,N_875,N_644);
nand U1442 (N_1442,N_980,N_975);
nand U1443 (N_1443,N_1057,N_987);
nor U1444 (N_1444,N_1185,N_822);
nor U1445 (N_1445,N_1182,N_834);
nand U1446 (N_1446,N_688,N_790);
nor U1447 (N_1447,N_804,N_1063);
or U1448 (N_1448,N_1010,N_732);
or U1449 (N_1449,N_761,N_854);
and U1450 (N_1450,N_1173,N_641);
nand U1451 (N_1451,N_1011,N_860);
and U1452 (N_1452,N_1079,N_880);
nor U1453 (N_1453,N_1084,N_652);
xnor U1454 (N_1454,N_812,N_1159);
nand U1455 (N_1455,N_623,N_755);
nor U1456 (N_1456,N_1039,N_986);
and U1457 (N_1457,N_894,N_758);
or U1458 (N_1458,N_600,N_1134);
nand U1459 (N_1459,N_874,N_1059);
or U1460 (N_1460,N_1140,N_609);
and U1461 (N_1461,N_736,N_794);
nor U1462 (N_1462,N_1042,N_689);
nor U1463 (N_1463,N_657,N_912);
nor U1464 (N_1464,N_1183,N_1198);
or U1465 (N_1465,N_855,N_779);
and U1466 (N_1466,N_686,N_699);
nand U1467 (N_1467,N_1196,N_748);
nand U1468 (N_1468,N_978,N_1136);
nor U1469 (N_1469,N_770,N_881);
nand U1470 (N_1470,N_862,N_1019);
xor U1471 (N_1471,N_928,N_1073);
or U1472 (N_1472,N_1044,N_1164);
nor U1473 (N_1473,N_1081,N_896);
nor U1474 (N_1474,N_1121,N_1129);
or U1475 (N_1475,N_776,N_921);
and U1476 (N_1476,N_1114,N_704);
nand U1477 (N_1477,N_867,N_941);
nor U1478 (N_1478,N_778,N_796);
nand U1479 (N_1479,N_607,N_948);
and U1480 (N_1480,N_840,N_760);
or U1481 (N_1481,N_891,N_999);
and U1482 (N_1482,N_615,N_654);
nand U1483 (N_1483,N_743,N_1021);
nor U1484 (N_1484,N_1169,N_668);
or U1485 (N_1485,N_870,N_944);
and U1486 (N_1486,N_1143,N_866);
nor U1487 (N_1487,N_1030,N_1124);
and U1488 (N_1488,N_1025,N_692);
nor U1489 (N_1489,N_612,N_695);
or U1490 (N_1490,N_799,N_1100);
nand U1491 (N_1491,N_1071,N_637);
nor U1492 (N_1492,N_1003,N_813);
nor U1493 (N_1493,N_824,N_1004);
nand U1494 (N_1494,N_649,N_783);
and U1495 (N_1495,N_1034,N_962);
and U1496 (N_1496,N_1177,N_937);
nand U1497 (N_1497,N_1172,N_1157);
nand U1498 (N_1498,N_953,N_611);
or U1499 (N_1499,N_1105,N_823);
xor U1500 (N_1500,N_675,N_1064);
nand U1501 (N_1501,N_1097,N_1006);
or U1502 (N_1502,N_744,N_731);
xnor U1503 (N_1503,N_755,N_827);
nand U1504 (N_1504,N_860,N_1158);
nor U1505 (N_1505,N_1164,N_1028);
xnor U1506 (N_1506,N_1009,N_686);
or U1507 (N_1507,N_1196,N_725);
nand U1508 (N_1508,N_803,N_1194);
xnor U1509 (N_1509,N_955,N_795);
nor U1510 (N_1510,N_930,N_1159);
or U1511 (N_1511,N_822,N_1053);
nand U1512 (N_1512,N_1068,N_1098);
nor U1513 (N_1513,N_1090,N_927);
nor U1514 (N_1514,N_1177,N_674);
or U1515 (N_1515,N_759,N_699);
nor U1516 (N_1516,N_1195,N_696);
xnor U1517 (N_1517,N_841,N_1072);
or U1518 (N_1518,N_644,N_764);
nand U1519 (N_1519,N_922,N_1126);
or U1520 (N_1520,N_881,N_1161);
or U1521 (N_1521,N_1136,N_771);
xnor U1522 (N_1522,N_1183,N_974);
nor U1523 (N_1523,N_972,N_709);
or U1524 (N_1524,N_925,N_1055);
nand U1525 (N_1525,N_882,N_700);
and U1526 (N_1526,N_683,N_961);
nand U1527 (N_1527,N_1198,N_688);
or U1528 (N_1528,N_1079,N_613);
nor U1529 (N_1529,N_1099,N_776);
and U1530 (N_1530,N_1157,N_1086);
and U1531 (N_1531,N_835,N_1170);
or U1532 (N_1532,N_1031,N_667);
nor U1533 (N_1533,N_1182,N_975);
nand U1534 (N_1534,N_926,N_725);
and U1535 (N_1535,N_1187,N_1073);
nor U1536 (N_1536,N_661,N_1032);
xor U1537 (N_1537,N_1174,N_864);
nand U1538 (N_1538,N_999,N_821);
nor U1539 (N_1539,N_864,N_1160);
or U1540 (N_1540,N_875,N_957);
nor U1541 (N_1541,N_1194,N_809);
nand U1542 (N_1542,N_825,N_889);
nand U1543 (N_1543,N_887,N_706);
and U1544 (N_1544,N_932,N_1118);
or U1545 (N_1545,N_1005,N_704);
nand U1546 (N_1546,N_825,N_790);
nand U1547 (N_1547,N_1041,N_839);
nor U1548 (N_1548,N_1186,N_976);
or U1549 (N_1549,N_783,N_1086);
or U1550 (N_1550,N_936,N_861);
or U1551 (N_1551,N_1052,N_1132);
nand U1552 (N_1552,N_1030,N_1026);
nand U1553 (N_1553,N_1158,N_880);
and U1554 (N_1554,N_665,N_859);
or U1555 (N_1555,N_624,N_704);
and U1556 (N_1556,N_1147,N_898);
and U1557 (N_1557,N_616,N_1159);
or U1558 (N_1558,N_1183,N_1029);
nand U1559 (N_1559,N_961,N_717);
and U1560 (N_1560,N_985,N_749);
or U1561 (N_1561,N_669,N_1122);
or U1562 (N_1562,N_964,N_948);
or U1563 (N_1563,N_696,N_1034);
nand U1564 (N_1564,N_1102,N_902);
nor U1565 (N_1565,N_1100,N_622);
nor U1566 (N_1566,N_833,N_793);
nand U1567 (N_1567,N_785,N_915);
or U1568 (N_1568,N_724,N_1111);
nor U1569 (N_1569,N_617,N_1116);
nor U1570 (N_1570,N_1072,N_1191);
xnor U1571 (N_1571,N_1179,N_705);
and U1572 (N_1572,N_974,N_1074);
xnor U1573 (N_1573,N_900,N_686);
nand U1574 (N_1574,N_1060,N_1029);
and U1575 (N_1575,N_1112,N_812);
nand U1576 (N_1576,N_1180,N_820);
and U1577 (N_1577,N_1077,N_1117);
nand U1578 (N_1578,N_830,N_851);
and U1579 (N_1579,N_623,N_811);
nand U1580 (N_1580,N_1069,N_837);
nand U1581 (N_1581,N_641,N_886);
or U1582 (N_1582,N_1185,N_788);
and U1583 (N_1583,N_1192,N_1108);
xnor U1584 (N_1584,N_830,N_665);
or U1585 (N_1585,N_936,N_930);
and U1586 (N_1586,N_885,N_705);
or U1587 (N_1587,N_845,N_812);
and U1588 (N_1588,N_707,N_807);
nor U1589 (N_1589,N_1160,N_1180);
or U1590 (N_1590,N_646,N_663);
nand U1591 (N_1591,N_873,N_1125);
or U1592 (N_1592,N_1187,N_964);
nand U1593 (N_1593,N_791,N_923);
or U1594 (N_1594,N_831,N_1127);
or U1595 (N_1595,N_836,N_984);
and U1596 (N_1596,N_663,N_944);
or U1597 (N_1597,N_1050,N_1091);
nor U1598 (N_1598,N_1058,N_643);
nor U1599 (N_1599,N_923,N_1061);
or U1600 (N_1600,N_900,N_709);
or U1601 (N_1601,N_734,N_1094);
nand U1602 (N_1602,N_1122,N_662);
nand U1603 (N_1603,N_690,N_821);
nand U1604 (N_1604,N_879,N_733);
nor U1605 (N_1605,N_916,N_940);
nor U1606 (N_1606,N_642,N_713);
and U1607 (N_1607,N_1192,N_1010);
nor U1608 (N_1608,N_1185,N_1159);
or U1609 (N_1609,N_986,N_874);
nor U1610 (N_1610,N_919,N_1076);
and U1611 (N_1611,N_666,N_1170);
and U1612 (N_1612,N_1090,N_612);
nor U1613 (N_1613,N_683,N_962);
or U1614 (N_1614,N_1198,N_806);
nand U1615 (N_1615,N_924,N_666);
nand U1616 (N_1616,N_1153,N_1130);
nand U1617 (N_1617,N_959,N_932);
and U1618 (N_1618,N_618,N_1044);
or U1619 (N_1619,N_860,N_1005);
or U1620 (N_1620,N_795,N_915);
and U1621 (N_1621,N_880,N_915);
nor U1622 (N_1622,N_1181,N_1073);
xnor U1623 (N_1623,N_1010,N_1173);
and U1624 (N_1624,N_910,N_698);
nand U1625 (N_1625,N_1141,N_987);
and U1626 (N_1626,N_757,N_992);
and U1627 (N_1627,N_975,N_1024);
nand U1628 (N_1628,N_1176,N_708);
nor U1629 (N_1629,N_744,N_1098);
or U1630 (N_1630,N_1043,N_615);
or U1631 (N_1631,N_1071,N_958);
nand U1632 (N_1632,N_850,N_1070);
nor U1633 (N_1633,N_952,N_711);
or U1634 (N_1634,N_1172,N_744);
nand U1635 (N_1635,N_631,N_922);
nand U1636 (N_1636,N_1125,N_1137);
nor U1637 (N_1637,N_759,N_750);
or U1638 (N_1638,N_958,N_999);
nand U1639 (N_1639,N_935,N_641);
and U1640 (N_1640,N_1126,N_855);
and U1641 (N_1641,N_658,N_1179);
nor U1642 (N_1642,N_1190,N_989);
and U1643 (N_1643,N_740,N_1060);
and U1644 (N_1644,N_1117,N_1188);
and U1645 (N_1645,N_854,N_689);
nand U1646 (N_1646,N_1186,N_674);
nor U1647 (N_1647,N_818,N_910);
nand U1648 (N_1648,N_848,N_898);
nand U1649 (N_1649,N_1010,N_788);
nor U1650 (N_1650,N_773,N_1172);
or U1651 (N_1651,N_963,N_947);
nor U1652 (N_1652,N_1177,N_627);
or U1653 (N_1653,N_1047,N_1033);
and U1654 (N_1654,N_907,N_1050);
nor U1655 (N_1655,N_739,N_999);
and U1656 (N_1656,N_867,N_982);
nor U1657 (N_1657,N_822,N_820);
and U1658 (N_1658,N_701,N_1150);
nor U1659 (N_1659,N_898,N_747);
nor U1660 (N_1660,N_781,N_887);
nand U1661 (N_1661,N_1189,N_783);
or U1662 (N_1662,N_1065,N_747);
and U1663 (N_1663,N_752,N_879);
and U1664 (N_1664,N_683,N_829);
nor U1665 (N_1665,N_982,N_727);
and U1666 (N_1666,N_1136,N_1129);
nor U1667 (N_1667,N_739,N_606);
and U1668 (N_1668,N_632,N_1141);
and U1669 (N_1669,N_1189,N_664);
nand U1670 (N_1670,N_934,N_953);
nor U1671 (N_1671,N_793,N_1043);
xor U1672 (N_1672,N_953,N_827);
nor U1673 (N_1673,N_785,N_1030);
nor U1674 (N_1674,N_831,N_961);
nor U1675 (N_1675,N_601,N_698);
nand U1676 (N_1676,N_753,N_1097);
and U1677 (N_1677,N_1038,N_746);
or U1678 (N_1678,N_772,N_605);
nor U1679 (N_1679,N_930,N_692);
and U1680 (N_1680,N_958,N_785);
or U1681 (N_1681,N_995,N_772);
and U1682 (N_1682,N_666,N_1065);
nand U1683 (N_1683,N_1183,N_760);
nand U1684 (N_1684,N_1082,N_924);
nand U1685 (N_1685,N_893,N_698);
nor U1686 (N_1686,N_743,N_631);
or U1687 (N_1687,N_789,N_878);
nor U1688 (N_1688,N_1169,N_650);
nor U1689 (N_1689,N_1178,N_678);
nand U1690 (N_1690,N_794,N_617);
or U1691 (N_1691,N_635,N_992);
and U1692 (N_1692,N_1122,N_696);
nand U1693 (N_1693,N_1173,N_847);
or U1694 (N_1694,N_922,N_1129);
nor U1695 (N_1695,N_1078,N_1131);
nor U1696 (N_1696,N_669,N_887);
nand U1697 (N_1697,N_947,N_625);
or U1698 (N_1698,N_699,N_799);
nand U1699 (N_1699,N_1014,N_615);
xnor U1700 (N_1700,N_1123,N_766);
or U1701 (N_1701,N_894,N_1153);
nand U1702 (N_1702,N_1133,N_922);
nor U1703 (N_1703,N_802,N_754);
or U1704 (N_1704,N_716,N_1013);
and U1705 (N_1705,N_766,N_881);
or U1706 (N_1706,N_1146,N_867);
and U1707 (N_1707,N_905,N_785);
nand U1708 (N_1708,N_934,N_1043);
or U1709 (N_1709,N_666,N_788);
and U1710 (N_1710,N_1089,N_717);
xor U1711 (N_1711,N_956,N_1141);
and U1712 (N_1712,N_845,N_1176);
and U1713 (N_1713,N_916,N_866);
xnor U1714 (N_1714,N_682,N_1040);
nand U1715 (N_1715,N_1097,N_995);
nand U1716 (N_1716,N_1104,N_874);
and U1717 (N_1717,N_665,N_1114);
or U1718 (N_1718,N_998,N_1171);
or U1719 (N_1719,N_798,N_728);
nor U1720 (N_1720,N_1164,N_1149);
and U1721 (N_1721,N_834,N_772);
and U1722 (N_1722,N_721,N_624);
or U1723 (N_1723,N_982,N_623);
nand U1724 (N_1724,N_603,N_983);
nor U1725 (N_1725,N_726,N_1008);
or U1726 (N_1726,N_1146,N_655);
nor U1727 (N_1727,N_803,N_1173);
nor U1728 (N_1728,N_794,N_1028);
nand U1729 (N_1729,N_732,N_615);
nor U1730 (N_1730,N_1004,N_794);
and U1731 (N_1731,N_1011,N_707);
and U1732 (N_1732,N_790,N_668);
and U1733 (N_1733,N_1104,N_1198);
nand U1734 (N_1734,N_979,N_853);
or U1735 (N_1735,N_1064,N_852);
nor U1736 (N_1736,N_1063,N_691);
and U1737 (N_1737,N_661,N_986);
or U1738 (N_1738,N_993,N_1174);
nor U1739 (N_1739,N_1063,N_856);
and U1740 (N_1740,N_694,N_847);
nor U1741 (N_1741,N_1106,N_754);
nor U1742 (N_1742,N_766,N_708);
or U1743 (N_1743,N_731,N_1030);
nand U1744 (N_1744,N_768,N_903);
nor U1745 (N_1745,N_1078,N_1003);
or U1746 (N_1746,N_634,N_967);
nor U1747 (N_1747,N_799,N_652);
xnor U1748 (N_1748,N_899,N_778);
or U1749 (N_1749,N_749,N_631);
nand U1750 (N_1750,N_642,N_1141);
nor U1751 (N_1751,N_979,N_700);
nor U1752 (N_1752,N_881,N_692);
nor U1753 (N_1753,N_936,N_712);
or U1754 (N_1754,N_779,N_985);
or U1755 (N_1755,N_786,N_1091);
or U1756 (N_1756,N_994,N_645);
nor U1757 (N_1757,N_675,N_710);
and U1758 (N_1758,N_911,N_917);
nor U1759 (N_1759,N_1021,N_644);
and U1760 (N_1760,N_719,N_903);
or U1761 (N_1761,N_654,N_1000);
nor U1762 (N_1762,N_1109,N_1045);
nand U1763 (N_1763,N_601,N_671);
nor U1764 (N_1764,N_955,N_1045);
and U1765 (N_1765,N_1081,N_689);
nor U1766 (N_1766,N_1111,N_1048);
nand U1767 (N_1767,N_1012,N_848);
nor U1768 (N_1768,N_858,N_1001);
or U1769 (N_1769,N_1002,N_684);
or U1770 (N_1770,N_1021,N_816);
or U1771 (N_1771,N_1058,N_965);
and U1772 (N_1772,N_910,N_855);
nand U1773 (N_1773,N_1034,N_1081);
nand U1774 (N_1774,N_1119,N_706);
nand U1775 (N_1775,N_745,N_772);
nand U1776 (N_1776,N_1186,N_1106);
and U1777 (N_1777,N_1055,N_622);
and U1778 (N_1778,N_1154,N_747);
and U1779 (N_1779,N_641,N_1087);
and U1780 (N_1780,N_975,N_819);
nand U1781 (N_1781,N_808,N_1023);
and U1782 (N_1782,N_1037,N_1087);
nor U1783 (N_1783,N_850,N_1102);
nand U1784 (N_1784,N_1036,N_1144);
or U1785 (N_1785,N_946,N_708);
or U1786 (N_1786,N_938,N_891);
nand U1787 (N_1787,N_962,N_758);
xor U1788 (N_1788,N_1025,N_812);
nor U1789 (N_1789,N_1004,N_828);
nand U1790 (N_1790,N_686,N_1099);
nand U1791 (N_1791,N_611,N_644);
nor U1792 (N_1792,N_952,N_981);
nand U1793 (N_1793,N_722,N_987);
nor U1794 (N_1794,N_787,N_966);
or U1795 (N_1795,N_971,N_1185);
nor U1796 (N_1796,N_1029,N_786);
nor U1797 (N_1797,N_768,N_1142);
or U1798 (N_1798,N_1090,N_638);
or U1799 (N_1799,N_837,N_799);
nand U1800 (N_1800,N_1477,N_1269);
xor U1801 (N_1801,N_1739,N_1323);
and U1802 (N_1802,N_1290,N_1251);
and U1803 (N_1803,N_1666,N_1671);
and U1804 (N_1804,N_1518,N_1472);
or U1805 (N_1805,N_1724,N_1276);
and U1806 (N_1806,N_1220,N_1210);
or U1807 (N_1807,N_1598,N_1591);
or U1808 (N_1808,N_1463,N_1437);
or U1809 (N_1809,N_1785,N_1252);
nand U1810 (N_1810,N_1315,N_1609);
or U1811 (N_1811,N_1539,N_1482);
xnor U1812 (N_1812,N_1688,N_1732);
nor U1813 (N_1813,N_1756,N_1730);
or U1814 (N_1814,N_1771,N_1744);
nor U1815 (N_1815,N_1774,N_1411);
and U1816 (N_1816,N_1381,N_1408);
or U1817 (N_1817,N_1259,N_1233);
or U1818 (N_1818,N_1726,N_1209);
nor U1819 (N_1819,N_1583,N_1594);
nand U1820 (N_1820,N_1500,N_1655);
nand U1821 (N_1821,N_1288,N_1424);
and U1822 (N_1822,N_1794,N_1721);
nand U1823 (N_1823,N_1585,N_1568);
nand U1824 (N_1824,N_1229,N_1257);
nand U1825 (N_1825,N_1275,N_1677);
or U1826 (N_1826,N_1641,N_1703);
or U1827 (N_1827,N_1738,N_1490);
and U1828 (N_1828,N_1452,N_1279);
or U1829 (N_1829,N_1234,N_1380);
nand U1830 (N_1830,N_1433,N_1772);
and U1831 (N_1831,N_1560,N_1619);
nand U1832 (N_1832,N_1610,N_1292);
or U1833 (N_1833,N_1617,N_1332);
nor U1834 (N_1834,N_1728,N_1551);
or U1835 (N_1835,N_1366,N_1543);
and U1836 (N_1836,N_1317,N_1314);
and U1837 (N_1837,N_1376,N_1662);
nand U1838 (N_1838,N_1696,N_1574);
nor U1839 (N_1839,N_1699,N_1328);
and U1840 (N_1840,N_1669,N_1658);
and U1841 (N_1841,N_1403,N_1531);
nor U1842 (N_1842,N_1468,N_1566);
nand U1843 (N_1843,N_1272,N_1430);
nand U1844 (N_1844,N_1534,N_1448);
nand U1845 (N_1845,N_1212,N_1420);
or U1846 (N_1846,N_1532,N_1710);
or U1847 (N_1847,N_1407,N_1797);
nor U1848 (N_1848,N_1608,N_1456);
and U1849 (N_1849,N_1321,N_1489);
or U1850 (N_1850,N_1384,N_1522);
or U1851 (N_1851,N_1659,N_1512);
nand U1852 (N_1852,N_1506,N_1559);
nand U1853 (N_1853,N_1254,N_1246);
nor U1854 (N_1854,N_1215,N_1258);
nand U1855 (N_1855,N_1673,N_1533);
and U1856 (N_1856,N_1438,N_1554);
nor U1857 (N_1857,N_1618,N_1752);
nand U1858 (N_1858,N_1647,N_1719);
nor U1859 (N_1859,N_1417,N_1218);
and U1860 (N_1860,N_1553,N_1747);
nand U1861 (N_1861,N_1341,N_1562);
or U1862 (N_1862,N_1379,N_1498);
and U1863 (N_1863,N_1602,N_1324);
nand U1864 (N_1864,N_1718,N_1701);
xor U1865 (N_1865,N_1410,N_1221);
nand U1866 (N_1866,N_1395,N_1651);
nand U1867 (N_1867,N_1383,N_1621);
nand U1868 (N_1868,N_1611,N_1636);
or U1869 (N_1869,N_1646,N_1670);
or U1870 (N_1870,N_1318,N_1309);
nand U1871 (N_1871,N_1654,N_1573);
or U1872 (N_1872,N_1765,N_1312);
and U1873 (N_1873,N_1557,N_1280);
nor U1874 (N_1874,N_1639,N_1453);
nor U1875 (N_1875,N_1331,N_1502);
and U1876 (N_1876,N_1465,N_1592);
xnor U1877 (N_1877,N_1773,N_1740);
and U1878 (N_1878,N_1492,N_1525);
and U1879 (N_1879,N_1255,N_1224);
nor U1880 (N_1880,N_1588,N_1386);
and U1881 (N_1881,N_1340,N_1289);
nor U1882 (N_1882,N_1799,N_1418);
or U1883 (N_1883,N_1577,N_1552);
nor U1884 (N_1884,N_1695,N_1550);
nor U1885 (N_1885,N_1788,N_1513);
or U1886 (N_1886,N_1741,N_1353);
nor U1887 (N_1887,N_1336,N_1729);
and U1888 (N_1888,N_1444,N_1682);
and U1889 (N_1889,N_1271,N_1450);
and U1890 (N_1890,N_1230,N_1347);
xor U1891 (N_1891,N_1627,N_1447);
nor U1892 (N_1892,N_1569,N_1389);
or U1893 (N_1893,N_1296,N_1645);
or U1894 (N_1894,N_1714,N_1293);
or U1895 (N_1895,N_1795,N_1443);
or U1896 (N_1896,N_1624,N_1634);
nor U1897 (N_1897,N_1571,N_1731);
nand U1898 (N_1898,N_1213,N_1364);
and U1899 (N_1899,N_1301,N_1432);
and U1900 (N_1900,N_1563,N_1733);
and U1901 (N_1901,N_1346,N_1576);
or U1902 (N_1902,N_1414,N_1235);
nand U1903 (N_1903,N_1322,N_1371);
xor U1904 (N_1904,N_1520,N_1690);
and U1905 (N_1905,N_1263,N_1613);
or U1906 (N_1906,N_1349,N_1205);
and U1907 (N_1907,N_1668,N_1387);
nand U1908 (N_1908,N_1762,N_1278);
nor U1909 (N_1909,N_1475,N_1697);
nand U1910 (N_1910,N_1337,N_1544);
and U1911 (N_1911,N_1684,N_1261);
and U1912 (N_1912,N_1285,N_1524);
and U1913 (N_1913,N_1567,N_1372);
or U1914 (N_1914,N_1495,N_1404);
nor U1915 (N_1915,N_1206,N_1491);
and U1916 (N_1916,N_1635,N_1273);
or U1917 (N_1917,N_1504,N_1743);
or U1918 (N_1918,N_1339,N_1485);
and U1919 (N_1919,N_1343,N_1734);
or U1920 (N_1920,N_1359,N_1793);
or U1921 (N_1921,N_1757,N_1558);
nor U1922 (N_1922,N_1750,N_1597);
or U1923 (N_1923,N_1222,N_1535);
nand U1924 (N_1924,N_1446,N_1326);
nor U1925 (N_1925,N_1219,N_1590);
nor U1926 (N_1926,N_1754,N_1413);
and U1927 (N_1927,N_1226,N_1792);
nand U1928 (N_1928,N_1615,N_1628);
nor U1929 (N_1929,N_1656,N_1589);
or U1930 (N_1930,N_1497,N_1297);
nand U1931 (N_1931,N_1427,N_1707);
and U1932 (N_1932,N_1236,N_1440);
nor U1933 (N_1933,N_1674,N_1382);
or U1934 (N_1934,N_1565,N_1333);
or U1935 (N_1935,N_1717,N_1545);
xor U1936 (N_1936,N_1361,N_1228);
nand U1937 (N_1937,N_1421,N_1607);
xnor U1938 (N_1938,N_1460,N_1758);
nand U1939 (N_1939,N_1434,N_1702);
nor U1940 (N_1940,N_1330,N_1334);
nor U1941 (N_1941,N_1516,N_1439);
and U1942 (N_1942,N_1377,N_1649);
or U1943 (N_1943,N_1536,N_1687);
or U1944 (N_1944,N_1678,N_1412);
and U1945 (N_1945,N_1601,N_1722);
xor U1946 (N_1946,N_1614,N_1307);
nor U1947 (N_1947,N_1537,N_1392);
nand U1948 (N_1948,N_1716,N_1685);
nor U1949 (N_1949,N_1705,N_1767);
and U1950 (N_1950,N_1352,N_1638);
nand U1951 (N_1951,N_1523,N_1399);
nor U1952 (N_1952,N_1599,N_1789);
and U1953 (N_1953,N_1470,N_1201);
nor U1954 (N_1954,N_1737,N_1342);
or U1955 (N_1955,N_1620,N_1373);
xor U1956 (N_1956,N_1640,N_1580);
nand U1957 (N_1957,N_1511,N_1249);
and U1958 (N_1958,N_1625,N_1239);
nand U1959 (N_1959,N_1692,N_1759);
nand U1960 (N_1960,N_1481,N_1686);
nor U1961 (N_1961,N_1242,N_1572);
nand U1962 (N_1962,N_1496,N_1355);
and U1963 (N_1963,N_1517,N_1704);
or U1964 (N_1964,N_1436,N_1268);
or U1965 (N_1965,N_1394,N_1760);
nand U1966 (N_1966,N_1422,N_1238);
and U1967 (N_1967,N_1781,N_1476);
nand U1968 (N_1968,N_1711,N_1473);
nor U1969 (N_1969,N_1391,N_1419);
nand U1970 (N_1970,N_1329,N_1316);
nor U1971 (N_1971,N_1350,N_1751);
nand U1972 (N_1972,N_1365,N_1600);
and U1973 (N_1973,N_1295,N_1466);
nand U1974 (N_1974,N_1214,N_1623);
nand U1975 (N_1975,N_1484,N_1510);
and U1976 (N_1976,N_1796,N_1631);
and U1977 (N_1977,N_1521,N_1786);
or U1978 (N_1978,N_1667,N_1713);
nand U1979 (N_1979,N_1277,N_1661);
or U1980 (N_1980,N_1266,N_1715);
nand U1981 (N_1981,N_1400,N_1304);
nand U1982 (N_1982,N_1325,N_1388);
and U1983 (N_1983,N_1435,N_1415);
nor U1984 (N_1984,N_1596,N_1459);
or U1985 (N_1985,N_1745,N_1256);
nor U1986 (N_1986,N_1274,N_1425);
or U1987 (N_1987,N_1327,N_1449);
nand U1988 (N_1988,N_1787,N_1308);
nor U1989 (N_1989,N_1547,N_1368);
nand U1990 (N_1990,N_1775,N_1556);
and U1991 (N_1991,N_1549,N_1783);
nand U1992 (N_1992,N_1454,N_1604);
and U1993 (N_1993,N_1612,N_1691);
nor U1994 (N_1994,N_1310,N_1727);
nor U1995 (N_1995,N_1445,N_1633);
nand U1996 (N_1996,N_1672,N_1225);
nand U1997 (N_1997,N_1519,N_1429);
nand U1998 (N_1998,N_1493,N_1302);
nand U1999 (N_1999,N_1363,N_1581);
and U2000 (N_2000,N_1299,N_1768);
nor U2001 (N_2001,N_1483,N_1709);
and U2002 (N_2002,N_1527,N_1338);
nand U2003 (N_2003,N_1385,N_1282);
or U2004 (N_2004,N_1622,N_1777);
nand U2005 (N_2005,N_1294,N_1305);
and U2006 (N_2006,N_1241,N_1480);
or U2007 (N_2007,N_1776,N_1753);
or U2008 (N_2008,N_1708,N_1455);
or U2009 (N_2009,N_1319,N_1243);
or U2010 (N_2010,N_1791,N_1766);
or U2011 (N_2011,N_1231,N_1575);
nor U2012 (N_2012,N_1593,N_1370);
or U2013 (N_2013,N_1528,N_1360);
or U2014 (N_2014,N_1644,N_1712);
nand U2015 (N_2015,N_1397,N_1451);
and U2016 (N_2016,N_1458,N_1579);
nor U2017 (N_2017,N_1461,N_1784);
and U2018 (N_2018,N_1770,N_1570);
nand U2019 (N_2019,N_1398,N_1664);
nor U2020 (N_2020,N_1507,N_1216);
or U2021 (N_2021,N_1508,N_1283);
nor U2022 (N_2022,N_1723,N_1603);
nand U2023 (N_2023,N_1313,N_1390);
nand U2024 (N_2024,N_1749,N_1291);
nor U2025 (N_2025,N_1260,N_1501);
nor U2026 (N_2026,N_1616,N_1605);
nor U2027 (N_2027,N_1681,N_1375);
nand U2028 (N_2028,N_1393,N_1642);
nand U2029 (N_2029,N_1200,N_1555);
or U2030 (N_2030,N_1736,N_1720);
nand U2031 (N_2031,N_1763,N_1345);
nor U2032 (N_2032,N_1428,N_1287);
and U2033 (N_2033,N_1650,N_1441);
xnor U2034 (N_2034,N_1300,N_1211);
nand U2035 (N_2035,N_1486,N_1725);
nor U2036 (N_2036,N_1262,N_1595);
and U2037 (N_2037,N_1790,N_1746);
and U2038 (N_2038,N_1402,N_1748);
xor U2039 (N_2039,N_1648,N_1735);
or U2040 (N_2040,N_1396,N_1742);
or U2041 (N_2041,N_1335,N_1679);
and U2042 (N_2042,N_1629,N_1227);
nand U2043 (N_2043,N_1653,N_1247);
or U2044 (N_2044,N_1764,N_1409);
nor U2045 (N_2045,N_1270,N_1494);
nand U2046 (N_2046,N_1462,N_1529);
and U2047 (N_2047,N_1405,N_1675);
or U2048 (N_2048,N_1362,N_1578);
or U2049 (N_2049,N_1546,N_1564);
and U2050 (N_2050,N_1487,N_1660);
or U2051 (N_2051,N_1298,N_1626);
nor U2052 (N_2052,N_1540,N_1245);
nand U2053 (N_2053,N_1354,N_1548);
nand U2054 (N_2054,N_1689,N_1311);
nand U2055 (N_2055,N_1207,N_1464);
nor U2056 (N_2056,N_1587,N_1478);
nand U2057 (N_2057,N_1369,N_1778);
nand U2058 (N_2058,N_1457,N_1515);
and U2059 (N_2059,N_1281,N_1683);
or U2060 (N_2060,N_1526,N_1374);
and U2061 (N_2061,N_1643,N_1351);
or U2062 (N_2062,N_1657,N_1503);
or U2063 (N_2063,N_1284,N_1240);
nand U2064 (N_2064,N_1442,N_1630);
nand U2065 (N_2065,N_1203,N_1250);
or U2066 (N_2066,N_1509,N_1505);
or U2067 (N_2067,N_1306,N_1244);
or U2068 (N_2068,N_1542,N_1204);
nor U2069 (N_2069,N_1780,N_1378);
and U2070 (N_2070,N_1652,N_1755);
and U2071 (N_2071,N_1248,N_1264);
and U2072 (N_2072,N_1663,N_1779);
and U2073 (N_2073,N_1700,N_1584);
or U2074 (N_2074,N_1356,N_1426);
and U2075 (N_2075,N_1530,N_1303);
or U2076 (N_2076,N_1232,N_1706);
and U2077 (N_2077,N_1586,N_1479);
nand U2078 (N_2078,N_1431,N_1223);
nand U2079 (N_2079,N_1693,N_1761);
and U2080 (N_2080,N_1488,N_1320);
and U2081 (N_2081,N_1208,N_1782);
and U2082 (N_2082,N_1676,N_1237);
and U2083 (N_2083,N_1344,N_1267);
or U2084 (N_2084,N_1423,N_1582);
nand U2085 (N_2085,N_1253,N_1798);
nor U2086 (N_2086,N_1694,N_1367);
nand U2087 (N_2087,N_1499,N_1286);
or U2088 (N_2088,N_1406,N_1632);
or U2089 (N_2089,N_1637,N_1561);
nand U2090 (N_2090,N_1538,N_1265);
and U2091 (N_2091,N_1202,N_1217);
nand U2092 (N_2092,N_1471,N_1474);
and U2093 (N_2093,N_1698,N_1401);
or U2094 (N_2094,N_1357,N_1348);
nand U2095 (N_2095,N_1680,N_1769);
nand U2096 (N_2096,N_1514,N_1416);
or U2097 (N_2097,N_1469,N_1358);
and U2098 (N_2098,N_1665,N_1467);
nand U2099 (N_2099,N_1606,N_1541);
nor U2100 (N_2100,N_1410,N_1622);
and U2101 (N_2101,N_1791,N_1255);
and U2102 (N_2102,N_1331,N_1792);
and U2103 (N_2103,N_1520,N_1601);
nand U2104 (N_2104,N_1373,N_1551);
xor U2105 (N_2105,N_1653,N_1422);
and U2106 (N_2106,N_1458,N_1287);
nor U2107 (N_2107,N_1738,N_1235);
or U2108 (N_2108,N_1554,N_1380);
and U2109 (N_2109,N_1411,N_1680);
and U2110 (N_2110,N_1296,N_1386);
nor U2111 (N_2111,N_1390,N_1751);
xnor U2112 (N_2112,N_1432,N_1527);
nor U2113 (N_2113,N_1368,N_1566);
nor U2114 (N_2114,N_1779,N_1719);
and U2115 (N_2115,N_1433,N_1728);
nor U2116 (N_2116,N_1765,N_1428);
nor U2117 (N_2117,N_1212,N_1513);
and U2118 (N_2118,N_1599,N_1515);
nor U2119 (N_2119,N_1238,N_1564);
nor U2120 (N_2120,N_1658,N_1420);
nand U2121 (N_2121,N_1616,N_1250);
or U2122 (N_2122,N_1684,N_1747);
and U2123 (N_2123,N_1571,N_1596);
nand U2124 (N_2124,N_1563,N_1610);
and U2125 (N_2125,N_1615,N_1247);
nand U2126 (N_2126,N_1233,N_1618);
or U2127 (N_2127,N_1304,N_1728);
nor U2128 (N_2128,N_1560,N_1521);
nand U2129 (N_2129,N_1418,N_1300);
nand U2130 (N_2130,N_1299,N_1245);
nor U2131 (N_2131,N_1519,N_1714);
nor U2132 (N_2132,N_1649,N_1601);
nor U2133 (N_2133,N_1439,N_1238);
or U2134 (N_2134,N_1260,N_1405);
xor U2135 (N_2135,N_1494,N_1555);
or U2136 (N_2136,N_1266,N_1319);
nand U2137 (N_2137,N_1725,N_1302);
and U2138 (N_2138,N_1641,N_1542);
or U2139 (N_2139,N_1215,N_1788);
nand U2140 (N_2140,N_1317,N_1771);
nand U2141 (N_2141,N_1306,N_1243);
or U2142 (N_2142,N_1711,N_1692);
or U2143 (N_2143,N_1299,N_1229);
nor U2144 (N_2144,N_1568,N_1546);
nand U2145 (N_2145,N_1744,N_1385);
and U2146 (N_2146,N_1267,N_1305);
and U2147 (N_2147,N_1454,N_1723);
nand U2148 (N_2148,N_1770,N_1683);
nor U2149 (N_2149,N_1577,N_1731);
nand U2150 (N_2150,N_1407,N_1241);
nor U2151 (N_2151,N_1687,N_1703);
or U2152 (N_2152,N_1572,N_1210);
xor U2153 (N_2153,N_1705,N_1492);
nand U2154 (N_2154,N_1423,N_1602);
nor U2155 (N_2155,N_1536,N_1796);
and U2156 (N_2156,N_1654,N_1570);
or U2157 (N_2157,N_1224,N_1465);
nor U2158 (N_2158,N_1734,N_1465);
or U2159 (N_2159,N_1635,N_1225);
nor U2160 (N_2160,N_1773,N_1260);
or U2161 (N_2161,N_1525,N_1796);
and U2162 (N_2162,N_1573,N_1264);
nand U2163 (N_2163,N_1763,N_1695);
nor U2164 (N_2164,N_1544,N_1799);
nor U2165 (N_2165,N_1638,N_1576);
nor U2166 (N_2166,N_1219,N_1511);
or U2167 (N_2167,N_1206,N_1397);
nand U2168 (N_2168,N_1447,N_1774);
nand U2169 (N_2169,N_1260,N_1558);
nand U2170 (N_2170,N_1626,N_1311);
nor U2171 (N_2171,N_1527,N_1315);
nand U2172 (N_2172,N_1316,N_1627);
xor U2173 (N_2173,N_1523,N_1316);
and U2174 (N_2174,N_1608,N_1407);
nor U2175 (N_2175,N_1476,N_1783);
nand U2176 (N_2176,N_1387,N_1679);
nor U2177 (N_2177,N_1531,N_1237);
nand U2178 (N_2178,N_1281,N_1660);
and U2179 (N_2179,N_1748,N_1409);
or U2180 (N_2180,N_1735,N_1379);
nor U2181 (N_2181,N_1533,N_1726);
nand U2182 (N_2182,N_1691,N_1572);
and U2183 (N_2183,N_1793,N_1520);
nor U2184 (N_2184,N_1706,N_1627);
and U2185 (N_2185,N_1641,N_1312);
and U2186 (N_2186,N_1410,N_1461);
nand U2187 (N_2187,N_1352,N_1762);
nand U2188 (N_2188,N_1259,N_1484);
or U2189 (N_2189,N_1754,N_1569);
and U2190 (N_2190,N_1345,N_1509);
and U2191 (N_2191,N_1643,N_1438);
nor U2192 (N_2192,N_1201,N_1677);
or U2193 (N_2193,N_1275,N_1326);
nand U2194 (N_2194,N_1785,N_1718);
or U2195 (N_2195,N_1739,N_1509);
nor U2196 (N_2196,N_1614,N_1707);
xor U2197 (N_2197,N_1370,N_1358);
and U2198 (N_2198,N_1481,N_1530);
or U2199 (N_2199,N_1411,N_1264);
nand U2200 (N_2200,N_1293,N_1596);
and U2201 (N_2201,N_1224,N_1504);
and U2202 (N_2202,N_1712,N_1708);
nand U2203 (N_2203,N_1611,N_1495);
nor U2204 (N_2204,N_1545,N_1763);
nor U2205 (N_2205,N_1302,N_1209);
nor U2206 (N_2206,N_1690,N_1755);
and U2207 (N_2207,N_1730,N_1388);
nand U2208 (N_2208,N_1629,N_1285);
or U2209 (N_2209,N_1275,N_1274);
and U2210 (N_2210,N_1285,N_1670);
nor U2211 (N_2211,N_1727,N_1304);
and U2212 (N_2212,N_1390,N_1524);
and U2213 (N_2213,N_1289,N_1474);
or U2214 (N_2214,N_1643,N_1357);
nor U2215 (N_2215,N_1454,N_1539);
and U2216 (N_2216,N_1776,N_1718);
nor U2217 (N_2217,N_1674,N_1712);
nand U2218 (N_2218,N_1632,N_1352);
nand U2219 (N_2219,N_1713,N_1535);
or U2220 (N_2220,N_1330,N_1528);
or U2221 (N_2221,N_1403,N_1430);
nor U2222 (N_2222,N_1343,N_1632);
nor U2223 (N_2223,N_1241,N_1369);
nand U2224 (N_2224,N_1423,N_1223);
and U2225 (N_2225,N_1206,N_1344);
and U2226 (N_2226,N_1769,N_1214);
and U2227 (N_2227,N_1217,N_1609);
nor U2228 (N_2228,N_1453,N_1389);
nor U2229 (N_2229,N_1789,N_1452);
nor U2230 (N_2230,N_1613,N_1627);
or U2231 (N_2231,N_1245,N_1711);
or U2232 (N_2232,N_1242,N_1241);
nor U2233 (N_2233,N_1705,N_1233);
nand U2234 (N_2234,N_1761,N_1239);
or U2235 (N_2235,N_1597,N_1331);
nand U2236 (N_2236,N_1335,N_1439);
nor U2237 (N_2237,N_1340,N_1724);
nand U2238 (N_2238,N_1540,N_1487);
nand U2239 (N_2239,N_1592,N_1492);
and U2240 (N_2240,N_1513,N_1372);
nor U2241 (N_2241,N_1705,N_1235);
nor U2242 (N_2242,N_1225,N_1690);
or U2243 (N_2243,N_1402,N_1221);
and U2244 (N_2244,N_1524,N_1622);
and U2245 (N_2245,N_1699,N_1633);
and U2246 (N_2246,N_1222,N_1260);
nand U2247 (N_2247,N_1612,N_1516);
nand U2248 (N_2248,N_1661,N_1332);
nand U2249 (N_2249,N_1754,N_1493);
nand U2250 (N_2250,N_1344,N_1443);
nand U2251 (N_2251,N_1688,N_1793);
or U2252 (N_2252,N_1272,N_1568);
or U2253 (N_2253,N_1317,N_1535);
or U2254 (N_2254,N_1759,N_1776);
nor U2255 (N_2255,N_1509,N_1475);
or U2256 (N_2256,N_1766,N_1704);
and U2257 (N_2257,N_1605,N_1698);
or U2258 (N_2258,N_1236,N_1489);
and U2259 (N_2259,N_1336,N_1794);
or U2260 (N_2260,N_1627,N_1652);
or U2261 (N_2261,N_1308,N_1654);
or U2262 (N_2262,N_1425,N_1351);
and U2263 (N_2263,N_1327,N_1605);
and U2264 (N_2264,N_1483,N_1304);
nand U2265 (N_2265,N_1688,N_1316);
or U2266 (N_2266,N_1340,N_1652);
and U2267 (N_2267,N_1428,N_1397);
and U2268 (N_2268,N_1513,N_1242);
and U2269 (N_2269,N_1464,N_1755);
nor U2270 (N_2270,N_1685,N_1240);
nand U2271 (N_2271,N_1422,N_1333);
or U2272 (N_2272,N_1368,N_1415);
and U2273 (N_2273,N_1446,N_1719);
and U2274 (N_2274,N_1418,N_1296);
or U2275 (N_2275,N_1537,N_1776);
nor U2276 (N_2276,N_1253,N_1297);
or U2277 (N_2277,N_1552,N_1560);
nand U2278 (N_2278,N_1514,N_1788);
or U2279 (N_2279,N_1365,N_1438);
nand U2280 (N_2280,N_1470,N_1306);
or U2281 (N_2281,N_1746,N_1466);
or U2282 (N_2282,N_1371,N_1259);
nand U2283 (N_2283,N_1216,N_1242);
or U2284 (N_2284,N_1451,N_1369);
nor U2285 (N_2285,N_1277,N_1701);
and U2286 (N_2286,N_1600,N_1493);
nor U2287 (N_2287,N_1739,N_1318);
and U2288 (N_2288,N_1223,N_1642);
nor U2289 (N_2289,N_1270,N_1484);
or U2290 (N_2290,N_1519,N_1293);
nand U2291 (N_2291,N_1401,N_1791);
and U2292 (N_2292,N_1536,N_1289);
nor U2293 (N_2293,N_1453,N_1595);
and U2294 (N_2294,N_1758,N_1278);
nor U2295 (N_2295,N_1362,N_1504);
nor U2296 (N_2296,N_1739,N_1676);
and U2297 (N_2297,N_1742,N_1728);
nand U2298 (N_2298,N_1679,N_1626);
nor U2299 (N_2299,N_1324,N_1399);
or U2300 (N_2300,N_1546,N_1764);
and U2301 (N_2301,N_1570,N_1649);
nand U2302 (N_2302,N_1266,N_1293);
nor U2303 (N_2303,N_1305,N_1245);
nor U2304 (N_2304,N_1704,N_1401);
nand U2305 (N_2305,N_1754,N_1255);
nor U2306 (N_2306,N_1413,N_1346);
or U2307 (N_2307,N_1633,N_1433);
xnor U2308 (N_2308,N_1746,N_1398);
nand U2309 (N_2309,N_1655,N_1504);
nand U2310 (N_2310,N_1441,N_1734);
nand U2311 (N_2311,N_1279,N_1640);
nand U2312 (N_2312,N_1645,N_1304);
or U2313 (N_2313,N_1442,N_1497);
nor U2314 (N_2314,N_1460,N_1730);
nor U2315 (N_2315,N_1267,N_1323);
nor U2316 (N_2316,N_1225,N_1639);
nand U2317 (N_2317,N_1501,N_1745);
and U2318 (N_2318,N_1536,N_1780);
or U2319 (N_2319,N_1350,N_1523);
or U2320 (N_2320,N_1624,N_1306);
or U2321 (N_2321,N_1403,N_1433);
or U2322 (N_2322,N_1205,N_1426);
or U2323 (N_2323,N_1526,N_1514);
and U2324 (N_2324,N_1443,N_1254);
and U2325 (N_2325,N_1786,N_1745);
nor U2326 (N_2326,N_1246,N_1637);
nor U2327 (N_2327,N_1404,N_1725);
nor U2328 (N_2328,N_1509,N_1436);
nand U2329 (N_2329,N_1613,N_1644);
nor U2330 (N_2330,N_1403,N_1357);
nand U2331 (N_2331,N_1246,N_1561);
nor U2332 (N_2332,N_1251,N_1318);
xor U2333 (N_2333,N_1749,N_1325);
or U2334 (N_2334,N_1206,N_1203);
or U2335 (N_2335,N_1673,N_1582);
and U2336 (N_2336,N_1724,N_1602);
and U2337 (N_2337,N_1318,N_1424);
nand U2338 (N_2338,N_1722,N_1572);
nand U2339 (N_2339,N_1725,N_1579);
or U2340 (N_2340,N_1618,N_1516);
nor U2341 (N_2341,N_1479,N_1449);
or U2342 (N_2342,N_1726,N_1338);
or U2343 (N_2343,N_1559,N_1755);
nand U2344 (N_2344,N_1504,N_1682);
and U2345 (N_2345,N_1732,N_1774);
nor U2346 (N_2346,N_1403,N_1446);
nor U2347 (N_2347,N_1701,N_1795);
nor U2348 (N_2348,N_1426,N_1667);
and U2349 (N_2349,N_1696,N_1766);
nor U2350 (N_2350,N_1549,N_1428);
and U2351 (N_2351,N_1351,N_1222);
nand U2352 (N_2352,N_1484,N_1611);
and U2353 (N_2353,N_1598,N_1253);
nand U2354 (N_2354,N_1291,N_1579);
nor U2355 (N_2355,N_1774,N_1665);
nand U2356 (N_2356,N_1393,N_1300);
nand U2357 (N_2357,N_1379,N_1266);
nor U2358 (N_2358,N_1626,N_1352);
nand U2359 (N_2359,N_1644,N_1296);
nand U2360 (N_2360,N_1651,N_1593);
and U2361 (N_2361,N_1764,N_1232);
or U2362 (N_2362,N_1600,N_1645);
xor U2363 (N_2363,N_1768,N_1727);
nor U2364 (N_2364,N_1302,N_1625);
and U2365 (N_2365,N_1285,N_1798);
or U2366 (N_2366,N_1464,N_1738);
nand U2367 (N_2367,N_1453,N_1700);
or U2368 (N_2368,N_1754,N_1539);
and U2369 (N_2369,N_1646,N_1534);
and U2370 (N_2370,N_1728,N_1572);
nor U2371 (N_2371,N_1464,N_1576);
and U2372 (N_2372,N_1572,N_1711);
nand U2373 (N_2373,N_1411,N_1623);
nand U2374 (N_2374,N_1648,N_1507);
and U2375 (N_2375,N_1330,N_1763);
and U2376 (N_2376,N_1472,N_1354);
nand U2377 (N_2377,N_1546,N_1716);
or U2378 (N_2378,N_1599,N_1252);
or U2379 (N_2379,N_1588,N_1263);
and U2380 (N_2380,N_1385,N_1419);
nor U2381 (N_2381,N_1587,N_1444);
nand U2382 (N_2382,N_1339,N_1250);
nor U2383 (N_2383,N_1759,N_1435);
or U2384 (N_2384,N_1763,N_1447);
nand U2385 (N_2385,N_1238,N_1693);
nand U2386 (N_2386,N_1448,N_1554);
nand U2387 (N_2387,N_1400,N_1608);
nand U2388 (N_2388,N_1398,N_1495);
and U2389 (N_2389,N_1598,N_1759);
nor U2390 (N_2390,N_1243,N_1501);
or U2391 (N_2391,N_1451,N_1554);
nand U2392 (N_2392,N_1461,N_1498);
xnor U2393 (N_2393,N_1416,N_1635);
nand U2394 (N_2394,N_1233,N_1413);
nand U2395 (N_2395,N_1381,N_1241);
nor U2396 (N_2396,N_1704,N_1620);
nand U2397 (N_2397,N_1675,N_1560);
nor U2398 (N_2398,N_1372,N_1289);
or U2399 (N_2399,N_1713,N_1510);
or U2400 (N_2400,N_2393,N_2323);
and U2401 (N_2401,N_2112,N_1810);
and U2402 (N_2402,N_2169,N_1897);
and U2403 (N_2403,N_2225,N_1952);
or U2404 (N_2404,N_2179,N_2298);
or U2405 (N_2405,N_1903,N_1981);
and U2406 (N_2406,N_2291,N_2153);
or U2407 (N_2407,N_2375,N_2265);
nor U2408 (N_2408,N_2226,N_2261);
nor U2409 (N_2409,N_2259,N_2084);
nand U2410 (N_2410,N_2145,N_2293);
nor U2411 (N_2411,N_2344,N_2369);
or U2412 (N_2412,N_2078,N_2223);
or U2413 (N_2413,N_2330,N_2041);
or U2414 (N_2414,N_2341,N_2386);
and U2415 (N_2415,N_2017,N_1912);
nor U2416 (N_2416,N_2029,N_1996);
and U2417 (N_2417,N_1926,N_2098);
and U2418 (N_2418,N_2103,N_1856);
nand U2419 (N_2419,N_2242,N_2068);
nor U2420 (N_2420,N_2154,N_2165);
or U2421 (N_2421,N_2244,N_1929);
or U2422 (N_2422,N_2326,N_2260);
nand U2423 (N_2423,N_2012,N_1852);
and U2424 (N_2424,N_2019,N_1917);
or U2425 (N_2425,N_2383,N_2340);
nor U2426 (N_2426,N_2020,N_1990);
nand U2427 (N_2427,N_1867,N_2137);
nor U2428 (N_2428,N_1971,N_2271);
and U2429 (N_2429,N_2127,N_1870);
or U2430 (N_2430,N_1828,N_1940);
nand U2431 (N_2431,N_2352,N_2274);
nand U2432 (N_2432,N_1838,N_1837);
or U2433 (N_2433,N_2364,N_1991);
and U2434 (N_2434,N_2363,N_2204);
nor U2435 (N_2435,N_2201,N_1920);
or U2436 (N_2436,N_2124,N_2117);
and U2437 (N_2437,N_2197,N_2027);
xnor U2438 (N_2438,N_1967,N_1899);
and U2439 (N_2439,N_2136,N_2356);
and U2440 (N_2440,N_2314,N_2105);
nand U2441 (N_2441,N_2186,N_2292);
or U2442 (N_2442,N_2138,N_1966);
or U2443 (N_2443,N_2106,N_2131);
nand U2444 (N_2444,N_2278,N_1829);
or U2445 (N_2445,N_2195,N_2241);
or U2446 (N_2446,N_1999,N_1827);
nand U2447 (N_2447,N_2193,N_1818);
nor U2448 (N_2448,N_1815,N_2316);
and U2449 (N_2449,N_2334,N_2245);
nor U2450 (N_2450,N_2272,N_1861);
or U2451 (N_2451,N_1879,N_1869);
or U2452 (N_2452,N_2228,N_1930);
or U2453 (N_2453,N_2142,N_2129);
or U2454 (N_2454,N_2171,N_2085);
nor U2455 (N_2455,N_1910,N_1922);
nand U2456 (N_2456,N_2328,N_2030);
and U2457 (N_2457,N_1942,N_2140);
nand U2458 (N_2458,N_1854,N_2066);
and U2459 (N_2459,N_2308,N_1863);
and U2460 (N_2460,N_2287,N_2174);
and U2461 (N_2461,N_1941,N_1975);
and U2462 (N_2462,N_2045,N_1892);
and U2463 (N_2463,N_2300,N_1979);
and U2464 (N_2464,N_1950,N_1878);
and U2465 (N_2465,N_2190,N_1821);
or U2466 (N_2466,N_2092,N_2229);
and U2467 (N_2467,N_2237,N_1946);
or U2468 (N_2468,N_2044,N_2094);
xor U2469 (N_2469,N_1889,N_2379);
nand U2470 (N_2470,N_2009,N_1898);
or U2471 (N_2471,N_2160,N_1935);
nor U2472 (N_2472,N_2203,N_2232);
or U2473 (N_2473,N_2047,N_2362);
or U2474 (N_2474,N_1953,N_2388);
nand U2475 (N_2475,N_1824,N_2152);
and U2476 (N_2476,N_2215,N_2310);
and U2477 (N_2477,N_1808,N_2216);
or U2478 (N_2478,N_2088,N_1846);
and U2479 (N_2479,N_2371,N_2309);
or U2480 (N_2480,N_1853,N_2162);
or U2481 (N_2481,N_2104,N_2376);
nand U2482 (N_2482,N_2266,N_1906);
or U2483 (N_2483,N_2317,N_2144);
or U2484 (N_2484,N_2024,N_1880);
nand U2485 (N_2485,N_2373,N_1924);
or U2486 (N_2486,N_1993,N_2346);
and U2487 (N_2487,N_2313,N_1944);
and U2488 (N_2488,N_2157,N_2285);
nor U2489 (N_2489,N_1948,N_2312);
nand U2490 (N_2490,N_2208,N_1812);
nand U2491 (N_2491,N_2374,N_2217);
nor U2492 (N_2492,N_2087,N_1890);
or U2493 (N_2493,N_1998,N_2176);
nor U2494 (N_2494,N_1862,N_2050);
nor U2495 (N_2495,N_2010,N_1978);
and U2496 (N_2496,N_2235,N_1961);
nor U2497 (N_2497,N_2108,N_2282);
nand U2498 (N_2498,N_2170,N_2167);
nand U2499 (N_2499,N_2339,N_1937);
nand U2500 (N_2500,N_2178,N_2290);
nand U2501 (N_2501,N_2355,N_2249);
nand U2502 (N_2502,N_2381,N_1848);
and U2503 (N_2503,N_2065,N_2099);
nor U2504 (N_2504,N_1801,N_2211);
or U2505 (N_2505,N_2018,N_2121);
nor U2506 (N_2506,N_2213,N_1908);
nor U2507 (N_2507,N_2306,N_1938);
and U2508 (N_2508,N_2380,N_2349);
nand U2509 (N_2509,N_2016,N_1809);
and U2510 (N_2510,N_2173,N_1825);
and U2511 (N_2511,N_2329,N_2276);
and U2512 (N_2512,N_2076,N_2311);
nand U2513 (N_2513,N_2342,N_2270);
or U2514 (N_2514,N_2135,N_2107);
nor U2515 (N_2515,N_1850,N_2033);
and U2516 (N_2516,N_1866,N_2296);
nor U2517 (N_2517,N_1987,N_2321);
nand U2518 (N_2518,N_2253,N_2224);
and U2519 (N_2519,N_2335,N_1921);
or U2520 (N_2520,N_2163,N_2281);
or U2521 (N_2521,N_2097,N_2149);
nor U2522 (N_2522,N_2366,N_1980);
nand U2523 (N_2523,N_1830,N_2187);
or U2524 (N_2524,N_1855,N_2234);
nor U2525 (N_2525,N_2268,N_2307);
or U2526 (N_2526,N_2230,N_2055);
or U2527 (N_2527,N_2015,N_2021);
or U2528 (N_2528,N_2166,N_1959);
nand U2529 (N_2529,N_2191,N_1883);
or U2530 (N_2530,N_2385,N_2331);
nor U2531 (N_2531,N_2196,N_2102);
nand U2532 (N_2532,N_1843,N_2052);
and U2533 (N_2533,N_2286,N_1976);
and U2534 (N_2534,N_2233,N_1826);
nand U2535 (N_2535,N_2370,N_1817);
or U2536 (N_2536,N_1988,N_1836);
or U2537 (N_2537,N_1943,N_2082);
and U2538 (N_2538,N_2014,N_2031);
or U2539 (N_2539,N_1877,N_2188);
and U2540 (N_2540,N_1939,N_1931);
and U2541 (N_2541,N_2059,N_2155);
or U2542 (N_2542,N_2389,N_2353);
or U2543 (N_2543,N_1845,N_2397);
and U2544 (N_2544,N_2199,N_1973);
and U2545 (N_2545,N_2354,N_2075);
nand U2546 (N_2546,N_2283,N_1907);
nor U2547 (N_2547,N_2175,N_1992);
nor U2548 (N_2548,N_2212,N_1945);
and U2549 (N_2549,N_2384,N_2156);
and U2550 (N_2550,N_2299,N_2183);
nand U2551 (N_2551,N_1813,N_2327);
and U2552 (N_2552,N_1805,N_2037);
nor U2553 (N_2553,N_2264,N_2001);
nor U2554 (N_2554,N_2113,N_1800);
and U2555 (N_2555,N_2148,N_1864);
and U2556 (N_2556,N_2238,N_2069);
and U2557 (N_2557,N_2011,N_2089);
or U2558 (N_2558,N_2036,N_1984);
or U2559 (N_2559,N_2302,N_2378);
nand U2560 (N_2560,N_2080,N_2267);
nor U2561 (N_2561,N_2119,N_2038);
or U2562 (N_2562,N_2141,N_1997);
or U2563 (N_2563,N_1820,N_1806);
xnor U2564 (N_2564,N_2218,N_1964);
and U2565 (N_2565,N_2043,N_2246);
or U2566 (N_2566,N_1936,N_2256);
nand U2567 (N_2567,N_1918,N_2109);
nor U2568 (N_2568,N_2301,N_2143);
and U2569 (N_2569,N_2251,N_2189);
nand U2570 (N_2570,N_2151,N_2116);
nor U2571 (N_2571,N_2122,N_2039);
and U2572 (N_2572,N_2398,N_2095);
nor U2573 (N_2573,N_1885,N_2134);
nand U2574 (N_2574,N_1804,N_1819);
or U2575 (N_2575,N_2064,N_2275);
or U2576 (N_2576,N_2358,N_1888);
nor U2577 (N_2577,N_1949,N_2128);
and U2578 (N_2578,N_1957,N_2248);
or U2579 (N_2579,N_2305,N_2194);
nor U2580 (N_2580,N_2114,N_2063);
or U2581 (N_2581,N_1954,N_1958);
xor U2582 (N_2582,N_2257,N_2284);
nor U2583 (N_2583,N_2372,N_1859);
or U2584 (N_2584,N_2395,N_2147);
nor U2585 (N_2585,N_2185,N_1893);
nand U2586 (N_2586,N_2336,N_2158);
nand U2587 (N_2587,N_2004,N_2255);
nand U2588 (N_2588,N_2240,N_1832);
nand U2589 (N_2589,N_2288,N_2247);
and U2590 (N_2590,N_2315,N_2222);
or U2591 (N_2591,N_1873,N_2118);
nor U2592 (N_2592,N_1871,N_2123);
nor U2593 (N_2593,N_2396,N_2184);
nand U2594 (N_2594,N_2219,N_2101);
nor U2595 (N_2595,N_2351,N_1934);
or U2596 (N_2596,N_2280,N_1902);
and U2597 (N_2597,N_2338,N_2126);
nor U2598 (N_2598,N_2221,N_2304);
nor U2599 (N_2599,N_2057,N_2289);
nor U2600 (N_2600,N_2046,N_2205);
or U2601 (N_2601,N_1842,N_1925);
or U2602 (N_2602,N_1896,N_2130);
nand U2603 (N_2603,N_2111,N_2210);
or U2604 (N_2604,N_1901,N_1844);
and U2605 (N_2605,N_2243,N_1956);
nor U2606 (N_2606,N_1977,N_2258);
and U2607 (N_2607,N_2172,N_2377);
or U2608 (N_2608,N_2003,N_2161);
nand U2609 (N_2609,N_1914,N_1816);
nor U2610 (N_2610,N_1822,N_1858);
and U2611 (N_2611,N_2180,N_1904);
or U2612 (N_2612,N_1811,N_2337);
or U2613 (N_2613,N_2079,N_2081);
nor U2614 (N_2614,N_1857,N_2008);
or U2615 (N_2615,N_2056,N_2006);
or U2616 (N_2616,N_1927,N_1839);
or U2617 (N_2617,N_1913,N_1947);
and U2618 (N_2618,N_2198,N_1968);
nor U2619 (N_2619,N_2382,N_2227);
and U2620 (N_2620,N_2177,N_2025);
or U2621 (N_2621,N_2034,N_2083);
or U2622 (N_2622,N_2345,N_1831);
and U2623 (N_2623,N_1995,N_2181);
nand U2624 (N_2624,N_2239,N_2214);
or U2625 (N_2625,N_2254,N_2125);
nor U2626 (N_2626,N_2399,N_1865);
and U2627 (N_2627,N_1974,N_1983);
nand U2628 (N_2628,N_2061,N_1982);
or U2629 (N_2629,N_2073,N_2071);
xnor U2630 (N_2630,N_2392,N_1915);
and U2631 (N_2631,N_2139,N_2100);
nor U2632 (N_2632,N_2263,N_2150);
nand U2633 (N_2633,N_1989,N_2347);
or U2634 (N_2634,N_2002,N_2028);
nand U2635 (N_2635,N_1994,N_2060);
or U2636 (N_2636,N_1891,N_2322);
nand U2637 (N_2637,N_2357,N_1872);
or U2638 (N_2638,N_2367,N_2077);
nand U2639 (N_2639,N_1814,N_1970);
and U2640 (N_2640,N_2042,N_2350);
nand U2641 (N_2641,N_2273,N_2324);
nor U2642 (N_2642,N_2394,N_2086);
or U2643 (N_2643,N_1923,N_2005);
nand U2644 (N_2644,N_2110,N_2325);
or U2645 (N_2645,N_1969,N_1876);
or U2646 (N_2646,N_2182,N_2074);
or U2647 (N_2647,N_1882,N_2368);
nor U2648 (N_2648,N_1874,N_1928);
nor U2649 (N_2649,N_2231,N_1985);
and U2650 (N_2650,N_2303,N_2051);
nand U2651 (N_2651,N_2343,N_1860);
nand U2652 (N_2652,N_2048,N_2159);
and U2653 (N_2653,N_2000,N_2202);
and U2654 (N_2654,N_2220,N_2070);
nor U2655 (N_2655,N_2277,N_1963);
or U2656 (N_2656,N_1886,N_2360);
nor U2657 (N_2657,N_1932,N_1823);
nor U2658 (N_2658,N_2013,N_2053);
nor U2659 (N_2659,N_1847,N_2192);
or U2660 (N_2660,N_2090,N_2361);
nor U2661 (N_2661,N_2391,N_2279);
or U2662 (N_2662,N_1802,N_1849);
nand U2663 (N_2663,N_2026,N_1911);
and U2664 (N_2664,N_1919,N_1834);
nor U2665 (N_2665,N_1955,N_1933);
and U2666 (N_2666,N_1851,N_1905);
or U2667 (N_2667,N_2318,N_2252);
nand U2668 (N_2668,N_1840,N_1965);
nor U2669 (N_2669,N_1875,N_2250);
nor U2670 (N_2670,N_2387,N_2359);
or U2671 (N_2671,N_2007,N_2262);
nor U2672 (N_2672,N_2032,N_2096);
nand U2673 (N_2673,N_2236,N_2209);
nor U2674 (N_2674,N_2072,N_2207);
nor U2675 (N_2675,N_2320,N_2133);
or U2676 (N_2676,N_2120,N_2023);
nor U2677 (N_2677,N_2022,N_2091);
nand U2678 (N_2678,N_2049,N_2146);
nor U2679 (N_2679,N_2348,N_1960);
or U2680 (N_2680,N_2168,N_1909);
and U2681 (N_2681,N_1894,N_1833);
nand U2682 (N_2682,N_2333,N_2332);
nor U2683 (N_2683,N_1916,N_2297);
and U2684 (N_2684,N_1986,N_2035);
nand U2685 (N_2685,N_2269,N_1868);
nor U2686 (N_2686,N_1951,N_2040);
nor U2687 (N_2687,N_2058,N_1884);
or U2688 (N_2688,N_1841,N_2062);
nor U2689 (N_2689,N_2390,N_2115);
nor U2690 (N_2690,N_2067,N_1803);
and U2691 (N_2691,N_2319,N_1972);
or U2692 (N_2692,N_2200,N_1835);
nand U2693 (N_2693,N_2206,N_1895);
and U2694 (N_2694,N_1887,N_2294);
or U2695 (N_2695,N_2295,N_2365);
or U2696 (N_2696,N_2093,N_1962);
nor U2697 (N_2697,N_2054,N_1807);
nor U2698 (N_2698,N_1900,N_2164);
nand U2699 (N_2699,N_1881,N_2132);
nand U2700 (N_2700,N_2277,N_1982);
nor U2701 (N_2701,N_1805,N_2398);
and U2702 (N_2702,N_2103,N_2396);
nor U2703 (N_2703,N_2337,N_1991);
or U2704 (N_2704,N_2179,N_2383);
and U2705 (N_2705,N_1941,N_1916);
and U2706 (N_2706,N_2362,N_2251);
or U2707 (N_2707,N_2172,N_2311);
nor U2708 (N_2708,N_1815,N_1800);
nor U2709 (N_2709,N_2217,N_2223);
and U2710 (N_2710,N_1862,N_2213);
or U2711 (N_2711,N_2045,N_2234);
or U2712 (N_2712,N_2310,N_2330);
or U2713 (N_2713,N_2100,N_2067);
nand U2714 (N_2714,N_1953,N_2332);
nor U2715 (N_2715,N_2162,N_2181);
nor U2716 (N_2716,N_2029,N_2296);
or U2717 (N_2717,N_2261,N_2149);
or U2718 (N_2718,N_1965,N_1959);
and U2719 (N_2719,N_2004,N_2145);
nor U2720 (N_2720,N_2161,N_2033);
or U2721 (N_2721,N_1864,N_1820);
or U2722 (N_2722,N_2004,N_2109);
nand U2723 (N_2723,N_2166,N_1899);
nor U2724 (N_2724,N_2282,N_2338);
nand U2725 (N_2725,N_1974,N_2160);
and U2726 (N_2726,N_2259,N_2388);
nor U2727 (N_2727,N_2225,N_2211);
nor U2728 (N_2728,N_2320,N_2391);
or U2729 (N_2729,N_2033,N_1949);
nor U2730 (N_2730,N_2384,N_2236);
and U2731 (N_2731,N_2214,N_2082);
nand U2732 (N_2732,N_2255,N_2283);
nor U2733 (N_2733,N_1880,N_2187);
or U2734 (N_2734,N_2036,N_1850);
nand U2735 (N_2735,N_2224,N_2067);
nand U2736 (N_2736,N_2380,N_2207);
nand U2737 (N_2737,N_2069,N_1863);
or U2738 (N_2738,N_2104,N_2177);
nand U2739 (N_2739,N_1970,N_2397);
or U2740 (N_2740,N_1985,N_2368);
and U2741 (N_2741,N_2103,N_2275);
and U2742 (N_2742,N_2270,N_2364);
and U2743 (N_2743,N_2027,N_1984);
nand U2744 (N_2744,N_2335,N_1802);
nand U2745 (N_2745,N_2047,N_2284);
nor U2746 (N_2746,N_2064,N_2068);
and U2747 (N_2747,N_2342,N_2137);
and U2748 (N_2748,N_1935,N_2166);
xnor U2749 (N_2749,N_2040,N_2310);
or U2750 (N_2750,N_2085,N_2261);
nand U2751 (N_2751,N_2340,N_1806);
or U2752 (N_2752,N_2210,N_2039);
xor U2753 (N_2753,N_2000,N_1920);
nand U2754 (N_2754,N_1818,N_2309);
nand U2755 (N_2755,N_2284,N_1862);
nand U2756 (N_2756,N_2260,N_1843);
or U2757 (N_2757,N_2055,N_2257);
nor U2758 (N_2758,N_1929,N_2037);
or U2759 (N_2759,N_1920,N_2023);
and U2760 (N_2760,N_2396,N_2083);
nand U2761 (N_2761,N_1942,N_2028);
nand U2762 (N_2762,N_2178,N_2208);
and U2763 (N_2763,N_2397,N_2080);
nor U2764 (N_2764,N_2174,N_2259);
or U2765 (N_2765,N_1896,N_2010);
and U2766 (N_2766,N_2340,N_1932);
or U2767 (N_2767,N_2349,N_2076);
or U2768 (N_2768,N_2235,N_2221);
and U2769 (N_2769,N_2322,N_2291);
nand U2770 (N_2770,N_2342,N_2325);
and U2771 (N_2771,N_1891,N_2372);
nor U2772 (N_2772,N_2260,N_2239);
xnor U2773 (N_2773,N_2059,N_1836);
and U2774 (N_2774,N_2030,N_2003);
and U2775 (N_2775,N_1869,N_2085);
and U2776 (N_2776,N_2066,N_2253);
or U2777 (N_2777,N_2148,N_1879);
nand U2778 (N_2778,N_1899,N_1920);
xnor U2779 (N_2779,N_2392,N_2377);
nor U2780 (N_2780,N_1810,N_2214);
and U2781 (N_2781,N_1951,N_1979);
or U2782 (N_2782,N_2254,N_2270);
nand U2783 (N_2783,N_1998,N_2370);
nor U2784 (N_2784,N_1994,N_2301);
nand U2785 (N_2785,N_2359,N_2061);
or U2786 (N_2786,N_2338,N_2071);
nand U2787 (N_2787,N_1816,N_1923);
and U2788 (N_2788,N_2242,N_2144);
or U2789 (N_2789,N_2083,N_2010);
and U2790 (N_2790,N_1834,N_2210);
or U2791 (N_2791,N_1951,N_2266);
nor U2792 (N_2792,N_2160,N_2370);
and U2793 (N_2793,N_2311,N_2007);
nor U2794 (N_2794,N_2254,N_1933);
and U2795 (N_2795,N_2251,N_1913);
and U2796 (N_2796,N_1898,N_1879);
or U2797 (N_2797,N_2279,N_2388);
and U2798 (N_2798,N_2307,N_1806);
and U2799 (N_2799,N_1802,N_2209);
nor U2800 (N_2800,N_2054,N_1909);
and U2801 (N_2801,N_2386,N_2322);
nor U2802 (N_2802,N_2047,N_1810);
or U2803 (N_2803,N_1908,N_2058);
nand U2804 (N_2804,N_2015,N_1833);
or U2805 (N_2805,N_2054,N_1889);
nand U2806 (N_2806,N_1918,N_2180);
or U2807 (N_2807,N_2099,N_1978);
nand U2808 (N_2808,N_2096,N_2128);
and U2809 (N_2809,N_2082,N_1927);
or U2810 (N_2810,N_1944,N_1984);
or U2811 (N_2811,N_2099,N_2149);
nand U2812 (N_2812,N_1878,N_1973);
and U2813 (N_2813,N_2290,N_2383);
and U2814 (N_2814,N_1914,N_2173);
nor U2815 (N_2815,N_2256,N_2287);
nor U2816 (N_2816,N_2330,N_2378);
or U2817 (N_2817,N_2360,N_2329);
or U2818 (N_2818,N_2095,N_1817);
nor U2819 (N_2819,N_2360,N_2022);
nand U2820 (N_2820,N_1929,N_1870);
nor U2821 (N_2821,N_2353,N_1838);
nor U2822 (N_2822,N_2190,N_2210);
and U2823 (N_2823,N_1884,N_2316);
nand U2824 (N_2824,N_1968,N_2205);
nand U2825 (N_2825,N_2292,N_2083);
nand U2826 (N_2826,N_2109,N_2039);
and U2827 (N_2827,N_2395,N_1988);
nor U2828 (N_2828,N_2393,N_2334);
and U2829 (N_2829,N_1962,N_1951);
or U2830 (N_2830,N_2326,N_2193);
nand U2831 (N_2831,N_2286,N_2376);
or U2832 (N_2832,N_2399,N_1910);
nand U2833 (N_2833,N_2104,N_2041);
and U2834 (N_2834,N_1802,N_2123);
nor U2835 (N_2835,N_1865,N_2268);
and U2836 (N_2836,N_2153,N_2227);
and U2837 (N_2837,N_2245,N_1986);
and U2838 (N_2838,N_1858,N_2382);
and U2839 (N_2839,N_2201,N_2397);
and U2840 (N_2840,N_2251,N_2093);
nand U2841 (N_2841,N_2348,N_1956);
nor U2842 (N_2842,N_1823,N_1802);
nor U2843 (N_2843,N_2108,N_2133);
or U2844 (N_2844,N_1863,N_2330);
or U2845 (N_2845,N_2112,N_2208);
nand U2846 (N_2846,N_1975,N_1875);
and U2847 (N_2847,N_2183,N_2317);
or U2848 (N_2848,N_2355,N_2379);
nor U2849 (N_2849,N_1817,N_2028);
or U2850 (N_2850,N_2391,N_2064);
nand U2851 (N_2851,N_2270,N_1872);
nor U2852 (N_2852,N_1994,N_2103);
or U2853 (N_2853,N_1963,N_2297);
and U2854 (N_2854,N_2242,N_2265);
nor U2855 (N_2855,N_2235,N_2009);
nand U2856 (N_2856,N_2240,N_2360);
nor U2857 (N_2857,N_2124,N_1843);
nor U2858 (N_2858,N_1815,N_2027);
nor U2859 (N_2859,N_2203,N_2317);
and U2860 (N_2860,N_1821,N_1948);
and U2861 (N_2861,N_1802,N_1982);
nor U2862 (N_2862,N_1863,N_1895);
nor U2863 (N_2863,N_2007,N_2145);
and U2864 (N_2864,N_2148,N_1839);
and U2865 (N_2865,N_2387,N_1960);
or U2866 (N_2866,N_1939,N_1878);
and U2867 (N_2867,N_2247,N_2332);
or U2868 (N_2868,N_1945,N_1884);
or U2869 (N_2869,N_1922,N_2373);
and U2870 (N_2870,N_1912,N_1974);
nand U2871 (N_2871,N_1851,N_2337);
nor U2872 (N_2872,N_2287,N_2307);
and U2873 (N_2873,N_2292,N_2337);
and U2874 (N_2874,N_2183,N_2115);
and U2875 (N_2875,N_2347,N_1901);
or U2876 (N_2876,N_2354,N_1928);
and U2877 (N_2877,N_2166,N_2187);
nor U2878 (N_2878,N_1898,N_2237);
nor U2879 (N_2879,N_1878,N_2276);
nor U2880 (N_2880,N_2020,N_2099);
or U2881 (N_2881,N_1949,N_1956);
or U2882 (N_2882,N_2247,N_1834);
nand U2883 (N_2883,N_2239,N_2204);
or U2884 (N_2884,N_1884,N_2388);
or U2885 (N_2885,N_2387,N_1884);
nor U2886 (N_2886,N_2095,N_2232);
or U2887 (N_2887,N_2029,N_1979);
nand U2888 (N_2888,N_1954,N_1813);
nor U2889 (N_2889,N_2148,N_2211);
and U2890 (N_2890,N_2001,N_1962);
nor U2891 (N_2891,N_1887,N_2227);
or U2892 (N_2892,N_2031,N_1902);
or U2893 (N_2893,N_2340,N_2000);
and U2894 (N_2894,N_1810,N_2288);
and U2895 (N_2895,N_1865,N_2005);
nand U2896 (N_2896,N_2075,N_1907);
or U2897 (N_2897,N_1903,N_2098);
nand U2898 (N_2898,N_1932,N_1810);
nand U2899 (N_2899,N_1823,N_2154);
nor U2900 (N_2900,N_1860,N_1844);
nor U2901 (N_2901,N_2074,N_1900);
or U2902 (N_2902,N_2283,N_1923);
and U2903 (N_2903,N_2119,N_2292);
nand U2904 (N_2904,N_2174,N_2089);
and U2905 (N_2905,N_2081,N_1914);
and U2906 (N_2906,N_2313,N_2244);
nand U2907 (N_2907,N_1841,N_2356);
or U2908 (N_2908,N_2040,N_2395);
nand U2909 (N_2909,N_2240,N_2276);
nand U2910 (N_2910,N_1971,N_2324);
nand U2911 (N_2911,N_2306,N_2235);
xor U2912 (N_2912,N_1952,N_1885);
nand U2913 (N_2913,N_2382,N_2370);
and U2914 (N_2914,N_2156,N_1891);
nor U2915 (N_2915,N_1866,N_2178);
nand U2916 (N_2916,N_1807,N_2107);
nand U2917 (N_2917,N_2190,N_1840);
nor U2918 (N_2918,N_2071,N_1868);
nor U2919 (N_2919,N_2037,N_1867);
nor U2920 (N_2920,N_1854,N_2227);
and U2921 (N_2921,N_1819,N_1866);
nor U2922 (N_2922,N_1839,N_2212);
nor U2923 (N_2923,N_2071,N_2108);
and U2924 (N_2924,N_1850,N_2167);
or U2925 (N_2925,N_2008,N_1881);
nand U2926 (N_2926,N_2138,N_2149);
and U2927 (N_2927,N_2181,N_2032);
or U2928 (N_2928,N_2238,N_2012);
or U2929 (N_2929,N_1890,N_2356);
nand U2930 (N_2930,N_2076,N_1990);
nand U2931 (N_2931,N_2117,N_2297);
or U2932 (N_2932,N_2066,N_2390);
nor U2933 (N_2933,N_2029,N_1868);
nor U2934 (N_2934,N_2308,N_2265);
nor U2935 (N_2935,N_1915,N_2136);
nand U2936 (N_2936,N_2233,N_2039);
nand U2937 (N_2937,N_2210,N_1957);
nor U2938 (N_2938,N_1970,N_1870);
nand U2939 (N_2939,N_1895,N_2378);
or U2940 (N_2940,N_2067,N_1932);
nor U2941 (N_2941,N_2395,N_2003);
nor U2942 (N_2942,N_2103,N_2061);
nand U2943 (N_2943,N_2049,N_2034);
and U2944 (N_2944,N_1842,N_2334);
or U2945 (N_2945,N_2184,N_1939);
xor U2946 (N_2946,N_2086,N_2139);
and U2947 (N_2947,N_2305,N_2107);
and U2948 (N_2948,N_2390,N_2045);
and U2949 (N_2949,N_2119,N_1866);
or U2950 (N_2950,N_2215,N_1977);
nand U2951 (N_2951,N_1803,N_2257);
nor U2952 (N_2952,N_2135,N_2145);
nor U2953 (N_2953,N_1920,N_2311);
nand U2954 (N_2954,N_1984,N_1939);
nand U2955 (N_2955,N_2246,N_1810);
and U2956 (N_2956,N_1941,N_2249);
nor U2957 (N_2957,N_2156,N_2356);
nor U2958 (N_2958,N_2268,N_1897);
nor U2959 (N_2959,N_2161,N_1831);
nor U2960 (N_2960,N_2156,N_1986);
nand U2961 (N_2961,N_2106,N_2230);
nand U2962 (N_2962,N_2307,N_2397);
nand U2963 (N_2963,N_1974,N_2334);
or U2964 (N_2964,N_1945,N_1941);
nand U2965 (N_2965,N_1977,N_2042);
or U2966 (N_2966,N_1908,N_2041);
or U2967 (N_2967,N_2259,N_2337);
nor U2968 (N_2968,N_2154,N_1871);
nand U2969 (N_2969,N_1920,N_2142);
or U2970 (N_2970,N_2215,N_1843);
nand U2971 (N_2971,N_2099,N_2121);
and U2972 (N_2972,N_1964,N_2198);
nor U2973 (N_2973,N_2187,N_1858);
and U2974 (N_2974,N_2244,N_2083);
and U2975 (N_2975,N_2329,N_2379);
and U2976 (N_2976,N_2103,N_2330);
or U2977 (N_2977,N_2164,N_2251);
and U2978 (N_2978,N_1906,N_1888);
and U2979 (N_2979,N_2132,N_2078);
nand U2980 (N_2980,N_2248,N_2236);
nor U2981 (N_2981,N_2160,N_1901);
nor U2982 (N_2982,N_2283,N_1816);
xor U2983 (N_2983,N_2203,N_2099);
nand U2984 (N_2984,N_2238,N_2328);
xor U2985 (N_2985,N_2220,N_1978);
nand U2986 (N_2986,N_2119,N_2227);
or U2987 (N_2987,N_1912,N_1875);
nor U2988 (N_2988,N_1990,N_2008);
and U2989 (N_2989,N_2299,N_2031);
or U2990 (N_2990,N_2170,N_2367);
nand U2991 (N_2991,N_1956,N_2068);
or U2992 (N_2992,N_2397,N_2243);
xor U2993 (N_2993,N_2180,N_1988);
nor U2994 (N_2994,N_1851,N_2352);
nor U2995 (N_2995,N_1950,N_2088);
nand U2996 (N_2996,N_2225,N_1832);
nor U2997 (N_2997,N_2203,N_2069);
xnor U2998 (N_2998,N_2089,N_2219);
nor U2999 (N_2999,N_2323,N_1951);
or UO_0 (O_0,N_2927,N_2431);
nand UO_1 (O_1,N_2713,N_2768);
or UO_2 (O_2,N_2847,N_2883);
nand UO_3 (O_3,N_2425,N_2512);
nor UO_4 (O_4,N_2962,N_2774);
and UO_5 (O_5,N_2554,N_2958);
nand UO_6 (O_6,N_2828,N_2858);
nand UO_7 (O_7,N_2954,N_2724);
and UO_8 (O_8,N_2445,N_2518);
nor UO_9 (O_9,N_2886,N_2878);
and UO_10 (O_10,N_2953,N_2563);
and UO_11 (O_11,N_2844,N_2460);
or UO_12 (O_12,N_2794,N_2461);
nand UO_13 (O_13,N_2432,N_2744);
nor UO_14 (O_14,N_2994,N_2814);
xnor UO_15 (O_15,N_2449,N_2764);
and UO_16 (O_16,N_2580,N_2625);
nor UO_17 (O_17,N_2682,N_2854);
and UO_18 (O_18,N_2675,N_2423);
nor UO_19 (O_19,N_2404,N_2598);
or UO_20 (O_20,N_2785,N_2827);
nand UO_21 (O_21,N_2813,N_2446);
nand UO_22 (O_22,N_2588,N_2624);
xnor UO_23 (O_23,N_2642,N_2907);
and UO_24 (O_24,N_2478,N_2718);
or UO_25 (O_25,N_2487,N_2899);
nor UO_26 (O_26,N_2811,N_2745);
and UO_27 (O_27,N_2699,N_2845);
nor UO_28 (O_28,N_2571,N_2535);
and UO_29 (O_29,N_2505,N_2916);
or UO_30 (O_30,N_2496,N_2918);
nand UO_31 (O_31,N_2417,N_2747);
or UO_32 (O_32,N_2541,N_2671);
and UO_33 (O_33,N_2822,N_2966);
nor UO_34 (O_34,N_2702,N_2705);
nand UO_35 (O_35,N_2611,N_2997);
or UO_36 (O_36,N_2412,N_2839);
nand UO_37 (O_37,N_2659,N_2495);
nor UO_38 (O_38,N_2829,N_2818);
nor UO_39 (O_39,N_2944,N_2645);
and UO_40 (O_40,N_2665,N_2762);
nor UO_41 (O_41,N_2416,N_2900);
and UO_42 (O_42,N_2630,N_2781);
and UO_43 (O_43,N_2974,N_2585);
or UO_44 (O_44,N_2867,N_2696);
and UO_45 (O_45,N_2434,N_2464);
nand UO_46 (O_46,N_2618,N_2415);
or UO_47 (O_47,N_2808,N_2977);
or UO_48 (O_48,N_2807,N_2567);
nor UO_49 (O_49,N_2855,N_2920);
nand UO_50 (O_50,N_2908,N_2952);
or UO_51 (O_51,N_2978,N_2592);
and UO_52 (O_52,N_2467,N_2532);
nand UO_53 (O_53,N_2629,N_2976);
nor UO_54 (O_54,N_2726,N_2892);
and UO_55 (O_55,N_2817,N_2519);
nor UO_56 (O_56,N_2683,N_2407);
or UO_57 (O_57,N_2775,N_2988);
nor UO_58 (O_58,N_2837,N_2778);
and UO_59 (O_59,N_2738,N_2693);
nand UO_60 (O_60,N_2689,N_2636);
nor UO_61 (O_61,N_2969,N_2812);
and UO_62 (O_62,N_2897,N_2427);
nand UO_63 (O_63,N_2825,N_2489);
nand UO_64 (O_64,N_2979,N_2426);
and UO_65 (O_65,N_2503,N_2928);
and UO_66 (O_66,N_2529,N_2457);
nand UO_67 (O_67,N_2819,N_2681);
or UO_68 (O_68,N_2465,N_2719);
nand UO_69 (O_69,N_2802,N_2943);
or UO_70 (O_70,N_2885,N_2947);
and UO_71 (O_71,N_2884,N_2485);
nand UO_72 (O_72,N_2413,N_2430);
nor UO_73 (O_73,N_2499,N_2428);
or UO_74 (O_74,N_2685,N_2609);
and UO_75 (O_75,N_2569,N_2720);
or UO_76 (O_76,N_2621,N_2964);
and UO_77 (O_77,N_2437,N_2779);
nor UO_78 (O_78,N_2664,N_2888);
xor UO_79 (O_79,N_2836,N_2882);
and UO_80 (O_80,N_2748,N_2587);
and UO_81 (O_81,N_2677,N_2450);
nor UO_82 (O_82,N_2546,N_2619);
nor UO_83 (O_83,N_2595,N_2850);
nand UO_84 (O_84,N_2482,N_2795);
nand UO_85 (O_85,N_2983,N_2872);
nand UO_86 (O_86,N_2521,N_2631);
nor UO_87 (O_87,N_2710,N_2753);
nor UO_88 (O_88,N_2655,N_2520);
or UO_89 (O_89,N_2833,N_2863);
nand UO_90 (O_90,N_2560,N_2422);
nor UO_91 (O_91,N_2627,N_2725);
or UO_92 (O_92,N_2590,N_2634);
or UO_93 (O_93,N_2763,N_2687);
nand UO_94 (O_94,N_2490,N_2824);
nor UO_95 (O_95,N_2670,N_2418);
nand UO_96 (O_96,N_2772,N_2477);
nand UO_97 (O_97,N_2454,N_2956);
nand UO_98 (O_98,N_2999,N_2647);
nor UO_99 (O_99,N_2408,N_2643);
nor UO_100 (O_100,N_2755,N_2965);
nor UO_101 (O_101,N_2919,N_2565);
and UO_102 (O_102,N_2946,N_2798);
nand UO_103 (O_103,N_2780,N_2934);
nor UO_104 (O_104,N_2752,N_2804);
and UO_105 (O_105,N_2514,N_2853);
nor UO_106 (O_106,N_2852,N_2501);
nor UO_107 (O_107,N_2568,N_2949);
and UO_108 (O_108,N_2517,N_2448);
and UO_109 (O_109,N_2701,N_2515);
nand UO_110 (O_110,N_2821,N_2690);
and UO_111 (O_111,N_2877,N_2424);
nand UO_112 (O_112,N_2938,N_2791);
nor UO_113 (O_113,N_2931,N_2547);
and UO_114 (O_114,N_2474,N_2623);
nor UO_115 (O_115,N_2576,N_2473);
nand UO_116 (O_116,N_2991,N_2589);
and UO_117 (O_117,N_2494,N_2522);
or UO_118 (O_118,N_2635,N_2471);
nand UO_119 (O_119,N_2507,N_2708);
or UO_120 (O_120,N_2572,N_2736);
nor UO_121 (O_121,N_2620,N_2536);
or UO_122 (O_122,N_2672,N_2865);
nand UO_123 (O_123,N_2714,N_2508);
nor UO_124 (O_124,N_2868,N_2816);
nand UO_125 (O_125,N_2472,N_2929);
or UO_126 (O_126,N_2806,N_2926);
nor UO_127 (O_127,N_2866,N_2901);
xnor UO_128 (O_128,N_2556,N_2729);
and UO_129 (O_129,N_2841,N_2746);
nand UO_130 (O_130,N_2948,N_2668);
and UO_131 (O_131,N_2530,N_2796);
nand UO_132 (O_132,N_2754,N_2993);
nand UO_133 (O_133,N_2443,N_2475);
or UO_134 (O_134,N_2578,N_2971);
nor UO_135 (O_135,N_2715,N_2596);
nor UO_136 (O_136,N_2638,N_2960);
xnor UO_137 (O_137,N_2469,N_2550);
and UO_138 (O_138,N_2921,N_2909);
nor UO_139 (O_139,N_2769,N_2455);
and UO_140 (O_140,N_2698,N_2923);
nor UO_141 (O_141,N_2980,N_2447);
and UO_142 (O_142,N_2653,N_2941);
nand UO_143 (O_143,N_2637,N_2893);
nand UO_144 (O_144,N_2728,N_2810);
nand UO_145 (O_145,N_2905,N_2711);
and UO_146 (O_146,N_2497,N_2722);
and UO_147 (O_147,N_2777,N_2986);
or UO_148 (O_148,N_2509,N_2786);
nand UO_149 (O_149,N_2996,N_2985);
nor UO_150 (O_150,N_2875,N_2442);
xor UO_151 (O_151,N_2959,N_2483);
nor UO_152 (O_152,N_2641,N_2933);
nor UO_153 (O_153,N_2502,N_2622);
and UO_154 (O_154,N_2771,N_2640);
nor UO_155 (O_155,N_2684,N_2930);
nand UO_156 (O_156,N_2479,N_2990);
nor UO_157 (O_157,N_2604,N_2743);
nand UO_158 (O_158,N_2680,N_2703);
nand UO_159 (O_159,N_2435,N_2616);
nor UO_160 (O_160,N_2552,N_2481);
nand UO_161 (O_161,N_2402,N_2906);
nand UO_162 (O_162,N_2770,N_2864);
nand UO_163 (O_163,N_2429,N_2626);
nand UO_164 (O_164,N_2995,N_2881);
and UO_165 (O_165,N_2871,N_2749);
or UO_166 (O_166,N_2876,N_2591);
nor UO_167 (O_167,N_2498,N_2543);
or UO_168 (O_168,N_2484,N_2527);
nand UO_169 (O_169,N_2932,N_2851);
and UO_170 (O_170,N_2524,N_2688);
nor UO_171 (O_171,N_2551,N_2444);
and UO_172 (O_172,N_2896,N_2579);
nand UO_173 (O_173,N_2523,N_2528);
and UO_174 (O_174,N_2712,N_2835);
nand UO_175 (O_175,N_2406,N_2678);
and UO_176 (O_176,N_2793,N_2451);
nor UO_177 (O_177,N_2697,N_2615);
nor UO_178 (O_178,N_2599,N_2957);
nor UO_179 (O_179,N_2555,N_2511);
nand UO_180 (O_180,N_2925,N_2717);
nand UO_181 (O_181,N_2666,N_2575);
nor UO_182 (O_182,N_2742,N_2767);
nand UO_183 (O_183,N_2913,N_2564);
nand UO_184 (O_184,N_2984,N_2648);
or UO_185 (O_185,N_2761,N_2750);
nand UO_186 (O_186,N_2758,N_2950);
nor UO_187 (O_187,N_2730,N_2727);
nand UO_188 (O_188,N_2662,N_2759);
and UO_189 (O_189,N_2739,N_2760);
and UO_190 (O_190,N_2776,N_2601);
nand UO_191 (O_191,N_2549,N_2911);
nor UO_192 (O_192,N_2751,N_2577);
nor UO_193 (O_193,N_2792,N_2782);
nand UO_194 (O_194,N_2452,N_2639);
and UO_195 (O_195,N_2438,N_2773);
and UO_196 (O_196,N_2797,N_2633);
nand UO_197 (O_197,N_2663,N_2721);
nand UO_198 (O_198,N_2973,N_2951);
and UO_199 (O_199,N_2910,N_2613);
and UO_200 (O_200,N_2686,N_2525);
or UO_201 (O_201,N_2963,N_2891);
nand UO_202 (O_202,N_2842,N_2840);
nor UO_203 (O_203,N_2492,N_2936);
nand UO_204 (O_204,N_2644,N_2832);
nor UO_205 (O_205,N_2573,N_2846);
nor UO_206 (O_206,N_2656,N_2940);
nand UO_207 (O_207,N_2981,N_2895);
or UO_208 (O_208,N_2924,N_2661);
or UO_209 (O_209,N_2790,N_2695);
nand UO_210 (O_210,N_2654,N_2676);
and UO_211 (O_211,N_2410,N_2470);
and UO_212 (O_212,N_2740,N_2400);
nor UO_213 (O_213,N_2539,N_2917);
xor UO_214 (O_214,N_2862,N_2800);
and UO_215 (O_215,N_2756,N_2561);
nand UO_216 (O_216,N_2405,N_2436);
or UO_217 (O_217,N_2998,N_2803);
nand UO_218 (O_218,N_2716,N_2510);
nand UO_219 (O_219,N_2935,N_2857);
nor UO_220 (O_220,N_2757,N_2433);
and UO_221 (O_221,N_2870,N_2830);
or UO_222 (O_222,N_2732,N_2922);
nor UO_223 (O_223,N_2879,N_2733);
or UO_224 (O_224,N_2904,N_2506);
or UO_225 (O_225,N_2513,N_2945);
or UO_226 (O_226,N_2860,N_2468);
or UO_227 (O_227,N_2600,N_2674);
nand UO_228 (O_228,N_2890,N_2788);
and UO_229 (O_229,N_2861,N_2440);
nand UO_230 (O_230,N_2784,N_2843);
and UO_231 (O_231,N_2669,N_2700);
nor UO_232 (O_232,N_2559,N_2657);
nor UO_233 (O_233,N_2838,N_2915);
nor UO_234 (O_234,N_2912,N_2799);
nand UO_235 (O_235,N_2741,N_2617);
and UO_236 (O_236,N_2462,N_2765);
and UO_237 (O_237,N_2570,N_2734);
or UO_238 (O_238,N_2558,N_2614);
nor UO_239 (O_239,N_2651,N_2859);
nand UO_240 (O_240,N_2874,N_2584);
xnor UO_241 (O_241,N_2608,N_2889);
or UO_242 (O_242,N_2658,N_2834);
or UO_243 (O_243,N_2602,N_2403);
or UO_244 (O_244,N_2610,N_2463);
nand UO_245 (O_245,N_2593,N_2419);
or UO_246 (O_246,N_2439,N_2731);
nand UO_247 (O_247,N_2476,N_2540);
nand UO_248 (O_248,N_2831,N_2970);
nand UO_249 (O_249,N_2414,N_2420);
nor UO_250 (O_250,N_2605,N_2537);
nand UO_251 (O_251,N_2491,N_2823);
nand UO_252 (O_252,N_2937,N_2486);
nor UO_253 (O_253,N_2694,N_2603);
xnor UO_254 (O_254,N_2989,N_2453);
nor UO_255 (O_255,N_2820,N_2704);
and UO_256 (O_256,N_2606,N_2488);
nor UO_257 (O_257,N_2707,N_2848);
nor UO_258 (O_258,N_2673,N_2516);
nor UO_259 (O_259,N_2667,N_2581);
nand UO_260 (O_260,N_2493,N_2809);
or UO_261 (O_261,N_2939,N_2456);
nand UO_262 (O_262,N_2480,N_2574);
and UO_263 (O_263,N_2914,N_2735);
nor UO_264 (O_264,N_2898,N_2982);
nand UO_265 (O_265,N_2805,N_2566);
nand UO_266 (O_266,N_2826,N_2894);
nand UO_267 (O_267,N_2500,N_2903);
xnor UO_268 (O_268,N_2801,N_2992);
nor UO_269 (O_269,N_2562,N_2504);
nand UO_270 (O_270,N_2538,N_2526);
xnor UO_271 (O_271,N_2545,N_2632);
nand UO_272 (O_272,N_2628,N_2534);
and UO_273 (O_273,N_2968,N_2869);
and UO_274 (O_274,N_2649,N_2955);
nand UO_275 (O_275,N_2975,N_2646);
and UO_276 (O_276,N_2548,N_2533);
nor UO_277 (O_277,N_2586,N_2542);
nand UO_278 (O_278,N_2607,N_2466);
nand UO_279 (O_279,N_2692,N_2582);
or UO_280 (O_280,N_2583,N_2679);
or UO_281 (O_281,N_2887,N_2660);
and UO_282 (O_282,N_2691,N_2652);
nor UO_283 (O_283,N_2459,N_2553);
or UO_284 (O_284,N_2612,N_2409);
or UO_285 (O_285,N_2815,N_2723);
nor UO_286 (O_286,N_2967,N_2458);
nand UO_287 (O_287,N_2987,N_2441);
nand UO_288 (O_288,N_2531,N_2709);
xor UO_289 (O_289,N_2597,N_2706);
and UO_290 (O_290,N_2789,N_2873);
and UO_291 (O_291,N_2594,N_2942);
xor UO_292 (O_292,N_2411,N_2972);
nand UO_293 (O_293,N_2544,N_2783);
and UO_294 (O_294,N_2766,N_2961);
nor UO_295 (O_295,N_2880,N_2557);
nand UO_296 (O_296,N_2737,N_2787);
and UO_297 (O_297,N_2650,N_2856);
xnor UO_298 (O_298,N_2849,N_2401);
and UO_299 (O_299,N_2902,N_2421);
and UO_300 (O_300,N_2610,N_2668);
nor UO_301 (O_301,N_2994,N_2839);
or UO_302 (O_302,N_2916,N_2577);
and UO_303 (O_303,N_2771,N_2500);
or UO_304 (O_304,N_2535,N_2724);
nand UO_305 (O_305,N_2911,N_2914);
nor UO_306 (O_306,N_2488,N_2588);
and UO_307 (O_307,N_2830,N_2523);
nand UO_308 (O_308,N_2659,N_2885);
nand UO_309 (O_309,N_2514,N_2757);
nor UO_310 (O_310,N_2998,N_2459);
nor UO_311 (O_311,N_2684,N_2417);
nand UO_312 (O_312,N_2830,N_2853);
nand UO_313 (O_313,N_2901,N_2841);
nand UO_314 (O_314,N_2469,N_2521);
nor UO_315 (O_315,N_2482,N_2660);
nor UO_316 (O_316,N_2898,N_2941);
xor UO_317 (O_317,N_2859,N_2605);
or UO_318 (O_318,N_2517,N_2540);
nand UO_319 (O_319,N_2908,N_2766);
or UO_320 (O_320,N_2944,N_2947);
or UO_321 (O_321,N_2614,N_2624);
and UO_322 (O_322,N_2590,N_2717);
or UO_323 (O_323,N_2403,N_2413);
nand UO_324 (O_324,N_2968,N_2851);
nand UO_325 (O_325,N_2495,N_2536);
or UO_326 (O_326,N_2958,N_2403);
nand UO_327 (O_327,N_2435,N_2935);
or UO_328 (O_328,N_2697,N_2888);
or UO_329 (O_329,N_2795,N_2751);
nor UO_330 (O_330,N_2846,N_2813);
and UO_331 (O_331,N_2975,N_2690);
nand UO_332 (O_332,N_2416,N_2644);
or UO_333 (O_333,N_2985,N_2557);
nand UO_334 (O_334,N_2851,N_2879);
or UO_335 (O_335,N_2442,N_2515);
or UO_336 (O_336,N_2843,N_2844);
nand UO_337 (O_337,N_2848,N_2467);
or UO_338 (O_338,N_2944,N_2973);
xor UO_339 (O_339,N_2490,N_2989);
and UO_340 (O_340,N_2550,N_2701);
and UO_341 (O_341,N_2627,N_2946);
or UO_342 (O_342,N_2984,N_2483);
nand UO_343 (O_343,N_2593,N_2824);
or UO_344 (O_344,N_2704,N_2430);
xor UO_345 (O_345,N_2660,N_2970);
nand UO_346 (O_346,N_2721,N_2699);
xnor UO_347 (O_347,N_2494,N_2606);
and UO_348 (O_348,N_2875,N_2467);
nor UO_349 (O_349,N_2797,N_2449);
nand UO_350 (O_350,N_2573,N_2458);
or UO_351 (O_351,N_2660,N_2739);
and UO_352 (O_352,N_2439,N_2678);
or UO_353 (O_353,N_2989,N_2824);
and UO_354 (O_354,N_2705,N_2917);
or UO_355 (O_355,N_2457,N_2753);
or UO_356 (O_356,N_2887,N_2545);
and UO_357 (O_357,N_2544,N_2878);
or UO_358 (O_358,N_2861,N_2905);
and UO_359 (O_359,N_2579,N_2494);
nor UO_360 (O_360,N_2533,N_2508);
nor UO_361 (O_361,N_2706,N_2816);
nor UO_362 (O_362,N_2697,N_2937);
xnor UO_363 (O_363,N_2663,N_2832);
nand UO_364 (O_364,N_2684,N_2538);
and UO_365 (O_365,N_2492,N_2455);
and UO_366 (O_366,N_2835,N_2814);
xor UO_367 (O_367,N_2975,N_2810);
or UO_368 (O_368,N_2972,N_2768);
nor UO_369 (O_369,N_2456,N_2593);
and UO_370 (O_370,N_2784,N_2921);
and UO_371 (O_371,N_2788,N_2627);
or UO_372 (O_372,N_2806,N_2828);
nand UO_373 (O_373,N_2435,N_2572);
nor UO_374 (O_374,N_2798,N_2490);
or UO_375 (O_375,N_2758,N_2631);
and UO_376 (O_376,N_2653,N_2647);
or UO_377 (O_377,N_2746,N_2485);
or UO_378 (O_378,N_2882,N_2991);
or UO_379 (O_379,N_2965,N_2837);
and UO_380 (O_380,N_2543,N_2823);
nor UO_381 (O_381,N_2796,N_2856);
nor UO_382 (O_382,N_2570,N_2510);
xnor UO_383 (O_383,N_2668,N_2430);
or UO_384 (O_384,N_2728,N_2563);
nor UO_385 (O_385,N_2530,N_2960);
or UO_386 (O_386,N_2524,N_2751);
nor UO_387 (O_387,N_2815,N_2555);
nor UO_388 (O_388,N_2447,N_2497);
and UO_389 (O_389,N_2721,N_2693);
or UO_390 (O_390,N_2750,N_2620);
nor UO_391 (O_391,N_2516,N_2996);
nand UO_392 (O_392,N_2740,N_2708);
or UO_393 (O_393,N_2760,N_2664);
and UO_394 (O_394,N_2616,N_2491);
nand UO_395 (O_395,N_2727,N_2570);
nor UO_396 (O_396,N_2588,N_2445);
nand UO_397 (O_397,N_2506,N_2955);
or UO_398 (O_398,N_2604,N_2791);
or UO_399 (O_399,N_2704,N_2613);
and UO_400 (O_400,N_2896,N_2649);
and UO_401 (O_401,N_2970,N_2545);
nor UO_402 (O_402,N_2670,N_2514);
xor UO_403 (O_403,N_2701,N_2608);
or UO_404 (O_404,N_2660,N_2917);
nand UO_405 (O_405,N_2962,N_2626);
or UO_406 (O_406,N_2949,N_2408);
or UO_407 (O_407,N_2456,N_2644);
and UO_408 (O_408,N_2421,N_2638);
nor UO_409 (O_409,N_2932,N_2882);
nand UO_410 (O_410,N_2807,N_2836);
and UO_411 (O_411,N_2428,N_2429);
nand UO_412 (O_412,N_2641,N_2521);
and UO_413 (O_413,N_2986,N_2727);
and UO_414 (O_414,N_2409,N_2734);
nand UO_415 (O_415,N_2828,N_2907);
or UO_416 (O_416,N_2917,N_2740);
and UO_417 (O_417,N_2725,N_2962);
or UO_418 (O_418,N_2563,N_2856);
nand UO_419 (O_419,N_2865,N_2657);
or UO_420 (O_420,N_2850,N_2825);
nand UO_421 (O_421,N_2644,N_2945);
or UO_422 (O_422,N_2826,N_2682);
nand UO_423 (O_423,N_2769,N_2456);
or UO_424 (O_424,N_2627,N_2848);
or UO_425 (O_425,N_2736,N_2983);
nor UO_426 (O_426,N_2826,N_2578);
and UO_427 (O_427,N_2806,N_2567);
or UO_428 (O_428,N_2583,N_2938);
nand UO_429 (O_429,N_2648,N_2440);
or UO_430 (O_430,N_2924,N_2999);
nand UO_431 (O_431,N_2577,N_2544);
xnor UO_432 (O_432,N_2799,N_2919);
or UO_433 (O_433,N_2671,N_2890);
nor UO_434 (O_434,N_2632,N_2798);
and UO_435 (O_435,N_2912,N_2987);
or UO_436 (O_436,N_2968,N_2425);
or UO_437 (O_437,N_2600,N_2830);
nand UO_438 (O_438,N_2461,N_2493);
or UO_439 (O_439,N_2521,N_2751);
nor UO_440 (O_440,N_2852,N_2553);
or UO_441 (O_441,N_2433,N_2901);
and UO_442 (O_442,N_2751,N_2559);
or UO_443 (O_443,N_2623,N_2974);
and UO_444 (O_444,N_2485,N_2465);
nand UO_445 (O_445,N_2784,N_2499);
nor UO_446 (O_446,N_2861,N_2935);
and UO_447 (O_447,N_2467,N_2934);
nor UO_448 (O_448,N_2673,N_2946);
and UO_449 (O_449,N_2745,N_2742);
and UO_450 (O_450,N_2518,N_2686);
nand UO_451 (O_451,N_2757,N_2454);
nor UO_452 (O_452,N_2956,N_2992);
nand UO_453 (O_453,N_2577,N_2472);
and UO_454 (O_454,N_2757,N_2682);
or UO_455 (O_455,N_2992,N_2537);
nand UO_456 (O_456,N_2428,N_2516);
and UO_457 (O_457,N_2943,N_2424);
nand UO_458 (O_458,N_2833,N_2986);
or UO_459 (O_459,N_2941,N_2493);
or UO_460 (O_460,N_2598,N_2602);
or UO_461 (O_461,N_2829,N_2827);
nor UO_462 (O_462,N_2430,N_2929);
xor UO_463 (O_463,N_2867,N_2897);
nor UO_464 (O_464,N_2863,N_2998);
or UO_465 (O_465,N_2466,N_2557);
or UO_466 (O_466,N_2831,N_2636);
or UO_467 (O_467,N_2660,N_2543);
nand UO_468 (O_468,N_2941,N_2592);
nor UO_469 (O_469,N_2733,N_2740);
or UO_470 (O_470,N_2994,N_2439);
or UO_471 (O_471,N_2491,N_2529);
nand UO_472 (O_472,N_2801,N_2663);
or UO_473 (O_473,N_2799,N_2830);
nor UO_474 (O_474,N_2859,N_2649);
nand UO_475 (O_475,N_2648,N_2929);
nor UO_476 (O_476,N_2581,N_2871);
nand UO_477 (O_477,N_2655,N_2999);
nor UO_478 (O_478,N_2870,N_2433);
nor UO_479 (O_479,N_2450,N_2818);
nor UO_480 (O_480,N_2858,N_2458);
nor UO_481 (O_481,N_2947,N_2572);
nand UO_482 (O_482,N_2506,N_2595);
and UO_483 (O_483,N_2645,N_2701);
nor UO_484 (O_484,N_2817,N_2694);
nor UO_485 (O_485,N_2871,N_2826);
nor UO_486 (O_486,N_2756,N_2406);
nor UO_487 (O_487,N_2873,N_2650);
and UO_488 (O_488,N_2901,N_2540);
or UO_489 (O_489,N_2851,N_2871);
nand UO_490 (O_490,N_2749,N_2613);
and UO_491 (O_491,N_2472,N_2913);
or UO_492 (O_492,N_2600,N_2948);
nand UO_493 (O_493,N_2626,N_2557);
and UO_494 (O_494,N_2998,N_2599);
or UO_495 (O_495,N_2484,N_2777);
nand UO_496 (O_496,N_2610,N_2552);
and UO_497 (O_497,N_2435,N_2415);
and UO_498 (O_498,N_2669,N_2705);
xor UO_499 (O_499,N_2932,N_2686);
endmodule