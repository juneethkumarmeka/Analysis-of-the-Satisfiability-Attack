module basic_2500_25000_3000_10_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_2045,In_1157);
nand U1 (N_1,In_1176,In_1291);
nand U2 (N_2,In_2059,In_1671);
nand U3 (N_3,In_2457,In_1325);
xnor U4 (N_4,In_1020,In_887);
nand U5 (N_5,In_1272,In_1760);
xnor U6 (N_6,In_2134,In_2246);
nand U7 (N_7,In_729,In_1452);
nand U8 (N_8,In_820,In_2399);
xor U9 (N_9,In_2170,In_971);
or U10 (N_10,In_1742,In_1113);
nor U11 (N_11,In_2097,In_476);
xnor U12 (N_12,In_1693,In_544);
nor U13 (N_13,In_1399,In_2112);
nor U14 (N_14,In_2317,In_1493);
or U15 (N_15,In_1567,In_1647);
nand U16 (N_16,In_648,In_842);
nor U17 (N_17,In_1966,In_1489);
nand U18 (N_18,In_854,In_1562);
xor U19 (N_19,In_2055,In_345);
xor U20 (N_20,In_2079,In_1215);
nand U21 (N_21,In_1505,In_1158);
and U22 (N_22,In_428,In_610);
xor U23 (N_23,In_1343,In_1889);
nand U24 (N_24,In_1495,In_808);
and U25 (N_25,In_756,In_2042);
nand U26 (N_26,In_167,In_970);
xnor U27 (N_27,In_2029,In_1858);
nand U28 (N_28,In_1256,In_1131);
nand U29 (N_29,In_165,In_1884);
nor U30 (N_30,In_1880,In_2220);
xnor U31 (N_31,In_1804,In_38);
nand U32 (N_32,In_456,In_1179);
or U33 (N_33,In_1756,In_1401);
nand U34 (N_34,In_1278,In_2251);
or U35 (N_35,In_653,In_1270);
xor U36 (N_36,In_1981,In_1682);
nor U37 (N_37,In_1108,In_1586);
nand U38 (N_38,In_241,In_1751);
and U39 (N_39,In_635,In_1826);
and U40 (N_40,In_2027,In_1442);
xnor U41 (N_41,In_251,In_1919);
xor U42 (N_42,In_154,In_1532);
nor U43 (N_43,In_2214,In_56);
nor U44 (N_44,In_291,In_677);
nand U45 (N_45,In_1873,In_1651);
and U46 (N_46,In_1725,In_2314);
and U47 (N_47,In_246,In_301);
or U48 (N_48,In_1887,In_238);
nor U49 (N_49,In_1095,In_2232);
or U50 (N_50,In_1320,In_2295);
nor U51 (N_51,In_1539,In_48);
nor U52 (N_52,In_464,In_1920);
xnor U53 (N_53,In_2224,In_614);
xnor U54 (N_54,In_2358,In_2233);
and U55 (N_55,In_1211,In_2350);
nor U56 (N_56,In_1890,In_2070);
nor U57 (N_57,In_906,In_181);
xor U58 (N_58,In_871,In_316);
or U59 (N_59,In_323,In_1746);
xor U60 (N_60,In_2156,In_2092);
nor U61 (N_61,In_829,In_58);
nand U62 (N_62,In_626,In_269);
and U63 (N_63,In_2162,In_1446);
or U64 (N_64,In_1697,In_1861);
nor U65 (N_65,In_2040,In_1555);
nand U66 (N_66,In_1012,In_1354);
nor U67 (N_67,In_795,In_1986);
xor U68 (N_68,In_2461,In_2274);
nor U69 (N_69,In_473,In_2261);
nand U70 (N_70,In_1909,In_72);
xor U71 (N_71,In_1512,In_333);
or U72 (N_72,In_1976,In_1075);
or U73 (N_73,In_2160,In_1266);
or U74 (N_74,In_2416,In_2106);
and U75 (N_75,In_1043,In_89);
xnor U76 (N_76,In_311,In_1249);
and U77 (N_77,In_2163,In_1750);
nand U78 (N_78,In_1772,In_1276);
and U79 (N_79,In_1968,In_805);
nor U80 (N_80,In_1246,In_1782);
nand U81 (N_81,In_1853,In_2094);
or U82 (N_82,In_2252,In_1662);
nand U83 (N_83,In_764,In_2436);
nand U84 (N_84,In_161,In_2310);
or U85 (N_85,In_1810,In_1953);
and U86 (N_86,In_368,In_1993);
xor U87 (N_87,In_617,In_500);
xnor U88 (N_88,In_1159,In_2153);
xnor U89 (N_89,In_1842,In_668);
xor U90 (N_90,In_1087,In_309);
or U91 (N_91,In_1921,In_1600);
and U92 (N_92,In_23,In_230);
nor U93 (N_93,In_200,In_1596);
or U94 (N_94,In_1235,In_1959);
or U95 (N_95,In_256,In_1857);
nand U96 (N_96,In_272,In_902);
or U97 (N_97,In_594,In_1002);
or U98 (N_98,In_217,In_1406);
xor U99 (N_99,In_460,In_1585);
and U100 (N_100,In_703,In_2419);
nor U101 (N_101,In_1089,In_117);
nand U102 (N_102,In_342,In_1488);
nor U103 (N_103,In_650,In_714);
or U104 (N_104,In_273,In_1508);
xnor U105 (N_105,In_352,In_262);
nor U106 (N_106,In_1450,In_107);
and U107 (N_107,In_2303,In_1797);
xnor U108 (N_108,In_2331,In_81);
xnor U109 (N_109,In_694,In_799);
xnor U110 (N_110,In_6,In_1269);
xnor U111 (N_111,In_454,In_576);
or U112 (N_112,In_1455,In_1244);
nor U113 (N_113,In_233,In_1286);
nand U114 (N_114,In_1610,In_2392);
nor U115 (N_115,In_914,In_1373);
nand U116 (N_116,In_2361,In_2101);
or U117 (N_117,In_671,In_13);
nand U118 (N_118,In_1118,In_1328);
or U119 (N_119,In_568,In_407);
xnor U120 (N_120,In_1901,In_1498);
xor U121 (N_121,In_2277,In_156);
xor U122 (N_122,In_1879,In_1552);
or U123 (N_123,In_402,In_227);
nand U124 (N_124,In_1622,In_1342);
nand U125 (N_125,In_410,In_1680);
xor U126 (N_126,In_511,In_2394);
nand U127 (N_127,In_2180,In_560);
or U128 (N_128,In_1597,In_478);
xor U129 (N_129,In_2213,In_2080);
nor U130 (N_130,In_1732,In_2406);
or U131 (N_131,In_27,In_2397);
xnor U132 (N_132,In_788,In_1308);
nand U133 (N_133,In_1471,In_1515);
xor U134 (N_134,In_494,In_191);
xor U135 (N_135,In_296,In_1413);
xor U136 (N_136,In_1188,In_1329);
nor U137 (N_137,In_1699,In_85);
or U138 (N_138,In_2169,In_840);
xnor U139 (N_139,In_125,In_639);
xnor U140 (N_140,In_681,In_78);
nor U141 (N_141,In_1056,In_986);
and U142 (N_142,In_1171,In_2304);
xnor U143 (N_143,In_87,In_212);
nor U144 (N_144,In_430,In_477);
or U145 (N_145,In_2328,In_841);
nor U146 (N_146,In_1007,In_451);
and U147 (N_147,In_2433,In_510);
nor U148 (N_148,In_1526,In_600);
xnor U149 (N_149,In_905,In_791);
nand U150 (N_150,In_395,In_2147);
nor U151 (N_151,In_1813,In_1685);
and U152 (N_152,In_858,In_2129);
and U153 (N_153,In_886,In_2119);
xnor U154 (N_154,In_1619,In_1008);
nand U155 (N_155,In_355,In_2105);
and U156 (N_156,In_935,In_818);
and U157 (N_157,In_1936,In_1423);
and U158 (N_158,In_1520,In_258);
nor U159 (N_159,In_1058,In_2004);
or U160 (N_160,In_526,In_114);
xnor U161 (N_161,In_1200,In_1883);
xor U162 (N_162,In_573,In_1633);
xor U163 (N_163,In_720,In_103);
xnor U164 (N_164,In_1740,In_972);
xor U165 (N_165,In_855,In_109);
and U166 (N_166,In_2276,In_376);
xor U167 (N_167,In_1061,In_2435);
nand U168 (N_168,In_1961,In_1963);
or U169 (N_169,In_226,In_1326);
or U170 (N_170,In_2269,In_2316);
xnor U171 (N_171,In_1848,In_1763);
nand U172 (N_172,In_540,In_2175);
nand U173 (N_173,In_1241,In_1440);
or U174 (N_174,In_969,In_1196);
or U175 (N_175,In_5,In_2149);
nand U176 (N_176,In_1777,In_1138);
nand U177 (N_177,In_1924,In_1709);
xnor U178 (N_178,In_659,In_961);
nand U179 (N_179,In_1482,In_913);
nor U180 (N_180,In_892,In_877);
xnor U181 (N_181,In_1139,In_1941);
xor U182 (N_182,In_2288,In_1033);
nor U183 (N_183,In_1727,In_197);
and U184 (N_184,In_2228,In_1353);
and U185 (N_185,In_2297,In_1823);
and U186 (N_186,In_2008,In_1566);
nand U187 (N_187,In_2302,In_1120);
nand U188 (N_188,In_189,In_960);
and U189 (N_189,In_926,In_2067);
nand U190 (N_190,In_784,In_1004);
nand U191 (N_191,In_1722,In_1467);
xor U192 (N_192,In_353,In_2155);
or U193 (N_193,In_1678,In_680);
and U194 (N_194,In_995,In_2352);
nor U195 (N_195,In_2061,In_849);
or U196 (N_196,In_1057,In_2192);
xor U197 (N_197,In_819,In_944);
or U198 (N_198,In_959,In_658);
and U199 (N_199,In_1458,In_664);
or U200 (N_200,In_900,In_257);
nand U201 (N_201,In_1184,In_437);
and U202 (N_202,In_925,In_1126);
or U203 (N_203,In_1666,In_1538);
or U204 (N_204,In_804,In_1821);
nor U205 (N_205,In_2211,In_1970);
xnor U206 (N_206,In_1793,In_2071);
nor U207 (N_207,In_1124,In_2474);
xor U208 (N_208,In_1192,In_991);
nand U209 (N_209,In_2076,In_555);
nand U210 (N_210,In_438,In_401);
and U211 (N_211,In_2482,In_1983);
xnor U212 (N_212,In_661,In_240);
xnor U213 (N_213,In_14,In_1207);
or U214 (N_214,In_1876,In_1389);
and U215 (N_215,In_457,In_2047);
xnor U216 (N_216,In_2410,In_380);
nand U217 (N_217,In_1477,In_259);
nand U218 (N_218,In_1845,In_1888);
nor U219 (N_219,In_973,In_274);
xor U220 (N_220,In_1439,In_2283);
xnor U221 (N_221,In_2108,In_2034);
or U222 (N_222,In_255,In_562);
and U223 (N_223,In_1726,In_351);
or U224 (N_224,In_119,In_807);
and U225 (N_225,In_232,In_2247);
xor U226 (N_226,In_751,In_597);
or U227 (N_227,In_1761,In_357);
nor U228 (N_228,In_2014,In_318);
and U229 (N_229,In_1815,In_498);
xnor U230 (N_230,In_1851,In_1136);
nor U231 (N_231,In_554,In_299);
xor U232 (N_232,In_243,In_1469);
or U233 (N_233,In_739,In_2370);
and U234 (N_234,In_2275,In_1205);
nor U235 (N_235,In_1754,In_493);
nor U236 (N_236,In_725,In_1724);
xor U237 (N_237,In_1836,In_1630);
and U238 (N_238,In_2376,In_2333);
nand U239 (N_239,In_1571,In_1068);
nand U240 (N_240,In_2087,In_63);
or U241 (N_241,In_2237,In_2238);
xnor U242 (N_242,In_1623,In_542);
nand U243 (N_243,In_1425,In_224);
xor U244 (N_244,In_1170,In_1965);
and U245 (N_245,In_2300,In_1369);
nor U246 (N_246,In_327,In_1400);
and U247 (N_247,In_1796,In_2496);
xor U248 (N_248,In_1510,In_1522);
nand U249 (N_249,In_2452,In_1214);
and U250 (N_250,In_2098,In_2064);
nor U251 (N_251,In_2033,In_1649);
or U252 (N_252,In_518,In_848);
or U253 (N_253,In_1799,In_1582);
xnor U254 (N_254,In_644,In_1577);
nand U255 (N_255,In_461,In_1317);
xor U256 (N_256,In_1125,In_1091);
nand U257 (N_257,In_2423,In_2017);
nor U258 (N_258,In_1368,In_264);
nor U259 (N_259,In_207,In_2073);
nor U260 (N_260,In_812,In_2168);
nor U261 (N_261,In_2332,In_1588);
nor U262 (N_262,In_1752,In_1860);
nand U263 (N_263,In_304,In_2414);
nand U264 (N_264,In_2479,In_2441);
xor U265 (N_265,In_1528,In_1589);
xnor U266 (N_266,In_435,In_1584);
nor U267 (N_267,In_1506,In_1658);
nor U268 (N_268,In_2009,In_1304);
nand U269 (N_269,In_507,In_162);
nor U270 (N_270,In_2466,In_1213);
nor U271 (N_271,In_1331,In_1429);
and U272 (N_272,In_1101,In_758);
nand U273 (N_273,In_669,In_1977);
nand U274 (N_274,In_1638,In_2194);
or U275 (N_275,In_1536,In_1947);
xor U276 (N_276,In_116,In_467);
and U277 (N_277,In_912,In_358);
and U278 (N_278,In_663,In_2336);
nand U279 (N_279,In_1110,In_1695);
nor U280 (N_280,In_1711,In_1173);
and U281 (N_281,In_2240,In_1607);
xnor U282 (N_282,In_1224,In_918);
and U283 (N_283,In_1995,In_867);
or U284 (N_284,In_1160,In_483);
nor U285 (N_285,In_1891,In_148);
or U286 (N_286,In_1978,In_1386);
nand U287 (N_287,In_1475,In_2325);
nand U288 (N_288,In_102,In_794);
or U289 (N_289,In_1587,In_646);
or U290 (N_290,In_1410,In_598);
nor U291 (N_291,In_2489,In_2151);
or U292 (N_292,In_1183,In_1453);
and U293 (N_293,In_252,In_182);
and U294 (N_294,In_846,In_365);
nand U295 (N_295,In_939,In_1850);
or U296 (N_296,In_1943,In_1805);
nand U297 (N_297,In_1785,In_2487);
nor U298 (N_298,In_180,In_2260);
nor U299 (N_299,In_850,In_377);
xor U300 (N_300,In_556,In_951);
xnor U301 (N_301,In_1042,In_261);
nand U302 (N_302,In_2030,In_422);
and U303 (N_303,In_984,In_2421);
or U304 (N_304,In_465,In_1461);
or U305 (N_305,In_415,In_621);
or U306 (N_306,In_1663,In_1019);
or U307 (N_307,In_1426,In_391);
xor U308 (N_308,In_463,In_816);
nand U309 (N_309,In_60,In_1409);
nand U310 (N_310,In_398,In_1164);
and U311 (N_311,In_2385,In_860);
or U312 (N_312,In_549,In_411);
or U313 (N_313,In_2286,In_1060);
or U314 (N_314,In_1152,In_2368);
nand U315 (N_315,In_814,In_2485);
xnor U316 (N_316,In_139,In_1491);
xor U317 (N_317,In_790,In_2424);
nand U318 (N_318,In_2491,In_1312);
nor U319 (N_319,In_567,In_1624);
or U320 (N_320,In_1690,In_1748);
xnor U321 (N_321,In_734,In_90);
xor U322 (N_322,In_1178,In_2090);
or U323 (N_323,In_1551,In_608);
or U324 (N_324,In_2308,In_1480);
or U325 (N_325,In_2124,In_130);
or U326 (N_326,In_1541,In_2103);
nand U327 (N_327,In_929,In_685);
xnor U328 (N_328,In_893,In_123);
and U329 (N_329,In_698,In_1545);
and U330 (N_330,In_993,In_1516);
and U331 (N_331,In_1064,In_830);
xnor U332 (N_332,In_40,In_177);
nand U333 (N_333,In_1870,In_1106);
or U334 (N_334,In_1172,In_1210);
nand U335 (N_335,In_824,In_1875);
nor U336 (N_336,In_1787,In_1017);
xnor U337 (N_337,In_131,In_1415);
and U338 (N_338,In_71,In_2375);
and U339 (N_339,In_470,In_1254);
nand U340 (N_340,In_838,In_440);
nand U341 (N_341,In_1411,In_54);
and U342 (N_342,In_1230,In_717);
nand U343 (N_343,In_1420,In_781);
or U344 (N_344,In_1239,In_836);
or U345 (N_345,In_1863,In_2315);
nor U346 (N_346,In_1611,In_396);
and U347 (N_347,In_2270,In_432);
nand U348 (N_348,In_1999,In_2340);
and U349 (N_349,In_413,In_1299);
nor U350 (N_350,In_2204,In_1313);
or U351 (N_351,In_1195,In_2467);
nand U352 (N_352,In_1825,In_66);
and U353 (N_353,In_688,In_689);
and U354 (N_354,In_444,In_1127);
nor U355 (N_355,In_2221,In_1010);
xor U356 (N_356,In_2038,In_295);
and U357 (N_357,In_1451,In_300);
or U358 (N_358,In_1397,In_1309);
nand U359 (N_359,In_2128,In_921);
and U360 (N_360,In_1543,In_937);
xor U361 (N_361,In_624,In_1757);
or U362 (N_362,In_1396,In_285);
and U363 (N_363,In_575,In_1497);
and U364 (N_364,In_2074,In_728);
nand U365 (N_365,In_426,In_2271);
or U366 (N_366,In_2455,In_1992);
xnor U367 (N_367,In_472,In_2182);
or U368 (N_368,In_948,In_1198);
or U369 (N_369,In_2422,In_2404);
xnor U370 (N_370,In_1071,In_1340);
xnor U371 (N_371,In_1783,In_707);
xor U372 (N_372,In_1513,In_1565);
and U373 (N_373,In_1533,In_213);
or U374 (N_374,In_619,In_2493);
xor U375 (N_375,In_235,In_2200);
and U376 (N_376,In_1980,In_1800);
nor U377 (N_377,In_2253,In_1000);
nor U378 (N_378,In_1496,In_1985);
or U379 (N_379,In_1706,In_2117);
or U380 (N_380,In_1387,In_1770);
xnor U381 (N_381,In_1578,In_1499);
or U382 (N_382,In_569,In_2443);
nor U383 (N_383,In_1688,In_1832);
nand U384 (N_384,In_1417,In_2039);
and U385 (N_385,In_2413,In_2309);
xnor U386 (N_386,In_1855,In_1122);
and U387 (N_387,In_915,In_1956);
nor U388 (N_388,In_220,In_828);
and U389 (N_389,In_1807,In_1692);
xnor U390 (N_390,In_953,In_364);
xor U391 (N_391,In_1689,In_2481);
nor U392 (N_392,In_1946,In_1114);
nor U393 (N_393,In_383,In_712);
xnor U394 (N_394,In_1203,In_2329);
or U395 (N_395,In_2227,In_2069);
nor U396 (N_396,In_686,In_733);
or U397 (N_397,In_651,In_800);
or U398 (N_398,In_101,In_897);
or U399 (N_399,In_1454,In_2028);
or U400 (N_400,In_1432,In_930);
xor U401 (N_401,In_1287,In_979);
nand U402 (N_402,In_852,In_825);
or U403 (N_403,In_2353,In_1581);
or U404 (N_404,In_350,In_1635);
nand U405 (N_405,In_2114,In_2141);
and U406 (N_406,In_1784,In_1872);
xor U407 (N_407,In_1606,In_150);
xor U408 (N_408,In_656,In_1938);
or U409 (N_409,In_421,In_533);
or U410 (N_410,In_745,In_1232);
xnor U411 (N_411,In_1657,In_1046);
nand U412 (N_412,In_700,In_1100);
and U413 (N_413,In_1443,In_360);
or U414 (N_414,In_715,In_2366);
xor U415 (N_415,In_459,In_520);
or U416 (N_416,In_471,In_179);
nor U417 (N_417,In_1402,In_997);
nor U418 (N_418,In_1228,In_2462);
xnor U419 (N_419,In_231,In_28);
xor U420 (N_420,In_936,In_337);
and U421 (N_421,In_205,In_1839);
and U422 (N_422,In_1238,In_505);
nor U423 (N_423,In_1655,In_370);
or U424 (N_424,In_1293,In_528);
xor U425 (N_425,In_2431,In_545);
nor U426 (N_426,In_1518,In_834);
xnor U427 (N_427,In_1758,In_865);
or U428 (N_428,In_1322,In_1816);
nor U429 (N_429,In_1242,In_2469);
xnor U430 (N_430,In_690,In_721);
or U431 (N_431,In_2239,In_1229);
xor U432 (N_432,In_1837,In_74);
and U433 (N_433,In_2006,In_1642);
and U434 (N_434,In_625,In_222);
nor U435 (N_435,In_2077,In_1145);
nand U436 (N_436,In_1935,In_1933);
xor U437 (N_437,In_420,In_332);
xnor U438 (N_438,In_412,In_7);
nand U439 (N_439,In_2454,In_596);
nor U440 (N_440,In_2085,In_1274);
nand U441 (N_441,In_118,In_2459);
or U442 (N_442,In_1323,In_2082);
and U443 (N_443,In_1133,In_704);
or U444 (N_444,In_779,In_777);
or U445 (N_445,In_956,In_1931);
and U446 (N_446,In_1421,In_552);
xor U447 (N_447,In_582,In_488);
or U448 (N_448,In_1954,In_26);
nor U449 (N_449,In_286,In_1519);
and U450 (N_450,In_684,In_1231);
or U451 (N_451,In_874,In_2245);
or U452 (N_452,In_943,In_2054);
xnor U453 (N_453,In_1253,In_302);
or U454 (N_454,In_379,In_492);
or U455 (N_455,In_2287,In_693);
nor U456 (N_456,In_2183,In_2035);
and U457 (N_457,In_1315,In_534);
nor U458 (N_458,In_641,In_2165);
xor U459 (N_459,In_12,In_97);
and U460 (N_460,In_1216,In_1081);
nor U461 (N_461,In_2116,In_2473);
xnor U462 (N_462,In_1219,In_966);
nand U463 (N_463,In_1896,In_2386);
xor U464 (N_464,In_1720,In_1592);
xnor U465 (N_465,In_1117,In_341);
nor U466 (N_466,In_530,In_324);
or U467 (N_467,In_479,In_1177);
and U468 (N_468,In_1026,In_976);
nand U469 (N_469,In_1779,In_697);
xor U470 (N_470,In_1803,In_19);
nor U471 (N_471,In_954,In_1161);
and U472 (N_472,In_1656,In_563);
nor U473 (N_473,In_1646,In_1031);
nand U474 (N_474,In_1557,In_1422);
xnor U475 (N_475,In_25,In_831);
and U476 (N_476,In_1570,In_623);
nand U477 (N_477,In_186,In_2312);
and U478 (N_478,In_1547,In_278);
nor U479 (N_479,In_111,In_1702);
nor U480 (N_480,In_1694,In_2344);
nand U481 (N_481,In_1653,In_888);
xnor U482 (N_482,In_769,In_2179);
and U483 (N_483,In_1032,In_2324);
nand U484 (N_484,In_95,In_1234);
nand U485 (N_485,In_1553,In_903);
nand U486 (N_486,In_2415,In_2378);
and U487 (N_487,In_2439,In_160);
or U488 (N_488,In_145,In_2046);
or U489 (N_489,In_2371,In_2161);
xor U490 (N_490,In_1072,In_1605);
xnor U491 (N_491,In_599,In_218);
and U492 (N_492,In_120,In_622);
xor U493 (N_493,In_1393,In_1137);
xnor U494 (N_494,In_168,In_1166);
or U495 (N_495,In_631,In_51);
nand U496 (N_496,In_37,In_1979);
or U497 (N_497,In_223,In_2057);
nor U498 (N_498,In_2041,In_1199);
xor U499 (N_499,In_1705,In_1701);
or U500 (N_500,In_147,In_2307);
nor U501 (N_501,In_1602,In_1673);
or U502 (N_502,In_1955,In_2338);
xor U503 (N_503,In_1733,In_861);
xor U504 (N_504,In_198,In_1794);
xor U505 (N_505,In_1362,In_209);
and U506 (N_506,In_2044,In_2468);
or U507 (N_507,In_1140,In_1301);
and U508 (N_508,In_2217,In_219);
and U509 (N_509,In_242,In_885);
and U510 (N_510,In_637,In_603);
nor U511 (N_511,In_1824,In_1868);
or U512 (N_512,In_216,In_91);
or U513 (N_513,In_1361,In_2465);
or U514 (N_514,In_482,In_2205);
xor U515 (N_515,In_1381,In_1268);
xor U516 (N_516,In_1053,In_2195);
and U517 (N_517,In_1465,In_952);
nand U518 (N_518,In_1460,In_1679);
nand U519 (N_519,In_927,In_1385);
nor U520 (N_520,In_32,In_676);
nor U521 (N_521,In_1405,In_2495);
xnor U522 (N_522,In_2250,In_388);
nor U523 (N_523,In_2208,In_2478);
nand U524 (N_524,In_2015,In_1206);
nand U525 (N_525,In_2362,In_601);
and U526 (N_526,In_506,In_2111);
nor U527 (N_527,In_8,In_919);
nor U528 (N_528,In_2427,In_1926);
nor U529 (N_529,In_1418,In_2197);
nand U530 (N_530,In_1485,In_796);
or U531 (N_531,In_1037,In_1352);
nor U532 (N_532,In_1365,In_538);
or U533 (N_533,In_590,In_307);
and U534 (N_534,In_2408,In_615);
and U535 (N_535,In_701,In_977);
or U536 (N_536,In_772,In_1221);
nor U537 (N_537,In_171,In_508);
nand U538 (N_538,In_331,In_361);
or U539 (N_539,In_2231,In_68);
nand U540 (N_540,In_1306,In_2321);
xnor U541 (N_541,In_86,In_2377);
xor U542 (N_542,In_983,In_1459);
and U543 (N_543,In_980,In_1382);
xnor U544 (N_544,In_1904,In_2096);
nor U545 (N_545,In_1065,In_2010);
xnor U546 (N_546,In_965,In_907);
or U547 (N_547,In_1257,In_1383);
nand U548 (N_548,In_2,In_1444);
nand U549 (N_549,In_1847,In_835);
or U550 (N_550,In_448,In_1094);
xor U551 (N_551,In_1906,In_667);
or U552 (N_552,In_1476,In_1237);
or U553 (N_553,In_940,In_325);
nand U554 (N_554,In_1038,In_1580);
or U555 (N_555,In_1059,In_2437);
or U556 (N_556,In_2456,In_2262);
nand U557 (N_557,In_1665,In_317);
nor U558 (N_558,In_868,In_155);
nand U559 (N_559,In_36,In_1082);
nand U560 (N_560,In_2490,In_762);
nand U561 (N_561,In_949,In_2159);
nand U562 (N_562,In_616,In_210);
xor U563 (N_563,In_1018,In_2292);
and U564 (N_564,In_2438,In_2018);
nand U565 (N_565,In_30,In_679);
nor U566 (N_566,In_1334,In_2137);
or U567 (N_567,In_1077,In_2174);
or U568 (N_568,In_1795,In_1358);
and U569 (N_569,In_122,In_1808);
nand U570 (N_570,In_367,In_1132);
nand U571 (N_571,In_416,In_2367);
nand U572 (N_572,In_1165,In_577);
nand U573 (N_573,In_297,In_1736);
nand U574 (N_574,In_2403,In_1903);
and U575 (N_575,In_2196,In_1554);
and U576 (N_576,In_536,In_2107);
and U577 (N_577,In_938,In_1414);
xor U578 (N_578,In_466,In_271);
nor U579 (N_579,In_339,In_917);
nor U580 (N_580,In_170,In_1835);
or U581 (N_581,In_485,In_2381);
and U582 (N_582,In_228,In_2395);
or U583 (N_583,In_2322,In_1084);
and U584 (N_584,In_780,In_967);
nand U585 (N_585,In_1672,In_1067);
or U586 (N_586,In_43,In_958);
or U587 (N_587,In_1424,In_2154);
nor U588 (N_588,In_570,In_390);
nand U589 (N_589,In_1509,In_1698);
nor U590 (N_590,In_691,In_1894);
xnor U591 (N_591,In_208,In_1831);
or U592 (N_592,In_1351,In_374);
nor U593 (N_593,In_1780,In_571);
nor U594 (N_594,In_1744,In_591);
xnor U595 (N_595,In_2343,In_988);
or U596 (N_596,In_1416,In_833);
or U597 (N_597,In_2301,In_250);
or U598 (N_598,In_821,In_2060);
nor U599 (N_599,In_673,In_1774);
or U600 (N_600,In_2110,In_1305);
and U601 (N_601,In_1503,In_773);
and U602 (N_602,In_1156,In_100);
xnor U603 (N_603,In_1376,In_2379);
or U604 (N_604,In_957,In_469);
and U605 (N_605,In_313,In_1934);
and U606 (N_606,In_1969,In_1817);
and U607 (N_607,In_2184,In_211);
nor U608 (N_608,In_1912,In_2255);
or U609 (N_609,In_1960,In_433);
nor U610 (N_610,In_687,In_1006);
xnor U611 (N_611,In_2345,In_1627);
xor U612 (N_612,In_2442,In_2382);
or U613 (N_613,In_484,In_996);
xor U614 (N_614,In_1186,In_737);
xor U615 (N_615,In_776,In_326);
nor U616 (N_616,In_950,In_1149);
or U617 (N_617,In_136,In_1871);
xnor U618 (N_618,In_826,In_225);
or U619 (N_619,In_1913,In_2460);
nor U620 (N_620,In_1975,In_329);
nor U621 (N_621,In_2498,In_1667);
nor U622 (N_622,In_632,In_1707);
nand U623 (N_623,In_692,In_654);
or U624 (N_624,In_2113,In_2430);
and U625 (N_625,In_1247,In_525);
or U626 (N_626,In_1016,In_1494);
nor U627 (N_627,In_1375,In_2463);
xor U628 (N_628,In_292,In_475);
nor U629 (N_629,In_203,In_1964);
or U630 (N_630,In_0,In_237);
or U631 (N_631,In_1648,In_845);
or U632 (N_632,In_1829,In_2072);
nor U633 (N_633,In_1811,In_24);
nor U634 (N_634,In_2475,In_2086);
or U635 (N_635,In_898,In_760);
or U636 (N_636,In_489,In_1045);
nor U637 (N_637,In_1511,In_2264);
nor U638 (N_638,In_1123,In_135);
or U639 (N_639,In_138,In_1462);
or U640 (N_640,In_2294,In_1996);
nand U641 (N_641,In_392,In_1079);
xor U642 (N_642,In_1737,In_890);
or U643 (N_643,In_2234,In_455);
nand U644 (N_644,In_748,In_736);
xor U645 (N_645,In_1005,In_2032);
or U646 (N_646,In_1590,In_2298);
or U647 (N_647,In_1967,In_495);
nor U648 (N_648,In_1144,In_2023);
xor U649 (N_649,In_1236,In_2356);
nand U650 (N_650,In_2150,In_348);
and U651 (N_651,In_875,In_1294);
nand U652 (N_652,In_1563,In_2120);
nand U653 (N_653,In_604,In_778);
and U654 (N_654,In_2360,In_1262);
xor U655 (N_655,In_110,In_1290);
nor U656 (N_656,In_153,In_2140);
nand U657 (N_657,In_827,In_1175);
and U658 (N_658,In_660,In_234);
xor U659 (N_659,In_843,In_1827);
or U660 (N_660,In_869,In_539);
xnor U661 (N_661,In_524,In_1771);
or U662 (N_662,In_1527,In_789);
or U663 (N_663,In_2143,In_1360);
or U664 (N_664,In_2118,In_1877);
nor U665 (N_665,In_239,In_1034);
nand U666 (N_666,In_2440,In_1277);
nor U667 (N_667,In_2145,In_2132);
nand U668 (N_668,In_1051,In_1820);
and U669 (N_669,In_1473,In_2102);
nand U670 (N_670,In_1609,In_1788);
xor U671 (N_671,In_2093,In_2313);
or U672 (N_672,In_2051,In_763);
xor U673 (N_673,In_1687,In_133);
and U674 (N_674,In_1631,In_2088);
nor U675 (N_675,In_747,In_785);
nor U676 (N_676,In_1478,In_1806);
nand U677 (N_677,In_336,In_1028);
and U678 (N_678,In_1279,In_1900);
nor U679 (N_679,In_1180,In_522);
or U680 (N_680,In_254,In_2235);
and U681 (N_681,In_1335,In_630);
or U682 (N_682,In_1074,In_1438);
xnor U683 (N_683,In_2203,In_894);
and U684 (N_684,In_2486,In_1898);
and U685 (N_685,In_46,In_268);
and U686 (N_686,In_1022,In_595);
or U687 (N_687,In_922,In_146);
xnor U688 (N_688,In_643,In_2226);
nand U689 (N_689,In_320,In_277);
nor U690 (N_690,In_1318,In_1621);
nand U691 (N_691,In_389,In_80);
and U692 (N_692,In_730,In_2449);
and U693 (N_693,In_1090,In_541);
xnor U694 (N_694,In_94,In_275);
and U695 (N_695,In_1989,In_1994);
nand U696 (N_696,In_431,In_706);
nor U697 (N_697,In_1828,In_1111);
and U698 (N_698,In_1338,In_1367);
and U699 (N_699,In_134,In_1350);
nor U700 (N_700,In_2230,In_2470);
xor U701 (N_701,In_866,In_1696);
nand U702 (N_702,In_1537,In_1972);
or U703 (N_703,In_1021,In_1412);
or U704 (N_704,In_1899,In_92);
and U705 (N_705,In_514,In_2402);
nand U706 (N_706,In_1715,In_711);
nor U707 (N_707,In_1991,In_1856);
and U708 (N_708,In_276,In_1854);
and U709 (N_709,In_1645,In_873);
xor U710 (N_710,In_2066,In_2104);
xor U711 (N_711,In_2337,In_20);
xnor U712 (N_712,In_1940,In_1251);
or U713 (N_713,In_584,In_1599);
xnor U714 (N_714,In_618,In_724);
nor U715 (N_715,In_2259,In_1713);
and U716 (N_716,In_1025,In_2158);
xnor U717 (N_717,In_862,In_480);
xnor U718 (N_718,In_2199,In_322);
nor U719 (N_719,In_1141,In_2254);
nor U720 (N_720,In_1483,In_638);
nand U721 (N_721,In_1029,In_2115);
xor U722 (N_722,In_588,In_1271);
nor U723 (N_723,In_2075,In_1115);
xor U724 (N_724,In_108,In_1289);
or U725 (N_725,In_310,In_34);
and U726 (N_726,In_2002,In_308);
nand U727 (N_727,In_2218,In_1288);
and U728 (N_728,In_1470,In_947);
and U729 (N_729,In_2444,In_1388);
nor U730 (N_730,In_1431,In_974);
xnor U731 (N_731,In_1468,In_1743);
xor U732 (N_732,In_83,In_1248);
and U733 (N_733,In_1573,In_1525);
or U734 (N_734,In_192,In_1735);
nor U735 (N_735,In_202,In_1500);
xnor U736 (N_736,In_369,In_387);
xnor U737 (N_737,In_1612,In_45);
xnor U738 (N_738,In_1275,In_1762);
nand U739 (N_739,In_882,In_452);
or U740 (N_740,In_981,In_2428);
and U741 (N_741,In_911,In_1834);
xnor U742 (N_742,In_1098,In_338);
xor U743 (N_743,In_2193,In_474);
and U744 (N_744,In_270,In_31);
nand U745 (N_745,In_2372,In_294);
xor U746 (N_746,In_1014,In_1830);
nor U747 (N_747,In_400,In_1486);
nand U748 (N_748,In_2056,In_1490);
nand U749 (N_749,In_434,In_481);
nor U750 (N_750,In_1227,In_1628);
xnor U751 (N_751,In_1790,In_248);
and U752 (N_752,In_42,In_340);
nor U753 (N_753,In_427,In_558);
xnor U754 (N_754,In_2306,In_1942);
nand U755 (N_755,In_1914,In_499);
nor U756 (N_756,In_458,In_2187);
or U757 (N_757,In_652,In_718);
nand U758 (N_758,In_2186,In_515);
nor U759 (N_759,In_1524,In_164);
or U760 (N_760,In_2464,In_2327);
or U761 (N_761,In_750,In_1945);
and U762 (N_762,In_786,In_1529);
or U763 (N_763,In_334,In_93);
nand U764 (N_764,In_2062,In_817);
and U765 (N_765,In_312,In_1049);
nor U766 (N_766,In_675,In_837);
and U767 (N_767,In_1759,In_363);
or U768 (N_768,In_1040,In_2063);
and U769 (N_769,In_35,In_503);
nand U770 (N_770,In_1364,In_738);
nand U771 (N_771,In_2290,In_535);
nor U772 (N_772,In_574,In_1867);
or U773 (N_773,In_229,In_206);
nor U774 (N_774,In_2348,In_548);
and U775 (N_775,In_1324,In_290);
nor U776 (N_776,In_129,In_1447);
nand U777 (N_777,In_2136,In_126);
nand U778 (N_778,In_281,In_832);
and U779 (N_779,In_1603,In_2164);
xor U780 (N_780,In_1674,In_409);
xor U781 (N_781,In_2447,In_999);
nor U782 (N_782,In_496,In_813);
nand U783 (N_783,In_1789,In_425);
or U784 (N_784,In_172,In_934);
xor U785 (N_785,In_1437,In_1282);
or U786 (N_786,In_2296,In_910);
xnor U787 (N_787,In_2279,In_2278);
nor U788 (N_788,In_1902,In_1895);
and U789 (N_789,In_746,In_1250);
xor U790 (N_790,In_305,In_1893);
nand U791 (N_791,In_1311,In_2177);
and U792 (N_792,In_2207,In_253);
xnor U793 (N_793,In_2225,In_732);
nand U794 (N_794,In_185,In_2100);
and U795 (N_795,In_605,In_314);
xnor U796 (N_796,In_1846,In_2139);
or U797 (N_797,In_1204,In_1548);
or U798 (N_798,In_10,In_1766);
or U799 (N_799,In_1096,In_2432);
xnor U800 (N_800,In_655,In_753);
xnor U801 (N_801,In_1997,In_1502);
nand U802 (N_802,In_1729,In_743);
nand U803 (N_803,In_1099,In_354);
xor U804 (N_804,In_2284,In_1083);
and U805 (N_805,In_2223,In_2241);
nor U806 (N_806,In_1718,In_580);
and U807 (N_807,In_1819,In_1728);
or U808 (N_808,In_1613,In_2011);
nor U809 (N_809,In_592,In_487);
and U810 (N_810,In_2273,In_247);
nor U811 (N_811,In_152,In_140);
nand U812 (N_812,In_945,In_344);
and U813 (N_813,In_113,In_1801);
and U814 (N_814,In_9,In_406);
and U815 (N_815,In_414,In_2429);
nor U816 (N_816,In_1550,In_1595);
nand U817 (N_817,In_1764,In_1739);
nand U818 (N_818,In_1374,In_2138);
and U819 (N_819,In_1911,In_2157);
nand U820 (N_820,In_502,In_1333);
nor U821 (N_821,In_774,In_1357);
and U822 (N_822,In_53,In_1574);
nand U823 (N_823,In_47,In_1844);
or U824 (N_824,In_620,In_2400);
xor U825 (N_825,In_178,In_1092);
nor U826 (N_826,In_1104,In_2215);
or U827 (N_827,In_1952,In_1243);
xor U828 (N_828,In_856,In_2188);
or U829 (N_829,In_2081,In_1833);
xnor U830 (N_830,In_1245,In_1463);
or U831 (N_831,In_1310,In_1148);
xnor U832 (N_832,In_1916,In_1191);
nor U833 (N_833,In_17,In_2122);
nor U834 (N_834,In_44,In_73);
xor U835 (N_835,In_2142,In_1190);
nor U836 (N_836,In_2243,In_1660);
and U837 (N_837,In_2198,In_1874);
xor U838 (N_838,In_1220,In_382);
and U839 (N_839,In_1910,In_1927);
xnor U840 (N_840,In_2007,In_2411);
nand U841 (N_841,In_1616,In_2494);
nor U842 (N_842,In_96,In_2152);
xnor U843 (N_843,In_1556,In_1719);
or U844 (N_844,In_1731,In_1472);
or U845 (N_845,In_287,In_2388);
nand U846 (N_846,In_761,In_719);
xor U847 (N_847,In_2206,In_1708);
nand U848 (N_848,In_1984,In_196);
nor U849 (N_849,In_1023,In_2359);
nand U850 (N_850,In_1741,In_442);
xor U851 (N_851,In_169,In_2000);
nand U852 (N_852,In_137,In_2026);
nor U853 (N_853,In_982,In_2266);
nand U854 (N_854,In_2472,In_1661);
xor U855 (N_855,In_2248,In_607);
or U856 (N_856,In_1949,In_289);
xor U857 (N_857,In_810,In_909);
xor U858 (N_858,In_16,In_2005);
xor U859 (N_859,In_1169,In_802);
nor U860 (N_860,In_88,In_166);
nor U861 (N_861,In_75,In_65);
nor U862 (N_862,In_2450,In_447);
nand U863 (N_863,In_2058,In_1380);
or U864 (N_864,In_490,In_2448);
or U865 (N_865,In_79,In_1650);
nand U866 (N_866,In_280,In_881);
and U867 (N_867,In_1121,In_1962);
and U868 (N_868,In_265,In_783);
or U869 (N_869,In_1066,In_2037);
nor U870 (N_870,In_429,In_1153);
or U871 (N_871,In_989,In_1225);
and U872 (N_872,In_904,In_1212);
and U873 (N_873,In_1601,In_1035);
nand U874 (N_874,In_1866,In_990);
nand U875 (N_875,In_2412,In_176);
nor U876 (N_876,In_359,In_319);
or U877 (N_877,In_1076,In_1330);
or U878 (N_878,In_1366,In_1973);
xnor U879 (N_879,In_445,In_2396);
or U880 (N_880,In_884,In_740);
or U881 (N_881,In_2380,In_923);
nor U882 (N_882,In_578,In_1427);
xnor U883 (N_883,In_851,In_550);
nor U884 (N_884,In_2282,In_33);
or U885 (N_885,In_2311,In_1542);
nand U886 (N_886,In_757,In_491);
xor U887 (N_887,In_1865,In_2257);
or U888 (N_888,In_1843,In_49);
nor U889 (N_889,In_1217,In_132);
nor U890 (N_890,In_2095,In_1174);
nor U891 (N_891,In_1723,In_2091);
xnor U892 (N_892,In_2236,In_1745);
xnor U893 (N_893,In_1116,In_1971);
xor U894 (N_894,In_1093,In_509);
and U895 (N_895,In_665,In_2222);
xor U896 (N_896,In_579,In_1939);
nand U897 (N_897,In_1925,In_349);
nor U898 (N_898,In_870,In_529);
nor U899 (N_899,In_1591,In_173);
nor U900 (N_900,In_787,In_2209);
nor U901 (N_901,In_215,In_1407);
xnor U902 (N_902,In_236,In_2065);
and U903 (N_903,In_18,In_1928);
or U904 (N_904,In_1721,In_2049);
or U905 (N_905,In_994,In_1013);
xnor U906 (N_906,In_1080,In_1765);
nor U907 (N_907,In_151,In_1134);
or U908 (N_908,In_547,In_609);
xnor U909 (N_909,In_857,In_1530);
nor U910 (N_910,In_15,In_397);
xnor U911 (N_911,In_1226,In_446);
nor U912 (N_912,In_1561,In_699);
nor U913 (N_913,In_1957,In_62);
and U914 (N_914,In_1062,In_735);
nor U915 (N_915,In_512,In_183);
nand U916 (N_916,In_59,In_749);
xor U917 (N_917,In_306,In_11);
or U918 (N_918,In_193,In_1107);
nor U919 (N_919,In_55,In_797);
nor U920 (N_920,In_1958,In_1892);
nand U921 (N_921,In_1208,In_1768);
and U922 (N_922,In_2126,In_916);
nand U923 (N_923,In_1456,In_589);
or U924 (N_924,In_2024,In_1307);
nor U925 (N_925,In_2291,In_144);
or U926 (N_926,In_1185,In_408);
nand U927 (N_927,In_1223,In_163);
xor U928 (N_928,In_878,In_1436);
and U929 (N_929,In_2016,In_1885);
nand U930 (N_930,In_441,In_321);
nor U931 (N_931,In_931,In_187);
nor U932 (N_932,In_1691,In_2068);
or U933 (N_933,In_649,In_1314);
or U934 (N_934,In_1052,In_941);
nand U935 (N_935,In_1484,In_798);
or U936 (N_936,In_628,In_1085);
or U937 (N_937,In_801,In_516);
nand U938 (N_938,In_1403,In_315);
nor U939 (N_939,In_611,In_1408);
nor U940 (N_940,In_928,In_1222);
xnor U941 (N_941,In_1265,In_806);
and U942 (N_942,In_1841,In_1344);
and U943 (N_943,In_1767,In_2146);
nand U944 (N_944,In_1404,In_1073);
and U945 (N_945,In_378,In_1950);
nand U946 (N_946,In_399,In_76);
nand U947 (N_947,In_504,In_1039);
or U948 (N_948,In_1747,In_2185);
or U949 (N_949,In_21,In_2458);
nand U950 (N_950,In_1088,In_2285);
nor U951 (N_951,In_2434,In_1346);
xor U952 (N_952,In_767,In_1918);
nand U953 (N_953,In_2099,In_1036);
nand U954 (N_954,In_201,In_403);
nor U955 (N_955,In_1298,In_2052);
and U956 (N_956,In_1990,In_770);
nand U957 (N_957,In_844,In_2210);
xnor U958 (N_958,In_1781,In_2121);
and U959 (N_959,In_1640,In_2355);
nand U960 (N_960,In_127,In_2384);
or U961 (N_961,In_1302,In_883);
nand U962 (N_962,In_486,In_1024);
nor U963 (N_963,In_859,In_1922);
xor U964 (N_964,In_462,In_2048);
or U965 (N_965,In_1923,In_1849);
xnor U966 (N_966,In_371,In_1112);
nor U967 (N_967,In_752,In_2341);
xor U968 (N_968,In_1684,In_955);
nand U969 (N_969,In_1753,In_1295);
and U970 (N_970,In_2299,In_1069);
and U971 (N_971,In_2330,In_1151);
xnor U972 (N_972,In_293,In_1791);
xor U973 (N_973,In_561,In_1755);
nor U974 (N_974,In_1457,In_1639);
xnor U975 (N_975,In_2125,In_1292);
and U976 (N_976,In_1348,In_2173);
xnor U977 (N_977,In_1730,In_2354);
nor U978 (N_978,In_1428,In_1738);
nor U979 (N_979,In_1189,In_57);
nand U980 (N_980,In_782,In_1128);
xor U981 (N_981,In_1775,In_1681);
nand U982 (N_982,In_1579,In_1063);
nor U983 (N_983,In_1637,In_1786);
nor U984 (N_984,In_1568,In_1818);
and U985 (N_985,In_2499,In_1704);
nor U986 (N_986,In_1197,In_2258);
nor U987 (N_987,In_386,In_2020);
nand U988 (N_988,In_204,In_1391);
nor U989 (N_989,In_2417,In_674);
and U990 (N_990,In_2216,In_975);
nand U991 (N_991,In_2497,In_124);
or U992 (N_992,In_1371,In_1987);
nor U993 (N_993,In_282,In_1332);
nand U994 (N_994,In_2178,In_104);
xor U995 (N_995,In_2172,In_1881);
or U996 (N_996,In_1598,In_1054);
and U997 (N_997,In_50,In_1433);
xnor U998 (N_998,In_1398,In_1209);
or U999 (N_999,In_1466,In_657);
or U1000 (N_1000,In_190,In_583);
nor U1001 (N_1001,In_1716,In_1252);
or U1002 (N_1002,In_266,In_1280);
xnor U1003 (N_1003,In_793,In_2084);
xor U1004 (N_1004,In_1944,In_1055);
or U1005 (N_1005,In_283,In_1201);
nand U1006 (N_1006,In_1261,In_1015);
and U1007 (N_1007,In_682,In_1143);
and U1008 (N_1008,In_121,In_1608);
and U1009 (N_1009,In_2420,In_2144);
xor U1010 (N_1010,In_1218,In_112);
nor U1011 (N_1011,In_1932,In_963);
xor U1012 (N_1012,In_99,In_2374);
nand U1013 (N_1013,In_1394,In_106);
nor U1014 (N_1014,In_2190,In_755);
nand U1015 (N_1015,In_1384,In_1009);
nand U1016 (N_1016,In_744,In_771);
or U1017 (N_1017,In_1564,In_1103);
nand U1018 (N_1018,In_1392,In_670);
and U1019 (N_1019,In_593,In_298);
nand U1020 (N_1020,In_1181,In_1620);
nand U1021 (N_1021,In_174,In_1285);
or U1022 (N_1022,In_942,In_417);
xor U1023 (N_1023,In_1625,In_1297);
or U1024 (N_1024,In_404,In_1372);
or U1025 (N_1025,In_1378,In_1163);
xor U1026 (N_1026,In_1862,In_1097);
nand U1027 (N_1027,In_1905,In_2001);
and U1028 (N_1028,In_1267,In_1948);
nand U1029 (N_1029,In_1263,In_2025);
nand U1030 (N_1030,In_1102,In_2019);
nor U1031 (N_1031,In_775,In_1864);
nand U1032 (N_1032,In_1534,In_647);
nand U1033 (N_1033,In_1915,In_2127);
xnor U1034 (N_1034,In_2320,In_2256);
or U1035 (N_1035,In_1130,In_998);
or U1036 (N_1036,In_2267,In_968);
nor U1037 (N_1037,In_2293,In_381);
xnor U1038 (N_1038,In_2171,In_2167);
or U1039 (N_1039,In_537,In_288);
nand U1040 (N_1040,In_67,In_1558);
nand U1041 (N_1041,In_2476,In_453);
or U1042 (N_1042,In_52,In_214);
xnor U1043 (N_1043,In_1441,In_1316);
and U1044 (N_1044,In_634,In_2021);
nand U1045 (N_1045,In_2148,In_962);
nor U1046 (N_1046,In_2272,In_159);
nor U1047 (N_1047,In_2305,In_1155);
or U1048 (N_1048,In_879,In_2387);
nor U1049 (N_1049,In_1676,In_1717);
nor U1050 (N_1050,In_449,In_1643);
nor U1051 (N_1051,In_901,In_1027);
or U1052 (N_1052,In_1041,In_1435);
and U1053 (N_1053,In_373,In_2281);
nand U1054 (N_1054,In_710,In_385);
or U1055 (N_1055,In_1769,In_423);
xnor U1056 (N_1056,In_1897,In_564);
nor U1057 (N_1057,In_1670,In_2229);
nor U1058 (N_1058,In_2369,In_2453);
xnor U1059 (N_1059,In_1356,In_1501);
or U1060 (N_1060,In_2131,In_895);
nand U1061 (N_1061,In_1576,In_1517);
or U1062 (N_1062,In_2265,In_184);
nand U1063 (N_1063,In_1930,In_384);
or U1064 (N_1064,In_245,In_84);
xor U1065 (N_1065,In_2339,In_2083);
xnor U1066 (N_1066,In_891,In_766);
nor U1067 (N_1067,In_39,In_1583);
or U1068 (N_1068,In_77,In_2013);
nand U1069 (N_1069,In_933,In_557);
xnor U1070 (N_1070,In_1878,In_1859);
and U1071 (N_1071,In_985,In_880);
or U1072 (N_1072,In_1535,In_666);
nor U1073 (N_1073,In_1050,In_2364);
nand U1074 (N_1074,In_705,In_517);
nand U1075 (N_1075,In_436,In_1734);
nand U1076 (N_1076,In_1434,In_2426);
or U1077 (N_1077,In_1147,In_1001);
nor U1078 (N_1078,In_1618,In_1559);
and U1079 (N_1079,In_1634,In_1838);
or U1080 (N_1080,In_2335,In_1540);
or U1081 (N_1081,In_1487,In_2202);
nor U1082 (N_1082,In_1654,In_1154);
nor U1083 (N_1083,In_853,In_1982);
or U1084 (N_1084,In_889,In_284);
nand U1085 (N_1085,In_809,In_815);
and U1086 (N_1086,In_1202,In_727);
or U1087 (N_1087,In_82,In_1142);
nand U1088 (N_1088,In_1544,In_3);
nand U1089 (N_1089,In_1710,In_188);
xnor U1090 (N_1090,In_1998,In_702);
xnor U1091 (N_1091,In_1504,In_2346);
or U1092 (N_1092,In_2373,In_1445);
nor U1093 (N_1093,In_759,In_1802);
nand U1094 (N_1094,In_2249,In_1714);
and U1095 (N_1095,In_1187,In_1390);
and U1096 (N_1096,In_2219,In_672);
and U1097 (N_1097,In_1776,In_115);
nand U1098 (N_1098,In_876,In_1569);
and U1099 (N_1099,In_2347,In_2357);
xor U1100 (N_1100,In_1129,In_678);
xnor U1101 (N_1101,In_2181,In_128);
nand U1102 (N_1102,In_2036,In_143);
or U1103 (N_1103,In_2409,In_613);
and U1104 (N_1104,In_978,In_1283);
nand U1105 (N_1105,In_2135,In_195);
or U1106 (N_1106,In_1882,In_1822);
or U1107 (N_1107,In_2492,In_328);
nor U1108 (N_1108,In_1479,In_194);
nor U1109 (N_1109,In_1886,In_1193);
nor U1110 (N_1110,In_22,In_532);
nor U1111 (N_1111,In_1321,In_2407);
and U1112 (N_1112,In_501,In_527);
nand U1113 (N_1113,In_362,In_519);
or U1114 (N_1114,In_765,In_2393);
nor U1115 (N_1115,In_393,In_2012);
nor U1116 (N_1116,In_1281,In_696);
nor U1117 (N_1117,In_1614,In_683);
nand U1118 (N_1118,In_612,In_602);
nor U1119 (N_1119,In_581,In_1255);
nand U1120 (N_1120,In_1703,In_1233);
nor U1121 (N_1121,In_1675,In_1641);
xor U1122 (N_1122,In_1349,In_754);
and U1123 (N_1123,In_157,In_424);
or U1124 (N_1124,In_1162,In_2263);
or U1125 (N_1125,In_768,In_2326);
xor U1126 (N_1126,In_70,In_2053);
nor U1127 (N_1127,In_1521,In_2133);
nor U1128 (N_1128,In_2166,In_1659);
nor U1129 (N_1129,In_2405,In_566);
nand U1130 (N_1130,In_1258,In_1937);
nor U1131 (N_1131,In_1168,In_1105);
nor U1132 (N_1132,In_1615,In_1677);
nand U1133 (N_1133,In_335,In_1355);
nor U1134 (N_1134,In_2022,In_2043);
nand U1135 (N_1135,In_920,In_356);
xnor U1136 (N_1136,In_1809,In_1146);
nand U1137 (N_1137,In_497,In_716);
and U1138 (N_1138,In_1531,In_1908);
nand U1139 (N_1139,In_633,In_1259);
nand U1140 (N_1140,In_468,In_1636);
nor U1141 (N_1141,In_41,In_731);
xnor U1142 (N_1142,In_4,In_2109);
or U1143 (N_1143,In_1988,In_1464);
or U1144 (N_1144,In_1575,In_1300);
and U1145 (N_1145,In_1341,In_1167);
nor U1146 (N_1146,In_565,In_2477);
xor U1147 (N_1147,In_1507,In_1560);
nand U1148 (N_1148,In_741,In_2445);
nor U1149 (N_1149,In_2488,In_1319);
nor U1150 (N_1150,In_2323,In_546);
and U1151 (N_1151,In_1549,In_2130);
xor U1152 (N_1152,In_1044,In_1047);
or U1153 (N_1153,In_1668,In_2365);
nor U1154 (N_1154,In_2342,In_375);
nand U1155 (N_1155,In_662,In_439);
xor U1156 (N_1156,In_722,In_1359);
and U1157 (N_1157,In_2089,In_69);
nor U1158 (N_1158,In_267,In_1812);
xor U1159 (N_1159,In_1395,In_199);
nor U1160 (N_1160,In_405,In_1449);
xnor U1161 (N_1161,In_142,In_2391);
nand U1162 (N_1162,In_629,In_249);
and U1163 (N_1163,In_839,In_1370);
or U1164 (N_1164,In_1852,In_2191);
nand U1165 (N_1165,In_29,In_523);
nand U1166 (N_1166,In_64,In_792);
xor U1167 (N_1167,In_1086,In_987);
or U1168 (N_1168,In_158,In_803);
nor U1169 (N_1169,In_1778,In_543);
xor U1170 (N_1170,In_1296,In_1419);
xnor U1171 (N_1171,In_636,In_1840);
xor U1172 (N_1172,In_2401,In_1481);
and U1173 (N_1173,In_2189,In_642);
xor U1174 (N_1174,In_2471,In_1974);
nor U1175 (N_1175,In_864,In_2389);
xor U1176 (N_1176,In_2050,In_1917);
nor U1177 (N_1177,In_175,In_872);
and U1178 (N_1178,In_1617,In_1347);
xnor U1179 (N_1179,In_1523,In_141);
xnor U1180 (N_1180,In_1264,In_2201);
nand U1181 (N_1181,In_899,In_863);
nor U1182 (N_1182,In_1379,In_2425);
or U1183 (N_1183,In_1604,In_1345);
or U1184 (N_1184,In_1907,In_2398);
and U1185 (N_1185,In_1869,In_1546);
xor U1186 (N_1186,In_330,In_551);
nor U1187 (N_1187,In_450,In_1336);
or U1188 (N_1188,In_2334,In_2390);
and U1189 (N_1189,In_1773,In_513);
and U1190 (N_1190,In_1669,In_2289);
xnor U1191 (N_1191,In_1749,In_1150);
xnor U1192 (N_1192,In_1700,In_1273);
xnor U1193 (N_1193,In_1929,In_346);
nor U1194 (N_1194,In_1327,In_847);
nand U1195 (N_1195,In_2031,In_61);
and U1196 (N_1196,In_1,In_645);
xnor U1197 (N_1197,In_1814,In_343);
nand U1198 (N_1198,In_2363,In_1284);
nor U1199 (N_1199,In_946,In_2349);
nor U1200 (N_1200,In_627,In_695);
nor U1201 (N_1201,In_419,In_1686);
nor U1202 (N_1202,In_2480,In_1048);
xnor U1203 (N_1203,In_587,In_964);
and U1204 (N_1204,In_1109,In_2244);
nor U1205 (N_1205,In_105,In_1632);
nor U1206 (N_1206,In_394,In_559);
or U1207 (N_1207,In_823,In_2484);
nand U1208 (N_1208,In_742,In_2212);
nor U1209 (N_1209,In_1594,In_303);
or U1210 (N_1210,In_1712,In_1240);
xnor U1211 (N_1211,In_2123,In_347);
and U1212 (N_1212,In_1430,In_553);
and U1213 (N_1213,In_1070,In_2418);
nor U1214 (N_1214,In_2351,In_531);
and U1215 (N_1215,In_366,In_1182);
nor U1216 (N_1216,In_1119,In_2280);
nor U1217 (N_1217,In_1492,In_992);
or U1218 (N_1218,In_1951,In_822);
nand U1219 (N_1219,In_723,In_2318);
nand U1220 (N_1220,In_2003,In_244);
or U1221 (N_1221,In_1664,In_709);
or U1222 (N_1222,In_1078,In_924);
or U1223 (N_1223,In_586,In_908);
or U1224 (N_1224,In_811,In_1798);
and U1225 (N_1225,In_1593,In_2451);
nand U1226 (N_1226,In_713,In_2176);
and U1227 (N_1227,In_1011,In_1448);
and U1228 (N_1228,In_372,In_640);
xnor U1229 (N_1229,In_1792,In_443);
nand U1230 (N_1230,In_149,In_606);
or U1231 (N_1231,In_221,In_1683);
xnor U1232 (N_1232,In_260,In_98);
or U1233 (N_1233,In_1003,In_418);
and U1234 (N_1234,In_2483,In_2078);
xor U1235 (N_1235,In_2319,In_1303);
nand U1236 (N_1236,In_585,In_2446);
or U1237 (N_1237,In_932,In_279);
xnor U1238 (N_1238,In_2268,In_1644);
and U1239 (N_1239,In_1629,In_1194);
nand U1240 (N_1240,In_1474,In_1626);
and U1241 (N_1241,In_1135,In_521);
or U1242 (N_1242,In_1363,In_572);
or U1243 (N_1243,In_2383,In_896);
or U1244 (N_1244,In_1652,In_1339);
nor U1245 (N_1245,In_1572,In_1337);
nand U1246 (N_1246,In_2242,In_1260);
xnor U1247 (N_1247,In_1377,In_1030);
nand U1248 (N_1248,In_1514,In_263);
and U1249 (N_1249,In_708,In_726);
nor U1250 (N_1250,In_1158,In_939);
nand U1251 (N_1251,In_1542,In_567);
nor U1252 (N_1252,In_1306,In_1171);
and U1253 (N_1253,In_1397,In_730);
nor U1254 (N_1254,In_1723,In_2003);
nand U1255 (N_1255,In_446,In_121);
xor U1256 (N_1256,In_1334,In_472);
nand U1257 (N_1257,In_1766,In_403);
or U1258 (N_1258,In_1233,In_37);
or U1259 (N_1259,In_1174,In_1957);
or U1260 (N_1260,In_777,In_1575);
nor U1261 (N_1261,In_1105,In_635);
and U1262 (N_1262,In_1791,In_1170);
nand U1263 (N_1263,In_1405,In_1554);
xor U1264 (N_1264,In_209,In_623);
nor U1265 (N_1265,In_355,In_1127);
and U1266 (N_1266,In_454,In_2331);
xnor U1267 (N_1267,In_2264,In_1984);
nand U1268 (N_1268,In_612,In_298);
nor U1269 (N_1269,In_398,In_215);
nand U1270 (N_1270,In_262,In_2079);
nor U1271 (N_1271,In_344,In_1881);
nand U1272 (N_1272,In_315,In_614);
and U1273 (N_1273,In_972,In_2454);
or U1274 (N_1274,In_2361,In_1829);
nor U1275 (N_1275,In_129,In_1937);
nor U1276 (N_1276,In_349,In_6);
nand U1277 (N_1277,In_1051,In_2167);
xnor U1278 (N_1278,In_1088,In_232);
nor U1279 (N_1279,In_1287,In_913);
and U1280 (N_1280,In_1095,In_1239);
or U1281 (N_1281,In_936,In_2387);
xor U1282 (N_1282,In_501,In_1273);
and U1283 (N_1283,In_230,In_794);
xor U1284 (N_1284,In_1331,In_743);
nor U1285 (N_1285,In_680,In_2316);
xnor U1286 (N_1286,In_1397,In_799);
xor U1287 (N_1287,In_222,In_1391);
nand U1288 (N_1288,In_1611,In_1826);
nor U1289 (N_1289,In_1570,In_1727);
or U1290 (N_1290,In_1017,In_113);
nand U1291 (N_1291,In_1237,In_947);
nor U1292 (N_1292,In_597,In_2167);
and U1293 (N_1293,In_901,In_1685);
xor U1294 (N_1294,In_340,In_2495);
or U1295 (N_1295,In_1452,In_1985);
or U1296 (N_1296,In_1926,In_1133);
xnor U1297 (N_1297,In_1681,In_1774);
and U1298 (N_1298,In_1045,In_50);
and U1299 (N_1299,In_530,In_757);
or U1300 (N_1300,In_1492,In_374);
nand U1301 (N_1301,In_1493,In_1248);
nand U1302 (N_1302,In_5,In_1624);
xor U1303 (N_1303,In_1340,In_1051);
nor U1304 (N_1304,In_2068,In_1104);
nor U1305 (N_1305,In_70,In_1545);
xor U1306 (N_1306,In_2081,In_1618);
or U1307 (N_1307,In_1794,In_1942);
or U1308 (N_1308,In_996,In_473);
nor U1309 (N_1309,In_740,In_2165);
nand U1310 (N_1310,In_1090,In_509);
nor U1311 (N_1311,In_1009,In_144);
nor U1312 (N_1312,In_118,In_2085);
nand U1313 (N_1313,In_2033,In_246);
nor U1314 (N_1314,In_2241,In_1748);
nor U1315 (N_1315,In_2124,In_852);
nor U1316 (N_1316,In_1455,In_1858);
nor U1317 (N_1317,In_177,In_1743);
xnor U1318 (N_1318,In_2335,In_1358);
and U1319 (N_1319,In_126,In_2202);
or U1320 (N_1320,In_1513,In_651);
nor U1321 (N_1321,In_1802,In_1979);
xnor U1322 (N_1322,In_2373,In_2291);
and U1323 (N_1323,In_1332,In_105);
and U1324 (N_1324,In_2049,In_2444);
nand U1325 (N_1325,In_2157,In_2255);
nor U1326 (N_1326,In_836,In_2103);
and U1327 (N_1327,In_1449,In_509);
xor U1328 (N_1328,In_1041,In_834);
nand U1329 (N_1329,In_834,In_1694);
and U1330 (N_1330,In_2164,In_1860);
xnor U1331 (N_1331,In_1618,In_1210);
xor U1332 (N_1332,In_2489,In_1082);
xnor U1333 (N_1333,In_669,In_1162);
xor U1334 (N_1334,In_2460,In_1066);
nand U1335 (N_1335,In_1400,In_2162);
nor U1336 (N_1336,In_1000,In_2021);
or U1337 (N_1337,In_592,In_546);
nor U1338 (N_1338,In_560,In_1315);
or U1339 (N_1339,In_373,In_1730);
nor U1340 (N_1340,In_1860,In_2429);
and U1341 (N_1341,In_375,In_1473);
xor U1342 (N_1342,In_1200,In_2001);
xnor U1343 (N_1343,In_228,In_125);
nand U1344 (N_1344,In_124,In_1923);
or U1345 (N_1345,In_1792,In_2242);
xor U1346 (N_1346,In_674,In_1862);
nor U1347 (N_1347,In_977,In_1961);
and U1348 (N_1348,In_747,In_2184);
nand U1349 (N_1349,In_1618,In_265);
nand U1350 (N_1350,In_1440,In_298);
xor U1351 (N_1351,In_818,In_1578);
nor U1352 (N_1352,In_1739,In_2482);
xnor U1353 (N_1353,In_1354,In_350);
nor U1354 (N_1354,In_2273,In_1585);
and U1355 (N_1355,In_1995,In_1318);
and U1356 (N_1356,In_2397,In_869);
xnor U1357 (N_1357,In_1914,In_1207);
xor U1358 (N_1358,In_372,In_2186);
nand U1359 (N_1359,In_2179,In_1285);
nand U1360 (N_1360,In_1399,In_1732);
and U1361 (N_1361,In_2061,In_1784);
and U1362 (N_1362,In_2084,In_1631);
nand U1363 (N_1363,In_2406,In_1993);
nor U1364 (N_1364,In_1007,In_2290);
and U1365 (N_1365,In_2447,In_1634);
xnor U1366 (N_1366,In_1360,In_747);
and U1367 (N_1367,In_143,In_2370);
nor U1368 (N_1368,In_1267,In_111);
xnor U1369 (N_1369,In_1626,In_747);
or U1370 (N_1370,In_765,In_762);
nor U1371 (N_1371,In_145,In_2026);
xor U1372 (N_1372,In_1913,In_394);
nand U1373 (N_1373,In_112,In_124);
nor U1374 (N_1374,In_2258,In_304);
or U1375 (N_1375,In_1965,In_960);
nand U1376 (N_1376,In_1892,In_1647);
nor U1377 (N_1377,In_685,In_268);
xnor U1378 (N_1378,In_93,In_719);
nand U1379 (N_1379,In_1659,In_654);
nor U1380 (N_1380,In_1075,In_2451);
nor U1381 (N_1381,In_1139,In_833);
nand U1382 (N_1382,In_842,In_1493);
and U1383 (N_1383,In_1939,In_582);
nor U1384 (N_1384,In_2341,In_2462);
xor U1385 (N_1385,In_661,In_100);
or U1386 (N_1386,In_2009,In_235);
or U1387 (N_1387,In_1189,In_1676);
nand U1388 (N_1388,In_754,In_1389);
or U1389 (N_1389,In_757,In_1268);
and U1390 (N_1390,In_1304,In_1575);
and U1391 (N_1391,In_2049,In_1917);
xnor U1392 (N_1392,In_715,In_2012);
or U1393 (N_1393,In_1121,In_1423);
or U1394 (N_1394,In_2054,In_1945);
nand U1395 (N_1395,In_935,In_763);
xor U1396 (N_1396,In_805,In_257);
nand U1397 (N_1397,In_1308,In_45);
xor U1398 (N_1398,In_1927,In_1539);
or U1399 (N_1399,In_2463,In_912);
nand U1400 (N_1400,In_841,In_676);
and U1401 (N_1401,In_146,In_1484);
nand U1402 (N_1402,In_1253,In_618);
nand U1403 (N_1403,In_1212,In_886);
and U1404 (N_1404,In_1429,In_717);
or U1405 (N_1405,In_682,In_698);
xor U1406 (N_1406,In_2083,In_253);
or U1407 (N_1407,In_1359,In_2025);
nand U1408 (N_1408,In_763,In_1835);
nand U1409 (N_1409,In_2170,In_97);
xnor U1410 (N_1410,In_1851,In_179);
or U1411 (N_1411,In_2450,In_2056);
nand U1412 (N_1412,In_121,In_1697);
nand U1413 (N_1413,In_286,In_1373);
xnor U1414 (N_1414,In_1300,In_1923);
nor U1415 (N_1415,In_1864,In_1865);
or U1416 (N_1416,In_1299,In_1472);
and U1417 (N_1417,In_2383,In_2181);
nand U1418 (N_1418,In_26,In_2290);
and U1419 (N_1419,In_460,In_992);
nand U1420 (N_1420,In_1321,In_1769);
xor U1421 (N_1421,In_132,In_187);
xnor U1422 (N_1422,In_730,In_856);
nor U1423 (N_1423,In_411,In_816);
or U1424 (N_1424,In_1349,In_25);
nor U1425 (N_1425,In_684,In_286);
xor U1426 (N_1426,In_2310,In_1305);
and U1427 (N_1427,In_399,In_916);
nand U1428 (N_1428,In_2020,In_442);
xnor U1429 (N_1429,In_354,In_2212);
and U1430 (N_1430,In_1627,In_658);
xnor U1431 (N_1431,In_722,In_1840);
nor U1432 (N_1432,In_361,In_2250);
and U1433 (N_1433,In_1586,In_1680);
nor U1434 (N_1434,In_88,In_2154);
xnor U1435 (N_1435,In_76,In_2149);
and U1436 (N_1436,In_1291,In_2015);
or U1437 (N_1437,In_2092,In_214);
nor U1438 (N_1438,In_597,In_1473);
nor U1439 (N_1439,In_2496,In_1757);
nor U1440 (N_1440,In_143,In_506);
xor U1441 (N_1441,In_1283,In_1841);
xor U1442 (N_1442,In_1994,In_1250);
xnor U1443 (N_1443,In_1429,In_2473);
and U1444 (N_1444,In_958,In_77);
nor U1445 (N_1445,In_217,In_1838);
or U1446 (N_1446,In_1169,In_1633);
and U1447 (N_1447,In_338,In_147);
or U1448 (N_1448,In_312,In_1029);
or U1449 (N_1449,In_128,In_1141);
nor U1450 (N_1450,In_771,In_152);
or U1451 (N_1451,In_2345,In_1686);
or U1452 (N_1452,In_755,In_739);
nand U1453 (N_1453,In_1091,In_2259);
and U1454 (N_1454,In_396,In_2404);
xor U1455 (N_1455,In_2485,In_1615);
or U1456 (N_1456,In_630,In_1082);
and U1457 (N_1457,In_175,In_891);
or U1458 (N_1458,In_1895,In_800);
nor U1459 (N_1459,In_2462,In_2298);
and U1460 (N_1460,In_1342,In_570);
xor U1461 (N_1461,In_2187,In_1467);
or U1462 (N_1462,In_1834,In_2173);
nand U1463 (N_1463,In_83,In_2081);
or U1464 (N_1464,In_2353,In_189);
nor U1465 (N_1465,In_721,In_768);
xnor U1466 (N_1466,In_2009,In_1741);
and U1467 (N_1467,In_2218,In_1073);
nor U1468 (N_1468,In_1873,In_158);
or U1469 (N_1469,In_20,In_2091);
nor U1470 (N_1470,In_446,In_1043);
or U1471 (N_1471,In_2075,In_2164);
nand U1472 (N_1472,In_2296,In_792);
xor U1473 (N_1473,In_418,In_48);
nand U1474 (N_1474,In_553,In_309);
xor U1475 (N_1475,In_2360,In_0);
or U1476 (N_1476,In_2493,In_1641);
nor U1477 (N_1477,In_1664,In_1189);
xnor U1478 (N_1478,In_1309,In_418);
xnor U1479 (N_1479,In_2137,In_2450);
nor U1480 (N_1480,In_1376,In_306);
xnor U1481 (N_1481,In_1588,In_61);
nand U1482 (N_1482,In_1576,In_2418);
xor U1483 (N_1483,In_516,In_701);
or U1484 (N_1484,In_2050,In_914);
nor U1485 (N_1485,In_826,In_767);
and U1486 (N_1486,In_666,In_1655);
xor U1487 (N_1487,In_469,In_537);
and U1488 (N_1488,In_608,In_912);
nand U1489 (N_1489,In_115,In_1090);
nand U1490 (N_1490,In_886,In_2441);
or U1491 (N_1491,In_433,In_1131);
nor U1492 (N_1492,In_947,In_0);
nor U1493 (N_1493,In_1291,In_2312);
and U1494 (N_1494,In_111,In_85);
xor U1495 (N_1495,In_2315,In_2258);
nand U1496 (N_1496,In_1769,In_1529);
xor U1497 (N_1497,In_965,In_554);
nand U1498 (N_1498,In_272,In_2186);
xor U1499 (N_1499,In_756,In_613);
nor U1500 (N_1500,In_359,In_846);
xnor U1501 (N_1501,In_189,In_282);
xnor U1502 (N_1502,In_2319,In_73);
or U1503 (N_1503,In_1798,In_1533);
nor U1504 (N_1504,In_1406,In_2495);
or U1505 (N_1505,In_214,In_1772);
and U1506 (N_1506,In_1002,In_293);
and U1507 (N_1507,In_228,In_2239);
nand U1508 (N_1508,In_2372,In_2296);
nor U1509 (N_1509,In_513,In_1311);
or U1510 (N_1510,In_218,In_1137);
and U1511 (N_1511,In_1336,In_1297);
xnor U1512 (N_1512,In_2053,In_2329);
nor U1513 (N_1513,In_1491,In_2321);
and U1514 (N_1514,In_182,In_29);
xor U1515 (N_1515,In_1695,In_2047);
nor U1516 (N_1516,In_1167,In_2055);
and U1517 (N_1517,In_2456,In_1486);
nor U1518 (N_1518,In_466,In_2468);
nor U1519 (N_1519,In_1626,In_1605);
or U1520 (N_1520,In_1198,In_1381);
nand U1521 (N_1521,In_2161,In_39);
nand U1522 (N_1522,In_860,In_501);
xnor U1523 (N_1523,In_2132,In_2331);
nand U1524 (N_1524,In_2404,In_2376);
nand U1525 (N_1525,In_320,In_2473);
and U1526 (N_1526,In_1155,In_1999);
nand U1527 (N_1527,In_438,In_2484);
and U1528 (N_1528,In_2042,In_19);
nand U1529 (N_1529,In_671,In_2336);
nor U1530 (N_1530,In_2051,In_1463);
xnor U1531 (N_1531,In_452,In_2099);
nor U1532 (N_1532,In_815,In_1897);
nor U1533 (N_1533,In_483,In_480);
xor U1534 (N_1534,In_1023,In_115);
and U1535 (N_1535,In_152,In_1726);
nand U1536 (N_1536,In_257,In_44);
or U1537 (N_1537,In_1386,In_760);
nand U1538 (N_1538,In_1499,In_2369);
nand U1539 (N_1539,In_1269,In_831);
or U1540 (N_1540,In_1714,In_1615);
nand U1541 (N_1541,In_774,In_1884);
xnor U1542 (N_1542,In_1833,In_817);
nor U1543 (N_1543,In_354,In_1861);
nand U1544 (N_1544,In_2199,In_136);
nand U1545 (N_1545,In_798,In_2340);
xnor U1546 (N_1546,In_372,In_276);
xor U1547 (N_1547,In_141,In_1427);
or U1548 (N_1548,In_457,In_679);
or U1549 (N_1549,In_1933,In_50);
and U1550 (N_1550,In_1066,In_237);
nor U1551 (N_1551,In_769,In_1670);
xnor U1552 (N_1552,In_2164,In_1923);
nor U1553 (N_1553,In_207,In_2407);
or U1554 (N_1554,In_50,In_1397);
xor U1555 (N_1555,In_936,In_12);
nand U1556 (N_1556,In_1103,In_2240);
xnor U1557 (N_1557,In_1042,In_684);
and U1558 (N_1558,In_2182,In_1395);
or U1559 (N_1559,In_1993,In_2487);
nor U1560 (N_1560,In_1295,In_1345);
or U1561 (N_1561,In_2103,In_1002);
nand U1562 (N_1562,In_2204,In_1866);
and U1563 (N_1563,In_1914,In_127);
nand U1564 (N_1564,In_1825,In_1092);
nand U1565 (N_1565,In_2101,In_592);
nand U1566 (N_1566,In_2164,In_1555);
xor U1567 (N_1567,In_661,In_1524);
xnor U1568 (N_1568,In_866,In_1637);
or U1569 (N_1569,In_528,In_748);
and U1570 (N_1570,In_221,In_2256);
nor U1571 (N_1571,In_517,In_268);
and U1572 (N_1572,In_765,In_2368);
nor U1573 (N_1573,In_819,In_144);
xor U1574 (N_1574,In_93,In_2239);
nor U1575 (N_1575,In_1897,In_248);
and U1576 (N_1576,In_793,In_1831);
nand U1577 (N_1577,In_1621,In_2056);
and U1578 (N_1578,In_1000,In_945);
xnor U1579 (N_1579,In_61,In_1058);
and U1580 (N_1580,In_850,In_284);
nor U1581 (N_1581,In_2216,In_558);
xnor U1582 (N_1582,In_1687,In_538);
or U1583 (N_1583,In_1038,In_1439);
xnor U1584 (N_1584,In_872,In_2052);
nor U1585 (N_1585,In_1122,In_2439);
and U1586 (N_1586,In_66,In_1405);
nor U1587 (N_1587,In_655,In_1126);
nand U1588 (N_1588,In_681,In_1256);
or U1589 (N_1589,In_1440,In_1050);
nor U1590 (N_1590,In_1708,In_498);
nor U1591 (N_1591,In_2117,In_544);
nand U1592 (N_1592,In_64,In_325);
or U1593 (N_1593,In_682,In_212);
and U1594 (N_1594,In_1996,In_674);
xnor U1595 (N_1595,In_2447,In_2427);
nor U1596 (N_1596,In_1338,In_419);
and U1597 (N_1597,In_1818,In_636);
and U1598 (N_1598,In_978,In_2027);
or U1599 (N_1599,In_2279,In_1256);
or U1600 (N_1600,In_813,In_803);
and U1601 (N_1601,In_2244,In_1106);
nand U1602 (N_1602,In_2159,In_1965);
nand U1603 (N_1603,In_1294,In_1103);
xor U1604 (N_1604,In_1532,In_2442);
nor U1605 (N_1605,In_2171,In_1561);
or U1606 (N_1606,In_1919,In_1041);
nor U1607 (N_1607,In_486,In_1343);
and U1608 (N_1608,In_1310,In_293);
nor U1609 (N_1609,In_1823,In_915);
xor U1610 (N_1610,In_1618,In_1527);
nor U1611 (N_1611,In_472,In_1653);
nor U1612 (N_1612,In_1828,In_199);
nor U1613 (N_1613,In_1600,In_229);
nand U1614 (N_1614,In_200,In_2221);
and U1615 (N_1615,In_1172,In_2218);
nor U1616 (N_1616,In_2454,In_355);
or U1617 (N_1617,In_285,In_2407);
or U1618 (N_1618,In_464,In_1579);
nor U1619 (N_1619,In_1098,In_1310);
or U1620 (N_1620,In_1092,In_360);
xor U1621 (N_1621,In_173,In_56);
xnor U1622 (N_1622,In_257,In_845);
nor U1623 (N_1623,In_545,In_1435);
nand U1624 (N_1624,In_107,In_300);
or U1625 (N_1625,In_72,In_2419);
nor U1626 (N_1626,In_84,In_773);
or U1627 (N_1627,In_516,In_1303);
nor U1628 (N_1628,In_199,In_363);
and U1629 (N_1629,In_251,In_2351);
nand U1630 (N_1630,In_1733,In_1618);
xor U1631 (N_1631,In_424,In_663);
nand U1632 (N_1632,In_772,In_379);
and U1633 (N_1633,In_1790,In_1996);
nand U1634 (N_1634,In_245,In_1087);
or U1635 (N_1635,In_2326,In_1161);
nand U1636 (N_1636,In_871,In_1808);
nand U1637 (N_1637,In_1572,In_907);
xnor U1638 (N_1638,In_729,In_320);
nand U1639 (N_1639,In_105,In_914);
nor U1640 (N_1640,In_44,In_50);
and U1641 (N_1641,In_2136,In_1808);
and U1642 (N_1642,In_2239,In_150);
xnor U1643 (N_1643,In_1795,In_2370);
or U1644 (N_1644,In_1635,In_205);
and U1645 (N_1645,In_1441,In_163);
nand U1646 (N_1646,In_1892,In_681);
or U1647 (N_1647,In_2368,In_1124);
and U1648 (N_1648,In_2162,In_686);
or U1649 (N_1649,In_2464,In_1466);
xnor U1650 (N_1650,In_194,In_2074);
nor U1651 (N_1651,In_1732,In_1617);
nand U1652 (N_1652,In_1414,In_456);
and U1653 (N_1653,In_1777,In_2173);
nand U1654 (N_1654,In_2433,In_1724);
xor U1655 (N_1655,In_1401,In_521);
xnor U1656 (N_1656,In_1096,In_873);
or U1657 (N_1657,In_1289,In_1886);
nor U1658 (N_1658,In_1003,In_1060);
nor U1659 (N_1659,In_522,In_925);
nand U1660 (N_1660,In_949,In_812);
nor U1661 (N_1661,In_1776,In_1055);
xnor U1662 (N_1662,In_87,In_2145);
nand U1663 (N_1663,In_1766,In_1482);
or U1664 (N_1664,In_1830,In_2078);
and U1665 (N_1665,In_1088,In_565);
or U1666 (N_1666,In_160,In_1557);
nand U1667 (N_1667,In_1614,In_2048);
or U1668 (N_1668,In_2269,In_2350);
nor U1669 (N_1669,In_1388,In_1892);
nor U1670 (N_1670,In_627,In_548);
nor U1671 (N_1671,In_1262,In_357);
nand U1672 (N_1672,In_1710,In_492);
nand U1673 (N_1673,In_824,In_2128);
nor U1674 (N_1674,In_1429,In_366);
nand U1675 (N_1675,In_1178,In_1276);
nor U1676 (N_1676,In_1903,In_1540);
nor U1677 (N_1677,In_582,In_378);
xnor U1678 (N_1678,In_829,In_391);
or U1679 (N_1679,In_1516,In_1319);
or U1680 (N_1680,In_333,In_1065);
and U1681 (N_1681,In_316,In_1545);
xnor U1682 (N_1682,In_1247,In_1053);
nand U1683 (N_1683,In_1612,In_1661);
nor U1684 (N_1684,In_1490,In_1899);
nand U1685 (N_1685,In_435,In_903);
or U1686 (N_1686,In_392,In_836);
xnor U1687 (N_1687,In_1305,In_813);
xnor U1688 (N_1688,In_684,In_2225);
and U1689 (N_1689,In_1900,In_2297);
nand U1690 (N_1690,In_1197,In_2303);
nor U1691 (N_1691,In_2116,In_1537);
or U1692 (N_1692,In_1006,In_2496);
or U1693 (N_1693,In_432,In_758);
nor U1694 (N_1694,In_987,In_2220);
or U1695 (N_1695,In_785,In_1916);
xor U1696 (N_1696,In_2234,In_686);
xor U1697 (N_1697,In_137,In_941);
or U1698 (N_1698,In_2211,In_411);
or U1699 (N_1699,In_346,In_1251);
or U1700 (N_1700,In_1397,In_805);
or U1701 (N_1701,In_61,In_1854);
nor U1702 (N_1702,In_1045,In_2313);
nor U1703 (N_1703,In_2412,In_662);
nor U1704 (N_1704,In_2102,In_831);
nor U1705 (N_1705,In_87,In_2223);
or U1706 (N_1706,In_2205,In_746);
xnor U1707 (N_1707,In_2174,In_1264);
and U1708 (N_1708,In_1942,In_488);
xor U1709 (N_1709,In_840,In_2202);
nand U1710 (N_1710,In_263,In_2106);
and U1711 (N_1711,In_2396,In_2052);
nand U1712 (N_1712,In_93,In_226);
and U1713 (N_1713,In_290,In_2434);
and U1714 (N_1714,In_1189,In_1148);
and U1715 (N_1715,In_1865,In_839);
nor U1716 (N_1716,In_2157,In_1962);
xnor U1717 (N_1717,In_310,In_257);
nor U1718 (N_1718,In_1310,In_1190);
or U1719 (N_1719,In_982,In_181);
or U1720 (N_1720,In_659,In_1574);
xor U1721 (N_1721,In_1462,In_1180);
and U1722 (N_1722,In_1159,In_779);
or U1723 (N_1723,In_981,In_1114);
nor U1724 (N_1724,In_1534,In_1704);
xnor U1725 (N_1725,In_1685,In_1549);
and U1726 (N_1726,In_2084,In_1375);
nand U1727 (N_1727,In_858,In_1093);
and U1728 (N_1728,In_2323,In_2403);
or U1729 (N_1729,In_585,In_1906);
nor U1730 (N_1730,In_1042,In_2341);
nand U1731 (N_1731,In_1438,In_813);
or U1732 (N_1732,In_1526,In_2110);
or U1733 (N_1733,In_1958,In_471);
nand U1734 (N_1734,In_2403,In_2476);
and U1735 (N_1735,In_1332,In_1948);
or U1736 (N_1736,In_1120,In_1386);
and U1737 (N_1737,In_252,In_521);
xnor U1738 (N_1738,In_481,In_1881);
xnor U1739 (N_1739,In_1973,In_2171);
xor U1740 (N_1740,In_1041,In_2388);
nor U1741 (N_1741,In_825,In_1547);
or U1742 (N_1742,In_294,In_2195);
and U1743 (N_1743,In_64,In_1460);
or U1744 (N_1744,In_1540,In_1121);
nor U1745 (N_1745,In_485,In_768);
nand U1746 (N_1746,In_1308,In_295);
nand U1747 (N_1747,In_223,In_2201);
nand U1748 (N_1748,In_2052,In_2372);
nor U1749 (N_1749,In_8,In_1129);
and U1750 (N_1750,In_806,In_1073);
xor U1751 (N_1751,In_896,In_13);
nand U1752 (N_1752,In_659,In_2161);
or U1753 (N_1753,In_1018,In_2118);
xnor U1754 (N_1754,In_964,In_2358);
nand U1755 (N_1755,In_1474,In_1613);
and U1756 (N_1756,In_565,In_560);
nand U1757 (N_1757,In_648,In_2073);
xor U1758 (N_1758,In_1239,In_554);
nor U1759 (N_1759,In_2218,In_2182);
nor U1760 (N_1760,In_34,In_277);
xnor U1761 (N_1761,In_2353,In_2306);
nand U1762 (N_1762,In_1460,In_628);
nor U1763 (N_1763,In_1625,In_39);
xnor U1764 (N_1764,In_1130,In_780);
or U1765 (N_1765,In_1717,In_333);
xnor U1766 (N_1766,In_191,In_251);
nor U1767 (N_1767,In_2228,In_1053);
nor U1768 (N_1768,In_2293,In_666);
xnor U1769 (N_1769,In_2113,In_1297);
nor U1770 (N_1770,In_2481,In_1284);
xnor U1771 (N_1771,In_2140,In_620);
or U1772 (N_1772,In_1220,In_1285);
nor U1773 (N_1773,In_963,In_1860);
nand U1774 (N_1774,In_917,In_1143);
or U1775 (N_1775,In_1859,In_1742);
nand U1776 (N_1776,In_729,In_1561);
nand U1777 (N_1777,In_1280,In_1330);
or U1778 (N_1778,In_1459,In_1094);
nand U1779 (N_1779,In_1611,In_30);
or U1780 (N_1780,In_1481,In_1026);
xnor U1781 (N_1781,In_1887,In_1030);
and U1782 (N_1782,In_222,In_2141);
or U1783 (N_1783,In_1665,In_1794);
xnor U1784 (N_1784,In_2159,In_1325);
xor U1785 (N_1785,In_1828,In_1891);
xor U1786 (N_1786,In_542,In_703);
or U1787 (N_1787,In_1246,In_1524);
and U1788 (N_1788,In_33,In_1678);
nor U1789 (N_1789,In_915,In_1802);
and U1790 (N_1790,In_2147,In_192);
xor U1791 (N_1791,In_746,In_1452);
or U1792 (N_1792,In_1,In_426);
and U1793 (N_1793,In_1335,In_1640);
nand U1794 (N_1794,In_813,In_1649);
and U1795 (N_1795,In_1403,In_1216);
xor U1796 (N_1796,In_1113,In_1715);
or U1797 (N_1797,In_1246,In_2244);
nand U1798 (N_1798,In_1136,In_2108);
nor U1799 (N_1799,In_263,In_877);
or U1800 (N_1800,In_560,In_2400);
nor U1801 (N_1801,In_1593,In_166);
xnor U1802 (N_1802,In_1325,In_1416);
nor U1803 (N_1803,In_610,In_132);
nor U1804 (N_1804,In_2251,In_1321);
and U1805 (N_1805,In_1729,In_1757);
xor U1806 (N_1806,In_1863,In_2188);
nor U1807 (N_1807,In_2074,In_2375);
or U1808 (N_1808,In_2261,In_1636);
nand U1809 (N_1809,In_2441,In_493);
xor U1810 (N_1810,In_1237,In_2291);
xor U1811 (N_1811,In_615,In_1442);
nand U1812 (N_1812,In_1324,In_1561);
nand U1813 (N_1813,In_562,In_469);
xnor U1814 (N_1814,In_2114,In_1099);
nand U1815 (N_1815,In_2412,In_1890);
and U1816 (N_1816,In_2437,In_2234);
xor U1817 (N_1817,In_1881,In_2135);
or U1818 (N_1818,In_425,In_1192);
nor U1819 (N_1819,In_602,In_550);
or U1820 (N_1820,In_1427,In_2011);
nor U1821 (N_1821,In_956,In_515);
or U1822 (N_1822,In_2297,In_1456);
or U1823 (N_1823,In_1994,In_1049);
or U1824 (N_1824,In_1694,In_1600);
or U1825 (N_1825,In_2027,In_1324);
nand U1826 (N_1826,In_1336,In_1996);
nor U1827 (N_1827,In_1614,In_1215);
nor U1828 (N_1828,In_1416,In_188);
xor U1829 (N_1829,In_1077,In_2485);
xnor U1830 (N_1830,In_238,In_210);
or U1831 (N_1831,In_1463,In_1702);
or U1832 (N_1832,In_1380,In_2234);
and U1833 (N_1833,In_1000,In_2133);
and U1834 (N_1834,In_1017,In_643);
or U1835 (N_1835,In_2327,In_160);
or U1836 (N_1836,In_1768,In_619);
and U1837 (N_1837,In_1427,In_1119);
and U1838 (N_1838,In_392,In_1410);
nand U1839 (N_1839,In_2303,In_1875);
nor U1840 (N_1840,In_35,In_728);
nor U1841 (N_1841,In_1242,In_64);
and U1842 (N_1842,In_550,In_705);
xnor U1843 (N_1843,In_1257,In_623);
nand U1844 (N_1844,In_2408,In_1232);
and U1845 (N_1845,In_1801,In_448);
xor U1846 (N_1846,In_844,In_2154);
xnor U1847 (N_1847,In_1575,In_632);
or U1848 (N_1848,In_144,In_1356);
xnor U1849 (N_1849,In_1584,In_743);
nor U1850 (N_1850,In_829,In_130);
nand U1851 (N_1851,In_2051,In_197);
and U1852 (N_1852,In_1397,In_1024);
and U1853 (N_1853,In_1443,In_80);
xnor U1854 (N_1854,In_1967,In_489);
xnor U1855 (N_1855,In_2144,In_1961);
xor U1856 (N_1856,In_1429,In_1843);
and U1857 (N_1857,In_1892,In_1146);
and U1858 (N_1858,In_1241,In_288);
or U1859 (N_1859,In_335,In_1002);
xor U1860 (N_1860,In_1504,In_2353);
or U1861 (N_1861,In_47,In_1921);
and U1862 (N_1862,In_1787,In_1190);
xor U1863 (N_1863,In_1490,In_2085);
xnor U1864 (N_1864,In_564,In_449);
nor U1865 (N_1865,In_1744,In_221);
xor U1866 (N_1866,In_1413,In_465);
nand U1867 (N_1867,In_1281,In_364);
xnor U1868 (N_1868,In_1621,In_378);
and U1869 (N_1869,In_2159,In_277);
xor U1870 (N_1870,In_2063,In_570);
or U1871 (N_1871,In_963,In_1677);
nor U1872 (N_1872,In_212,In_744);
nor U1873 (N_1873,In_1328,In_1524);
or U1874 (N_1874,In_111,In_288);
and U1875 (N_1875,In_2095,In_1438);
xnor U1876 (N_1876,In_446,In_157);
xor U1877 (N_1877,In_1804,In_278);
and U1878 (N_1878,In_899,In_1582);
and U1879 (N_1879,In_880,In_1860);
or U1880 (N_1880,In_1365,In_1507);
nor U1881 (N_1881,In_1757,In_2188);
and U1882 (N_1882,In_1323,In_1022);
xnor U1883 (N_1883,In_576,In_1923);
nor U1884 (N_1884,In_467,In_1754);
and U1885 (N_1885,In_1469,In_2430);
and U1886 (N_1886,In_691,In_716);
nand U1887 (N_1887,In_2284,In_1146);
and U1888 (N_1888,In_970,In_1343);
or U1889 (N_1889,In_2354,In_2179);
nand U1890 (N_1890,In_17,In_2486);
nand U1891 (N_1891,In_1354,In_484);
or U1892 (N_1892,In_335,In_1483);
and U1893 (N_1893,In_1738,In_2291);
nor U1894 (N_1894,In_1507,In_1721);
or U1895 (N_1895,In_1230,In_1710);
or U1896 (N_1896,In_2150,In_164);
xnor U1897 (N_1897,In_2476,In_101);
or U1898 (N_1898,In_1826,In_1339);
and U1899 (N_1899,In_1878,In_2);
or U1900 (N_1900,In_625,In_1693);
and U1901 (N_1901,In_593,In_384);
xnor U1902 (N_1902,In_1628,In_786);
xor U1903 (N_1903,In_2364,In_1626);
nor U1904 (N_1904,In_1410,In_1767);
nor U1905 (N_1905,In_123,In_924);
and U1906 (N_1906,In_2139,In_1279);
and U1907 (N_1907,In_1821,In_198);
nor U1908 (N_1908,In_1684,In_2030);
and U1909 (N_1909,In_643,In_716);
nand U1910 (N_1910,In_603,In_1034);
nor U1911 (N_1911,In_1462,In_1970);
and U1912 (N_1912,In_1151,In_1688);
nor U1913 (N_1913,In_2448,In_332);
and U1914 (N_1914,In_713,In_518);
and U1915 (N_1915,In_1394,In_1136);
or U1916 (N_1916,In_47,In_392);
and U1917 (N_1917,In_1667,In_846);
and U1918 (N_1918,In_2289,In_998);
nor U1919 (N_1919,In_2268,In_1721);
or U1920 (N_1920,In_2255,In_257);
nand U1921 (N_1921,In_1892,In_710);
nand U1922 (N_1922,In_1436,In_228);
and U1923 (N_1923,In_509,In_305);
xor U1924 (N_1924,In_937,In_1867);
xnor U1925 (N_1925,In_956,In_1802);
nor U1926 (N_1926,In_1752,In_1037);
or U1927 (N_1927,In_1289,In_522);
or U1928 (N_1928,In_2160,In_525);
or U1929 (N_1929,In_1966,In_2178);
or U1930 (N_1930,In_401,In_873);
and U1931 (N_1931,In_1462,In_1066);
and U1932 (N_1932,In_1505,In_810);
or U1933 (N_1933,In_120,In_1378);
and U1934 (N_1934,In_998,In_489);
or U1935 (N_1935,In_781,In_1914);
xor U1936 (N_1936,In_2361,In_1932);
or U1937 (N_1937,In_2455,In_203);
xor U1938 (N_1938,In_167,In_97);
nor U1939 (N_1939,In_1162,In_1597);
nand U1940 (N_1940,In_968,In_1243);
or U1941 (N_1941,In_1801,In_1595);
nor U1942 (N_1942,In_1955,In_2152);
xor U1943 (N_1943,In_2207,In_303);
nor U1944 (N_1944,In_117,In_1558);
nand U1945 (N_1945,In_1322,In_2289);
nand U1946 (N_1946,In_1951,In_2351);
xnor U1947 (N_1947,In_42,In_1770);
or U1948 (N_1948,In_1034,In_401);
nand U1949 (N_1949,In_414,In_736);
xor U1950 (N_1950,In_807,In_279);
nand U1951 (N_1951,In_1421,In_523);
xnor U1952 (N_1952,In_2403,In_1980);
nor U1953 (N_1953,In_640,In_1058);
xnor U1954 (N_1954,In_191,In_1777);
nand U1955 (N_1955,In_226,In_2151);
and U1956 (N_1956,In_1552,In_1282);
nand U1957 (N_1957,In_225,In_710);
nor U1958 (N_1958,In_253,In_303);
xnor U1959 (N_1959,In_1452,In_1790);
or U1960 (N_1960,In_2181,In_2037);
or U1961 (N_1961,In_1861,In_175);
or U1962 (N_1962,In_729,In_993);
xor U1963 (N_1963,In_96,In_1454);
xnor U1964 (N_1964,In_1699,In_1266);
nor U1965 (N_1965,In_415,In_2278);
nor U1966 (N_1966,In_1111,In_2083);
or U1967 (N_1967,In_702,In_1292);
nand U1968 (N_1968,In_2458,In_534);
nand U1969 (N_1969,In_992,In_1460);
and U1970 (N_1970,In_676,In_2415);
nor U1971 (N_1971,In_201,In_547);
or U1972 (N_1972,In_489,In_785);
xnor U1973 (N_1973,In_1436,In_974);
xnor U1974 (N_1974,In_540,In_1460);
nand U1975 (N_1975,In_845,In_271);
and U1976 (N_1976,In_1923,In_2160);
xnor U1977 (N_1977,In_949,In_1157);
xnor U1978 (N_1978,In_2043,In_1672);
xnor U1979 (N_1979,In_1022,In_235);
nor U1980 (N_1980,In_652,In_971);
nand U1981 (N_1981,In_1126,In_1925);
and U1982 (N_1982,In_603,In_537);
xnor U1983 (N_1983,In_1661,In_1077);
or U1984 (N_1984,In_1526,In_384);
nand U1985 (N_1985,In_2456,In_243);
and U1986 (N_1986,In_1196,In_1605);
xor U1987 (N_1987,In_1483,In_821);
or U1988 (N_1988,In_1949,In_1533);
or U1989 (N_1989,In_1617,In_317);
and U1990 (N_1990,In_1895,In_2466);
or U1991 (N_1991,In_889,In_431);
and U1992 (N_1992,In_406,In_262);
nand U1993 (N_1993,In_1876,In_2443);
nand U1994 (N_1994,In_1665,In_1496);
xor U1995 (N_1995,In_223,In_232);
nand U1996 (N_1996,In_1632,In_940);
xor U1997 (N_1997,In_1182,In_2063);
and U1998 (N_1998,In_397,In_426);
or U1999 (N_1999,In_2118,In_1079);
nand U2000 (N_2000,In_1977,In_1204);
nor U2001 (N_2001,In_996,In_2224);
nand U2002 (N_2002,In_973,In_1061);
or U2003 (N_2003,In_319,In_2424);
and U2004 (N_2004,In_327,In_481);
xnor U2005 (N_2005,In_1042,In_1530);
nand U2006 (N_2006,In_890,In_63);
nand U2007 (N_2007,In_1615,In_811);
nand U2008 (N_2008,In_395,In_2351);
and U2009 (N_2009,In_1418,In_2411);
and U2010 (N_2010,In_2262,In_1651);
or U2011 (N_2011,In_1150,In_865);
and U2012 (N_2012,In_807,In_2184);
xor U2013 (N_2013,In_115,In_897);
or U2014 (N_2014,In_603,In_1639);
and U2015 (N_2015,In_1385,In_1983);
nand U2016 (N_2016,In_793,In_154);
and U2017 (N_2017,In_1348,In_1429);
nand U2018 (N_2018,In_1235,In_2293);
xnor U2019 (N_2019,In_280,In_1507);
or U2020 (N_2020,In_1159,In_1911);
or U2021 (N_2021,In_648,In_1790);
or U2022 (N_2022,In_1693,In_386);
or U2023 (N_2023,In_727,In_1865);
or U2024 (N_2024,In_1019,In_2326);
or U2025 (N_2025,In_231,In_2110);
or U2026 (N_2026,In_101,In_1725);
nor U2027 (N_2027,In_2102,In_2237);
xor U2028 (N_2028,In_1168,In_276);
xnor U2029 (N_2029,In_567,In_1175);
xnor U2030 (N_2030,In_1144,In_5);
xor U2031 (N_2031,In_811,In_246);
and U2032 (N_2032,In_2040,In_590);
nor U2033 (N_2033,In_495,In_516);
or U2034 (N_2034,In_1544,In_234);
or U2035 (N_2035,In_2080,In_1718);
nand U2036 (N_2036,In_534,In_1701);
nand U2037 (N_2037,In_1550,In_1321);
and U2038 (N_2038,In_2363,In_725);
and U2039 (N_2039,In_1960,In_297);
or U2040 (N_2040,In_1235,In_1208);
or U2041 (N_2041,In_2067,In_1149);
and U2042 (N_2042,In_1057,In_1419);
nor U2043 (N_2043,In_2135,In_163);
and U2044 (N_2044,In_1034,In_2110);
nor U2045 (N_2045,In_680,In_2343);
or U2046 (N_2046,In_2300,In_2073);
nor U2047 (N_2047,In_2085,In_2318);
or U2048 (N_2048,In_393,In_428);
and U2049 (N_2049,In_1455,In_2336);
nand U2050 (N_2050,In_1734,In_1656);
or U2051 (N_2051,In_90,In_414);
or U2052 (N_2052,In_1999,In_1492);
nand U2053 (N_2053,In_1609,In_2164);
nor U2054 (N_2054,In_21,In_280);
or U2055 (N_2055,In_767,In_638);
xnor U2056 (N_2056,In_1585,In_559);
nand U2057 (N_2057,In_2065,In_947);
nand U2058 (N_2058,In_30,In_2382);
and U2059 (N_2059,In_191,In_2026);
nand U2060 (N_2060,In_2289,In_2045);
nor U2061 (N_2061,In_2016,In_439);
or U2062 (N_2062,In_532,In_206);
and U2063 (N_2063,In_1007,In_1165);
xor U2064 (N_2064,In_2364,In_1313);
nand U2065 (N_2065,In_1180,In_1688);
xor U2066 (N_2066,In_1750,In_1200);
xnor U2067 (N_2067,In_1182,In_1481);
xor U2068 (N_2068,In_760,In_108);
nor U2069 (N_2069,In_1366,In_301);
nand U2070 (N_2070,In_575,In_2332);
xor U2071 (N_2071,In_2169,In_1971);
and U2072 (N_2072,In_797,In_1714);
nand U2073 (N_2073,In_2455,In_495);
xor U2074 (N_2074,In_610,In_1470);
and U2075 (N_2075,In_1225,In_219);
xnor U2076 (N_2076,In_1670,In_758);
and U2077 (N_2077,In_2027,In_1522);
and U2078 (N_2078,In_1837,In_2053);
nor U2079 (N_2079,In_1624,In_1373);
xor U2080 (N_2080,In_225,In_174);
or U2081 (N_2081,In_1428,In_24);
and U2082 (N_2082,In_1791,In_1322);
nor U2083 (N_2083,In_1153,In_1974);
and U2084 (N_2084,In_1769,In_1066);
and U2085 (N_2085,In_148,In_1523);
and U2086 (N_2086,In_1033,In_576);
and U2087 (N_2087,In_908,In_1511);
nor U2088 (N_2088,In_684,In_344);
nor U2089 (N_2089,In_2310,In_260);
nand U2090 (N_2090,In_1804,In_718);
nor U2091 (N_2091,In_2021,In_1881);
nor U2092 (N_2092,In_302,In_2230);
nand U2093 (N_2093,In_673,In_494);
and U2094 (N_2094,In_665,In_2163);
nand U2095 (N_2095,In_1619,In_1296);
nand U2096 (N_2096,In_797,In_652);
and U2097 (N_2097,In_68,In_830);
or U2098 (N_2098,In_661,In_750);
nor U2099 (N_2099,In_1970,In_1859);
nand U2100 (N_2100,In_771,In_9);
xnor U2101 (N_2101,In_1404,In_1358);
or U2102 (N_2102,In_1830,In_974);
nor U2103 (N_2103,In_952,In_1035);
nor U2104 (N_2104,In_2318,In_1881);
xor U2105 (N_2105,In_637,In_2377);
nor U2106 (N_2106,In_1977,In_2232);
nand U2107 (N_2107,In_1978,In_1821);
and U2108 (N_2108,In_1721,In_1756);
nor U2109 (N_2109,In_1880,In_2269);
nor U2110 (N_2110,In_1149,In_1890);
or U2111 (N_2111,In_635,In_1404);
xor U2112 (N_2112,In_1077,In_2031);
and U2113 (N_2113,In_801,In_1124);
xor U2114 (N_2114,In_433,In_1158);
xor U2115 (N_2115,In_1661,In_1902);
nand U2116 (N_2116,In_2366,In_1691);
or U2117 (N_2117,In_1134,In_2128);
xnor U2118 (N_2118,In_679,In_2489);
or U2119 (N_2119,In_1064,In_2193);
xor U2120 (N_2120,In_1986,In_405);
nor U2121 (N_2121,In_2000,In_1491);
nor U2122 (N_2122,In_2285,In_425);
nand U2123 (N_2123,In_1059,In_1060);
nand U2124 (N_2124,In_317,In_714);
nor U2125 (N_2125,In_1108,In_1829);
xor U2126 (N_2126,In_1618,In_1105);
xnor U2127 (N_2127,In_2044,In_1695);
or U2128 (N_2128,In_364,In_1745);
xor U2129 (N_2129,In_849,In_903);
and U2130 (N_2130,In_693,In_413);
xor U2131 (N_2131,In_1637,In_181);
nand U2132 (N_2132,In_2379,In_139);
nand U2133 (N_2133,In_234,In_1666);
nand U2134 (N_2134,In_2298,In_161);
or U2135 (N_2135,In_1636,In_1297);
or U2136 (N_2136,In_2412,In_1731);
xor U2137 (N_2137,In_2178,In_2084);
xor U2138 (N_2138,In_708,In_2094);
nand U2139 (N_2139,In_1359,In_152);
and U2140 (N_2140,In_1771,In_877);
nor U2141 (N_2141,In_2228,In_954);
nor U2142 (N_2142,In_1360,In_764);
nand U2143 (N_2143,In_1932,In_841);
xnor U2144 (N_2144,In_1295,In_1888);
nor U2145 (N_2145,In_502,In_280);
nor U2146 (N_2146,In_1750,In_472);
nor U2147 (N_2147,In_1761,In_2214);
xnor U2148 (N_2148,In_136,In_1261);
or U2149 (N_2149,In_2186,In_2361);
nor U2150 (N_2150,In_827,In_1490);
xnor U2151 (N_2151,In_1873,In_544);
xnor U2152 (N_2152,In_1554,In_2192);
and U2153 (N_2153,In_1600,In_923);
or U2154 (N_2154,In_1311,In_969);
and U2155 (N_2155,In_772,In_1345);
nor U2156 (N_2156,In_2336,In_1286);
nand U2157 (N_2157,In_1788,In_1893);
and U2158 (N_2158,In_2153,In_276);
or U2159 (N_2159,In_1748,In_2364);
nand U2160 (N_2160,In_1815,In_481);
xnor U2161 (N_2161,In_1418,In_1003);
and U2162 (N_2162,In_562,In_2371);
or U2163 (N_2163,In_535,In_216);
or U2164 (N_2164,In_1319,In_257);
nor U2165 (N_2165,In_345,In_680);
xnor U2166 (N_2166,In_1695,In_578);
nand U2167 (N_2167,In_584,In_1204);
xnor U2168 (N_2168,In_351,In_1473);
nand U2169 (N_2169,In_806,In_1066);
nand U2170 (N_2170,In_582,In_552);
nor U2171 (N_2171,In_1681,In_1946);
nand U2172 (N_2172,In_869,In_1652);
xnor U2173 (N_2173,In_1925,In_329);
xor U2174 (N_2174,In_664,In_2469);
or U2175 (N_2175,In_32,In_1917);
nor U2176 (N_2176,In_1384,In_39);
and U2177 (N_2177,In_1939,In_163);
or U2178 (N_2178,In_841,In_487);
nor U2179 (N_2179,In_2446,In_516);
or U2180 (N_2180,In_2415,In_636);
nor U2181 (N_2181,In_414,In_1820);
and U2182 (N_2182,In_1042,In_1907);
xnor U2183 (N_2183,In_1552,In_1515);
xor U2184 (N_2184,In_1765,In_1048);
and U2185 (N_2185,In_1054,In_1779);
nand U2186 (N_2186,In_422,In_2353);
nand U2187 (N_2187,In_517,In_1014);
or U2188 (N_2188,In_928,In_2241);
or U2189 (N_2189,In_1421,In_1812);
nor U2190 (N_2190,In_1441,In_1980);
or U2191 (N_2191,In_825,In_2226);
or U2192 (N_2192,In_1198,In_1606);
or U2193 (N_2193,In_1774,In_485);
and U2194 (N_2194,In_335,In_1122);
or U2195 (N_2195,In_1765,In_1536);
nand U2196 (N_2196,In_774,In_2112);
and U2197 (N_2197,In_1319,In_85);
xor U2198 (N_2198,In_1409,In_1913);
nor U2199 (N_2199,In_2449,In_1069);
xnor U2200 (N_2200,In_2285,In_1018);
nand U2201 (N_2201,In_325,In_2119);
or U2202 (N_2202,In_2328,In_984);
or U2203 (N_2203,In_2369,In_2140);
nor U2204 (N_2204,In_1817,In_1144);
xor U2205 (N_2205,In_213,In_2036);
or U2206 (N_2206,In_481,In_870);
xnor U2207 (N_2207,In_200,In_2307);
nand U2208 (N_2208,In_964,In_1383);
or U2209 (N_2209,In_43,In_63);
or U2210 (N_2210,In_403,In_1543);
and U2211 (N_2211,In_1195,In_97);
and U2212 (N_2212,In_908,In_2275);
xnor U2213 (N_2213,In_1673,In_577);
nor U2214 (N_2214,In_1606,In_1131);
nor U2215 (N_2215,In_644,In_1472);
nand U2216 (N_2216,In_1166,In_203);
and U2217 (N_2217,In_455,In_382);
nor U2218 (N_2218,In_1750,In_2235);
or U2219 (N_2219,In_24,In_2433);
xnor U2220 (N_2220,In_564,In_1001);
nor U2221 (N_2221,In_1867,In_801);
nand U2222 (N_2222,In_2102,In_2394);
nor U2223 (N_2223,In_1337,In_1859);
and U2224 (N_2224,In_802,In_661);
and U2225 (N_2225,In_633,In_2285);
nand U2226 (N_2226,In_1146,In_921);
or U2227 (N_2227,In_1977,In_1371);
or U2228 (N_2228,In_677,In_1353);
nor U2229 (N_2229,In_1648,In_526);
nor U2230 (N_2230,In_1181,In_196);
xor U2231 (N_2231,In_1213,In_29);
nor U2232 (N_2232,In_1758,In_1145);
and U2233 (N_2233,In_534,In_2415);
xor U2234 (N_2234,In_165,In_345);
nor U2235 (N_2235,In_280,In_2268);
or U2236 (N_2236,In_2358,In_2157);
or U2237 (N_2237,In_838,In_695);
or U2238 (N_2238,In_1590,In_2047);
or U2239 (N_2239,In_2232,In_899);
nand U2240 (N_2240,In_1344,In_155);
and U2241 (N_2241,In_1032,In_1918);
nand U2242 (N_2242,In_546,In_345);
nand U2243 (N_2243,In_532,In_590);
nor U2244 (N_2244,In_330,In_2128);
or U2245 (N_2245,In_1422,In_432);
xor U2246 (N_2246,In_2193,In_2316);
and U2247 (N_2247,In_1251,In_542);
xor U2248 (N_2248,In_1715,In_2369);
nand U2249 (N_2249,In_1977,In_1208);
nor U2250 (N_2250,In_1819,In_1875);
nor U2251 (N_2251,In_2462,In_2253);
and U2252 (N_2252,In_2170,In_2357);
and U2253 (N_2253,In_2232,In_1644);
or U2254 (N_2254,In_71,In_2303);
nand U2255 (N_2255,In_1531,In_419);
nand U2256 (N_2256,In_1789,In_1275);
and U2257 (N_2257,In_919,In_632);
nor U2258 (N_2258,In_972,In_155);
nor U2259 (N_2259,In_790,In_1068);
nand U2260 (N_2260,In_210,In_2207);
or U2261 (N_2261,In_407,In_1683);
xnor U2262 (N_2262,In_1012,In_1078);
or U2263 (N_2263,In_2442,In_956);
xor U2264 (N_2264,In_639,In_532);
or U2265 (N_2265,In_550,In_2080);
nand U2266 (N_2266,In_1546,In_593);
xnor U2267 (N_2267,In_2439,In_2225);
xnor U2268 (N_2268,In_921,In_488);
and U2269 (N_2269,In_1108,In_644);
or U2270 (N_2270,In_512,In_1069);
nand U2271 (N_2271,In_553,In_1276);
nand U2272 (N_2272,In_2448,In_356);
and U2273 (N_2273,In_1079,In_928);
or U2274 (N_2274,In_506,In_1986);
nor U2275 (N_2275,In_1356,In_125);
and U2276 (N_2276,In_226,In_1836);
or U2277 (N_2277,In_2272,In_552);
nand U2278 (N_2278,In_1856,In_1939);
nor U2279 (N_2279,In_457,In_2125);
or U2280 (N_2280,In_803,In_280);
nor U2281 (N_2281,In_1233,In_1477);
xor U2282 (N_2282,In_144,In_1622);
or U2283 (N_2283,In_2178,In_2206);
and U2284 (N_2284,In_1850,In_1412);
nand U2285 (N_2285,In_2499,In_1000);
nand U2286 (N_2286,In_488,In_2375);
and U2287 (N_2287,In_1219,In_799);
and U2288 (N_2288,In_1123,In_2239);
nor U2289 (N_2289,In_1993,In_2228);
nor U2290 (N_2290,In_1843,In_2129);
nand U2291 (N_2291,In_1842,In_1406);
nand U2292 (N_2292,In_975,In_808);
nor U2293 (N_2293,In_1715,In_376);
nand U2294 (N_2294,In_1779,In_1790);
xor U2295 (N_2295,In_2348,In_148);
nand U2296 (N_2296,In_2176,In_1570);
nand U2297 (N_2297,In_1474,In_1000);
or U2298 (N_2298,In_1077,In_1640);
nand U2299 (N_2299,In_121,In_2321);
nand U2300 (N_2300,In_1063,In_197);
or U2301 (N_2301,In_1189,In_833);
nor U2302 (N_2302,In_1688,In_411);
xnor U2303 (N_2303,In_2166,In_929);
nand U2304 (N_2304,In_1877,In_1030);
or U2305 (N_2305,In_132,In_1300);
and U2306 (N_2306,In_610,In_1792);
nand U2307 (N_2307,In_1841,In_541);
or U2308 (N_2308,In_146,In_869);
nand U2309 (N_2309,In_1428,In_1844);
nor U2310 (N_2310,In_1992,In_1633);
nor U2311 (N_2311,In_914,In_854);
xnor U2312 (N_2312,In_265,In_1211);
nand U2313 (N_2313,In_2122,In_1456);
xnor U2314 (N_2314,In_1594,In_1494);
nand U2315 (N_2315,In_251,In_1944);
or U2316 (N_2316,In_1069,In_1406);
nor U2317 (N_2317,In_1156,In_460);
nor U2318 (N_2318,In_864,In_247);
xnor U2319 (N_2319,In_731,In_1776);
and U2320 (N_2320,In_1630,In_1706);
or U2321 (N_2321,In_957,In_1718);
nor U2322 (N_2322,In_1000,In_2372);
or U2323 (N_2323,In_2069,In_2253);
or U2324 (N_2324,In_1653,In_1997);
xnor U2325 (N_2325,In_1885,In_1332);
and U2326 (N_2326,In_2423,In_2106);
nand U2327 (N_2327,In_1432,In_1173);
nand U2328 (N_2328,In_1176,In_1118);
nor U2329 (N_2329,In_2205,In_1997);
and U2330 (N_2330,In_691,In_1606);
nand U2331 (N_2331,In_224,In_1862);
nand U2332 (N_2332,In_761,In_2088);
xnor U2333 (N_2333,In_390,In_110);
or U2334 (N_2334,In_435,In_2377);
xnor U2335 (N_2335,In_2155,In_586);
and U2336 (N_2336,In_1502,In_187);
nand U2337 (N_2337,In_488,In_1383);
and U2338 (N_2338,In_1732,In_562);
xor U2339 (N_2339,In_888,In_603);
nor U2340 (N_2340,In_830,In_1419);
or U2341 (N_2341,In_1406,In_971);
xor U2342 (N_2342,In_683,In_2118);
nor U2343 (N_2343,In_692,In_536);
nor U2344 (N_2344,In_1109,In_2372);
xnor U2345 (N_2345,In_169,In_1708);
xor U2346 (N_2346,In_1521,In_146);
xor U2347 (N_2347,In_1725,In_2333);
and U2348 (N_2348,In_798,In_2355);
or U2349 (N_2349,In_2331,In_874);
and U2350 (N_2350,In_779,In_563);
xnor U2351 (N_2351,In_2171,In_2033);
xor U2352 (N_2352,In_1671,In_1328);
or U2353 (N_2353,In_203,In_1727);
nand U2354 (N_2354,In_2485,In_2493);
nand U2355 (N_2355,In_1290,In_2158);
and U2356 (N_2356,In_1836,In_1095);
or U2357 (N_2357,In_908,In_2308);
nand U2358 (N_2358,In_975,In_149);
xor U2359 (N_2359,In_1647,In_2440);
and U2360 (N_2360,In_1423,In_870);
or U2361 (N_2361,In_1516,In_1469);
nand U2362 (N_2362,In_1220,In_863);
nor U2363 (N_2363,In_300,In_1014);
nand U2364 (N_2364,In_1797,In_750);
or U2365 (N_2365,In_662,In_2034);
and U2366 (N_2366,In_1449,In_926);
nor U2367 (N_2367,In_1617,In_150);
or U2368 (N_2368,In_954,In_979);
and U2369 (N_2369,In_1132,In_82);
nor U2370 (N_2370,In_1204,In_186);
xnor U2371 (N_2371,In_80,In_1192);
or U2372 (N_2372,In_325,In_2328);
nand U2373 (N_2373,In_2393,In_293);
and U2374 (N_2374,In_1547,In_803);
nor U2375 (N_2375,In_1349,In_858);
and U2376 (N_2376,In_1520,In_90);
or U2377 (N_2377,In_2033,In_398);
and U2378 (N_2378,In_2053,In_2383);
and U2379 (N_2379,In_678,In_1731);
nor U2380 (N_2380,In_1523,In_2204);
or U2381 (N_2381,In_1104,In_2077);
nand U2382 (N_2382,In_2288,In_448);
or U2383 (N_2383,In_1592,In_1734);
nor U2384 (N_2384,In_579,In_310);
or U2385 (N_2385,In_533,In_338);
nor U2386 (N_2386,In_1492,In_1355);
nor U2387 (N_2387,In_1245,In_1436);
nand U2388 (N_2388,In_2130,In_1373);
nand U2389 (N_2389,In_299,In_1479);
and U2390 (N_2390,In_2458,In_950);
nor U2391 (N_2391,In_1368,In_2477);
nor U2392 (N_2392,In_1904,In_1854);
xor U2393 (N_2393,In_2360,In_2157);
or U2394 (N_2394,In_920,In_112);
nand U2395 (N_2395,In_1687,In_122);
xor U2396 (N_2396,In_1422,In_1195);
xnor U2397 (N_2397,In_96,In_2319);
or U2398 (N_2398,In_1206,In_1661);
nor U2399 (N_2399,In_59,In_140);
or U2400 (N_2400,In_697,In_463);
nand U2401 (N_2401,In_930,In_1829);
xor U2402 (N_2402,In_2383,In_2104);
nand U2403 (N_2403,In_1395,In_1282);
xor U2404 (N_2404,In_537,In_41);
nand U2405 (N_2405,In_2101,In_2302);
xnor U2406 (N_2406,In_2044,In_2001);
nor U2407 (N_2407,In_579,In_2021);
and U2408 (N_2408,In_1825,In_141);
and U2409 (N_2409,In_1877,In_1098);
or U2410 (N_2410,In_407,In_1253);
xor U2411 (N_2411,In_1171,In_1020);
or U2412 (N_2412,In_503,In_2025);
nor U2413 (N_2413,In_583,In_561);
and U2414 (N_2414,In_1070,In_2035);
xor U2415 (N_2415,In_2239,In_598);
xnor U2416 (N_2416,In_838,In_546);
xnor U2417 (N_2417,In_1856,In_1269);
or U2418 (N_2418,In_398,In_1981);
or U2419 (N_2419,In_1083,In_341);
nor U2420 (N_2420,In_64,In_1689);
or U2421 (N_2421,In_724,In_600);
nor U2422 (N_2422,In_2053,In_896);
nand U2423 (N_2423,In_366,In_2399);
and U2424 (N_2424,In_387,In_2178);
and U2425 (N_2425,In_1089,In_1284);
and U2426 (N_2426,In_1693,In_230);
nand U2427 (N_2427,In_1705,In_452);
or U2428 (N_2428,In_1520,In_1562);
nand U2429 (N_2429,In_1575,In_1647);
nor U2430 (N_2430,In_1382,In_8);
and U2431 (N_2431,In_336,In_55);
and U2432 (N_2432,In_2327,In_932);
xnor U2433 (N_2433,In_542,In_871);
or U2434 (N_2434,In_297,In_1174);
xor U2435 (N_2435,In_1662,In_1266);
and U2436 (N_2436,In_148,In_328);
or U2437 (N_2437,In_701,In_1496);
nor U2438 (N_2438,In_2182,In_30);
nand U2439 (N_2439,In_2221,In_1212);
nand U2440 (N_2440,In_1395,In_1095);
nand U2441 (N_2441,In_2468,In_1346);
nor U2442 (N_2442,In_2311,In_1840);
or U2443 (N_2443,In_2244,In_614);
xor U2444 (N_2444,In_336,In_43);
and U2445 (N_2445,In_1400,In_1688);
or U2446 (N_2446,In_1583,In_2125);
and U2447 (N_2447,In_989,In_1042);
and U2448 (N_2448,In_1452,In_1353);
nor U2449 (N_2449,In_1249,In_328);
nor U2450 (N_2450,In_2016,In_1208);
or U2451 (N_2451,In_1613,In_830);
or U2452 (N_2452,In_1221,In_2137);
nor U2453 (N_2453,In_2046,In_955);
and U2454 (N_2454,In_1648,In_1198);
nor U2455 (N_2455,In_1498,In_1436);
or U2456 (N_2456,In_2380,In_2093);
nor U2457 (N_2457,In_1428,In_1532);
nor U2458 (N_2458,In_1482,In_1946);
and U2459 (N_2459,In_2330,In_1326);
xnor U2460 (N_2460,In_2477,In_2441);
nor U2461 (N_2461,In_1211,In_2267);
or U2462 (N_2462,In_767,In_2303);
and U2463 (N_2463,In_227,In_2065);
xor U2464 (N_2464,In_2175,In_1299);
and U2465 (N_2465,In_615,In_1347);
nand U2466 (N_2466,In_2326,In_2110);
nand U2467 (N_2467,In_2319,In_171);
nor U2468 (N_2468,In_2086,In_1015);
or U2469 (N_2469,In_2027,In_216);
xor U2470 (N_2470,In_887,In_196);
xor U2471 (N_2471,In_1166,In_1604);
nor U2472 (N_2472,In_2474,In_1525);
nand U2473 (N_2473,In_1496,In_1895);
nand U2474 (N_2474,In_798,In_1621);
nand U2475 (N_2475,In_1074,In_1793);
xor U2476 (N_2476,In_367,In_2008);
nand U2477 (N_2477,In_542,In_1362);
nand U2478 (N_2478,In_1916,In_833);
or U2479 (N_2479,In_2151,In_1926);
or U2480 (N_2480,In_1498,In_1388);
nand U2481 (N_2481,In_1504,In_1087);
and U2482 (N_2482,In_2083,In_756);
xor U2483 (N_2483,In_2442,In_1842);
xor U2484 (N_2484,In_1201,In_1018);
nor U2485 (N_2485,In_1833,In_1656);
nor U2486 (N_2486,In_2098,In_2391);
or U2487 (N_2487,In_1276,In_1014);
nor U2488 (N_2488,In_1152,In_2453);
and U2489 (N_2489,In_534,In_2474);
nand U2490 (N_2490,In_10,In_2079);
or U2491 (N_2491,In_1682,In_1258);
or U2492 (N_2492,In_2429,In_418);
nor U2493 (N_2493,In_1565,In_1226);
xnor U2494 (N_2494,In_923,In_1130);
and U2495 (N_2495,In_401,In_860);
and U2496 (N_2496,In_1436,In_439);
nand U2497 (N_2497,In_1316,In_248);
xor U2498 (N_2498,In_915,In_1283);
or U2499 (N_2499,In_467,In_437);
and U2500 (N_2500,N_303,N_2324);
and U2501 (N_2501,N_1650,N_681);
and U2502 (N_2502,N_2250,N_1518);
xor U2503 (N_2503,N_985,N_1005);
and U2504 (N_2504,N_2355,N_119);
or U2505 (N_2505,N_2288,N_1155);
or U2506 (N_2506,N_798,N_37);
or U2507 (N_2507,N_2212,N_1078);
or U2508 (N_2508,N_2376,N_2310);
nor U2509 (N_2509,N_1238,N_1751);
or U2510 (N_2510,N_520,N_598);
nor U2511 (N_2511,N_478,N_941);
nand U2512 (N_2512,N_1033,N_1489);
and U2513 (N_2513,N_1815,N_2369);
or U2514 (N_2514,N_2478,N_1353);
xor U2515 (N_2515,N_2373,N_674);
nand U2516 (N_2516,N_559,N_2088);
xnor U2517 (N_2517,N_99,N_51);
nand U2518 (N_2518,N_2239,N_318);
or U2519 (N_2519,N_626,N_169);
nand U2520 (N_2520,N_352,N_515);
nand U2521 (N_2521,N_1955,N_963);
nand U2522 (N_2522,N_368,N_1121);
xnor U2523 (N_2523,N_1800,N_2110);
or U2524 (N_2524,N_2447,N_469);
nor U2525 (N_2525,N_1550,N_886);
xor U2526 (N_2526,N_347,N_2096);
nand U2527 (N_2527,N_842,N_1529);
nor U2528 (N_2528,N_2125,N_2368);
xnor U2529 (N_2529,N_1417,N_7);
and U2530 (N_2530,N_1723,N_1652);
and U2531 (N_2531,N_2022,N_1185);
and U2532 (N_2532,N_821,N_1318);
nor U2533 (N_2533,N_526,N_1705);
and U2534 (N_2534,N_808,N_2344);
nand U2535 (N_2535,N_498,N_2409);
nor U2536 (N_2536,N_796,N_760);
or U2537 (N_2537,N_2488,N_2198);
and U2538 (N_2538,N_1180,N_1835);
and U2539 (N_2539,N_2177,N_2440);
nor U2540 (N_2540,N_1172,N_1854);
xor U2541 (N_2541,N_1971,N_1767);
nand U2542 (N_2542,N_1341,N_115);
nand U2543 (N_2543,N_1631,N_841);
or U2544 (N_2544,N_1623,N_2282);
nand U2545 (N_2545,N_1153,N_1739);
and U2546 (N_2546,N_2021,N_1345);
or U2547 (N_2547,N_656,N_1308);
and U2548 (N_2548,N_191,N_1612);
and U2549 (N_2549,N_969,N_1448);
and U2550 (N_2550,N_256,N_132);
xor U2551 (N_2551,N_94,N_793);
or U2552 (N_2552,N_953,N_1268);
nor U2553 (N_2553,N_732,N_903);
or U2554 (N_2554,N_447,N_121);
and U2555 (N_2555,N_1614,N_1899);
and U2556 (N_2556,N_1516,N_2422);
xnor U2557 (N_2557,N_390,N_788);
nor U2558 (N_2558,N_822,N_1259);
xor U2559 (N_2559,N_2170,N_1405);
nor U2560 (N_2560,N_1343,N_2001);
xnor U2561 (N_2561,N_2060,N_2487);
or U2562 (N_2562,N_1449,N_1936);
or U2563 (N_2563,N_1289,N_1138);
or U2564 (N_2564,N_1775,N_1560);
nor U2565 (N_2565,N_1179,N_66);
nand U2566 (N_2566,N_2073,N_1588);
xnor U2567 (N_2567,N_262,N_1726);
and U2568 (N_2568,N_48,N_301);
and U2569 (N_2569,N_255,N_646);
xnor U2570 (N_2570,N_464,N_1194);
or U2571 (N_2571,N_769,N_415);
nor U2572 (N_2572,N_1535,N_906);
or U2573 (N_2573,N_1748,N_600);
nor U2574 (N_2574,N_1821,N_1255);
or U2575 (N_2575,N_1166,N_2009);
or U2576 (N_2576,N_1544,N_1036);
and U2577 (N_2577,N_25,N_652);
nand U2578 (N_2578,N_828,N_2240);
nor U2579 (N_2579,N_980,N_1670);
xnor U2580 (N_2580,N_1840,N_1896);
nand U2581 (N_2581,N_2248,N_2492);
nand U2582 (N_2582,N_1541,N_1611);
xnor U2583 (N_2583,N_2499,N_1870);
xor U2584 (N_2584,N_2237,N_706);
nand U2585 (N_2585,N_649,N_1431);
nor U2586 (N_2586,N_915,N_166);
nand U2587 (N_2587,N_2404,N_89);
and U2588 (N_2588,N_1037,N_1380);
or U2589 (N_2589,N_845,N_581);
and U2590 (N_2590,N_235,N_1260);
nand U2591 (N_2591,N_2421,N_1659);
or U2592 (N_2592,N_1433,N_1591);
nand U2593 (N_2593,N_183,N_42);
or U2594 (N_2594,N_1864,N_217);
xor U2595 (N_2595,N_203,N_727);
xnor U2596 (N_2596,N_533,N_2143);
nor U2597 (N_2597,N_468,N_370);
nor U2598 (N_2598,N_647,N_2062);
xor U2599 (N_2599,N_1646,N_1326);
nor U2600 (N_2600,N_1735,N_445);
or U2601 (N_2601,N_1359,N_1447);
or U2602 (N_2602,N_2216,N_2093);
nand U2603 (N_2603,N_2168,N_2393);
xnor U2604 (N_2604,N_297,N_2272);
or U2605 (N_2605,N_1609,N_1104);
nor U2606 (N_2606,N_504,N_146);
xnor U2607 (N_2607,N_1182,N_1630);
nor U2608 (N_2608,N_2238,N_1527);
nor U2609 (N_2609,N_2337,N_429);
and U2610 (N_2610,N_1521,N_46);
or U2611 (N_2611,N_344,N_1797);
nand U2612 (N_2612,N_1437,N_1025);
and U2613 (N_2613,N_2194,N_2446);
or U2614 (N_2614,N_147,N_1613);
and U2615 (N_2615,N_112,N_438);
nor U2616 (N_2616,N_2327,N_1910);
or U2617 (N_2617,N_1214,N_313);
or U2618 (N_2618,N_157,N_1678);
and U2619 (N_2619,N_59,N_2275);
or U2620 (N_2620,N_2353,N_852);
nand U2621 (N_2621,N_2121,N_1388);
or U2622 (N_2622,N_215,N_2476);
or U2623 (N_2623,N_230,N_2006);
nor U2624 (N_2624,N_2289,N_1070);
and U2625 (N_2625,N_1196,N_1265);
or U2626 (N_2626,N_1770,N_1965);
and U2627 (N_2627,N_1200,N_1615);
or U2628 (N_2628,N_630,N_596);
nor U2629 (N_2629,N_1998,N_1158);
or U2630 (N_2630,N_1204,N_2114);
nor U2631 (N_2631,N_16,N_20);
xor U2632 (N_2632,N_2280,N_994);
and U2633 (N_2633,N_2158,N_1993);
nand U2634 (N_2634,N_1974,N_1366);
xnor U2635 (N_2635,N_1703,N_509);
nand U2636 (N_2636,N_864,N_87);
nor U2637 (N_2637,N_1410,N_2196);
and U2638 (N_2638,N_323,N_759);
or U2639 (N_2639,N_1892,N_584);
xnor U2640 (N_2640,N_420,N_1378);
and U2641 (N_2641,N_1583,N_1634);
or U2642 (N_2642,N_333,N_1478);
and U2643 (N_2643,N_1243,N_618);
or U2644 (N_2644,N_1576,N_1163);
and U2645 (N_2645,N_1118,N_668);
and U2646 (N_2646,N_2396,N_1487);
nand U2647 (N_2647,N_1868,N_1392);
or U2648 (N_2648,N_529,N_2258);
or U2649 (N_2649,N_1977,N_627);
or U2650 (N_2650,N_439,N_314);
and U2651 (N_2651,N_2483,N_1917);
xnor U2652 (N_2652,N_1708,N_371);
nor U2653 (N_2653,N_1477,N_1444);
nor U2654 (N_2654,N_718,N_1212);
xnor U2655 (N_2655,N_1768,N_1465);
and U2656 (N_2656,N_862,N_1334);
xnor U2657 (N_2657,N_2246,N_2261);
xor U2658 (N_2658,N_856,N_180);
nor U2659 (N_2659,N_1125,N_1696);
and U2660 (N_2660,N_1428,N_446);
xnor U2661 (N_2661,N_699,N_1666);
xor U2662 (N_2662,N_340,N_1145);
xnor U2663 (N_2663,N_1862,N_1842);
xor U2664 (N_2664,N_1788,N_1024);
nand U2665 (N_2665,N_1566,N_1371);
nand U2666 (N_2666,N_461,N_1173);
nand U2667 (N_2667,N_560,N_2103);
and U2668 (N_2668,N_1843,N_477);
and U2669 (N_2669,N_1504,N_847);
or U2670 (N_2670,N_155,N_1450);
nand U2671 (N_2671,N_1498,N_551);
xnor U2672 (N_2672,N_1873,N_1803);
or U2673 (N_2673,N_2406,N_1783);
or U2674 (N_2674,N_1397,N_1727);
nand U2675 (N_2675,N_624,N_1745);
or U2676 (N_2676,N_2397,N_810);
and U2677 (N_2677,N_41,N_1299);
or U2678 (N_2678,N_1990,N_2226);
nor U2679 (N_2679,N_827,N_1338);
or U2680 (N_2680,N_1470,N_761);
xnor U2681 (N_2681,N_1658,N_372);
nand U2682 (N_2682,N_2047,N_518);
xor U2683 (N_2683,N_939,N_1324);
nand U2684 (N_2684,N_1097,N_1963);
or U2685 (N_2685,N_1314,N_790);
nand U2686 (N_2686,N_224,N_547);
xor U2687 (N_2687,N_825,N_2259);
nor U2688 (N_2688,N_1635,N_36);
nand U2689 (N_2689,N_399,N_1626);
and U2690 (N_2690,N_1301,N_1344);
nor U2691 (N_2691,N_654,N_265);
nand U2692 (N_2692,N_1556,N_936);
and U2693 (N_2693,N_1710,N_558);
nor U2694 (N_2694,N_752,N_1459);
and U2695 (N_2695,N_250,N_1045);
nand U2696 (N_2696,N_252,N_909);
nand U2697 (N_2697,N_33,N_164);
or U2698 (N_2698,N_1011,N_1589);
or U2699 (N_2699,N_385,N_2140);
or U2700 (N_2700,N_1628,N_24);
nor U2701 (N_2701,N_2438,N_1075);
nor U2702 (N_2702,N_2274,N_454);
nor U2703 (N_2703,N_1510,N_400);
xnor U2704 (N_2704,N_2350,N_1547);
and U2705 (N_2705,N_640,N_1230);
nand U2706 (N_2706,N_588,N_156);
nand U2707 (N_2707,N_615,N_1931);
or U2708 (N_2708,N_2025,N_1453);
nor U2709 (N_2709,N_182,N_108);
xnor U2710 (N_2710,N_2020,N_197);
xor U2711 (N_2711,N_643,N_660);
nand U2712 (N_2712,N_290,N_979);
nand U2713 (N_2713,N_1831,N_1199);
nand U2714 (N_2714,N_218,N_67);
or U2715 (N_2715,N_337,N_1575);
nor U2716 (N_2716,N_2149,N_103);
nor U2717 (N_2717,N_667,N_2081);
nand U2718 (N_2718,N_809,N_1016);
or U2719 (N_2719,N_1935,N_1622);
xor U2720 (N_2720,N_1570,N_925);
and U2721 (N_2721,N_2163,N_64);
or U2722 (N_2722,N_1536,N_234);
or U2723 (N_2723,N_1606,N_2308);
and U2724 (N_2724,N_1240,N_1332);
and U2725 (N_2725,N_432,N_1164);
and U2726 (N_2726,N_1539,N_1534);
and U2727 (N_2727,N_8,N_2122);
nor U2728 (N_2728,N_1916,N_1773);
or U2729 (N_2729,N_1406,N_1063);
xor U2730 (N_2730,N_1056,N_2144);
xnor U2731 (N_2731,N_2207,N_1485);
xor U2732 (N_2732,N_677,N_1123);
nor U2733 (N_2733,N_2391,N_311);
xor U2734 (N_2734,N_2323,N_1330);
nor U2735 (N_2735,N_1643,N_2162);
nand U2736 (N_2736,N_1430,N_720);
nand U2737 (N_2737,N_834,N_1017);
and U2738 (N_2738,N_1263,N_848);
and U2739 (N_2739,N_1262,N_1673);
xor U2740 (N_2740,N_2070,N_2413);
or U2741 (N_2741,N_383,N_875);
nand U2742 (N_2742,N_1236,N_2039);
nand U2743 (N_2743,N_1227,N_872);
nand U2744 (N_2744,N_516,N_136);
nand U2745 (N_2745,N_525,N_916);
or U2746 (N_2746,N_1595,N_353);
xnor U2747 (N_2747,N_1718,N_927);
and U2748 (N_2748,N_2235,N_733);
or U2749 (N_2749,N_1348,N_2416);
or U2750 (N_2750,N_359,N_1554);
or U2751 (N_2751,N_1632,N_416);
or U2752 (N_2752,N_641,N_201);
and U2753 (N_2753,N_1007,N_2042);
or U2754 (N_2754,N_871,N_1960);
and U2755 (N_2755,N_1789,N_958);
xnor U2756 (N_2756,N_2155,N_675);
xnor U2757 (N_2757,N_1151,N_700);
and U2758 (N_2758,N_418,N_1538);
and U2759 (N_2759,N_657,N_2470);
and U2760 (N_2760,N_2467,N_1697);
xnor U2761 (N_2761,N_709,N_1598);
and U2762 (N_2762,N_830,N_1372);
xor U2763 (N_2763,N_1969,N_1526);
nor U2764 (N_2764,N_2139,N_2091);
xnor U2765 (N_2765,N_1913,N_734);
xor U2766 (N_2766,N_405,N_229);
or U2767 (N_2767,N_1169,N_1368);
or U2768 (N_2768,N_2108,N_2307);
or U2769 (N_2769,N_635,N_1711);
nor U2770 (N_2770,N_737,N_1776);
nand U2771 (N_2771,N_1493,N_145);
nand U2772 (N_2772,N_307,N_2418);
xor U2773 (N_2773,N_1225,N_1374);
nor U2774 (N_2774,N_986,N_1999);
nor U2775 (N_2775,N_482,N_72);
xnor U2776 (N_2776,N_1686,N_2490);
nand U2777 (N_2777,N_1919,N_2112);
nand U2778 (N_2778,N_1569,N_549);
xor U2779 (N_2779,N_1537,N_728);
nor U2780 (N_2780,N_736,N_437);
or U2781 (N_2781,N_1580,N_2043);
nand U2782 (N_2782,N_2400,N_1724);
and U2783 (N_2783,N_1581,N_2460);
nor U2784 (N_2784,N_1810,N_1191);
nor U2785 (N_2785,N_137,N_1655);
or U2786 (N_2786,N_680,N_611);
or U2787 (N_2787,N_1462,N_269);
xor U2788 (N_2788,N_2389,N_1687);
nor U2789 (N_2789,N_874,N_1393);
and U2790 (N_2790,N_320,N_373);
nand U2791 (N_2791,N_2375,N_2315);
and U2792 (N_2792,N_1765,N_1672);
or U2793 (N_2793,N_1205,N_2429);
and U2794 (N_2794,N_1813,N_1699);
nand U2795 (N_2795,N_2431,N_1805);
nand U2796 (N_2796,N_1725,N_1226);
or U2797 (N_2797,N_1908,N_1853);
or U2798 (N_2798,N_2102,N_263);
nor U2799 (N_2799,N_1423,N_1064);
nand U2800 (N_2800,N_159,N_1052);
or U2801 (N_2801,N_705,N_91);
nand U2802 (N_2802,N_396,N_476);
or U2803 (N_2803,N_55,N_208);
xnor U2804 (N_2804,N_1074,N_165);
and U2805 (N_2805,N_616,N_2343);
xnor U2806 (N_2806,N_86,N_757);
and U2807 (N_2807,N_329,N_1736);
or U2808 (N_2808,N_238,N_1439);
or U2809 (N_2809,N_754,N_459);
nor U2810 (N_2810,N_711,N_1080);
or U2811 (N_2811,N_1925,N_716);
xnor U2812 (N_2812,N_81,N_1716);
nand U2813 (N_2813,N_910,N_1914);
and U2814 (N_2814,N_186,N_972);
nand U2815 (N_2815,N_152,N_1340);
xnor U2816 (N_2816,N_1427,N_1738);
nand U2817 (N_2817,N_731,N_2094);
nor U2818 (N_2818,N_729,N_2281);
or U2819 (N_2819,N_2129,N_777);
nor U2820 (N_2820,N_648,N_1491);
nand U2821 (N_2821,N_687,N_712);
and U2822 (N_2822,N_623,N_1039);
and U2823 (N_2823,N_15,N_1249);
xnor U2824 (N_2824,N_1071,N_912);
xnor U2825 (N_2825,N_2420,N_111);
and U2826 (N_2826,N_1188,N_2165);
nor U2827 (N_2827,N_2301,N_1384);
and U2828 (N_2828,N_690,N_1675);
nor U2829 (N_2829,N_655,N_332);
nor U2830 (N_2830,N_2267,N_1790);
xnor U2831 (N_2831,N_682,N_1203);
nand U2832 (N_2832,N_639,N_1261);
xnor U2833 (N_2833,N_316,N_2491);
and U2834 (N_2834,N_1316,N_1975);
and U2835 (N_2835,N_2031,N_1949);
and U2836 (N_2836,N_2286,N_838);
nand U2837 (N_2837,N_1277,N_1764);
nand U2838 (N_2838,N_948,N_1664);
nand U2839 (N_2839,N_1859,N_2424);
xor U2840 (N_2840,N_349,N_1252);
nand U2841 (N_2841,N_2152,N_1046);
xnor U2842 (N_2842,N_1144,N_1545);
nor U2843 (N_2843,N_2097,N_1273);
nand U2844 (N_2844,N_695,N_1302);
and U2845 (N_2845,N_2189,N_1432);
and U2846 (N_2846,N_1293,N_2321);
nand U2847 (N_2847,N_2182,N_1654);
nand U2848 (N_2848,N_1496,N_1929);
and U2849 (N_2849,N_2331,N_2033);
nand U2850 (N_2850,N_110,N_998);
or U2851 (N_2851,N_450,N_441);
or U2852 (N_2852,N_283,N_2494);
or U2853 (N_2853,N_1210,N_2256);
nand U2854 (N_2854,N_595,N_328);
or U2855 (N_2855,N_869,N_686);
and U2856 (N_2856,N_1010,N_2298);
or U2857 (N_2857,N_1540,N_1733);
nand U2858 (N_2858,N_859,N_548);
or U2859 (N_2859,N_68,N_409);
xor U2860 (N_2860,N_343,N_943);
xor U2861 (N_2861,N_932,N_342);
and U2862 (N_2862,N_688,N_13);
or U2863 (N_2863,N_2290,N_800);
and U2864 (N_2864,N_378,N_2450);
or U2865 (N_2865,N_2383,N_486);
nand U2866 (N_2866,N_1031,N_995);
and U2867 (N_2867,N_692,N_488);
nand U2868 (N_2868,N_1375,N_1605);
nand U2869 (N_2869,N_2356,N_23);
nor U2870 (N_2870,N_277,N_122);
nor U2871 (N_2871,N_1514,N_713);
and U2872 (N_2872,N_1044,N_2489);
or U2873 (N_2873,N_1898,N_1661);
xnor U2874 (N_2874,N_497,N_877);
xnor U2875 (N_2875,N_1952,N_507);
nor U2876 (N_2876,N_501,N_211);
xnor U2877 (N_2877,N_1223,N_779);
nand U2878 (N_2878,N_1972,N_2219);
and U2879 (N_2879,N_105,N_1245);
nand U2880 (N_2880,N_950,N_1774);
and U2881 (N_2881,N_38,N_1181);
xnor U2882 (N_2882,N_1532,N_665);
nor U2883 (N_2883,N_523,N_2099);
nor U2884 (N_2884,N_1363,N_1662);
nor U2885 (N_2885,N_2179,N_19);
nor U2886 (N_2886,N_2241,N_1548);
xor U2887 (N_2887,N_1127,N_1120);
nand U2888 (N_2888,N_98,N_1246);
or U2889 (N_2889,N_740,N_2051);
nor U2890 (N_2890,N_1717,N_61);
and U2891 (N_2891,N_1481,N_2380);
xnor U2892 (N_2892,N_1331,N_1020);
and U2893 (N_2893,N_1928,N_1455);
nor U2894 (N_2894,N_1985,N_2319);
nor U2895 (N_2895,N_988,N_1844);
nand U2896 (N_2896,N_1701,N_983);
nand U2897 (N_2897,N_52,N_707);
and U2898 (N_2898,N_1440,N_173);
nand U2899 (N_2899,N_39,N_1508);
nor U2900 (N_2900,N_236,N_1306);
nor U2901 (N_2901,N_2451,N_2045);
and U2902 (N_2902,N_2195,N_1677);
xnor U2903 (N_2903,N_607,N_719);
nor U2904 (N_2904,N_921,N_1256);
nor U2905 (N_2905,N_1117,N_1869);
xor U2906 (N_2906,N_1827,N_970);
xnor U2907 (N_2907,N_1313,N_367);
or U2908 (N_2908,N_975,N_1676);
nor U2909 (N_2909,N_1795,N_1055);
and U2910 (N_2910,N_9,N_1032);
or U2911 (N_2911,N_1105,N_1746);
xor U2912 (N_2912,N_1712,N_1207);
nand U2913 (N_2913,N_1004,N_602);
xor U2914 (N_2914,N_1891,N_1412);
nand U2915 (N_2915,N_151,N_2074);
nand U2916 (N_2916,N_2167,N_2063);
or U2917 (N_2917,N_747,N_532);
or U2918 (N_2918,N_2046,N_617);
nor U2919 (N_2919,N_176,N_566);
or U2920 (N_2920,N_1415,N_2215);
or U2921 (N_2921,N_118,N_2126);
or U2922 (N_2922,N_673,N_2474);
or U2923 (N_2923,N_776,N_2065);
or U2924 (N_2924,N_604,N_1679);
nand U2925 (N_2925,N_1729,N_2077);
nand U2926 (N_2926,N_1291,N_578);
nor U2927 (N_2927,N_2263,N_1553);
and U2928 (N_2928,N_569,N_1355);
or U2929 (N_2929,N_781,N_2318);
nand U2930 (N_2930,N_1093,N_2232);
nand U2931 (N_2931,N_1793,N_2132);
nand U2932 (N_2932,N_1861,N_1441);
and U2933 (N_2933,N_2457,N_1102);
nand U2934 (N_2934,N_421,N_1012);
or U2935 (N_2935,N_88,N_2078);
nand U2936 (N_2936,N_892,N_356);
xnor U2937 (N_2937,N_774,N_1107);
and U2938 (N_2938,N_2486,N_2436);
nand U2939 (N_2939,N_1087,N_1546);
nand U2940 (N_2940,N_43,N_413);
or U2941 (N_2941,N_2221,N_448);
nor U2942 (N_2942,N_633,N_913);
xor U2943 (N_2943,N_276,N_2066);
and U2944 (N_2944,N_1244,N_2480);
nor U2945 (N_2945,N_65,N_1193);
nor U2946 (N_2946,N_484,N_653);
xnor U2947 (N_2947,N_35,N_694);
nand U2948 (N_2948,N_1407,N_404);
or U2949 (N_2949,N_1280,N_601);
xor U2950 (N_2950,N_1798,N_1709);
and U2951 (N_2951,N_2087,N_851);
xnor U2952 (N_2952,N_1177,N_907);
or U2953 (N_2953,N_503,N_483);
nor U2954 (N_2954,N_2076,N_550);
nand U2955 (N_2955,N_1351,N_1274);
nor U2956 (N_2956,N_1571,N_2026);
and U2957 (N_2957,N_1992,N_2178);
nand U2958 (N_2958,N_955,N_47);
xnor U2959 (N_2959,N_1059,N_2079);
nand U2960 (N_2960,N_381,N_2015);
xnor U2961 (N_2961,N_806,N_1513);
nor U2962 (N_2962,N_663,N_2111);
and U2963 (N_2963,N_1620,N_1694);
xnor U2964 (N_2964,N_104,N_801);
xor U2965 (N_2965,N_2305,N_519);
and U2966 (N_2966,N_1877,N_844);
xor U2967 (N_2967,N_2269,N_260);
nor U2968 (N_2968,N_1649,N_2445);
or U2969 (N_2969,N_1192,N_45);
nor U2970 (N_2970,N_1001,N_2496);
xor U2971 (N_2971,N_114,N_193);
or U2972 (N_2972,N_914,N_1939);
xor U2973 (N_2973,N_553,N_2271);
nor U2974 (N_2974,N_557,N_967);
and U2975 (N_2975,N_1888,N_487);
nand U2976 (N_2976,N_622,N_1644);
nor U2977 (N_2977,N_1799,N_1000);
nor U2978 (N_2978,N_1116,N_1515);
or U2979 (N_2979,N_2161,N_1023);
xor U2980 (N_2980,N_768,N_2090);
or U2981 (N_2981,N_1836,N_2202);
xnor U2982 (N_2982,N_1053,N_1567);
xor U2983 (N_2983,N_2037,N_567);
nand U2984 (N_2984,N_937,N_2357);
nand U2985 (N_2985,N_1483,N_325);
nand U2986 (N_2986,N_1109,N_944);
xor U2987 (N_2987,N_194,N_1275);
xnor U2988 (N_2988,N_956,N_2018);
nor U2989 (N_2989,N_113,N_393);
nor U2990 (N_2990,N_280,N_198);
xnor U2991 (N_2991,N_1988,N_1856);
nand U2992 (N_2992,N_1966,N_2294);
xnor U2993 (N_2993,N_2234,N_1336);
nand U2994 (N_2994,N_401,N_1394);
nand U2995 (N_2995,N_1241,N_1119);
and U2996 (N_2996,N_2381,N_2471);
and U2997 (N_2997,N_1257,N_949);
xor U2998 (N_2998,N_1841,N_2302);
nor U2999 (N_2999,N_605,N_21);
xor U3000 (N_3000,N_1195,N_1176);
or U3001 (N_3001,N_258,N_295);
nor U3002 (N_3002,N_964,N_2367);
and U3003 (N_3003,N_811,N_49);
nor U3004 (N_3004,N_1923,N_2201);
or U3005 (N_3005,N_977,N_1463);
or U3006 (N_3006,N_141,N_1135);
nor U3007 (N_3007,N_1160,N_931);
nor U3008 (N_3008,N_1413,N_1845);
nor U3009 (N_3009,N_1390,N_1989);
or U3010 (N_3010,N_1747,N_60);
nand U3011 (N_3011,N_452,N_552);
and U3012 (N_3012,N_1915,N_82);
nand U3013 (N_3013,N_1497,N_1134);
and U3014 (N_3014,N_69,N_984);
xor U3015 (N_3015,N_1984,N_2151);
nor U3016 (N_3016,N_693,N_1148);
nand U3017 (N_3017,N_580,N_2419);
or U3018 (N_3018,N_403,N_2303);
nor U3019 (N_3019,N_1587,N_535);
nor U3020 (N_3020,N_1784,N_1197);
nor U3021 (N_3021,N_2448,N_2055);
and U3022 (N_3022,N_563,N_1629);
nand U3023 (N_3023,N_590,N_163);
xor U3024 (N_3024,N_1681,N_228);
nor U3025 (N_3025,N_2218,N_1713);
or U3026 (N_3026,N_174,N_1579);
nand U3027 (N_3027,N_2316,N_2200);
and U3028 (N_3028,N_846,N_2137);
nor U3029 (N_3029,N_742,N_1731);
nand U3030 (N_3030,N_397,N_435);
nand U3031 (N_3031,N_1286,N_457);
nor U3032 (N_3032,N_1253,N_2402);
and U3033 (N_3033,N_1954,N_1389);
xor U3034 (N_3034,N_1584,N_882);
xnor U3035 (N_3035,N_1596,N_1607);
nor U3036 (N_3036,N_1633,N_453);
nor U3037 (N_3037,N_1346,N_1271);
nand U3038 (N_3038,N_2224,N_1174);
nand U3039 (N_3039,N_574,N_2329);
and U3040 (N_3040,N_1749,N_298);
nor U3041 (N_3041,N_481,N_2101);
nand U3042 (N_3042,N_1013,N_1980);
and U3043 (N_3043,N_2192,N_2386);
xnor U3044 (N_3044,N_1617,N_1543);
nand U3045 (N_3045,N_1250,N_2186);
xor U3046 (N_3046,N_540,N_1752);
or U3047 (N_3047,N_703,N_1691);
or U3048 (N_3048,N_1549,N_1754);
nand U3049 (N_3049,N_947,N_310);
nor U3050 (N_3050,N_1771,N_213);
and U3051 (N_3051,N_794,N_1221);
and U3052 (N_3052,N_1582,N_918);
xnor U3053 (N_3053,N_29,N_2325);
or U3054 (N_3054,N_27,N_1517);
xnor U3055 (N_3055,N_2003,N_30);
or U3056 (N_3056,N_527,N_2222);
xor U3057 (N_3057,N_243,N_2333);
nor U3058 (N_3058,N_896,N_1402);
nor U3059 (N_3059,N_860,N_586);
xnor U3060 (N_3060,N_392,N_375);
nor U3061 (N_3061,N_335,N_109);
nor U3062 (N_3062,N_2415,N_582);
and U3063 (N_3063,N_2395,N_1944);
xor U3064 (N_3064,N_162,N_222);
xor U3065 (N_3065,N_2257,N_2128);
nor U3066 (N_3066,N_339,N_2306);
or U3067 (N_3067,N_1298,N_1295);
or U3068 (N_3068,N_2214,N_456);
xnor U3069 (N_3069,N_2169,N_139);
xnor U3070 (N_3070,N_2203,N_1466);
nand U3071 (N_3071,N_1342,N_2159);
xnor U3072 (N_3072,N_2228,N_289);
nor U3073 (N_3073,N_664,N_539);
nand U3074 (N_3074,N_1068,N_645);
xnor U3075 (N_3075,N_1700,N_2085);
or U3076 (N_3076,N_717,N_1141);
nor U3077 (N_3077,N_1851,N_1222);
nand U3078 (N_3078,N_1884,N_2233);
nand U3079 (N_3079,N_899,N_1152);
xnor U3080 (N_3080,N_1715,N_1616);
nor U3081 (N_3081,N_829,N_2285);
xnor U3082 (N_3082,N_1577,N_2131);
nand U3083 (N_3083,N_725,N_1471);
nand U3084 (N_3084,N_1401,N_2390);
xnor U3085 (N_3085,N_2459,N_1801);
xor U3086 (N_3086,N_2387,N_1284);
nand U3087 (N_3087,N_1420,N_154);
xor U3088 (N_3088,N_573,N_2057);
and U3089 (N_3089,N_571,N_2370);
nor U3090 (N_3090,N_989,N_2292);
xnor U3091 (N_3091,N_2401,N_1647);
xnor U3092 (N_3092,N_300,N_1041);
or U3093 (N_3093,N_1435,N_2273);
nor U3094 (N_3094,N_1034,N_1624);
or U3095 (N_3095,N_2084,N_175);
or U3096 (N_3096,N_2069,N_1834);
xnor U3097 (N_3097,N_50,N_264);
or U3098 (N_3098,N_1573,N_221);
nor U3099 (N_3099,N_366,N_158);
nor U3100 (N_3100,N_704,N_1668);
nand U3101 (N_3101,N_1356,N_2209);
xor U3102 (N_3102,N_1695,N_826);
and U3103 (N_3103,N_1132,N_90);
or U3104 (N_3104,N_1015,N_1290);
nor U3105 (N_3105,N_974,N_2453);
and U3106 (N_3106,N_1885,N_2034);
and U3107 (N_3107,N_1889,N_904);
or U3108 (N_3108,N_167,N_556);
nand U3109 (N_3109,N_784,N_678);
or U3110 (N_3110,N_1436,N_1822);
and U3111 (N_3111,N_374,N_270);
and U3112 (N_3112,N_93,N_749);
xnor U3113 (N_3113,N_1552,N_148);
and U3114 (N_3114,N_942,N_795);
or U3115 (N_3115,N_2107,N_436);
and U3116 (N_3116,N_267,N_782);
nor U3117 (N_3117,N_2243,N_765);
or U3118 (N_3118,N_2468,N_517);
and U3119 (N_3119,N_1669,N_2231);
xor U3120 (N_3120,N_2035,N_58);
xor U3121 (N_3121,N_1426,N_1706);
and U3122 (N_3122,N_2495,N_766);
nor U3123 (N_3123,N_524,N_952);
and U3124 (N_3124,N_2268,N_505);
xnor U3125 (N_3125,N_2029,N_1464);
and U3126 (N_3126,N_1641,N_1874);
nor U3127 (N_3127,N_358,N_1021);
nand U3128 (N_3128,N_1317,N_1186);
or U3129 (N_3129,N_2276,N_2314);
xnor U3130 (N_3130,N_417,N_2142);
nor U3131 (N_3131,N_1796,N_888);
xor U3132 (N_3132,N_2399,N_1918);
xor U3133 (N_3133,N_2105,N_576);
and U3134 (N_3134,N_2408,N_1114);
xor U3135 (N_3135,N_990,N_1008);
and U3136 (N_3136,N_2054,N_1320);
xnor U3137 (N_3137,N_107,N_572);
and U3138 (N_3138,N_466,N_272);
nand U3139 (N_3139,N_758,N_908);
nor U3140 (N_3140,N_101,N_1398);
or U3141 (N_3141,N_77,N_1802);
nor U3142 (N_3142,N_1101,N_160);
nand U3143 (N_3143,N_1335,N_423);
xnor U3144 (N_3144,N_962,N_178);
or U3145 (N_3145,N_933,N_676);
nand U3146 (N_3146,N_968,N_1364);
or U3147 (N_3147,N_406,N_127);
nand U3148 (N_3148,N_976,N_723);
xor U3149 (N_3149,N_982,N_1347);
nor U3150 (N_3150,N_1894,N_510);
nor U3151 (N_3151,N_1930,N_1882);
and U3152 (N_3152,N_1395,N_1867);
nor U3153 (N_3153,N_1294,N_2064);
nor U3154 (N_3154,N_74,N_1086);
or U3155 (N_3155,N_209,N_386);
or U3156 (N_3156,N_44,N_1325);
nor U3157 (N_3157,N_204,N_1461);
or U3158 (N_3158,N_959,N_1339);
or U3159 (N_3159,N_1111,N_1809);
nor U3160 (N_3160,N_1714,N_1385);
nor U3161 (N_3161,N_895,N_181);
nand U3162 (N_3162,N_1599,N_473);
and U3163 (N_3163,N_1136,N_783);
xnor U3164 (N_3164,N_853,N_1737);
nor U3165 (N_3165,N_2469,N_1637);
xor U3166 (N_3166,N_818,N_879);
and U3167 (N_3167,N_1947,N_1829);
nand U3168 (N_3168,N_669,N_1905);
nand U3169 (N_3169,N_1996,N_2184);
or U3170 (N_3170,N_1542,N_1211);
nand U3171 (N_3171,N_1379,N_1830);
and U3172 (N_3172,N_661,N_636);
or U3173 (N_3173,N_1565,N_1076);
or U3174 (N_3174,N_422,N_1772);
and U3175 (N_3175,N_940,N_2378);
and U3176 (N_3176,N_6,N_2210);
nor U3177 (N_3177,N_1400,N_511);
xnor U3178 (N_3178,N_537,N_1458);
xor U3179 (N_3179,N_599,N_1759);
xnor U3180 (N_3180,N_2465,N_2147);
nor U3181 (N_3181,N_5,N_724);
and U3182 (N_3182,N_350,N_568);
and U3183 (N_3183,N_331,N_642);
nand U3184 (N_3184,N_2430,N_1171);
nor U3185 (N_3185,N_2245,N_2141);
xnor U3186 (N_3186,N_1365,N_2036);
nor U3187 (N_3187,N_2106,N_889);
or U3188 (N_3188,N_2145,N_2156);
nand U3189 (N_3189,N_1264,N_85);
xnor U3190 (N_3190,N_268,N_1886);
and U3191 (N_3191,N_144,N_394);
and U3192 (N_3192,N_18,N_2254);
xor U3193 (N_3193,N_2384,N_1247);
nand U3194 (N_3194,N_1920,N_1707);
nand U3195 (N_3195,N_522,N_701);
xor U3196 (N_3196,N_2452,N_1962);
xor U3197 (N_3197,N_1585,N_1030);
xor U3198 (N_3198,N_945,N_254);
and U3199 (N_3199,N_2411,N_1040);
nor U3200 (N_3200,N_837,N_80);
nand U3201 (N_3201,N_1893,N_628);
nor U3202 (N_3202,N_1826,N_1807);
or U3203 (N_3203,N_1533,N_128);
or U3204 (N_3204,N_2403,N_2164);
or U3205 (N_3205,N_190,N_1865);
nor U3206 (N_3206,N_1476,N_2109);
xnor U3207 (N_3207,N_1901,N_632);
xor U3208 (N_3208,N_207,N_992);
nor U3209 (N_3209,N_1422,N_1358);
nand U3210 (N_3210,N_273,N_1645);
and U3211 (N_3211,N_410,N_1309);
nor U3212 (N_3212,N_75,N_1610);
xnor U3213 (N_3213,N_1467,N_321);
and U3214 (N_3214,N_1740,N_1239);
nand U3215 (N_3215,N_2287,N_2358);
or U3216 (N_3216,N_492,N_419);
nand U3217 (N_3217,N_1112,N_1049);
xor U3218 (N_3218,N_923,N_1297);
xor U3219 (N_3219,N_1603,N_129);
or U3220 (N_3220,N_1572,N_1561);
nand U3221 (N_3221,N_131,N_1228);
xnor U3222 (N_3222,N_1551,N_1354);
and U3223 (N_3223,N_1147,N_751);
or U3224 (N_3224,N_341,N_1029);
or U3225 (N_3225,N_890,N_1251);
nand U3226 (N_3226,N_2270,N_2127);
or U3227 (N_3227,N_135,N_735);
nand U3228 (N_3228,N_541,N_2174);
xor U3229 (N_3229,N_965,N_2089);
nor U3230 (N_3230,N_651,N_1213);
nor U3231 (N_3231,N_1073,N_2493);
or U3232 (N_3232,N_1943,N_1557);
xor U3233 (N_3233,N_1206,N_629);
or U3234 (N_3234,N_245,N_32);
or U3235 (N_3235,N_2188,N_772);
nand U3236 (N_3236,N_1067,N_2100);
xor U3237 (N_3237,N_2364,N_2392);
or U3238 (N_3238,N_1942,N_2052);
nand U3239 (N_3239,N_840,N_1982);
nor U3240 (N_3240,N_1806,N_1756);
nand U3241 (N_3241,N_816,N_1103);
or U3242 (N_3242,N_444,N_324);
nor U3243 (N_3243,N_603,N_2426);
and U3244 (N_3244,N_2098,N_411);
xnor U3245 (N_3245,N_1184,N_2095);
or U3246 (N_3246,N_2136,N_1474);
xor U3247 (N_3247,N_770,N_2423);
nor U3248 (N_3248,N_1229,N_1946);
nand U3249 (N_3249,N_996,N_62);
and U3250 (N_3250,N_1369,N_184);
nor U3251 (N_3251,N_2362,N_721);
nand U3252 (N_3252,N_1593,N_843);
nor U3253 (N_3253,N_1502,N_2173);
nand U3254 (N_3254,N_1048,N_427);
xnor U3255 (N_3255,N_1209,N_249);
or U3256 (N_3256,N_1162,N_1625);
or U3257 (N_3257,N_1983,N_2071);
or U3258 (N_3258,N_819,N_867);
or U3259 (N_3259,N_935,N_1322);
and U3260 (N_3260,N_594,N_142);
or U3261 (N_3261,N_1242,N_451);
and U3262 (N_3262,N_1501,N_1373);
nand U3263 (N_3263,N_2072,N_1656);
xnor U3264 (N_3264,N_1887,N_291);
and U3265 (N_3265,N_1311,N_542);
xnor U3266 (N_3266,N_1600,N_824);
xnor U3267 (N_3267,N_1006,N_1702);
xnor U3268 (N_3268,N_426,N_1077);
and U3269 (N_3269,N_2010,N_2252);
nor U3270 (N_3270,N_2197,N_1051);
nor U3271 (N_3271,N_1098,N_1932);
nor U3272 (N_3272,N_1846,N_2019);
nand U3273 (N_3273,N_2116,N_1421);
nor U3274 (N_3274,N_1578,N_1875);
xnor U3275 (N_3275,N_1505,N_748);
nand U3276 (N_3276,N_1137,N_2040);
or U3277 (N_3277,N_402,N_565);
xor U3278 (N_3278,N_855,N_917);
and U3279 (N_3279,N_741,N_2264);
xnor U3280 (N_3280,N_534,N_70);
nand U3281 (N_3281,N_946,N_1900);
xnor U3282 (N_3282,N_407,N_266);
nand U3283 (N_3283,N_1159,N_1860);
nand U3284 (N_3284,N_330,N_1961);
or U3285 (N_3285,N_884,N_433);
and U3286 (N_3286,N_858,N_1909);
nand U3287 (N_3287,N_619,N_1953);
nand U3288 (N_3288,N_1857,N_1321);
nor U3289 (N_3289,N_1352,N_143);
nand U3290 (N_3290,N_762,N_2120);
nand U3291 (N_3291,N_2008,N_1978);
and U3292 (N_3292,N_697,N_1763);
nand U3293 (N_3293,N_1512,N_2115);
and U3294 (N_3294,N_1079,N_1956);
xnor U3295 (N_3295,N_2083,N_95);
or U3296 (N_3296,N_1639,N_924);
nor U3297 (N_3297,N_1520,N_1667);
xnor U3298 (N_3298,N_84,N_1113);
nor U3299 (N_3299,N_885,N_1558);
or U3300 (N_3300,N_225,N_1208);
or U3301 (N_3301,N_56,N_1224);
or U3302 (N_3302,N_1927,N_2277);
or U3303 (N_3303,N_1941,N_1602);
nor U3304 (N_3304,N_2092,N_465);
or U3305 (N_3305,N_170,N_614);
and U3306 (N_3306,N_780,N_2317);
nand U3307 (N_3307,N_279,N_1528);
nand U3308 (N_3308,N_1133,N_2181);
nor U3309 (N_3309,N_804,N_1559);
nand U3310 (N_3310,N_1814,N_177);
nand U3311 (N_3311,N_2032,N_1220);
or U3312 (N_3312,N_1912,N_2148);
xor U3313 (N_3313,N_1060,N_1108);
xor U3314 (N_3314,N_231,N_919);
and U3315 (N_3315,N_1457,N_1175);
nand U3316 (N_3316,N_561,N_1638);
or U3317 (N_3317,N_854,N_894);
nand U3318 (N_3318,N_1126,N_2299);
nand U3319 (N_3319,N_1880,N_1376);
and U3320 (N_3320,N_2185,N_1750);
or U3321 (N_3321,N_216,N_514);
nor U3322 (N_3322,N_2227,N_2374);
nor U3323 (N_3323,N_14,N_2193);
nor U3324 (N_3324,N_1621,N_1035);
or U3325 (N_3325,N_2472,N_1110);
xnor U3326 (N_3326,N_1054,N_2366);
or U3327 (N_3327,N_361,N_696);
or U3328 (N_3328,N_1362,N_1387);
nand U3329 (N_3329,N_1276,N_1642);
or U3330 (N_3330,N_1769,N_857);
nand U3331 (N_3331,N_2482,N_531);
nor U3332 (N_3332,N_389,N_1131);
and U3333 (N_3333,N_2191,N_1494);
xor U3334 (N_3334,N_2385,N_1315);
xnor U3335 (N_3335,N_2005,N_237);
nand U3336 (N_3336,N_1704,N_708);
or U3337 (N_3337,N_833,N_1081);
nor U3338 (N_3338,N_2172,N_738);
nor U3339 (N_3339,N_1486,N_2497);
nor U3340 (N_3340,N_799,N_2253);
and U3341 (N_3341,N_2278,N_179);
xnor U3342 (N_3342,N_187,N_1312);
nor U3343 (N_3343,N_312,N_930);
and U3344 (N_3344,N_360,N_666);
nor U3345 (N_3345,N_336,N_502);
nor U3346 (N_3346,N_2291,N_1069);
xor U3347 (N_3347,N_1484,N_2176);
nor U3348 (N_3348,N_2335,N_2427);
nor U3349 (N_3349,N_1926,N_442);
or U3350 (N_3350,N_315,N_430);
nor U3351 (N_3351,N_282,N_999);
nor U3352 (N_3352,N_1525,N_1660);
nor U3353 (N_3353,N_1879,N_1762);
xnor U3354 (N_3354,N_1933,N_778);
nor U3355 (N_3355,N_1468,N_662);
xnor U3356 (N_3356,N_891,N_863);
and U3357 (N_3357,N_658,N_1636);
xnor U3358 (N_3358,N_881,N_319);
nand U3359 (N_3359,N_898,N_1088);
xnor U3360 (N_3360,N_1719,N_1812);
or U3361 (N_3361,N_309,N_2041);
xor U3362 (N_3362,N_1734,N_1043);
nand U3363 (N_3363,N_1149,N_1418);
nand U3364 (N_3364,N_1743,N_412);
and U3365 (N_3365,N_1452,N_587);
or U3366 (N_3366,N_545,N_345);
xnor U3367 (N_3367,N_2334,N_866);
or U3368 (N_3368,N_2223,N_97);
nor U3369 (N_3369,N_1456,N_1042);
nand U3370 (N_3370,N_911,N_495);
nor U3371 (N_3371,N_878,N_1663);
or U3372 (N_3372,N_1028,N_2410);
nor U3373 (N_3373,N_1488,N_1142);
xnor U3374 (N_3374,N_1511,N_278);
xnor U3375 (N_3375,N_583,N_1479);
or U3376 (N_3376,N_1590,N_1816);
xnor U3377 (N_3377,N_388,N_1732);
and U3378 (N_3378,N_870,N_1876);
nand U3379 (N_3379,N_233,N_1777);
xnor U3380 (N_3380,N_192,N_2439);
xor U3381 (N_3381,N_247,N_1791);
nand U3382 (N_3382,N_1266,N_739);
nand U3383 (N_3383,N_902,N_1269);
and U3384 (N_3384,N_608,N_391);
nor U3385 (N_3385,N_512,N_2014);
nor U3386 (N_3386,N_813,N_2432);
or U3387 (N_3387,N_960,N_2016);
and U3388 (N_3388,N_2086,N_2477);
xnor U3389 (N_3389,N_650,N_613);
and U3390 (N_3390,N_536,N_1755);
and U3391 (N_3391,N_1608,N_577);
nor U3392 (N_3392,N_1099,N_1409);
nor U3393 (N_3393,N_1597,N_2048);
nand U3394 (N_3394,N_2326,N_294);
and U3395 (N_3395,N_2135,N_1360);
and U3396 (N_3396,N_900,N_634);
or U3397 (N_3397,N_865,N_1414);
nor U3398 (N_3398,N_1089,N_1248);
or U3399 (N_3399,N_2428,N_1720);
xnor U3400 (N_3400,N_1530,N_638);
nand U3401 (N_3401,N_2328,N_261);
nor U3402 (N_3402,N_440,N_1657);
and U3403 (N_3403,N_756,N_961);
nand U3404 (N_3404,N_2498,N_1047);
or U3405 (N_3405,N_2360,N_644);
xor U3406 (N_3406,N_2382,N_382);
nor U3407 (N_3407,N_12,N_2044);
xnor U3408 (N_3408,N_1187,N_538);
and U3409 (N_3409,N_2304,N_1922);
nand U3410 (N_3410,N_555,N_1818);
and U3411 (N_3411,N_1948,N_2229);
and U3412 (N_3412,N_2080,N_722);
nand U3413 (N_3413,N_934,N_2425);
nand U3414 (N_3414,N_835,N_2311);
nor U3415 (N_3415,N_1895,N_1303);
nand U3416 (N_3416,N_1091,N_868);
and U3417 (N_3417,N_1823,N_2180);
xnor U3418 (N_3418,N_1500,N_1482);
xnor U3419 (N_3419,N_1058,N_287);
and U3420 (N_3420,N_1753,N_2458);
and U3421 (N_3421,N_880,N_1);
or U3422 (N_3422,N_791,N_188);
nor U3423 (N_3423,N_304,N_22);
xor U3424 (N_3424,N_130,N_1555);
or U3425 (N_3425,N_365,N_2372);
or U3426 (N_3426,N_1618,N_1973);
or U3427 (N_3427,N_1416,N_1396);
and U3428 (N_3428,N_1741,N_978);
nand U3429 (N_3429,N_1178,N_2434);
and U3430 (N_3430,N_2068,N_1328);
nor U3431 (N_3431,N_1146,N_1839);
xor U3432 (N_3432,N_348,N_1568);
nand U3433 (N_3433,N_2484,N_2296);
nor U3434 (N_3434,N_1124,N_684);
nand U3435 (N_3435,N_241,N_1690);
or U3436 (N_3436,N_1698,N_275);
or U3437 (N_3437,N_1100,N_299);
or U3438 (N_3438,N_803,N_1878);
or U3439 (N_3439,N_317,N_1319);
nor U3440 (N_3440,N_820,N_1951);
nor U3441 (N_3441,N_2394,N_922);
and U3442 (N_3442,N_1082,N_715);
nand U3443 (N_3443,N_659,N_1627);
and U3444 (N_3444,N_351,N_1991);
nand U3445 (N_3445,N_189,N_327);
xor U3446 (N_3446,N_460,N_1278);
and U3447 (N_3447,N_1574,N_1445);
xnor U3448 (N_3448,N_893,N_185);
nand U3449 (N_3449,N_212,N_2417);
and U3450 (N_3450,N_610,N_1522);
nor U3451 (N_3451,N_2002,N_491);
nor U3452 (N_3452,N_53,N_1967);
nand U3453 (N_3453,N_1333,N_528);
and U3454 (N_3454,N_1653,N_1472);
or U3455 (N_3455,N_2354,N_2388);
xor U3456 (N_3456,N_2166,N_2359);
or U3457 (N_3457,N_102,N_805);
nand U3458 (N_3458,N_2464,N_1849);
xor U3459 (N_3459,N_883,N_2336);
and U3460 (N_3460,N_679,N_2441);
or U3461 (N_3461,N_1442,N_1183);
xor U3462 (N_3462,N_338,N_214);
xor U3463 (N_3463,N_521,N_2183);
nand U3464 (N_3464,N_609,N_199);
and U3465 (N_3465,N_2435,N_792);
or U3466 (N_3466,N_271,N_1085);
and U3467 (N_3467,N_1115,N_1744);
xnor U3468 (N_3468,N_2190,N_554);
xor U3469 (N_3469,N_54,N_815);
xor U3470 (N_3470,N_196,N_2365);
and U3471 (N_3471,N_2187,N_31);
nand U3472 (N_3472,N_993,N_380);
or U3473 (N_3473,N_750,N_592);
and U3474 (N_3474,N_2442,N_286);
or U3475 (N_3475,N_1027,N_1460);
nor U3476 (N_3476,N_116,N_106);
nand U3477 (N_3477,N_1237,N_1824);
or U3478 (N_3478,N_1411,N_1760);
or U3479 (N_3479,N_226,N_938);
xnor U3480 (N_3480,N_2455,N_1350);
nor U3481 (N_3481,N_2379,N_424);
or U3482 (N_3482,N_220,N_1161);
or U3483 (N_3483,N_2322,N_585);
or U3484 (N_3484,N_1092,N_398);
or U3485 (N_3485,N_1828,N_1847);
nand U3486 (N_3486,N_887,N_981);
xor U3487 (N_3487,N_1391,N_726);
nand U3488 (N_3488,N_1904,N_2053);
and U3489 (N_3489,N_920,N_2123);
and U3490 (N_3490,N_2398,N_1586);
xnor U3491 (N_3491,N_929,N_2208);
nor U3492 (N_3492,N_785,N_202);
nor U3493 (N_3493,N_434,N_1217);
or U3494 (N_3494,N_1285,N_1940);
nand U3495 (N_3495,N_1361,N_2363);
nor U3496 (N_3496,N_2138,N_3);
nor U3497 (N_3497,N_2061,N_100);
xnor U3498 (N_3498,N_285,N_1066);
nand U3499 (N_3499,N_2004,N_2260);
nand U3500 (N_3500,N_966,N_2462);
and U3501 (N_3501,N_1758,N_2220);
nand U3502 (N_3502,N_2414,N_242);
nand U3503 (N_3503,N_34,N_1156);
nand U3504 (N_3504,N_1959,N_546);
or U3505 (N_3505,N_292,N_1399);
nand U3506 (N_3506,N_414,N_2171);
or U3507 (N_3507,N_2330,N_210);
and U3508 (N_3508,N_1282,N_251);
and U3509 (N_3509,N_73,N_83);
or U3510 (N_3510,N_1674,N_2017);
and U3511 (N_3511,N_1026,N_2449);
nand U3512 (N_3512,N_2351,N_2242);
nor U3513 (N_3513,N_274,N_2443);
xor U3514 (N_3514,N_2341,N_2444);
xnor U3515 (N_3515,N_745,N_1995);
nand U3516 (N_3516,N_1837,N_1848);
or U3517 (N_3517,N_1524,N_1693);
and U3518 (N_3518,N_384,N_957);
and U3519 (N_3519,N_63,N_589);
xnor U3520 (N_3520,N_1685,N_637);
and U3521 (N_3521,N_954,N_463);
or U3522 (N_3522,N_1454,N_1507);
nor U3523 (N_3523,N_2225,N_802);
and U3524 (N_3524,N_1327,N_1057);
nor U3525 (N_3525,N_773,N_1671);
or U3526 (N_3526,N_2150,N_1451);
or U3527 (N_3527,N_544,N_472);
nor U3528 (N_3528,N_714,N_987);
or U3529 (N_3529,N_1651,N_1050);
nand U3530 (N_3530,N_2153,N_1425);
xor U3531 (N_3531,N_305,N_138);
nand U3532 (N_3532,N_1202,N_2454);
and U3533 (N_3533,N_1682,N_1757);
xnor U3534 (N_3534,N_1304,N_1523);
nand U3535 (N_3535,N_1231,N_2157);
xor U3536 (N_3536,N_471,N_26);
or U3537 (N_3537,N_485,N_1150);
xnor U3538 (N_3538,N_1531,N_232);
xor U3539 (N_3539,N_500,N_1872);
or U3540 (N_3540,N_2104,N_1038);
and U3541 (N_3541,N_2050,N_4);
nand U3542 (N_3542,N_814,N_1883);
nor U3543 (N_3543,N_530,N_621);
nor U3544 (N_3544,N_2024,N_257);
and U3545 (N_3545,N_928,N_1003);
nor U3546 (N_3546,N_1281,N_428);
and U3547 (N_3547,N_206,N_1934);
and U3548 (N_3548,N_671,N_2075);
xnor U3549 (N_3549,N_1902,N_1825);
xnor U3550 (N_3550,N_2481,N_1787);
and U3551 (N_3551,N_2466,N_1688);
or U3552 (N_3552,N_357,N_395);
xnor U3553 (N_3553,N_296,N_2463);
or U3554 (N_3554,N_1072,N_499);
or U3555 (N_3555,N_470,N_240);
nand U3556 (N_3556,N_124,N_1219);
or U3557 (N_3557,N_1009,N_79);
and U3558 (N_3558,N_789,N_1811);
and U3559 (N_3559,N_1792,N_1945);
or U3560 (N_3560,N_1911,N_973);
and U3561 (N_3561,N_346,N_730);
and U3562 (N_3562,N_839,N_2056);
nand U3563 (N_3563,N_1234,N_1981);
and U3564 (N_3564,N_379,N_1903);
nor U3565 (N_3565,N_253,N_1002);
xor U3566 (N_3566,N_562,N_775);
nand U3567 (N_3567,N_1167,N_579);
nor U3568 (N_3568,N_612,N_1168);
or U3569 (N_3569,N_2347,N_1780);
and U3570 (N_3570,N_951,N_1438);
nand U3571 (N_3571,N_2284,N_2309);
nor U3572 (N_3572,N_369,N_1680);
or U3573 (N_3573,N_1866,N_1782);
or U3574 (N_3574,N_1403,N_1804);
or U3575 (N_3575,N_474,N_205);
or U3576 (N_3576,N_376,N_620);
nand U3577 (N_3577,N_1871,N_746);
nand U3578 (N_3578,N_494,N_1562);
or U3579 (N_3579,N_1305,N_1684);
and U3580 (N_3580,N_506,N_1083);
and U3581 (N_3581,N_1189,N_117);
or U3582 (N_3582,N_2117,N_1604);
nand U3583 (N_3583,N_2244,N_2340);
and U3584 (N_3584,N_408,N_832);
nor U3585 (N_3585,N_1761,N_2011);
nor U3586 (N_3586,N_489,N_2199);
or U3587 (N_3587,N_1480,N_836);
xor U3588 (N_3588,N_354,N_2412);
xnor U3589 (N_3589,N_334,N_1958);
nor U3590 (N_3590,N_1018,N_140);
nor U3591 (N_3591,N_496,N_2332);
xor U3592 (N_3592,N_302,N_1950);
nor U3593 (N_3593,N_873,N_1594);
or U3594 (N_3594,N_2023,N_1509);
nor U3595 (N_3595,N_2067,N_767);
xor U3596 (N_3596,N_1938,N_797);
or U3597 (N_3597,N_1288,N_1890);
nor U3598 (N_3598,N_1964,N_849);
xor U3599 (N_3599,N_2247,N_2312);
xnor U3600 (N_3600,N_2433,N_901);
or U3601 (N_3601,N_76,N_1094);
or U3602 (N_3602,N_2146,N_1519);
nor U3603 (N_3603,N_1858,N_120);
nand U3604 (N_3604,N_1267,N_281);
nor U3605 (N_3605,N_150,N_1446);
nor U3606 (N_3606,N_2007,N_593);
and U3607 (N_3607,N_1096,N_2352);
or U3608 (N_3608,N_971,N_2012);
nor U3609 (N_3609,N_1808,N_493);
and U3610 (N_3610,N_2283,N_1065);
or U3611 (N_3611,N_467,N_1404);
or U3612 (N_3612,N_1233,N_1235);
nor U3613 (N_3613,N_631,N_817);
and U3614 (N_3614,N_1258,N_1469);
and U3615 (N_3615,N_1349,N_1986);
nand U3616 (N_3616,N_1506,N_1019);
and U3617 (N_3617,N_1924,N_570);
nor U3618 (N_3618,N_2479,N_2013);
xnor U3619 (N_3619,N_1022,N_698);
nor U3620 (N_3620,N_823,N_2320);
nor U3621 (N_3621,N_1976,N_172);
or U3622 (N_3622,N_326,N_812);
nand U3623 (N_3623,N_2000,N_2255);
nor U3624 (N_3624,N_1062,N_2345);
and U3625 (N_3625,N_1492,N_1863);
and U3626 (N_3626,N_1689,N_1157);
or U3627 (N_3627,N_876,N_1722);
nor U3628 (N_3628,N_161,N_831);
or U3629 (N_3629,N_1307,N_2030);
or U3630 (N_3630,N_2230,N_223);
nor U3631 (N_3631,N_1323,N_2342);
xor U3632 (N_3632,N_1968,N_2);
or U3633 (N_3633,N_1781,N_2213);
nor U3634 (N_3634,N_1563,N_259);
and U3635 (N_3635,N_2346,N_2124);
or U3636 (N_3636,N_1128,N_1090);
nor U3637 (N_3637,N_1778,N_1495);
nor U3638 (N_3638,N_0,N_1490);
xor U3639 (N_3639,N_195,N_1994);
or U3640 (N_3640,N_807,N_125);
nand U3641 (N_3641,N_1434,N_1819);
or U3642 (N_3642,N_2313,N_1216);
nand U3643 (N_3643,N_1143,N_1838);
or U3644 (N_3644,N_991,N_1785);
or U3645 (N_3645,N_2485,N_1721);
or U3646 (N_3646,N_248,N_40);
or U3647 (N_3647,N_2262,N_543);
or U3648 (N_3648,N_1640,N_1429);
xor U3649 (N_3649,N_11,N_2206);
or U3650 (N_3650,N_1215,N_126);
nand U3651 (N_3651,N_1287,N_1014);
or U3652 (N_3652,N_513,N_458);
nand U3653 (N_3653,N_1337,N_1832);
xnor U3654 (N_3654,N_1283,N_689);
nand U3655 (N_3655,N_1270,N_1061);
or U3656 (N_3656,N_1692,N_377);
xor U3657 (N_3657,N_71,N_2217);
and U3658 (N_3658,N_2339,N_771);
and U3659 (N_3659,N_670,N_786);
and U3660 (N_3660,N_1367,N_2265);
and U3661 (N_3661,N_1084,N_1499);
and U3662 (N_3662,N_861,N_431);
and U3663 (N_3663,N_743,N_92);
and U3664 (N_3664,N_362,N_2295);
nand U3665 (N_3665,N_2249,N_1564);
and U3666 (N_3666,N_1218,N_308);
and U3667 (N_3667,N_1140,N_134);
nand U3668 (N_3668,N_850,N_455);
or U3669 (N_3669,N_219,N_1921);
nand U3670 (N_3670,N_1881,N_2461);
or U3671 (N_3671,N_1987,N_480);
nand U3672 (N_3672,N_1473,N_1794);
nand U3673 (N_3673,N_2175,N_1382);
xor U3674 (N_3674,N_2361,N_1619);
nand U3675 (N_3675,N_2266,N_2211);
nand U3676 (N_3676,N_246,N_284);
and U3677 (N_3677,N_200,N_764);
nand U3678 (N_3678,N_1601,N_2405);
nor U3679 (N_3679,N_2300,N_171);
nand U3680 (N_3680,N_575,N_244);
or U3681 (N_3681,N_1979,N_239);
or U3682 (N_3682,N_1683,N_685);
nand U3683 (N_3683,N_1833,N_1728);
and U3684 (N_3684,N_1907,N_1310);
xor U3685 (N_3685,N_123,N_1106);
nor U3686 (N_3686,N_2160,N_1139);
nor U3687 (N_3687,N_1279,N_306);
and U3688 (N_3688,N_1906,N_133);
nor U3689 (N_3689,N_2338,N_1408);
nand U3690 (N_3690,N_2473,N_1122);
nand U3691 (N_3691,N_1296,N_2130);
nor U3692 (N_3692,N_2251,N_1377);
nand U3693 (N_3693,N_1381,N_691);
xor U3694 (N_3694,N_1779,N_1997);
nor U3695 (N_3695,N_2456,N_2027);
nor U3696 (N_3696,N_57,N_1957);
nor U3697 (N_3697,N_364,N_625);
nand U3698 (N_3698,N_2204,N_710);
xor U3699 (N_3699,N_1329,N_443);
nand U3700 (N_3700,N_1730,N_787);
xnor U3701 (N_3701,N_1165,N_744);
nor U3702 (N_3702,N_755,N_425);
nor U3703 (N_3703,N_1592,N_1357);
nor U3704 (N_3704,N_2349,N_78);
nand U3705 (N_3705,N_2293,N_2205);
xnor U3706 (N_3706,N_2407,N_2279);
nand U3707 (N_3707,N_1443,N_2049);
and U3708 (N_3708,N_10,N_905);
or U3709 (N_3709,N_1386,N_1424);
nand U3710 (N_3710,N_1170,N_1820);
and U3711 (N_3711,N_355,N_2437);
nand U3712 (N_3712,N_96,N_606);
or U3713 (N_3713,N_1850,N_363);
nand U3714 (N_3714,N_1154,N_2118);
or U3715 (N_3715,N_1855,N_926);
or U3716 (N_3716,N_2134,N_2058);
nor U3717 (N_3717,N_28,N_2371);
or U3718 (N_3718,N_17,N_1300);
or U3719 (N_3719,N_1766,N_2113);
or U3720 (N_3720,N_479,N_462);
nand U3721 (N_3721,N_597,N_763);
xor U3722 (N_3722,N_288,N_2038);
or U3723 (N_3723,N_1475,N_2028);
nand U3724 (N_3724,N_1129,N_702);
nand U3725 (N_3725,N_293,N_1095);
nand U3726 (N_3726,N_1383,N_508);
or U3727 (N_3727,N_2059,N_997);
nor U3728 (N_3728,N_1503,N_683);
or U3729 (N_3729,N_1970,N_1130);
and U3730 (N_3730,N_490,N_449);
xor U3731 (N_3731,N_149,N_753);
xor U3732 (N_3732,N_168,N_897);
nand U3733 (N_3733,N_1190,N_1665);
xnor U3734 (N_3734,N_1742,N_1852);
nor U3735 (N_3735,N_1254,N_1201);
nor U3736 (N_3736,N_2119,N_2297);
and U3737 (N_3737,N_1419,N_2475);
and U3738 (N_3738,N_1817,N_475);
nand U3739 (N_3739,N_227,N_564);
xor U3740 (N_3740,N_2236,N_2133);
nor U3741 (N_3741,N_2154,N_1897);
or U3742 (N_3742,N_1370,N_2377);
nand U3743 (N_3743,N_1272,N_322);
and U3744 (N_3744,N_1648,N_1198);
xnor U3745 (N_3745,N_153,N_1232);
xor U3746 (N_3746,N_2082,N_591);
or U3747 (N_3747,N_1786,N_2348);
nand U3748 (N_3748,N_1292,N_387);
and U3749 (N_3749,N_672,N_1937);
xnor U3750 (N_3750,N_2390,N_2177);
or U3751 (N_3751,N_434,N_1781);
or U3752 (N_3752,N_124,N_1039);
xor U3753 (N_3753,N_777,N_841);
or U3754 (N_3754,N_599,N_2160);
and U3755 (N_3755,N_2400,N_531);
nor U3756 (N_3756,N_1986,N_1598);
and U3757 (N_3757,N_483,N_663);
and U3758 (N_3758,N_1008,N_1819);
xnor U3759 (N_3759,N_1183,N_1726);
nand U3760 (N_3760,N_1973,N_2123);
and U3761 (N_3761,N_2334,N_1785);
or U3762 (N_3762,N_2327,N_1047);
xnor U3763 (N_3763,N_1552,N_1844);
nor U3764 (N_3764,N_1788,N_1902);
nand U3765 (N_3765,N_1031,N_2371);
nor U3766 (N_3766,N_365,N_789);
nand U3767 (N_3767,N_1151,N_210);
xor U3768 (N_3768,N_402,N_2446);
nor U3769 (N_3769,N_670,N_1609);
or U3770 (N_3770,N_2276,N_580);
nand U3771 (N_3771,N_1092,N_508);
nor U3772 (N_3772,N_2264,N_1265);
nor U3773 (N_3773,N_1212,N_1354);
nor U3774 (N_3774,N_2088,N_694);
xor U3775 (N_3775,N_480,N_1026);
or U3776 (N_3776,N_975,N_1543);
or U3777 (N_3777,N_223,N_969);
nor U3778 (N_3778,N_781,N_108);
nand U3779 (N_3779,N_1926,N_1057);
nor U3780 (N_3780,N_1472,N_718);
and U3781 (N_3781,N_777,N_2241);
nor U3782 (N_3782,N_2231,N_608);
and U3783 (N_3783,N_1594,N_1336);
nor U3784 (N_3784,N_648,N_1771);
or U3785 (N_3785,N_751,N_2386);
and U3786 (N_3786,N_560,N_257);
xnor U3787 (N_3787,N_424,N_2151);
nand U3788 (N_3788,N_607,N_1075);
and U3789 (N_3789,N_1066,N_1);
nand U3790 (N_3790,N_1358,N_2288);
nor U3791 (N_3791,N_278,N_1009);
xnor U3792 (N_3792,N_2274,N_1053);
and U3793 (N_3793,N_966,N_2405);
or U3794 (N_3794,N_2108,N_470);
nand U3795 (N_3795,N_683,N_2422);
or U3796 (N_3796,N_1794,N_288);
nor U3797 (N_3797,N_319,N_1981);
and U3798 (N_3798,N_2384,N_1615);
nor U3799 (N_3799,N_1308,N_382);
nor U3800 (N_3800,N_1998,N_446);
nor U3801 (N_3801,N_384,N_939);
nand U3802 (N_3802,N_1133,N_1720);
and U3803 (N_3803,N_1033,N_659);
xnor U3804 (N_3804,N_1111,N_1135);
and U3805 (N_3805,N_1806,N_1182);
nand U3806 (N_3806,N_1567,N_423);
and U3807 (N_3807,N_753,N_2086);
and U3808 (N_3808,N_1341,N_1659);
and U3809 (N_3809,N_1438,N_370);
nand U3810 (N_3810,N_1098,N_1384);
or U3811 (N_3811,N_2351,N_801);
nand U3812 (N_3812,N_589,N_397);
xnor U3813 (N_3813,N_1972,N_911);
or U3814 (N_3814,N_1727,N_642);
or U3815 (N_3815,N_2495,N_201);
or U3816 (N_3816,N_1595,N_498);
and U3817 (N_3817,N_267,N_126);
and U3818 (N_3818,N_325,N_885);
nor U3819 (N_3819,N_645,N_2138);
nor U3820 (N_3820,N_1651,N_1212);
and U3821 (N_3821,N_1264,N_622);
and U3822 (N_3822,N_1575,N_621);
xor U3823 (N_3823,N_653,N_386);
xor U3824 (N_3824,N_1538,N_200);
nor U3825 (N_3825,N_269,N_1089);
xnor U3826 (N_3826,N_339,N_1016);
xor U3827 (N_3827,N_154,N_556);
nor U3828 (N_3828,N_7,N_487);
or U3829 (N_3829,N_2077,N_921);
and U3830 (N_3830,N_2023,N_984);
nor U3831 (N_3831,N_681,N_1849);
or U3832 (N_3832,N_2277,N_138);
nand U3833 (N_3833,N_1969,N_2497);
or U3834 (N_3834,N_635,N_1880);
or U3835 (N_3835,N_580,N_362);
and U3836 (N_3836,N_442,N_1594);
nor U3837 (N_3837,N_2120,N_676);
nor U3838 (N_3838,N_630,N_604);
xnor U3839 (N_3839,N_1125,N_989);
nand U3840 (N_3840,N_1531,N_1396);
nand U3841 (N_3841,N_2456,N_131);
xnor U3842 (N_3842,N_1659,N_2193);
and U3843 (N_3843,N_1740,N_1907);
or U3844 (N_3844,N_1218,N_625);
nand U3845 (N_3845,N_695,N_1456);
nor U3846 (N_3846,N_2260,N_2007);
nand U3847 (N_3847,N_796,N_1360);
nor U3848 (N_3848,N_1726,N_134);
nand U3849 (N_3849,N_1072,N_2365);
and U3850 (N_3850,N_492,N_756);
xnor U3851 (N_3851,N_790,N_825);
nand U3852 (N_3852,N_1078,N_1412);
nand U3853 (N_3853,N_2395,N_1751);
nand U3854 (N_3854,N_914,N_2044);
and U3855 (N_3855,N_1486,N_1777);
and U3856 (N_3856,N_2379,N_905);
nor U3857 (N_3857,N_575,N_1580);
and U3858 (N_3858,N_2333,N_527);
nand U3859 (N_3859,N_1282,N_525);
and U3860 (N_3860,N_2174,N_93);
nor U3861 (N_3861,N_2161,N_2071);
nand U3862 (N_3862,N_1777,N_996);
and U3863 (N_3863,N_2472,N_1187);
or U3864 (N_3864,N_588,N_153);
or U3865 (N_3865,N_163,N_343);
and U3866 (N_3866,N_2102,N_756);
xnor U3867 (N_3867,N_1925,N_937);
and U3868 (N_3868,N_758,N_289);
and U3869 (N_3869,N_1686,N_1687);
nor U3870 (N_3870,N_1455,N_600);
nand U3871 (N_3871,N_1246,N_32);
or U3872 (N_3872,N_964,N_87);
and U3873 (N_3873,N_702,N_206);
nand U3874 (N_3874,N_2019,N_800);
nand U3875 (N_3875,N_1800,N_741);
nand U3876 (N_3876,N_1885,N_85);
nor U3877 (N_3877,N_1764,N_1767);
nand U3878 (N_3878,N_39,N_16);
nor U3879 (N_3879,N_389,N_1755);
nor U3880 (N_3880,N_746,N_1022);
and U3881 (N_3881,N_1389,N_1837);
or U3882 (N_3882,N_1354,N_1775);
nor U3883 (N_3883,N_1624,N_927);
or U3884 (N_3884,N_1599,N_1866);
nand U3885 (N_3885,N_708,N_619);
or U3886 (N_3886,N_277,N_1231);
nor U3887 (N_3887,N_267,N_1924);
or U3888 (N_3888,N_2157,N_1134);
and U3889 (N_3889,N_2475,N_1320);
or U3890 (N_3890,N_898,N_2433);
xor U3891 (N_3891,N_708,N_566);
xor U3892 (N_3892,N_348,N_2306);
or U3893 (N_3893,N_1189,N_912);
xor U3894 (N_3894,N_259,N_1463);
and U3895 (N_3895,N_58,N_833);
and U3896 (N_3896,N_775,N_1169);
nand U3897 (N_3897,N_2448,N_2315);
and U3898 (N_3898,N_836,N_981);
and U3899 (N_3899,N_2472,N_2461);
nand U3900 (N_3900,N_1853,N_1779);
nand U3901 (N_3901,N_2078,N_170);
and U3902 (N_3902,N_588,N_2251);
or U3903 (N_3903,N_546,N_1691);
or U3904 (N_3904,N_2364,N_1937);
and U3905 (N_3905,N_2356,N_1241);
and U3906 (N_3906,N_922,N_2070);
nand U3907 (N_3907,N_763,N_72);
xnor U3908 (N_3908,N_1500,N_934);
xor U3909 (N_3909,N_2067,N_133);
and U3910 (N_3910,N_103,N_1189);
and U3911 (N_3911,N_596,N_1028);
and U3912 (N_3912,N_1066,N_1052);
or U3913 (N_3913,N_2000,N_1417);
xor U3914 (N_3914,N_2084,N_1696);
nor U3915 (N_3915,N_988,N_520);
xor U3916 (N_3916,N_62,N_1721);
nand U3917 (N_3917,N_2344,N_1612);
and U3918 (N_3918,N_591,N_2240);
and U3919 (N_3919,N_1220,N_1769);
xor U3920 (N_3920,N_431,N_907);
nor U3921 (N_3921,N_1907,N_2162);
or U3922 (N_3922,N_2275,N_1481);
or U3923 (N_3923,N_989,N_219);
xnor U3924 (N_3924,N_190,N_1634);
nand U3925 (N_3925,N_1773,N_2167);
or U3926 (N_3926,N_1592,N_1964);
xor U3927 (N_3927,N_248,N_363);
xnor U3928 (N_3928,N_95,N_146);
and U3929 (N_3929,N_123,N_2365);
xnor U3930 (N_3930,N_1751,N_1746);
nand U3931 (N_3931,N_1875,N_769);
and U3932 (N_3932,N_2257,N_418);
xnor U3933 (N_3933,N_2346,N_2359);
nor U3934 (N_3934,N_1094,N_1575);
xnor U3935 (N_3935,N_1396,N_708);
nor U3936 (N_3936,N_785,N_1952);
nor U3937 (N_3937,N_1935,N_2184);
xor U3938 (N_3938,N_1918,N_2196);
nor U3939 (N_3939,N_2244,N_274);
or U3940 (N_3940,N_990,N_1499);
and U3941 (N_3941,N_324,N_1595);
nor U3942 (N_3942,N_734,N_469);
nor U3943 (N_3943,N_147,N_288);
nor U3944 (N_3944,N_652,N_1006);
and U3945 (N_3945,N_54,N_57);
or U3946 (N_3946,N_1037,N_1971);
nor U3947 (N_3947,N_2173,N_2021);
nor U3948 (N_3948,N_1014,N_1634);
and U3949 (N_3949,N_1431,N_263);
or U3950 (N_3950,N_464,N_2435);
or U3951 (N_3951,N_1507,N_243);
or U3952 (N_3952,N_565,N_1805);
and U3953 (N_3953,N_1510,N_663);
or U3954 (N_3954,N_2230,N_1923);
or U3955 (N_3955,N_337,N_2138);
xnor U3956 (N_3956,N_966,N_591);
or U3957 (N_3957,N_714,N_1574);
and U3958 (N_3958,N_548,N_2165);
xor U3959 (N_3959,N_1812,N_2234);
or U3960 (N_3960,N_222,N_6);
or U3961 (N_3961,N_1929,N_2434);
nor U3962 (N_3962,N_587,N_1658);
nor U3963 (N_3963,N_2331,N_1584);
nor U3964 (N_3964,N_533,N_789);
nand U3965 (N_3965,N_625,N_235);
nor U3966 (N_3966,N_812,N_1349);
or U3967 (N_3967,N_794,N_543);
and U3968 (N_3968,N_1022,N_2411);
xnor U3969 (N_3969,N_1518,N_636);
nor U3970 (N_3970,N_136,N_1226);
and U3971 (N_3971,N_2397,N_111);
nor U3972 (N_3972,N_11,N_2236);
or U3973 (N_3973,N_2207,N_1635);
and U3974 (N_3974,N_703,N_1039);
xor U3975 (N_3975,N_546,N_435);
or U3976 (N_3976,N_1495,N_1948);
nor U3977 (N_3977,N_1381,N_1086);
xor U3978 (N_3978,N_737,N_1963);
or U3979 (N_3979,N_2007,N_910);
xor U3980 (N_3980,N_1309,N_945);
nor U3981 (N_3981,N_1899,N_538);
xnor U3982 (N_3982,N_1880,N_176);
nand U3983 (N_3983,N_563,N_972);
nand U3984 (N_3984,N_158,N_1274);
or U3985 (N_3985,N_613,N_1780);
and U3986 (N_3986,N_2200,N_437);
or U3987 (N_3987,N_1073,N_1985);
or U3988 (N_3988,N_963,N_2397);
xnor U3989 (N_3989,N_1603,N_990);
nor U3990 (N_3990,N_1455,N_859);
and U3991 (N_3991,N_509,N_936);
nand U3992 (N_3992,N_1581,N_667);
or U3993 (N_3993,N_1785,N_2035);
nor U3994 (N_3994,N_1838,N_2262);
xor U3995 (N_3995,N_109,N_45);
and U3996 (N_3996,N_1566,N_615);
nor U3997 (N_3997,N_653,N_373);
xnor U3998 (N_3998,N_249,N_2437);
xnor U3999 (N_3999,N_642,N_198);
and U4000 (N_4000,N_1664,N_2495);
or U4001 (N_4001,N_1644,N_323);
nor U4002 (N_4002,N_1334,N_39);
nand U4003 (N_4003,N_2397,N_2108);
nor U4004 (N_4004,N_1061,N_1845);
or U4005 (N_4005,N_99,N_2250);
and U4006 (N_4006,N_1065,N_64);
nor U4007 (N_4007,N_2024,N_837);
and U4008 (N_4008,N_1627,N_444);
nand U4009 (N_4009,N_487,N_1411);
nand U4010 (N_4010,N_481,N_2212);
nand U4011 (N_4011,N_1029,N_2136);
or U4012 (N_4012,N_455,N_1402);
nand U4013 (N_4013,N_801,N_550);
nor U4014 (N_4014,N_257,N_1284);
nand U4015 (N_4015,N_774,N_1204);
or U4016 (N_4016,N_1679,N_1273);
and U4017 (N_4017,N_2387,N_1521);
and U4018 (N_4018,N_482,N_1703);
and U4019 (N_4019,N_1275,N_1);
or U4020 (N_4020,N_546,N_973);
nand U4021 (N_4021,N_1461,N_534);
nor U4022 (N_4022,N_1682,N_1685);
or U4023 (N_4023,N_1702,N_1842);
nor U4024 (N_4024,N_548,N_1700);
xor U4025 (N_4025,N_1757,N_1921);
nor U4026 (N_4026,N_777,N_1357);
xor U4027 (N_4027,N_58,N_998);
or U4028 (N_4028,N_1582,N_668);
or U4029 (N_4029,N_358,N_1615);
and U4030 (N_4030,N_2280,N_1324);
and U4031 (N_4031,N_1470,N_1909);
or U4032 (N_4032,N_933,N_818);
and U4033 (N_4033,N_998,N_1399);
or U4034 (N_4034,N_1398,N_2468);
or U4035 (N_4035,N_80,N_209);
nor U4036 (N_4036,N_2134,N_922);
nor U4037 (N_4037,N_856,N_1839);
or U4038 (N_4038,N_515,N_1212);
or U4039 (N_4039,N_391,N_2123);
and U4040 (N_4040,N_1567,N_2217);
nand U4041 (N_4041,N_953,N_2238);
nand U4042 (N_4042,N_1171,N_672);
nor U4043 (N_4043,N_2032,N_863);
xor U4044 (N_4044,N_2298,N_75);
nand U4045 (N_4045,N_1423,N_1556);
xor U4046 (N_4046,N_1521,N_1288);
nand U4047 (N_4047,N_324,N_1051);
or U4048 (N_4048,N_448,N_1314);
or U4049 (N_4049,N_906,N_2231);
nor U4050 (N_4050,N_998,N_538);
nor U4051 (N_4051,N_653,N_1282);
nor U4052 (N_4052,N_1612,N_620);
or U4053 (N_4053,N_320,N_2081);
and U4054 (N_4054,N_2396,N_2402);
nor U4055 (N_4055,N_1308,N_262);
and U4056 (N_4056,N_1456,N_812);
or U4057 (N_4057,N_669,N_233);
and U4058 (N_4058,N_1456,N_1792);
xor U4059 (N_4059,N_489,N_2268);
nor U4060 (N_4060,N_2404,N_2148);
or U4061 (N_4061,N_814,N_2375);
and U4062 (N_4062,N_1891,N_2397);
nand U4063 (N_4063,N_2091,N_1665);
and U4064 (N_4064,N_566,N_815);
xor U4065 (N_4065,N_936,N_1215);
xnor U4066 (N_4066,N_2399,N_2015);
xor U4067 (N_4067,N_1364,N_642);
xor U4068 (N_4068,N_328,N_1824);
and U4069 (N_4069,N_180,N_1142);
or U4070 (N_4070,N_152,N_258);
xnor U4071 (N_4071,N_1287,N_1967);
nand U4072 (N_4072,N_1003,N_1941);
xnor U4073 (N_4073,N_1730,N_2106);
xor U4074 (N_4074,N_2268,N_2340);
and U4075 (N_4075,N_992,N_1711);
nor U4076 (N_4076,N_1531,N_1965);
nor U4077 (N_4077,N_1076,N_576);
or U4078 (N_4078,N_414,N_509);
xor U4079 (N_4079,N_596,N_1053);
or U4080 (N_4080,N_839,N_328);
and U4081 (N_4081,N_134,N_63);
nand U4082 (N_4082,N_2194,N_1855);
and U4083 (N_4083,N_724,N_230);
and U4084 (N_4084,N_2449,N_189);
and U4085 (N_4085,N_1974,N_2046);
and U4086 (N_4086,N_473,N_8);
and U4087 (N_4087,N_223,N_1161);
or U4088 (N_4088,N_2216,N_2267);
nand U4089 (N_4089,N_184,N_451);
nand U4090 (N_4090,N_592,N_1725);
xnor U4091 (N_4091,N_1158,N_635);
xor U4092 (N_4092,N_1503,N_341);
nand U4093 (N_4093,N_1059,N_200);
nor U4094 (N_4094,N_801,N_2211);
xor U4095 (N_4095,N_2211,N_1002);
nand U4096 (N_4096,N_845,N_2445);
nor U4097 (N_4097,N_412,N_795);
and U4098 (N_4098,N_2481,N_2303);
xnor U4099 (N_4099,N_533,N_1588);
and U4100 (N_4100,N_1363,N_1545);
nor U4101 (N_4101,N_2327,N_2435);
nor U4102 (N_4102,N_69,N_1860);
nor U4103 (N_4103,N_285,N_1737);
or U4104 (N_4104,N_1632,N_1575);
and U4105 (N_4105,N_2379,N_2011);
and U4106 (N_4106,N_668,N_1807);
and U4107 (N_4107,N_2278,N_1803);
xor U4108 (N_4108,N_197,N_294);
and U4109 (N_4109,N_896,N_356);
xor U4110 (N_4110,N_999,N_467);
nand U4111 (N_4111,N_740,N_1782);
or U4112 (N_4112,N_1910,N_2035);
and U4113 (N_4113,N_2156,N_2249);
xor U4114 (N_4114,N_2499,N_1888);
xnor U4115 (N_4115,N_2434,N_2457);
or U4116 (N_4116,N_2475,N_404);
xor U4117 (N_4117,N_1416,N_1261);
nor U4118 (N_4118,N_2486,N_1201);
nor U4119 (N_4119,N_821,N_232);
nor U4120 (N_4120,N_2309,N_2119);
nand U4121 (N_4121,N_546,N_1039);
and U4122 (N_4122,N_952,N_1942);
nand U4123 (N_4123,N_177,N_797);
xor U4124 (N_4124,N_2145,N_897);
or U4125 (N_4125,N_112,N_461);
and U4126 (N_4126,N_1679,N_589);
xor U4127 (N_4127,N_1624,N_942);
xnor U4128 (N_4128,N_204,N_2117);
xnor U4129 (N_4129,N_265,N_1759);
nor U4130 (N_4130,N_1294,N_1239);
xor U4131 (N_4131,N_218,N_1101);
nand U4132 (N_4132,N_819,N_2028);
xor U4133 (N_4133,N_570,N_2455);
or U4134 (N_4134,N_1714,N_61);
and U4135 (N_4135,N_376,N_742);
xnor U4136 (N_4136,N_42,N_1732);
nand U4137 (N_4137,N_1193,N_2457);
xnor U4138 (N_4138,N_1056,N_2283);
or U4139 (N_4139,N_1557,N_484);
and U4140 (N_4140,N_399,N_529);
xnor U4141 (N_4141,N_1369,N_1154);
and U4142 (N_4142,N_208,N_2044);
and U4143 (N_4143,N_1787,N_770);
or U4144 (N_4144,N_1813,N_1880);
and U4145 (N_4145,N_1233,N_1070);
xor U4146 (N_4146,N_1180,N_267);
nand U4147 (N_4147,N_671,N_1735);
nand U4148 (N_4148,N_1417,N_1768);
and U4149 (N_4149,N_2063,N_1796);
and U4150 (N_4150,N_704,N_78);
nor U4151 (N_4151,N_1983,N_1270);
xnor U4152 (N_4152,N_521,N_1031);
and U4153 (N_4153,N_85,N_1254);
and U4154 (N_4154,N_2419,N_2052);
nand U4155 (N_4155,N_2134,N_196);
or U4156 (N_4156,N_1961,N_515);
nor U4157 (N_4157,N_1177,N_1837);
or U4158 (N_4158,N_2232,N_981);
nand U4159 (N_4159,N_2304,N_2195);
and U4160 (N_4160,N_325,N_1937);
xnor U4161 (N_4161,N_797,N_198);
nand U4162 (N_4162,N_2350,N_884);
nand U4163 (N_4163,N_44,N_833);
and U4164 (N_4164,N_2322,N_408);
and U4165 (N_4165,N_899,N_217);
or U4166 (N_4166,N_1076,N_2489);
and U4167 (N_4167,N_2142,N_1054);
xnor U4168 (N_4168,N_964,N_1842);
and U4169 (N_4169,N_1421,N_1650);
xor U4170 (N_4170,N_1226,N_313);
or U4171 (N_4171,N_499,N_2251);
or U4172 (N_4172,N_949,N_1062);
nand U4173 (N_4173,N_1265,N_1240);
nor U4174 (N_4174,N_745,N_274);
nor U4175 (N_4175,N_1039,N_1707);
xor U4176 (N_4176,N_313,N_677);
nand U4177 (N_4177,N_485,N_2150);
and U4178 (N_4178,N_2074,N_1703);
xnor U4179 (N_4179,N_1479,N_1341);
nor U4180 (N_4180,N_1209,N_1234);
nand U4181 (N_4181,N_888,N_1929);
or U4182 (N_4182,N_1274,N_306);
nand U4183 (N_4183,N_1341,N_1509);
nand U4184 (N_4184,N_979,N_1847);
nand U4185 (N_4185,N_2047,N_1366);
xor U4186 (N_4186,N_2162,N_320);
and U4187 (N_4187,N_1551,N_934);
nand U4188 (N_4188,N_1797,N_249);
or U4189 (N_4189,N_2416,N_667);
nor U4190 (N_4190,N_1825,N_1058);
xnor U4191 (N_4191,N_1555,N_1208);
xor U4192 (N_4192,N_390,N_1827);
nor U4193 (N_4193,N_41,N_1885);
nand U4194 (N_4194,N_2293,N_1058);
xor U4195 (N_4195,N_25,N_990);
nand U4196 (N_4196,N_427,N_1221);
nor U4197 (N_4197,N_93,N_1061);
nand U4198 (N_4198,N_1158,N_67);
or U4199 (N_4199,N_2198,N_1380);
xnor U4200 (N_4200,N_1824,N_1120);
nor U4201 (N_4201,N_1931,N_145);
xor U4202 (N_4202,N_2155,N_393);
or U4203 (N_4203,N_288,N_1003);
xnor U4204 (N_4204,N_2219,N_1578);
nand U4205 (N_4205,N_688,N_1699);
nand U4206 (N_4206,N_1674,N_1383);
xnor U4207 (N_4207,N_2152,N_1510);
and U4208 (N_4208,N_1392,N_978);
nand U4209 (N_4209,N_2137,N_2138);
nand U4210 (N_4210,N_1334,N_424);
nand U4211 (N_4211,N_2035,N_2053);
nand U4212 (N_4212,N_1000,N_1115);
and U4213 (N_4213,N_235,N_1856);
and U4214 (N_4214,N_2284,N_869);
xor U4215 (N_4215,N_263,N_2290);
nand U4216 (N_4216,N_2264,N_268);
nor U4217 (N_4217,N_697,N_834);
or U4218 (N_4218,N_97,N_676);
xnor U4219 (N_4219,N_2008,N_2188);
nand U4220 (N_4220,N_146,N_985);
nand U4221 (N_4221,N_2023,N_419);
xor U4222 (N_4222,N_1244,N_368);
or U4223 (N_4223,N_2333,N_87);
or U4224 (N_4224,N_447,N_180);
nand U4225 (N_4225,N_1691,N_688);
nor U4226 (N_4226,N_1624,N_2358);
and U4227 (N_4227,N_39,N_730);
xnor U4228 (N_4228,N_539,N_2220);
xor U4229 (N_4229,N_1850,N_250);
nand U4230 (N_4230,N_2453,N_1967);
and U4231 (N_4231,N_2006,N_1053);
nand U4232 (N_4232,N_419,N_1959);
and U4233 (N_4233,N_2396,N_1967);
and U4234 (N_4234,N_1928,N_1567);
nor U4235 (N_4235,N_1784,N_1668);
xnor U4236 (N_4236,N_481,N_2409);
and U4237 (N_4237,N_1747,N_1246);
xor U4238 (N_4238,N_1835,N_2068);
nand U4239 (N_4239,N_1055,N_1063);
xnor U4240 (N_4240,N_501,N_850);
and U4241 (N_4241,N_1903,N_2231);
and U4242 (N_4242,N_2495,N_1859);
and U4243 (N_4243,N_1381,N_2492);
nand U4244 (N_4244,N_1579,N_1443);
and U4245 (N_4245,N_1873,N_988);
or U4246 (N_4246,N_2116,N_1476);
nor U4247 (N_4247,N_1675,N_703);
and U4248 (N_4248,N_91,N_1624);
xor U4249 (N_4249,N_1925,N_1862);
nor U4250 (N_4250,N_2010,N_2308);
xnor U4251 (N_4251,N_493,N_1520);
nand U4252 (N_4252,N_264,N_670);
or U4253 (N_4253,N_1456,N_382);
nor U4254 (N_4254,N_1220,N_1898);
xnor U4255 (N_4255,N_29,N_812);
nand U4256 (N_4256,N_336,N_1545);
nand U4257 (N_4257,N_467,N_138);
and U4258 (N_4258,N_411,N_103);
or U4259 (N_4259,N_1293,N_160);
nand U4260 (N_4260,N_836,N_815);
or U4261 (N_4261,N_1307,N_540);
or U4262 (N_4262,N_2114,N_1640);
nand U4263 (N_4263,N_1164,N_1223);
and U4264 (N_4264,N_561,N_828);
xnor U4265 (N_4265,N_897,N_1834);
or U4266 (N_4266,N_871,N_824);
nor U4267 (N_4267,N_202,N_1074);
nor U4268 (N_4268,N_141,N_693);
xor U4269 (N_4269,N_1231,N_1946);
nand U4270 (N_4270,N_1782,N_1147);
and U4271 (N_4271,N_2407,N_435);
or U4272 (N_4272,N_810,N_920);
nor U4273 (N_4273,N_1276,N_847);
and U4274 (N_4274,N_2457,N_1913);
xor U4275 (N_4275,N_578,N_1959);
xnor U4276 (N_4276,N_802,N_1465);
xnor U4277 (N_4277,N_1488,N_2005);
and U4278 (N_4278,N_459,N_2167);
or U4279 (N_4279,N_1946,N_1222);
and U4280 (N_4280,N_126,N_748);
nand U4281 (N_4281,N_1157,N_286);
xnor U4282 (N_4282,N_266,N_593);
nand U4283 (N_4283,N_2489,N_1998);
nor U4284 (N_4284,N_1207,N_390);
nor U4285 (N_4285,N_1629,N_1828);
xnor U4286 (N_4286,N_644,N_149);
and U4287 (N_4287,N_2211,N_22);
nand U4288 (N_4288,N_456,N_1556);
or U4289 (N_4289,N_2143,N_275);
or U4290 (N_4290,N_2303,N_1317);
and U4291 (N_4291,N_1276,N_410);
nor U4292 (N_4292,N_898,N_415);
nand U4293 (N_4293,N_1526,N_1678);
xor U4294 (N_4294,N_129,N_1878);
and U4295 (N_4295,N_1094,N_2193);
and U4296 (N_4296,N_1503,N_1212);
nor U4297 (N_4297,N_1625,N_380);
nand U4298 (N_4298,N_2058,N_870);
and U4299 (N_4299,N_2498,N_560);
or U4300 (N_4300,N_312,N_1640);
xor U4301 (N_4301,N_778,N_2095);
nand U4302 (N_4302,N_1191,N_310);
xnor U4303 (N_4303,N_299,N_1107);
and U4304 (N_4304,N_975,N_904);
xnor U4305 (N_4305,N_2089,N_877);
xnor U4306 (N_4306,N_1101,N_2127);
or U4307 (N_4307,N_1263,N_385);
and U4308 (N_4308,N_229,N_514);
or U4309 (N_4309,N_1443,N_651);
or U4310 (N_4310,N_1890,N_2014);
xor U4311 (N_4311,N_1602,N_1433);
xnor U4312 (N_4312,N_595,N_2042);
xor U4313 (N_4313,N_694,N_1021);
nand U4314 (N_4314,N_2360,N_1280);
or U4315 (N_4315,N_1411,N_1578);
or U4316 (N_4316,N_1302,N_678);
and U4317 (N_4317,N_1741,N_1089);
xor U4318 (N_4318,N_398,N_2384);
nor U4319 (N_4319,N_1216,N_1267);
nand U4320 (N_4320,N_2143,N_138);
nand U4321 (N_4321,N_1615,N_2360);
nand U4322 (N_4322,N_1994,N_1125);
nor U4323 (N_4323,N_1732,N_1743);
xnor U4324 (N_4324,N_416,N_2286);
xnor U4325 (N_4325,N_2041,N_1033);
and U4326 (N_4326,N_234,N_1259);
nor U4327 (N_4327,N_1168,N_2334);
and U4328 (N_4328,N_1481,N_518);
and U4329 (N_4329,N_2159,N_1388);
and U4330 (N_4330,N_1775,N_1644);
xnor U4331 (N_4331,N_563,N_1630);
or U4332 (N_4332,N_1924,N_1222);
nor U4333 (N_4333,N_1336,N_1948);
and U4334 (N_4334,N_461,N_2366);
nand U4335 (N_4335,N_1544,N_508);
nor U4336 (N_4336,N_4,N_1150);
xnor U4337 (N_4337,N_2346,N_613);
xnor U4338 (N_4338,N_695,N_1467);
or U4339 (N_4339,N_129,N_214);
xor U4340 (N_4340,N_1198,N_489);
nand U4341 (N_4341,N_2153,N_2254);
xnor U4342 (N_4342,N_339,N_1757);
xor U4343 (N_4343,N_39,N_1602);
or U4344 (N_4344,N_1131,N_1005);
nor U4345 (N_4345,N_1026,N_1863);
xnor U4346 (N_4346,N_1691,N_1483);
and U4347 (N_4347,N_1758,N_497);
or U4348 (N_4348,N_1491,N_2051);
or U4349 (N_4349,N_1047,N_699);
nor U4350 (N_4350,N_1562,N_181);
nor U4351 (N_4351,N_1677,N_408);
nor U4352 (N_4352,N_326,N_277);
nand U4353 (N_4353,N_584,N_2169);
nor U4354 (N_4354,N_144,N_689);
nor U4355 (N_4355,N_1301,N_432);
or U4356 (N_4356,N_383,N_1199);
xnor U4357 (N_4357,N_807,N_2154);
and U4358 (N_4358,N_1512,N_1719);
and U4359 (N_4359,N_1916,N_1980);
xnor U4360 (N_4360,N_836,N_963);
and U4361 (N_4361,N_805,N_983);
nand U4362 (N_4362,N_149,N_2033);
nand U4363 (N_4363,N_2041,N_1997);
nor U4364 (N_4364,N_763,N_1053);
nor U4365 (N_4365,N_1891,N_824);
and U4366 (N_4366,N_282,N_398);
nor U4367 (N_4367,N_986,N_1685);
or U4368 (N_4368,N_729,N_609);
nand U4369 (N_4369,N_237,N_404);
or U4370 (N_4370,N_1454,N_1978);
nand U4371 (N_4371,N_2492,N_492);
nor U4372 (N_4372,N_2018,N_1509);
or U4373 (N_4373,N_710,N_181);
nor U4374 (N_4374,N_433,N_1948);
and U4375 (N_4375,N_140,N_1773);
nand U4376 (N_4376,N_1135,N_747);
or U4377 (N_4377,N_1386,N_76);
and U4378 (N_4378,N_314,N_902);
nor U4379 (N_4379,N_28,N_1733);
and U4380 (N_4380,N_1712,N_2426);
nand U4381 (N_4381,N_1440,N_712);
nor U4382 (N_4382,N_1638,N_693);
xor U4383 (N_4383,N_2372,N_118);
or U4384 (N_4384,N_294,N_2136);
xnor U4385 (N_4385,N_2381,N_876);
or U4386 (N_4386,N_1382,N_2132);
xnor U4387 (N_4387,N_1060,N_1386);
nor U4388 (N_4388,N_1465,N_2023);
and U4389 (N_4389,N_1353,N_1061);
nand U4390 (N_4390,N_847,N_1435);
or U4391 (N_4391,N_2395,N_1515);
xor U4392 (N_4392,N_683,N_1432);
or U4393 (N_4393,N_2373,N_1796);
or U4394 (N_4394,N_732,N_1910);
xor U4395 (N_4395,N_2433,N_1135);
nand U4396 (N_4396,N_817,N_334);
nand U4397 (N_4397,N_2032,N_1453);
xnor U4398 (N_4398,N_1278,N_1402);
nor U4399 (N_4399,N_715,N_1418);
or U4400 (N_4400,N_684,N_1881);
nand U4401 (N_4401,N_2404,N_1031);
xnor U4402 (N_4402,N_2122,N_93);
xnor U4403 (N_4403,N_1132,N_1472);
and U4404 (N_4404,N_202,N_294);
xor U4405 (N_4405,N_2323,N_1356);
nand U4406 (N_4406,N_1635,N_2490);
nor U4407 (N_4407,N_671,N_1609);
or U4408 (N_4408,N_2213,N_884);
or U4409 (N_4409,N_1932,N_1138);
or U4410 (N_4410,N_1118,N_1002);
xnor U4411 (N_4411,N_601,N_1420);
and U4412 (N_4412,N_821,N_402);
and U4413 (N_4413,N_2064,N_110);
and U4414 (N_4414,N_2015,N_795);
xnor U4415 (N_4415,N_883,N_1710);
nand U4416 (N_4416,N_2330,N_145);
or U4417 (N_4417,N_1345,N_64);
xnor U4418 (N_4418,N_930,N_2261);
and U4419 (N_4419,N_1879,N_1593);
and U4420 (N_4420,N_1817,N_1498);
nor U4421 (N_4421,N_2067,N_1105);
and U4422 (N_4422,N_2478,N_60);
and U4423 (N_4423,N_1535,N_2379);
and U4424 (N_4424,N_408,N_2004);
xnor U4425 (N_4425,N_1614,N_2236);
or U4426 (N_4426,N_945,N_2252);
and U4427 (N_4427,N_456,N_1960);
nor U4428 (N_4428,N_223,N_1655);
nor U4429 (N_4429,N_1291,N_31);
or U4430 (N_4430,N_42,N_318);
and U4431 (N_4431,N_977,N_1872);
xnor U4432 (N_4432,N_1282,N_1738);
nor U4433 (N_4433,N_583,N_1464);
xor U4434 (N_4434,N_627,N_1090);
nor U4435 (N_4435,N_803,N_2259);
xor U4436 (N_4436,N_1003,N_597);
or U4437 (N_4437,N_223,N_1920);
or U4438 (N_4438,N_1947,N_2112);
xor U4439 (N_4439,N_553,N_1564);
nor U4440 (N_4440,N_1946,N_821);
nor U4441 (N_4441,N_2317,N_812);
or U4442 (N_4442,N_2177,N_1676);
xor U4443 (N_4443,N_48,N_1235);
or U4444 (N_4444,N_2102,N_1363);
nand U4445 (N_4445,N_1976,N_53);
and U4446 (N_4446,N_1585,N_1683);
or U4447 (N_4447,N_1826,N_1214);
nor U4448 (N_4448,N_1393,N_1781);
and U4449 (N_4449,N_320,N_288);
xnor U4450 (N_4450,N_818,N_2396);
nand U4451 (N_4451,N_2246,N_1239);
xor U4452 (N_4452,N_112,N_161);
and U4453 (N_4453,N_177,N_1609);
nand U4454 (N_4454,N_1649,N_1519);
or U4455 (N_4455,N_583,N_1275);
and U4456 (N_4456,N_2374,N_579);
or U4457 (N_4457,N_228,N_2418);
nor U4458 (N_4458,N_1733,N_289);
nand U4459 (N_4459,N_140,N_2025);
nand U4460 (N_4460,N_501,N_843);
nand U4461 (N_4461,N_1707,N_1096);
xnor U4462 (N_4462,N_2382,N_1895);
nand U4463 (N_4463,N_332,N_1120);
nor U4464 (N_4464,N_1378,N_1169);
nor U4465 (N_4465,N_1630,N_1980);
or U4466 (N_4466,N_2319,N_1236);
nor U4467 (N_4467,N_982,N_2485);
nor U4468 (N_4468,N_2264,N_2376);
nor U4469 (N_4469,N_380,N_928);
nand U4470 (N_4470,N_2253,N_692);
nor U4471 (N_4471,N_1761,N_875);
and U4472 (N_4472,N_2071,N_112);
nand U4473 (N_4473,N_1850,N_1148);
and U4474 (N_4474,N_2293,N_62);
nand U4475 (N_4475,N_822,N_2457);
nor U4476 (N_4476,N_802,N_989);
nand U4477 (N_4477,N_2007,N_740);
xor U4478 (N_4478,N_797,N_431);
xnor U4479 (N_4479,N_1305,N_906);
and U4480 (N_4480,N_1355,N_1672);
nand U4481 (N_4481,N_2077,N_176);
or U4482 (N_4482,N_1551,N_384);
or U4483 (N_4483,N_2121,N_1934);
nand U4484 (N_4484,N_240,N_830);
nand U4485 (N_4485,N_2062,N_476);
nor U4486 (N_4486,N_82,N_2400);
xnor U4487 (N_4487,N_2286,N_2427);
nand U4488 (N_4488,N_1581,N_1707);
xor U4489 (N_4489,N_1632,N_1913);
xor U4490 (N_4490,N_1811,N_2362);
nor U4491 (N_4491,N_1985,N_2020);
nor U4492 (N_4492,N_2312,N_1867);
nor U4493 (N_4493,N_2431,N_1074);
nor U4494 (N_4494,N_1592,N_407);
and U4495 (N_4495,N_754,N_1975);
nor U4496 (N_4496,N_2072,N_973);
xor U4497 (N_4497,N_42,N_189);
xnor U4498 (N_4498,N_1277,N_406);
nor U4499 (N_4499,N_424,N_1240);
or U4500 (N_4500,N_2145,N_1671);
xor U4501 (N_4501,N_1777,N_86);
xnor U4502 (N_4502,N_1625,N_1773);
nand U4503 (N_4503,N_2109,N_2374);
or U4504 (N_4504,N_2385,N_320);
nor U4505 (N_4505,N_2278,N_1730);
or U4506 (N_4506,N_300,N_352);
nor U4507 (N_4507,N_1136,N_960);
or U4508 (N_4508,N_2316,N_743);
nor U4509 (N_4509,N_228,N_1719);
nand U4510 (N_4510,N_180,N_942);
nor U4511 (N_4511,N_557,N_372);
nor U4512 (N_4512,N_1886,N_1440);
or U4513 (N_4513,N_2368,N_1812);
nand U4514 (N_4514,N_1579,N_1450);
xnor U4515 (N_4515,N_106,N_991);
and U4516 (N_4516,N_931,N_87);
nand U4517 (N_4517,N_73,N_82);
and U4518 (N_4518,N_1355,N_378);
nor U4519 (N_4519,N_26,N_2354);
nand U4520 (N_4520,N_1675,N_946);
xor U4521 (N_4521,N_1989,N_2325);
or U4522 (N_4522,N_1128,N_2003);
or U4523 (N_4523,N_2164,N_727);
nor U4524 (N_4524,N_68,N_896);
and U4525 (N_4525,N_269,N_2144);
nand U4526 (N_4526,N_1450,N_1527);
or U4527 (N_4527,N_1229,N_1206);
xor U4528 (N_4528,N_1052,N_1447);
and U4529 (N_4529,N_116,N_1682);
and U4530 (N_4530,N_1165,N_298);
or U4531 (N_4531,N_329,N_209);
and U4532 (N_4532,N_948,N_651);
xor U4533 (N_4533,N_1115,N_70);
or U4534 (N_4534,N_2320,N_564);
and U4535 (N_4535,N_915,N_1827);
nand U4536 (N_4536,N_844,N_1261);
nor U4537 (N_4537,N_339,N_1795);
or U4538 (N_4538,N_2154,N_708);
nor U4539 (N_4539,N_691,N_229);
nor U4540 (N_4540,N_395,N_2413);
nand U4541 (N_4541,N_2448,N_1352);
xor U4542 (N_4542,N_664,N_179);
xor U4543 (N_4543,N_2047,N_1702);
and U4544 (N_4544,N_1300,N_2282);
or U4545 (N_4545,N_698,N_294);
nand U4546 (N_4546,N_1419,N_1996);
nand U4547 (N_4547,N_139,N_1729);
nor U4548 (N_4548,N_1522,N_153);
nand U4549 (N_4549,N_1275,N_1948);
nor U4550 (N_4550,N_1408,N_1079);
and U4551 (N_4551,N_1984,N_1330);
xnor U4552 (N_4552,N_1415,N_1501);
nor U4553 (N_4553,N_541,N_1869);
and U4554 (N_4554,N_527,N_2166);
or U4555 (N_4555,N_2046,N_2069);
xor U4556 (N_4556,N_988,N_874);
nand U4557 (N_4557,N_891,N_2303);
xor U4558 (N_4558,N_1390,N_2259);
nand U4559 (N_4559,N_1186,N_907);
nor U4560 (N_4560,N_360,N_2110);
nand U4561 (N_4561,N_1739,N_2076);
and U4562 (N_4562,N_2206,N_0);
and U4563 (N_4563,N_509,N_622);
xor U4564 (N_4564,N_1559,N_2459);
and U4565 (N_4565,N_2363,N_654);
nand U4566 (N_4566,N_2240,N_1550);
xor U4567 (N_4567,N_7,N_1562);
nand U4568 (N_4568,N_1620,N_1064);
nor U4569 (N_4569,N_1110,N_445);
or U4570 (N_4570,N_1173,N_437);
and U4571 (N_4571,N_686,N_733);
and U4572 (N_4572,N_36,N_1047);
and U4573 (N_4573,N_221,N_723);
nor U4574 (N_4574,N_35,N_387);
xnor U4575 (N_4575,N_2169,N_468);
or U4576 (N_4576,N_1653,N_231);
nand U4577 (N_4577,N_1468,N_2470);
xor U4578 (N_4578,N_2348,N_131);
and U4579 (N_4579,N_161,N_2125);
nor U4580 (N_4580,N_2022,N_2285);
xor U4581 (N_4581,N_1553,N_1463);
or U4582 (N_4582,N_1392,N_1816);
and U4583 (N_4583,N_41,N_498);
nor U4584 (N_4584,N_968,N_459);
or U4585 (N_4585,N_1855,N_2335);
nand U4586 (N_4586,N_1877,N_669);
xor U4587 (N_4587,N_1783,N_335);
xnor U4588 (N_4588,N_1140,N_1014);
nand U4589 (N_4589,N_1000,N_2356);
nand U4590 (N_4590,N_960,N_302);
nor U4591 (N_4591,N_199,N_464);
xor U4592 (N_4592,N_2013,N_469);
or U4593 (N_4593,N_993,N_843);
xnor U4594 (N_4594,N_1742,N_1277);
xnor U4595 (N_4595,N_1918,N_455);
and U4596 (N_4596,N_25,N_2370);
xor U4597 (N_4597,N_1568,N_1373);
and U4598 (N_4598,N_1126,N_1013);
nor U4599 (N_4599,N_21,N_340);
xor U4600 (N_4600,N_2171,N_1285);
nor U4601 (N_4601,N_1480,N_1074);
xor U4602 (N_4602,N_1757,N_2187);
and U4603 (N_4603,N_1456,N_235);
and U4604 (N_4604,N_1328,N_605);
xnor U4605 (N_4605,N_1507,N_1212);
xnor U4606 (N_4606,N_475,N_41);
xnor U4607 (N_4607,N_1913,N_793);
and U4608 (N_4608,N_950,N_1878);
and U4609 (N_4609,N_1429,N_986);
and U4610 (N_4610,N_414,N_1022);
or U4611 (N_4611,N_1889,N_2472);
and U4612 (N_4612,N_955,N_2148);
nor U4613 (N_4613,N_1275,N_523);
or U4614 (N_4614,N_1646,N_696);
and U4615 (N_4615,N_1365,N_297);
nand U4616 (N_4616,N_1819,N_684);
and U4617 (N_4617,N_2267,N_1189);
xnor U4618 (N_4618,N_1775,N_2357);
nor U4619 (N_4619,N_1273,N_1142);
nor U4620 (N_4620,N_1759,N_848);
or U4621 (N_4621,N_264,N_1805);
or U4622 (N_4622,N_1872,N_2471);
xnor U4623 (N_4623,N_349,N_1024);
and U4624 (N_4624,N_636,N_55);
and U4625 (N_4625,N_627,N_1138);
nor U4626 (N_4626,N_1210,N_1112);
or U4627 (N_4627,N_1414,N_857);
xnor U4628 (N_4628,N_1835,N_1401);
or U4629 (N_4629,N_354,N_1615);
and U4630 (N_4630,N_235,N_2167);
or U4631 (N_4631,N_236,N_1697);
and U4632 (N_4632,N_2155,N_2459);
nor U4633 (N_4633,N_339,N_241);
xor U4634 (N_4634,N_1291,N_922);
nor U4635 (N_4635,N_206,N_2453);
and U4636 (N_4636,N_828,N_1365);
nand U4637 (N_4637,N_996,N_1058);
xnor U4638 (N_4638,N_681,N_62);
nand U4639 (N_4639,N_1630,N_1943);
and U4640 (N_4640,N_1774,N_1887);
nand U4641 (N_4641,N_1573,N_1842);
nand U4642 (N_4642,N_1036,N_1563);
nand U4643 (N_4643,N_1864,N_2104);
or U4644 (N_4644,N_1625,N_1385);
and U4645 (N_4645,N_984,N_1373);
nor U4646 (N_4646,N_950,N_309);
and U4647 (N_4647,N_699,N_1029);
xor U4648 (N_4648,N_1732,N_1619);
xor U4649 (N_4649,N_127,N_791);
or U4650 (N_4650,N_1128,N_1893);
or U4651 (N_4651,N_79,N_1943);
nand U4652 (N_4652,N_748,N_1639);
or U4653 (N_4653,N_1594,N_1444);
nand U4654 (N_4654,N_315,N_1617);
and U4655 (N_4655,N_2219,N_905);
and U4656 (N_4656,N_811,N_801);
and U4657 (N_4657,N_401,N_1910);
nand U4658 (N_4658,N_1904,N_2415);
and U4659 (N_4659,N_1867,N_1816);
xnor U4660 (N_4660,N_911,N_309);
and U4661 (N_4661,N_2404,N_972);
nand U4662 (N_4662,N_1927,N_221);
nand U4663 (N_4663,N_61,N_1501);
and U4664 (N_4664,N_1686,N_2481);
nand U4665 (N_4665,N_1871,N_516);
or U4666 (N_4666,N_1797,N_1035);
nand U4667 (N_4667,N_492,N_125);
nand U4668 (N_4668,N_1929,N_638);
nand U4669 (N_4669,N_6,N_1237);
nand U4670 (N_4670,N_1249,N_941);
and U4671 (N_4671,N_738,N_423);
or U4672 (N_4672,N_1593,N_490);
nor U4673 (N_4673,N_2263,N_1285);
or U4674 (N_4674,N_1507,N_1566);
or U4675 (N_4675,N_1287,N_1419);
and U4676 (N_4676,N_1523,N_735);
and U4677 (N_4677,N_1092,N_183);
nor U4678 (N_4678,N_2219,N_1229);
or U4679 (N_4679,N_427,N_1656);
or U4680 (N_4680,N_2003,N_351);
xor U4681 (N_4681,N_1694,N_2449);
nand U4682 (N_4682,N_762,N_1247);
xnor U4683 (N_4683,N_229,N_2215);
or U4684 (N_4684,N_1094,N_1685);
nand U4685 (N_4685,N_540,N_284);
xnor U4686 (N_4686,N_1569,N_1559);
nor U4687 (N_4687,N_2011,N_2169);
xnor U4688 (N_4688,N_482,N_2130);
nor U4689 (N_4689,N_281,N_1784);
and U4690 (N_4690,N_314,N_1204);
nand U4691 (N_4691,N_1223,N_2322);
nor U4692 (N_4692,N_527,N_2291);
xnor U4693 (N_4693,N_1657,N_498);
or U4694 (N_4694,N_1155,N_2203);
and U4695 (N_4695,N_1660,N_390);
nand U4696 (N_4696,N_1031,N_2035);
or U4697 (N_4697,N_714,N_1892);
xor U4698 (N_4698,N_1191,N_4);
nor U4699 (N_4699,N_2272,N_1527);
nand U4700 (N_4700,N_16,N_1546);
nor U4701 (N_4701,N_1478,N_821);
xor U4702 (N_4702,N_2481,N_316);
or U4703 (N_4703,N_2331,N_218);
xnor U4704 (N_4704,N_1655,N_1324);
or U4705 (N_4705,N_1322,N_971);
and U4706 (N_4706,N_573,N_771);
or U4707 (N_4707,N_1118,N_1217);
or U4708 (N_4708,N_1121,N_302);
nor U4709 (N_4709,N_223,N_2164);
nor U4710 (N_4710,N_1524,N_39);
and U4711 (N_4711,N_503,N_1126);
xnor U4712 (N_4712,N_2380,N_2456);
nor U4713 (N_4713,N_163,N_1286);
xor U4714 (N_4714,N_1960,N_531);
or U4715 (N_4715,N_1748,N_2435);
xor U4716 (N_4716,N_2490,N_1646);
and U4717 (N_4717,N_761,N_1161);
nor U4718 (N_4718,N_1684,N_2491);
nand U4719 (N_4719,N_2488,N_347);
nand U4720 (N_4720,N_88,N_1108);
and U4721 (N_4721,N_2338,N_98);
nor U4722 (N_4722,N_2415,N_158);
xnor U4723 (N_4723,N_820,N_2065);
nor U4724 (N_4724,N_331,N_2006);
xor U4725 (N_4725,N_1093,N_2477);
xor U4726 (N_4726,N_1713,N_2067);
or U4727 (N_4727,N_1303,N_181);
or U4728 (N_4728,N_386,N_1150);
and U4729 (N_4729,N_1427,N_155);
xor U4730 (N_4730,N_1675,N_2165);
nor U4731 (N_4731,N_606,N_1758);
and U4732 (N_4732,N_2001,N_1179);
xor U4733 (N_4733,N_2211,N_309);
and U4734 (N_4734,N_900,N_1042);
and U4735 (N_4735,N_2154,N_962);
and U4736 (N_4736,N_2479,N_1127);
and U4737 (N_4737,N_351,N_17);
xor U4738 (N_4738,N_1767,N_345);
xor U4739 (N_4739,N_658,N_1172);
or U4740 (N_4740,N_1871,N_742);
or U4741 (N_4741,N_399,N_1771);
nand U4742 (N_4742,N_2037,N_2110);
xnor U4743 (N_4743,N_1356,N_838);
nand U4744 (N_4744,N_605,N_966);
xor U4745 (N_4745,N_186,N_368);
and U4746 (N_4746,N_455,N_1384);
nand U4747 (N_4747,N_1569,N_2019);
nand U4748 (N_4748,N_1095,N_2420);
nand U4749 (N_4749,N_1956,N_1089);
and U4750 (N_4750,N_1879,N_1365);
or U4751 (N_4751,N_1463,N_1675);
xor U4752 (N_4752,N_908,N_1241);
xnor U4753 (N_4753,N_2287,N_2305);
and U4754 (N_4754,N_1941,N_1798);
nor U4755 (N_4755,N_1253,N_1460);
xor U4756 (N_4756,N_704,N_157);
nor U4757 (N_4757,N_928,N_2132);
xor U4758 (N_4758,N_370,N_707);
or U4759 (N_4759,N_2239,N_568);
nor U4760 (N_4760,N_1616,N_373);
nand U4761 (N_4761,N_35,N_1212);
and U4762 (N_4762,N_1897,N_1075);
nand U4763 (N_4763,N_1435,N_1215);
or U4764 (N_4764,N_1576,N_2432);
or U4765 (N_4765,N_1460,N_1744);
and U4766 (N_4766,N_658,N_253);
nor U4767 (N_4767,N_564,N_906);
nor U4768 (N_4768,N_1303,N_597);
nor U4769 (N_4769,N_275,N_1185);
or U4770 (N_4770,N_2275,N_2082);
xor U4771 (N_4771,N_91,N_1001);
nor U4772 (N_4772,N_2155,N_2014);
nand U4773 (N_4773,N_438,N_2147);
or U4774 (N_4774,N_662,N_2465);
and U4775 (N_4775,N_2117,N_2247);
and U4776 (N_4776,N_1974,N_415);
xor U4777 (N_4777,N_2334,N_375);
and U4778 (N_4778,N_2025,N_1721);
nor U4779 (N_4779,N_2001,N_2473);
or U4780 (N_4780,N_2267,N_1447);
or U4781 (N_4781,N_1332,N_404);
and U4782 (N_4782,N_1557,N_1642);
nor U4783 (N_4783,N_266,N_1166);
and U4784 (N_4784,N_224,N_1674);
or U4785 (N_4785,N_1043,N_489);
xor U4786 (N_4786,N_2099,N_973);
nor U4787 (N_4787,N_1266,N_350);
nand U4788 (N_4788,N_862,N_652);
or U4789 (N_4789,N_205,N_1082);
xnor U4790 (N_4790,N_798,N_1876);
xor U4791 (N_4791,N_319,N_2137);
and U4792 (N_4792,N_2448,N_684);
xor U4793 (N_4793,N_500,N_2139);
xor U4794 (N_4794,N_1583,N_1434);
nand U4795 (N_4795,N_1436,N_960);
nand U4796 (N_4796,N_2352,N_1716);
and U4797 (N_4797,N_74,N_282);
and U4798 (N_4798,N_1604,N_1471);
nand U4799 (N_4799,N_738,N_492);
or U4800 (N_4800,N_822,N_2258);
or U4801 (N_4801,N_1265,N_1551);
or U4802 (N_4802,N_1072,N_595);
or U4803 (N_4803,N_1025,N_665);
xor U4804 (N_4804,N_2421,N_792);
xnor U4805 (N_4805,N_967,N_76);
or U4806 (N_4806,N_1098,N_742);
nor U4807 (N_4807,N_2285,N_1516);
or U4808 (N_4808,N_2405,N_2184);
xor U4809 (N_4809,N_204,N_283);
xor U4810 (N_4810,N_1666,N_2286);
and U4811 (N_4811,N_692,N_1712);
and U4812 (N_4812,N_1725,N_2498);
nor U4813 (N_4813,N_2457,N_372);
nor U4814 (N_4814,N_2456,N_1050);
nand U4815 (N_4815,N_463,N_1972);
or U4816 (N_4816,N_1644,N_921);
or U4817 (N_4817,N_1516,N_648);
or U4818 (N_4818,N_774,N_629);
nand U4819 (N_4819,N_446,N_2184);
nor U4820 (N_4820,N_16,N_272);
and U4821 (N_4821,N_1793,N_25);
or U4822 (N_4822,N_1735,N_1292);
or U4823 (N_4823,N_1028,N_2363);
nand U4824 (N_4824,N_1880,N_2114);
or U4825 (N_4825,N_1917,N_1220);
or U4826 (N_4826,N_1461,N_1157);
nand U4827 (N_4827,N_1461,N_762);
and U4828 (N_4828,N_174,N_1422);
or U4829 (N_4829,N_1082,N_2108);
nor U4830 (N_4830,N_335,N_391);
and U4831 (N_4831,N_2,N_1208);
nand U4832 (N_4832,N_1863,N_1137);
nand U4833 (N_4833,N_2110,N_898);
and U4834 (N_4834,N_1551,N_2318);
and U4835 (N_4835,N_1679,N_897);
nor U4836 (N_4836,N_1784,N_367);
and U4837 (N_4837,N_1122,N_904);
or U4838 (N_4838,N_993,N_368);
xnor U4839 (N_4839,N_1021,N_902);
and U4840 (N_4840,N_2095,N_732);
and U4841 (N_4841,N_2328,N_765);
nand U4842 (N_4842,N_662,N_738);
xnor U4843 (N_4843,N_841,N_927);
nand U4844 (N_4844,N_2016,N_2476);
and U4845 (N_4845,N_1637,N_1544);
xnor U4846 (N_4846,N_1812,N_2478);
nand U4847 (N_4847,N_245,N_1868);
or U4848 (N_4848,N_905,N_681);
nand U4849 (N_4849,N_316,N_1067);
xor U4850 (N_4850,N_396,N_1873);
nor U4851 (N_4851,N_365,N_1322);
nand U4852 (N_4852,N_929,N_60);
and U4853 (N_4853,N_1124,N_784);
xor U4854 (N_4854,N_508,N_1000);
nor U4855 (N_4855,N_308,N_666);
xor U4856 (N_4856,N_466,N_1165);
nand U4857 (N_4857,N_11,N_490);
nand U4858 (N_4858,N_599,N_1583);
nand U4859 (N_4859,N_1459,N_1712);
xnor U4860 (N_4860,N_1963,N_2470);
nor U4861 (N_4861,N_227,N_2322);
xnor U4862 (N_4862,N_2439,N_314);
nor U4863 (N_4863,N_584,N_1756);
and U4864 (N_4864,N_827,N_1763);
or U4865 (N_4865,N_1863,N_403);
or U4866 (N_4866,N_1822,N_96);
nand U4867 (N_4867,N_1635,N_833);
or U4868 (N_4868,N_255,N_771);
and U4869 (N_4869,N_2056,N_171);
xor U4870 (N_4870,N_1031,N_682);
and U4871 (N_4871,N_360,N_1413);
or U4872 (N_4872,N_670,N_994);
nor U4873 (N_4873,N_710,N_881);
or U4874 (N_4874,N_1132,N_302);
nor U4875 (N_4875,N_393,N_1519);
and U4876 (N_4876,N_1867,N_627);
or U4877 (N_4877,N_674,N_2131);
xor U4878 (N_4878,N_128,N_1781);
or U4879 (N_4879,N_422,N_1537);
or U4880 (N_4880,N_1369,N_1117);
xnor U4881 (N_4881,N_2439,N_2190);
or U4882 (N_4882,N_730,N_1728);
and U4883 (N_4883,N_1173,N_1159);
nand U4884 (N_4884,N_763,N_166);
and U4885 (N_4885,N_1385,N_2337);
nand U4886 (N_4886,N_8,N_7);
nand U4887 (N_4887,N_137,N_604);
or U4888 (N_4888,N_2375,N_1459);
and U4889 (N_4889,N_2394,N_12);
nand U4890 (N_4890,N_805,N_2478);
nand U4891 (N_4891,N_991,N_278);
and U4892 (N_4892,N_1960,N_2428);
nor U4893 (N_4893,N_1591,N_2204);
or U4894 (N_4894,N_1842,N_2473);
nand U4895 (N_4895,N_803,N_1583);
or U4896 (N_4896,N_1749,N_450);
nor U4897 (N_4897,N_682,N_1007);
nor U4898 (N_4898,N_1792,N_2067);
or U4899 (N_4899,N_2441,N_1897);
xnor U4900 (N_4900,N_1815,N_824);
and U4901 (N_4901,N_920,N_1449);
nor U4902 (N_4902,N_8,N_1866);
nand U4903 (N_4903,N_1298,N_1621);
nand U4904 (N_4904,N_144,N_1487);
nand U4905 (N_4905,N_2239,N_754);
nor U4906 (N_4906,N_315,N_1305);
nand U4907 (N_4907,N_1230,N_2189);
or U4908 (N_4908,N_1455,N_1642);
or U4909 (N_4909,N_778,N_2435);
nand U4910 (N_4910,N_803,N_987);
nor U4911 (N_4911,N_1274,N_1821);
nor U4912 (N_4912,N_488,N_953);
and U4913 (N_4913,N_1202,N_1938);
and U4914 (N_4914,N_2156,N_1421);
or U4915 (N_4915,N_588,N_445);
nand U4916 (N_4916,N_893,N_1379);
nor U4917 (N_4917,N_1188,N_933);
xor U4918 (N_4918,N_1359,N_721);
and U4919 (N_4919,N_2079,N_2390);
xor U4920 (N_4920,N_1163,N_1374);
xor U4921 (N_4921,N_1541,N_735);
or U4922 (N_4922,N_2246,N_501);
nand U4923 (N_4923,N_1832,N_2033);
and U4924 (N_4924,N_446,N_1086);
nand U4925 (N_4925,N_325,N_490);
and U4926 (N_4926,N_2084,N_2234);
nand U4927 (N_4927,N_942,N_1304);
nand U4928 (N_4928,N_1710,N_2219);
nor U4929 (N_4929,N_804,N_1641);
and U4930 (N_4930,N_764,N_938);
xnor U4931 (N_4931,N_1853,N_2047);
nand U4932 (N_4932,N_2160,N_2175);
and U4933 (N_4933,N_1918,N_2487);
and U4934 (N_4934,N_2057,N_2127);
xnor U4935 (N_4935,N_587,N_102);
or U4936 (N_4936,N_1019,N_0);
or U4937 (N_4937,N_1056,N_657);
nand U4938 (N_4938,N_1247,N_2411);
and U4939 (N_4939,N_700,N_1826);
or U4940 (N_4940,N_391,N_169);
nand U4941 (N_4941,N_231,N_1907);
nor U4942 (N_4942,N_1713,N_1096);
nand U4943 (N_4943,N_1737,N_1575);
or U4944 (N_4944,N_1143,N_258);
xor U4945 (N_4945,N_944,N_1588);
nor U4946 (N_4946,N_1947,N_1681);
or U4947 (N_4947,N_2288,N_748);
nor U4948 (N_4948,N_1708,N_2188);
and U4949 (N_4949,N_2414,N_909);
nor U4950 (N_4950,N_72,N_1021);
and U4951 (N_4951,N_765,N_2319);
xor U4952 (N_4952,N_15,N_2169);
or U4953 (N_4953,N_893,N_933);
or U4954 (N_4954,N_2420,N_2273);
and U4955 (N_4955,N_1163,N_955);
or U4956 (N_4956,N_1056,N_533);
nor U4957 (N_4957,N_186,N_884);
xnor U4958 (N_4958,N_1715,N_2278);
and U4959 (N_4959,N_891,N_628);
nand U4960 (N_4960,N_1377,N_282);
or U4961 (N_4961,N_355,N_2277);
nor U4962 (N_4962,N_1543,N_2365);
xor U4963 (N_4963,N_551,N_1996);
nand U4964 (N_4964,N_1530,N_763);
nor U4965 (N_4965,N_1739,N_167);
or U4966 (N_4966,N_7,N_1180);
nor U4967 (N_4967,N_224,N_211);
or U4968 (N_4968,N_128,N_894);
xnor U4969 (N_4969,N_668,N_952);
nand U4970 (N_4970,N_486,N_450);
xnor U4971 (N_4971,N_2059,N_2305);
xor U4972 (N_4972,N_883,N_2108);
nor U4973 (N_4973,N_612,N_1002);
and U4974 (N_4974,N_1949,N_1505);
and U4975 (N_4975,N_304,N_834);
xor U4976 (N_4976,N_1923,N_961);
nand U4977 (N_4977,N_1673,N_1573);
and U4978 (N_4978,N_397,N_151);
nor U4979 (N_4979,N_1752,N_1610);
and U4980 (N_4980,N_1859,N_732);
nand U4981 (N_4981,N_49,N_67);
and U4982 (N_4982,N_355,N_320);
or U4983 (N_4983,N_1943,N_80);
nand U4984 (N_4984,N_123,N_1283);
and U4985 (N_4985,N_1205,N_2086);
and U4986 (N_4986,N_451,N_584);
or U4987 (N_4987,N_2467,N_171);
nand U4988 (N_4988,N_1858,N_2129);
or U4989 (N_4989,N_2274,N_760);
and U4990 (N_4990,N_63,N_1725);
or U4991 (N_4991,N_494,N_2035);
xor U4992 (N_4992,N_1348,N_1251);
or U4993 (N_4993,N_1981,N_1041);
xor U4994 (N_4994,N_283,N_1726);
and U4995 (N_4995,N_1227,N_1807);
xor U4996 (N_4996,N_652,N_224);
or U4997 (N_4997,N_1298,N_2493);
nand U4998 (N_4998,N_2223,N_24);
or U4999 (N_4999,N_2238,N_327);
and U5000 (N_5000,N_4941,N_4651);
xnor U5001 (N_5001,N_4442,N_4504);
nor U5002 (N_5002,N_4301,N_4893);
nor U5003 (N_5003,N_4699,N_2719);
or U5004 (N_5004,N_4053,N_4878);
and U5005 (N_5005,N_2546,N_3155);
nand U5006 (N_5006,N_4282,N_4915);
and U5007 (N_5007,N_3739,N_4805);
xor U5008 (N_5008,N_2600,N_4338);
nand U5009 (N_5009,N_4686,N_3250);
xnor U5010 (N_5010,N_2873,N_3227);
or U5011 (N_5011,N_4593,N_4585);
nand U5012 (N_5012,N_3210,N_3955);
or U5013 (N_5013,N_3008,N_4355);
or U5014 (N_5014,N_2889,N_2895);
or U5015 (N_5015,N_4302,N_3132);
or U5016 (N_5016,N_3542,N_2678);
nor U5017 (N_5017,N_3658,N_4682);
and U5018 (N_5018,N_3574,N_3017);
or U5019 (N_5019,N_4044,N_2589);
nor U5020 (N_5020,N_4503,N_3254);
or U5021 (N_5021,N_3539,N_3570);
or U5022 (N_5022,N_4760,N_4165);
xor U5023 (N_5023,N_3727,N_4909);
xnor U5024 (N_5024,N_4020,N_3631);
or U5025 (N_5025,N_2676,N_4841);
and U5026 (N_5026,N_4179,N_4101);
nand U5027 (N_5027,N_4074,N_2721);
or U5028 (N_5028,N_3908,N_3113);
or U5029 (N_5029,N_4931,N_2745);
or U5030 (N_5030,N_3255,N_3364);
xor U5031 (N_5031,N_4641,N_4278);
nand U5032 (N_5032,N_3275,N_2919);
or U5033 (N_5033,N_3597,N_4709);
nor U5034 (N_5034,N_2624,N_3147);
xnor U5035 (N_5035,N_3737,N_3645);
nand U5036 (N_5036,N_3029,N_3318);
nand U5037 (N_5037,N_2630,N_4266);
xnor U5038 (N_5038,N_4605,N_4362);
xnor U5039 (N_5039,N_4779,N_3948);
xnor U5040 (N_5040,N_2775,N_3891);
and U5041 (N_5041,N_3368,N_4449);
or U5042 (N_5042,N_4528,N_4057);
or U5043 (N_5043,N_4562,N_2541);
xor U5044 (N_5044,N_3315,N_3386);
xnor U5045 (N_5045,N_3650,N_3199);
or U5046 (N_5046,N_4914,N_4412);
and U5047 (N_5047,N_2901,N_4293);
and U5048 (N_5048,N_4437,N_3712);
and U5049 (N_5049,N_3102,N_4444);
and U5050 (N_5050,N_4396,N_4778);
xnor U5051 (N_5051,N_4887,N_3095);
xor U5052 (N_5052,N_3310,N_4588);
and U5053 (N_5053,N_3377,N_2662);
xnor U5054 (N_5054,N_2864,N_3871);
or U5055 (N_5055,N_2565,N_4537);
xnor U5056 (N_5056,N_2569,N_3897);
nor U5057 (N_5057,N_4352,N_3838);
and U5058 (N_5058,N_4190,N_4256);
xor U5059 (N_5059,N_4094,N_3163);
and U5060 (N_5060,N_4481,N_2759);
and U5061 (N_5061,N_3634,N_3917);
and U5062 (N_5062,N_2982,N_4617);
nand U5063 (N_5063,N_3929,N_4634);
nor U5064 (N_5064,N_4785,N_3359);
nand U5065 (N_5065,N_4730,N_3333);
and U5066 (N_5066,N_3054,N_4988);
nand U5067 (N_5067,N_4400,N_4142);
nor U5068 (N_5068,N_2968,N_4843);
or U5069 (N_5069,N_2900,N_4246);
and U5070 (N_5070,N_3313,N_2955);
xnor U5071 (N_5071,N_4599,N_3282);
nand U5072 (N_5072,N_3443,N_4765);
xnor U5073 (N_5073,N_2620,N_3938);
or U5074 (N_5074,N_3477,N_3679);
or U5075 (N_5075,N_4243,N_3060);
or U5076 (N_5076,N_4073,N_4337);
or U5077 (N_5077,N_3793,N_4918);
nand U5078 (N_5078,N_2707,N_3661);
nand U5079 (N_5079,N_2844,N_4772);
xor U5080 (N_5080,N_4536,N_4509);
nor U5081 (N_5081,N_3302,N_4812);
nor U5082 (N_5082,N_3503,N_3910);
and U5083 (N_5083,N_2856,N_2553);
nor U5084 (N_5084,N_4786,N_4761);
or U5085 (N_5085,N_3669,N_4114);
nand U5086 (N_5086,N_4565,N_4307);
xnor U5087 (N_5087,N_4674,N_4450);
nand U5088 (N_5088,N_4203,N_3906);
xnor U5089 (N_5089,N_4678,N_3374);
and U5090 (N_5090,N_2803,N_3342);
or U5091 (N_5091,N_3493,N_2796);
nand U5092 (N_5092,N_4006,N_2659);
xor U5093 (N_5093,N_2785,N_2742);
nor U5094 (N_5094,N_3206,N_4410);
nand U5095 (N_5095,N_3211,N_3852);
and U5096 (N_5096,N_3492,N_3235);
or U5097 (N_5097,N_3200,N_4137);
nand U5098 (N_5098,N_4220,N_4152);
xnor U5099 (N_5099,N_2886,N_3548);
nand U5100 (N_5100,N_3144,N_3077);
nor U5101 (N_5101,N_4622,N_3516);
xnor U5102 (N_5102,N_4694,N_3911);
and U5103 (N_5103,N_4126,N_4557);
nor U5104 (N_5104,N_3828,N_3191);
nor U5105 (N_5105,N_4616,N_3401);
xnor U5106 (N_5106,N_3009,N_3428);
nor U5107 (N_5107,N_3587,N_4321);
and U5108 (N_5108,N_4801,N_4047);
nand U5109 (N_5109,N_3786,N_4609);
nand U5110 (N_5110,N_4866,N_3016);
nor U5111 (N_5111,N_3784,N_2501);
or U5112 (N_5112,N_4690,N_4718);
nor U5113 (N_5113,N_4592,N_3892);
and U5114 (N_5114,N_3532,N_2523);
xnor U5115 (N_5115,N_3125,N_4341);
nor U5116 (N_5116,N_2947,N_3084);
nand U5117 (N_5117,N_4862,N_3152);
and U5118 (N_5118,N_4929,N_3940);
nor U5119 (N_5119,N_3703,N_4034);
or U5120 (N_5120,N_4574,N_4568);
or U5121 (N_5121,N_4238,N_3521);
and U5122 (N_5122,N_3243,N_2545);
or U5123 (N_5123,N_4250,N_2787);
xor U5124 (N_5124,N_3788,N_2832);
nand U5125 (N_5125,N_3139,N_2894);
nor U5126 (N_5126,N_4430,N_2792);
nor U5127 (N_5127,N_3482,N_4195);
nand U5128 (N_5128,N_3068,N_4169);
nand U5129 (N_5129,N_2995,N_4883);
nor U5130 (N_5130,N_4743,N_4349);
nor U5131 (N_5131,N_3122,N_3137);
nor U5132 (N_5132,N_4206,N_4403);
nor U5133 (N_5133,N_3510,N_4305);
and U5134 (N_5134,N_3716,N_4214);
or U5135 (N_5135,N_4998,N_2664);
nand U5136 (N_5136,N_3439,N_4832);
or U5137 (N_5137,N_3462,N_4040);
xor U5138 (N_5138,N_2506,N_4813);
xor U5139 (N_5139,N_2524,N_4484);
nand U5140 (N_5140,N_4402,N_4242);
and U5141 (N_5141,N_4212,N_2652);
or U5142 (N_5142,N_3434,N_4050);
or U5143 (N_5143,N_2790,N_2608);
xnor U5144 (N_5144,N_2926,N_3148);
and U5145 (N_5145,N_4940,N_4086);
xnor U5146 (N_5146,N_2529,N_3965);
and U5147 (N_5147,N_3995,N_3288);
xor U5148 (N_5148,N_2503,N_3070);
and U5149 (N_5149,N_3001,N_2776);
xnor U5150 (N_5150,N_3624,N_3447);
nor U5151 (N_5151,N_3878,N_3279);
nor U5152 (N_5152,N_3706,N_3805);
xor U5153 (N_5153,N_3021,N_4953);
nand U5154 (N_5154,N_3361,N_2964);
xnor U5155 (N_5155,N_4640,N_2879);
and U5156 (N_5156,N_4994,N_4932);
or U5157 (N_5157,N_3662,N_3641);
and U5158 (N_5158,N_3923,N_4700);
nor U5159 (N_5159,N_2944,N_2599);
nand U5160 (N_5160,N_2839,N_4719);
and U5161 (N_5161,N_3037,N_3138);
or U5162 (N_5162,N_4098,N_2603);
nand U5163 (N_5163,N_2680,N_3019);
nand U5164 (N_5164,N_2841,N_4092);
nor U5165 (N_5165,N_4561,N_3287);
nand U5166 (N_5166,N_3049,N_4159);
or U5167 (N_5167,N_2720,N_4625);
or U5168 (N_5168,N_4175,N_2863);
nor U5169 (N_5169,N_4933,N_4334);
nor U5170 (N_5170,N_4667,N_2799);
or U5171 (N_5171,N_4973,N_4011);
or U5172 (N_5172,N_4168,N_4067);
xnor U5173 (N_5173,N_2640,N_4435);
xnor U5174 (N_5174,N_2667,N_4836);
nand U5175 (N_5175,N_4368,N_4041);
nor U5176 (N_5176,N_3162,N_3689);
or U5177 (N_5177,N_4249,N_4657);
xnor U5178 (N_5178,N_4264,N_4748);
or U5179 (N_5179,N_2925,N_4001);
or U5180 (N_5180,N_3336,N_4023);
xnor U5181 (N_5181,N_3925,N_4543);
xor U5182 (N_5182,N_3142,N_3421);
or U5183 (N_5183,N_4636,N_4826);
nand U5184 (N_5184,N_2770,N_2713);
xor U5185 (N_5185,N_3329,N_4263);
and U5186 (N_5186,N_4583,N_4937);
and U5187 (N_5187,N_3502,N_3649);
nor U5188 (N_5188,N_4372,N_3121);
or U5189 (N_5189,N_4601,N_3856);
or U5190 (N_5190,N_3422,N_2972);
or U5191 (N_5191,N_3347,N_3754);
nor U5192 (N_5192,N_4275,N_3585);
or U5193 (N_5193,N_4178,N_3725);
nand U5194 (N_5194,N_2959,N_2625);
xor U5195 (N_5195,N_2973,N_3000);
and U5196 (N_5196,N_4698,N_3559);
nand U5197 (N_5197,N_4116,N_4790);
xnor U5198 (N_5198,N_3094,N_2960);
xor U5199 (N_5199,N_3078,N_2507);
nor U5200 (N_5200,N_4395,N_4376);
nor U5201 (N_5201,N_4834,N_4202);
nor U5202 (N_5202,N_3639,N_3403);
nor U5203 (N_5203,N_4024,N_3399);
nand U5204 (N_5204,N_3913,N_4956);
nand U5205 (N_5205,N_4774,N_4642);
nor U5206 (N_5206,N_4840,N_4298);
or U5207 (N_5207,N_2809,N_4677);
nor U5208 (N_5208,N_4594,N_4365);
xor U5209 (N_5209,N_4889,N_4324);
and U5210 (N_5210,N_4051,N_4144);
and U5211 (N_5211,N_3159,N_2617);
or U5212 (N_5212,N_4666,N_3905);
nand U5213 (N_5213,N_4174,N_4630);
xnor U5214 (N_5214,N_3337,N_3695);
nor U5215 (N_5215,N_4756,N_2533);
or U5216 (N_5216,N_4139,N_2797);
nor U5217 (N_5217,N_4611,N_4967);
xor U5218 (N_5218,N_3033,N_4343);
nand U5219 (N_5219,N_4469,N_3220);
or U5220 (N_5220,N_3415,N_4835);
or U5221 (N_5221,N_3188,N_2635);
and U5222 (N_5222,N_3978,N_4963);
and U5223 (N_5223,N_2777,N_2906);
nor U5224 (N_5224,N_3231,N_2666);
or U5225 (N_5225,N_4755,N_3013);
nand U5226 (N_5226,N_2717,N_4661);
nor U5227 (N_5227,N_4248,N_4171);
nor U5228 (N_5228,N_3629,N_3660);
or U5229 (N_5229,N_4035,N_4529);
nand U5230 (N_5230,N_3804,N_4415);
or U5231 (N_5231,N_4502,N_3221);
nor U5232 (N_5232,N_4229,N_3473);
xor U5233 (N_5233,N_3979,N_4454);
or U5234 (N_5234,N_4770,N_3762);
and U5235 (N_5235,N_4614,N_3930);
and U5236 (N_5236,N_3893,N_3406);
and U5237 (N_5237,N_2606,N_3463);
and U5238 (N_5238,N_3633,N_3869);
xor U5239 (N_5239,N_4042,N_3562);
xor U5240 (N_5240,N_3888,N_4087);
xnor U5241 (N_5241,N_2967,N_2774);
xnor U5242 (N_5242,N_4069,N_3720);
xor U5243 (N_5243,N_2696,N_4132);
nor U5244 (N_5244,N_3203,N_4428);
nor U5245 (N_5245,N_3396,N_2949);
or U5246 (N_5246,N_4377,N_4827);
xor U5247 (N_5247,N_4319,N_2527);
nor U5248 (N_5248,N_2808,N_3229);
or U5249 (N_5249,N_4673,N_4125);
or U5250 (N_5250,N_4331,N_4367);
nor U5251 (N_5251,N_4347,N_4946);
and U5252 (N_5252,N_2862,N_3207);
or U5253 (N_5253,N_2897,N_3290);
and U5254 (N_5254,N_3438,N_4104);
nor U5255 (N_5255,N_2851,N_4759);
and U5256 (N_5256,N_3698,N_4039);
xor U5257 (N_5257,N_2510,N_3922);
nand U5258 (N_5258,N_4731,N_3289);
or U5259 (N_5259,N_3536,N_3360);
nand U5260 (N_5260,N_3946,N_2534);
nand U5261 (N_5261,N_2555,N_3519);
nor U5262 (N_5262,N_3175,N_2789);
or U5263 (N_5263,N_2556,N_2561);
and U5264 (N_5264,N_3820,N_4131);
and U5265 (N_5265,N_4890,N_4160);
nand U5266 (N_5266,N_3864,N_3063);
nor U5267 (N_5267,N_3441,N_4392);
nand U5268 (N_5268,N_4850,N_3111);
nand U5269 (N_5269,N_3848,N_4971);
nor U5270 (N_5270,N_4414,N_4378);
and U5271 (N_5271,N_4794,N_4527);
nor U5272 (N_5272,N_4888,N_3092);
and U5273 (N_5273,N_3557,N_2802);
nor U5274 (N_5274,N_3205,N_3372);
nor U5275 (N_5275,N_3529,N_2725);
xor U5276 (N_5276,N_4285,N_2996);
or U5277 (N_5277,N_3857,N_4628);
nor U5278 (N_5278,N_4598,N_2899);
or U5279 (N_5279,N_3495,N_4992);
nor U5280 (N_5280,N_3304,N_2548);
xor U5281 (N_5281,N_4102,N_2638);
nand U5282 (N_5282,N_4310,N_4121);
or U5283 (N_5283,N_4486,N_3128);
nand U5284 (N_5284,N_4891,N_2761);
or U5285 (N_5285,N_2647,N_3116);
or U5286 (N_5286,N_3269,N_4383);
nand U5287 (N_5287,N_2512,N_3161);
nand U5288 (N_5288,N_2714,N_2646);
xnor U5289 (N_5289,N_4512,N_3627);
or U5290 (N_5290,N_2724,N_2869);
xnor U5291 (N_5291,N_3755,N_4236);
xor U5292 (N_5292,N_3898,N_3792);
and U5293 (N_5293,N_2557,N_3759);
nand U5294 (N_5294,N_2650,N_4209);
nor U5295 (N_5295,N_4123,N_3846);
nand U5296 (N_5296,N_2674,N_3385);
and U5297 (N_5297,N_2602,N_2665);
nand U5298 (N_5298,N_3974,N_4300);
and U5299 (N_5299,N_3829,N_3305);
and U5300 (N_5300,N_3050,N_2817);
xnor U5301 (N_5301,N_3872,N_2554);
xor U5302 (N_5302,N_3540,N_2609);
and U5303 (N_5303,N_4079,N_2757);
nor U5304 (N_5304,N_4446,N_3611);
nand U5305 (N_5305,N_4531,N_3520);
nor U5306 (N_5306,N_4255,N_3988);
xnor U5307 (N_5307,N_3990,N_3150);
or U5308 (N_5308,N_3547,N_2627);
nand U5309 (N_5309,N_4800,N_4422);
nor U5310 (N_5310,N_3284,N_4492);
or U5311 (N_5311,N_4675,N_4004);
nand U5312 (N_5312,N_3405,N_4222);
nor U5313 (N_5313,N_2835,N_3815);
and U5314 (N_5314,N_2651,N_4656);
and U5315 (N_5315,N_3416,N_4578);
nor U5316 (N_5316,N_3022,N_4689);
and U5317 (N_5317,N_3187,N_4618);
nand U5318 (N_5318,N_3959,N_3004);
or U5319 (N_5319,N_3193,N_3697);
or U5320 (N_5320,N_3992,N_4398);
nand U5321 (N_5321,N_2870,N_2623);
xor U5322 (N_5322,N_4751,N_4182);
or U5323 (N_5323,N_3072,N_3655);
and U5324 (N_5324,N_4257,N_3819);
nor U5325 (N_5325,N_2692,N_4729);
xor U5326 (N_5326,N_3732,N_3354);
nor U5327 (N_5327,N_3485,N_3334);
nor U5328 (N_5328,N_3902,N_2961);
nand U5329 (N_5329,N_2539,N_3430);
nor U5330 (N_5330,N_2850,N_2830);
or U5331 (N_5331,N_4853,N_4672);
nor U5332 (N_5332,N_3603,N_3041);
xnor U5333 (N_5333,N_2801,N_4518);
nor U5334 (N_5334,N_3300,N_3293);
nand U5335 (N_5335,N_3295,N_2567);
or U5336 (N_5336,N_4096,N_3919);
and U5337 (N_5337,N_2880,N_4693);
nand U5338 (N_5338,N_4192,N_4393);
and U5339 (N_5339,N_4013,N_4949);
and U5340 (N_5340,N_3771,N_4776);
nor U5341 (N_5341,N_2709,N_4259);
or U5342 (N_5342,N_2928,N_2679);
or U5343 (N_5343,N_3937,N_3555);
and U5344 (N_5344,N_3174,N_3920);
and U5345 (N_5345,N_4360,N_4854);
or U5346 (N_5346,N_4564,N_4350);
and U5347 (N_5347,N_2752,N_4107);
nor U5348 (N_5348,N_4576,N_3517);
nand U5349 (N_5349,N_2866,N_3380);
nand U5350 (N_5350,N_3475,N_3451);
nor U5351 (N_5351,N_4647,N_3876);
nor U5352 (N_5352,N_3103,N_4455);
xor U5353 (N_5353,N_3038,N_2758);
and U5354 (N_5354,N_3171,N_4077);
nor U5355 (N_5355,N_4373,N_3143);
nand U5356 (N_5356,N_3093,N_3666);
nand U5357 (N_5357,N_2582,N_2578);
and U5358 (N_5358,N_4582,N_3785);
and U5359 (N_5359,N_3608,N_2977);
nor U5360 (N_5360,N_4620,N_2610);
or U5361 (N_5361,N_4669,N_3672);
nand U5362 (N_5362,N_3332,N_3899);
xor U5363 (N_5363,N_4272,N_4317);
nor U5364 (N_5364,N_3470,N_3226);
nor U5365 (N_5365,N_3181,N_4205);
and U5366 (N_5366,N_3259,N_4007);
nor U5367 (N_5367,N_4438,N_3061);
nor U5368 (N_5368,N_4002,N_4613);
xor U5369 (N_5369,N_4911,N_3170);
xor U5370 (N_5370,N_2860,N_3348);
xnor U5371 (N_5371,N_3246,N_2922);
and U5372 (N_5372,N_3825,N_3970);
nor U5373 (N_5373,N_3831,N_2907);
and U5374 (N_5374,N_2857,N_3836);
or U5375 (N_5375,N_4817,N_3015);
or U5376 (N_5376,N_4838,N_4787);
xnor U5377 (N_5377,N_2950,N_4627);
xor U5378 (N_5378,N_3760,N_2951);
and U5379 (N_5379,N_4510,N_4186);
nor U5380 (N_5380,N_3756,N_3816);
nor U5381 (N_5381,N_3257,N_3465);
or U5382 (N_5382,N_4980,N_2882);
nor U5383 (N_5383,N_4149,N_4409);
nor U5384 (N_5384,N_2945,N_4985);
and U5385 (N_5385,N_4379,N_3971);
nand U5386 (N_5386,N_4181,N_2645);
and U5387 (N_5387,N_4551,N_3803);
xor U5388 (N_5388,N_4173,N_4737);
nor U5389 (N_5389,N_4567,N_4919);
xor U5390 (N_5390,N_4900,N_3708);
and U5391 (N_5391,N_3391,N_3117);
nand U5392 (N_5392,N_3593,N_4873);
nor U5393 (N_5393,N_4722,N_3127);
and U5394 (N_5394,N_3184,N_3091);
and U5395 (N_5395,N_3081,N_2601);
nand U5396 (N_5396,N_4468,N_2974);
nand U5397 (N_5397,N_2791,N_4767);
and U5398 (N_5398,N_4138,N_4608);
nand U5399 (N_5399,N_3747,N_3594);
and U5400 (N_5400,N_2994,N_4783);
nor U5401 (N_5401,N_4905,N_4947);
xnor U5402 (N_5402,N_4969,N_3030);
xor U5403 (N_5403,N_3524,N_3323);
nand U5404 (N_5404,N_3404,N_4391);
xnor U5405 (N_5405,N_4717,N_4712);
nand U5406 (N_5406,N_3455,N_4394);
or U5407 (N_5407,N_4329,N_2671);
or U5408 (N_5408,N_2747,N_4299);
xor U5409 (N_5409,N_3615,N_2502);
nand U5410 (N_5410,N_3886,N_4984);
or U5411 (N_5411,N_3249,N_2537);
xnor U5412 (N_5412,N_3076,N_2508);
xnor U5413 (N_5413,N_4844,N_4258);
and U5414 (N_5414,N_4872,N_3146);
nor U5415 (N_5415,N_4108,N_4981);
xnor U5416 (N_5416,N_3256,N_3607);
nand U5417 (N_5417,N_3023,N_2827);
and U5418 (N_5418,N_4032,N_3994);
nand U5419 (N_5419,N_4254,N_3487);
xnor U5420 (N_5420,N_3583,N_4653);
xor U5421 (N_5421,N_4676,N_3976);
and U5422 (N_5422,N_2905,N_3789);
nand U5423 (N_5423,N_4099,N_3653);
or U5424 (N_5424,N_3400,N_4831);
or U5425 (N_5425,N_3367,N_4027);
xnor U5426 (N_5426,N_4433,N_3479);
nor U5427 (N_5427,N_4429,N_3251);
and U5428 (N_5428,N_3357,N_2735);
and U5429 (N_5429,N_4494,N_3692);
xnor U5430 (N_5430,N_4701,N_3794);
nor U5431 (N_5431,N_2682,N_3518);
and U5432 (N_5432,N_4015,N_2936);
and U5433 (N_5433,N_2954,N_2980);
and U5434 (N_5434,N_4133,N_3036);
or U5435 (N_5435,N_3201,N_4999);
or U5436 (N_5436,N_4789,N_3136);
xor U5437 (N_5437,N_3702,N_3052);
and U5438 (N_5438,N_4474,N_3528);
nor U5439 (N_5439,N_4271,N_2673);
nand U5440 (N_5440,N_2748,N_4530);
or U5441 (N_5441,N_2685,N_4210);
xor U5442 (N_5442,N_4081,N_3343);
nand U5443 (N_5443,N_3039,N_2631);
nand U5444 (N_5444,N_4277,N_3134);
nor U5445 (N_5445,N_3527,N_2657);
nor U5446 (N_5446,N_3779,N_4063);
nor U5447 (N_5447,N_3308,N_3873);
xnor U5448 (N_5448,N_2815,N_4668);
nand U5449 (N_5449,N_4026,N_4581);
nor U5450 (N_5450,N_3606,N_4912);
or U5451 (N_5451,N_4803,N_3713);
and U5452 (N_5452,N_3932,N_2636);
nor U5453 (N_5453,N_4858,N_3715);
nand U5454 (N_5454,N_3933,N_3821);
nand U5455 (N_5455,N_3325,N_2616);
xor U5456 (N_5456,N_4112,N_4521);
or U5457 (N_5457,N_4679,N_2822);
xnor U5458 (N_5458,N_3590,N_3665);
and U5459 (N_5459,N_2511,N_4837);
nor U5460 (N_5460,N_4629,N_4539);
nand U5461 (N_5461,N_2971,N_4573);
xor U5462 (N_5462,N_2948,N_4579);
or U5463 (N_5463,N_3972,N_3240);
xor U5464 (N_5464,N_3297,N_4809);
nor U5465 (N_5465,N_3035,N_2596);
xnor U5466 (N_5466,N_3237,N_4631);
xnor U5467 (N_5467,N_2910,N_3306);
nand U5468 (N_5468,N_4535,N_2924);
and U5469 (N_5469,N_2978,N_2908);
nand U5470 (N_5470,N_3185,N_4920);
nand U5471 (N_5471,N_3307,N_4344);
nand U5472 (N_5472,N_2923,N_2612);
xor U5473 (N_5473,N_4707,N_4003);
xnor U5474 (N_5474,N_4268,N_3750);
xor U5475 (N_5475,N_4456,N_3945);
or U5476 (N_5476,N_2522,N_4348);
nor U5477 (N_5477,N_3281,N_2644);
nor U5478 (N_5478,N_3417,N_2591);
nor U5479 (N_5479,N_3654,N_4875);
xor U5480 (N_5480,N_4172,N_4059);
xor U5481 (N_5481,N_4216,N_3951);
nand U5482 (N_5482,N_4660,N_2969);
nor U5483 (N_5483,N_3273,N_4496);
nand U5484 (N_5484,N_4150,N_4775);
nand U5485 (N_5485,N_3676,N_3884);
and U5486 (N_5486,N_4655,N_3673);
and U5487 (N_5487,N_4824,N_4118);
or U5488 (N_5488,N_4749,N_4279);
and U5489 (N_5489,N_4610,N_3425);
nand U5490 (N_5490,N_4276,N_4166);
nand U5491 (N_5491,N_4085,N_3027);
nand U5492 (N_5492,N_2992,N_4607);
nor U5493 (N_5493,N_3253,N_2504);
nor U5494 (N_5494,N_2584,N_3817);
xor U5495 (N_5495,N_2571,N_3228);
nor U5496 (N_5496,N_2654,N_2788);
xor U5497 (N_5497,N_2999,N_4418);
xor U5498 (N_5498,N_3894,N_3602);
or U5499 (N_5499,N_4524,N_4136);
and U5500 (N_5500,N_2838,N_4990);
nor U5501 (N_5501,N_2766,N_4037);
xnor U5502 (N_5502,N_2962,N_3213);
and U5503 (N_5503,N_4076,N_2622);
nor U5504 (N_5504,N_4284,N_4559);
and U5505 (N_5505,N_3694,N_4370);
nand U5506 (N_5506,N_3133,N_2867);
nand U5507 (N_5507,N_4333,N_4857);
nand U5508 (N_5508,N_3717,N_2693);
and U5509 (N_5509,N_4874,N_4600);
or U5510 (N_5510,N_4713,N_3285);
and U5511 (N_5511,N_3667,N_2812);
nand U5512 (N_5512,N_4811,N_4061);
and U5513 (N_5513,N_3675,N_3445);
nand U5514 (N_5514,N_4241,N_2751);
xor U5515 (N_5515,N_4369,N_3296);
or U5516 (N_5516,N_3935,N_4477);
or U5517 (N_5517,N_2698,N_4151);
and U5518 (N_5518,N_4645,N_3044);
nand U5519 (N_5519,N_3936,N_4322);
or U5520 (N_5520,N_3340,N_3413);
nor U5521 (N_5521,N_4198,N_3239);
xnor U5522 (N_5522,N_2687,N_2749);
nor U5523 (N_5523,N_2542,N_3059);
xor U5524 (N_5524,N_3392,N_4532);
xor U5525 (N_5525,N_3543,N_3619);
or U5526 (N_5526,N_4315,N_2594);
and U5527 (N_5527,N_4017,N_3344);
nor U5528 (N_5528,N_4554,N_2935);
nor U5529 (N_5529,N_3459,N_3355);
nor U5530 (N_5530,N_3806,N_3761);
or U5531 (N_5531,N_4606,N_2818);
and U5532 (N_5532,N_3861,N_4421);
nand U5533 (N_5533,N_4586,N_4736);
nor U5534 (N_5534,N_3149,N_3778);
nand U5535 (N_5535,N_2753,N_3839);
nor U5536 (N_5536,N_2518,N_3108);
nand U5537 (N_5537,N_2932,N_3944);
nand U5538 (N_5538,N_2691,N_3458);
and U5539 (N_5539,N_4445,N_3985);
and U5540 (N_5540,N_3748,N_4867);
nand U5541 (N_5541,N_4080,N_4938);
nand U5542 (N_5542,N_3693,N_3048);
nor U5543 (N_5543,N_3066,N_3683);
xor U5544 (N_5544,N_4541,N_3471);
nor U5545 (N_5545,N_4461,N_2669);
nor U5546 (N_5546,N_4335,N_3166);
nand U5547 (N_5547,N_3729,N_4806);
nand U5548 (N_5548,N_4795,N_4955);
nor U5549 (N_5549,N_3464,N_3560);
or U5550 (N_5550,N_2750,N_3800);
xor U5551 (N_5551,N_4545,N_4991);
xnor U5552 (N_5552,N_3073,N_4120);
nor U5553 (N_5553,N_3467,N_4232);
nand U5554 (N_5554,N_2681,N_4522);
xor U5555 (N_5555,N_2976,N_3212);
and U5556 (N_5556,N_4711,N_4066);
nand U5557 (N_5557,N_3082,N_4566);
xnor U5558 (N_5558,N_3115,N_3671);
or U5559 (N_5559,N_4773,N_3565);
nand U5560 (N_5560,N_3278,N_4028);
nand U5561 (N_5561,N_4745,N_3997);
nor U5562 (N_5562,N_4604,N_4879);
nor U5563 (N_5563,N_4043,N_3832);
nor U5564 (N_5564,N_3599,N_2800);
and U5565 (N_5565,N_3087,N_3005);
or U5566 (N_5566,N_3659,N_3882);
or U5567 (N_5567,N_3842,N_4382);
and U5568 (N_5568,N_2842,N_2605);
nor U5569 (N_5569,N_3040,N_3709);
nor U5570 (N_5570,N_3034,N_4830);
xnor U5571 (N_5571,N_3339,N_2514);
nand U5572 (N_5572,N_3494,N_4320);
nor U5573 (N_5573,N_2878,N_4847);
or U5574 (N_5574,N_3682,N_2816);
or U5575 (N_5575,N_3769,N_2829);
nand U5576 (N_5576,N_3907,N_3774);
and U5577 (N_5577,N_4978,N_3469);
xor U5578 (N_5578,N_3018,N_4122);
nor U5579 (N_5579,N_4458,N_2806);
or U5580 (N_5580,N_4763,N_3582);
nand U5581 (N_5581,N_3773,N_2595);
nand U5582 (N_5582,N_3969,N_4194);
nand U5583 (N_5583,N_4820,N_2965);
and U5584 (N_5584,N_3544,N_2639);
xnor U5585 (N_5585,N_2733,N_3840);
nand U5586 (N_5586,N_4880,N_2585);
nor U5587 (N_5587,N_2990,N_4798);
or U5588 (N_5588,N_4744,N_2987);
or U5589 (N_5589,N_2580,N_2550);
and U5590 (N_5590,N_4726,N_4917);
nand U5591 (N_5591,N_3956,N_4359);
nand U5592 (N_5592,N_3609,N_2739);
or U5593 (N_5593,N_3365,N_4519);
nand U5594 (N_5594,N_3763,N_3379);
or U5595 (N_5595,N_4167,N_3918);
and U5596 (N_5596,N_4500,N_4808);
nor U5597 (N_5597,N_3025,N_4036);
nand U5598 (N_5598,N_3489,N_3424);
and U5599 (N_5599,N_3787,N_4134);
nand U5600 (N_5600,N_2500,N_4860);
xor U5601 (N_5601,N_4762,N_2756);
and U5602 (N_5602,N_4654,N_2942);
or U5603 (N_5603,N_3074,N_4463);
or U5604 (N_5604,N_4547,N_3757);
nand U5605 (N_5605,N_4452,N_4735);
and U5606 (N_5606,N_3798,N_3903);
or U5607 (N_5607,N_2614,N_3126);
nor U5608 (N_5608,N_2769,N_4062);
or U5609 (N_5609,N_3991,N_4064);
nor U5610 (N_5610,N_4312,N_4472);
nor U5611 (N_5611,N_3818,N_2598);
xor U5612 (N_5612,N_3772,N_3576);
nor U5613 (N_5613,N_4239,N_3157);
and U5614 (N_5614,N_4979,N_4234);
xor U5615 (N_5615,N_2904,N_3432);
xnor U5616 (N_5616,N_3690,N_2549);
or U5617 (N_5617,N_3862,N_3501);
nor U5618 (N_5618,N_2934,N_4056);
and U5619 (N_5619,N_3914,N_4842);
xor U5620 (N_5620,N_3065,N_3604);
xnor U5621 (N_5621,N_2765,N_2834);
nor U5622 (N_5622,N_2985,N_3963);
xnor U5623 (N_5623,N_4624,N_4501);
nor U5624 (N_5624,N_3640,N_4091);
or U5625 (N_5625,N_3320,N_3026);
nand U5626 (N_5626,N_4750,N_3277);
and U5627 (N_5627,N_3114,N_3567);
or U5628 (N_5628,N_4154,N_4870);
nand U5629 (N_5629,N_4296,N_3363);
xor U5630 (N_5630,N_3217,N_4218);
and U5631 (N_5631,N_4727,N_2940);
or U5632 (N_5632,N_4211,N_4265);
nor U5633 (N_5633,N_3904,N_2909);
xor U5634 (N_5634,N_3442,N_3851);
nand U5635 (N_5635,N_3209,N_4327);
xnor U5636 (N_5636,N_3984,N_3766);
or U5637 (N_5637,N_3656,N_3558);
and U5638 (N_5638,N_3097,N_3651);
and U5639 (N_5639,N_3316,N_3681);
and U5640 (N_5640,N_3849,N_3234);
and U5641 (N_5641,N_3423,N_3169);
or U5642 (N_5642,N_3499,N_3575);
nor U5643 (N_5643,N_4071,N_3939);
nand U5644 (N_5644,N_4478,N_3014);
nand U5645 (N_5645,N_4952,N_4714);
and U5646 (N_5646,N_4240,N_3584);
nand U5647 (N_5647,N_4742,N_2649);
xnor U5648 (N_5648,N_3067,N_3621);
nor U5649 (N_5649,N_3768,N_4340);
nor U5650 (N_5650,N_4397,N_4052);
or U5651 (N_5651,N_4068,N_4771);
nand U5652 (N_5652,N_4596,N_3887);
nand U5653 (N_5653,N_4164,N_4100);
or U5654 (N_5654,N_3195,N_2697);
xor U5655 (N_5655,N_3924,N_4489);
xor U5656 (N_5656,N_3346,N_2970);
xnor U5657 (N_5657,N_4643,N_4336);
and U5658 (N_5658,N_3260,N_2988);
nand U5659 (N_5659,N_2558,N_3674);
nor U5660 (N_5660,N_3192,N_4637);
nor U5661 (N_5661,N_2648,N_3173);
xnor U5662 (N_5662,N_2521,N_3738);
nor U5663 (N_5663,N_3811,N_3418);
xnor U5664 (N_5664,N_3827,N_4000);
xor U5665 (N_5665,N_3506,N_2613);
or U5666 (N_5666,N_3198,N_4796);
nor U5667 (N_5667,N_3177,N_4498);
nor U5668 (N_5668,N_3895,N_4384);
nor U5669 (N_5669,N_4253,N_3085);
and U5670 (N_5670,N_2858,N_4797);
xnor U5671 (N_5671,N_3896,N_4930);
or U5672 (N_5672,N_4499,N_3523);
and U5673 (N_5673,N_4413,N_3637);
nor U5674 (N_5674,N_3370,N_3744);
and U5675 (N_5675,N_4290,N_4670);
and U5676 (N_5676,N_3531,N_2819);
nor U5677 (N_5677,N_3145,N_4544);
or U5678 (N_5678,N_3783,N_2740);
nand U5679 (N_5679,N_3124,N_3223);
xnor U5680 (N_5680,N_3507,N_4652);
xnor U5681 (N_5681,N_4558,N_4534);
or U5682 (N_5682,N_2913,N_4280);
xnor U5683 (N_5683,N_3456,N_3268);
xnor U5684 (N_5684,N_4408,N_2868);
xnor U5685 (N_5685,N_2798,N_3452);
or U5686 (N_5686,N_3299,N_4411);
nand U5687 (N_5687,N_3964,N_3740);
nor U5688 (N_5688,N_3541,N_3734);
xnor U5689 (N_5689,N_3020,N_3841);
nor U5690 (N_5690,N_3183,N_4473);
and U5691 (N_5691,N_3472,N_4148);
and U5692 (N_5692,N_3182,N_4960);
or U5693 (N_5693,N_4016,N_4704);
xnor U5694 (N_5694,N_4908,N_3813);
or U5695 (N_5695,N_2849,N_3801);
nand U5696 (N_5696,N_2738,N_4155);
xnor U5697 (N_5697,N_3488,N_2520);
xnor U5698 (N_5698,N_2888,N_4295);
or U5699 (N_5699,N_3514,N_4517);
nand U5700 (N_5700,N_4286,N_4323);
or U5701 (N_5701,N_3197,N_4869);
xnor U5702 (N_5702,N_2780,N_3533);
or U5703 (N_5703,N_4665,N_3691);
or U5704 (N_5704,N_3180,N_4513);
nand U5705 (N_5705,N_4683,N_3409);
and U5706 (N_5706,N_3319,N_4140);
nand U5707 (N_5707,N_4025,N_3500);
or U5708 (N_5708,N_4570,N_4995);
nand U5709 (N_5709,N_3099,N_2695);
nand U5710 (N_5710,N_3795,N_4487);
and U5711 (N_5711,N_2618,N_3577);
xnor U5712 (N_5712,N_2577,N_3758);
and U5713 (N_5713,N_2861,N_4128);
nor U5714 (N_5714,N_3387,N_3915);
nor U5715 (N_5715,N_4363,N_3341);
nand U5716 (N_5716,N_4959,N_4306);
and U5717 (N_5717,N_3436,N_4584);
and U5718 (N_5718,N_4520,N_4633);
nand U5719 (N_5719,N_3283,N_4939);
and U5720 (N_5720,N_3552,N_2871);
xnor U5721 (N_5721,N_3954,N_3468);
xnor U5722 (N_5722,N_3934,N_2525);
nor U5723 (N_5723,N_3003,N_4177);
xnor U5724 (N_5724,N_2804,N_3865);
nor U5725 (N_5725,N_3158,N_4381);
xnor U5726 (N_5726,N_4111,N_2628);
nand U5727 (N_5727,N_4260,N_4078);
nand U5728 (N_5728,N_3598,N_4987);
nor U5729 (N_5729,N_4038,N_2813);
xor U5730 (N_5730,N_3002,N_2767);
nand U5731 (N_5731,N_4725,N_3550);
and U5732 (N_5732,N_4684,N_4127);
nor U5733 (N_5733,N_4845,N_3643);
nor U5734 (N_5734,N_3190,N_3854);
or U5735 (N_5735,N_3537,N_4441);
or U5736 (N_5736,N_2760,N_3810);
xnor U5737 (N_5737,N_4590,N_3314);
or U5738 (N_5738,N_2754,N_4859);
nor U5739 (N_5739,N_2865,N_4791);
nor U5740 (N_5740,N_3885,N_2579);
or U5741 (N_5741,N_4124,N_4311);
xor U5742 (N_5742,N_3433,N_3414);
nor U5743 (N_5743,N_4922,N_3110);
nand U5744 (N_5744,N_3204,N_2683);
nor U5745 (N_5745,N_3941,N_3294);
and U5746 (N_5746,N_2807,N_2731);
nand U5747 (N_5747,N_4815,N_3652);
nand U5748 (N_5748,N_2737,N_3796);
nand U5749 (N_5749,N_4591,N_4885);
nor U5750 (N_5750,N_3481,N_4215);
or U5751 (N_5751,N_3687,N_4217);
nor U5752 (N_5752,N_4308,N_3156);
nand U5753 (N_5753,N_2956,N_4420);
and U5754 (N_5754,N_3561,N_2734);
and U5755 (N_5755,N_4728,N_4436);
nor U5756 (N_5756,N_4130,N_3596);
and U5757 (N_5757,N_4924,N_3626);
or U5758 (N_5758,N_3618,N_3511);
or U5759 (N_5759,N_3830,N_4464);
or U5760 (N_5760,N_2937,N_2828);
or U5761 (N_5761,N_3616,N_4515);
or U5762 (N_5762,N_4225,N_4833);
xor U5763 (N_5763,N_2551,N_4351);
or U5764 (N_5764,N_3311,N_3677);
xor U5765 (N_5765,N_2505,N_3266);
or U5766 (N_5766,N_4710,N_4734);
and U5767 (N_5767,N_4303,N_3595);
nand U5768 (N_5768,N_3101,N_4153);
xor U5769 (N_5769,N_4170,N_2872);
xnor U5770 (N_5770,N_3484,N_3402);
xor U5771 (N_5771,N_2704,N_2986);
or U5772 (N_5772,N_3298,N_3429);
nand U5773 (N_5773,N_4353,N_4696);
nor U5774 (N_5774,N_3309,N_4560);
or U5775 (N_5775,N_2795,N_3731);
or U5776 (N_5776,N_2744,N_3522);
nor U5777 (N_5777,N_2586,N_2535);
or U5778 (N_5778,N_4715,N_4886);
or U5779 (N_5779,N_4427,N_2686);
nor U5780 (N_5780,N_4219,N_4597);
and U5781 (N_5781,N_3265,N_4029);
nor U5782 (N_5782,N_3427,N_3880);
xnor U5783 (N_5783,N_4221,N_3610);
nand U5784 (N_5784,N_2728,N_4580);
nand U5785 (N_5785,N_4426,N_4325);
nor U5786 (N_5786,N_4419,N_4852);
xor U5787 (N_5787,N_4405,N_2703);
xnor U5788 (N_5788,N_4358,N_3165);
xor U5789 (N_5789,N_4401,N_3480);
xnor U5790 (N_5790,N_4213,N_4864);
nor U5791 (N_5791,N_3875,N_3345);
nor U5792 (N_5792,N_4162,N_3107);
and U5793 (N_5793,N_3554,N_4720);
xor U5794 (N_5794,N_3710,N_4848);
nor U5795 (N_5795,N_4207,N_4288);
xnor U5796 (N_5796,N_3850,N_3454);
or U5797 (N_5797,N_3330,N_4493);
xnor U5798 (N_5798,N_4916,N_4287);
or U5799 (N_5799,N_2778,N_3823);
nand U5800 (N_5800,N_3966,N_2927);
or U5801 (N_5801,N_3981,N_3461);
nand U5802 (N_5802,N_2689,N_3408);
nand U5803 (N_5803,N_3244,N_3168);
nor U5804 (N_5804,N_2592,N_2660);
xnor U5805 (N_5805,N_3853,N_4662);
xnor U5806 (N_5806,N_4671,N_4741);
nand U5807 (N_5807,N_4996,N_4200);
nand U5808 (N_5808,N_3312,N_4145);
nor U5809 (N_5809,N_4819,N_3628);
nor U5810 (N_5810,N_3086,N_3047);
xnor U5811 (N_5811,N_3496,N_4975);
or U5812 (N_5812,N_4964,N_4644);
nand U5813 (N_5813,N_2914,N_3216);
or U5814 (N_5814,N_4406,N_3721);
nand U5815 (N_5815,N_2573,N_2675);
or U5816 (N_5816,N_4332,N_4119);
and U5817 (N_5817,N_2845,N_3440);
nand U5818 (N_5818,N_2946,N_4289);
and U5819 (N_5819,N_3680,N_3877);
nor U5820 (N_5820,N_4687,N_3508);
nand U5821 (N_5821,N_3620,N_4022);
nand U5822 (N_5822,N_4951,N_3644);
xor U5823 (N_5823,N_3509,N_3696);
xor U5824 (N_5824,N_4443,N_2513);
xnor U5825 (N_5825,N_3245,N_4846);
or U5826 (N_5826,N_4928,N_3647);
or U5827 (N_5827,N_4188,N_4184);
xor U5828 (N_5828,N_2543,N_4507);
xnor U5829 (N_5829,N_4799,N_4595);
or U5830 (N_5830,N_3196,N_4465);
nor U5831 (N_5831,N_2916,N_3090);
nor U5832 (N_5832,N_2824,N_2629);
or U5833 (N_5833,N_4863,N_2840);
nand U5834 (N_5834,N_4009,N_4049);
xor U5835 (N_5835,N_3350,N_4899);
xor U5836 (N_5836,N_4910,N_4199);
or U5837 (N_5837,N_3879,N_4865);
nor U5838 (N_5838,N_3371,N_3642);
xor U5839 (N_5839,N_3612,N_2997);
or U5840 (N_5840,N_3578,N_3684);
and U5841 (N_5841,N_4270,N_3701);
and U5842 (N_5842,N_3028,N_3967);
nor U5843 (N_5843,N_4183,N_3538);
and U5844 (N_5844,N_4161,N_2854);
or U5845 (N_5845,N_4060,N_4230);
nand U5846 (N_5846,N_4623,N_3352);
and U5847 (N_5847,N_4577,N_3222);
nand U5848 (N_5848,N_3328,N_2825);
or U5849 (N_5849,N_4462,N_3733);
nor U5850 (N_5850,N_4861,N_3855);
or U5851 (N_5851,N_2794,N_4482);
xor U5852 (N_5852,N_3711,N_3096);
or U5853 (N_5853,N_3743,N_2773);
or U5854 (N_5854,N_4485,N_4746);
nor U5855 (N_5855,N_2741,N_3749);
and U5856 (N_5856,N_3389,N_2633);
nand U5857 (N_5857,N_2957,N_4708);
and U5858 (N_5858,N_4208,N_2688);
nand U5859 (N_5859,N_4506,N_3724);
nand U5860 (N_5860,N_2587,N_4855);
xor U5861 (N_5861,N_4318,N_3635);
xor U5862 (N_5862,N_4993,N_2763);
and U5863 (N_5863,N_3474,N_2517);
xnor U5864 (N_5864,N_2619,N_4768);
nand U5865 (N_5865,N_3261,N_3699);
xor U5866 (N_5866,N_4638,N_3622);
or U5867 (N_5867,N_4480,N_4664);
nor U5868 (N_5868,N_3230,N_3767);
xor U5869 (N_5869,N_4309,N_2581);
nor U5870 (N_5870,N_3863,N_3977);
and U5871 (N_5871,N_4021,N_4505);
nand U5872 (N_5872,N_3926,N_4983);
or U5873 (N_5873,N_3663,N_4802);
nand U5874 (N_5874,N_4902,N_3075);
xnor U5875 (N_5875,N_2764,N_3569);
or U5876 (N_5876,N_2626,N_2710);
or U5877 (N_5877,N_2576,N_3782);
xnor U5878 (N_5878,N_4156,N_4357);
and U5879 (N_5879,N_2831,N_3563);
and U5880 (N_5880,N_4935,N_3356);
xor U5881 (N_5881,N_2783,N_4158);
nor U5882 (N_5882,N_3581,N_4828);
xnor U5883 (N_5883,N_4511,N_4471);
and U5884 (N_5884,N_3426,N_4466);
nand U5885 (N_5885,N_4723,N_3949);
or U5886 (N_5886,N_3069,N_4375);
nor U5887 (N_5887,N_2516,N_2903);
and U5888 (N_5888,N_3194,N_4818);
nor U5889 (N_5889,N_3780,N_4146);
and U5890 (N_5890,N_4934,N_3781);
nor U5891 (N_5891,N_3623,N_3351);
nand U5892 (N_5892,N_2705,N_4330);
nor U5893 (N_5893,N_3921,N_3381);
nand U5894 (N_5894,N_4550,N_3045);
and U5895 (N_5895,N_3505,N_2898);
xnor U5896 (N_5896,N_2852,N_3215);
nand U5897 (N_5897,N_4780,N_4926);
xor U5898 (N_5898,N_4945,N_2736);
nor U5899 (N_5899,N_2708,N_2732);
nand U5900 (N_5900,N_3119,N_3808);
nand U5901 (N_5901,N_2991,N_3591);
and U5902 (N_5902,N_3225,N_4758);
or U5903 (N_5903,N_3545,N_3130);
or U5904 (N_5904,N_3057,N_4706);
or U5905 (N_5905,N_4459,N_3916);
nand U5906 (N_5906,N_3987,N_4523);
xnor U5907 (N_5907,N_4884,N_3395);
xnor U5908 (N_5908,N_4747,N_3588);
nand U5909 (N_5909,N_4048,N_3457);
xnor U5910 (N_5910,N_3617,N_3006);
or U5911 (N_5911,N_4388,N_4943);
nand U5912 (N_5912,N_4448,N_4781);
xnor U5913 (N_5913,N_4389,N_3247);
or U5914 (N_5914,N_4479,N_4115);
nand U5915 (N_5915,N_4825,N_3847);
or U5916 (N_5916,N_3664,N_4944);
and U5917 (N_5917,N_3397,N_2876);
and U5918 (N_5918,N_3601,N_4269);
nor U5919 (N_5919,N_4233,N_4497);
xor U5920 (N_5920,N_2998,N_3998);
or U5921 (N_5921,N_3973,N_3055);
or U5922 (N_5922,N_4476,N_3079);
nor U5923 (N_5923,N_4814,N_4297);
nand U5924 (N_5924,N_2723,N_3398);
or U5925 (N_5925,N_3214,N_2607);
xnor U5926 (N_5926,N_3999,N_3614);
or U5927 (N_5927,N_4058,N_4228);
nand U5928 (N_5928,N_4457,N_4816);
nor U5929 (N_5929,N_3530,N_4223);
xnor U5930 (N_5930,N_2509,N_4538);
nand U5931 (N_5931,N_2820,N_3912);
xnor U5932 (N_5932,N_3889,N_3688);
or U5933 (N_5933,N_2874,N_3579);
nor U5934 (N_5934,N_3497,N_3007);
nor U5935 (N_5935,N_2716,N_3549);
or U5936 (N_5936,N_4226,N_2772);
nor U5937 (N_5937,N_2981,N_3176);
xnor U5938 (N_5938,N_4876,N_2670);
xnor U5939 (N_5939,N_4740,N_3167);
nor U5940 (N_5940,N_3046,N_3291);
and U5941 (N_5941,N_4065,N_4516);
nor U5942 (N_5942,N_2966,N_3638);
xnor U5943 (N_5943,N_3264,N_2726);
nor U5944 (N_5944,N_4793,N_3625);
xor U5945 (N_5945,N_4105,N_2570);
nand U5946 (N_5946,N_3534,N_4877);
xnor U5947 (N_5947,N_3233,N_2846);
or U5948 (N_5948,N_2859,N_4822);
nor U5949 (N_5949,N_4724,N_4354);
nand U5950 (N_5950,N_4097,N_3589);
and U5951 (N_5951,N_2702,N_4508);
nand U5952 (N_5952,N_4075,N_4103);
nor U5953 (N_5953,N_2779,N_3866);
and U5954 (N_5954,N_2784,N_4626);
nand U5955 (N_5955,N_3900,N_3648);
nand U5956 (N_5956,N_4012,N_2700);
nor U5957 (N_5957,N_3366,N_4982);
or U5958 (N_5958,N_3151,N_4434);
nand U5959 (N_5959,N_2615,N_3301);
and U5960 (N_5960,N_3327,N_3512);
nor U5961 (N_5961,N_4892,N_4881);
and U5962 (N_5962,N_4014,N_2684);
nand U5963 (N_5963,N_2921,N_4084);
xor U5964 (N_5964,N_4235,N_3728);
and U5965 (N_5965,N_4440,N_3384);
nor U5966 (N_5966,N_4702,N_4777);
nand U5967 (N_5967,N_4010,N_3083);
or U5968 (N_5968,N_2715,N_3751);
or U5969 (N_5969,N_3860,N_2699);
nand U5970 (N_5970,N_2847,N_3431);
xor U5971 (N_5971,N_4283,N_2559);
xnor U5972 (N_5972,N_3286,N_2540);
nand U5973 (N_5973,N_3722,N_3491);
xnor U5974 (N_5974,N_3613,N_3931);
nor U5975 (N_5975,N_2963,N_4423);
xor U5976 (N_5976,N_3258,N_3807);
or U5977 (N_5977,N_3600,N_4361);
and U5978 (N_5978,N_3353,N_4936);
or U5979 (N_5979,N_4907,N_2536);
and U5980 (N_5980,N_4589,N_3412);
nor U5981 (N_5981,N_4095,N_2564);
nor U5982 (N_5982,N_4526,N_4898);
or U5983 (N_5983,N_2892,N_3868);
or U5984 (N_5984,N_3962,N_3953);
nor U5985 (N_5985,N_4345,N_3928);
xnor U5986 (N_5986,N_4894,N_4109);
nand U5987 (N_5987,N_4697,N_3824);
xnor U5988 (N_5988,N_4033,N_3670);
nor U5989 (N_5989,N_4328,N_4273);
and U5990 (N_5990,N_3338,N_3446);
nand U5991 (N_5991,N_4163,N_2655);
xor U5992 (N_5992,N_3745,N_3267);
nand U5993 (N_5993,N_2526,N_2933);
nor U5994 (N_5994,N_3131,N_4681);
nor U5995 (N_5995,N_4346,N_4632);
or U5996 (N_5996,N_3753,N_2643);
xnor U5997 (N_5997,N_4691,N_4839);
nor U5998 (N_5998,N_3051,N_4090);
or U5999 (N_5999,N_3719,N_4031);
and U6000 (N_6000,N_4602,N_2572);
or U6001 (N_6001,N_3123,N_3450);
xnor U6002 (N_6002,N_3636,N_2701);
and U6003 (N_6003,N_4187,N_4143);
nand U6004 (N_6004,N_2727,N_3874);
nand U6005 (N_6005,N_2637,N_4088);
nand U6006 (N_6006,N_2746,N_2755);
or U6007 (N_6007,N_2718,N_4314);
and U6008 (N_6008,N_4575,N_4197);
and U6009 (N_6009,N_3980,N_4970);
or U6010 (N_6010,N_4475,N_4685);
or U6011 (N_6011,N_4019,N_3274);
nand U6012 (N_6012,N_2552,N_3105);
or U6013 (N_6013,N_4572,N_2519);
xor U6014 (N_6014,N_2590,N_2544);
and U6015 (N_6015,N_3444,N_3100);
xor U6016 (N_6016,N_2989,N_3490);
nand U6017 (N_6017,N_4868,N_3777);
and U6018 (N_6018,N_3383,N_4556);
or U6019 (N_6019,N_3390,N_4546);
nand U6020 (N_6020,N_4364,N_3420);
nand U6021 (N_6021,N_2621,N_2663);
nand U6022 (N_6022,N_4180,N_2583);
nand U6023 (N_6023,N_2593,N_4895);
or U6024 (N_6024,N_4294,N_3178);
nand U6025 (N_6025,N_4548,N_4901);
and U6026 (N_6026,N_3632,N_3513);
nand U6027 (N_6027,N_3407,N_4635);
xnor U6028 (N_6028,N_3098,N_3564);
nor U6029 (N_6029,N_3262,N_4555);
nand U6030 (N_6030,N_4965,N_3568);
or U6031 (N_6031,N_3515,N_4552);
xor U6032 (N_6032,N_2722,N_2711);
xor U6033 (N_6033,N_4821,N_4757);
xor U6034 (N_6034,N_3986,N_3053);
and U6035 (N_6035,N_2661,N_3478);
nand U6036 (N_6036,N_3566,N_4387);
and U6037 (N_6037,N_3292,N_4495);
or U6038 (N_6038,N_3476,N_4968);
xor U6039 (N_6039,N_3551,N_4650);
xnor U6040 (N_6040,N_3845,N_4196);
nor U6041 (N_6041,N_2694,N_4639);
nor U6042 (N_6042,N_2855,N_4542);
and U6043 (N_6043,N_3411,N_3172);
xnor U6044 (N_6044,N_4733,N_3448);
nand U6045 (N_6045,N_2893,N_4792);
xnor U6046 (N_6046,N_3592,N_4972);
or U6047 (N_6047,N_4054,N_4431);
or U6048 (N_6048,N_3678,N_3375);
or U6049 (N_6049,N_2712,N_2743);
xor U6050 (N_6050,N_3449,N_4407);
or U6051 (N_6051,N_4261,N_2877);
nand U6052 (N_6052,N_4176,N_3393);
or U6053 (N_6053,N_4703,N_4304);
nand U6054 (N_6054,N_2528,N_2826);
nor U6055 (N_6055,N_4680,N_2848);
xor U6056 (N_6056,N_3726,N_2677);
and U6057 (N_6057,N_4716,N_4008);
and U6058 (N_6058,N_3410,N_2821);
or U6059 (N_6059,N_2729,N_3844);
and U6060 (N_6060,N_3242,N_2563);
and U6061 (N_6061,N_3272,N_3752);
or U6062 (N_6062,N_4204,N_4267);
nor U6063 (N_6063,N_3483,N_4371);
nor U6064 (N_6064,N_4005,N_4721);
and U6065 (N_6065,N_4117,N_4754);
or U6066 (N_6066,N_4082,N_4615);
nor U6067 (N_6067,N_4829,N_3942);
nor U6068 (N_6068,N_4055,N_3089);
and U6069 (N_6069,N_2793,N_4374);
xnor U6070 (N_6070,N_2530,N_4470);
nand U6071 (N_6071,N_4070,N_3605);
or U6072 (N_6072,N_3859,N_3322);
nor U6073 (N_6073,N_4491,N_3668);
nor U6074 (N_6074,N_2979,N_3968);
nor U6075 (N_6075,N_3843,N_4089);
or U6076 (N_6076,N_4986,N_3776);
xor U6077 (N_6077,N_4921,N_4262);
and U6078 (N_6078,N_3858,N_3993);
and U6079 (N_6079,N_3270,N_2958);
xnor U6080 (N_6080,N_4925,N_4961);
nor U6081 (N_6081,N_4451,N_2611);
and U6082 (N_6082,N_3280,N_4648);
xnor U6083 (N_6083,N_3362,N_4385);
nand U6084 (N_6084,N_3791,N_2984);
xnor U6085 (N_6085,N_4856,N_2931);
nand U6086 (N_6086,N_4113,N_4784);
nand U6087 (N_6087,N_3657,N_4326);
nand U6088 (N_6088,N_2918,N_3704);
nor U6089 (N_6089,N_4766,N_4292);
and U6090 (N_6090,N_4404,N_3943);
nand U6091 (N_6091,N_2566,N_2515);
nor U6092 (N_6092,N_2768,N_4483);
xnor U6093 (N_6093,N_3996,N_3271);
or U6094 (N_6094,N_3765,N_3062);
nand U6095 (N_6095,N_4447,N_2930);
or U6096 (N_6096,N_3317,N_3140);
or U6097 (N_6097,N_3388,N_3011);
nor U6098 (N_6098,N_3707,N_3770);
or U6099 (N_6099,N_3331,N_4356);
and U6100 (N_6100,N_2993,N_3901);
nor U6101 (N_6101,N_2911,N_2952);
xnor U6102 (N_6102,N_2881,N_4659);
xnor U6103 (N_6103,N_3024,N_2836);
nor U6104 (N_6104,N_4882,N_4110);
or U6105 (N_6105,N_3909,N_3822);
nor U6106 (N_6106,N_3746,N_2814);
or U6107 (N_6107,N_4366,N_2730);
nor U6108 (N_6108,N_4453,N_3419);
xnor U6109 (N_6109,N_3546,N_4764);
nor U6110 (N_6110,N_3950,N_3032);
and U6111 (N_6111,N_2538,N_4849);
and U6112 (N_6112,N_3252,N_3241);
or U6113 (N_6113,N_2975,N_3833);
or U6114 (N_6114,N_3263,N_3058);
xor U6115 (N_6115,N_3042,N_4274);
nand U6116 (N_6116,N_3118,N_4231);
or U6117 (N_6117,N_4962,N_2672);
nand U6118 (N_6118,N_2853,N_4201);
or U6119 (N_6119,N_3630,N_2575);
xor U6120 (N_6120,N_4291,N_2547);
xnor U6121 (N_6121,N_4903,N_3088);
xor U6122 (N_6122,N_2843,N_3525);
nand U6123 (N_6123,N_3870,N_2604);
xnor U6124 (N_6124,N_4424,N_4185);
or U6125 (N_6125,N_4488,N_3723);
nor U6126 (N_6126,N_3112,N_3153);
and U6127 (N_6127,N_3927,N_3730);
nand U6128 (N_6128,N_4823,N_3010);
or U6129 (N_6129,N_2917,N_2568);
xor U6130 (N_6130,N_4927,N_4244);
nor U6131 (N_6131,N_3556,N_2912);
and U6132 (N_6132,N_3957,N_3881);
nand U6133 (N_6133,N_4810,N_3435);
and U6134 (N_6134,N_4688,N_3358);
nand U6135 (N_6135,N_3238,N_4966);
nor U6136 (N_6136,N_2902,N_3571);
and U6137 (N_6137,N_4619,N_3790);
nor U6138 (N_6138,N_3012,N_4252);
and U6139 (N_6139,N_4997,N_3526);
or U6140 (N_6140,N_2811,N_2782);
xor U6141 (N_6141,N_4621,N_4732);
xor U6142 (N_6142,N_3947,N_4977);
nand U6143 (N_6143,N_2656,N_3373);
and U6144 (N_6144,N_3802,N_4417);
nand U6145 (N_6145,N_4692,N_2896);
and U6146 (N_6146,N_3129,N_4193);
or U6147 (N_6147,N_2562,N_2883);
nor U6148 (N_6148,N_4569,N_3580);
nand U6149 (N_6149,N_4514,N_4851);
and U6150 (N_6150,N_3989,N_2668);
xnor U6151 (N_6151,N_3186,N_3764);
nor U6152 (N_6152,N_3809,N_4553);
nor U6153 (N_6153,N_3826,N_3553);
or U6154 (N_6154,N_4045,N_2953);
xor U6155 (N_6155,N_4490,N_2983);
nor U6156 (N_6156,N_2943,N_2588);
xor U6157 (N_6157,N_4018,N_3686);
or U6158 (N_6158,N_2941,N_4807);
or U6159 (N_6159,N_3236,N_2634);
nor U6160 (N_6160,N_3056,N_2823);
and U6161 (N_6161,N_3498,N_4942);
and U6162 (N_6162,N_3775,N_2762);
or U6163 (N_6163,N_3164,N_3466);
and U6164 (N_6164,N_3572,N_3961);
xor U6165 (N_6165,N_3160,N_3189);
nand U6166 (N_6166,N_4913,N_2642);
and U6167 (N_6167,N_3705,N_3276);
nand U6168 (N_6168,N_3883,N_3349);
and U6169 (N_6169,N_4467,N_3742);
nand U6170 (N_6170,N_2531,N_2833);
nand U6171 (N_6171,N_4141,N_4906);
or U6172 (N_6172,N_4904,N_2920);
nor U6173 (N_6173,N_3799,N_4191);
or U6174 (N_6174,N_3960,N_3834);
and U6175 (N_6175,N_4313,N_3104);
xor U6176 (N_6176,N_4030,N_3324);
or U6177 (N_6177,N_2786,N_4316);
and U6178 (N_6178,N_2658,N_3837);
and U6179 (N_6179,N_3106,N_4948);
and U6180 (N_6180,N_3179,N_3248);
or U6181 (N_6181,N_2890,N_2929);
and U6182 (N_6182,N_3735,N_3394);
xor U6183 (N_6183,N_2532,N_2805);
nor U6184 (N_6184,N_4923,N_4129);
or U6185 (N_6185,N_3460,N_3573);
nor U6186 (N_6186,N_2781,N_3326);
and U6187 (N_6187,N_3535,N_3064);
nand U6188 (N_6188,N_2915,N_4342);
xnor U6189 (N_6189,N_4958,N_3382);
xnor U6190 (N_6190,N_4663,N_4739);
nor U6191 (N_6191,N_3646,N_3736);
xnor U6192 (N_6192,N_4237,N_3208);
or U6193 (N_6193,N_3043,N_3586);
nand U6194 (N_6194,N_4147,N_3376);
nand U6195 (N_6195,N_4251,N_3975);
nand U6196 (N_6196,N_4954,N_2706);
nand U6197 (N_6197,N_3958,N_3814);
xor U6198 (N_6198,N_4897,N_4695);
and U6199 (N_6199,N_4399,N_2887);
nand U6200 (N_6200,N_3071,N_2574);
and U6201 (N_6201,N_4386,N_4046);
nand U6202 (N_6202,N_4245,N_4525);
nor U6203 (N_6203,N_4658,N_4106);
or U6204 (N_6204,N_3031,N_3321);
nand U6205 (N_6205,N_4390,N_4549);
nand U6206 (N_6206,N_4587,N_4093);
nand U6207 (N_6207,N_4135,N_2597);
nand U6208 (N_6208,N_3080,N_3224);
xor U6209 (N_6209,N_4227,N_3219);
nand U6210 (N_6210,N_3109,N_4612);
and U6211 (N_6211,N_2884,N_4603);
nor U6212 (N_6212,N_4416,N_3154);
and U6213 (N_6213,N_4871,N_3335);
xnor U6214 (N_6214,N_2641,N_3718);
and U6215 (N_6215,N_4247,N_4769);
xor U6216 (N_6216,N_4957,N_4083);
and U6217 (N_6217,N_4738,N_3369);
nand U6218 (N_6218,N_3202,N_4752);
nor U6219 (N_6219,N_3835,N_4705);
nand U6220 (N_6220,N_4804,N_3797);
xnor U6221 (N_6221,N_4460,N_4224);
nor U6222 (N_6222,N_3486,N_2632);
xnor U6223 (N_6223,N_4976,N_2837);
nor U6224 (N_6224,N_2939,N_4432);
and U6225 (N_6225,N_4649,N_3303);
and U6226 (N_6226,N_2690,N_3232);
nor U6227 (N_6227,N_4563,N_4974);
nor U6228 (N_6228,N_3120,N_2560);
and U6229 (N_6229,N_3714,N_4646);
and U6230 (N_6230,N_2885,N_4896);
xor U6231 (N_6231,N_4189,N_4989);
nand U6232 (N_6232,N_3812,N_2938);
nor U6233 (N_6233,N_2771,N_4788);
nor U6234 (N_6234,N_3437,N_4950);
or U6235 (N_6235,N_4281,N_3685);
and U6236 (N_6236,N_3890,N_4157);
and U6237 (N_6237,N_3982,N_4339);
or U6238 (N_6238,N_3504,N_3378);
and U6239 (N_6239,N_4753,N_2875);
nand U6240 (N_6240,N_3867,N_4380);
nor U6241 (N_6241,N_3952,N_4072);
or U6242 (N_6242,N_4533,N_3700);
or U6243 (N_6243,N_4571,N_4782);
nor U6244 (N_6244,N_3135,N_2891);
xor U6245 (N_6245,N_2653,N_4439);
nand U6246 (N_6246,N_3983,N_3453);
and U6247 (N_6247,N_2810,N_4540);
and U6248 (N_6248,N_3741,N_4425);
xnor U6249 (N_6249,N_3218,N_3141);
nand U6250 (N_6250,N_3396,N_4595);
nor U6251 (N_6251,N_3978,N_4181);
nor U6252 (N_6252,N_3578,N_2649);
xnor U6253 (N_6253,N_4529,N_3457);
and U6254 (N_6254,N_3958,N_4289);
nor U6255 (N_6255,N_3764,N_2719);
xnor U6256 (N_6256,N_2947,N_2991);
nand U6257 (N_6257,N_4692,N_4940);
xor U6258 (N_6258,N_4667,N_2777);
or U6259 (N_6259,N_3175,N_3355);
nor U6260 (N_6260,N_4516,N_3185);
nor U6261 (N_6261,N_4901,N_4954);
nor U6262 (N_6262,N_2980,N_2938);
nor U6263 (N_6263,N_4497,N_4829);
xnor U6264 (N_6264,N_4212,N_3858);
nand U6265 (N_6265,N_3044,N_3563);
and U6266 (N_6266,N_2671,N_4665);
or U6267 (N_6267,N_2972,N_3738);
and U6268 (N_6268,N_3743,N_3062);
xor U6269 (N_6269,N_3799,N_4584);
xor U6270 (N_6270,N_3093,N_4808);
and U6271 (N_6271,N_2803,N_4103);
nor U6272 (N_6272,N_3549,N_4062);
and U6273 (N_6273,N_4480,N_4382);
nand U6274 (N_6274,N_2619,N_3824);
or U6275 (N_6275,N_3122,N_3577);
xnor U6276 (N_6276,N_3936,N_4591);
or U6277 (N_6277,N_2962,N_4055);
xor U6278 (N_6278,N_4459,N_4246);
nor U6279 (N_6279,N_2951,N_4127);
and U6280 (N_6280,N_3338,N_2750);
nand U6281 (N_6281,N_3640,N_4795);
and U6282 (N_6282,N_4180,N_3825);
and U6283 (N_6283,N_3465,N_2612);
xor U6284 (N_6284,N_2599,N_2956);
nand U6285 (N_6285,N_4715,N_4932);
xnor U6286 (N_6286,N_4614,N_4306);
and U6287 (N_6287,N_3952,N_4702);
or U6288 (N_6288,N_4548,N_4329);
nand U6289 (N_6289,N_3669,N_3152);
nor U6290 (N_6290,N_3479,N_4755);
or U6291 (N_6291,N_4502,N_4007);
nand U6292 (N_6292,N_3097,N_4968);
nor U6293 (N_6293,N_2630,N_4071);
nand U6294 (N_6294,N_4224,N_2995);
nand U6295 (N_6295,N_3892,N_2790);
xor U6296 (N_6296,N_4271,N_4629);
and U6297 (N_6297,N_3488,N_3060);
and U6298 (N_6298,N_3951,N_4485);
and U6299 (N_6299,N_2917,N_3625);
nor U6300 (N_6300,N_4700,N_3574);
or U6301 (N_6301,N_4039,N_3459);
or U6302 (N_6302,N_2677,N_4001);
and U6303 (N_6303,N_4843,N_4011);
nand U6304 (N_6304,N_3213,N_2812);
and U6305 (N_6305,N_2881,N_4334);
or U6306 (N_6306,N_4173,N_3778);
and U6307 (N_6307,N_3738,N_3037);
nor U6308 (N_6308,N_4354,N_3354);
nor U6309 (N_6309,N_4043,N_4890);
or U6310 (N_6310,N_4088,N_3326);
nor U6311 (N_6311,N_2806,N_3579);
or U6312 (N_6312,N_3447,N_2940);
xnor U6313 (N_6313,N_3293,N_4013);
nor U6314 (N_6314,N_3800,N_4878);
or U6315 (N_6315,N_4646,N_4829);
xor U6316 (N_6316,N_2697,N_4896);
xor U6317 (N_6317,N_4371,N_3511);
xnor U6318 (N_6318,N_4701,N_4407);
and U6319 (N_6319,N_3513,N_3740);
or U6320 (N_6320,N_4970,N_4861);
and U6321 (N_6321,N_4850,N_3052);
nor U6322 (N_6322,N_3476,N_3292);
nor U6323 (N_6323,N_4825,N_4338);
or U6324 (N_6324,N_4992,N_3128);
xnor U6325 (N_6325,N_3549,N_2720);
xor U6326 (N_6326,N_4274,N_4444);
xnor U6327 (N_6327,N_3377,N_3423);
nand U6328 (N_6328,N_4883,N_3958);
or U6329 (N_6329,N_2673,N_3972);
nor U6330 (N_6330,N_4732,N_3964);
nand U6331 (N_6331,N_3976,N_3781);
nor U6332 (N_6332,N_3104,N_4415);
xnor U6333 (N_6333,N_3603,N_4902);
xor U6334 (N_6334,N_3091,N_3787);
or U6335 (N_6335,N_3993,N_3463);
or U6336 (N_6336,N_3747,N_3828);
nand U6337 (N_6337,N_3512,N_3525);
nor U6338 (N_6338,N_4291,N_3433);
xnor U6339 (N_6339,N_2737,N_4694);
or U6340 (N_6340,N_4119,N_4724);
or U6341 (N_6341,N_4045,N_3595);
nor U6342 (N_6342,N_4985,N_4279);
and U6343 (N_6343,N_4755,N_3417);
nor U6344 (N_6344,N_2758,N_2710);
nand U6345 (N_6345,N_3994,N_2864);
xnor U6346 (N_6346,N_3047,N_2812);
nand U6347 (N_6347,N_3079,N_3481);
nor U6348 (N_6348,N_3997,N_4054);
and U6349 (N_6349,N_2669,N_3939);
and U6350 (N_6350,N_4595,N_4935);
and U6351 (N_6351,N_2614,N_3544);
xnor U6352 (N_6352,N_4864,N_3449);
xor U6353 (N_6353,N_3639,N_4993);
or U6354 (N_6354,N_3450,N_3876);
xnor U6355 (N_6355,N_3629,N_4271);
xnor U6356 (N_6356,N_2964,N_4460);
and U6357 (N_6357,N_4039,N_4578);
nand U6358 (N_6358,N_3909,N_2806);
xnor U6359 (N_6359,N_3724,N_3571);
nor U6360 (N_6360,N_3707,N_3551);
and U6361 (N_6361,N_3674,N_4809);
nor U6362 (N_6362,N_3450,N_3808);
nand U6363 (N_6363,N_3114,N_4401);
or U6364 (N_6364,N_3754,N_4194);
nand U6365 (N_6365,N_4079,N_4208);
or U6366 (N_6366,N_3404,N_2549);
or U6367 (N_6367,N_4866,N_2747);
nand U6368 (N_6368,N_3990,N_4632);
or U6369 (N_6369,N_3177,N_4100);
nor U6370 (N_6370,N_3983,N_4019);
and U6371 (N_6371,N_3191,N_3597);
nor U6372 (N_6372,N_3638,N_4940);
and U6373 (N_6373,N_3614,N_3501);
or U6374 (N_6374,N_4138,N_4793);
or U6375 (N_6375,N_4072,N_4042);
and U6376 (N_6376,N_2825,N_3824);
and U6377 (N_6377,N_4619,N_3542);
or U6378 (N_6378,N_4480,N_2836);
nor U6379 (N_6379,N_2785,N_3832);
or U6380 (N_6380,N_3303,N_4812);
or U6381 (N_6381,N_3918,N_3541);
xor U6382 (N_6382,N_2642,N_4186);
xnor U6383 (N_6383,N_4908,N_4961);
and U6384 (N_6384,N_4156,N_3904);
and U6385 (N_6385,N_4718,N_3249);
or U6386 (N_6386,N_3911,N_3433);
or U6387 (N_6387,N_4763,N_3036);
xor U6388 (N_6388,N_4959,N_3269);
nand U6389 (N_6389,N_4451,N_4387);
xor U6390 (N_6390,N_4600,N_3225);
and U6391 (N_6391,N_3653,N_4521);
nand U6392 (N_6392,N_3229,N_4378);
or U6393 (N_6393,N_3075,N_4174);
and U6394 (N_6394,N_4095,N_2950);
nand U6395 (N_6395,N_4221,N_3580);
or U6396 (N_6396,N_3019,N_2716);
xnor U6397 (N_6397,N_4982,N_3331);
nor U6398 (N_6398,N_3706,N_4795);
nor U6399 (N_6399,N_4804,N_3525);
or U6400 (N_6400,N_2722,N_3166);
nor U6401 (N_6401,N_4961,N_4074);
xnor U6402 (N_6402,N_4481,N_4227);
nor U6403 (N_6403,N_3134,N_3386);
nand U6404 (N_6404,N_4876,N_2816);
nand U6405 (N_6405,N_4761,N_3000);
xor U6406 (N_6406,N_3299,N_2528);
or U6407 (N_6407,N_2512,N_3771);
or U6408 (N_6408,N_2938,N_4695);
and U6409 (N_6409,N_3554,N_4098);
xnor U6410 (N_6410,N_4777,N_4482);
or U6411 (N_6411,N_2922,N_3805);
xor U6412 (N_6412,N_3316,N_3843);
nand U6413 (N_6413,N_3470,N_3189);
xnor U6414 (N_6414,N_4751,N_3284);
nor U6415 (N_6415,N_4306,N_4438);
nand U6416 (N_6416,N_4379,N_4894);
xor U6417 (N_6417,N_2548,N_2658);
and U6418 (N_6418,N_4791,N_4345);
nand U6419 (N_6419,N_4080,N_4123);
nor U6420 (N_6420,N_3950,N_2516);
nor U6421 (N_6421,N_2598,N_3981);
nand U6422 (N_6422,N_2614,N_3356);
nand U6423 (N_6423,N_4895,N_4125);
nor U6424 (N_6424,N_3758,N_4303);
xnor U6425 (N_6425,N_3033,N_4654);
and U6426 (N_6426,N_4085,N_3940);
and U6427 (N_6427,N_2549,N_4016);
xor U6428 (N_6428,N_3629,N_2810);
or U6429 (N_6429,N_2836,N_3666);
or U6430 (N_6430,N_4268,N_3399);
nor U6431 (N_6431,N_2985,N_3099);
and U6432 (N_6432,N_3215,N_4791);
nand U6433 (N_6433,N_3199,N_3059);
and U6434 (N_6434,N_3017,N_3488);
nor U6435 (N_6435,N_4045,N_2762);
nand U6436 (N_6436,N_4517,N_4350);
and U6437 (N_6437,N_2893,N_4621);
and U6438 (N_6438,N_3388,N_2976);
xnor U6439 (N_6439,N_3446,N_2551);
xor U6440 (N_6440,N_2567,N_4659);
xor U6441 (N_6441,N_4001,N_3587);
nor U6442 (N_6442,N_2772,N_2854);
or U6443 (N_6443,N_3084,N_4016);
or U6444 (N_6444,N_3979,N_3060);
or U6445 (N_6445,N_3910,N_2793);
and U6446 (N_6446,N_2694,N_4711);
xor U6447 (N_6447,N_4353,N_3949);
and U6448 (N_6448,N_3658,N_3054);
xor U6449 (N_6449,N_3444,N_3224);
and U6450 (N_6450,N_2992,N_3636);
nand U6451 (N_6451,N_4474,N_3038);
nand U6452 (N_6452,N_4125,N_4238);
nand U6453 (N_6453,N_4844,N_3025);
and U6454 (N_6454,N_4736,N_2978);
nand U6455 (N_6455,N_3103,N_2800);
and U6456 (N_6456,N_3615,N_4393);
nand U6457 (N_6457,N_4876,N_2744);
nand U6458 (N_6458,N_4560,N_4411);
nand U6459 (N_6459,N_3821,N_3114);
and U6460 (N_6460,N_4192,N_4213);
or U6461 (N_6461,N_3742,N_3246);
nand U6462 (N_6462,N_4399,N_4726);
or U6463 (N_6463,N_4730,N_2548);
or U6464 (N_6464,N_3208,N_2811);
xnor U6465 (N_6465,N_4252,N_3888);
or U6466 (N_6466,N_4627,N_2881);
or U6467 (N_6467,N_3428,N_3781);
nor U6468 (N_6468,N_2766,N_4197);
nand U6469 (N_6469,N_4733,N_4432);
or U6470 (N_6470,N_3158,N_4089);
and U6471 (N_6471,N_2932,N_3164);
nand U6472 (N_6472,N_2809,N_3241);
or U6473 (N_6473,N_3601,N_4659);
and U6474 (N_6474,N_4849,N_4224);
xor U6475 (N_6475,N_3587,N_4079);
and U6476 (N_6476,N_4082,N_3379);
or U6477 (N_6477,N_2552,N_2780);
and U6478 (N_6478,N_2919,N_2876);
and U6479 (N_6479,N_3937,N_4920);
xnor U6480 (N_6480,N_2660,N_4074);
and U6481 (N_6481,N_4612,N_4546);
nand U6482 (N_6482,N_3077,N_3107);
nand U6483 (N_6483,N_3536,N_3616);
xnor U6484 (N_6484,N_4989,N_4347);
or U6485 (N_6485,N_3516,N_2777);
or U6486 (N_6486,N_2583,N_4139);
and U6487 (N_6487,N_3885,N_4257);
or U6488 (N_6488,N_3342,N_3553);
nand U6489 (N_6489,N_2648,N_3554);
nor U6490 (N_6490,N_4015,N_4989);
or U6491 (N_6491,N_3812,N_3383);
or U6492 (N_6492,N_4014,N_4086);
xor U6493 (N_6493,N_3464,N_3211);
and U6494 (N_6494,N_4916,N_3753);
nand U6495 (N_6495,N_4794,N_3628);
nand U6496 (N_6496,N_2700,N_2677);
and U6497 (N_6497,N_4953,N_4856);
and U6498 (N_6498,N_3511,N_4569);
nor U6499 (N_6499,N_3690,N_4674);
nand U6500 (N_6500,N_3202,N_3987);
nand U6501 (N_6501,N_3899,N_4974);
or U6502 (N_6502,N_3292,N_2506);
and U6503 (N_6503,N_2708,N_2935);
and U6504 (N_6504,N_3379,N_3652);
or U6505 (N_6505,N_4079,N_3571);
or U6506 (N_6506,N_3378,N_2814);
or U6507 (N_6507,N_4537,N_3809);
or U6508 (N_6508,N_3756,N_4767);
nand U6509 (N_6509,N_4386,N_3942);
or U6510 (N_6510,N_4081,N_3986);
and U6511 (N_6511,N_2523,N_3738);
or U6512 (N_6512,N_2806,N_3194);
or U6513 (N_6513,N_3305,N_2670);
and U6514 (N_6514,N_3303,N_4354);
or U6515 (N_6515,N_4149,N_3301);
nand U6516 (N_6516,N_4804,N_2578);
nand U6517 (N_6517,N_2988,N_4647);
xnor U6518 (N_6518,N_3860,N_4646);
and U6519 (N_6519,N_4377,N_2762);
nand U6520 (N_6520,N_3987,N_2632);
and U6521 (N_6521,N_4111,N_2600);
nor U6522 (N_6522,N_4159,N_4643);
xor U6523 (N_6523,N_3066,N_3540);
and U6524 (N_6524,N_4953,N_4469);
and U6525 (N_6525,N_3877,N_4936);
and U6526 (N_6526,N_4206,N_2518);
and U6527 (N_6527,N_3230,N_2916);
and U6528 (N_6528,N_2502,N_3265);
or U6529 (N_6529,N_4961,N_3046);
nor U6530 (N_6530,N_2513,N_4420);
nor U6531 (N_6531,N_4261,N_2508);
xnor U6532 (N_6532,N_2986,N_3702);
xnor U6533 (N_6533,N_3054,N_2907);
and U6534 (N_6534,N_3212,N_3898);
nor U6535 (N_6535,N_3258,N_3808);
or U6536 (N_6536,N_4815,N_3691);
nor U6537 (N_6537,N_2930,N_4910);
xnor U6538 (N_6538,N_4502,N_4260);
xnor U6539 (N_6539,N_3217,N_3158);
and U6540 (N_6540,N_3298,N_3692);
and U6541 (N_6541,N_3818,N_3530);
and U6542 (N_6542,N_2733,N_4919);
nor U6543 (N_6543,N_2735,N_4070);
or U6544 (N_6544,N_2732,N_3738);
nor U6545 (N_6545,N_3820,N_3857);
nand U6546 (N_6546,N_3812,N_3501);
and U6547 (N_6547,N_2532,N_3227);
and U6548 (N_6548,N_4934,N_3247);
nor U6549 (N_6549,N_2562,N_2974);
nor U6550 (N_6550,N_2684,N_3258);
nand U6551 (N_6551,N_3306,N_3580);
and U6552 (N_6552,N_4373,N_4487);
or U6553 (N_6553,N_4031,N_2854);
or U6554 (N_6554,N_4233,N_4808);
and U6555 (N_6555,N_3837,N_4557);
nand U6556 (N_6556,N_2695,N_4125);
or U6557 (N_6557,N_2582,N_4493);
and U6558 (N_6558,N_4744,N_4855);
and U6559 (N_6559,N_3236,N_3372);
or U6560 (N_6560,N_2630,N_4888);
nor U6561 (N_6561,N_3854,N_2582);
xor U6562 (N_6562,N_3794,N_4425);
nand U6563 (N_6563,N_4368,N_4004);
nand U6564 (N_6564,N_4357,N_4683);
and U6565 (N_6565,N_4578,N_3674);
nand U6566 (N_6566,N_3676,N_4000);
nor U6567 (N_6567,N_2519,N_4058);
nor U6568 (N_6568,N_2843,N_3636);
or U6569 (N_6569,N_4914,N_2539);
nor U6570 (N_6570,N_3074,N_3438);
or U6571 (N_6571,N_4471,N_3409);
xnor U6572 (N_6572,N_3356,N_4262);
xor U6573 (N_6573,N_4127,N_3429);
nand U6574 (N_6574,N_2756,N_4923);
nand U6575 (N_6575,N_4012,N_4955);
xnor U6576 (N_6576,N_3374,N_4415);
nand U6577 (N_6577,N_3388,N_3937);
and U6578 (N_6578,N_4520,N_2713);
nand U6579 (N_6579,N_4458,N_2511);
xnor U6580 (N_6580,N_3652,N_4765);
xor U6581 (N_6581,N_2907,N_4037);
nand U6582 (N_6582,N_4595,N_3086);
or U6583 (N_6583,N_4628,N_4998);
or U6584 (N_6584,N_3353,N_4361);
and U6585 (N_6585,N_3485,N_3809);
and U6586 (N_6586,N_3850,N_3276);
nor U6587 (N_6587,N_4108,N_3870);
or U6588 (N_6588,N_4125,N_4864);
xor U6589 (N_6589,N_2661,N_4484);
nor U6590 (N_6590,N_3838,N_3376);
and U6591 (N_6591,N_4256,N_3759);
xor U6592 (N_6592,N_2761,N_2577);
nand U6593 (N_6593,N_3593,N_4087);
or U6594 (N_6594,N_3645,N_3958);
and U6595 (N_6595,N_3539,N_2711);
nand U6596 (N_6596,N_4379,N_3742);
or U6597 (N_6597,N_3780,N_3044);
or U6598 (N_6598,N_4496,N_2541);
and U6599 (N_6599,N_3440,N_2892);
and U6600 (N_6600,N_3225,N_4259);
nor U6601 (N_6601,N_4976,N_4332);
xnor U6602 (N_6602,N_3895,N_3968);
xor U6603 (N_6603,N_2646,N_2692);
and U6604 (N_6604,N_4956,N_2851);
xnor U6605 (N_6605,N_2654,N_3813);
nor U6606 (N_6606,N_3986,N_4684);
or U6607 (N_6607,N_4332,N_4334);
or U6608 (N_6608,N_3416,N_3603);
nand U6609 (N_6609,N_2910,N_4948);
and U6610 (N_6610,N_2665,N_3610);
nor U6611 (N_6611,N_4288,N_3233);
nor U6612 (N_6612,N_3953,N_4929);
xor U6613 (N_6613,N_4185,N_3348);
nor U6614 (N_6614,N_4125,N_2505);
or U6615 (N_6615,N_2502,N_4064);
nor U6616 (N_6616,N_2965,N_4477);
or U6617 (N_6617,N_3537,N_3195);
and U6618 (N_6618,N_3580,N_4420);
nand U6619 (N_6619,N_4933,N_2659);
nor U6620 (N_6620,N_3527,N_3413);
nand U6621 (N_6621,N_3696,N_2576);
xor U6622 (N_6622,N_4303,N_4579);
nand U6623 (N_6623,N_3199,N_4516);
nand U6624 (N_6624,N_4966,N_4347);
nor U6625 (N_6625,N_3357,N_3609);
or U6626 (N_6626,N_3635,N_3394);
xor U6627 (N_6627,N_2561,N_4810);
xnor U6628 (N_6628,N_2515,N_3140);
xnor U6629 (N_6629,N_4421,N_4239);
or U6630 (N_6630,N_3221,N_4836);
nor U6631 (N_6631,N_3093,N_3942);
nor U6632 (N_6632,N_4792,N_4904);
xor U6633 (N_6633,N_4453,N_2616);
or U6634 (N_6634,N_4776,N_2990);
xor U6635 (N_6635,N_3713,N_4113);
nand U6636 (N_6636,N_3812,N_4892);
and U6637 (N_6637,N_3603,N_2860);
xor U6638 (N_6638,N_4152,N_3868);
and U6639 (N_6639,N_3214,N_2506);
and U6640 (N_6640,N_4472,N_3952);
or U6641 (N_6641,N_3940,N_2827);
and U6642 (N_6642,N_2705,N_3172);
and U6643 (N_6643,N_4599,N_2538);
nand U6644 (N_6644,N_4688,N_2546);
xnor U6645 (N_6645,N_3228,N_3966);
and U6646 (N_6646,N_4475,N_3200);
nor U6647 (N_6647,N_3850,N_3556);
and U6648 (N_6648,N_2525,N_4168);
nand U6649 (N_6649,N_3344,N_3124);
xor U6650 (N_6650,N_4233,N_4142);
xnor U6651 (N_6651,N_3474,N_3606);
and U6652 (N_6652,N_3685,N_4711);
nor U6653 (N_6653,N_2684,N_4983);
nor U6654 (N_6654,N_3508,N_3241);
or U6655 (N_6655,N_2896,N_4388);
or U6656 (N_6656,N_4225,N_3825);
and U6657 (N_6657,N_4816,N_3989);
nand U6658 (N_6658,N_4395,N_4644);
nor U6659 (N_6659,N_4366,N_4092);
and U6660 (N_6660,N_3072,N_4765);
xnor U6661 (N_6661,N_2913,N_4200);
or U6662 (N_6662,N_2972,N_4668);
xnor U6663 (N_6663,N_2919,N_3632);
nand U6664 (N_6664,N_2934,N_4039);
nor U6665 (N_6665,N_3658,N_3356);
xor U6666 (N_6666,N_4904,N_3987);
xnor U6667 (N_6667,N_3941,N_4189);
xor U6668 (N_6668,N_4827,N_3294);
or U6669 (N_6669,N_2657,N_3529);
xnor U6670 (N_6670,N_2710,N_2994);
nand U6671 (N_6671,N_3715,N_4756);
or U6672 (N_6672,N_4244,N_4133);
xor U6673 (N_6673,N_4860,N_4294);
and U6674 (N_6674,N_4562,N_4560);
xnor U6675 (N_6675,N_4121,N_3879);
nor U6676 (N_6676,N_2790,N_3385);
nor U6677 (N_6677,N_2842,N_3074);
or U6678 (N_6678,N_2644,N_3860);
and U6679 (N_6679,N_4157,N_4165);
or U6680 (N_6680,N_3497,N_4317);
xnor U6681 (N_6681,N_4196,N_2796);
or U6682 (N_6682,N_3429,N_2638);
nand U6683 (N_6683,N_3725,N_2997);
xor U6684 (N_6684,N_4700,N_4275);
and U6685 (N_6685,N_3449,N_3842);
and U6686 (N_6686,N_4563,N_3490);
xnor U6687 (N_6687,N_3486,N_4369);
and U6688 (N_6688,N_2602,N_3069);
xnor U6689 (N_6689,N_4566,N_4086);
nand U6690 (N_6690,N_3322,N_4462);
or U6691 (N_6691,N_4487,N_2629);
or U6692 (N_6692,N_4648,N_3383);
nand U6693 (N_6693,N_4081,N_3646);
nor U6694 (N_6694,N_3210,N_4602);
or U6695 (N_6695,N_4391,N_4923);
xor U6696 (N_6696,N_3314,N_4536);
xnor U6697 (N_6697,N_4223,N_4919);
nor U6698 (N_6698,N_3217,N_4758);
and U6699 (N_6699,N_3433,N_4337);
nor U6700 (N_6700,N_3359,N_2876);
or U6701 (N_6701,N_2778,N_4741);
nor U6702 (N_6702,N_3261,N_4800);
xnor U6703 (N_6703,N_3362,N_4972);
nor U6704 (N_6704,N_3975,N_4657);
xnor U6705 (N_6705,N_4032,N_3872);
or U6706 (N_6706,N_3209,N_4045);
nand U6707 (N_6707,N_4226,N_2822);
or U6708 (N_6708,N_3314,N_4985);
nand U6709 (N_6709,N_3439,N_2593);
nor U6710 (N_6710,N_4792,N_2613);
or U6711 (N_6711,N_2629,N_4147);
and U6712 (N_6712,N_4311,N_3340);
nand U6713 (N_6713,N_2869,N_4774);
nor U6714 (N_6714,N_2891,N_4972);
nor U6715 (N_6715,N_2762,N_4177);
nand U6716 (N_6716,N_2713,N_3267);
nand U6717 (N_6717,N_4133,N_2580);
xor U6718 (N_6718,N_4153,N_2606);
nor U6719 (N_6719,N_3813,N_3097);
nand U6720 (N_6720,N_4905,N_3047);
and U6721 (N_6721,N_4082,N_2515);
or U6722 (N_6722,N_4918,N_3142);
and U6723 (N_6723,N_3519,N_3706);
nand U6724 (N_6724,N_3256,N_4118);
or U6725 (N_6725,N_3241,N_4047);
or U6726 (N_6726,N_3501,N_2994);
and U6727 (N_6727,N_2547,N_3863);
or U6728 (N_6728,N_3050,N_2734);
nor U6729 (N_6729,N_4069,N_3238);
nor U6730 (N_6730,N_4836,N_2817);
or U6731 (N_6731,N_4380,N_2937);
xor U6732 (N_6732,N_2852,N_4590);
and U6733 (N_6733,N_3270,N_4665);
xor U6734 (N_6734,N_4783,N_4272);
and U6735 (N_6735,N_3786,N_3717);
xor U6736 (N_6736,N_4620,N_2830);
or U6737 (N_6737,N_3756,N_3943);
and U6738 (N_6738,N_2729,N_4035);
nor U6739 (N_6739,N_3835,N_4622);
nor U6740 (N_6740,N_3505,N_2583);
and U6741 (N_6741,N_2973,N_4249);
nand U6742 (N_6742,N_3012,N_4907);
nor U6743 (N_6743,N_4011,N_2608);
and U6744 (N_6744,N_4148,N_4344);
and U6745 (N_6745,N_2833,N_4309);
nand U6746 (N_6746,N_4770,N_2615);
or U6747 (N_6747,N_2970,N_3447);
or U6748 (N_6748,N_3586,N_3286);
or U6749 (N_6749,N_4090,N_3080);
nand U6750 (N_6750,N_3949,N_3553);
or U6751 (N_6751,N_4756,N_2536);
xor U6752 (N_6752,N_2891,N_2631);
nand U6753 (N_6753,N_4271,N_3191);
xor U6754 (N_6754,N_3198,N_4694);
and U6755 (N_6755,N_4734,N_3851);
nor U6756 (N_6756,N_3690,N_3199);
and U6757 (N_6757,N_2999,N_3360);
xor U6758 (N_6758,N_4054,N_2989);
and U6759 (N_6759,N_3780,N_2579);
nand U6760 (N_6760,N_3323,N_3276);
or U6761 (N_6761,N_3663,N_4409);
nor U6762 (N_6762,N_2614,N_4771);
and U6763 (N_6763,N_3547,N_3402);
xnor U6764 (N_6764,N_4202,N_4552);
or U6765 (N_6765,N_3295,N_4895);
or U6766 (N_6766,N_3799,N_4094);
and U6767 (N_6767,N_3419,N_4241);
or U6768 (N_6768,N_4530,N_2567);
nand U6769 (N_6769,N_2915,N_2935);
or U6770 (N_6770,N_3081,N_2734);
and U6771 (N_6771,N_3656,N_4843);
xnor U6772 (N_6772,N_4810,N_4195);
nor U6773 (N_6773,N_4745,N_4430);
nand U6774 (N_6774,N_4470,N_2842);
and U6775 (N_6775,N_4935,N_2715);
nand U6776 (N_6776,N_4601,N_3960);
and U6777 (N_6777,N_4756,N_4243);
nand U6778 (N_6778,N_3262,N_4290);
xor U6779 (N_6779,N_2635,N_2621);
or U6780 (N_6780,N_4473,N_4042);
and U6781 (N_6781,N_4362,N_4002);
nand U6782 (N_6782,N_3065,N_3813);
nor U6783 (N_6783,N_4055,N_4066);
nor U6784 (N_6784,N_4156,N_4687);
nand U6785 (N_6785,N_3510,N_3452);
and U6786 (N_6786,N_4458,N_3514);
xor U6787 (N_6787,N_3894,N_3717);
xor U6788 (N_6788,N_2901,N_4601);
or U6789 (N_6789,N_3630,N_3628);
nor U6790 (N_6790,N_3000,N_4110);
nor U6791 (N_6791,N_3564,N_4748);
nor U6792 (N_6792,N_3162,N_3831);
and U6793 (N_6793,N_4554,N_3496);
and U6794 (N_6794,N_2637,N_4134);
nand U6795 (N_6795,N_2690,N_3195);
nor U6796 (N_6796,N_2520,N_4087);
nand U6797 (N_6797,N_4931,N_3073);
nand U6798 (N_6798,N_3622,N_3011);
nor U6799 (N_6799,N_3055,N_4744);
nor U6800 (N_6800,N_4848,N_4748);
or U6801 (N_6801,N_4017,N_4578);
nand U6802 (N_6802,N_2683,N_4953);
nor U6803 (N_6803,N_4617,N_3176);
and U6804 (N_6804,N_4147,N_4699);
or U6805 (N_6805,N_2740,N_2993);
or U6806 (N_6806,N_3085,N_3938);
and U6807 (N_6807,N_4985,N_2776);
and U6808 (N_6808,N_2506,N_4644);
nor U6809 (N_6809,N_2602,N_3787);
or U6810 (N_6810,N_4332,N_3363);
nor U6811 (N_6811,N_4313,N_4102);
or U6812 (N_6812,N_4782,N_4704);
and U6813 (N_6813,N_3894,N_4068);
or U6814 (N_6814,N_3187,N_2692);
nand U6815 (N_6815,N_4958,N_4304);
xnor U6816 (N_6816,N_3953,N_3936);
nand U6817 (N_6817,N_3650,N_4367);
nand U6818 (N_6818,N_3855,N_3770);
nand U6819 (N_6819,N_3097,N_2524);
nor U6820 (N_6820,N_3976,N_2524);
and U6821 (N_6821,N_4755,N_4291);
xor U6822 (N_6822,N_3031,N_3132);
nand U6823 (N_6823,N_4580,N_4864);
nand U6824 (N_6824,N_3033,N_4280);
xnor U6825 (N_6825,N_3446,N_4378);
xnor U6826 (N_6826,N_2846,N_3880);
nand U6827 (N_6827,N_3239,N_3999);
or U6828 (N_6828,N_3317,N_3663);
and U6829 (N_6829,N_3670,N_2872);
nor U6830 (N_6830,N_4503,N_2792);
xor U6831 (N_6831,N_2901,N_4741);
xor U6832 (N_6832,N_4767,N_3997);
xnor U6833 (N_6833,N_4226,N_4033);
xor U6834 (N_6834,N_4879,N_3834);
nand U6835 (N_6835,N_3405,N_2975);
and U6836 (N_6836,N_3823,N_4780);
nor U6837 (N_6837,N_2653,N_4583);
xor U6838 (N_6838,N_2875,N_3130);
nor U6839 (N_6839,N_4118,N_4753);
xor U6840 (N_6840,N_4679,N_3414);
and U6841 (N_6841,N_3333,N_2826);
nand U6842 (N_6842,N_3415,N_2574);
or U6843 (N_6843,N_3788,N_4954);
and U6844 (N_6844,N_3792,N_3311);
nor U6845 (N_6845,N_4384,N_3144);
or U6846 (N_6846,N_4650,N_4699);
nand U6847 (N_6847,N_4077,N_4719);
xor U6848 (N_6848,N_3203,N_2752);
or U6849 (N_6849,N_4786,N_3063);
nand U6850 (N_6850,N_4313,N_4747);
nor U6851 (N_6851,N_3859,N_3005);
nand U6852 (N_6852,N_4896,N_4093);
nand U6853 (N_6853,N_3011,N_3245);
nand U6854 (N_6854,N_2577,N_2525);
nor U6855 (N_6855,N_3175,N_3602);
xor U6856 (N_6856,N_4589,N_4354);
xnor U6857 (N_6857,N_4838,N_4521);
nor U6858 (N_6858,N_3231,N_4578);
and U6859 (N_6859,N_2976,N_3209);
or U6860 (N_6860,N_4939,N_3364);
nand U6861 (N_6861,N_4878,N_3955);
xnor U6862 (N_6862,N_4164,N_4561);
xnor U6863 (N_6863,N_4909,N_2847);
nand U6864 (N_6864,N_4070,N_2679);
nand U6865 (N_6865,N_2821,N_4642);
and U6866 (N_6866,N_2719,N_3369);
or U6867 (N_6867,N_3804,N_3685);
nand U6868 (N_6868,N_4585,N_4942);
or U6869 (N_6869,N_2956,N_3096);
xnor U6870 (N_6870,N_4980,N_4632);
nand U6871 (N_6871,N_3775,N_3008);
or U6872 (N_6872,N_3745,N_3474);
nand U6873 (N_6873,N_2939,N_3213);
nand U6874 (N_6874,N_4380,N_4937);
and U6875 (N_6875,N_4291,N_4244);
nand U6876 (N_6876,N_2622,N_3313);
and U6877 (N_6877,N_4859,N_4267);
xnor U6878 (N_6878,N_4269,N_3163);
and U6879 (N_6879,N_4957,N_3308);
and U6880 (N_6880,N_4774,N_3540);
xor U6881 (N_6881,N_4388,N_4236);
xor U6882 (N_6882,N_2937,N_4731);
or U6883 (N_6883,N_3327,N_4531);
or U6884 (N_6884,N_3977,N_2506);
nand U6885 (N_6885,N_2999,N_3893);
nand U6886 (N_6886,N_2824,N_4983);
and U6887 (N_6887,N_4519,N_3371);
and U6888 (N_6888,N_2858,N_4598);
nand U6889 (N_6889,N_2991,N_4748);
xor U6890 (N_6890,N_3809,N_4288);
xor U6891 (N_6891,N_3807,N_2820);
nand U6892 (N_6892,N_2764,N_4459);
xor U6893 (N_6893,N_4355,N_3707);
nand U6894 (N_6894,N_4392,N_4669);
xor U6895 (N_6895,N_3565,N_3147);
or U6896 (N_6896,N_4423,N_3375);
xnor U6897 (N_6897,N_4312,N_4509);
xor U6898 (N_6898,N_4526,N_4145);
or U6899 (N_6899,N_3750,N_4543);
nand U6900 (N_6900,N_2857,N_3378);
or U6901 (N_6901,N_2553,N_3068);
nor U6902 (N_6902,N_3011,N_3891);
xnor U6903 (N_6903,N_2568,N_3546);
or U6904 (N_6904,N_4707,N_3783);
nor U6905 (N_6905,N_4326,N_3506);
xor U6906 (N_6906,N_2970,N_3722);
or U6907 (N_6907,N_2538,N_3090);
and U6908 (N_6908,N_2673,N_3454);
nor U6909 (N_6909,N_3417,N_3594);
nor U6910 (N_6910,N_4649,N_4656);
or U6911 (N_6911,N_4365,N_4020);
nand U6912 (N_6912,N_3285,N_2806);
nand U6913 (N_6913,N_3816,N_3296);
nand U6914 (N_6914,N_3497,N_4825);
nand U6915 (N_6915,N_4723,N_3004);
nor U6916 (N_6916,N_3392,N_4260);
or U6917 (N_6917,N_4579,N_3173);
xnor U6918 (N_6918,N_4657,N_3325);
xor U6919 (N_6919,N_3605,N_4972);
nand U6920 (N_6920,N_3351,N_3259);
xnor U6921 (N_6921,N_4703,N_4647);
or U6922 (N_6922,N_4172,N_2639);
xnor U6923 (N_6923,N_4350,N_4471);
and U6924 (N_6924,N_3074,N_3840);
nor U6925 (N_6925,N_3645,N_4082);
xnor U6926 (N_6926,N_2978,N_3072);
nand U6927 (N_6927,N_2706,N_2718);
nor U6928 (N_6928,N_3210,N_3418);
or U6929 (N_6929,N_4377,N_4633);
nand U6930 (N_6930,N_2583,N_4473);
nor U6931 (N_6931,N_4659,N_3458);
nand U6932 (N_6932,N_4488,N_3208);
xor U6933 (N_6933,N_4080,N_4103);
nor U6934 (N_6934,N_4223,N_3282);
nand U6935 (N_6935,N_3397,N_4858);
nor U6936 (N_6936,N_4201,N_3140);
or U6937 (N_6937,N_3011,N_2580);
nand U6938 (N_6938,N_3070,N_2989);
xor U6939 (N_6939,N_4676,N_3836);
nand U6940 (N_6940,N_3488,N_3259);
xor U6941 (N_6941,N_4442,N_3965);
and U6942 (N_6942,N_4176,N_3294);
xor U6943 (N_6943,N_4651,N_4458);
and U6944 (N_6944,N_4952,N_3729);
xnor U6945 (N_6945,N_2687,N_2545);
and U6946 (N_6946,N_2707,N_3360);
nand U6947 (N_6947,N_2998,N_4368);
nand U6948 (N_6948,N_3700,N_3134);
nor U6949 (N_6949,N_3911,N_3642);
xor U6950 (N_6950,N_3489,N_3319);
and U6951 (N_6951,N_3373,N_3085);
xnor U6952 (N_6952,N_4204,N_4815);
and U6953 (N_6953,N_4330,N_4515);
xor U6954 (N_6954,N_4332,N_4410);
and U6955 (N_6955,N_2876,N_3533);
xnor U6956 (N_6956,N_4861,N_4452);
nor U6957 (N_6957,N_3537,N_2629);
xnor U6958 (N_6958,N_3900,N_3480);
xor U6959 (N_6959,N_4638,N_3534);
nor U6960 (N_6960,N_4701,N_4138);
nand U6961 (N_6961,N_3559,N_4153);
or U6962 (N_6962,N_3815,N_4739);
nand U6963 (N_6963,N_3462,N_4390);
xor U6964 (N_6964,N_4748,N_2954);
or U6965 (N_6965,N_3428,N_2827);
or U6966 (N_6966,N_2739,N_4770);
nand U6967 (N_6967,N_4216,N_2859);
or U6968 (N_6968,N_2726,N_2568);
nand U6969 (N_6969,N_4844,N_3895);
nand U6970 (N_6970,N_3603,N_3877);
nor U6971 (N_6971,N_3113,N_4530);
nand U6972 (N_6972,N_4954,N_3158);
xnor U6973 (N_6973,N_3040,N_4659);
or U6974 (N_6974,N_2580,N_4729);
xnor U6975 (N_6975,N_4914,N_4927);
nor U6976 (N_6976,N_4440,N_3466);
or U6977 (N_6977,N_3297,N_4679);
xor U6978 (N_6978,N_4703,N_3133);
and U6979 (N_6979,N_3209,N_4482);
or U6980 (N_6980,N_2932,N_2996);
xnor U6981 (N_6981,N_3439,N_4315);
xnor U6982 (N_6982,N_4023,N_4161);
nor U6983 (N_6983,N_3812,N_3413);
or U6984 (N_6984,N_3862,N_3688);
xor U6985 (N_6985,N_3574,N_4684);
or U6986 (N_6986,N_3580,N_3084);
nand U6987 (N_6987,N_3822,N_4414);
nand U6988 (N_6988,N_3382,N_4673);
nor U6989 (N_6989,N_3601,N_2879);
and U6990 (N_6990,N_3669,N_3177);
xor U6991 (N_6991,N_4463,N_4962);
or U6992 (N_6992,N_2820,N_2507);
xnor U6993 (N_6993,N_4762,N_2524);
nand U6994 (N_6994,N_4348,N_4968);
nor U6995 (N_6995,N_3036,N_4569);
nor U6996 (N_6996,N_3617,N_4556);
nand U6997 (N_6997,N_4889,N_3055);
nor U6998 (N_6998,N_4574,N_4976);
nand U6999 (N_6999,N_3387,N_3070);
xor U7000 (N_7000,N_2899,N_3009);
xnor U7001 (N_7001,N_4693,N_3081);
and U7002 (N_7002,N_4903,N_4729);
and U7003 (N_7003,N_4817,N_4700);
nand U7004 (N_7004,N_3879,N_4859);
or U7005 (N_7005,N_4647,N_3490);
xnor U7006 (N_7006,N_4137,N_3509);
or U7007 (N_7007,N_3133,N_2539);
xor U7008 (N_7008,N_3250,N_3620);
nor U7009 (N_7009,N_3132,N_4898);
and U7010 (N_7010,N_4223,N_2526);
nor U7011 (N_7011,N_4784,N_3939);
nor U7012 (N_7012,N_4837,N_4601);
and U7013 (N_7013,N_3362,N_3280);
xnor U7014 (N_7014,N_2950,N_3807);
xor U7015 (N_7015,N_4090,N_2668);
and U7016 (N_7016,N_3402,N_4924);
and U7017 (N_7017,N_4138,N_4751);
and U7018 (N_7018,N_3669,N_3006);
and U7019 (N_7019,N_4414,N_4284);
or U7020 (N_7020,N_3249,N_3017);
or U7021 (N_7021,N_2585,N_4910);
nand U7022 (N_7022,N_4685,N_4782);
and U7023 (N_7023,N_4606,N_4827);
and U7024 (N_7024,N_2823,N_3785);
xnor U7025 (N_7025,N_3742,N_3066);
nor U7026 (N_7026,N_2662,N_3820);
or U7027 (N_7027,N_4818,N_4192);
nor U7028 (N_7028,N_4834,N_3971);
nand U7029 (N_7029,N_4247,N_4303);
xnor U7030 (N_7030,N_2905,N_4095);
nor U7031 (N_7031,N_3547,N_2891);
and U7032 (N_7032,N_3807,N_3765);
nor U7033 (N_7033,N_2977,N_2931);
or U7034 (N_7034,N_3950,N_3363);
nor U7035 (N_7035,N_3633,N_4527);
nand U7036 (N_7036,N_3215,N_3611);
and U7037 (N_7037,N_2597,N_2939);
or U7038 (N_7038,N_4681,N_3387);
and U7039 (N_7039,N_2889,N_3347);
and U7040 (N_7040,N_3924,N_3414);
or U7041 (N_7041,N_2558,N_2919);
nor U7042 (N_7042,N_4518,N_2800);
or U7043 (N_7043,N_4784,N_4821);
and U7044 (N_7044,N_3520,N_3294);
nor U7045 (N_7045,N_3099,N_3923);
xor U7046 (N_7046,N_3053,N_4102);
nand U7047 (N_7047,N_4692,N_3696);
xnor U7048 (N_7048,N_4691,N_3706);
and U7049 (N_7049,N_2801,N_3565);
nor U7050 (N_7050,N_2525,N_2738);
and U7051 (N_7051,N_3373,N_4655);
nor U7052 (N_7052,N_4602,N_4914);
or U7053 (N_7053,N_2539,N_4739);
xor U7054 (N_7054,N_4317,N_3516);
nand U7055 (N_7055,N_3294,N_3848);
or U7056 (N_7056,N_4530,N_4479);
or U7057 (N_7057,N_4022,N_3932);
nor U7058 (N_7058,N_3555,N_3966);
or U7059 (N_7059,N_4694,N_4724);
or U7060 (N_7060,N_2567,N_2702);
and U7061 (N_7061,N_2533,N_3640);
and U7062 (N_7062,N_3203,N_4058);
and U7063 (N_7063,N_2555,N_4047);
and U7064 (N_7064,N_4346,N_3674);
and U7065 (N_7065,N_4043,N_3709);
nor U7066 (N_7066,N_3801,N_4071);
nand U7067 (N_7067,N_3868,N_3073);
or U7068 (N_7068,N_4938,N_4248);
nand U7069 (N_7069,N_2917,N_2843);
xnor U7070 (N_7070,N_3772,N_3045);
xor U7071 (N_7071,N_4857,N_3741);
xor U7072 (N_7072,N_3289,N_3668);
or U7073 (N_7073,N_4576,N_3124);
nor U7074 (N_7074,N_3478,N_4444);
nor U7075 (N_7075,N_4436,N_4939);
and U7076 (N_7076,N_2905,N_3991);
nor U7077 (N_7077,N_2872,N_3071);
and U7078 (N_7078,N_4845,N_4034);
nor U7079 (N_7079,N_3628,N_2940);
and U7080 (N_7080,N_3027,N_4742);
and U7081 (N_7081,N_2547,N_2864);
xnor U7082 (N_7082,N_2858,N_3587);
xor U7083 (N_7083,N_3873,N_3070);
nor U7084 (N_7084,N_2750,N_3878);
nand U7085 (N_7085,N_2549,N_3334);
xor U7086 (N_7086,N_4481,N_3932);
nor U7087 (N_7087,N_4424,N_3808);
or U7088 (N_7088,N_2562,N_3088);
xnor U7089 (N_7089,N_3785,N_3790);
nor U7090 (N_7090,N_2530,N_4966);
nand U7091 (N_7091,N_4712,N_4982);
nand U7092 (N_7092,N_4136,N_3262);
and U7093 (N_7093,N_4788,N_4092);
nor U7094 (N_7094,N_4571,N_4891);
nand U7095 (N_7095,N_3962,N_3135);
and U7096 (N_7096,N_3362,N_3621);
and U7097 (N_7097,N_4925,N_2595);
or U7098 (N_7098,N_4962,N_3587);
xnor U7099 (N_7099,N_4307,N_4300);
or U7100 (N_7100,N_4450,N_3231);
xnor U7101 (N_7101,N_4633,N_2658);
xnor U7102 (N_7102,N_3291,N_4304);
or U7103 (N_7103,N_4091,N_3006);
or U7104 (N_7104,N_3166,N_3738);
nand U7105 (N_7105,N_3347,N_3939);
nor U7106 (N_7106,N_3855,N_2742);
and U7107 (N_7107,N_4587,N_3076);
xor U7108 (N_7108,N_4764,N_3577);
nor U7109 (N_7109,N_3933,N_4735);
or U7110 (N_7110,N_4349,N_3151);
and U7111 (N_7111,N_3324,N_2574);
or U7112 (N_7112,N_3149,N_3703);
xnor U7113 (N_7113,N_2918,N_4332);
and U7114 (N_7114,N_3979,N_3728);
and U7115 (N_7115,N_2827,N_3137);
and U7116 (N_7116,N_3204,N_3062);
nor U7117 (N_7117,N_4903,N_4674);
nand U7118 (N_7118,N_3289,N_3454);
nor U7119 (N_7119,N_4421,N_2971);
or U7120 (N_7120,N_4444,N_3679);
nor U7121 (N_7121,N_3243,N_3860);
and U7122 (N_7122,N_3260,N_3865);
and U7123 (N_7123,N_4358,N_2843);
nor U7124 (N_7124,N_3782,N_4846);
nand U7125 (N_7125,N_4951,N_4868);
nor U7126 (N_7126,N_2893,N_2583);
or U7127 (N_7127,N_3591,N_2644);
xor U7128 (N_7128,N_3226,N_3024);
and U7129 (N_7129,N_4104,N_3305);
or U7130 (N_7130,N_3397,N_4108);
or U7131 (N_7131,N_4120,N_3682);
nand U7132 (N_7132,N_2993,N_4104);
or U7133 (N_7133,N_3830,N_4395);
nand U7134 (N_7134,N_3308,N_4030);
xor U7135 (N_7135,N_3834,N_4068);
nand U7136 (N_7136,N_3325,N_3096);
nand U7137 (N_7137,N_4230,N_4229);
nand U7138 (N_7138,N_3105,N_2690);
xnor U7139 (N_7139,N_4252,N_3599);
nand U7140 (N_7140,N_4522,N_4277);
or U7141 (N_7141,N_3622,N_3275);
nor U7142 (N_7142,N_4963,N_3805);
or U7143 (N_7143,N_3452,N_4395);
and U7144 (N_7144,N_3597,N_3523);
nand U7145 (N_7145,N_3593,N_4160);
and U7146 (N_7146,N_3596,N_3995);
or U7147 (N_7147,N_3379,N_4034);
xor U7148 (N_7148,N_3266,N_4068);
nand U7149 (N_7149,N_2886,N_2661);
nand U7150 (N_7150,N_4664,N_2834);
and U7151 (N_7151,N_3117,N_3650);
xor U7152 (N_7152,N_3605,N_4727);
xor U7153 (N_7153,N_4108,N_3521);
nand U7154 (N_7154,N_3723,N_3709);
xnor U7155 (N_7155,N_3114,N_3098);
xor U7156 (N_7156,N_3520,N_4924);
xnor U7157 (N_7157,N_4321,N_2582);
xor U7158 (N_7158,N_3179,N_3665);
or U7159 (N_7159,N_2765,N_3222);
nand U7160 (N_7160,N_4046,N_2732);
and U7161 (N_7161,N_3510,N_4653);
nor U7162 (N_7162,N_3426,N_3762);
nor U7163 (N_7163,N_3988,N_4847);
and U7164 (N_7164,N_4557,N_3398);
xnor U7165 (N_7165,N_2607,N_4914);
nand U7166 (N_7166,N_3629,N_4666);
xnor U7167 (N_7167,N_3606,N_2764);
nand U7168 (N_7168,N_4119,N_4211);
xor U7169 (N_7169,N_4293,N_3081);
or U7170 (N_7170,N_3681,N_3384);
nor U7171 (N_7171,N_3540,N_3444);
nor U7172 (N_7172,N_3362,N_3697);
and U7173 (N_7173,N_4827,N_3439);
nor U7174 (N_7174,N_4023,N_4861);
or U7175 (N_7175,N_3663,N_4136);
and U7176 (N_7176,N_4749,N_4682);
nor U7177 (N_7177,N_3720,N_4317);
nand U7178 (N_7178,N_4215,N_2673);
or U7179 (N_7179,N_2892,N_3968);
or U7180 (N_7180,N_4408,N_2915);
nor U7181 (N_7181,N_3461,N_4763);
and U7182 (N_7182,N_4030,N_4516);
nand U7183 (N_7183,N_3944,N_3122);
xnor U7184 (N_7184,N_2873,N_4779);
or U7185 (N_7185,N_3172,N_3191);
nor U7186 (N_7186,N_2913,N_2768);
or U7187 (N_7187,N_4899,N_2671);
and U7188 (N_7188,N_4653,N_3789);
xnor U7189 (N_7189,N_4437,N_3793);
nor U7190 (N_7190,N_4291,N_3429);
and U7191 (N_7191,N_3818,N_4570);
nor U7192 (N_7192,N_4922,N_2993);
or U7193 (N_7193,N_4229,N_3143);
nand U7194 (N_7194,N_3075,N_4774);
nand U7195 (N_7195,N_3924,N_3493);
nand U7196 (N_7196,N_4441,N_3662);
or U7197 (N_7197,N_3514,N_3613);
or U7198 (N_7198,N_3014,N_4046);
nand U7199 (N_7199,N_2690,N_4034);
nor U7200 (N_7200,N_4326,N_3789);
xnor U7201 (N_7201,N_3955,N_3747);
or U7202 (N_7202,N_4387,N_4840);
nand U7203 (N_7203,N_4218,N_2589);
nand U7204 (N_7204,N_4893,N_4649);
nand U7205 (N_7205,N_4069,N_2765);
or U7206 (N_7206,N_2534,N_4305);
nor U7207 (N_7207,N_2934,N_3100);
and U7208 (N_7208,N_2605,N_3877);
xnor U7209 (N_7209,N_2997,N_4522);
or U7210 (N_7210,N_4380,N_4664);
and U7211 (N_7211,N_3993,N_3451);
nand U7212 (N_7212,N_3599,N_3702);
nand U7213 (N_7213,N_3479,N_2665);
or U7214 (N_7214,N_2749,N_3403);
nor U7215 (N_7215,N_2943,N_3507);
xor U7216 (N_7216,N_4448,N_3302);
xnor U7217 (N_7217,N_4594,N_2895);
or U7218 (N_7218,N_3116,N_3536);
xor U7219 (N_7219,N_2737,N_2989);
and U7220 (N_7220,N_3816,N_4339);
or U7221 (N_7221,N_4471,N_3353);
xor U7222 (N_7222,N_3466,N_4220);
and U7223 (N_7223,N_3578,N_4644);
nand U7224 (N_7224,N_3016,N_2889);
or U7225 (N_7225,N_2753,N_3006);
or U7226 (N_7226,N_4857,N_2987);
or U7227 (N_7227,N_3950,N_3112);
nand U7228 (N_7228,N_3834,N_3568);
xor U7229 (N_7229,N_4070,N_4681);
nand U7230 (N_7230,N_4717,N_2801);
nor U7231 (N_7231,N_4175,N_3176);
nand U7232 (N_7232,N_4090,N_2890);
and U7233 (N_7233,N_4043,N_3895);
xnor U7234 (N_7234,N_3555,N_4490);
or U7235 (N_7235,N_4614,N_4240);
nor U7236 (N_7236,N_4704,N_4497);
or U7237 (N_7237,N_3210,N_3770);
nand U7238 (N_7238,N_4129,N_3521);
or U7239 (N_7239,N_3964,N_3958);
nor U7240 (N_7240,N_4355,N_3427);
nand U7241 (N_7241,N_4187,N_4638);
xor U7242 (N_7242,N_4157,N_4389);
or U7243 (N_7243,N_4981,N_4103);
and U7244 (N_7244,N_4557,N_3246);
nor U7245 (N_7245,N_3794,N_2622);
xnor U7246 (N_7246,N_2514,N_3603);
or U7247 (N_7247,N_3357,N_4439);
or U7248 (N_7248,N_3097,N_3318);
nand U7249 (N_7249,N_4316,N_4937);
nor U7250 (N_7250,N_4383,N_4904);
nor U7251 (N_7251,N_4310,N_4309);
and U7252 (N_7252,N_3943,N_3687);
nand U7253 (N_7253,N_3517,N_2638);
and U7254 (N_7254,N_4121,N_4162);
xor U7255 (N_7255,N_2651,N_4119);
nand U7256 (N_7256,N_2522,N_4001);
xnor U7257 (N_7257,N_4241,N_3109);
nor U7258 (N_7258,N_2612,N_2947);
or U7259 (N_7259,N_3223,N_4364);
nor U7260 (N_7260,N_2512,N_4007);
xor U7261 (N_7261,N_3139,N_4796);
nand U7262 (N_7262,N_4612,N_4956);
or U7263 (N_7263,N_3969,N_3497);
nand U7264 (N_7264,N_4199,N_4617);
nor U7265 (N_7265,N_2914,N_2971);
and U7266 (N_7266,N_4840,N_4242);
xnor U7267 (N_7267,N_3805,N_2971);
nor U7268 (N_7268,N_3862,N_3166);
nor U7269 (N_7269,N_2668,N_4972);
nand U7270 (N_7270,N_3791,N_4157);
or U7271 (N_7271,N_4537,N_4520);
xor U7272 (N_7272,N_4765,N_2699);
and U7273 (N_7273,N_4515,N_4154);
xor U7274 (N_7274,N_4624,N_3462);
nor U7275 (N_7275,N_2527,N_3628);
xor U7276 (N_7276,N_3436,N_3581);
nor U7277 (N_7277,N_4945,N_3901);
xnor U7278 (N_7278,N_4518,N_2954);
and U7279 (N_7279,N_4314,N_4614);
xnor U7280 (N_7280,N_4118,N_4861);
xnor U7281 (N_7281,N_4116,N_3342);
nand U7282 (N_7282,N_3631,N_4035);
and U7283 (N_7283,N_3584,N_3488);
and U7284 (N_7284,N_3498,N_4480);
or U7285 (N_7285,N_3652,N_4021);
or U7286 (N_7286,N_2865,N_4633);
xor U7287 (N_7287,N_2676,N_4647);
nor U7288 (N_7288,N_3860,N_3213);
nor U7289 (N_7289,N_3662,N_4841);
or U7290 (N_7290,N_4279,N_4953);
nand U7291 (N_7291,N_4114,N_4412);
nor U7292 (N_7292,N_2995,N_3293);
nor U7293 (N_7293,N_2539,N_3270);
xnor U7294 (N_7294,N_4008,N_2665);
xor U7295 (N_7295,N_3074,N_4525);
nand U7296 (N_7296,N_3269,N_4546);
nand U7297 (N_7297,N_4141,N_4745);
nor U7298 (N_7298,N_3993,N_3367);
and U7299 (N_7299,N_4608,N_3896);
nor U7300 (N_7300,N_3530,N_4117);
nor U7301 (N_7301,N_3574,N_3444);
nand U7302 (N_7302,N_2771,N_3761);
nand U7303 (N_7303,N_3146,N_4349);
nand U7304 (N_7304,N_2504,N_3358);
and U7305 (N_7305,N_3308,N_2834);
xor U7306 (N_7306,N_4039,N_2943);
and U7307 (N_7307,N_2951,N_3443);
nor U7308 (N_7308,N_2707,N_4870);
and U7309 (N_7309,N_4691,N_4125);
and U7310 (N_7310,N_3580,N_3646);
and U7311 (N_7311,N_3798,N_4807);
nand U7312 (N_7312,N_2888,N_3162);
or U7313 (N_7313,N_4654,N_4972);
nand U7314 (N_7314,N_3221,N_4480);
and U7315 (N_7315,N_3151,N_4482);
nor U7316 (N_7316,N_4742,N_4198);
nand U7317 (N_7317,N_3561,N_3712);
or U7318 (N_7318,N_4682,N_3655);
or U7319 (N_7319,N_2554,N_2539);
or U7320 (N_7320,N_4990,N_4905);
xnor U7321 (N_7321,N_2861,N_2922);
nand U7322 (N_7322,N_4885,N_4486);
nor U7323 (N_7323,N_4544,N_3380);
nor U7324 (N_7324,N_4502,N_2871);
or U7325 (N_7325,N_2861,N_2663);
xor U7326 (N_7326,N_3269,N_3790);
xnor U7327 (N_7327,N_2578,N_4767);
xor U7328 (N_7328,N_4325,N_4892);
nand U7329 (N_7329,N_4672,N_4015);
xor U7330 (N_7330,N_3222,N_2518);
xnor U7331 (N_7331,N_2862,N_3254);
xnor U7332 (N_7332,N_4440,N_4083);
nor U7333 (N_7333,N_4894,N_4873);
xor U7334 (N_7334,N_3546,N_2574);
xnor U7335 (N_7335,N_3496,N_3509);
nor U7336 (N_7336,N_4309,N_2628);
or U7337 (N_7337,N_4895,N_3109);
or U7338 (N_7338,N_3791,N_4653);
and U7339 (N_7339,N_2556,N_3726);
or U7340 (N_7340,N_2557,N_2681);
nand U7341 (N_7341,N_3515,N_4455);
and U7342 (N_7342,N_4739,N_4612);
nor U7343 (N_7343,N_4462,N_2569);
nand U7344 (N_7344,N_2797,N_4453);
nand U7345 (N_7345,N_2838,N_3881);
or U7346 (N_7346,N_2826,N_4292);
and U7347 (N_7347,N_3842,N_4341);
nand U7348 (N_7348,N_2606,N_2560);
or U7349 (N_7349,N_3160,N_2519);
or U7350 (N_7350,N_3957,N_4451);
and U7351 (N_7351,N_3114,N_4224);
xor U7352 (N_7352,N_4697,N_4006);
nand U7353 (N_7353,N_3157,N_4688);
nand U7354 (N_7354,N_2821,N_2766);
nor U7355 (N_7355,N_3927,N_3585);
or U7356 (N_7356,N_3000,N_4215);
or U7357 (N_7357,N_3691,N_4490);
nor U7358 (N_7358,N_3377,N_3203);
nand U7359 (N_7359,N_2872,N_3362);
nand U7360 (N_7360,N_2759,N_4165);
nand U7361 (N_7361,N_2810,N_2604);
and U7362 (N_7362,N_3195,N_3716);
nor U7363 (N_7363,N_3387,N_4523);
xor U7364 (N_7364,N_4929,N_2644);
and U7365 (N_7365,N_4069,N_4731);
or U7366 (N_7366,N_3252,N_3815);
xnor U7367 (N_7367,N_3059,N_4010);
xor U7368 (N_7368,N_3117,N_4027);
nor U7369 (N_7369,N_3314,N_4957);
or U7370 (N_7370,N_4205,N_4624);
or U7371 (N_7371,N_4604,N_3443);
and U7372 (N_7372,N_2529,N_4512);
and U7373 (N_7373,N_4517,N_2958);
nand U7374 (N_7374,N_3913,N_2649);
and U7375 (N_7375,N_2978,N_4360);
and U7376 (N_7376,N_4756,N_2691);
or U7377 (N_7377,N_3310,N_4610);
and U7378 (N_7378,N_2536,N_3206);
nor U7379 (N_7379,N_4380,N_4551);
and U7380 (N_7380,N_3624,N_3780);
or U7381 (N_7381,N_4589,N_3930);
xor U7382 (N_7382,N_3766,N_2702);
nor U7383 (N_7383,N_4040,N_3450);
nor U7384 (N_7384,N_2987,N_2535);
xnor U7385 (N_7385,N_3593,N_4268);
or U7386 (N_7386,N_3859,N_3466);
and U7387 (N_7387,N_4464,N_3582);
nand U7388 (N_7388,N_3705,N_3794);
nor U7389 (N_7389,N_2865,N_3102);
xnor U7390 (N_7390,N_4918,N_3444);
nand U7391 (N_7391,N_3336,N_3504);
and U7392 (N_7392,N_2702,N_4636);
xnor U7393 (N_7393,N_3094,N_3496);
or U7394 (N_7394,N_4028,N_3051);
nand U7395 (N_7395,N_3280,N_3660);
nor U7396 (N_7396,N_3401,N_4768);
and U7397 (N_7397,N_4726,N_2958);
or U7398 (N_7398,N_3311,N_3257);
or U7399 (N_7399,N_4648,N_3967);
nand U7400 (N_7400,N_3510,N_4189);
and U7401 (N_7401,N_2775,N_4845);
xor U7402 (N_7402,N_4695,N_4319);
xnor U7403 (N_7403,N_3830,N_2916);
or U7404 (N_7404,N_4669,N_4752);
nand U7405 (N_7405,N_3998,N_3739);
nand U7406 (N_7406,N_4425,N_3290);
and U7407 (N_7407,N_3799,N_3744);
xor U7408 (N_7408,N_3751,N_3736);
and U7409 (N_7409,N_4557,N_4751);
nand U7410 (N_7410,N_4915,N_4866);
nor U7411 (N_7411,N_4218,N_4340);
nor U7412 (N_7412,N_4737,N_3590);
or U7413 (N_7413,N_3077,N_3784);
nor U7414 (N_7414,N_4854,N_2744);
and U7415 (N_7415,N_3292,N_2508);
or U7416 (N_7416,N_4088,N_3084);
or U7417 (N_7417,N_3082,N_4624);
and U7418 (N_7418,N_3271,N_4660);
and U7419 (N_7419,N_3455,N_4333);
or U7420 (N_7420,N_4406,N_2743);
xnor U7421 (N_7421,N_4496,N_3645);
nor U7422 (N_7422,N_4821,N_4337);
xor U7423 (N_7423,N_3825,N_3587);
or U7424 (N_7424,N_2971,N_4583);
or U7425 (N_7425,N_3014,N_3843);
xnor U7426 (N_7426,N_2539,N_4083);
and U7427 (N_7427,N_4453,N_4058);
and U7428 (N_7428,N_3562,N_3402);
nand U7429 (N_7429,N_4583,N_3899);
nand U7430 (N_7430,N_4769,N_4557);
xor U7431 (N_7431,N_4732,N_3201);
xnor U7432 (N_7432,N_4086,N_3405);
and U7433 (N_7433,N_3101,N_4915);
xnor U7434 (N_7434,N_4213,N_3583);
nor U7435 (N_7435,N_4518,N_3438);
nor U7436 (N_7436,N_4175,N_4517);
nand U7437 (N_7437,N_4520,N_4599);
xnor U7438 (N_7438,N_3689,N_4938);
xnor U7439 (N_7439,N_2698,N_3589);
or U7440 (N_7440,N_2818,N_3290);
nand U7441 (N_7441,N_3444,N_3722);
nor U7442 (N_7442,N_4713,N_4412);
xnor U7443 (N_7443,N_4958,N_4313);
nor U7444 (N_7444,N_3604,N_4087);
xor U7445 (N_7445,N_4899,N_3534);
or U7446 (N_7446,N_2684,N_3713);
xnor U7447 (N_7447,N_4284,N_4937);
or U7448 (N_7448,N_3868,N_4695);
and U7449 (N_7449,N_2974,N_2760);
and U7450 (N_7450,N_4557,N_3276);
xnor U7451 (N_7451,N_3997,N_4454);
xnor U7452 (N_7452,N_2664,N_3935);
or U7453 (N_7453,N_3421,N_3484);
nor U7454 (N_7454,N_4441,N_3141);
xnor U7455 (N_7455,N_4232,N_4119);
or U7456 (N_7456,N_2932,N_4949);
nand U7457 (N_7457,N_4601,N_3336);
xnor U7458 (N_7458,N_4063,N_4279);
or U7459 (N_7459,N_3168,N_3218);
and U7460 (N_7460,N_2679,N_4599);
nand U7461 (N_7461,N_3417,N_3409);
nor U7462 (N_7462,N_2656,N_4811);
and U7463 (N_7463,N_3851,N_4140);
xnor U7464 (N_7464,N_3137,N_2875);
nand U7465 (N_7465,N_3799,N_3911);
or U7466 (N_7466,N_3311,N_2913);
xor U7467 (N_7467,N_3078,N_3380);
and U7468 (N_7468,N_4488,N_4804);
nor U7469 (N_7469,N_3401,N_3805);
xor U7470 (N_7470,N_3919,N_3022);
xnor U7471 (N_7471,N_3376,N_3333);
or U7472 (N_7472,N_4451,N_4649);
and U7473 (N_7473,N_3961,N_3651);
or U7474 (N_7474,N_4316,N_4769);
and U7475 (N_7475,N_4384,N_3698);
nand U7476 (N_7476,N_3128,N_2681);
or U7477 (N_7477,N_3581,N_4463);
and U7478 (N_7478,N_3257,N_2961);
and U7479 (N_7479,N_4702,N_2687);
or U7480 (N_7480,N_3162,N_2533);
nor U7481 (N_7481,N_3549,N_2752);
nor U7482 (N_7482,N_3703,N_4789);
xnor U7483 (N_7483,N_3910,N_4284);
nor U7484 (N_7484,N_3933,N_4178);
nor U7485 (N_7485,N_2631,N_3802);
nor U7486 (N_7486,N_3922,N_2594);
or U7487 (N_7487,N_3264,N_2651);
nand U7488 (N_7488,N_3653,N_3804);
and U7489 (N_7489,N_3415,N_2615);
nor U7490 (N_7490,N_3375,N_4707);
nand U7491 (N_7491,N_3370,N_3540);
or U7492 (N_7492,N_3248,N_3673);
nor U7493 (N_7493,N_3856,N_2788);
xnor U7494 (N_7494,N_2532,N_2716);
nand U7495 (N_7495,N_4571,N_4220);
nor U7496 (N_7496,N_3732,N_2522);
and U7497 (N_7497,N_2770,N_4070);
nor U7498 (N_7498,N_3082,N_2784);
nor U7499 (N_7499,N_4936,N_3791);
or U7500 (N_7500,N_6963,N_5889);
nor U7501 (N_7501,N_7346,N_5490);
nand U7502 (N_7502,N_7050,N_6482);
nor U7503 (N_7503,N_6329,N_6349);
or U7504 (N_7504,N_6340,N_5437);
nand U7505 (N_7505,N_5439,N_6268);
xor U7506 (N_7506,N_6111,N_7147);
nor U7507 (N_7507,N_6899,N_5545);
and U7508 (N_7508,N_5680,N_6562);
nor U7509 (N_7509,N_7066,N_5152);
and U7510 (N_7510,N_7159,N_5890);
nand U7511 (N_7511,N_7443,N_7136);
and U7512 (N_7512,N_5268,N_5223);
and U7513 (N_7513,N_6447,N_5238);
nor U7514 (N_7514,N_7177,N_5380);
xnor U7515 (N_7515,N_6394,N_6816);
xor U7516 (N_7516,N_7111,N_6998);
nand U7517 (N_7517,N_5556,N_6885);
xnor U7518 (N_7518,N_7377,N_6121);
nor U7519 (N_7519,N_7055,N_6265);
nand U7520 (N_7520,N_7202,N_7208);
nor U7521 (N_7521,N_7024,N_7408);
and U7522 (N_7522,N_6664,N_7426);
or U7523 (N_7523,N_6529,N_5245);
and U7524 (N_7524,N_5704,N_6148);
nand U7525 (N_7525,N_5633,N_5289);
nor U7526 (N_7526,N_5730,N_6160);
or U7527 (N_7527,N_6947,N_5685);
or U7528 (N_7528,N_6218,N_5902);
xor U7529 (N_7529,N_5322,N_6175);
and U7530 (N_7530,N_6569,N_7071);
nor U7531 (N_7531,N_7458,N_5251);
nor U7532 (N_7532,N_7387,N_7382);
and U7533 (N_7533,N_6366,N_5084);
xnor U7534 (N_7534,N_6464,N_6993);
and U7535 (N_7535,N_7467,N_6927);
xnor U7536 (N_7536,N_7252,N_6603);
or U7537 (N_7537,N_6370,N_5495);
and U7538 (N_7538,N_6581,N_6258);
and U7539 (N_7539,N_5724,N_6708);
xor U7540 (N_7540,N_6656,N_7432);
nor U7541 (N_7541,N_5412,N_6991);
nand U7542 (N_7542,N_7155,N_5977);
nand U7543 (N_7543,N_7306,N_6004);
nor U7544 (N_7544,N_5781,N_5079);
nand U7545 (N_7545,N_6086,N_5710);
nand U7546 (N_7546,N_6235,N_5608);
or U7547 (N_7547,N_5331,N_6772);
nor U7548 (N_7548,N_6929,N_7180);
xor U7549 (N_7549,N_7279,N_5513);
nor U7550 (N_7550,N_6161,N_5302);
nor U7551 (N_7551,N_5837,N_5930);
nor U7552 (N_7552,N_7470,N_6645);
xnor U7553 (N_7553,N_5792,N_6653);
xnor U7554 (N_7554,N_5498,N_6026);
nand U7555 (N_7555,N_6870,N_7120);
and U7556 (N_7556,N_5903,N_5611);
and U7557 (N_7557,N_5367,N_5709);
and U7558 (N_7558,N_6391,N_5448);
or U7559 (N_7559,N_6251,N_6986);
and U7560 (N_7560,N_7313,N_5594);
and U7561 (N_7561,N_6295,N_6304);
xor U7562 (N_7562,N_6669,N_5697);
nor U7563 (N_7563,N_7474,N_7295);
or U7564 (N_7564,N_6844,N_6262);
nor U7565 (N_7565,N_6321,N_6454);
nor U7566 (N_7566,N_7182,N_5879);
nor U7567 (N_7567,N_6410,N_6977);
nor U7568 (N_7568,N_5241,N_6889);
nor U7569 (N_7569,N_6956,N_5688);
or U7570 (N_7570,N_6650,N_5215);
nand U7571 (N_7571,N_5395,N_6017);
nand U7572 (N_7572,N_6516,N_5392);
or U7573 (N_7573,N_7047,N_7199);
xor U7574 (N_7574,N_5012,N_6784);
and U7575 (N_7575,N_6663,N_7283);
xnor U7576 (N_7576,N_7016,N_6078);
nor U7577 (N_7577,N_5428,N_5122);
or U7578 (N_7578,N_5993,N_5404);
nand U7579 (N_7579,N_6139,N_5487);
xor U7580 (N_7580,N_5727,N_5725);
nand U7581 (N_7581,N_7378,N_6876);
and U7582 (N_7582,N_5071,N_5209);
or U7583 (N_7583,N_6856,N_6584);
and U7584 (N_7584,N_5884,N_6032);
or U7585 (N_7585,N_7434,N_6125);
and U7586 (N_7586,N_7475,N_6101);
nand U7587 (N_7587,N_7076,N_6085);
nand U7588 (N_7588,N_6731,N_6705);
nand U7589 (N_7589,N_7414,N_6848);
or U7590 (N_7590,N_7300,N_6310);
nor U7591 (N_7591,N_5098,N_6021);
and U7592 (N_7592,N_5352,N_6460);
or U7593 (N_7593,N_5329,N_6932);
or U7594 (N_7594,N_6071,N_5198);
xnor U7595 (N_7595,N_6113,N_6577);
and U7596 (N_7596,N_7369,N_5693);
xor U7597 (N_7597,N_7341,N_6944);
xnor U7598 (N_7598,N_5869,N_6594);
xnor U7599 (N_7599,N_5908,N_5808);
or U7600 (N_7600,N_6002,N_5916);
nand U7601 (N_7601,N_5783,N_5973);
nor U7602 (N_7602,N_6419,N_7082);
xnor U7603 (N_7603,N_5178,N_5876);
nor U7604 (N_7604,N_7130,N_6589);
nand U7605 (N_7605,N_7026,N_6165);
nor U7606 (N_7606,N_7203,N_6520);
nor U7607 (N_7607,N_5267,N_6171);
xnor U7608 (N_7608,N_6005,N_7256);
nand U7609 (N_7609,N_6193,N_6623);
or U7610 (N_7610,N_7342,N_5381);
nor U7611 (N_7611,N_6392,N_6754);
nor U7612 (N_7612,N_7222,N_6335);
or U7613 (N_7613,N_6771,N_7035);
and U7614 (N_7614,N_6999,N_6324);
or U7615 (N_7615,N_6477,N_5682);
and U7616 (N_7616,N_5488,N_6903);
and U7617 (N_7617,N_5151,N_6363);
nor U7618 (N_7618,N_5140,N_7077);
xor U7619 (N_7619,N_6158,N_6008);
and U7620 (N_7620,N_5541,N_7109);
or U7621 (N_7621,N_5828,N_7296);
or U7622 (N_7622,N_5833,N_5628);
and U7623 (N_7623,N_7193,N_6990);
nor U7624 (N_7624,N_5192,N_5443);
and U7625 (N_7625,N_6415,N_6895);
nor U7626 (N_7626,N_6658,N_5265);
nand U7627 (N_7627,N_6475,N_5899);
xor U7628 (N_7628,N_5044,N_5176);
xnor U7629 (N_7629,N_7488,N_7008);
nor U7630 (N_7630,N_7268,N_7194);
or U7631 (N_7631,N_7463,N_6197);
or U7632 (N_7632,N_5831,N_5575);
and U7633 (N_7633,N_5610,N_6434);
or U7634 (N_7634,N_6812,N_6504);
xnor U7635 (N_7635,N_6127,N_7438);
nand U7636 (N_7636,N_6961,N_5957);
and U7637 (N_7637,N_7116,N_5982);
xor U7638 (N_7638,N_5738,N_5306);
nor U7639 (N_7639,N_5967,N_5637);
or U7640 (N_7640,N_5978,N_5410);
nor U7641 (N_7641,N_6323,N_5130);
and U7642 (N_7642,N_5764,N_7200);
nor U7643 (N_7643,N_5384,N_6906);
nand U7644 (N_7644,N_5021,N_7015);
nand U7645 (N_7645,N_7046,N_6893);
and U7646 (N_7646,N_7166,N_5801);
and U7647 (N_7647,N_6887,N_5600);
nand U7648 (N_7648,N_6972,N_6431);
and U7649 (N_7649,N_6588,N_5868);
xor U7650 (N_7650,N_5980,N_6219);
and U7651 (N_7651,N_7479,N_7105);
xor U7652 (N_7652,N_5444,N_5548);
or U7653 (N_7653,N_5325,N_6718);
or U7654 (N_7654,N_6845,N_7053);
nor U7655 (N_7655,N_7437,N_5963);
nor U7656 (N_7656,N_6606,N_6390);
xnor U7657 (N_7657,N_5171,N_6354);
nor U7658 (N_7658,N_6747,N_7093);
or U7659 (N_7659,N_5670,N_6888);
and U7660 (N_7660,N_6337,N_7362);
nand U7661 (N_7661,N_5460,N_5749);
or U7662 (N_7662,N_6621,N_6339);
nor U7663 (N_7663,N_5970,N_5737);
nor U7664 (N_7664,N_6808,N_5587);
or U7665 (N_7665,N_5403,N_6300);
nand U7666 (N_7666,N_6980,N_6683);
xor U7667 (N_7667,N_6328,N_6609);
or U7668 (N_7668,N_5865,N_6655);
xor U7669 (N_7669,N_6692,N_6401);
and U7670 (N_7670,N_6847,N_7406);
and U7671 (N_7671,N_5974,N_5270);
or U7672 (N_7672,N_5374,N_5386);
xnor U7673 (N_7673,N_5298,N_5851);
and U7674 (N_7674,N_6874,N_5585);
nor U7675 (N_7675,N_7392,N_5421);
xnor U7676 (N_7676,N_6369,N_5187);
or U7677 (N_7677,N_6863,N_6676);
xor U7678 (N_7678,N_5701,N_6129);
xnor U7679 (N_7679,N_7397,N_6629);
nor U7680 (N_7680,N_5888,N_7267);
nand U7681 (N_7681,N_5128,N_6221);
xor U7682 (N_7682,N_7269,N_5845);
or U7683 (N_7683,N_6615,N_5093);
nor U7684 (N_7684,N_7049,N_6319);
or U7685 (N_7685,N_7302,N_6740);
nor U7686 (N_7686,N_6823,N_5305);
nand U7687 (N_7687,N_5842,N_5641);
nand U7688 (N_7688,N_5220,N_5489);
or U7689 (N_7689,N_6924,N_7245);
nand U7690 (N_7690,N_6413,N_6398);
or U7691 (N_7691,N_6247,N_5172);
and U7692 (N_7692,N_6459,N_5847);
nor U7693 (N_7693,N_7454,N_5820);
and U7694 (N_7694,N_6696,N_5167);
or U7695 (N_7695,N_5160,N_6546);
nor U7696 (N_7696,N_6048,N_5123);
or U7697 (N_7697,N_5986,N_5274);
or U7698 (N_7698,N_5043,N_5962);
xnor U7699 (N_7699,N_5365,N_6060);
or U7700 (N_7700,N_7061,N_6837);
and U7701 (N_7701,N_7373,N_6836);
xor U7702 (N_7702,N_5371,N_5087);
nand U7703 (N_7703,N_6439,N_6182);
or U7704 (N_7704,N_7229,N_5006);
nand U7705 (N_7705,N_6450,N_5583);
and U7706 (N_7706,N_5001,N_7052);
xnor U7707 (N_7707,N_6662,N_5227);
xnor U7708 (N_7708,N_6470,N_6979);
and U7709 (N_7709,N_6719,N_5330);
xor U7710 (N_7710,N_7103,N_7175);
nand U7711 (N_7711,N_6850,N_7368);
or U7712 (N_7712,N_5987,N_7181);
or U7713 (N_7713,N_5214,N_6519);
nand U7714 (N_7714,N_5674,N_7223);
and U7715 (N_7715,N_6442,N_5399);
or U7716 (N_7716,N_6451,N_6496);
nor U7717 (N_7717,N_7080,N_5275);
nand U7718 (N_7718,N_7030,N_6612);
or U7719 (N_7719,N_7335,N_6178);
xor U7720 (N_7720,N_5625,N_6509);
and U7721 (N_7721,N_5651,N_6809);
and U7722 (N_7722,N_6495,N_5383);
or U7723 (N_7723,N_5387,N_6146);
xnor U7724 (N_7724,N_7044,N_7259);
nand U7725 (N_7725,N_6087,N_5033);
nor U7726 (N_7726,N_5683,N_6671);
xor U7727 (N_7727,N_6526,N_5148);
nor U7728 (N_7728,N_6695,N_6521);
nand U7729 (N_7729,N_6025,N_7492);
or U7730 (N_7730,N_6560,N_5508);
xor U7731 (N_7731,N_5811,N_5592);
and U7732 (N_7732,N_5005,N_5185);
and U7733 (N_7733,N_5059,N_5994);
nor U7734 (N_7734,N_6643,N_7249);
nand U7735 (N_7735,N_5332,N_6834);
or U7736 (N_7736,N_5702,N_6079);
xnor U7737 (N_7737,N_6040,N_7151);
xnor U7738 (N_7738,N_5959,N_6810);
xnor U7739 (N_7739,N_6617,N_6780);
nor U7740 (N_7740,N_5664,N_6648);
or U7741 (N_7741,N_6142,N_7452);
nor U7742 (N_7742,N_7243,N_7304);
nor U7743 (N_7743,N_5037,N_6232);
and U7744 (N_7744,N_5003,N_6039);
or U7745 (N_7745,N_6535,N_5173);
and U7746 (N_7746,N_7083,N_5455);
nand U7747 (N_7747,N_7308,N_5264);
nand U7748 (N_7748,N_7402,N_7340);
xor U7749 (N_7749,N_6992,N_7025);
and U7750 (N_7750,N_6367,N_6128);
or U7751 (N_7751,N_5008,N_7237);
nand U7752 (N_7752,N_6839,N_5112);
nand U7753 (N_7753,N_5675,N_6371);
nand U7754 (N_7754,N_6649,N_6841);
or U7755 (N_7755,N_5396,N_5233);
and U7756 (N_7756,N_6877,N_5613);
xnor U7757 (N_7757,N_6498,N_7000);
or U7758 (N_7758,N_5124,N_5434);
nor U7759 (N_7759,N_5925,N_7228);
nor U7760 (N_7760,N_6170,N_6982);
or U7761 (N_7761,N_5166,N_5789);
xor U7762 (N_7762,N_7446,N_5110);
xor U7763 (N_7763,N_5426,N_5321);
and U7764 (N_7764,N_6095,N_7090);
xnor U7765 (N_7765,N_6716,N_6420);
xnor U7766 (N_7766,N_6252,N_6514);
xnor U7767 (N_7767,N_5424,N_6965);
xor U7768 (N_7768,N_6618,N_5142);
nand U7769 (N_7769,N_6666,N_5323);
or U7770 (N_7770,N_6717,N_5234);
and U7771 (N_7771,N_5626,N_5662);
nand U7772 (N_7772,N_6897,N_5663);
nand U7773 (N_7773,N_7301,N_6978);
or U7774 (N_7774,N_6124,N_5972);
or U7775 (N_7775,N_5866,N_6236);
xor U7776 (N_7776,N_5870,N_7032);
nand U7777 (N_7777,N_6345,N_7466);
nor U7778 (N_7778,N_6802,N_6417);
nor U7779 (N_7779,N_5644,N_5077);
xor U7780 (N_7780,N_5984,N_6657);
xor U7781 (N_7781,N_7419,N_5307);
xnor U7782 (N_7782,N_5753,N_7084);
nor U7783 (N_7783,N_5537,N_6134);
xor U7784 (N_7784,N_6901,N_6303);
and U7785 (N_7785,N_5373,N_6455);
or U7786 (N_7786,N_5825,N_6852);
xor U7787 (N_7787,N_5589,N_7435);
and U7788 (N_7788,N_5024,N_5327);
nor U7789 (N_7789,N_6123,N_5956);
xor U7790 (N_7790,N_5258,N_6619);
nand U7791 (N_7791,N_7043,N_6380);
nand U7792 (N_7792,N_6920,N_6973);
and U7793 (N_7793,N_5824,N_7086);
or U7794 (N_7794,N_5207,N_5486);
xnor U7795 (N_7795,N_6082,N_6385);
nand U7796 (N_7796,N_5765,N_6725);
nor U7797 (N_7797,N_5072,N_5518);
or U7798 (N_7798,N_5741,N_7323);
xnor U7799 (N_7799,N_6800,N_5914);
xnor U7800 (N_7800,N_5108,N_6548);
or U7801 (N_7801,N_7439,N_5939);
and U7802 (N_7802,N_7074,N_6285);
nor U7803 (N_7803,N_5841,N_5791);
or U7804 (N_7804,N_5131,N_6566);
or U7805 (N_7805,N_6141,N_7487);
or U7806 (N_7806,N_7298,N_7126);
nor U7807 (N_7807,N_7135,N_6234);
or U7808 (N_7808,N_6189,N_7004);
or U7809 (N_7809,N_7211,N_5347);
or U7810 (N_7810,N_6365,N_7178);
or U7811 (N_7811,N_6216,N_6813);
xnor U7812 (N_7812,N_7113,N_5189);
nand U7813 (N_7813,N_6625,N_6274);
and U7814 (N_7814,N_6883,N_5926);
xor U7815 (N_7815,N_7236,N_7484);
xor U7816 (N_7816,N_6690,N_5068);
nand U7817 (N_7817,N_7089,N_7002);
nor U7818 (N_7818,N_6376,N_6631);
nand U7819 (N_7819,N_6827,N_5966);
xor U7820 (N_7820,N_5375,N_5253);
nor U7821 (N_7821,N_7210,N_5810);
and U7822 (N_7822,N_7418,N_7065);
or U7823 (N_7823,N_7101,N_6188);
xnor U7824 (N_7824,N_5767,N_6254);
xor U7825 (N_7825,N_7413,N_6037);
nor U7826 (N_7826,N_5062,N_6389);
and U7827 (N_7827,N_7311,N_5905);
nand U7828 (N_7828,N_5063,N_7363);
nand U7829 (N_7829,N_7185,N_7213);
nor U7830 (N_7830,N_5555,N_7179);
nor U7831 (N_7831,N_5565,N_5768);
xnor U7832 (N_7832,N_6547,N_6787);
or U7833 (N_7833,N_5948,N_5419);
xnor U7834 (N_7834,N_5221,N_7230);
or U7835 (N_7835,N_5504,N_6361);
xnor U7836 (N_7836,N_7345,N_5423);
nand U7837 (N_7837,N_6730,N_6144);
xnor U7838 (N_7838,N_6091,N_7013);
nand U7839 (N_7839,N_7227,N_6374);
nand U7840 (N_7840,N_5362,N_5576);
xnor U7841 (N_7841,N_5304,N_7144);
and U7842 (N_7842,N_6033,N_5127);
and U7843 (N_7843,N_5679,N_5017);
nand U7844 (N_7844,N_6412,N_6151);
nor U7845 (N_7845,N_5822,N_6478);
xnor U7846 (N_7846,N_6660,N_6767);
nand U7847 (N_7847,N_7410,N_7100);
nand U7848 (N_7848,N_7197,N_7070);
or U7849 (N_7849,N_7483,N_6159);
or U7850 (N_7850,N_5244,N_7033);
xor U7851 (N_7851,N_6733,N_6120);
xnor U7852 (N_7852,N_5468,N_6407);
and U7853 (N_7853,N_5479,N_6036);
xnor U7854 (N_7854,N_6131,N_5475);
nor U7855 (N_7855,N_7158,N_5200);
or U7856 (N_7856,N_6953,N_5678);
nor U7857 (N_7857,N_6900,N_5429);
and U7858 (N_7858,N_5402,N_7085);
nor U7859 (N_7859,N_5250,N_6396);
xnor U7860 (N_7860,N_6034,N_5883);
or U7861 (N_7861,N_6777,N_7293);
and U7862 (N_7862,N_5010,N_5642);
nor U7863 (N_7863,N_5070,N_6822);
xnor U7864 (N_7864,N_5053,N_7314);
and U7865 (N_7865,N_5619,N_5609);
and U7866 (N_7866,N_5717,N_5687);
and U7867 (N_7867,N_6923,N_5105);
nand U7868 (N_7868,N_6425,N_5928);
or U7869 (N_7869,N_5955,N_6106);
nand U7870 (N_7870,N_5909,N_6473);
or U7871 (N_7871,N_6568,N_5534);
nand U7872 (N_7872,N_6818,N_5850);
and U7873 (N_7873,N_5635,N_5170);
nand U7874 (N_7874,N_5586,N_7328);
or U7875 (N_7875,N_7472,N_5296);
nor U7876 (N_7876,N_6281,N_5547);
nand U7877 (N_7877,N_5368,N_6987);
and U7878 (N_7878,N_6534,N_5470);
xnor U7879 (N_7879,N_5137,N_7272);
nand U7880 (N_7880,N_6443,N_6208);
nand U7881 (N_7881,N_5927,N_7031);
xor U7882 (N_7882,N_6769,N_5536);
or U7883 (N_7883,N_6384,N_5469);
xor U7884 (N_7884,N_6640,N_6186);
or U7885 (N_7885,N_5111,N_5535);
and U7886 (N_7886,N_5595,N_7481);
nand U7887 (N_7887,N_6075,N_6513);
nor U7888 (N_7888,N_6860,N_7195);
nor U7889 (N_7889,N_5356,N_6076);
nor U7890 (N_7890,N_5100,N_5540);
and U7891 (N_7891,N_7491,N_6344);
nand U7892 (N_7892,N_6287,N_6312);
xor U7893 (N_7893,N_6405,N_5665);
xor U7894 (N_7894,N_7358,N_5848);
and U7895 (N_7895,N_6068,N_5333);
nand U7896 (N_7896,N_6273,N_7097);
xor U7897 (N_7897,N_5653,N_6143);
nor U7898 (N_7898,N_5278,N_6253);
nand U7899 (N_7899,N_5853,N_6018);
or U7900 (N_7900,N_6884,N_7292);
xnor U7901 (N_7901,N_6156,N_7427);
xnor U7902 (N_7902,N_7352,N_6064);
or U7903 (N_7903,N_7216,N_6421);
nand U7904 (N_7904,N_6222,N_7020);
or U7905 (N_7905,N_7133,N_7198);
or U7906 (N_7906,N_5856,N_5559);
xor U7907 (N_7907,N_7496,N_5466);
xnor U7908 (N_7908,N_6647,N_5666);
xnor U7909 (N_7909,N_6342,N_7495);
and U7910 (N_7910,N_6430,N_6047);
or U7911 (N_7911,N_6796,N_5722);
nor U7912 (N_7912,N_5398,N_5568);
xnor U7913 (N_7913,N_5237,N_5126);
nand U7914 (N_7914,N_5211,N_6402);
xnor U7915 (N_7915,N_6579,N_6684);
nand U7916 (N_7916,N_6493,N_6084);
nor U7917 (N_7917,N_5300,N_7416);
nor U7918 (N_7918,N_5188,N_6433);
xnor U7919 (N_7919,N_7280,N_6333);
and U7920 (N_7920,N_6819,N_6622);
or U7921 (N_7921,N_6766,N_7164);
nor U7922 (N_7922,N_5210,N_5430);
or U7923 (N_7923,N_6092,N_6437);
nor U7924 (N_7924,N_7478,N_5953);
xnor U7925 (N_7925,N_7232,N_6824);
and U7926 (N_7926,N_6867,N_5569);
nand U7927 (N_7927,N_7367,N_7212);
and U7928 (N_7928,N_6515,N_5389);
nor U7929 (N_7929,N_5938,N_6061);
nor U7930 (N_7930,N_6561,N_5219);
xnor U7931 (N_7931,N_5511,N_6072);
nand U7932 (N_7932,N_6379,N_7398);
nor U7933 (N_7933,N_6729,N_6373);
or U7934 (N_7934,N_5951,N_7457);
nand U7935 (N_7935,N_6712,N_6317);
nand U7936 (N_7936,N_6706,N_6697);
nor U7937 (N_7937,N_6331,N_5671);
and U7938 (N_7938,N_7238,N_5415);
or U7939 (N_7939,N_7054,N_6104);
or U7940 (N_7940,N_5983,N_7494);
xnor U7941 (N_7941,N_6549,N_7121);
nor U7942 (N_7942,N_5136,N_7117);
nor U7943 (N_7943,N_7285,N_6489);
xnor U7944 (N_7944,N_5648,N_6267);
nor U7945 (N_7945,N_5055,N_5880);
nor U7946 (N_7946,N_5533,N_6890);
nor U7947 (N_7947,N_5996,N_7465);
or U7948 (N_7948,N_6926,N_5164);
and U7949 (N_7949,N_6461,N_6330);
and U7950 (N_7950,N_6630,N_6913);
nor U7951 (N_7951,N_6116,N_7220);
nand U7952 (N_7952,N_6423,N_6593);
and U7953 (N_7953,N_6613,N_6908);
nand U7954 (N_7954,N_5472,N_6830);
nor U7955 (N_7955,N_7331,N_5580);
nand U7956 (N_7956,N_6959,N_7493);
xnor U7957 (N_7957,N_6751,N_7365);
nor U7958 (N_7958,N_5999,N_5638);
nand U7959 (N_7959,N_6152,N_6550);
or U7960 (N_7960,N_6567,N_5769);
xor U7961 (N_7961,N_6167,N_7123);
and U7962 (N_7962,N_6756,N_6030);
or U7963 (N_7963,N_6934,N_6907);
xnor U7964 (N_7964,N_5558,N_5370);
or U7965 (N_7965,N_7273,N_6642);
nand U7966 (N_7966,N_7260,N_7343);
or U7967 (N_7967,N_7183,N_5520);
nor U7968 (N_7968,N_6203,N_6735);
xnor U7969 (N_7969,N_7442,N_6743);
or U7970 (N_7970,N_5803,N_7330);
xnor U7971 (N_7971,N_5525,N_6024);
xnor U7972 (N_7972,N_5058,N_5915);
xor U7973 (N_7973,N_5015,N_6387);
nand U7974 (N_7974,N_7385,N_5819);
xnor U7975 (N_7975,N_6685,N_7337);
and U7976 (N_7976,N_7067,N_6172);
or U7977 (N_7977,N_6245,N_5643);
nor U7978 (N_7978,N_7316,N_5684);
or U7979 (N_7979,N_5627,N_5875);
or U7980 (N_7980,N_6792,N_5288);
xnor U7981 (N_7981,N_6654,N_6051);
and U7982 (N_7982,N_6954,N_5573);
nand U7983 (N_7983,N_5965,N_7012);
xor U7984 (N_7984,N_6806,N_7455);
xnor U7985 (N_7985,N_6173,N_5800);
and U7986 (N_7986,N_6456,N_5532);
and U7987 (N_7987,N_5262,N_5163);
nor U7988 (N_7988,N_6322,N_5186);
nand U7989 (N_7989,N_6108,N_6744);
and U7990 (N_7990,N_6191,N_6467);
nand U7991 (N_7991,N_6540,N_5603);
nor U7992 (N_7992,N_7137,N_6851);
nor U7993 (N_7993,N_6166,N_6503);
xnor U7994 (N_7994,N_6937,N_5457);
nand U7995 (N_7995,N_6416,N_6497);
nand U7996 (N_7996,N_7235,N_6558);
or U7997 (N_7997,N_6016,N_7134);
and U7998 (N_7998,N_6872,N_5636);
xor U7999 (N_7999,N_6190,N_5528);
or U8000 (N_8000,N_5981,N_5588);
nor U8001 (N_8001,N_5579,N_6055);
or U8002 (N_8002,N_6403,N_6964);
and U8003 (N_8003,N_5836,N_5090);
nor U8004 (N_8004,N_6555,N_5968);
xnor U8005 (N_8005,N_5357,N_5952);
and U8006 (N_8006,N_7125,N_5358);
nand U8007 (N_8007,N_5074,N_5623);
xnor U8008 (N_8008,N_5155,N_5440);
nand U8009 (N_8009,N_6791,N_5794);
nand U8010 (N_8010,N_5584,N_6049);
xnor U8011 (N_8011,N_5135,N_7165);
nand U8012 (N_8012,N_6163,N_5858);
nand U8013 (N_8013,N_5591,N_5432);
or U8014 (N_8014,N_5046,N_5624);
or U8015 (N_8015,N_5852,N_5156);
nand U8016 (N_8016,N_7417,N_6501);
and U8017 (N_8017,N_6833,N_6453);
nand U8018 (N_8018,N_7157,N_6372);
and U8019 (N_8019,N_6013,N_6511);
nand U8020 (N_8020,N_6704,N_5277);
nor U8021 (N_8021,N_6878,N_5658);
and U8022 (N_8022,N_6195,N_5607);
nand U8023 (N_8023,N_7264,N_5775);
nor U8024 (N_8024,N_7440,N_6749);
and U8025 (N_8025,N_7196,N_6089);
nor U8026 (N_8026,N_6228,N_5338);
xnor U8027 (N_8027,N_5121,N_6636);
and U8028 (N_8028,N_6452,N_6522);
nand U8029 (N_8029,N_5385,N_6846);
and U8030 (N_8030,N_7266,N_6424);
and U8031 (N_8031,N_7407,N_7124);
nor U8032 (N_8032,N_5523,N_5256);
nor U8033 (N_8033,N_7310,N_7056);
xnor U8034 (N_8034,N_5144,N_6554);
xnor U8035 (N_8035,N_6432,N_6399);
nor U8036 (N_8036,N_5311,N_7353);
nor U8037 (N_8037,N_5259,N_7286);
nand U8038 (N_8038,N_5078,N_5004);
xnor U8039 (N_8039,N_6278,N_6610);
xnor U8040 (N_8040,N_6912,N_6103);
and U8041 (N_8041,N_5028,N_6518);
nand U8042 (N_8042,N_6798,N_7209);
or U8043 (N_8043,N_6598,N_5349);
xnor U8044 (N_8044,N_6294,N_7336);
and U8045 (N_8045,N_5409,N_6115);
or U8046 (N_8046,N_7099,N_6093);
nand U8047 (N_8047,N_6682,N_6270);
nand U8048 (N_8048,N_7167,N_7386);
nand U8049 (N_8049,N_5141,N_7045);
nor U8050 (N_8050,N_6821,N_7349);
nand U8051 (N_8051,N_7303,N_5067);
xor U8052 (N_8052,N_6817,N_7250);
and U8053 (N_8053,N_6677,N_5691);
nand U8054 (N_8054,N_5652,N_5463);
and U8055 (N_8055,N_6794,N_6559);
nor U8056 (N_8056,N_6320,N_7058);
and U8057 (N_8057,N_5407,N_6378);
and U8058 (N_8058,N_5254,N_5334);
xor U8059 (N_8059,N_6038,N_6626);
xor U8060 (N_8060,N_7350,N_5807);
nor U8061 (N_8061,N_5025,N_5075);
nand U8062 (N_8062,N_6020,N_5692);
or U8063 (N_8063,N_5041,N_5125);
nand U8064 (N_8064,N_6699,N_7497);
nand U8065 (N_8065,N_6462,N_5213);
xnor U8066 (N_8066,N_5991,N_6576);
nand U8067 (N_8067,N_6723,N_6727);
nand U8068 (N_8068,N_6183,N_7436);
nand U8069 (N_8069,N_6763,N_6411);
or U8070 (N_8070,N_6517,N_6523);
or U8071 (N_8071,N_6006,N_6572);
xnor U8072 (N_8072,N_6255,N_7078);
xnor U8073 (N_8073,N_6917,N_5208);
nand U8074 (N_8074,N_6224,N_5193);
nor U8075 (N_8075,N_6620,N_5835);
or U8076 (N_8076,N_6343,N_6512);
xnor U8077 (N_8077,N_5871,N_5734);
xor U8078 (N_8078,N_7057,N_5681);
xnor U8079 (N_8079,N_6905,N_6275);
and U8080 (N_8080,N_5290,N_6616);
and U8081 (N_8081,N_5695,N_6177);
or U8082 (N_8082,N_6446,N_7247);
or U8083 (N_8083,N_5799,N_6499);
and U8084 (N_8084,N_6201,N_5085);
and U8085 (N_8085,N_5089,N_5507);
nor U8086 (N_8086,N_5042,N_6951);
nor U8087 (N_8087,N_5571,N_5921);
xor U8088 (N_8088,N_5766,N_5620);
nand U8089 (N_8089,N_5777,N_6797);
nor U8090 (N_8090,N_5034,N_5045);
and U8091 (N_8091,N_6785,N_6122);
xnor U8092 (N_8092,N_5711,N_6261);
nor U8093 (N_8093,N_6046,N_5433);
xnor U8094 (N_8094,N_7422,N_6738);
and U8095 (N_8095,N_5496,N_5922);
or U8096 (N_8096,N_6911,N_5197);
or U8097 (N_8097,N_6137,N_6181);
nor U8098 (N_8098,N_5550,N_6637);
and U8099 (N_8099,N_5199,N_5894);
nand U8100 (N_8100,N_5920,N_7277);
or U8101 (N_8101,N_7261,N_7184);
nand U8102 (N_8102,N_6217,N_5750);
nand U8103 (N_8103,N_6942,N_5478);
nor U8104 (N_8104,N_7370,N_5119);
nand U8105 (N_8105,N_7149,N_7319);
nor U8106 (N_8106,N_6056,N_5312);
or U8107 (N_8107,N_7281,N_7242);
nand U8108 (N_8108,N_5026,N_5343);
and U8109 (N_8109,N_5802,N_6710);
or U8110 (N_8110,N_5933,N_5397);
xnor U8111 (N_8111,N_6135,N_5570);
and U8112 (N_8112,N_5351,N_5821);
nand U8113 (N_8113,N_6360,N_5009);
or U8114 (N_8114,N_5097,N_7490);
or U8115 (N_8115,N_6428,N_6634);
nand U8116 (N_8116,N_7499,N_6601);
xor U8117 (N_8117,N_5563,N_7214);
nand U8118 (N_8118,N_6553,N_5785);
and U8119 (N_8119,N_5514,N_7464);
nand U8120 (N_8120,N_6840,N_7219);
nand U8121 (N_8121,N_5049,N_6703);
xor U8122 (N_8122,N_7169,N_5562);
nand U8123 (N_8123,N_6632,N_6722);
xor U8124 (N_8124,N_5031,N_6313);
nand U8125 (N_8125,N_6975,N_5517);
or U8126 (N_8126,N_6679,N_5061);
nand U8127 (N_8127,N_6212,N_6938);
or U8128 (N_8128,N_6272,N_6269);
or U8129 (N_8129,N_6861,N_6145);
nand U8130 (N_8130,N_5877,N_7122);
and U8131 (N_8131,N_6280,N_6946);
and U8132 (N_8132,N_7399,N_7092);
xnor U8133 (N_8133,N_5318,N_5759);
nor U8134 (N_8134,N_6592,N_5640);
nand U8135 (N_8135,N_7156,N_5650);
xor U8136 (N_8136,N_5988,N_6918);
nand U8137 (N_8137,N_5266,N_6149);
and U8138 (N_8138,N_6578,N_6069);
xnor U8139 (N_8139,N_5743,N_6943);
or U8140 (N_8140,N_5669,N_6441);
or U8141 (N_8141,N_5634,N_7073);
xor U8142 (N_8142,N_5924,N_7023);
and U8143 (N_8143,N_7448,N_7460);
or U8144 (N_8144,N_5590,N_5095);
nand U8145 (N_8145,N_6935,N_6480);
xor U8146 (N_8146,N_7449,N_6849);
and U8147 (N_8147,N_5169,N_7361);
or U8148 (N_8148,N_5113,N_6701);
or U8149 (N_8149,N_6814,N_6675);
nand U8150 (N_8150,N_5815,N_6117);
nand U8151 (N_8151,N_6571,N_6318);
or U8152 (N_8152,N_6305,N_7376);
and U8153 (N_8153,N_5900,N_6799);
nand U8154 (N_8154,N_5231,N_6205);
or U8155 (N_8155,N_7096,N_6066);
and U8156 (N_8156,N_5761,N_7405);
or U8157 (N_8157,N_6099,N_6220);
or U8158 (N_8158,N_7005,N_6429);
nand U8159 (N_8159,N_5016,N_5526);
or U8160 (N_8160,N_5599,N_6418);
and U8161 (N_8161,N_6481,N_6494);
or U8162 (N_8162,N_6788,N_6914);
xnor U8163 (N_8163,N_5104,N_6962);
nor U8164 (N_8164,N_5276,N_5790);
or U8165 (N_8165,N_5280,N_6291);
xnor U8166 (N_8166,N_5225,N_6311);
and U8167 (N_8167,N_5601,N_6882);
and U8168 (N_8168,N_6752,N_6873);
xor U8169 (N_8169,N_5204,N_7003);
nor U8170 (N_8170,N_6297,N_7451);
xnor U8171 (N_8171,N_5174,N_6673);
and U8172 (N_8172,N_5316,N_5561);
nand U8173 (N_8173,N_6638,N_5752);
and U8174 (N_8174,N_5138,N_6243);
and U8175 (N_8175,N_7409,N_6940);
xnor U8176 (N_8176,N_5932,N_5366);
nand U8177 (N_8177,N_5872,N_5893);
nor U8178 (N_8178,N_6358,N_6393);
xor U8179 (N_8179,N_5597,N_6492);
and U8180 (N_8180,N_5546,N_5917);
and U8181 (N_8181,N_6326,N_6563);
nand U8182 (N_8182,N_7028,N_5906);
xnor U8183 (N_8183,N_5645,N_6691);
or U8184 (N_8184,N_5065,N_6179);
and U8185 (N_8185,N_7276,N_6408);
xnor U8186 (N_8186,N_5639,N_5284);
nand U8187 (N_8187,N_6600,N_6575);
nor U8188 (N_8188,N_6996,N_5942);
or U8189 (N_8189,N_6353,N_5891);
and U8190 (N_8190,N_6628,N_7039);
or U8191 (N_8191,N_5066,N_6674);
xnor U8192 (N_8192,N_5328,N_6551);
and U8193 (N_8193,N_6608,N_6855);
nor U8194 (N_8194,N_5762,N_6074);
xnor U8195 (N_8195,N_7041,N_6256);
or U8196 (N_8196,N_6011,N_7042);
or U8197 (N_8197,N_5226,N_5660);
nor U8198 (N_8198,N_5694,N_6597);
nand U8199 (N_8199,N_6073,N_5716);
and U8200 (N_8200,N_5002,N_7132);
or U8201 (N_8201,N_5949,N_7431);
or U8202 (N_8202,N_5855,N_7430);
nor U8203 (N_8203,N_6750,N_6154);
and U8204 (N_8204,N_6400,N_5462);
or U8205 (N_8205,N_7107,N_5796);
or U8206 (N_8206,N_7290,N_7258);
nand U8207 (N_8207,N_6090,N_5557);
nand U8208 (N_8208,N_5830,N_5285);
xor U8209 (N_8209,N_7265,N_7244);
and U8210 (N_8210,N_5236,N_6527);
or U8211 (N_8211,N_6933,N_7379);
xnor U8212 (N_8212,N_6916,N_6260);
or U8213 (N_8213,N_5708,N_5778);
xnor U8214 (N_8214,N_6012,N_5435);
nor U8215 (N_8215,N_5438,N_6044);
nor U8216 (N_8216,N_5018,N_6031);
xnor U8217 (N_8217,N_7444,N_6970);
or U8218 (N_8218,N_5997,N_6042);
nor U8219 (N_8219,N_5896,N_5604);
nand U8220 (N_8220,N_6029,N_5094);
or U8221 (N_8221,N_7381,N_6215);
nand U8222 (N_8222,N_7139,N_5503);
and U8223 (N_8223,N_6556,N_5157);
nand U8224 (N_8224,N_5919,N_6533);
or U8225 (N_8225,N_7075,N_6960);
or U8226 (N_8226,N_6225,N_6668);
xnor U8227 (N_8227,N_5782,N_7215);
and U8228 (N_8228,N_5758,N_6605);
nor U8229 (N_8229,N_6388,N_6721);
nor U8230 (N_8230,N_7441,N_7391);
nor U8231 (N_8231,N_5461,N_5196);
nand U8232 (N_8232,N_5606,N_6854);
nand U8233 (N_8233,N_6332,N_7476);
nor U8234 (N_8234,N_5816,N_6707);
nand U8235 (N_8235,N_7396,N_5696);
nand U8236 (N_8236,N_6043,N_7226);
nor U8237 (N_8237,N_7324,N_6505);
and U8238 (N_8238,N_6804,N_7355);
nor U8239 (N_8239,N_5360,N_6528);
nand U8240 (N_8240,N_5413,N_5497);
xor U8241 (N_8241,N_6966,N_6815);
nand U8242 (N_8242,N_7334,N_5934);
xnor U8243 (N_8243,N_6022,N_7318);
or U8244 (N_8244,N_7143,N_5022);
or U8245 (N_8245,N_5499,N_5282);
xnor U8246 (N_8246,N_7469,N_7010);
xnor U8247 (N_8247,N_6939,N_6476);
and U8248 (N_8248,N_5849,N_5971);
nand U8249 (N_8249,N_6404,N_6457);
xnor U8250 (N_8250,N_6868,N_6138);
nor U8251 (N_8251,N_5441,N_6014);
nor U8252 (N_8252,N_7326,N_5101);
xnor U8253 (N_8253,N_7471,N_7224);
and U8254 (N_8254,N_6080,N_6984);
nor U8255 (N_8255,N_6880,N_5912);
nand U8256 (N_8256,N_5324,N_6237);
and U8257 (N_8257,N_6053,N_5255);
nor U8258 (N_8258,N_5205,N_6760);
nand U8259 (N_8259,N_6805,N_6891);
or U8260 (N_8260,N_7064,N_5361);
or U8261 (N_8261,N_6644,N_5840);
and U8262 (N_8262,N_7019,N_6768);
nor U8263 (N_8263,N_7189,N_6857);
and U8264 (N_8264,N_5279,N_6542);
nand U8265 (N_8265,N_6422,N_5656);
or U8266 (N_8266,N_5809,N_5340);
xor U8267 (N_8267,N_5260,N_5632);
nor U8268 (N_8268,N_6180,N_6843);
and U8269 (N_8269,N_6536,N_6826);
nor U8270 (N_8270,N_6257,N_5393);
nand U8271 (N_8271,N_7017,N_7240);
nor U8272 (N_8272,N_5713,N_5076);
and U8273 (N_8273,N_7404,N_5787);
xnor U8274 (N_8274,N_5247,N_6096);
nand U8275 (N_8275,N_7063,N_5572);
or U8276 (N_8276,N_6646,N_7278);
or U8277 (N_8277,N_6007,N_7138);
or U8278 (N_8278,N_5501,N_6651);
or U8279 (N_8279,N_5346,N_5667);
and U8280 (N_8280,N_6035,N_7450);
and U8281 (N_8281,N_5408,N_6746);
xnor U8282 (N_8282,N_7006,N_7486);
xor U8283 (N_8283,N_6694,N_6102);
nand U8284 (N_8284,N_5382,N_7153);
nor U8285 (N_8285,N_5153,N_7140);
nor U8286 (N_8286,N_6713,N_6150);
nor U8287 (N_8287,N_6758,N_5735);
nor U8288 (N_8288,N_5720,N_5774);
xnor U8289 (N_8289,N_6614,N_7119);
and U8290 (N_8290,N_6742,N_6538);
or U8291 (N_8291,N_5615,N_7339);
or U8292 (N_8292,N_6241,N_5491);
nor U8293 (N_8293,N_7059,N_6702);
and U8294 (N_8294,N_5447,N_7289);
nand U8295 (N_8295,N_6602,N_6119);
nor U8296 (N_8296,N_5027,N_5175);
nor U8297 (N_8297,N_7351,N_6835);
or U8298 (N_8298,N_6687,N_5829);
nor U8299 (N_8299,N_6282,N_7321);
and U8300 (N_8300,N_5574,N_5731);
xnor U8301 (N_8301,N_5088,N_5292);
nand U8302 (N_8302,N_6375,N_5315);
xor U8303 (N_8303,N_5180,N_6244);
nor U8304 (N_8304,N_5964,N_5235);
and U8305 (N_8305,N_5446,N_5907);
and U8306 (N_8306,N_5985,N_5476);
or U8307 (N_8307,N_6807,N_6338);
xnor U8308 (N_8308,N_5147,N_6449);
or U8309 (N_8309,N_7048,N_5335);
xnor U8310 (N_8310,N_7423,N_5786);
or U8311 (N_8311,N_6136,N_5773);
nor U8312 (N_8312,N_7098,N_6782);
and U8313 (N_8313,N_5391,N_7411);
or U8314 (N_8314,N_5109,N_7190);
and U8315 (N_8315,N_7480,N_7309);
nor U8316 (N_8316,N_6357,N_6383);
nor U8317 (N_8317,N_7221,N_5294);
or U8318 (N_8318,N_5149,N_5654);
xor U8319 (N_8319,N_5165,N_5301);
nand U8320 (N_8320,N_6928,N_6168);
or U8321 (N_8321,N_6155,N_5672);
nand U8322 (N_8322,N_5477,N_5484);
nor U8323 (N_8323,N_5936,N_6466);
xnor U8324 (N_8324,N_6448,N_6296);
xnor U8325 (N_8325,N_5388,N_6661);
xor U8326 (N_8326,N_5494,N_6829);
or U8327 (N_8327,N_5106,N_6865);
or U8328 (N_8328,N_5689,N_6263);
xor U8329 (N_8329,N_5817,N_6530);
and U8330 (N_8330,N_7160,N_5179);
nand U8331 (N_8331,N_5229,N_5252);
nand U8332 (N_8332,N_6298,N_7348);
or U8333 (N_8333,N_5317,N_6196);
xor U8334 (N_8334,N_7114,N_5826);
xor U8335 (N_8335,N_7271,N_7161);
xnor U8336 (N_8336,N_5659,N_5935);
and U8337 (N_8337,N_6582,N_5246);
or U8338 (N_8338,N_5023,N_5728);
and U8339 (N_8339,N_5976,N_7091);
nor U8340 (N_8340,N_5542,N_6869);
nor U8341 (N_8341,N_7069,N_6974);
nor U8342 (N_8342,N_5291,N_7498);
nor U8343 (N_8343,N_5598,N_6284);
or U8344 (N_8344,N_5493,N_6734);
or U8345 (N_8345,N_6226,N_5715);
nor U8346 (N_8346,N_5183,N_5240);
or U8347 (N_8347,N_6997,N_6315);
nor U8348 (N_8348,N_5319,N_6336);
and U8349 (N_8349,N_5771,N_5788);
xor U8350 (N_8350,N_6325,N_5394);
or U8351 (N_8351,N_6599,N_7394);
xnor U8352 (N_8352,N_6097,N_7364);
nor U8353 (N_8353,N_5339,N_5464);
nor U8354 (N_8354,N_5551,N_5673);
nor U8355 (N_8355,N_5116,N_6715);
xnor U8356 (N_8356,N_7459,N_5212);
nand U8357 (N_8357,N_7485,N_5032);
xnor U8358 (N_8358,N_5892,N_5863);
nor U8359 (N_8359,N_6543,N_7275);
nand U8360 (N_8360,N_6789,N_5293);
nor U8361 (N_8361,N_5732,N_5117);
nand U8362 (N_8362,N_5158,N_5755);
or U8363 (N_8363,N_5377,N_5239);
nor U8364 (N_8364,N_5083,N_6130);
and U8365 (N_8365,N_6776,N_7145);
and U8366 (N_8366,N_7192,N_7270);
nor U8367 (N_8367,N_5940,N_5677);
or U8368 (N_8368,N_5539,N_6438);
or U8369 (N_8369,N_5502,N_6242);
and U8370 (N_8370,N_7374,N_5605);
xnor U8371 (N_8371,N_6688,N_5797);
nand U8372 (N_8372,N_6479,N_6957);
nor U8373 (N_8373,N_6248,N_5543);
nand U8374 (N_8374,N_6299,N_5261);
nor U8375 (N_8375,N_5616,N_5459);
or U8376 (N_8376,N_6709,N_6853);
nor U8377 (N_8377,N_6983,N_5485);
nand U8378 (N_8378,N_5950,N_5243);
nor U8379 (N_8379,N_6967,N_5030);
nand U8380 (N_8380,N_6875,N_7425);
xor U8381 (N_8381,N_5712,N_6539);
and U8382 (N_8382,N_5617,N_5354);
and U8383 (N_8383,N_6490,N_7287);
and U8384 (N_8384,N_5263,N_5744);
or U8385 (N_8385,N_6436,N_5772);
and U8386 (N_8386,N_6063,N_6341);
nor U8387 (N_8387,N_6083,N_5272);
xor U8388 (N_8388,N_7233,N_6348);
and U8389 (N_8389,N_5353,N_5390);
nand U8390 (N_8390,N_5287,N_5947);
or U8391 (N_8391,N_5465,N_7011);
nand U8392 (N_8392,N_5056,N_6356);
nor U8393 (N_8393,N_5480,N_6187);
and U8394 (N_8394,N_7315,N_7393);
and U8395 (N_8395,N_5581,N_6133);
or U8396 (N_8396,N_5454,N_5516);
and U8397 (N_8397,N_6286,N_5804);
and U8398 (N_8398,N_5946,N_5115);
and U8399 (N_8399,N_5416,N_7127);
or U8400 (N_8400,N_6067,N_5629);
nand U8401 (N_8401,N_6206,N_6686);
nor U8402 (N_8402,N_6355,N_6239);
nand U8403 (N_8403,N_6487,N_6010);
nand U8404 (N_8404,N_6027,N_5522);
and U8405 (N_8405,N_5931,N_7205);
nand U8406 (N_8406,N_7389,N_7014);
and U8407 (N_8407,N_6545,N_6184);
or U8408 (N_8408,N_6762,N_6409);
nor U8409 (N_8409,N_7253,N_6334);
nand U8410 (N_8410,N_6969,N_7251);
xnor U8411 (N_8411,N_5177,N_7390);
nor U8412 (N_8412,N_6803,N_5379);
nand U8413 (N_8413,N_7307,N_6350);
and U8414 (N_8414,N_5886,N_6635);
nand U8415 (N_8415,N_5714,N_7388);
or U8416 (N_8416,N_5195,N_7453);
xnor U8417 (N_8417,N_6444,N_5057);
or U8418 (N_8418,N_7060,N_5699);
or U8419 (N_8419,N_5182,N_6842);
xnor U8420 (N_8420,N_6828,N_6386);
and U8421 (N_8421,N_6486,N_6077);
xnor U8422 (N_8422,N_7129,N_5102);
nand U8423 (N_8423,N_5647,N_5202);
or U8424 (N_8424,N_7104,N_6607);
and U8425 (N_8425,N_5161,N_6544);
and U8426 (N_8426,N_5793,N_7072);
or U8427 (N_8427,N_7354,N_5745);
nor U8428 (N_8428,N_7338,N_7380);
nor U8429 (N_8429,N_6936,N_5566);
or U8430 (N_8430,N_5612,N_6639);
nand U8431 (N_8431,N_5355,N_7037);
nor U8432 (N_8432,N_7001,N_6015);
or U8433 (N_8433,N_6720,N_5707);
nand U8434 (N_8434,N_6028,N_5184);
and U8435 (N_8435,N_7170,N_6126);
and U8436 (N_8436,N_6070,N_5064);
xor U8437 (N_8437,N_6753,N_6790);
nand U8438 (N_8438,N_6395,N_5029);
and U8439 (N_8439,N_6468,N_5118);
and U8440 (N_8440,N_5943,N_6580);
and U8441 (N_8441,N_5431,N_7429);
or U8442 (N_8442,N_6811,N_5411);
nand U8443 (N_8443,N_5913,N_7257);
nand U8444 (N_8444,N_5885,N_7246);
or U8445 (N_8445,N_6898,N_5748);
or U8446 (N_8446,N_5897,N_5107);
and U8447 (N_8447,N_5129,N_5602);
xor U8448 (N_8448,N_6950,N_6624);
and U8449 (N_8449,N_5860,N_5336);
and U8450 (N_8450,N_5929,N_6795);
nand U8451 (N_8451,N_5369,N_7201);
nand U8452 (N_8452,N_6525,N_7021);
nor U8453 (N_8453,N_5832,N_6000);
nand U8454 (N_8454,N_7282,N_6755);
or U8455 (N_8455,N_7087,N_5222);
nor U8456 (N_8456,N_6700,N_5553);
xnor U8457 (N_8457,N_6088,N_7187);
xnor U8458 (N_8458,N_6825,N_5014);
xnor U8459 (N_8459,N_5417,N_5019);
or U8460 (N_8460,N_6922,N_5217);
xnor U8461 (N_8461,N_5979,N_5854);
nand U8462 (N_8462,N_6307,N_6406);
and U8463 (N_8463,N_7274,N_6506);
xnor U8464 (N_8464,N_6059,N_5086);
and U8465 (N_8465,N_6301,N_6347);
and U8466 (N_8466,N_7433,N_6831);
nor U8467 (N_8467,N_6971,N_5567);
xnor U8468 (N_8468,N_6552,N_5544);
nor U8469 (N_8469,N_6793,N_7152);
xor U8470 (N_8470,N_6264,N_6488);
and U8471 (N_8471,N_7375,N_6770);
xnor U8472 (N_8472,N_6359,N_6541);
or U8473 (N_8473,N_5740,N_7225);
xnor U8474 (N_8474,N_5257,N_7288);
or U8475 (N_8475,N_6052,N_6292);
nor U8476 (N_8476,N_6192,N_5007);
nor U8477 (N_8477,N_5596,N_5901);
nand U8478 (N_8478,N_7468,N_5676);
and U8479 (N_8479,N_5700,N_5846);
nand U8480 (N_8480,N_5941,N_6465);
nand U8481 (N_8481,N_6665,N_7036);
nand U8482 (N_8482,N_6352,N_6739);
xnor U8483 (N_8483,N_6507,N_6881);
nand U8484 (N_8484,N_5047,N_5705);
nor U8485 (N_8485,N_7347,N_5052);
and U8486 (N_8486,N_5998,N_5474);
xnor U8487 (N_8487,N_5882,N_7359);
xnor U8488 (N_8488,N_5812,N_7317);
nand U8489 (N_8489,N_5881,N_5564);
nor U8490 (N_8490,N_7108,N_6157);
nor U8491 (N_8491,N_7305,N_6081);
or U8492 (N_8492,N_5092,N_7400);
xnor U8493 (N_8493,N_6057,N_7263);
and U8494 (N_8494,N_5228,N_6233);
xor U8495 (N_8495,N_6838,N_6283);
and U8496 (N_8496,N_5898,N_5309);
nor U8497 (N_8497,N_6198,N_5698);
or U8498 (N_8498,N_6864,N_6910);
xnor U8499 (N_8499,N_5631,N_6065);
xor U8500 (N_8500,N_6213,N_5453);
nand U8501 (N_8501,N_5726,N_6435);
or U8502 (N_8502,N_5798,N_6164);
nor U8503 (N_8503,N_5646,N_5048);
xnor U8504 (N_8504,N_5281,N_7142);
or U8505 (N_8505,N_6174,N_7040);
xnor U8506 (N_8506,N_5834,N_5910);
xnor U8507 (N_8507,N_6949,N_6832);
or U8508 (N_8508,N_5000,N_7168);
nor U8509 (N_8509,N_7106,N_7329);
xnor U8510 (N_8510,N_6989,N_6050);
xor U8511 (N_8511,N_6941,N_6368);
xor U8512 (N_8512,N_7007,N_5286);
xor U8513 (N_8513,N_5757,N_5990);
nand U8514 (N_8514,N_5401,N_6362);
xnor U8515 (N_8515,N_6659,N_5827);
xnor U8516 (N_8516,N_6210,N_5746);
nor U8517 (N_8517,N_6469,N_5721);
nand U8518 (N_8518,N_5776,N_5506);
nand U8519 (N_8519,N_7174,N_5420);
xnor U8520 (N_8520,N_6667,N_6976);
or U8521 (N_8521,N_5181,N_6211);
and U8522 (N_8522,N_6302,N_5400);
nand U8523 (N_8523,N_6672,N_6327);
xor U8524 (N_8524,N_6153,N_5806);
or U8525 (N_8525,N_5838,N_6223);
nor U8526 (N_8526,N_5364,N_5114);
xor U8527 (N_8527,N_7110,N_7009);
xor U8528 (N_8528,N_5481,N_6246);
and U8529 (N_8529,N_7403,N_5344);
nand U8530 (N_8530,N_5857,N_6537);
and U8531 (N_8531,N_5719,N_6204);
and U8532 (N_8532,N_5073,N_6231);
nor U8533 (N_8533,N_5668,N_5425);
nand U8534 (N_8534,N_7027,N_6214);
xor U8535 (N_8535,N_7051,N_5937);
nor U8536 (N_8536,N_5132,N_5341);
or U8537 (N_8537,N_7312,N_5560);
xor U8538 (N_8538,N_6693,N_7262);
nor U8539 (N_8539,N_6985,N_5283);
and U8540 (N_8540,N_7094,N_5458);
nand U8541 (N_8541,N_6565,N_6745);
or U8542 (N_8542,N_7022,N_7477);
xor U8543 (N_8543,N_5452,N_6009);
xnor U8544 (N_8544,N_5206,N_5873);
nor U8545 (N_8545,N_5011,N_6484);
and U8546 (N_8546,N_5780,N_7146);
nor U8547 (N_8547,N_6801,N_6587);
xor U8548 (N_8548,N_5527,N_5861);
xor U8549 (N_8549,N_6001,N_5054);
nor U8550 (N_8550,N_5405,N_6381);
nand U8551 (N_8551,N_6227,N_5904);
xor U8552 (N_8552,N_5150,N_6781);
xnor U8553 (N_8553,N_6314,N_6871);
nor U8554 (N_8554,N_5249,N_7383);
and U8555 (N_8555,N_5630,N_5756);
and U8556 (N_8556,N_6309,N_6596);
and U8557 (N_8557,N_7150,N_5975);
and U8558 (N_8558,N_5154,N_6382);
or U8559 (N_8559,N_6879,N_5843);
nand U8560 (N_8560,N_5500,N_6230);
nand U8561 (N_8561,N_6277,N_5303);
nor U8562 (N_8562,N_7333,N_5505);
xor U8563 (N_8563,N_5145,N_7148);
nand U8564 (N_8564,N_5190,N_5051);
xnor U8565 (N_8565,N_6783,N_6958);
xnor U8566 (N_8566,N_7291,N_6207);
or U8567 (N_8567,N_5867,N_6892);
xor U8568 (N_8568,N_5538,N_5297);
nand U8569 (N_8569,N_6109,N_6915);
nand U8570 (N_8570,N_6604,N_6585);
and U8571 (N_8571,N_7325,N_5295);
nand U8572 (N_8572,N_6200,N_6948);
nand U8573 (N_8573,N_6732,N_6583);
nand U8574 (N_8574,N_7171,N_7115);
nor U8575 (N_8575,N_7415,N_5039);
nor U8576 (N_8576,N_6574,N_5690);
and U8577 (N_8577,N_5313,N_7034);
xor U8578 (N_8578,N_5814,N_5622);
or U8579 (N_8579,N_6524,N_6931);
xor U8580 (N_8580,N_5299,N_5961);
nor U8581 (N_8581,N_6862,N_6779);
or U8582 (N_8582,N_6748,N_7322);
nor U8583 (N_8583,N_5969,N_6866);
and U8584 (N_8584,N_5218,N_6100);
nand U8585 (N_8585,N_5242,N_5954);
nand U8586 (N_8586,N_7068,N_6573);
or U8587 (N_8587,N_6023,N_7102);
nand U8588 (N_8588,N_6351,N_6110);
nor U8589 (N_8589,N_7372,N_6414);
nand U8590 (N_8590,N_7095,N_6162);
nor U8591 (N_8591,N_5751,N_5337);
nor U8592 (N_8592,N_5779,N_5418);
xor U8593 (N_8593,N_5168,N_5248);
xnor U8594 (N_8594,N_7489,N_5060);
xnor U8595 (N_8595,N_6652,N_6238);
nor U8596 (N_8596,N_6773,N_5482);
xor U8597 (N_8597,N_6471,N_5989);
nor U8598 (N_8598,N_6564,N_5473);
and U8599 (N_8599,N_6681,N_7079);
or U8600 (N_8600,N_6176,N_6397);
nand U8601 (N_8601,N_5308,N_5139);
xor U8602 (N_8602,N_6590,N_5747);
xor U8603 (N_8603,N_6737,N_6114);
nor U8604 (N_8604,N_5718,N_5483);
or U8605 (N_8605,N_5050,N_5406);
or U8606 (N_8606,N_6988,N_6316);
nand U8607 (N_8607,N_7241,N_6202);
and U8608 (N_8608,N_6474,N_5230);
or U8609 (N_8609,N_5069,N_5512);
xnor U8610 (N_8610,N_6279,N_6364);
and U8611 (N_8611,N_5162,N_5091);
nand U8612 (N_8612,N_5378,N_7447);
and U8613 (N_8613,N_6595,N_5103);
nand U8614 (N_8614,N_5686,N_5320);
and U8615 (N_8615,N_5554,N_5859);
nand U8616 (N_8616,N_5878,N_6458);
nor U8617 (N_8617,N_5372,N_5733);
or U8618 (N_8618,N_5577,N_6736);
xor U8619 (N_8619,N_7128,N_5080);
nand U8620 (N_8620,N_5960,N_5593);
xnor U8621 (N_8621,N_6930,N_7038);
and U8622 (N_8622,N_5655,N_6062);
and U8623 (N_8623,N_5345,N_7473);
and U8624 (N_8624,N_5739,N_5035);
and U8625 (N_8625,N_5350,N_5376);
or U8626 (N_8626,N_5099,N_5895);
and U8627 (N_8627,N_7412,N_6293);
or U8628 (N_8628,N_6485,N_5451);
nor U8629 (N_8629,N_6994,N_6491);
or U8630 (N_8630,N_6570,N_6041);
xor U8631 (N_8631,N_5944,N_6054);
nor U8632 (N_8632,N_5992,N_6249);
nand U8633 (N_8633,N_7461,N_5143);
and U8634 (N_8634,N_5445,N_5271);
and U8635 (N_8635,N_5436,N_6633);
xnor U8636 (N_8636,N_5621,N_5515);
nor U8637 (N_8637,N_7395,N_7112);
nand U8638 (N_8638,N_7234,N_7344);
nand U8639 (N_8639,N_6955,N_5760);
nand U8640 (N_8640,N_5706,N_6968);
xnor U8641 (N_8641,N_5958,N_6952);
or U8642 (N_8642,N_7248,N_5945);
nand U8643 (N_8643,N_6266,N_6711);
nor U8644 (N_8644,N_5096,N_5864);
or U8645 (N_8645,N_5427,N_7320);
nand U8646 (N_8646,N_7366,N_7206);
xnor U8647 (N_8647,N_5529,N_6306);
xor U8648 (N_8648,N_5549,N_6240);
and U8649 (N_8649,N_5795,N_5348);
xnor U8650 (N_8650,N_6886,N_6698);
nor U8651 (N_8651,N_6229,N_5578);
xor U8652 (N_8652,N_6346,N_5649);
and U8653 (N_8653,N_5442,N_6764);
and U8654 (N_8654,N_6726,N_7445);
nor U8655 (N_8655,N_6289,N_6775);
and U8656 (N_8656,N_6194,N_5918);
and U8657 (N_8657,N_5509,N_5450);
nor U8658 (N_8658,N_7384,N_5082);
and U8659 (N_8659,N_5203,N_5770);
xnor U8660 (N_8660,N_5146,N_6500);
or U8661 (N_8661,N_5359,N_6118);
nor U8662 (N_8662,N_6045,N_7207);
and U8663 (N_8663,N_6894,N_7401);
or U8664 (N_8664,N_5736,N_6925);
and U8665 (N_8665,N_6445,N_5224);
nand U8666 (N_8666,N_5310,N_7294);
xnor U8667 (N_8667,N_6724,N_5887);
xor U8668 (N_8668,N_7204,N_5519);
nand U8669 (N_8669,N_7421,N_5521);
nor U8670 (N_8670,N_5159,N_6761);
and U8671 (N_8671,N_7131,N_6557);
nor U8672 (N_8672,N_7424,N_5530);
xnor U8673 (N_8673,N_6765,N_6591);
nor U8674 (N_8674,N_6757,N_5805);
xor U8675 (N_8675,N_7191,N_6508);
xnor U8676 (N_8676,N_6502,N_5191);
xor U8677 (N_8677,N_6896,N_5661);
or U8678 (N_8678,N_7239,N_5911);
or U8679 (N_8679,N_6250,N_6680);
or U8680 (N_8680,N_6586,N_7172);
and U8681 (N_8681,N_7118,N_5844);
or U8682 (N_8682,N_6820,N_7188);
and U8683 (N_8683,N_6510,N_6778);
nor U8684 (N_8684,N_5013,N_6463);
nand U8685 (N_8685,N_7163,N_6140);
xor U8686 (N_8686,N_5618,N_5729);
nand U8687 (N_8687,N_6308,N_6107);
and U8688 (N_8688,N_6440,N_6902);
nand U8689 (N_8689,N_6909,N_6185);
or U8690 (N_8690,N_7141,N_6098);
or U8691 (N_8691,N_5582,N_5038);
nand U8692 (N_8692,N_6741,N_7462);
or U8693 (N_8693,N_5754,N_5449);
xor U8694 (N_8694,N_7176,N_7173);
xor U8695 (N_8695,N_5456,N_6427);
and U8696 (N_8696,N_5040,N_5314);
or U8697 (N_8697,N_6774,N_5269);
nor U8698 (N_8698,N_6611,N_6531);
or U8699 (N_8699,N_7154,N_5742);
or U8700 (N_8700,N_5703,N_6981);
and U8701 (N_8701,N_5614,N_5232);
and U8702 (N_8702,N_6276,N_7254);
xnor U8703 (N_8703,N_6641,N_6288);
nor U8704 (N_8704,N_6377,N_7088);
nor U8705 (N_8705,N_5823,N_6483);
or U8706 (N_8706,N_6627,N_7162);
or U8707 (N_8707,N_6689,N_5471);
and U8708 (N_8708,N_5763,N_6678);
xnor U8709 (N_8709,N_6259,N_7357);
nand U8710 (N_8710,N_5342,N_6169);
or U8711 (N_8711,N_5874,N_5120);
nand U8712 (N_8712,N_5422,N_7081);
or U8713 (N_8713,N_7217,N_6786);
and U8714 (N_8714,N_6472,N_5081);
nor U8715 (N_8715,N_6209,N_6426);
xor U8716 (N_8716,N_5201,N_6058);
and U8717 (N_8717,N_7299,N_6859);
and U8718 (N_8718,N_5524,N_5194);
nor U8719 (N_8719,N_6003,N_7029);
nand U8720 (N_8720,N_6019,N_7327);
nor U8721 (N_8721,N_7420,N_6105);
and U8722 (N_8722,N_7332,N_6919);
xnor U8723 (N_8723,N_7428,N_6728);
nand U8724 (N_8724,N_7186,N_6904);
and U8725 (N_8725,N_6921,N_5818);
xnor U8726 (N_8726,N_5813,N_7356);
or U8727 (N_8727,N_6995,N_5036);
nor U8728 (N_8728,N_7360,N_6132);
nand U8729 (N_8729,N_7218,N_6858);
and U8730 (N_8730,N_5363,N_5216);
and U8731 (N_8731,N_7231,N_5134);
xor U8732 (N_8732,N_6532,N_5510);
and U8733 (N_8733,N_5414,N_5862);
or U8734 (N_8734,N_7371,N_6094);
and U8735 (N_8735,N_6271,N_5467);
or U8736 (N_8736,N_6199,N_7062);
nand U8737 (N_8737,N_5020,N_5923);
nand U8738 (N_8738,N_7284,N_5723);
or U8739 (N_8739,N_6945,N_6112);
nand U8740 (N_8740,N_5133,N_5995);
nor U8741 (N_8741,N_5552,N_5492);
and U8742 (N_8742,N_5273,N_5531);
nand U8743 (N_8743,N_7018,N_7255);
nand U8744 (N_8744,N_6759,N_5784);
xnor U8745 (N_8745,N_6147,N_6714);
nand U8746 (N_8746,N_5657,N_6290);
xnor U8747 (N_8747,N_7456,N_7482);
nand U8748 (N_8748,N_5326,N_7297);
xor U8749 (N_8749,N_6670,N_5839);
or U8750 (N_8750,N_6351,N_7270);
and U8751 (N_8751,N_5030,N_5365);
nand U8752 (N_8752,N_5747,N_6830);
xor U8753 (N_8753,N_5455,N_5494);
xor U8754 (N_8754,N_7208,N_5776);
nand U8755 (N_8755,N_5506,N_6379);
xnor U8756 (N_8756,N_6920,N_7292);
and U8757 (N_8757,N_5869,N_5675);
or U8758 (N_8758,N_6410,N_7214);
nor U8759 (N_8759,N_5952,N_6602);
or U8760 (N_8760,N_6207,N_5468);
nand U8761 (N_8761,N_6926,N_7320);
xnor U8762 (N_8762,N_5946,N_6410);
or U8763 (N_8763,N_6288,N_6476);
nor U8764 (N_8764,N_7302,N_7368);
nor U8765 (N_8765,N_7137,N_5593);
or U8766 (N_8766,N_6971,N_5403);
xor U8767 (N_8767,N_6294,N_7461);
xnor U8768 (N_8768,N_7372,N_5529);
nand U8769 (N_8769,N_6360,N_7229);
nor U8770 (N_8770,N_7217,N_6325);
xor U8771 (N_8771,N_6676,N_7382);
xnor U8772 (N_8772,N_7493,N_7188);
nor U8773 (N_8773,N_6471,N_7007);
and U8774 (N_8774,N_5523,N_6855);
and U8775 (N_8775,N_5131,N_6002);
xor U8776 (N_8776,N_5756,N_6806);
and U8777 (N_8777,N_5197,N_5699);
nand U8778 (N_8778,N_5811,N_6977);
xnor U8779 (N_8779,N_6419,N_6074);
xnor U8780 (N_8780,N_5334,N_7214);
nand U8781 (N_8781,N_7295,N_7377);
xor U8782 (N_8782,N_6926,N_5459);
nand U8783 (N_8783,N_7099,N_5001);
or U8784 (N_8784,N_5607,N_5709);
and U8785 (N_8785,N_6639,N_7238);
or U8786 (N_8786,N_7086,N_5016);
and U8787 (N_8787,N_6195,N_7320);
or U8788 (N_8788,N_6090,N_5951);
or U8789 (N_8789,N_5290,N_5312);
xnor U8790 (N_8790,N_6387,N_5653);
and U8791 (N_8791,N_7095,N_6279);
and U8792 (N_8792,N_6084,N_5268);
or U8793 (N_8793,N_6649,N_7419);
nand U8794 (N_8794,N_5582,N_6530);
xor U8795 (N_8795,N_6247,N_6717);
and U8796 (N_8796,N_6442,N_7068);
xnor U8797 (N_8797,N_5037,N_7423);
nor U8798 (N_8798,N_6130,N_5651);
nor U8799 (N_8799,N_5951,N_6414);
or U8800 (N_8800,N_5246,N_6613);
nand U8801 (N_8801,N_5624,N_6643);
or U8802 (N_8802,N_5832,N_7497);
xnor U8803 (N_8803,N_5720,N_5934);
nand U8804 (N_8804,N_6687,N_7311);
and U8805 (N_8805,N_6570,N_6239);
xnor U8806 (N_8806,N_5680,N_6121);
xnor U8807 (N_8807,N_6287,N_7464);
xnor U8808 (N_8808,N_6078,N_5475);
and U8809 (N_8809,N_5993,N_7093);
nand U8810 (N_8810,N_5704,N_5154);
and U8811 (N_8811,N_5406,N_7337);
and U8812 (N_8812,N_6282,N_5299);
xnor U8813 (N_8813,N_6078,N_7404);
nand U8814 (N_8814,N_7287,N_6466);
and U8815 (N_8815,N_5851,N_5832);
xor U8816 (N_8816,N_5514,N_7063);
or U8817 (N_8817,N_7128,N_5904);
xnor U8818 (N_8818,N_6374,N_5272);
or U8819 (N_8819,N_6030,N_6235);
nand U8820 (N_8820,N_6092,N_6452);
or U8821 (N_8821,N_6878,N_6245);
or U8822 (N_8822,N_7175,N_5229);
or U8823 (N_8823,N_5813,N_6074);
or U8824 (N_8824,N_6662,N_5877);
and U8825 (N_8825,N_6848,N_7350);
nand U8826 (N_8826,N_7199,N_5709);
and U8827 (N_8827,N_6044,N_5032);
xor U8828 (N_8828,N_7218,N_6914);
and U8829 (N_8829,N_6863,N_5534);
and U8830 (N_8830,N_6992,N_7404);
xnor U8831 (N_8831,N_7052,N_7348);
and U8832 (N_8832,N_5537,N_6558);
nand U8833 (N_8833,N_6703,N_6895);
nor U8834 (N_8834,N_5673,N_6254);
xnor U8835 (N_8835,N_6724,N_7195);
nor U8836 (N_8836,N_5100,N_7076);
and U8837 (N_8837,N_5652,N_6775);
nand U8838 (N_8838,N_7089,N_5968);
nand U8839 (N_8839,N_6709,N_7174);
or U8840 (N_8840,N_5421,N_5582);
xnor U8841 (N_8841,N_7417,N_5226);
or U8842 (N_8842,N_7341,N_7300);
or U8843 (N_8843,N_6542,N_5762);
or U8844 (N_8844,N_6525,N_6313);
xnor U8845 (N_8845,N_5501,N_5970);
and U8846 (N_8846,N_6017,N_6764);
and U8847 (N_8847,N_5921,N_5599);
or U8848 (N_8848,N_5540,N_5125);
or U8849 (N_8849,N_6578,N_5044);
nand U8850 (N_8850,N_5849,N_6594);
nand U8851 (N_8851,N_5248,N_6398);
xor U8852 (N_8852,N_5349,N_6813);
and U8853 (N_8853,N_5653,N_7170);
xnor U8854 (N_8854,N_6735,N_5077);
nor U8855 (N_8855,N_6729,N_6830);
nand U8856 (N_8856,N_5053,N_6056);
nor U8857 (N_8857,N_6422,N_6280);
nor U8858 (N_8858,N_5571,N_6650);
nor U8859 (N_8859,N_7007,N_6823);
and U8860 (N_8860,N_6745,N_6939);
or U8861 (N_8861,N_6386,N_5420);
nor U8862 (N_8862,N_6685,N_6462);
xor U8863 (N_8863,N_5972,N_5277);
nand U8864 (N_8864,N_5602,N_6284);
xnor U8865 (N_8865,N_6683,N_6346);
xor U8866 (N_8866,N_7455,N_6577);
nand U8867 (N_8867,N_5167,N_7405);
nand U8868 (N_8868,N_7295,N_5647);
nand U8869 (N_8869,N_6703,N_6425);
nand U8870 (N_8870,N_6170,N_7499);
or U8871 (N_8871,N_7326,N_5816);
and U8872 (N_8872,N_5360,N_6412);
xnor U8873 (N_8873,N_6209,N_6542);
nor U8874 (N_8874,N_6401,N_6896);
or U8875 (N_8875,N_6411,N_6967);
or U8876 (N_8876,N_6502,N_5715);
or U8877 (N_8877,N_5287,N_7178);
nand U8878 (N_8878,N_5607,N_5285);
and U8879 (N_8879,N_6637,N_5267);
nor U8880 (N_8880,N_7181,N_6163);
xor U8881 (N_8881,N_7446,N_6699);
and U8882 (N_8882,N_7488,N_7394);
or U8883 (N_8883,N_7019,N_6204);
or U8884 (N_8884,N_6955,N_7265);
nor U8885 (N_8885,N_6686,N_5862);
nor U8886 (N_8886,N_6717,N_5264);
nand U8887 (N_8887,N_5710,N_7043);
and U8888 (N_8888,N_7482,N_7438);
or U8889 (N_8889,N_5894,N_5156);
and U8890 (N_8890,N_6857,N_7098);
xnor U8891 (N_8891,N_5770,N_6058);
nand U8892 (N_8892,N_6701,N_6870);
nand U8893 (N_8893,N_6353,N_6669);
and U8894 (N_8894,N_5914,N_5349);
nor U8895 (N_8895,N_6888,N_6325);
nor U8896 (N_8896,N_6582,N_5973);
nor U8897 (N_8897,N_5329,N_5295);
or U8898 (N_8898,N_5829,N_6382);
or U8899 (N_8899,N_7082,N_7077);
nor U8900 (N_8900,N_6283,N_5182);
and U8901 (N_8901,N_7211,N_5703);
and U8902 (N_8902,N_6973,N_6665);
or U8903 (N_8903,N_6321,N_5921);
nand U8904 (N_8904,N_5790,N_7465);
nand U8905 (N_8905,N_6224,N_5684);
nand U8906 (N_8906,N_7479,N_5623);
and U8907 (N_8907,N_5216,N_5615);
or U8908 (N_8908,N_6871,N_6579);
or U8909 (N_8909,N_5409,N_5109);
xor U8910 (N_8910,N_7146,N_7370);
or U8911 (N_8911,N_7044,N_6560);
or U8912 (N_8912,N_5838,N_5663);
nand U8913 (N_8913,N_5771,N_6406);
or U8914 (N_8914,N_6285,N_5724);
or U8915 (N_8915,N_7277,N_5900);
and U8916 (N_8916,N_6078,N_5722);
and U8917 (N_8917,N_6056,N_6946);
or U8918 (N_8918,N_7067,N_5830);
or U8919 (N_8919,N_6009,N_7201);
and U8920 (N_8920,N_7374,N_5279);
xnor U8921 (N_8921,N_5479,N_5338);
or U8922 (N_8922,N_7415,N_7160);
nor U8923 (N_8923,N_5535,N_6677);
xor U8924 (N_8924,N_7039,N_5119);
or U8925 (N_8925,N_5098,N_7300);
or U8926 (N_8926,N_5203,N_5241);
and U8927 (N_8927,N_5037,N_5757);
nand U8928 (N_8928,N_5002,N_7343);
and U8929 (N_8929,N_5284,N_5233);
nand U8930 (N_8930,N_6052,N_6633);
xnor U8931 (N_8931,N_5378,N_6344);
or U8932 (N_8932,N_6722,N_6275);
nand U8933 (N_8933,N_6587,N_6380);
nand U8934 (N_8934,N_6622,N_6479);
nor U8935 (N_8935,N_5054,N_5386);
or U8936 (N_8936,N_5495,N_5069);
nand U8937 (N_8937,N_7290,N_5995);
nand U8938 (N_8938,N_6343,N_5041);
nor U8939 (N_8939,N_6795,N_5358);
xor U8940 (N_8940,N_5046,N_6241);
xnor U8941 (N_8941,N_5848,N_7311);
nand U8942 (N_8942,N_6999,N_7330);
and U8943 (N_8943,N_5973,N_5904);
nor U8944 (N_8944,N_6897,N_5736);
xnor U8945 (N_8945,N_6521,N_5062);
nor U8946 (N_8946,N_7442,N_5373);
nor U8947 (N_8947,N_6252,N_6312);
or U8948 (N_8948,N_7127,N_5595);
and U8949 (N_8949,N_7156,N_6012);
and U8950 (N_8950,N_6510,N_7111);
nand U8951 (N_8951,N_6674,N_7141);
nor U8952 (N_8952,N_7375,N_5472);
or U8953 (N_8953,N_7211,N_6681);
xnor U8954 (N_8954,N_7074,N_6143);
nor U8955 (N_8955,N_5758,N_6166);
xnor U8956 (N_8956,N_6183,N_6453);
nor U8957 (N_8957,N_6972,N_6909);
xnor U8958 (N_8958,N_5376,N_6283);
xor U8959 (N_8959,N_6371,N_5768);
nand U8960 (N_8960,N_7030,N_6758);
xor U8961 (N_8961,N_7259,N_6276);
or U8962 (N_8962,N_6813,N_5908);
nand U8963 (N_8963,N_5736,N_7279);
nor U8964 (N_8964,N_6825,N_6513);
nor U8965 (N_8965,N_6822,N_7002);
nand U8966 (N_8966,N_5021,N_5929);
nand U8967 (N_8967,N_5007,N_5221);
and U8968 (N_8968,N_5623,N_5729);
nand U8969 (N_8969,N_5345,N_5423);
or U8970 (N_8970,N_5636,N_5691);
xnor U8971 (N_8971,N_6615,N_6158);
and U8972 (N_8972,N_6850,N_6233);
or U8973 (N_8973,N_6720,N_5365);
or U8974 (N_8974,N_5961,N_6314);
and U8975 (N_8975,N_7379,N_6562);
xnor U8976 (N_8976,N_7354,N_5677);
nand U8977 (N_8977,N_7135,N_6719);
nor U8978 (N_8978,N_6922,N_5208);
xnor U8979 (N_8979,N_6329,N_5089);
or U8980 (N_8980,N_6348,N_6460);
nand U8981 (N_8981,N_6172,N_6011);
nor U8982 (N_8982,N_5936,N_5788);
xnor U8983 (N_8983,N_6425,N_6438);
nand U8984 (N_8984,N_6725,N_7336);
nand U8985 (N_8985,N_7071,N_6396);
and U8986 (N_8986,N_7013,N_5063);
nor U8987 (N_8987,N_5539,N_5643);
xor U8988 (N_8988,N_5041,N_5129);
nand U8989 (N_8989,N_6555,N_6583);
and U8990 (N_8990,N_5852,N_5925);
nor U8991 (N_8991,N_6994,N_5903);
and U8992 (N_8992,N_7165,N_7229);
xnor U8993 (N_8993,N_5482,N_7041);
and U8994 (N_8994,N_5062,N_6851);
or U8995 (N_8995,N_5776,N_5332);
nor U8996 (N_8996,N_6269,N_5437);
or U8997 (N_8997,N_5643,N_7463);
xor U8998 (N_8998,N_5702,N_6296);
xnor U8999 (N_8999,N_5215,N_6530);
nor U9000 (N_9000,N_5505,N_6426);
xor U9001 (N_9001,N_5478,N_7482);
xnor U9002 (N_9002,N_6625,N_6786);
or U9003 (N_9003,N_6460,N_6202);
or U9004 (N_9004,N_6031,N_5682);
or U9005 (N_9005,N_5773,N_6138);
or U9006 (N_9006,N_7381,N_6044);
xor U9007 (N_9007,N_5451,N_5660);
and U9008 (N_9008,N_5460,N_6224);
or U9009 (N_9009,N_6892,N_6574);
and U9010 (N_9010,N_6618,N_5828);
nor U9011 (N_9011,N_6364,N_6898);
and U9012 (N_9012,N_6905,N_6964);
nor U9013 (N_9013,N_7012,N_5666);
nand U9014 (N_9014,N_7359,N_6135);
and U9015 (N_9015,N_5766,N_6462);
xor U9016 (N_9016,N_6031,N_6228);
or U9017 (N_9017,N_7077,N_5877);
nor U9018 (N_9018,N_6077,N_6140);
xnor U9019 (N_9019,N_5503,N_6917);
nand U9020 (N_9020,N_6884,N_7362);
xnor U9021 (N_9021,N_6202,N_6770);
nor U9022 (N_9022,N_6194,N_6095);
nor U9023 (N_9023,N_6225,N_6612);
nand U9024 (N_9024,N_6852,N_5539);
nor U9025 (N_9025,N_5287,N_7032);
nor U9026 (N_9026,N_6991,N_5922);
nand U9027 (N_9027,N_5055,N_6505);
nor U9028 (N_9028,N_7247,N_6029);
nor U9029 (N_9029,N_7419,N_7096);
nor U9030 (N_9030,N_5693,N_5512);
and U9031 (N_9031,N_7201,N_6277);
and U9032 (N_9032,N_7281,N_6635);
or U9033 (N_9033,N_6925,N_5411);
nor U9034 (N_9034,N_5456,N_6347);
nor U9035 (N_9035,N_5844,N_7373);
nand U9036 (N_9036,N_5689,N_5324);
xor U9037 (N_9037,N_5942,N_5372);
nor U9038 (N_9038,N_7253,N_7236);
xnor U9039 (N_9039,N_7452,N_7073);
and U9040 (N_9040,N_6264,N_5427);
nand U9041 (N_9041,N_5683,N_5235);
or U9042 (N_9042,N_5087,N_5312);
xnor U9043 (N_9043,N_5329,N_6847);
xor U9044 (N_9044,N_6047,N_6213);
xor U9045 (N_9045,N_5442,N_5254);
xor U9046 (N_9046,N_6469,N_5357);
nor U9047 (N_9047,N_7298,N_5827);
nand U9048 (N_9048,N_5499,N_5820);
and U9049 (N_9049,N_5518,N_7200);
nand U9050 (N_9050,N_6375,N_5317);
or U9051 (N_9051,N_6235,N_5130);
nor U9052 (N_9052,N_7107,N_5879);
nor U9053 (N_9053,N_6652,N_6615);
nor U9054 (N_9054,N_5523,N_7453);
nand U9055 (N_9055,N_7228,N_5151);
xnor U9056 (N_9056,N_5786,N_7178);
and U9057 (N_9057,N_5574,N_6258);
nor U9058 (N_9058,N_5051,N_7392);
nand U9059 (N_9059,N_7468,N_7394);
xor U9060 (N_9060,N_6652,N_7330);
or U9061 (N_9061,N_5005,N_5779);
nand U9062 (N_9062,N_7242,N_5769);
nor U9063 (N_9063,N_6800,N_6912);
nand U9064 (N_9064,N_6369,N_5712);
nor U9065 (N_9065,N_6057,N_6665);
nor U9066 (N_9066,N_5355,N_7124);
nor U9067 (N_9067,N_5411,N_6599);
xnor U9068 (N_9068,N_6248,N_6678);
or U9069 (N_9069,N_6421,N_7462);
and U9070 (N_9070,N_6305,N_5471);
nand U9071 (N_9071,N_6254,N_5711);
and U9072 (N_9072,N_5180,N_7016);
or U9073 (N_9073,N_5322,N_5949);
nand U9074 (N_9074,N_5754,N_6022);
nand U9075 (N_9075,N_5430,N_6457);
or U9076 (N_9076,N_5931,N_6181);
or U9077 (N_9077,N_7167,N_7156);
nor U9078 (N_9078,N_5334,N_6156);
nor U9079 (N_9079,N_6649,N_6729);
and U9080 (N_9080,N_5714,N_6661);
or U9081 (N_9081,N_5469,N_6927);
and U9082 (N_9082,N_6054,N_6296);
nor U9083 (N_9083,N_5502,N_5565);
nor U9084 (N_9084,N_5503,N_5895);
or U9085 (N_9085,N_7343,N_6067);
nand U9086 (N_9086,N_5670,N_5718);
or U9087 (N_9087,N_6550,N_7478);
and U9088 (N_9088,N_7316,N_5109);
nand U9089 (N_9089,N_5509,N_6983);
and U9090 (N_9090,N_6337,N_6919);
nor U9091 (N_9091,N_5666,N_6894);
nand U9092 (N_9092,N_6151,N_7435);
nor U9093 (N_9093,N_6849,N_6945);
nand U9094 (N_9094,N_7375,N_5730);
and U9095 (N_9095,N_6069,N_5173);
nand U9096 (N_9096,N_6276,N_7219);
and U9097 (N_9097,N_6293,N_6924);
and U9098 (N_9098,N_5927,N_6803);
nand U9099 (N_9099,N_5800,N_6828);
xor U9100 (N_9100,N_5743,N_5508);
nand U9101 (N_9101,N_6629,N_6475);
and U9102 (N_9102,N_7369,N_5459);
xnor U9103 (N_9103,N_5505,N_5617);
nor U9104 (N_9104,N_6074,N_6594);
xor U9105 (N_9105,N_6873,N_5232);
xor U9106 (N_9106,N_6774,N_6000);
nand U9107 (N_9107,N_6604,N_6507);
nor U9108 (N_9108,N_7288,N_6632);
xor U9109 (N_9109,N_5989,N_6035);
nand U9110 (N_9110,N_5350,N_7342);
nand U9111 (N_9111,N_5446,N_5145);
nor U9112 (N_9112,N_6729,N_5982);
and U9113 (N_9113,N_7244,N_6304);
or U9114 (N_9114,N_5088,N_7251);
and U9115 (N_9115,N_5621,N_6625);
nor U9116 (N_9116,N_7224,N_7305);
or U9117 (N_9117,N_7113,N_5474);
or U9118 (N_9118,N_6295,N_6261);
and U9119 (N_9119,N_6532,N_5001);
nor U9120 (N_9120,N_6971,N_7263);
and U9121 (N_9121,N_6471,N_7072);
or U9122 (N_9122,N_5982,N_6792);
or U9123 (N_9123,N_5685,N_6563);
xnor U9124 (N_9124,N_5318,N_6472);
nor U9125 (N_9125,N_5008,N_7157);
nor U9126 (N_9126,N_5963,N_6477);
xnor U9127 (N_9127,N_7241,N_6813);
or U9128 (N_9128,N_6443,N_7189);
xor U9129 (N_9129,N_5626,N_6616);
and U9130 (N_9130,N_5094,N_6176);
xor U9131 (N_9131,N_5154,N_6992);
xor U9132 (N_9132,N_5509,N_7142);
xnor U9133 (N_9133,N_7443,N_6063);
and U9134 (N_9134,N_5635,N_6220);
xnor U9135 (N_9135,N_6548,N_6609);
nand U9136 (N_9136,N_6367,N_5541);
and U9137 (N_9137,N_5582,N_6342);
xor U9138 (N_9138,N_5984,N_7342);
nand U9139 (N_9139,N_6567,N_6635);
or U9140 (N_9140,N_6040,N_7469);
xnor U9141 (N_9141,N_6198,N_6854);
and U9142 (N_9142,N_5888,N_5592);
nand U9143 (N_9143,N_5303,N_5519);
or U9144 (N_9144,N_5453,N_6994);
nand U9145 (N_9145,N_5609,N_5986);
xnor U9146 (N_9146,N_6544,N_5364);
nand U9147 (N_9147,N_6375,N_7115);
or U9148 (N_9148,N_6475,N_7311);
or U9149 (N_9149,N_6251,N_5063);
nand U9150 (N_9150,N_6142,N_6028);
and U9151 (N_9151,N_6604,N_6497);
and U9152 (N_9152,N_5725,N_5108);
nor U9153 (N_9153,N_5812,N_6559);
and U9154 (N_9154,N_6124,N_5742);
nor U9155 (N_9155,N_5254,N_6675);
nor U9156 (N_9156,N_6319,N_5643);
nor U9157 (N_9157,N_7406,N_7193);
xnor U9158 (N_9158,N_7319,N_5526);
and U9159 (N_9159,N_5599,N_5581);
or U9160 (N_9160,N_6652,N_7248);
nor U9161 (N_9161,N_6787,N_6638);
and U9162 (N_9162,N_6954,N_6851);
nand U9163 (N_9163,N_5472,N_7236);
nand U9164 (N_9164,N_6278,N_6895);
nor U9165 (N_9165,N_6332,N_7016);
nand U9166 (N_9166,N_5723,N_6051);
or U9167 (N_9167,N_5644,N_5627);
or U9168 (N_9168,N_5203,N_6474);
xor U9169 (N_9169,N_5879,N_7402);
nor U9170 (N_9170,N_5220,N_6884);
nor U9171 (N_9171,N_6334,N_5643);
nor U9172 (N_9172,N_7400,N_7446);
and U9173 (N_9173,N_5240,N_7280);
xnor U9174 (N_9174,N_5380,N_5672);
nand U9175 (N_9175,N_5117,N_7073);
nor U9176 (N_9176,N_6662,N_6416);
nand U9177 (N_9177,N_6205,N_5114);
and U9178 (N_9178,N_6247,N_7201);
nand U9179 (N_9179,N_5521,N_6484);
or U9180 (N_9180,N_5196,N_6086);
xor U9181 (N_9181,N_6112,N_6931);
nand U9182 (N_9182,N_6866,N_5135);
nand U9183 (N_9183,N_6664,N_5635);
and U9184 (N_9184,N_5043,N_6238);
and U9185 (N_9185,N_6119,N_5844);
xnor U9186 (N_9186,N_5694,N_6857);
nor U9187 (N_9187,N_5107,N_5706);
nor U9188 (N_9188,N_5381,N_6462);
xnor U9189 (N_9189,N_5678,N_6159);
nand U9190 (N_9190,N_6943,N_6368);
nand U9191 (N_9191,N_6518,N_5921);
or U9192 (N_9192,N_5511,N_7046);
nor U9193 (N_9193,N_6534,N_7251);
nand U9194 (N_9194,N_6651,N_6777);
and U9195 (N_9195,N_6106,N_5221);
nor U9196 (N_9196,N_7341,N_7136);
and U9197 (N_9197,N_5277,N_7273);
xnor U9198 (N_9198,N_6051,N_7032);
xnor U9199 (N_9199,N_7294,N_5961);
xnor U9200 (N_9200,N_5088,N_5194);
nand U9201 (N_9201,N_6057,N_5490);
or U9202 (N_9202,N_7247,N_7291);
and U9203 (N_9203,N_6514,N_6938);
nand U9204 (N_9204,N_5723,N_6751);
nand U9205 (N_9205,N_6096,N_7434);
nand U9206 (N_9206,N_5543,N_7285);
nand U9207 (N_9207,N_7237,N_5047);
or U9208 (N_9208,N_5181,N_6669);
nand U9209 (N_9209,N_5808,N_6799);
xnor U9210 (N_9210,N_6829,N_5091);
nor U9211 (N_9211,N_7127,N_7483);
and U9212 (N_9212,N_7481,N_6197);
and U9213 (N_9213,N_7113,N_6254);
xnor U9214 (N_9214,N_6892,N_6918);
nand U9215 (N_9215,N_6786,N_6885);
or U9216 (N_9216,N_5576,N_5126);
nand U9217 (N_9217,N_6826,N_5685);
nor U9218 (N_9218,N_7460,N_6022);
nand U9219 (N_9219,N_7239,N_6763);
or U9220 (N_9220,N_7206,N_7169);
nand U9221 (N_9221,N_7390,N_7454);
xnor U9222 (N_9222,N_5111,N_6248);
nand U9223 (N_9223,N_6754,N_6138);
and U9224 (N_9224,N_6768,N_5556);
and U9225 (N_9225,N_5262,N_5198);
and U9226 (N_9226,N_5754,N_6307);
nand U9227 (N_9227,N_5905,N_5813);
xor U9228 (N_9228,N_6473,N_6155);
nor U9229 (N_9229,N_6260,N_7222);
and U9230 (N_9230,N_5815,N_5811);
nand U9231 (N_9231,N_5763,N_5424);
and U9232 (N_9232,N_6610,N_5095);
or U9233 (N_9233,N_5347,N_5407);
nand U9234 (N_9234,N_6991,N_6792);
nand U9235 (N_9235,N_5823,N_6029);
nand U9236 (N_9236,N_6858,N_5600);
xor U9237 (N_9237,N_6775,N_6049);
xor U9238 (N_9238,N_6049,N_5379);
and U9239 (N_9239,N_5538,N_5521);
xor U9240 (N_9240,N_5334,N_6427);
nor U9241 (N_9241,N_5027,N_5335);
xor U9242 (N_9242,N_5229,N_5827);
nor U9243 (N_9243,N_6401,N_5446);
xor U9244 (N_9244,N_7122,N_7068);
xnor U9245 (N_9245,N_7101,N_5846);
nor U9246 (N_9246,N_5093,N_5670);
nand U9247 (N_9247,N_5164,N_7244);
nand U9248 (N_9248,N_5009,N_6681);
and U9249 (N_9249,N_5620,N_6128);
xnor U9250 (N_9250,N_6775,N_5412);
or U9251 (N_9251,N_6026,N_6292);
or U9252 (N_9252,N_5726,N_6833);
nand U9253 (N_9253,N_7288,N_6886);
and U9254 (N_9254,N_5187,N_7470);
and U9255 (N_9255,N_7409,N_5590);
nor U9256 (N_9256,N_7204,N_6938);
or U9257 (N_9257,N_6581,N_5951);
xor U9258 (N_9258,N_6870,N_6244);
xnor U9259 (N_9259,N_6318,N_6615);
nor U9260 (N_9260,N_5124,N_6879);
or U9261 (N_9261,N_6256,N_7091);
nor U9262 (N_9262,N_5209,N_6335);
xnor U9263 (N_9263,N_5746,N_5923);
xnor U9264 (N_9264,N_7468,N_6655);
nand U9265 (N_9265,N_5903,N_7090);
or U9266 (N_9266,N_6929,N_5497);
nand U9267 (N_9267,N_5275,N_5337);
nor U9268 (N_9268,N_5246,N_6700);
xnor U9269 (N_9269,N_5894,N_5776);
nor U9270 (N_9270,N_6746,N_5630);
nor U9271 (N_9271,N_6897,N_5139);
nand U9272 (N_9272,N_6599,N_5788);
nand U9273 (N_9273,N_6287,N_5585);
xor U9274 (N_9274,N_7101,N_7179);
nand U9275 (N_9275,N_6671,N_7477);
xnor U9276 (N_9276,N_6552,N_5155);
and U9277 (N_9277,N_6916,N_5404);
nand U9278 (N_9278,N_7317,N_7047);
nand U9279 (N_9279,N_6058,N_6299);
nor U9280 (N_9280,N_5775,N_5727);
nand U9281 (N_9281,N_6599,N_7416);
and U9282 (N_9282,N_6589,N_7327);
xor U9283 (N_9283,N_6127,N_6457);
nand U9284 (N_9284,N_5375,N_6095);
xnor U9285 (N_9285,N_7124,N_5385);
nand U9286 (N_9286,N_7338,N_6892);
and U9287 (N_9287,N_6578,N_5698);
and U9288 (N_9288,N_6158,N_5691);
xnor U9289 (N_9289,N_6595,N_5524);
xor U9290 (N_9290,N_7109,N_6107);
or U9291 (N_9291,N_7358,N_6532);
or U9292 (N_9292,N_5620,N_5833);
nor U9293 (N_9293,N_5474,N_5270);
or U9294 (N_9294,N_5147,N_6065);
xnor U9295 (N_9295,N_7204,N_5000);
nand U9296 (N_9296,N_6870,N_7183);
or U9297 (N_9297,N_6437,N_5456);
or U9298 (N_9298,N_5597,N_5281);
nand U9299 (N_9299,N_5886,N_5266);
nor U9300 (N_9300,N_6339,N_7167);
nor U9301 (N_9301,N_7291,N_6563);
xor U9302 (N_9302,N_6893,N_7227);
nand U9303 (N_9303,N_7475,N_6668);
nand U9304 (N_9304,N_6257,N_6101);
nor U9305 (N_9305,N_6347,N_7174);
nand U9306 (N_9306,N_7265,N_5476);
and U9307 (N_9307,N_7360,N_6759);
and U9308 (N_9308,N_5224,N_5919);
or U9309 (N_9309,N_5892,N_5385);
nand U9310 (N_9310,N_6955,N_6077);
or U9311 (N_9311,N_5509,N_6660);
nand U9312 (N_9312,N_6845,N_7241);
nor U9313 (N_9313,N_7084,N_6668);
or U9314 (N_9314,N_7467,N_7382);
or U9315 (N_9315,N_5699,N_6233);
nor U9316 (N_9316,N_5579,N_6078);
and U9317 (N_9317,N_5061,N_5553);
and U9318 (N_9318,N_7149,N_7153);
nor U9319 (N_9319,N_6450,N_6014);
xor U9320 (N_9320,N_7404,N_5577);
nand U9321 (N_9321,N_6096,N_5029);
nor U9322 (N_9322,N_6082,N_6655);
nand U9323 (N_9323,N_6984,N_6860);
and U9324 (N_9324,N_7186,N_7285);
xnor U9325 (N_9325,N_6560,N_6815);
xor U9326 (N_9326,N_5774,N_7338);
and U9327 (N_9327,N_7307,N_5554);
and U9328 (N_9328,N_6700,N_7449);
or U9329 (N_9329,N_7025,N_5925);
and U9330 (N_9330,N_5128,N_7301);
nor U9331 (N_9331,N_6290,N_6704);
nor U9332 (N_9332,N_6235,N_6398);
nor U9333 (N_9333,N_6963,N_5650);
or U9334 (N_9334,N_6584,N_6009);
nand U9335 (N_9335,N_6585,N_5385);
and U9336 (N_9336,N_5508,N_7252);
nand U9337 (N_9337,N_6086,N_6905);
and U9338 (N_9338,N_7361,N_5090);
xor U9339 (N_9339,N_5359,N_6658);
nand U9340 (N_9340,N_7303,N_5389);
and U9341 (N_9341,N_5950,N_6897);
or U9342 (N_9342,N_5685,N_7454);
and U9343 (N_9343,N_6616,N_5827);
nand U9344 (N_9344,N_5775,N_5625);
nand U9345 (N_9345,N_6362,N_7244);
nor U9346 (N_9346,N_5008,N_5098);
nand U9347 (N_9347,N_6223,N_7290);
and U9348 (N_9348,N_7434,N_6462);
and U9349 (N_9349,N_5386,N_5039);
nand U9350 (N_9350,N_5831,N_5980);
and U9351 (N_9351,N_5424,N_6737);
and U9352 (N_9352,N_5578,N_6447);
nand U9353 (N_9353,N_5885,N_6652);
or U9354 (N_9354,N_7009,N_7183);
and U9355 (N_9355,N_6491,N_5612);
and U9356 (N_9356,N_6472,N_6358);
xnor U9357 (N_9357,N_6581,N_5980);
and U9358 (N_9358,N_6420,N_7152);
and U9359 (N_9359,N_6136,N_6446);
nand U9360 (N_9360,N_5640,N_7084);
xor U9361 (N_9361,N_6173,N_5136);
xnor U9362 (N_9362,N_6131,N_6728);
or U9363 (N_9363,N_7089,N_7338);
nor U9364 (N_9364,N_6862,N_7085);
xnor U9365 (N_9365,N_6112,N_6738);
and U9366 (N_9366,N_6925,N_6601);
or U9367 (N_9367,N_5380,N_7453);
nor U9368 (N_9368,N_6972,N_7321);
nand U9369 (N_9369,N_7103,N_7227);
and U9370 (N_9370,N_5704,N_6428);
and U9371 (N_9371,N_6096,N_6986);
or U9372 (N_9372,N_5632,N_5785);
xor U9373 (N_9373,N_5396,N_5357);
or U9374 (N_9374,N_6326,N_5680);
xnor U9375 (N_9375,N_6344,N_6728);
or U9376 (N_9376,N_7356,N_5612);
and U9377 (N_9377,N_7124,N_7081);
and U9378 (N_9378,N_6803,N_6813);
nand U9379 (N_9379,N_5093,N_5005);
xor U9380 (N_9380,N_7074,N_6107);
xor U9381 (N_9381,N_5696,N_5142);
or U9382 (N_9382,N_7473,N_5106);
and U9383 (N_9383,N_6150,N_6448);
and U9384 (N_9384,N_5677,N_6668);
nand U9385 (N_9385,N_5248,N_6491);
nor U9386 (N_9386,N_6764,N_5668);
or U9387 (N_9387,N_7222,N_6078);
xor U9388 (N_9388,N_7106,N_5094);
nand U9389 (N_9389,N_6719,N_7111);
xor U9390 (N_9390,N_6766,N_7390);
or U9391 (N_9391,N_5686,N_6790);
xor U9392 (N_9392,N_7438,N_5119);
nand U9393 (N_9393,N_7316,N_7026);
nor U9394 (N_9394,N_6698,N_5609);
xnor U9395 (N_9395,N_5532,N_6877);
and U9396 (N_9396,N_5674,N_6096);
nor U9397 (N_9397,N_5964,N_7231);
xnor U9398 (N_9398,N_6723,N_5437);
nand U9399 (N_9399,N_7207,N_5306);
or U9400 (N_9400,N_5658,N_6371);
nand U9401 (N_9401,N_5806,N_7379);
nor U9402 (N_9402,N_5903,N_7399);
nand U9403 (N_9403,N_5588,N_5986);
and U9404 (N_9404,N_5755,N_6118);
xor U9405 (N_9405,N_5127,N_6349);
and U9406 (N_9406,N_6998,N_5771);
or U9407 (N_9407,N_6936,N_6383);
xor U9408 (N_9408,N_6062,N_6707);
and U9409 (N_9409,N_5078,N_6023);
nand U9410 (N_9410,N_6240,N_6539);
xor U9411 (N_9411,N_6094,N_5159);
xnor U9412 (N_9412,N_6747,N_5918);
or U9413 (N_9413,N_6663,N_6461);
or U9414 (N_9414,N_7073,N_5974);
xor U9415 (N_9415,N_6472,N_6244);
and U9416 (N_9416,N_6286,N_7493);
nand U9417 (N_9417,N_6188,N_5079);
and U9418 (N_9418,N_5335,N_5619);
and U9419 (N_9419,N_5824,N_5869);
nor U9420 (N_9420,N_6098,N_6379);
xor U9421 (N_9421,N_6968,N_7307);
nand U9422 (N_9422,N_6701,N_5213);
or U9423 (N_9423,N_7220,N_5390);
nand U9424 (N_9424,N_6884,N_7397);
nor U9425 (N_9425,N_5723,N_6068);
nor U9426 (N_9426,N_5791,N_5941);
xnor U9427 (N_9427,N_6468,N_7191);
xor U9428 (N_9428,N_6121,N_6099);
nand U9429 (N_9429,N_7274,N_5051);
xor U9430 (N_9430,N_6474,N_6492);
or U9431 (N_9431,N_7184,N_6286);
xnor U9432 (N_9432,N_7245,N_5201);
xnor U9433 (N_9433,N_6580,N_5897);
xor U9434 (N_9434,N_6538,N_6026);
nor U9435 (N_9435,N_6401,N_5256);
or U9436 (N_9436,N_7171,N_5103);
nor U9437 (N_9437,N_5887,N_7301);
or U9438 (N_9438,N_6396,N_7291);
or U9439 (N_9439,N_5369,N_6264);
and U9440 (N_9440,N_6234,N_5635);
nor U9441 (N_9441,N_7422,N_6056);
xor U9442 (N_9442,N_6894,N_5902);
nand U9443 (N_9443,N_5322,N_5474);
or U9444 (N_9444,N_5194,N_6394);
and U9445 (N_9445,N_5259,N_6736);
nand U9446 (N_9446,N_6404,N_7098);
and U9447 (N_9447,N_6707,N_6757);
nand U9448 (N_9448,N_6512,N_5760);
xnor U9449 (N_9449,N_7236,N_7231);
and U9450 (N_9450,N_5926,N_5276);
xnor U9451 (N_9451,N_6247,N_6313);
nor U9452 (N_9452,N_5648,N_6983);
nor U9453 (N_9453,N_5040,N_6828);
nor U9454 (N_9454,N_7067,N_5366);
xor U9455 (N_9455,N_5220,N_5419);
xnor U9456 (N_9456,N_6726,N_6668);
xor U9457 (N_9457,N_6199,N_5783);
and U9458 (N_9458,N_6095,N_7410);
nand U9459 (N_9459,N_7254,N_6116);
nand U9460 (N_9460,N_5053,N_6092);
and U9461 (N_9461,N_5993,N_7135);
or U9462 (N_9462,N_5329,N_5134);
or U9463 (N_9463,N_5899,N_6004);
and U9464 (N_9464,N_7000,N_6739);
or U9465 (N_9465,N_5029,N_6849);
and U9466 (N_9466,N_5527,N_7230);
nor U9467 (N_9467,N_5477,N_6850);
xnor U9468 (N_9468,N_6354,N_5344);
and U9469 (N_9469,N_6509,N_5072);
nor U9470 (N_9470,N_6890,N_5056);
or U9471 (N_9471,N_6534,N_6231);
or U9472 (N_9472,N_7135,N_7257);
and U9473 (N_9473,N_6239,N_6689);
and U9474 (N_9474,N_6393,N_6744);
and U9475 (N_9475,N_6068,N_6292);
xnor U9476 (N_9476,N_5816,N_5783);
nand U9477 (N_9477,N_6581,N_6485);
nor U9478 (N_9478,N_6667,N_6697);
nand U9479 (N_9479,N_5667,N_7292);
nand U9480 (N_9480,N_6616,N_5838);
nor U9481 (N_9481,N_6125,N_5854);
and U9482 (N_9482,N_5749,N_5710);
nand U9483 (N_9483,N_6429,N_7070);
and U9484 (N_9484,N_7362,N_5339);
or U9485 (N_9485,N_7268,N_7178);
and U9486 (N_9486,N_5655,N_5026);
nor U9487 (N_9487,N_5552,N_6811);
nand U9488 (N_9488,N_5991,N_6637);
nor U9489 (N_9489,N_5097,N_5399);
nor U9490 (N_9490,N_5051,N_6878);
or U9491 (N_9491,N_6072,N_5338);
xnor U9492 (N_9492,N_6735,N_7275);
nor U9493 (N_9493,N_6224,N_5280);
or U9494 (N_9494,N_6454,N_6693);
and U9495 (N_9495,N_5249,N_6220);
and U9496 (N_9496,N_5194,N_7380);
nor U9497 (N_9497,N_6277,N_6608);
nor U9498 (N_9498,N_7014,N_6541);
nand U9499 (N_9499,N_6390,N_5685);
and U9500 (N_9500,N_5386,N_6651);
nor U9501 (N_9501,N_5418,N_6767);
xor U9502 (N_9502,N_5421,N_5019);
nor U9503 (N_9503,N_5722,N_7191);
and U9504 (N_9504,N_6987,N_6107);
nor U9505 (N_9505,N_6079,N_6471);
xor U9506 (N_9506,N_6877,N_7208);
xnor U9507 (N_9507,N_6655,N_6596);
nor U9508 (N_9508,N_7146,N_6873);
nor U9509 (N_9509,N_6971,N_6074);
and U9510 (N_9510,N_5745,N_7033);
nor U9511 (N_9511,N_7330,N_6863);
nand U9512 (N_9512,N_5133,N_6383);
or U9513 (N_9513,N_6518,N_5140);
and U9514 (N_9514,N_6258,N_5881);
nand U9515 (N_9515,N_6927,N_5359);
or U9516 (N_9516,N_5217,N_5848);
or U9517 (N_9517,N_6212,N_5415);
nand U9518 (N_9518,N_5741,N_5675);
or U9519 (N_9519,N_6402,N_6001);
nand U9520 (N_9520,N_6382,N_5247);
and U9521 (N_9521,N_6440,N_6411);
and U9522 (N_9522,N_6915,N_5990);
or U9523 (N_9523,N_6584,N_5974);
nor U9524 (N_9524,N_6988,N_5878);
xor U9525 (N_9525,N_7261,N_6900);
nor U9526 (N_9526,N_5809,N_6376);
nand U9527 (N_9527,N_7145,N_7466);
nand U9528 (N_9528,N_5825,N_5813);
or U9529 (N_9529,N_6829,N_5240);
xnor U9530 (N_9530,N_5823,N_6396);
and U9531 (N_9531,N_6421,N_6563);
nor U9532 (N_9532,N_7417,N_7141);
and U9533 (N_9533,N_7181,N_7414);
and U9534 (N_9534,N_6027,N_5807);
xor U9535 (N_9535,N_5630,N_5642);
or U9536 (N_9536,N_6245,N_5044);
nor U9537 (N_9537,N_6465,N_6411);
nand U9538 (N_9538,N_5670,N_7334);
or U9539 (N_9539,N_5068,N_6695);
or U9540 (N_9540,N_5167,N_6972);
or U9541 (N_9541,N_5055,N_7123);
nor U9542 (N_9542,N_5921,N_5878);
or U9543 (N_9543,N_5868,N_7428);
or U9544 (N_9544,N_6902,N_5593);
or U9545 (N_9545,N_6632,N_6125);
nor U9546 (N_9546,N_5754,N_6681);
and U9547 (N_9547,N_5772,N_6773);
xnor U9548 (N_9548,N_5563,N_6472);
nor U9549 (N_9549,N_7369,N_5900);
xor U9550 (N_9550,N_5090,N_6057);
and U9551 (N_9551,N_6594,N_5216);
nand U9552 (N_9552,N_5110,N_5872);
xor U9553 (N_9553,N_5161,N_5707);
xnor U9554 (N_9554,N_5845,N_6947);
xor U9555 (N_9555,N_7126,N_6161);
and U9556 (N_9556,N_5220,N_5997);
or U9557 (N_9557,N_7214,N_6166);
and U9558 (N_9558,N_5612,N_6003);
nor U9559 (N_9559,N_7470,N_7217);
nand U9560 (N_9560,N_5499,N_6917);
or U9561 (N_9561,N_6213,N_5426);
nand U9562 (N_9562,N_6032,N_7466);
and U9563 (N_9563,N_6106,N_6940);
nand U9564 (N_9564,N_6075,N_6012);
and U9565 (N_9565,N_5585,N_7253);
and U9566 (N_9566,N_6661,N_7391);
nand U9567 (N_9567,N_5419,N_6744);
xnor U9568 (N_9568,N_5416,N_7076);
and U9569 (N_9569,N_6939,N_5013);
nand U9570 (N_9570,N_6104,N_5818);
nor U9571 (N_9571,N_5348,N_6118);
or U9572 (N_9572,N_6329,N_5601);
or U9573 (N_9573,N_7361,N_5220);
xnor U9574 (N_9574,N_7487,N_5982);
or U9575 (N_9575,N_5451,N_5078);
nand U9576 (N_9576,N_5003,N_7066);
nor U9577 (N_9577,N_7071,N_5025);
and U9578 (N_9578,N_5146,N_5332);
nand U9579 (N_9579,N_6590,N_6239);
xor U9580 (N_9580,N_6178,N_5439);
nand U9581 (N_9581,N_7397,N_7243);
xnor U9582 (N_9582,N_6362,N_7078);
nand U9583 (N_9583,N_6400,N_6425);
and U9584 (N_9584,N_6315,N_6370);
nand U9585 (N_9585,N_5290,N_6601);
xnor U9586 (N_9586,N_5764,N_5646);
nand U9587 (N_9587,N_6681,N_7460);
xnor U9588 (N_9588,N_6022,N_5037);
xnor U9589 (N_9589,N_7380,N_6024);
xnor U9590 (N_9590,N_7006,N_6387);
nand U9591 (N_9591,N_5896,N_7463);
xnor U9592 (N_9592,N_6670,N_6283);
nor U9593 (N_9593,N_5992,N_7480);
nor U9594 (N_9594,N_5334,N_5950);
nand U9595 (N_9595,N_5471,N_5742);
or U9596 (N_9596,N_6474,N_5868);
nor U9597 (N_9597,N_5657,N_5302);
and U9598 (N_9598,N_6029,N_5925);
nand U9599 (N_9599,N_5059,N_6480);
nand U9600 (N_9600,N_5790,N_5346);
or U9601 (N_9601,N_5754,N_6528);
and U9602 (N_9602,N_7043,N_7459);
nor U9603 (N_9603,N_6170,N_7342);
xnor U9604 (N_9604,N_6196,N_5884);
and U9605 (N_9605,N_6394,N_5871);
nand U9606 (N_9606,N_5437,N_7389);
and U9607 (N_9607,N_6863,N_5317);
nand U9608 (N_9608,N_5101,N_6548);
nand U9609 (N_9609,N_7411,N_5182);
and U9610 (N_9610,N_5990,N_5308);
or U9611 (N_9611,N_6525,N_6786);
nand U9612 (N_9612,N_7036,N_5636);
nor U9613 (N_9613,N_5313,N_5044);
or U9614 (N_9614,N_5235,N_7140);
nand U9615 (N_9615,N_5005,N_5249);
xor U9616 (N_9616,N_6807,N_7048);
nor U9617 (N_9617,N_5828,N_7029);
and U9618 (N_9618,N_6343,N_6474);
nand U9619 (N_9619,N_7089,N_7067);
xor U9620 (N_9620,N_6494,N_6360);
nand U9621 (N_9621,N_5327,N_6922);
nor U9622 (N_9622,N_6373,N_6849);
nor U9623 (N_9623,N_6444,N_7081);
nor U9624 (N_9624,N_7456,N_6343);
or U9625 (N_9625,N_5904,N_5125);
or U9626 (N_9626,N_7359,N_7440);
nor U9627 (N_9627,N_7187,N_6262);
or U9628 (N_9628,N_5413,N_6109);
nand U9629 (N_9629,N_6640,N_7332);
and U9630 (N_9630,N_6694,N_5599);
xor U9631 (N_9631,N_5889,N_6664);
or U9632 (N_9632,N_7122,N_5300);
and U9633 (N_9633,N_5647,N_5956);
nor U9634 (N_9634,N_6225,N_5256);
or U9635 (N_9635,N_6379,N_6091);
xnor U9636 (N_9636,N_5684,N_7267);
and U9637 (N_9637,N_5314,N_7437);
and U9638 (N_9638,N_5699,N_5296);
nor U9639 (N_9639,N_5432,N_6077);
xnor U9640 (N_9640,N_5935,N_5013);
nand U9641 (N_9641,N_5769,N_5353);
xor U9642 (N_9642,N_6643,N_5334);
xnor U9643 (N_9643,N_7290,N_6475);
and U9644 (N_9644,N_7346,N_6173);
or U9645 (N_9645,N_6429,N_6290);
nor U9646 (N_9646,N_6353,N_5391);
or U9647 (N_9647,N_5538,N_6087);
xnor U9648 (N_9648,N_5661,N_5349);
nand U9649 (N_9649,N_7146,N_6332);
and U9650 (N_9650,N_5969,N_5057);
nor U9651 (N_9651,N_5401,N_6564);
nand U9652 (N_9652,N_7462,N_6650);
and U9653 (N_9653,N_5006,N_6628);
and U9654 (N_9654,N_7133,N_6123);
or U9655 (N_9655,N_5214,N_7469);
nand U9656 (N_9656,N_6233,N_7482);
and U9657 (N_9657,N_6318,N_5045);
or U9658 (N_9658,N_5686,N_6247);
nor U9659 (N_9659,N_7103,N_5777);
and U9660 (N_9660,N_5700,N_5510);
nor U9661 (N_9661,N_5978,N_5059);
xnor U9662 (N_9662,N_7200,N_7108);
nor U9663 (N_9663,N_5622,N_5361);
xnor U9664 (N_9664,N_5901,N_7283);
nor U9665 (N_9665,N_5914,N_6934);
xnor U9666 (N_9666,N_7009,N_6570);
nand U9667 (N_9667,N_6868,N_6873);
xnor U9668 (N_9668,N_6915,N_5125);
and U9669 (N_9669,N_5080,N_6793);
and U9670 (N_9670,N_6996,N_5269);
nand U9671 (N_9671,N_6208,N_7313);
and U9672 (N_9672,N_5910,N_6449);
or U9673 (N_9673,N_7027,N_6657);
and U9674 (N_9674,N_6935,N_6859);
xnor U9675 (N_9675,N_5007,N_7333);
or U9676 (N_9676,N_7332,N_7361);
or U9677 (N_9677,N_6540,N_6583);
nand U9678 (N_9678,N_6277,N_6264);
nor U9679 (N_9679,N_5306,N_5118);
or U9680 (N_9680,N_7290,N_6203);
or U9681 (N_9681,N_5913,N_5036);
nand U9682 (N_9682,N_7415,N_5124);
nand U9683 (N_9683,N_5734,N_6228);
xor U9684 (N_9684,N_6604,N_5180);
nand U9685 (N_9685,N_6046,N_7371);
or U9686 (N_9686,N_7409,N_5527);
nor U9687 (N_9687,N_5571,N_5188);
or U9688 (N_9688,N_5461,N_5391);
or U9689 (N_9689,N_5484,N_5190);
nor U9690 (N_9690,N_6599,N_6297);
xnor U9691 (N_9691,N_7247,N_5962);
nor U9692 (N_9692,N_7399,N_7197);
or U9693 (N_9693,N_5939,N_5020);
or U9694 (N_9694,N_6574,N_7400);
nor U9695 (N_9695,N_6628,N_6085);
nand U9696 (N_9696,N_6956,N_6368);
nor U9697 (N_9697,N_7393,N_6371);
and U9698 (N_9698,N_5042,N_5113);
nor U9699 (N_9699,N_5037,N_6380);
nand U9700 (N_9700,N_5129,N_7195);
or U9701 (N_9701,N_5786,N_7027);
xnor U9702 (N_9702,N_5531,N_5573);
nand U9703 (N_9703,N_6774,N_6885);
and U9704 (N_9704,N_7077,N_5713);
and U9705 (N_9705,N_6420,N_5708);
and U9706 (N_9706,N_7139,N_6921);
xor U9707 (N_9707,N_6953,N_5024);
or U9708 (N_9708,N_7146,N_7396);
and U9709 (N_9709,N_7099,N_7472);
or U9710 (N_9710,N_7153,N_6899);
and U9711 (N_9711,N_5005,N_6747);
or U9712 (N_9712,N_7238,N_5257);
xor U9713 (N_9713,N_5636,N_5771);
and U9714 (N_9714,N_5930,N_7085);
xnor U9715 (N_9715,N_7369,N_5629);
and U9716 (N_9716,N_5898,N_7497);
or U9717 (N_9717,N_6580,N_5017);
xnor U9718 (N_9718,N_5818,N_5343);
or U9719 (N_9719,N_7324,N_6549);
xnor U9720 (N_9720,N_7032,N_6480);
nand U9721 (N_9721,N_6925,N_6285);
or U9722 (N_9722,N_7309,N_6359);
or U9723 (N_9723,N_5260,N_6130);
nor U9724 (N_9724,N_5107,N_5265);
nand U9725 (N_9725,N_5429,N_6954);
nand U9726 (N_9726,N_5425,N_5140);
nor U9727 (N_9727,N_5395,N_6249);
xor U9728 (N_9728,N_7055,N_6329);
nand U9729 (N_9729,N_6223,N_6614);
nand U9730 (N_9730,N_5994,N_5703);
nor U9731 (N_9731,N_6095,N_5379);
or U9732 (N_9732,N_5134,N_5005);
nor U9733 (N_9733,N_6152,N_6083);
xnor U9734 (N_9734,N_7214,N_5255);
or U9735 (N_9735,N_7287,N_6209);
and U9736 (N_9736,N_5558,N_5178);
and U9737 (N_9737,N_6502,N_5411);
xnor U9738 (N_9738,N_7006,N_5706);
nand U9739 (N_9739,N_6547,N_5016);
or U9740 (N_9740,N_5141,N_6097);
or U9741 (N_9741,N_6900,N_5512);
and U9742 (N_9742,N_5028,N_7277);
xnor U9743 (N_9743,N_7021,N_6968);
xnor U9744 (N_9744,N_5805,N_6730);
or U9745 (N_9745,N_5834,N_5450);
nand U9746 (N_9746,N_7330,N_5320);
and U9747 (N_9747,N_6006,N_6747);
nand U9748 (N_9748,N_5168,N_6599);
nor U9749 (N_9749,N_7017,N_7355);
xor U9750 (N_9750,N_5971,N_6088);
or U9751 (N_9751,N_6593,N_5439);
and U9752 (N_9752,N_6798,N_5398);
nand U9753 (N_9753,N_5601,N_5929);
xor U9754 (N_9754,N_6008,N_7148);
xor U9755 (N_9755,N_5809,N_6658);
xor U9756 (N_9756,N_5820,N_7239);
or U9757 (N_9757,N_7245,N_5814);
or U9758 (N_9758,N_7246,N_5197);
and U9759 (N_9759,N_7032,N_7037);
nand U9760 (N_9760,N_6440,N_6079);
and U9761 (N_9761,N_7299,N_6628);
xnor U9762 (N_9762,N_7429,N_6778);
xor U9763 (N_9763,N_7179,N_6442);
and U9764 (N_9764,N_6499,N_5266);
nor U9765 (N_9765,N_6983,N_5883);
or U9766 (N_9766,N_6877,N_5460);
nor U9767 (N_9767,N_5723,N_6261);
nor U9768 (N_9768,N_6932,N_6915);
xnor U9769 (N_9769,N_6449,N_7237);
xnor U9770 (N_9770,N_6954,N_6559);
xnor U9771 (N_9771,N_6462,N_6976);
nor U9772 (N_9772,N_7303,N_6870);
nand U9773 (N_9773,N_6601,N_7356);
nor U9774 (N_9774,N_6177,N_7359);
nor U9775 (N_9775,N_5341,N_6502);
nand U9776 (N_9776,N_6889,N_5668);
and U9777 (N_9777,N_5041,N_7403);
and U9778 (N_9778,N_6233,N_6290);
xnor U9779 (N_9779,N_5989,N_5533);
xor U9780 (N_9780,N_5260,N_7136);
or U9781 (N_9781,N_7264,N_5104);
nor U9782 (N_9782,N_6897,N_6250);
nand U9783 (N_9783,N_6074,N_6983);
or U9784 (N_9784,N_6099,N_5128);
or U9785 (N_9785,N_5317,N_6869);
and U9786 (N_9786,N_6718,N_6598);
nor U9787 (N_9787,N_6999,N_6199);
xor U9788 (N_9788,N_5843,N_5821);
nor U9789 (N_9789,N_6241,N_5188);
or U9790 (N_9790,N_6855,N_5627);
or U9791 (N_9791,N_5852,N_5995);
and U9792 (N_9792,N_7493,N_5822);
or U9793 (N_9793,N_7151,N_5072);
nand U9794 (N_9794,N_5560,N_6867);
nand U9795 (N_9795,N_6085,N_5143);
nand U9796 (N_9796,N_5202,N_5799);
nor U9797 (N_9797,N_6401,N_5456);
or U9798 (N_9798,N_6359,N_6220);
xnor U9799 (N_9799,N_5992,N_7151);
or U9800 (N_9800,N_6741,N_5994);
or U9801 (N_9801,N_6405,N_5251);
and U9802 (N_9802,N_5274,N_6842);
and U9803 (N_9803,N_5350,N_6979);
nor U9804 (N_9804,N_6893,N_7476);
and U9805 (N_9805,N_7289,N_6533);
nand U9806 (N_9806,N_6039,N_7255);
and U9807 (N_9807,N_6810,N_6585);
xor U9808 (N_9808,N_5784,N_6963);
xor U9809 (N_9809,N_6152,N_6449);
nand U9810 (N_9810,N_7032,N_7242);
or U9811 (N_9811,N_6950,N_7469);
xor U9812 (N_9812,N_5770,N_5191);
or U9813 (N_9813,N_5017,N_5610);
or U9814 (N_9814,N_5908,N_5014);
or U9815 (N_9815,N_6563,N_6095);
nor U9816 (N_9816,N_5081,N_6129);
and U9817 (N_9817,N_6635,N_7371);
nor U9818 (N_9818,N_6442,N_6009);
xor U9819 (N_9819,N_6494,N_6466);
xnor U9820 (N_9820,N_7159,N_7337);
and U9821 (N_9821,N_6646,N_7154);
and U9822 (N_9822,N_7091,N_6340);
and U9823 (N_9823,N_5533,N_7408);
or U9824 (N_9824,N_6951,N_7121);
nand U9825 (N_9825,N_5391,N_7190);
nor U9826 (N_9826,N_7224,N_6449);
and U9827 (N_9827,N_6679,N_5979);
nor U9828 (N_9828,N_7205,N_6920);
or U9829 (N_9829,N_6155,N_6645);
nor U9830 (N_9830,N_6102,N_7006);
nand U9831 (N_9831,N_5617,N_5238);
and U9832 (N_9832,N_7096,N_5778);
nor U9833 (N_9833,N_6488,N_6880);
or U9834 (N_9834,N_6513,N_7183);
and U9835 (N_9835,N_6573,N_6719);
or U9836 (N_9836,N_6806,N_6715);
xor U9837 (N_9837,N_5893,N_5740);
or U9838 (N_9838,N_6788,N_6415);
xor U9839 (N_9839,N_6858,N_5283);
or U9840 (N_9840,N_5130,N_6468);
or U9841 (N_9841,N_7292,N_6640);
nand U9842 (N_9842,N_5434,N_5150);
and U9843 (N_9843,N_6450,N_6044);
nand U9844 (N_9844,N_5628,N_6465);
xnor U9845 (N_9845,N_5137,N_5612);
and U9846 (N_9846,N_5661,N_5645);
xor U9847 (N_9847,N_6583,N_6475);
nand U9848 (N_9848,N_6660,N_5062);
or U9849 (N_9849,N_5793,N_5944);
nand U9850 (N_9850,N_5777,N_5103);
and U9851 (N_9851,N_6917,N_5726);
nor U9852 (N_9852,N_5430,N_6214);
xor U9853 (N_9853,N_5737,N_7018);
nor U9854 (N_9854,N_5740,N_6805);
and U9855 (N_9855,N_6146,N_7233);
nor U9856 (N_9856,N_7252,N_6972);
nor U9857 (N_9857,N_7365,N_5267);
or U9858 (N_9858,N_5457,N_6281);
and U9859 (N_9859,N_6157,N_7112);
nor U9860 (N_9860,N_5566,N_5636);
or U9861 (N_9861,N_7424,N_6791);
xor U9862 (N_9862,N_7126,N_6810);
nand U9863 (N_9863,N_6389,N_7030);
and U9864 (N_9864,N_7434,N_5944);
nor U9865 (N_9865,N_7096,N_6790);
nand U9866 (N_9866,N_6742,N_5491);
or U9867 (N_9867,N_5056,N_5491);
or U9868 (N_9868,N_6417,N_5395);
nand U9869 (N_9869,N_5548,N_5033);
nand U9870 (N_9870,N_7149,N_5589);
nor U9871 (N_9871,N_5158,N_5353);
nand U9872 (N_9872,N_5053,N_7383);
nand U9873 (N_9873,N_5902,N_6260);
xnor U9874 (N_9874,N_6257,N_6335);
xnor U9875 (N_9875,N_5700,N_6854);
nand U9876 (N_9876,N_6106,N_5341);
or U9877 (N_9877,N_5999,N_6935);
xnor U9878 (N_9878,N_6113,N_5709);
nand U9879 (N_9879,N_5454,N_5534);
and U9880 (N_9880,N_5942,N_7150);
xor U9881 (N_9881,N_5686,N_6712);
nand U9882 (N_9882,N_5531,N_6331);
or U9883 (N_9883,N_5239,N_6721);
xor U9884 (N_9884,N_7427,N_5780);
nor U9885 (N_9885,N_5916,N_6854);
xor U9886 (N_9886,N_7307,N_5164);
nor U9887 (N_9887,N_6669,N_6292);
or U9888 (N_9888,N_5792,N_6133);
nor U9889 (N_9889,N_6431,N_6019);
and U9890 (N_9890,N_7114,N_5808);
nor U9891 (N_9891,N_7069,N_6098);
nand U9892 (N_9892,N_7138,N_7184);
xnor U9893 (N_9893,N_6691,N_6066);
and U9894 (N_9894,N_5387,N_5578);
nand U9895 (N_9895,N_6148,N_5231);
or U9896 (N_9896,N_5726,N_7455);
nor U9897 (N_9897,N_6557,N_7368);
xor U9898 (N_9898,N_5843,N_6012);
or U9899 (N_9899,N_6975,N_7235);
nor U9900 (N_9900,N_6896,N_5047);
nand U9901 (N_9901,N_7068,N_6793);
xor U9902 (N_9902,N_5072,N_6718);
and U9903 (N_9903,N_7284,N_5732);
xor U9904 (N_9904,N_5596,N_5732);
xor U9905 (N_9905,N_6051,N_6972);
nor U9906 (N_9906,N_5525,N_5905);
nand U9907 (N_9907,N_5476,N_6207);
nor U9908 (N_9908,N_5295,N_5558);
and U9909 (N_9909,N_5450,N_5493);
nand U9910 (N_9910,N_6764,N_6823);
or U9911 (N_9911,N_7223,N_5913);
and U9912 (N_9912,N_5853,N_5467);
and U9913 (N_9913,N_7163,N_5611);
xnor U9914 (N_9914,N_6253,N_5303);
or U9915 (N_9915,N_5904,N_5711);
nor U9916 (N_9916,N_7183,N_6079);
and U9917 (N_9917,N_5671,N_7324);
nand U9918 (N_9918,N_6355,N_6987);
or U9919 (N_9919,N_6161,N_6926);
nand U9920 (N_9920,N_5833,N_6591);
and U9921 (N_9921,N_5308,N_6490);
nor U9922 (N_9922,N_5452,N_7183);
and U9923 (N_9923,N_5834,N_6595);
xnor U9924 (N_9924,N_6669,N_6778);
or U9925 (N_9925,N_7223,N_5849);
nand U9926 (N_9926,N_5070,N_5430);
nor U9927 (N_9927,N_6868,N_6799);
and U9928 (N_9928,N_6851,N_6626);
xor U9929 (N_9929,N_6701,N_5743);
and U9930 (N_9930,N_6302,N_6493);
nor U9931 (N_9931,N_6857,N_6006);
xnor U9932 (N_9932,N_6750,N_6309);
and U9933 (N_9933,N_6227,N_5487);
nor U9934 (N_9934,N_5445,N_6844);
and U9935 (N_9935,N_7011,N_5769);
and U9936 (N_9936,N_7274,N_6163);
or U9937 (N_9937,N_6999,N_6715);
xor U9938 (N_9938,N_5086,N_7068);
and U9939 (N_9939,N_6886,N_5248);
nor U9940 (N_9940,N_5486,N_7338);
nor U9941 (N_9941,N_6147,N_6286);
or U9942 (N_9942,N_5866,N_5432);
and U9943 (N_9943,N_5614,N_5759);
xnor U9944 (N_9944,N_6379,N_6027);
and U9945 (N_9945,N_6984,N_6402);
and U9946 (N_9946,N_7338,N_6655);
and U9947 (N_9947,N_6889,N_5159);
nor U9948 (N_9948,N_7373,N_5718);
nand U9949 (N_9949,N_5136,N_5874);
xor U9950 (N_9950,N_5856,N_5257);
xor U9951 (N_9951,N_5511,N_7107);
or U9952 (N_9952,N_5281,N_5452);
nor U9953 (N_9953,N_6935,N_6406);
nor U9954 (N_9954,N_7273,N_5783);
nor U9955 (N_9955,N_5111,N_6516);
nand U9956 (N_9956,N_6087,N_6289);
xor U9957 (N_9957,N_5766,N_6709);
or U9958 (N_9958,N_7385,N_6678);
and U9959 (N_9959,N_5959,N_7316);
or U9960 (N_9960,N_6894,N_6012);
or U9961 (N_9961,N_5883,N_6556);
or U9962 (N_9962,N_6082,N_5879);
or U9963 (N_9963,N_5171,N_5614);
nor U9964 (N_9964,N_6538,N_6846);
xor U9965 (N_9965,N_6933,N_6955);
xor U9966 (N_9966,N_6448,N_5297);
xor U9967 (N_9967,N_5547,N_5665);
nand U9968 (N_9968,N_5065,N_5135);
or U9969 (N_9969,N_6935,N_6869);
nand U9970 (N_9970,N_7058,N_5316);
and U9971 (N_9971,N_6870,N_7268);
and U9972 (N_9972,N_6515,N_6043);
nor U9973 (N_9973,N_7266,N_6247);
nand U9974 (N_9974,N_5162,N_5171);
nor U9975 (N_9975,N_5880,N_6470);
nand U9976 (N_9976,N_5997,N_7305);
xnor U9977 (N_9977,N_6399,N_5223);
or U9978 (N_9978,N_6622,N_5612);
or U9979 (N_9979,N_6641,N_5614);
nor U9980 (N_9980,N_6901,N_6096);
xnor U9981 (N_9981,N_5754,N_7426);
or U9982 (N_9982,N_5716,N_5152);
nor U9983 (N_9983,N_5338,N_5183);
and U9984 (N_9984,N_5855,N_6545);
nand U9985 (N_9985,N_6465,N_6241);
or U9986 (N_9986,N_5412,N_5307);
or U9987 (N_9987,N_5966,N_7129);
xnor U9988 (N_9988,N_6259,N_5816);
and U9989 (N_9989,N_5309,N_5762);
and U9990 (N_9990,N_7487,N_6780);
nor U9991 (N_9991,N_5047,N_5417);
xnor U9992 (N_9992,N_6718,N_6867);
xor U9993 (N_9993,N_5523,N_6748);
nand U9994 (N_9994,N_6194,N_5000);
or U9995 (N_9995,N_7445,N_7359);
or U9996 (N_9996,N_7195,N_5594);
nor U9997 (N_9997,N_6418,N_7139);
and U9998 (N_9998,N_6836,N_6390);
nand U9999 (N_9999,N_7403,N_7106);
xnor U10000 (N_10000,N_8938,N_9616);
xor U10001 (N_10001,N_7922,N_8344);
xnor U10002 (N_10002,N_8851,N_8150);
nand U10003 (N_10003,N_9638,N_8961);
or U10004 (N_10004,N_9433,N_9354);
xnor U10005 (N_10005,N_7977,N_8746);
nand U10006 (N_10006,N_9088,N_8117);
and U10007 (N_10007,N_8881,N_7889);
or U10008 (N_10008,N_8037,N_7806);
and U10009 (N_10009,N_9317,N_8358);
xor U10010 (N_10010,N_8660,N_8108);
or U10011 (N_10011,N_9807,N_7856);
nand U10012 (N_10012,N_8917,N_7942);
nand U10013 (N_10013,N_8871,N_8270);
nand U10014 (N_10014,N_9056,N_7907);
xnor U10015 (N_10015,N_8352,N_9707);
nor U10016 (N_10016,N_7507,N_9199);
and U10017 (N_10017,N_7840,N_9685);
nor U10018 (N_10018,N_9168,N_9187);
xor U10019 (N_10019,N_9725,N_8217);
xor U10020 (N_10020,N_8130,N_9206);
xnor U10021 (N_10021,N_7800,N_8215);
nand U10022 (N_10022,N_7620,N_7743);
xor U10023 (N_10023,N_9784,N_8387);
or U10024 (N_10024,N_9870,N_8191);
xor U10025 (N_10025,N_9937,N_9138);
nand U10026 (N_10026,N_7905,N_7625);
nand U10027 (N_10027,N_8714,N_8866);
nor U10028 (N_10028,N_8870,N_8311);
and U10029 (N_10029,N_9182,N_7923);
nand U10030 (N_10030,N_9911,N_8452);
nand U10031 (N_10031,N_8659,N_9126);
nand U10032 (N_10032,N_8098,N_8619);
nand U10033 (N_10033,N_8239,N_7698);
or U10034 (N_10034,N_9779,N_9503);
xor U10035 (N_10035,N_7647,N_9236);
nor U10036 (N_10036,N_7991,N_8367);
nand U10037 (N_10037,N_9452,N_9595);
or U10038 (N_10038,N_8213,N_9411);
nand U10039 (N_10039,N_9566,N_9408);
nand U10040 (N_10040,N_9170,N_9618);
nand U10041 (N_10041,N_9901,N_7906);
or U10042 (N_10042,N_8821,N_9283);
or U10043 (N_10043,N_7848,N_8374);
or U10044 (N_10044,N_9254,N_9607);
xor U10045 (N_10045,N_8815,N_7535);
or U10046 (N_10046,N_9213,N_8685);
xnor U10047 (N_10047,N_8987,N_9373);
nor U10048 (N_10048,N_7694,N_9844);
or U10049 (N_10049,N_8470,N_7682);
nand U10050 (N_10050,N_9415,N_9293);
nor U10051 (N_10051,N_7758,N_8722);
nor U10052 (N_10052,N_8805,N_8534);
xor U10053 (N_10053,N_9852,N_8835);
or U10054 (N_10054,N_8644,N_7735);
and U10055 (N_10055,N_9800,N_7777);
xor U10056 (N_10056,N_8400,N_8365);
nand U10057 (N_10057,N_8043,N_9387);
xnor U10058 (N_10058,N_8364,N_9572);
xor U10059 (N_10059,N_9322,N_9127);
nor U10060 (N_10060,N_9396,N_8186);
and U10061 (N_10061,N_8732,N_7787);
xnor U10062 (N_10062,N_9392,N_8554);
nand U10063 (N_10063,N_9550,N_8220);
or U10064 (N_10064,N_7861,N_8710);
nand U10065 (N_10065,N_7669,N_8002);
nor U10066 (N_10066,N_7707,N_8971);
nand U10067 (N_10067,N_8095,N_8583);
nor U10068 (N_10068,N_9027,N_9704);
and U10069 (N_10069,N_8692,N_8886);
nor U10070 (N_10070,N_8234,N_9274);
and U10071 (N_10071,N_7830,N_7614);
or U10072 (N_10072,N_9519,N_8636);
xnor U10073 (N_10073,N_7641,N_9553);
xor U10074 (N_10074,N_9804,N_8308);
and U10075 (N_10075,N_8051,N_8676);
or U10076 (N_10076,N_9172,N_8891);
and U10077 (N_10077,N_7703,N_9637);
nand U10078 (N_10078,N_8544,N_9710);
nand U10079 (N_10079,N_7779,N_9507);
or U10080 (N_10080,N_7846,N_8582);
nor U10081 (N_10081,N_8836,N_8492);
and U10082 (N_10082,N_8459,N_7926);
nand U10083 (N_10083,N_9668,N_8229);
or U10084 (N_10084,N_7911,N_9690);
and U10085 (N_10085,N_9526,N_9301);
or U10086 (N_10086,N_8696,N_9313);
xnor U10087 (N_10087,N_8376,N_9218);
or U10088 (N_10088,N_8238,N_9399);
nand U10089 (N_10089,N_9070,N_9255);
or U10090 (N_10090,N_9693,N_8713);
nand U10091 (N_10091,N_9863,N_8741);
or U10092 (N_10092,N_7594,N_8740);
or U10093 (N_10093,N_8324,N_7757);
and U10094 (N_10094,N_7900,N_7903);
or U10095 (N_10095,N_8353,N_9688);
xnor U10096 (N_10096,N_8859,N_8794);
nor U10097 (N_10097,N_8342,N_7933);
xor U10098 (N_10098,N_8883,N_8813);
and U10099 (N_10099,N_8826,N_8251);
and U10100 (N_10100,N_7601,N_9555);
xnor U10101 (N_10101,N_9895,N_8960);
xnor U10102 (N_10102,N_8514,N_7695);
nand U10103 (N_10103,N_8924,N_9980);
nor U10104 (N_10104,N_7710,N_7638);
nand U10105 (N_10105,N_7585,N_8911);
and U10106 (N_10106,N_9906,N_8857);
and U10107 (N_10107,N_8996,N_9943);
or U10108 (N_10108,N_8314,N_7843);
xor U10109 (N_10109,N_8372,N_9936);
xnor U10110 (N_10110,N_9064,N_8418);
and U10111 (N_10111,N_9613,N_7578);
and U10112 (N_10112,N_9682,N_9259);
nand U10113 (N_10113,N_7804,N_8417);
or U10114 (N_10114,N_9952,N_9375);
or U10115 (N_10115,N_9588,N_9402);
or U10116 (N_10116,N_7718,N_8793);
xor U10117 (N_10117,N_8007,N_9820);
or U10118 (N_10118,N_8904,N_8948);
xnor U10119 (N_10119,N_7603,N_9278);
nor U10120 (N_10120,N_8884,N_9294);
xor U10121 (N_10121,N_9040,N_9030);
nand U10122 (N_10122,N_8631,N_9081);
nand U10123 (N_10123,N_9038,N_8188);
and U10124 (N_10124,N_9381,N_9847);
and U10125 (N_10125,N_7720,N_7755);
nand U10126 (N_10126,N_8466,N_8716);
nor U10127 (N_10127,N_9031,N_9380);
xnor U10128 (N_10128,N_9496,N_7795);
nor U10129 (N_10129,N_8966,N_8927);
or U10130 (N_10130,N_9851,N_7870);
or U10131 (N_10131,N_9224,N_8548);
and U10132 (N_10132,N_9769,N_9882);
and U10133 (N_10133,N_8993,N_9592);
nand U10134 (N_10134,N_8616,N_9214);
nor U10135 (N_10135,N_8183,N_9403);
or U10136 (N_10136,N_9926,N_8882);
nor U10137 (N_10137,N_8686,N_9540);
and U10138 (N_10138,N_9664,N_8280);
nor U10139 (N_10139,N_7636,N_8428);
and U10140 (N_10140,N_9130,N_8590);
nor U10141 (N_10141,N_9098,N_8675);
or U10142 (N_10142,N_8061,N_9875);
and U10143 (N_10143,N_8091,N_8345);
and U10144 (N_10144,N_8945,N_9709);
and U10145 (N_10145,N_8446,N_9228);
xor U10146 (N_10146,N_7765,N_9086);
nand U10147 (N_10147,N_7910,N_9110);
and U10148 (N_10148,N_9476,N_8808);
nor U10149 (N_10149,N_8063,N_9145);
nand U10150 (N_10150,N_9775,N_9961);
nor U10151 (N_10151,N_7640,N_9249);
and U10152 (N_10152,N_9866,N_8954);
or U10153 (N_10153,N_8187,N_9985);
xnor U10154 (N_10154,N_9343,N_8320);
or U10155 (N_10155,N_8106,N_7521);
or U10156 (N_10156,N_9956,N_8918);
nor U10157 (N_10157,N_8972,N_8723);
nor U10158 (N_10158,N_8463,N_9619);
nor U10159 (N_10159,N_9369,N_7874);
xor U10160 (N_10160,N_8254,N_9517);
xor U10161 (N_10161,N_9651,N_8760);
and U10162 (N_10162,N_9609,N_9571);
nand U10163 (N_10163,N_8067,N_8507);
nand U10164 (N_10164,N_9159,N_7925);
nor U10165 (N_10165,N_7737,N_9243);
or U10166 (N_10166,N_8082,N_9568);
and U10167 (N_10167,N_9312,N_8397);
or U10168 (N_10168,N_7687,N_8440);
nor U10169 (N_10169,N_9597,N_8245);
nor U10170 (N_10170,N_7617,N_7862);
nor U10171 (N_10171,N_9049,N_8946);
xor U10172 (N_10172,N_8936,N_8623);
and U10173 (N_10173,N_9449,N_9564);
nand U10174 (N_10174,N_8385,N_8873);
nor U10175 (N_10175,N_7833,N_7868);
nand U10176 (N_10176,N_8368,N_8286);
and U10177 (N_10177,N_9994,N_8877);
and U10178 (N_10178,N_8756,N_9835);
nand U10179 (N_10179,N_7767,N_9843);
xnor U10180 (N_10180,N_8610,N_8856);
xor U10181 (N_10181,N_8465,N_7835);
and U10182 (N_10182,N_9347,N_7891);
and U10183 (N_10183,N_9802,N_8453);
and U10184 (N_10184,N_9995,N_9378);
xor U10185 (N_10185,N_8216,N_8281);
xor U10186 (N_10186,N_9441,N_9438);
xor U10187 (N_10187,N_8609,N_8173);
or U10188 (N_10188,N_8337,N_9205);
nor U10189 (N_10189,N_7685,N_8162);
xnor U10190 (N_10190,N_8858,N_8155);
and U10191 (N_10191,N_8399,N_7668);
and U10192 (N_10192,N_9511,N_7709);
xor U10193 (N_10193,N_9394,N_9115);
and U10194 (N_10194,N_9101,N_9535);
nor U10195 (N_10195,N_7637,N_8435);
and U10196 (N_10196,N_8131,N_8252);
and U10197 (N_10197,N_8690,N_7932);
xor U10198 (N_10198,N_7766,N_8197);
and U10199 (N_10199,N_9909,N_9385);
xnor U10200 (N_10200,N_9736,N_7985);
and U10201 (N_10201,N_8831,N_7834);
and U10202 (N_10202,N_7505,N_8903);
or U10203 (N_10203,N_8983,N_8908);
and U10204 (N_10204,N_8824,N_7542);
and U10205 (N_10205,N_9979,N_7930);
or U10206 (N_10206,N_8271,N_9796);
nand U10207 (N_10207,N_9220,N_9608);
or U10208 (N_10208,N_9792,N_9950);
nor U10209 (N_10209,N_7885,N_9017);
or U10210 (N_10210,N_9041,N_8982);
and U10211 (N_10211,N_8331,N_8218);
nand U10212 (N_10212,N_8253,N_9084);
or U10213 (N_10213,N_8336,N_9593);
nand U10214 (N_10214,N_8672,N_9495);
nor U10215 (N_10215,N_9014,N_7631);
nand U10216 (N_10216,N_9284,N_8839);
xnor U10217 (N_10217,N_9148,N_9927);
nor U10218 (N_10218,N_8750,N_8485);
xor U10219 (N_10219,N_7956,N_7852);
xnor U10220 (N_10220,N_9247,N_8712);
nor U10221 (N_10221,N_8673,N_9512);
and U10222 (N_10222,N_8158,N_8260);
or U10223 (N_10223,N_8121,N_9591);
or U10224 (N_10224,N_8975,N_8768);
xnor U10225 (N_10225,N_8880,N_9203);
nor U10226 (N_10226,N_8295,N_9417);
nor U10227 (N_10227,N_9741,N_9035);
and U10228 (N_10228,N_9850,N_7722);
nand U10229 (N_10229,N_9718,N_7530);
nor U10230 (N_10230,N_7656,N_9193);
and U10231 (N_10231,N_8231,N_9768);
nor U10232 (N_10232,N_9587,N_9235);
nor U10233 (N_10233,N_8290,N_8436);
nor U10234 (N_10234,N_8152,N_7621);
nand U10235 (N_10235,N_7602,N_9337);
xor U10236 (N_10236,N_9878,N_7534);
or U10237 (N_10237,N_9002,N_8930);
nand U10238 (N_10238,N_8315,N_8471);
or U10239 (N_10239,N_8762,N_7917);
or U10240 (N_10240,N_7527,N_7963);
xnor U10241 (N_10241,N_7524,N_9341);
xor U10242 (N_10242,N_9154,N_9893);
xor U10243 (N_10243,N_7763,N_9240);
or U10244 (N_10244,N_8089,N_8594);
nor U10245 (N_10245,N_8497,N_8167);
nand U10246 (N_10246,N_8994,N_8834);
nand U10247 (N_10247,N_8481,N_8677);
nand U10248 (N_10248,N_9482,N_8810);
nand U10249 (N_10249,N_8057,N_8034);
nand U10250 (N_10250,N_8309,N_7597);
and U10251 (N_10251,N_9504,N_8041);
nand U10252 (N_10252,N_8112,N_7775);
or U10253 (N_10253,N_9429,N_9061);
nor U10254 (N_10254,N_9012,N_9414);
nor U10255 (N_10255,N_8107,N_8506);
nand U10256 (N_10256,N_9432,N_8820);
xor U10257 (N_10257,N_8292,N_9633);
nor U10258 (N_10258,N_8472,N_7897);
and U10259 (N_10259,N_7973,N_8450);
nand U10260 (N_10260,N_8643,N_9241);
or U10261 (N_10261,N_9716,N_9972);
xor U10262 (N_10262,N_8640,N_8444);
xor U10263 (N_10263,N_8247,N_8373);
and U10264 (N_10264,N_8703,N_8235);
nand U10265 (N_10265,N_7512,N_9569);
nor U10266 (N_10266,N_9260,N_9303);
xor U10267 (N_10267,N_9376,N_9462);
and U10268 (N_10268,N_8670,N_7877);
and U10269 (N_10269,N_8144,N_7708);
and U10270 (N_10270,N_7705,N_9627);
or U10271 (N_10271,N_9100,N_8088);
xnor U10272 (N_10272,N_7600,N_8460);
xor U10273 (N_10273,N_9421,N_8600);
xnor U10274 (N_10274,N_8495,N_9246);
nand U10275 (N_10275,N_9773,N_9457);
or U10276 (N_10276,N_8906,N_7970);
and U10277 (N_10277,N_8599,N_9678);
or U10278 (N_10278,N_8734,N_8598);
and U10279 (N_10279,N_9036,N_8141);
and U10280 (N_10280,N_7649,N_9386);
nand U10281 (N_10281,N_7577,N_9756);
or U10282 (N_10282,N_8384,N_9112);
xor U10283 (N_10283,N_8763,N_9836);
xor U10284 (N_10284,N_9219,N_9470);
nor U10285 (N_10285,N_8161,N_8093);
and U10286 (N_10286,N_8556,N_9005);
nand U10287 (N_10287,N_9812,N_8114);
nor U10288 (N_10288,N_8123,N_7946);
xnor U10289 (N_10289,N_8897,N_9671);
nor U10290 (N_10290,N_8745,N_9382);
nand U10291 (N_10291,N_7934,N_8687);
or U10292 (N_10292,N_7522,N_9239);
xnor U10293 (N_10293,N_8928,N_8389);
and U10294 (N_10294,N_9781,N_7635);
xor U10295 (N_10295,N_8626,N_9121);
xnor U10296 (N_10296,N_9719,N_8689);
nand U10297 (N_10297,N_8099,N_7878);
or U10298 (N_10298,N_8981,N_8707);
and U10299 (N_10299,N_7915,N_8738);
xor U10300 (N_10300,N_9102,N_8596);
nand U10301 (N_10301,N_9400,N_9819);
nand U10302 (N_10302,N_8953,N_9493);
xnor U10303 (N_10303,N_8962,N_7898);
nor U10304 (N_10304,N_9302,N_7745);
and U10305 (N_10305,N_8242,N_8584);
or U10306 (N_10306,N_9541,N_7776);
nand U10307 (N_10307,N_9596,N_7756);
nand U10308 (N_10308,N_8893,N_7583);
xor U10309 (N_10309,N_9022,N_7947);
and U10310 (N_10310,N_8761,N_9352);
nand U10311 (N_10311,N_9497,N_8869);
xor U10312 (N_10312,N_9448,N_8748);
nor U10313 (N_10313,N_7873,N_8299);
and U10314 (N_10314,N_9748,N_9024);
nor U10315 (N_10315,N_8553,N_8416);
nand U10316 (N_10316,N_7580,N_9065);
or U10317 (N_10317,N_9184,N_9874);
xor U10318 (N_10318,N_9039,N_9516);
nand U10319 (N_10319,N_9771,N_7789);
nand U10320 (N_10320,N_9643,N_8663);
and U10321 (N_10321,N_7884,N_9894);
nor U10322 (N_10322,N_7510,N_8731);
nand U10323 (N_10323,N_7725,N_9295);
nor U10324 (N_10324,N_7960,N_8978);
xor U10325 (N_10325,N_9848,N_9991);
nand U10326 (N_10326,N_9749,N_9478);
xnor U10327 (N_10327,N_7842,N_9885);
or U10328 (N_10328,N_7676,N_9237);
nand U10329 (N_10329,N_8500,N_7860);
and U10330 (N_10330,N_9296,N_8874);
nor U10331 (N_10331,N_9873,N_9288);
xnor U10332 (N_10332,N_8124,N_9599);
nor U10333 (N_10333,N_8825,N_7784);
or U10334 (N_10334,N_9700,N_8525);
nor U10335 (N_10335,N_9267,N_8661);
or U10336 (N_10336,N_9589,N_9965);
xor U10337 (N_10337,N_8044,N_9131);
xor U10338 (N_10338,N_9188,N_8040);
and U10339 (N_10339,N_9058,N_7634);
nand U10340 (N_10340,N_9854,N_9356);
or U10341 (N_10341,N_8795,N_9363);
or U10342 (N_10342,N_8351,N_8457);
xor U10343 (N_10343,N_7540,N_8375);
xnor U10344 (N_10344,N_9522,N_8070);
nand U10345 (N_10345,N_8058,N_9395);
nor U10346 (N_10346,N_8861,N_9862);
and U10347 (N_10347,N_9125,N_9045);
nand U10348 (N_10348,N_8575,N_8468);
and U10349 (N_10349,N_9348,N_9492);
xnor U10350 (N_10350,N_7882,N_8879);
xnor U10351 (N_10351,N_7672,N_7837);
nor U10352 (N_10352,N_8822,N_9310);
xor U10353 (N_10353,N_8023,N_9562);
nand U10354 (N_10354,N_9028,N_8570);
or U10355 (N_10355,N_7734,N_9534);
nand U10356 (N_10356,N_8862,N_7805);
and U10357 (N_10357,N_9477,N_9645);
and U10358 (N_10358,N_8048,N_8050);
and U10359 (N_10359,N_8885,N_9320);
xor U10360 (N_10360,N_7751,N_9451);
nor U10361 (N_10361,N_8766,N_7890);
nor U10362 (N_10362,N_8175,N_7714);
or U10363 (N_10363,N_9136,N_9113);
and U10364 (N_10364,N_9672,N_9015);
or U10365 (N_10365,N_7772,N_7531);
nand U10366 (N_10366,N_8390,N_8411);
nor U10367 (N_10367,N_8285,N_8289);
nand U10368 (N_10368,N_7626,N_8977);
xor U10369 (N_10369,N_8441,N_7717);
nor U10370 (N_10370,N_9905,N_9270);
and U10371 (N_10371,N_8066,N_7579);
nor U10372 (N_10372,N_7517,N_7954);
and U10373 (N_10373,N_7536,N_7630);
or U10374 (N_10374,N_9471,N_9106);
or U10375 (N_10375,N_9500,N_9439);
xnor U10376 (N_10376,N_8012,N_9244);
xor U10377 (N_10377,N_9649,N_8156);
nand U10378 (N_10378,N_8101,N_9305);
nor U10379 (N_10379,N_8394,N_9368);
nand U10380 (N_10380,N_7727,N_8684);
or U10381 (N_10381,N_8038,N_9839);
or U10382 (N_10382,N_7914,N_8473);
or U10383 (N_10383,N_9958,N_9173);
or U10384 (N_10384,N_9232,N_8282);
or U10385 (N_10385,N_8184,N_9147);
xnor U10386 (N_10386,N_8257,N_8042);
or U10387 (N_10387,N_7814,N_9578);
or U10388 (N_10388,N_9581,N_7742);
and U10389 (N_10389,N_9584,N_9225);
nor U10390 (N_10390,N_7568,N_8611);
nand U10391 (N_10391,N_8147,N_7622);
and U10392 (N_10392,N_8724,N_7659);
nand U10393 (N_10393,N_7901,N_8736);
or U10394 (N_10394,N_8475,N_8651);
xor U10395 (N_10395,N_7681,N_7908);
xor U10396 (N_10396,N_9297,N_8438);
xnor U10397 (N_10397,N_9289,N_9810);
or U10398 (N_10398,N_9811,N_8542);
nor U10399 (N_10399,N_9610,N_8550);
or U10400 (N_10400,N_8637,N_8297);
or U10401 (N_10401,N_8014,N_8146);
xnor U10402 (N_10402,N_9953,N_8404);
nand U10403 (N_10403,N_9050,N_9881);
nor U10404 (N_10404,N_8642,N_7984);
nor U10405 (N_10405,N_7724,N_9212);
and U10406 (N_10406,N_9883,N_9648);
or U10407 (N_10407,N_9475,N_8226);
or U10408 (N_10408,N_8476,N_9941);
xor U10409 (N_10409,N_7895,N_8728);
xor U10410 (N_10410,N_9520,N_8221);
and U10411 (N_10411,N_7969,N_8382);
xnor U10412 (N_10412,N_8803,N_7972);
nand U10413 (N_10413,N_9197,N_8018);
nand U10414 (N_10414,N_8432,N_7616);
nand U10415 (N_10415,N_8633,N_9080);
and U10416 (N_10416,N_9673,N_8852);
xnor U10417 (N_10417,N_9712,N_7693);
xnor U10418 (N_10418,N_8786,N_8778);
or U10419 (N_10419,N_9276,N_8595);
xor U10420 (N_10420,N_9787,N_8787);
nand U10421 (N_10421,N_9407,N_7674);
nor U10422 (N_10422,N_9345,N_8137);
or U10423 (N_10423,N_9242,N_8287);
nor U10424 (N_10424,N_9984,N_9198);
nand U10425 (N_10425,N_8464,N_9715);
and U10426 (N_10426,N_9653,N_8076);
nor U10427 (N_10427,N_9546,N_9349);
and U10428 (N_10428,N_9099,N_9308);
and U10429 (N_10429,N_8629,N_9545);
nor U10430 (N_10430,N_9877,N_8343);
xnor U10431 (N_10431,N_9207,N_7988);
and U10432 (N_10432,N_7753,N_9964);
xnor U10433 (N_10433,N_7989,N_8838);
nor U10434 (N_10434,N_9391,N_8817);
xor U10435 (N_10435,N_9180,N_8843);
and U10436 (N_10436,N_9264,N_8228);
xnor U10437 (N_10437,N_9669,N_9765);
or U10438 (N_10438,N_8895,N_8135);
and U10439 (N_10439,N_9279,N_7831);
nor U10440 (N_10440,N_7995,N_8293);
nand U10441 (N_10441,N_8313,N_8201);
or U10442 (N_10442,N_9754,N_8192);
nand U10443 (N_10443,N_9738,N_9124);
nor U10444 (N_10444,N_9268,N_7528);
nor U10445 (N_10445,N_9215,N_9123);
and U10446 (N_10446,N_8539,N_7516);
and U10447 (N_10447,N_7918,N_8347);
and U10448 (N_10448,N_9861,N_7962);
and U10449 (N_10449,N_8065,N_8721);
xnor U10450 (N_10450,N_9766,N_9614);
nor U10451 (N_10451,N_7666,N_7713);
nor U10452 (N_10452,N_8456,N_7605);
or U10453 (N_10453,N_9939,N_8984);
or U10454 (N_10454,N_9120,N_7539);
nor U10455 (N_10455,N_9751,N_7570);
nor U10456 (N_10456,N_7587,N_9932);
or U10457 (N_10457,N_8937,N_9933);
nor U10458 (N_10458,N_8172,N_7808);
xor U10459 (N_10459,N_8420,N_9063);
nor U10460 (N_10460,N_7606,N_8486);
xnor U10461 (N_10461,N_9079,N_7935);
nor U10462 (N_10462,N_8126,N_8046);
or U10463 (N_10463,N_7957,N_8319);
nand U10464 (N_10464,N_7955,N_9632);
and U10465 (N_10465,N_8361,N_7994);
xor U10466 (N_10466,N_7683,N_9988);
and U10467 (N_10467,N_7980,N_8036);
nor U10468 (N_10468,N_9947,N_7648);
xnor U10469 (N_10469,N_9983,N_9582);
nand U10470 (N_10470,N_8491,N_9158);
xnor U10471 (N_10471,N_7850,N_8649);
nand U10472 (N_10472,N_8537,N_7558);
nand U10473 (N_10473,N_9730,N_9372);
xnor U10474 (N_10474,N_8222,N_8205);
xor U10475 (N_10475,N_8209,N_9001);
and U10476 (N_10476,N_8853,N_8952);
or U10477 (N_10477,N_7823,N_9480);
xnor U10478 (N_10478,N_9763,N_8109);
xor U10479 (N_10479,N_7997,N_9731);
xor U10480 (N_10480,N_8800,N_9579);
nor U10481 (N_10481,N_8900,N_9355);
nor U10482 (N_10482,N_8022,N_8198);
or U10483 (N_10483,N_9074,N_9362);
nand U10484 (N_10484,N_7978,N_7770);
or U10485 (N_10485,N_8033,N_9304);
nor U10486 (N_10486,N_8693,N_8828);
xnor U10487 (N_10487,N_9023,N_8017);
nand U10488 (N_10488,N_9004,N_8846);
nor U10489 (N_10489,N_8097,N_8206);
nand U10490 (N_10490,N_9324,N_7798);
xnor U10491 (N_10491,N_8434,N_8711);
or U10492 (N_10492,N_8415,N_9339);
or U10493 (N_10493,N_7658,N_7520);
and U10494 (N_10494,N_9502,N_9271);
xor U10495 (N_10495,N_9903,N_8225);
xor U10496 (N_10496,N_7919,N_9805);
nand U10497 (N_10497,N_9221,N_9361);
xnor U10498 (N_10498,N_8567,N_9216);
nand U10499 (N_10499,N_9251,N_9666);
xnor U10500 (N_10500,N_8772,N_9698);
or U10501 (N_10501,N_7999,N_7596);
nor U10502 (N_10502,N_7607,N_7826);
or U10503 (N_10503,N_8274,N_9151);
nand U10504 (N_10504,N_9948,N_9944);
or U10505 (N_10505,N_9694,N_9160);
nand U10506 (N_10506,N_9641,N_8968);
or U10507 (N_10507,N_8933,N_8160);
or U10508 (N_10508,N_8530,N_9670);
xnor U10509 (N_10509,N_8455,N_7552);
nand U10510 (N_10510,N_7939,N_8988);
nand U10511 (N_10511,N_8749,N_7712);
nand U10512 (N_10512,N_9547,N_9560);
and U10513 (N_10513,N_9019,N_7686);
nor U10514 (N_10514,N_9824,N_8547);
nand U10515 (N_10515,N_8402,N_9105);
xor U10516 (N_10516,N_9155,N_7886);
or U10517 (N_10517,N_9436,N_9574);
or U10518 (N_10518,N_9186,N_8340);
nor U10519 (N_10519,N_8237,N_7700);
or U10520 (N_10520,N_8096,N_8910);
and U10521 (N_10521,N_9367,N_7642);
nand U10522 (N_10522,N_9307,N_9865);
nor U10523 (N_10523,N_8484,N_9838);
xnor U10524 (N_10524,N_8601,N_9257);
nand U10525 (N_10525,N_7741,N_9636);
and U10526 (N_10526,N_9963,N_9563);
nand U10527 (N_10527,N_8868,N_8812);
nand U10528 (N_10528,N_8605,N_8136);
and U10529 (N_10529,N_8443,N_9938);
nand U10530 (N_10530,N_9652,N_8110);
and U10531 (N_10531,N_9490,N_8671);
and U10532 (N_10532,N_9816,N_9067);
xor U10533 (N_10533,N_9623,N_7711);
xor U10534 (N_10534,N_9795,N_7888);
or U10535 (N_10535,N_7559,N_9726);
and U10536 (N_10536,N_8516,N_7943);
nor U10537 (N_10537,N_7588,N_8422);
nor U10538 (N_10538,N_8275,N_8602);
nor U10539 (N_10539,N_8625,N_9258);
or U10540 (N_10540,N_9798,N_9328);
or U10541 (N_10541,N_8758,N_9879);
nor U10542 (N_10542,N_9423,N_9739);
nor U10543 (N_10543,N_7863,N_8923);
nand U10544 (N_10544,N_9116,N_9007);
nor U10545 (N_10545,N_8512,N_9602);
and U10546 (N_10546,N_9479,N_8262);
nand U10547 (N_10547,N_7748,N_9889);
xor U10548 (N_10548,N_9142,N_9447);
or U10549 (N_10549,N_9097,N_7797);
xor U10550 (N_10550,N_7543,N_8377);
nor U10551 (N_10551,N_9498,N_8383);
or U10552 (N_10552,N_9853,N_7781);
and U10553 (N_10553,N_7665,N_7785);
and U10554 (N_10554,N_9444,N_8538);
nor U10555 (N_10555,N_9857,N_8439);
nand U10556 (N_10556,N_9141,N_7662);
nor U10557 (N_10557,N_9483,N_9639);
nor U10558 (N_10558,N_7819,N_9190);
xnor U10559 (N_10559,N_9860,N_8572);
nor U10560 (N_10560,N_7555,N_9424);
and U10561 (N_10561,N_9764,N_8127);
and U10562 (N_10562,N_8504,N_7750);
xor U10563 (N_10563,N_9277,N_9683);
xnor U10564 (N_10564,N_9508,N_9734);
and U10565 (N_10565,N_8887,N_9531);
nor U10566 (N_10566,N_7818,N_9450);
or U10567 (N_10567,N_8641,N_8739);
or U10568 (N_10568,N_8224,N_9931);
xor U10569 (N_10569,N_8726,N_9412);
nand U10570 (N_10570,N_9679,N_8312);
nand U10571 (N_10571,N_8779,N_7887);
and U10572 (N_10572,N_8326,N_9179);
xnor U10573 (N_10573,N_8769,N_7660);
nor U10574 (N_10574,N_9077,N_8785);
or U10575 (N_10575,N_9405,N_7786);
or U10576 (N_10576,N_8263,N_8341);
nand U10577 (N_10577,N_7582,N_8635);
and U10578 (N_10578,N_7618,N_8378);
and U10579 (N_10579,N_9897,N_8719);
or U10580 (N_10580,N_9156,N_8489);
or U10581 (N_10581,N_9946,N_8301);
and U10582 (N_10582,N_9606,N_8026);
nor U10583 (N_10583,N_9855,N_8490);
xnor U10584 (N_10584,N_9431,N_8102);
nor U10585 (N_10585,N_8913,N_9042);
xnor U10586 (N_10586,N_7774,N_9465);
or U10587 (N_10587,N_8875,N_9311);
nor U10588 (N_10588,N_7913,N_9223);
nor U10589 (N_10589,N_7557,N_9467);
or U10590 (N_10590,N_8190,N_8360);
xor U10591 (N_10591,N_9923,N_8627);
nor U10592 (N_10592,N_7858,N_8129);
nand U10593 (N_10593,N_7747,N_7793);
nor U10594 (N_10594,N_9675,N_8273);
nor U10595 (N_10595,N_8024,N_8030);
nor U10596 (N_10596,N_9822,N_8560);
nand U10597 (N_10597,N_8219,N_8979);
or U10598 (N_10598,N_9955,N_8833);
or U10599 (N_10599,N_8919,N_8009);
xor U10600 (N_10600,N_9515,N_8305);
xor U10601 (N_10601,N_8356,N_8348);
nand U10602 (N_10602,N_7839,N_8612);
nor U10603 (N_10603,N_8566,N_8591);
and U10604 (N_10604,N_8593,N_8277);
nand U10605 (N_10605,N_9434,N_8549);
or U10606 (N_10606,N_8433,N_8170);
nand U10607 (N_10607,N_9506,N_8149);
or U10608 (N_10608,N_9696,N_9181);
or U10609 (N_10609,N_8832,N_9997);
and U10610 (N_10610,N_7810,N_8568);
nand U10611 (N_10611,N_9073,N_9152);
nand U10612 (N_10612,N_8458,N_8501);
and U10613 (N_10613,N_7575,N_8533);
and U10614 (N_10614,N_7813,N_9868);
and U10615 (N_10615,N_9780,N_9728);
and U10616 (N_10616,N_9252,N_9573);
xnor U10617 (N_10617,N_8143,N_7729);
xor U10618 (N_10618,N_8515,N_8699);
or U10619 (N_10619,N_9003,N_8330);
and U10620 (N_10620,N_9891,N_9025);
nor U10621 (N_10621,N_9743,N_8581);
nor U10622 (N_10622,N_7768,N_8743);
or U10623 (N_10623,N_8119,N_9542);
nor U10624 (N_10624,N_8545,N_9913);
nand U10625 (N_10625,N_8752,N_8379);
nor U10626 (N_10626,N_9650,N_7696);
nor U10627 (N_10627,N_9999,N_7701);
or U10628 (N_10628,N_8448,N_7953);
nor U10629 (N_10629,N_8084,N_7692);
or U10630 (N_10630,N_9020,N_7792);
nand U10631 (N_10631,N_7822,N_9622);
or U10632 (N_10632,N_7836,N_9841);
or U10633 (N_10633,N_8957,N_7938);
nor U10634 (N_10634,N_9803,N_7553);
and U10635 (N_10635,N_7723,N_7663);
and U10636 (N_10636,N_9150,N_9194);
and U10637 (N_10637,N_7967,N_7998);
or U10638 (N_10638,N_9548,N_8059);
xnor U10639 (N_10639,N_8789,N_8157);
or U10640 (N_10640,N_8510,N_7556);
or U10641 (N_10641,N_9122,N_9556);
nand U10642 (N_10642,N_8614,N_8480);
nand U10643 (N_10643,N_9009,N_8196);
and U10644 (N_10644,N_9175,N_9018);
nor U10645 (N_10645,N_7993,N_9292);
xor U10646 (N_10646,N_8698,N_8942);
xnor U10647 (N_10647,N_8682,N_7562);
nor U10648 (N_10648,N_9358,N_8970);
or U10649 (N_10649,N_8483,N_7547);
and U10650 (N_10650,N_8288,N_9786);
nand U10651 (N_10651,N_9982,N_8797);
and U10652 (N_10652,N_8276,N_7538);
nand U10653 (N_10653,N_8780,N_8250);
or U10654 (N_10654,N_8317,N_9344);
nor U10655 (N_10655,N_7628,N_7549);
or U10656 (N_10656,N_8060,N_7651);
xor U10657 (N_10657,N_7802,N_7644);
nor U10658 (N_10658,N_9418,N_8969);
and U10659 (N_10659,N_7876,N_8306);
and U10660 (N_10660,N_9072,N_8565);
nor U10661 (N_10661,N_7688,N_9708);
nand U10662 (N_10662,N_7982,N_9149);
xnor U10663 (N_10663,N_9817,N_8303);
xnor U10664 (N_10664,N_8630,N_8876);
nand U10665 (N_10665,N_8248,N_8437);
or U10666 (N_10666,N_9060,N_7719);
nor U10667 (N_10667,N_9724,N_7574);
or U10668 (N_10668,N_8381,N_9699);
and U10669 (N_10669,N_8705,N_9667);
xnor U10670 (N_10670,N_8159,N_7533);
nand U10671 (N_10671,N_8425,N_9428);
and U10672 (N_10672,N_9717,N_9489);
or U10673 (N_10673,N_8648,N_8944);
nand U10674 (N_10674,N_9806,N_8055);
xor U10675 (N_10675,N_8115,N_9353);
xor U10676 (N_10676,N_8487,N_9974);
or U10677 (N_10677,N_8767,N_7761);
or U10678 (N_10678,N_9185,N_8680);
nor U10679 (N_10679,N_8081,N_9351);
nand U10680 (N_10680,N_9513,N_7545);
or U10681 (N_10681,N_8943,N_9549);
nor U10682 (N_10682,N_7788,N_7646);
xnor U10683 (N_10683,N_8922,N_7744);
or U10684 (N_10684,N_7853,N_7563);
nand U10685 (N_10685,N_9420,N_9887);
or U10686 (N_10686,N_8811,N_7892);
nand U10687 (N_10687,N_7859,N_8462);
or U10688 (N_10688,N_8298,N_9799);
nand U10689 (N_10689,N_9740,N_8087);
or U10690 (N_10690,N_7847,N_8335);
nor U10691 (N_10691,N_8008,N_9907);
and U10692 (N_10692,N_9275,N_8860);
nor U10693 (N_10693,N_8809,N_8540);
xnor U10694 (N_10694,N_9880,N_7619);
xnor U10695 (N_10695,N_8956,N_8355);
and U10696 (N_10696,N_9642,N_9998);
nor U10697 (N_10697,N_8939,N_8607);
nor U10698 (N_10698,N_9539,N_9189);
nor U10699 (N_10699,N_9318,N_7503);
nand U10700 (N_10700,N_9654,N_9455);
nand U10701 (N_10701,N_9954,N_9069);
nor U10702 (N_10702,N_7902,N_7824);
nand U10703 (N_10703,N_7624,N_9401);
xor U10704 (N_10704,N_8424,N_9309);
or U10705 (N_10705,N_8733,N_8255);
nor U10706 (N_10706,N_9196,N_8423);
and U10707 (N_10707,N_9750,N_8751);
xor U10708 (N_10708,N_7975,N_9332);
and U10709 (N_10709,N_8620,N_9969);
xor U10710 (N_10710,N_9487,N_9248);
xor U10711 (N_10711,N_9744,N_8163);
xnor U10712 (N_10712,N_8523,N_9200);
xor U10713 (N_10713,N_9404,N_9229);
xor U10714 (N_10714,N_9524,N_9285);
xnor U10715 (N_10715,N_8264,N_9048);
nand U10716 (N_10716,N_8431,N_9419);
xnor U10717 (N_10717,N_9869,N_8045);
or U10718 (N_10718,N_8980,N_7740);
and U10719 (N_10719,N_9829,N_7829);
or U10720 (N_10720,N_7523,N_7820);
nand U10721 (N_10721,N_9262,N_9008);
nand U10722 (N_10722,N_7731,N_7880);
xor U10723 (N_10723,N_9864,N_7506);
or U10724 (N_10724,N_8442,N_9426);
or U10725 (N_10725,N_8935,N_8177);
or U10726 (N_10726,N_9192,N_7508);
or U10727 (N_10727,N_7699,N_8715);
nor U10728 (N_10728,N_7732,N_9090);
and U10729 (N_10729,N_9327,N_7645);
xor U10730 (N_10730,N_8369,N_9975);
or U10731 (N_10731,N_8010,N_7794);
nand U10732 (N_10732,N_9697,N_7571);
or U10733 (N_10733,N_8896,N_7857);
and U10734 (N_10734,N_8182,N_9888);
nor U10735 (N_10735,N_8818,N_8709);
nand U10736 (N_10736,N_8211,N_9989);
and U10737 (N_10737,N_8559,N_8079);
or U10738 (N_10738,N_8246,N_9902);
nor U10739 (N_10739,N_7551,N_9144);
and U10740 (N_10740,N_9117,N_7780);
or U10741 (N_10741,N_9253,N_8717);
xor U10742 (N_10742,N_8603,N_9559);
nor U10743 (N_10743,N_9701,N_9057);
and U10744 (N_10744,N_8080,N_9986);
xnor U10745 (N_10745,N_7611,N_8474);
or U10746 (N_10746,N_7615,N_9778);
nor U10747 (N_10747,N_9640,N_8915);
or U10748 (N_10748,N_9557,N_8655);
nor U10749 (N_10749,N_9443,N_7951);
nand U10750 (N_10750,N_9458,N_9942);
or U10751 (N_10751,N_8000,N_8429);
nor U10752 (N_10752,N_8639,N_7736);
xor U10753 (N_10753,N_9665,N_8174);
and U10754 (N_10754,N_8855,N_8086);
xnor U10755 (N_10755,N_8771,N_9842);
nor U10756 (N_10756,N_8799,N_8658);
and U10757 (N_10757,N_7796,N_7610);
or U10758 (N_10758,N_8477,N_8517);
nor U10759 (N_10759,N_9440,N_9107);
or U10760 (N_10760,N_9809,N_9876);
nand U10761 (N_10761,N_9335,N_8258);
xor U10762 (N_10762,N_9217,N_7609);
nor U10763 (N_10763,N_7762,N_9977);
nor U10764 (N_10764,N_8116,N_9917);
and U10765 (N_10765,N_8393,N_9825);
nand U10766 (N_10766,N_7537,N_7799);
nand U10767 (N_10767,N_8419,N_9821);
nor U10768 (N_10768,N_9808,N_7949);
nand U10769 (N_10769,N_8359,N_8656);
and U10770 (N_10770,N_7971,N_9379);
nand U10771 (N_10771,N_8574,N_9286);
and U10772 (N_10772,N_9171,N_8624);
nand U10773 (N_10773,N_9397,N_9630);
and U10774 (N_10774,N_8232,N_8194);
nand U10775 (N_10775,N_9266,N_7961);
nor U10776 (N_10776,N_7670,N_9245);
or U10777 (N_10777,N_8138,N_9227);
nand U10778 (N_10778,N_8256,N_7673);
nand U10779 (N_10779,N_7738,N_8140);
nand U10780 (N_10780,N_9054,N_7684);
nor U10781 (N_10781,N_9957,N_7667);
and U10782 (N_10782,N_7629,N_9552);
nor U10783 (N_10783,N_9454,N_9059);
nand U10784 (N_10784,N_7894,N_8310);
nand U10785 (N_10785,N_9598,N_9919);
nor U10786 (N_10786,N_8518,N_9066);
nor U10787 (N_10787,N_9706,N_8111);
and U10788 (N_10788,N_8072,N_8467);
and U10789 (N_10789,N_8204,N_8973);
nor U10790 (N_10790,N_9233,N_7548);
nor U10791 (N_10791,N_8113,N_7976);
nand U10792 (N_10792,N_7945,N_8139);
or U10793 (N_10793,N_9898,N_8078);
nand U10794 (N_10794,N_9762,N_9949);
nor U10795 (N_10795,N_9167,N_9453);
xor U10796 (N_10796,N_9910,N_9968);
nor U10797 (N_10797,N_9576,N_8410);
nor U10798 (N_10798,N_9747,N_8505);
nor U10799 (N_10799,N_8951,N_9132);
nor U10800 (N_10800,N_8318,N_9357);
or U10801 (N_10801,N_7657,N_7879);
nand U10802 (N_10802,N_9723,N_9727);
nand U10803 (N_10803,N_7613,N_8576);
xnor U10804 (N_10804,N_8850,N_8181);
and U10805 (N_10805,N_9053,N_7746);
or U10806 (N_10806,N_8564,N_9319);
nand U10807 (N_10807,N_8180,N_9435);
nor U10808 (N_10808,N_9713,N_9692);
nand U10809 (N_10809,N_7643,N_8774);
xor U10810 (N_10810,N_9210,N_9103);
and U10811 (N_10811,N_7927,N_9460);
xor U10812 (N_10812,N_9827,N_8451);
nor U10813 (N_10813,N_9990,N_9300);
or U10814 (N_10814,N_9316,N_9374);
or U10815 (N_10815,N_9006,N_8819);
nor U10816 (N_10816,N_8199,N_8865);
or U10817 (N_10817,N_8907,N_9076);
nor U10818 (N_10818,N_8552,N_8508);
and U10819 (N_10819,N_9051,N_7529);
xnor U10820 (N_10820,N_8765,N_9393);
or U10821 (N_10821,N_7948,N_9306);
xor U10822 (N_10822,N_7502,N_8445);
nor U10823 (N_10823,N_7875,N_8796);
nand U10824 (N_10824,N_9899,N_9128);
and U10825 (N_10825,N_9095,N_8902);
xor U10826 (N_10826,N_7992,N_9191);
nor U10827 (N_10827,N_8588,N_9409);
nand U10828 (N_10828,N_7650,N_8029);
nor U10829 (N_10829,N_8864,N_8398);
nor U10830 (N_10830,N_7896,N_9745);
nor U10831 (N_10831,N_8279,N_8498);
nand U10832 (N_10832,N_8321,N_9010);
nand U10833 (N_10833,N_9759,N_8999);
nor U10834 (N_10834,N_7584,N_9859);
and U10835 (N_10835,N_9644,N_8208);
or U10836 (N_10836,N_8125,N_8019);
and U10837 (N_10837,N_8662,N_7983);
or U10838 (N_10838,N_8001,N_8562);
and U10839 (N_10839,N_7827,N_8718);
or U10840 (N_10840,N_8346,N_9735);
and U10841 (N_10841,N_8151,N_9331);
and U10842 (N_10842,N_8744,N_9705);
xnor U10843 (N_10843,N_8837,N_8959);
xor U10844 (N_10844,N_9600,N_8804);
or U10845 (N_10845,N_8997,N_9840);
nor U10846 (N_10846,N_7608,N_7845);
xor U10847 (N_10847,N_8628,N_9340);
nand U10848 (N_10848,N_7560,N_8334);
and U10849 (N_10849,N_8240,N_9663);
nand U10850 (N_10850,N_9761,N_9612);
and U10851 (N_10851,N_9000,N_8214);
and U10852 (N_10852,N_9326,N_9265);
nand U10853 (N_10853,N_8267,N_8062);
and U10854 (N_10854,N_8412,N_9996);
nor U10855 (N_10855,N_8664,N_7803);
or U10856 (N_10856,N_9791,N_8541);
nor U10857 (N_10857,N_7893,N_9966);
or U10858 (N_10858,N_9427,N_8006);
or U10859 (N_10859,N_8947,N_7721);
nor U10860 (N_10860,N_9442,N_8697);
nand U10861 (N_10861,N_9580,N_8386);
xnor U10862 (N_10862,N_9767,N_8929);
nor U10863 (N_10863,N_7855,N_8571);
xnor U10864 (N_10864,N_7764,N_9753);
nor U10865 (N_10865,N_8669,N_8985);
nor U10866 (N_10866,N_8754,N_9398);
and U10867 (N_10867,N_8168,N_8210);
nand U10868 (N_10868,N_8569,N_8587);
xor U10869 (N_10869,N_9945,N_9062);
xnor U10870 (N_10870,N_8531,N_8323);
xor U10871 (N_10871,N_8154,N_9746);
and U10872 (N_10872,N_8878,N_9577);
nand U10873 (N_10873,N_9583,N_9788);
and U10874 (N_10874,N_9684,N_8653);
nand U10875 (N_10875,N_9760,N_8546);
nand U10876 (N_10876,N_7654,N_9129);
nand U10877 (N_10877,N_9537,N_9164);
nor U10878 (N_10878,N_9801,N_8027);
xor U10879 (N_10879,N_8284,N_8666);
and U10880 (N_10880,N_9410,N_7509);
nand U10881 (N_10881,N_8934,N_7912);
or U10882 (N_10882,N_9603,N_9789);
nand U10883 (N_10883,N_8647,N_9920);
xnor U10884 (N_10884,N_9729,N_8737);
and U10885 (N_10885,N_8499,N_8589);
xor U10886 (N_10886,N_8841,N_9973);
nor U10887 (N_10887,N_8300,N_8528);
and U10888 (N_10888,N_8781,N_7730);
xor U10889 (N_10889,N_7773,N_8261);
xnor U10890 (N_10890,N_7664,N_9273);
and U10891 (N_10891,N_9445,N_8195);
and U10892 (N_10892,N_9094,N_7778);
nor U10893 (N_10893,N_8729,N_9463);
xnor U10894 (N_10894,N_9703,N_8133);
and U10895 (N_10895,N_9951,N_8557);
and U10896 (N_10896,N_7899,N_9166);
and U10897 (N_10897,N_7541,N_8322);
or U10898 (N_10898,N_8145,N_9091);
or U10899 (N_10899,N_7974,N_9621);
nand U10900 (N_10900,N_8854,N_8621);
nor U10901 (N_10901,N_9833,N_9929);
and U10902 (N_10902,N_8816,N_9231);
nor U10903 (N_10903,N_8304,N_7760);
nor U10904 (N_10904,N_8678,N_9456);
or U10905 (N_10905,N_8788,N_8783);
or U10906 (N_10906,N_9752,N_8203);
nor U10907 (N_10907,N_8925,N_9960);
and U10908 (N_10908,N_8950,N_9677);
nand U10909 (N_10909,N_8802,N_9532);
nand U10910 (N_10910,N_8622,N_8995);
nor U10911 (N_10911,N_8695,N_8998);
and U10912 (N_10912,N_7791,N_9163);
nor U10913 (N_10913,N_9201,N_7864);
or U10914 (N_10914,N_7801,N_8294);
nor U10915 (N_10915,N_8122,N_8223);
or U10916 (N_10916,N_7950,N_8403);
xnor U10917 (N_10917,N_8683,N_7511);
nor U10918 (N_10918,N_8679,N_7844);
nand U10919 (N_10919,N_7981,N_9987);
xnor U10920 (N_10920,N_9605,N_8667);
nor U10921 (N_10921,N_8069,N_9388);
nand U10922 (N_10922,N_8867,N_8077);
and U10923 (N_10923,N_8176,N_7576);
nand U10924 (N_10924,N_8401,N_9830);
nand U10925 (N_10925,N_8563,N_9282);
or U10926 (N_10926,N_7952,N_8202);
nor U10927 (N_10927,N_9867,N_9346);
and U10928 (N_10928,N_8327,N_9656);
or U10929 (N_10929,N_9390,N_9543);
nor U10930 (N_10930,N_9104,N_8488);
nand U10931 (N_10931,N_7817,N_8094);
nor U10932 (N_10932,N_8847,N_9230);
xor U10933 (N_10933,N_8329,N_8668);
nand U10934 (N_10934,N_8503,N_9620);
nor U10935 (N_10935,N_7593,N_9342);
and U10936 (N_10936,N_8701,N_8075);
or U10937 (N_10937,N_9370,N_8171);
or U10938 (N_10938,N_8396,N_9377);
or U10939 (N_10939,N_9256,N_7715);
and U10940 (N_10940,N_7759,N_8513);
or U10941 (N_10941,N_9208,N_9384);
nor U10942 (N_10942,N_9733,N_7728);
nor U10943 (N_10943,N_7500,N_7940);
and U10944 (N_10944,N_8296,N_9509);
and U10945 (N_10945,N_8958,N_8406);
xor U10946 (N_10946,N_9935,N_8259);
and U10947 (N_10947,N_9567,N_9797);
or U10948 (N_10948,N_8153,N_8461);
nand U10949 (N_10949,N_9604,N_9481);
and U10950 (N_10950,N_9702,N_8888);
or U10951 (N_10951,N_7680,N_9940);
or U10952 (N_10952,N_8617,N_9055);
xnor U10953 (N_10953,N_9089,N_9016);
nand U10954 (N_10954,N_7832,N_8519);
nor U10955 (N_10955,N_7807,N_7851);
and U10956 (N_10956,N_8268,N_8244);
or U10957 (N_10957,N_9554,N_8148);
xor U10958 (N_10958,N_9992,N_9558);
xor U10959 (N_10959,N_8920,N_7661);
nand U10960 (N_10960,N_8328,N_8700);
or U10961 (N_10961,N_8608,N_9772);
and U10962 (N_10962,N_9137,N_8028);
and U10963 (N_10963,N_8005,N_8645);
nand U10964 (N_10964,N_7564,N_8179);
or U10965 (N_10965,N_8083,N_7572);
xnor U10966 (N_10966,N_8964,N_9518);
nor U10967 (N_10967,N_8543,N_9291);
nor U10968 (N_10968,N_7590,N_8790);
and U10969 (N_10969,N_9134,N_9092);
xnor U10970 (N_10970,N_9365,N_8278);
nand U10971 (N_10971,N_9635,N_8720);
and U10972 (N_10972,N_8727,N_8708);
and U10973 (N_10973,N_9790,N_7921);
and U10974 (N_10974,N_8178,N_7733);
nand U10975 (N_10975,N_9770,N_7904);
nor U10976 (N_10976,N_7920,N_9366);
nor U10977 (N_10977,N_9626,N_7841);
or U10978 (N_10978,N_8827,N_9528);
xor U10979 (N_10979,N_9068,N_9631);
xor U10980 (N_10980,N_8967,N_8974);
xor U10981 (N_10981,N_7532,N_8391);
xnor U10982 (N_10982,N_9586,N_7592);
nor U10983 (N_10983,N_8773,N_7702);
xnor U10984 (N_10984,N_8349,N_9174);
nor U10985 (N_10985,N_8899,N_8777);
or U10986 (N_10986,N_8169,N_9299);
xor U10987 (N_10987,N_7671,N_9527);
xor U10988 (N_10988,N_9135,N_8302);
xnor U10989 (N_10989,N_9083,N_7544);
nand U10990 (N_10990,N_9011,N_9111);
or U10991 (N_10991,N_7958,N_9314);
xnor U10992 (N_10992,N_9930,N_8333);
and U10993 (N_10993,N_7573,N_7909);
nor U10994 (N_10994,N_8770,N_9321);
xnor U10995 (N_10995,N_9662,N_9858);
nand U10996 (N_10996,N_9269,N_8283);
nor U10997 (N_10997,N_9287,N_8706);
and U10998 (N_10998,N_9658,N_8020);
nor U10999 (N_10999,N_7979,N_8527);
xor U11000 (N_11000,N_7986,N_9657);
or U11001 (N_11001,N_9601,N_9783);
nor U11002 (N_11002,N_9281,N_8522);
or U11003 (N_11003,N_7501,N_8047);
nand U11004 (N_11004,N_8449,N_7677);
nand U11005 (N_11005,N_8889,N_8909);
and U11006 (N_11006,N_8561,N_9695);
and U11007 (N_11007,N_7726,N_9334);
or U11008 (N_11008,N_7871,N_7883);
and U11009 (N_11009,N_9133,N_9918);
or U11010 (N_11010,N_8388,N_9681);
nand U11011 (N_11011,N_7867,N_9834);
nand U11012 (N_11012,N_8965,N_8370);
xor U11013 (N_11013,N_8207,N_8035);
xnor U11014 (N_11014,N_7518,N_9529);
or U11015 (N_11015,N_8558,N_8634);
or U11016 (N_11016,N_8784,N_8426);
nand U11017 (N_11017,N_7546,N_7632);
and U11018 (N_11018,N_8586,N_9336);
nand U11019 (N_11019,N_8430,N_9561);
and U11020 (N_11020,N_8269,N_8227);
nor U11021 (N_11021,N_8577,N_9469);
nand U11022 (N_11022,N_9691,N_9459);
and U11023 (N_11023,N_9521,N_9333);
and U11024 (N_11024,N_8872,N_7514);
nor U11025 (N_11025,N_9721,N_9794);
xnor U11026 (N_11026,N_9828,N_8316);
and U11027 (N_11027,N_8118,N_8053);
xnor U11028 (N_11028,N_8120,N_7679);
or U11029 (N_11029,N_8013,N_8652);
xnor U11030 (N_11030,N_9013,N_8704);
nand U11031 (N_11031,N_8103,N_8395);
or U11032 (N_11032,N_8363,N_8791);
nand U11033 (N_11033,N_8249,N_9924);
and U11034 (N_11034,N_9928,N_9976);
and U11035 (N_11035,N_7783,N_9437);
nor U11036 (N_11036,N_8747,N_9485);
or U11037 (N_11037,N_9211,N_8016);
nor U11038 (N_11038,N_8730,N_9085);
xor U11039 (N_11039,N_8332,N_9338);
nand U11040 (N_11040,N_9845,N_9466);
nor U11041 (N_11041,N_8236,N_8949);
nor U11042 (N_11042,N_9046,N_8357);
xnor U11043 (N_11043,N_8478,N_7866);
nor U11044 (N_11044,N_8842,N_8742);
or U11045 (N_11045,N_9676,N_7990);
xnor U11046 (N_11046,N_8092,N_8646);
and U11047 (N_11047,N_9021,N_8578);
xnor U11048 (N_11048,N_9590,N_8976);
or U11049 (N_11049,N_8074,N_8806);
and U11050 (N_11050,N_8407,N_9494);
nand U11051 (N_11051,N_8916,N_9714);
nor U11052 (N_11052,N_9818,N_9912);
nor U11053 (N_11053,N_8392,N_9849);
xnor U11054 (N_11054,N_9565,N_9034);
xor U11055 (N_11055,N_8990,N_8521);
and U11056 (N_11056,N_7838,N_9585);
or U11057 (N_11057,N_7706,N_9501);
and U11058 (N_11058,N_8164,N_8801);
and U11059 (N_11059,N_9525,N_7809);
or U11060 (N_11060,N_9646,N_9360);
and U11061 (N_11061,N_7849,N_8691);
nand U11062 (N_11062,N_8764,N_8380);
xnor U11063 (N_11063,N_9364,N_8955);
nand U11064 (N_11064,N_9037,N_9934);
nor U11065 (N_11065,N_9472,N_9491);
and U11066 (N_11066,N_9461,N_9962);
nand U11067 (N_11067,N_9140,N_9915);
nand U11068 (N_11068,N_8454,N_8128);
and U11069 (N_11069,N_7586,N_8052);
nand U11070 (N_11070,N_9872,N_9538);
and U11071 (N_11071,N_7513,N_9114);
nor U11072 (N_11072,N_9793,N_8890);
nand U11073 (N_11073,N_9777,N_7515);
or U11074 (N_11074,N_8681,N_8921);
nor U11075 (N_11075,N_7525,N_9474);
and U11076 (N_11076,N_8665,N_7581);
or U11077 (N_11077,N_7595,N_9143);
nor U11078 (N_11078,N_7964,N_9659);
and U11079 (N_11079,N_8071,N_9425);
or U11080 (N_11080,N_8233,N_7739);
and U11081 (N_11081,N_8551,N_8914);
nand U11082 (N_11082,N_8654,N_9359);
nand U11083 (N_11083,N_9925,N_8339);
and U11084 (N_11084,N_9488,N_7881);
nor U11085 (N_11085,N_9959,N_8782);
nor U11086 (N_11086,N_9446,N_8073);
and U11087 (N_11087,N_9096,N_9389);
and U11088 (N_11088,N_7929,N_9536);
and U11089 (N_11089,N_9505,N_9890);
nor U11090 (N_11090,N_8986,N_8165);
xor U11091 (N_11091,N_9026,N_9575);
or U11092 (N_11092,N_8604,N_9776);
and U11093 (N_11093,N_7865,N_8753);
or U11094 (N_11094,N_9075,N_7690);
and U11095 (N_11095,N_7565,N_7996);
or U11096 (N_11096,N_8408,N_9468);
nand U11097 (N_11097,N_8011,N_8004);
and U11098 (N_11098,N_9422,N_9161);
and U11099 (N_11099,N_8863,N_9178);
and U11100 (N_11100,N_8792,N_9033);
nor U11101 (N_11101,N_9499,N_9530);
or U11102 (N_11102,N_8526,N_8735);
xor U11103 (N_11103,N_8798,N_9165);
nand U11104 (N_11104,N_9209,N_9263);
or U11105 (N_11105,N_7754,N_9087);
nand U11106 (N_11106,N_7959,N_8963);
nor U11107 (N_11107,N_7675,N_7598);
xnor U11108 (N_11108,N_9758,N_8941);
nand U11109 (N_11109,N_9720,N_7916);
xnor U11110 (N_11110,N_9687,N_8585);
xor U11111 (N_11111,N_7924,N_9109);
and U11112 (N_11112,N_9350,N_8898);
xnor U11113 (N_11113,N_9813,N_9484);
xnor U11114 (N_11114,N_8496,N_8266);
xnor U11115 (N_11115,N_9234,N_8511);
or U11116 (N_11116,N_7811,N_9226);
xnor U11117 (N_11117,N_8350,N_7655);
and U11118 (N_11118,N_8845,N_7854);
nand U11119 (N_11119,N_7941,N_8265);
nand U11120 (N_11120,N_9514,N_7937);
and U11121 (N_11121,N_7604,N_8090);
nor U11122 (N_11122,N_8524,N_9900);
nand U11123 (N_11123,N_9272,N_9413);
xor U11124 (N_11124,N_8849,N_9922);
or U11125 (N_11125,N_9044,N_7716);
and U11126 (N_11126,N_9153,N_8366);
and U11127 (N_11127,N_8166,N_8049);
nor U11128 (N_11128,N_9371,N_8291);
nor U11129 (N_11129,N_8650,N_8932);
xor U11130 (N_11130,N_8775,N_8325);
or U11131 (N_11131,N_9078,N_9416);
or U11132 (N_11132,N_9523,N_8992);
or U11133 (N_11133,N_8021,N_9162);
nand U11134 (N_11134,N_9406,N_9108);
or U11135 (N_11135,N_7567,N_8991);
nor U11136 (N_11136,N_9686,N_9628);
or U11137 (N_11137,N_7633,N_7561);
and U11138 (N_11138,N_9473,N_9886);
nor U11139 (N_11139,N_8405,N_9832);
and U11140 (N_11140,N_9856,N_9329);
and U11141 (N_11141,N_7815,N_7944);
xor U11142 (N_11142,N_8015,N_9647);
or U11143 (N_11143,N_9815,N_9967);
nand U11144 (N_11144,N_7623,N_8580);
xnor U11145 (N_11145,N_8613,N_9204);
nand U11146 (N_11146,N_9826,N_9551);
nand U11147 (N_11147,N_9325,N_7653);
xnor U11148 (N_11148,N_9202,N_8032);
nand U11149 (N_11149,N_9814,N_8354);
nand U11150 (N_11150,N_9831,N_8529);
or U11151 (N_11151,N_9774,N_9298);
or U11152 (N_11152,N_9634,N_7591);
and U11153 (N_11153,N_9782,N_9846);
nor U11154 (N_11154,N_7569,N_8494);
nand U11155 (N_11155,N_9981,N_7968);
nand U11156 (N_11156,N_9510,N_7966);
nand U11157 (N_11157,N_8892,N_8414);
nor U11158 (N_11158,N_7691,N_9290);
or U11159 (N_11159,N_8054,N_7639);
and U11160 (N_11160,N_9169,N_9892);
or U11161 (N_11161,N_9655,N_7697);
and U11162 (N_11162,N_7782,N_8193);
nor U11163 (N_11163,N_7554,N_7550);
nand U11164 (N_11164,N_9238,N_9464);
xnor U11165 (N_11165,N_7749,N_9978);
or U11166 (N_11166,N_8132,N_8912);
nor U11167 (N_11167,N_8807,N_8413);
and U11168 (N_11168,N_8479,N_9871);
xnor U11169 (N_11169,N_9970,N_8814);
nand U11170 (N_11170,N_8776,N_8243);
or U11171 (N_11171,N_9904,N_9914);
nor U11172 (N_11172,N_8421,N_9533);
or U11173 (N_11173,N_8757,N_7965);
and U11174 (N_11174,N_9222,N_9052);
nor U11175 (N_11175,N_9029,N_9157);
nand U11176 (N_11176,N_8573,N_8694);
nor U11177 (N_11177,N_8535,N_9742);
nor U11178 (N_11178,N_8536,N_8447);
or U11179 (N_11179,N_9624,N_8100);
xnor U11180 (N_11180,N_9486,N_7931);
and U11181 (N_11181,N_7704,N_9993);
or U11182 (N_11182,N_9323,N_7821);
or U11183 (N_11183,N_8940,N_9195);
xnor U11184 (N_11184,N_7566,N_8469);
nor U11185 (N_11185,N_7589,N_8830);
or U11186 (N_11186,N_9047,N_9660);
and U11187 (N_11187,N_7652,N_8844);
xnor U11188 (N_11188,N_8200,N_8056);
nand U11189 (N_11189,N_8185,N_8493);
nand U11190 (N_11190,N_8615,N_8502);
nand U11191 (N_11191,N_8003,N_7504);
nor U11192 (N_11192,N_8618,N_7769);
or U11193 (N_11193,N_9757,N_9430);
nor U11194 (N_11194,N_8338,N_9737);
xnor U11195 (N_11195,N_9711,N_8409);
xor U11196 (N_11196,N_7816,N_8555);
and U11197 (N_11197,N_9896,N_9661);
nand U11198 (N_11198,N_7526,N_8894);
xnor U11199 (N_11199,N_9544,N_8427);
nor U11200 (N_11200,N_9617,N_8674);
and U11201 (N_11201,N_8212,N_9383);
nand U11202 (N_11202,N_9177,N_9176);
nand U11203 (N_11203,N_8848,N_8068);
or U11204 (N_11204,N_8371,N_7872);
xor U11205 (N_11205,N_9884,N_8230);
nand U11206 (N_11206,N_7987,N_9680);
xnor U11207 (N_11207,N_7627,N_8272);
and U11208 (N_11208,N_7825,N_9315);
nor U11209 (N_11209,N_8104,N_9082);
or U11210 (N_11210,N_9330,N_9732);
xnor U11211 (N_11211,N_9250,N_8823);
or U11212 (N_11212,N_9280,N_8362);
and U11213 (N_11213,N_8702,N_8520);
xor U11214 (N_11214,N_8905,N_8755);
nor U11215 (N_11215,N_9071,N_8597);
and U11216 (N_11216,N_8901,N_7936);
xnor U11217 (N_11217,N_8931,N_9093);
xnor U11218 (N_11218,N_8759,N_8638);
nand U11219 (N_11219,N_9594,N_7599);
xnor U11220 (N_11220,N_8632,N_8241);
xnor U11221 (N_11221,N_9625,N_8031);
xnor U11222 (N_11222,N_8307,N_7812);
and U11223 (N_11223,N_9921,N_9971);
nand U11224 (N_11224,N_9118,N_8989);
xor U11225 (N_11225,N_9146,N_9261);
nor U11226 (N_11226,N_9139,N_9823);
or U11227 (N_11227,N_8579,N_9043);
xor U11228 (N_11228,N_7928,N_9611);
nand U11229 (N_11229,N_9722,N_9916);
xor U11230 (N_11230,N_7771,N_7752);
and U11231 (N_11231,N_7519,N_9689);
or U11232 (N_11232,N_8657,N_9119);
nor U11233 (N_11233,N_9570,N_8509);
or U11234 (N_11234,N_9908,N_9785);
xor U11235 (N_11235,N_9032,N_9629);
or U11236 (N_11236,N_8840,N_7689);
nand U11237 (N_11237,N_9615,N_8064);
or U11238 (N_11238,N_9755,N_8085);
or U11239 (N_11239,N_8688,N_8482);
and U11240 (N_11240,N_8829,N_8025);
or U11241 (N_11241,N_7790,N_8725);
and U11242 (N_11242,N_9837,N_8189);
xnor U11243 (N_11243,N_8606,N_7828);
nand U11244 (N_11244,N_8926,N_8039);
xnor U11245 (N_11245,N_8142,N_7678);
nor U11246 (N_11246,N_8105,N_7612);
nor U11247 (N_11247,N_8592,N_8134);
nand U11248 (N_11248,N_7869,N_9183);
and U11249 (N_11249,N_9674,N_8532);
and U11250 (N_11250,N_9413,N_8303);
nor U11251 (N_11251,N_9634,N_9323);
nor U11252 (N_11252,N_9560,N_7690);
nand U11253 (N_11253,N_8688,N_9816);
nand U11254 (N_11254,N_7853,N_8033);
or U11255 (N_11255,N_9694,N_9310);
and U11256 (N_11256,N_7757,N_8559);
nand U11257 (N_11257,N_9640,N_7912);
nand U11258 (N_11258,N_9080,N_8953);
or U11259 (N_11259,N_8309,N_8122);
xor U11260 (N_11260,N_8144,N_8687);
nand U11261 (N_11261,N_7922,N_9430);
nor U11262 (N_11262,N_9193,N_8214);
or U11263 (N_11263,N_7950,N_8809);
or U11264 (N_11264,N_9564,N_8559);
xnor U11265 (N_11265,N_9349,N_8714);
nor U11266 (N_11266,N_9110,N_8246);
nor U11267 (N_11267,N_7828,N_8156);
or U11268 (N_11268,N_9566,N_7965);
nor U11269 (N_11269,N_9492,N_9907);
xnor U11270 (N_11270,N_7666,N_9417);
or U11271 (N_11271,N_8355,N_8110);
or U11272 (N_11272,N_7940,N_7502);
and U11273 (N_11273,N_9922,N_8868);
or U11274 (N_11274,N_9143,N_9117);
nand U11275 (N_11275,N_9383,N_8814);
xor U11276 (N_11276,N_8400,N_8104);
and U11277 (N_11277,N_8518,N_7696);
nand U11278 (N_11278,N_8043,N_9656);
or U11279 (N_11279,N_8801,N_9232);
or U11280 (N_11280,N_9214,N_8759);
and U11281 (N_11281,N_9676,N_9821);
or U11282 (N_11282,N_8705,N_7521);
or U11283 (N_11283,N_9780,N_9708);
or U11284 (N_11284,N_8365,N_7566);
or U11285 (N_11285,N_9182,N_9605);
and U11286 (N_11286,N_7880,N_8275);
and U11287 (N_11287,N_9397,N_9051);
nor U11288 (N_11288,N_8327,N_9026);
or U11289 (N_11289,N_8673,N_8925);
xnor U11290 (N_11290,N_9369,N_8131);
nand U11291 (N_11291,N_8237,N_9498);
nand U11292 (N_11292,N_9310,N_8897);
nor U11293 (N_11293,N_9266,N_8722);
and U11294 (N_11294,N_7798,N_9539);
xnor U11295 (N_11295,N_8026,N_8402);
xnor U11296 (N_11296,N_8995,N_7914);
xnor U11297 (N_11297,N_9507,N_9172);
and U11298 (N_11298,N_7976,N_8313);
or U11299 (N_11299,N_8137,N_8023);
or U11300 (N_11300,N_9967,N_8232);
and U11301 (N_11301,N_8130,N_7749);
or U11302 (N_11302,N_9988,N_8691);
or U11303 (N_11303,N_9101,N_8798);
xnor U11304 (N_11304,N_9312,N_9669);
nor U11305 (N_11305,N_8529,N_9586);
nand U11306 (N_11306,N_8818,N_7683);
xor U11307 (N_11307,N_8350,N_8471);
or U11308 (N_11308,N_8133,N_8735);
or U11309 (N_11309,N_9534,N_9011);
and U11310 (N_11310,N_9744,N_9003);
and U11311 (N_11311,N_8734,N_9098);
nor U11312 (N_11312,N_8895,N_8938);
or U11313 (N_11313,N_8558,N_8402);
or U11314 (N_11314,N_7736,N_8998);
nand U11315 (N_11315,N_9142,N_7688);
xnor U11316 (N_11316,N_8937,N_7935);
nor U11317 (N_11317,N_7743,N_8935);
nor U11318 (N_11318,N_9816,N_7830);
or U11319 (N_11319,N_9075,N_7800);
nor U11320 (N_11320,N_8973,N_7625);
nand U11321 (N_11321,N_8833,N_8257);
xnor U11322 (N_11322,N_8537,N_7822);
nand U11323 (N_11323,N_7855,N_9735);
nor U11324 (N_11324,N_7829,N_9234);
and U11325 (N_11325,N_9880,N_8299);
xnor U11326 (N_11326,N_8000,N_8294);
or U11327 (N_11327,N_9319,N_7708);
and U11328 (N_11328,N_7818,N_7849);
or U11329 (N_11329,N_8482,N_7573);
and U11330 (N_11330,N_8183,N_9337);
and U11331 (N_11331,N_9008,N_7761);
or U11332 (N_11332,N_7860,N_8065);
or U11333 (N_11333,N_8799,N_8899);
nor U11334 (N_11334,N_9622,N_9889);
xnor U11335 (N_11335,N_9780,N_7848);
or U11336 (N_11336,N_9364,N_8763);
nand U11337 (N_11337,N_8184,N_9782);
xor U11338 (N_11338,N_9835,N_9573);
nand U11339 (N_11339,N_9461,N_7988);
and U11340 (N_11340,N_9907,N_8971);
or U11341 (N_11341,N_9040,N_9085);
nor U11342 (N_11342,N_7689,N_9412);
xor U11343 (N_11343,N_8508,N_9880);
nand U11344 (N_11344,N_9791,N_7740);
and U11345 (N_11345,N_9875,N_9589);
nor U11346 (N_11346,N_9429,N_9153);
and U11347 (N_11347,N_7624,N_8718);
or U11348 (N_11348,N_8196,N_8316);
xnor U11349 (N_11349,N_9761,N_8403);
or U11350 (N_11350,N_7632,N_7841);
or U11351 (N_11351,N_9584,N_7637);
nor U11352 (N_11352,N_9396,N_8323);
nor U11353 (N_11353,N_8507,N_7994);
and U11354 (N_11354,N_9149,N_9083);
nand U11355 (N_11355,N_9333,N_8693);
nor U11356 (N_11356,N_8235,N_8048);
nand U11357 (N_11357,N_9050,N_8866);
and U11358 (N_11358,N_9215,N_9571);
xor U11359 (N_11359,N_7984,N_9760);
nand U11360 (N_11360,N_9420,N_8325);
and U11361 (N_11361,N_9516,N_9463);
nand U11362 (N_11362,N_9779,N_9443);
or U11363 (N_11363,N_7835,N_8517);
nor U11364 (N_11364,N_7839,N_9826);
or U11365 (N_11365,N_9768,N_8103);
nand U11366 (N_11366,N_8915,N_8298);
nand U11367 (N_11367,N_8929,N_7782);
xor U11368 (N_11368,N_9152,N_9515);
and U11369 (N_11369,N_8117,N_7766);
nor U11370 (N_11370,N_8281,N_8157);
and U11371 (N_11371,N_9570,N_8220);
and U11372 (N_11372,N_8080,N_8384);
and U11373 (N_11373,N_8674,N_9954);
nand U11374 (N_11374,N_7688,N_8345);
or U11375 (N_11375,N_8718,N_8067);
nor U11376 (N_11376,N_9316,N_9447);
or U11377 (N_11377,N_8409,N_8291);
nor U11378 (N_11378,N_7524,N_7936);
and U11379 (N_11379,N_7988,N_7738);
xor U11380 (N_11380,N_9496,N_8064);
nor U11381 (N_11381,N_8900,N_7831);
and U11382 (N_11382,N_9314,N_8756);
xor U11383 (N_11383,N_9298,N_7758);
and U11384 (N_11384,N_9289,N_9115);
or U11385 (N_11385,N_9284,N_9545);
or U11386 (N_11386,N_9851,N_8472);
nand U11387 (N_11387,N_8042,N_8299);
or U11388 (N_11388,N_8819,N_8410);
nand U11389 (N_11389,N_8419,N_8435);
or U11390 (N_11390,N_8869,N_8740);
nand U11391 (N_11391,N_8400,N_9180);
nor U11392 (N_11392,N_8344,N_7670);
nand U11393 (N_11393,N_8944,N_8472);
or U11394 (N_11394,N_8541,N_9254);
nor U11395 (N_11395,N_9134,N_8229);
nand U11396 (N_11396,N_9384,N_9210);
xor U11397 (N_11397,N_9124,N_9694);
nand U11398 (N_11398,N_9345,N_8203);
nor U11399 (N_11399,N_8771,N_8433);
nor U11400 (N_11400,N_9023,N_9434);
nor U11401 (N_11401,N_9336,N_9536);
xor U11402 (N_11402,N_8509,N_8287);
nor U11403 (N_11403,N_9233,N_7524);
nor U11404 (N_11404,N_9234,N_9995);
nor U11405 (N_11405,N_8141,N_9526);
nand U11406 (N_11406,N_8708,N_9975);
xnor U11407 (N_11407,N_8087,N_8095);
or U11408 (N_11408,N_9067,N_8090);
or U11409 (N_11409,N_8302,N_8513);
and U11410 (N_11410,N_7736,N_8169);
or U11411 (N_11411,N_7851,N_8911);
xor U11412 (N_11412,N_9402,N_9141);
nand U11413 (N_11413,N_8014,N_9991);
xor U11414 (N_11414,N_8419,N_9385);
or U11415 (N_11415,N_9427,N_8254);
and U11416 (N_11416,N_9989,N_8079);
nand U11417 (N_11417,N_8940,N_9489);
nand U11418 (N_11418,N_7971,N_8772);
xor U11419 (N_11419,N_9968,N_8800);
nor U11420 (N_11420,N_8794,N_7713);
nor U11421 (N_11421,N_9481,N_9614);
xnor U11422 (N_11422,N_8556,N_8509);
nor U11423 (N_11423,N_9064,N_7877);
xor U11424 (N_11424,N_9221,N_8722);
nand U11425 (N_11425,N_8889,N_9267);
nor U11426 (N_11426,N_8870,N_7669);
or U11427 (N_11427,N_8211,N_8649);
nand U11428 (N_11428,N_9144,N_8900);
or U11429 (N_11429,N_7761,N_9275);
and U11430 (N_11430,N_9978,N_9135);
nand U11431 (N_11431,N_8104,N_8279);
and U11432 (N_11432,N_8030,N_8401);
nor U11433 (N_11433,N_8522,N_7710);
nor U11434 (N_11434,N_9565,N_9436);
or U11435 (N_11435,N_7928,N_8138);
nand U11436 (N_11436,N_8516,N_9875);
or U11437 (N_11437,N_8063,N_8088);
and U11438 (N_11438,N_8795,N_9803);
or U11439 (N_11439,N_9575,N_8341);
nand U11440 (N_11440,N_7526,N_9065);
and U11441 (N_11441,N_7942,N_9562);
or U11442 (N_11442,N_7785,N_9943);
nand U11443 (N_11443,N_8700,N_7926);
nand U11444 (N_11444,N_8232,N_8655);
xor U11445 (N_11445,N_9589,N_8686);
nor U11446 (N_11446,N_9286,N_8783);
xnor U11447 (N_11447,N_9031,N_8089);
nand U11448 (N_11448,N_9278,N_8613);
nor U11449 (N_11449,N_9394,N_8572);
xnor U11450 (N_11450,N_7951,N_8899);
nand U11451 (N_11451,N_9225,N_8272);
nand U11452 (N_11452,N_8742,N_9359);
and U11453 (N_11453,N_8190,N_7568);
xor U11454 (N_11454,N_9247,N_8501);
nor U11455 (N_11455,N_8537,N_8635);
nor U11456 (N_11456,N_8071,N_9197);
nor U11457 (N_11457,N_9922,N_9245);
nor U11458 (N_11458,N_8601,N_9697);
xnor U11459 (N_11459,N_8352,N_9612);
nand U11460 (N_11460,N_8567,N_7969);
nand U11461 (N_11461,N_9795,N_9003);
xnor U11462 (N_11462,N_9425,N_9548);
nand U11463 (N_11463,N_7870,N_8545);
or U11464 (N_11464,N_8847,N_8953);
or U11465 (N_11465,N_8511,N_7654);
nor U11466 (N_11466,N_7975,N_7967);
nand U11467 (N_11467,N_9925,N_9561);
and U11468 (N_11468,N_8255,N_8186);
and U11469 (N_11469,N_9580,N_9758);
nand U11470 (N_11470,N_8239,N_7840);
xor U11471 (N_11471,N_8666,N_8363);
nand U11472 (N_11472,N_7592,N_8652);
nor U11473 (N_11473,N_9997,N_9427);
nor U11474 (N_11474,N_7886,N_8847);
and U11475 (N_11475,N_9028,N_8360);
xnor U11476 (N_11476,N_9041,N_8930);
and U11477 (N_11477,N_7661,N_8245);
nand U11478 (N_11478,N_8575,N_9046);
nand U11479 (N_11479,N_9966,N_7747);
xnor U11480 (N_11480,N_9036,N_9307);
and U11481 (N_11481,N_8715,N_7619);
and U11482 (N_11482,N_9931,N_9544);
or U11483 (N_11483,N_8375,N_8336);
and U11484 (N_11484,N_9594,N_9993);
xor U11485 (N_11485,N_9912,N_9086);
xnor U11486 (N_11486,N_7513,N_7808);
nand U11487 (N_11487,N_8073,N_9071);
and U11488 (N_11488,N_9078,N_7809);
nor U11489 (N_11489,N_9683,N_8274);
xnor U11490 (N_11490,N_9808,N_8030);
and U11491 (N_11491,N_8538,N_8288);
and U11492 (N_11492,N_9075,N_8514);
xor U11493 (N_11493,N_9376,N_9020);
and U11494 (N_11494,N_8795,N_8561);
nand U11495 (N_11495,N_8087,N_9530);
xnor U11496 (N_11496,N_8560,N_9417);
and U11497 (N_11497,N_9958,N_7867);
and U11498 (N_11498,N_9485,N_9794);
or U11499 (N_11499,N_9406,N_9940);
and U11500 (N_11500,N_9473,N_7509);
xor U11501 (N_11501,N_8212,N_8649);
nor U11502 (N_11502,N_9166,N_8680);
or U11503 (N_11503,N_8054,N_9575);
xor U11504 (N_11504,N_8018,N_7502);
nor U11505 (N_11505,N_7560,N_9343);
or U11506 (N_11506,N_8894,N_8441);
nand U11507 (N_11507,N_9093,N_7969);
or U11508 (N_11508,N_9880,N_9540);
or U11509 (N_11509,N_9928,N_8928);
and U11510 (N_11510,N_8561,N_7889);
nand U11511 (N_11511,N_8896,N_9953);
nor U11512 (N_11512,N_8633,N_9902);
xnor U11513 (N_11513,N_9440,N_8841);
nor U11514 (N_11514,N_9276,N_8554);
xor U11515 (N_11515,N_9970,N_9050);
nand U11516 (N_11516,N_8310,N_9233);
nand U11517 (N_11517,N_8141,N_9833);
xnor U11518 (N_11518,N_8868,N_7913);
xor U11519 (N_11519,N_8995,N_9077);
nand U11520 (N_11520,N_9199,N_8858);
and U11521 (N_11521,N_8834,N_9928);
and U11522 (N_11522,N_9283,N_9923);
xnor U11523 (N_11523,N_9954,N_9645);
or U11524 (N_11524,N_7542,N_9611);
xor U11525 (N_11525,N_8384,N_9930);
and U11526 (N_11526,N_9874,N_9871);
nor U11527 (N_11527,N_8615,N_7812);
or U11528 (N_11528,N_9765,N_8860);
xor U11529 (N_11529,N_8048,N_8003);
nor U11530 (N_11530,N_8571,N_7540);
and U11531 (N_11531,N_7572,N_8010);
or U11532 (N_11532,N_7593,N_7664);
nor U11533 (N_11533,N_9707,N_7772);
and U11534 (N_11534,N_8579,N_7914);
and U11535 (N_11535,N_8047,N_8029);
and U11536 (N_11536,N_9223,N_7897);
nor U11537 (N_11537,N_9528,N_8245);
nand U11538 (N_11538,N_8096,N_8578);
xor U11539 (N_11539,N_8044,N_8896);
or U11540 (N_11540,N_9118,N_8190);
and U11541 (N_11541,N_8419,N_7638);
xnor U11542 (N_11542,N_7924,N_8324);
nor U11543 (N_11543,N_9239,N_8617);
xor U11544 (N_11544,N_8622,N_8605);
and U11545 (N_11545,N_7956,N_8431);
nand U11546 (N_11546,N_9559,N_9194);
or U11547 (N_11547,N_9286,N_9729);
and U11548 (N_11548,N_8627,N_7687);
xor U11549 (N_11549,N_7659,N_8022);
nand U11550 (N_11550,N_7707,N_8412);
nand U11551 (N_11551,N_9537,N_8729);
nand U11552 (N_11552,N_9704,N_9076);
and U11553 (N_11553,N_9167,N_9063);
nand U11554 (N_11554,N_8006,N_8851);
nand U11555 (N_11555,N_8453,N_9658);
or U11556 (N_11556,N_9373,N_8158);
and U11557 (N_11557,N_9343,N_8766);
xnor U11558 (N_11558,N_8855,N_8479);
nor U11559 (N_11559,N_9439,N_8564);
or U11560 (N_11560,N_9674,N_8707);
or U11561 (N_11561,N_9974,N_9055);
nor U11562 (N_11562,N_8150,N_9909);
or U11563 (N_11563,N_7955,N_8013);
and U11564 (N_11564,N_7500,N_8114);
nand U11565 (N_11565,N_8303,N_9851);
nand U11566 (N_11566,N_7966,N_8543);
nor U11567 (N_11567,N_9335,N_8287);
xor U11568 (N_11568,N_8326,N_8885);
nor U11569 (N_11569,N_7894,N_7504);
and U11570 (N_11570,N_9115,N_8049);
xor U11571 (N_11571,N_9659,N_9182);
xor U11572 (N_11572,N_8552,N_7998);
or U11573 (N_11573,N_9608,N_9141);
nor U11574 (N_11574,N_9019,N_8900);
or U11575 (N_11575,N_8313,N_7712);
and U11576 (N_11576,N_7629,N_7908);
nor U11577 (N_11577,N_8660,N_9796);
or U11578 (N_11578,N_7657,N_9931);
nor U11579 (N_11579,N_9304,N_8517);
nand U11580 (N_11580,N_9483,N_7960);
nor U11581 (N_11581,N_7688,N_8185);
xnor U11582 (N_11582,N_8017,N_8545);
and U11583 (N_11583,N_8633,N_8905);
nand U11584 (N_11584,N_7510,N_7799);
xor U11585 (N_11585,N_8451,N_8743);
and U11586 (N_11586,N_9598,N_9043);
or U11587 (N_11587,N_8369,N_7518);
nor U11588 (N_11588,N_9674,N_8514);
nand U11589 (N_11589,N_8684,N_9655);
and U11590 (N_11590,N_8123,N_9724);
and U11591 (N_11591,N_9468,N_8661);
and U11592 (N_11592,N_8940,N_9480);
nand U11593 (N_11593,N_8717,N_7690);
nor U11594 (N_11594,N_8178,N_8371);
nand U11595 (N_11595,N_8664,N_9088);
and U11596 (N_11596,N_9288,N_9084);
xnor U11597 (N_11597,N_8210,N_9393);
and U11598 (N_11598,N_7965,N_7590);
and U11599 (N_11599,N_9031,N_7842);
and U11600 (N_11600,N_9730,N_7554);
xor U11601 (N_11601,N_8978,N_8434);
xnor U11602 (N_11602,N_9549,N_8958);
and U11603 (N_11603,N_8839,N_8246);
or U11604 (N_11604,N_8674,N_8947);
nand U11605 (N_11605,N_8414,N_8625);
nand U11606 (N_11606,N_8856,N_7756);
or U11607 (N_11607,N_7715,N_8003);
nor U11608 (N_11608,N_9463,N_7605);
nand U11609 (N_11609,N_7596,N_7756);
nand U11610 (N_11610,N_9064,N_8037);
or U11611 (N_11611,N_8508,N_9286);
xnor U11612 (N_11612,N_8335,N_9764);
or U11613 (N_11613,N_9586,N_9605);
or U11614 (N_11614,N_8916,N_7955);
nor U11615 (N_11615,N_8985,N_8164);
nor U11616 (N_11616,N_9159,N_7833);
xor U11617 (N_11617,N_8477,N_7535);
nor U11618 (N_11618,N_9532,N_7530);
nor U11619 (N_11619,N_8117,N_9505);
nand U11620 (N_11620,N_9882,N_8501);
or U11621 (N_11621,N_7724,N_9472);
xnor U11622 (N_11622,N_9936,N_7546);
or U11623 (N_11623,N_8234,N_9225);
and U11624 (N_11624,N_9100,N_9643);
xor U11625 (N_11625,N_9838,N_8961);
nand U11626 (N_11626,N_9577,N_8292);
or U11627 (N_11627,N_8321,N_8891);
or U11628 (N_11628,N_9938,N_7817);
xnor U11629 (N_11629,N_8812,N_7685);
nand U11630 (N_11630,N_8045,N_8545);
nor U11631 (N_11631,N_9642,N_8720);
xnor U11632 (N_11632,N_8718,N_8256);
nor U11633 (N_11633,N_8145,N_8126);
nor U11634 (N_11634,N_9010,N_8020);
xor U11635 (N_11635,N_9575,N_9934);
xor U11636 (N_11636,N_8868,N_9251);
nor U11637 (N_11637,N_8622,N_9096);
xnor U11638 (N_11638,N_9406,N_8091);
or U11639 (N_11639,N_9579,N_7517);
and U11640 (N_11640,N_8130,N_9406);
xor U11641 (N_11641,N_7664,N_8353);
or U11642 (N_11642,N_9766,N_8664);
and U11643 (N_11643,N_7963,N_8016);
or U11644 (N_11644,N_9695,N_8971);
nand U11645 (N_11645,N_9430,N_7738);
or U11646 (N_11646,N_9640,N_8580);
nand U11647 (N_11647,N_9435,N_7659);
nor U11648 (N_11648,N_9423,N_9672);
xnor U11649 (N_11649,N_8642,N_9755);
xnor U11650 (N_11650,N_8675,N_9094);
and U11651 (N_11651,N_7624,N_8848);
and U11652 (N_11652,N_8625,N_7928);
or U11653 (N_11653,N_8342,N_9325);
nor U11654 (N_11654,N_9160,N_8273);
nand U11655 (N_11655,N_8871,N_8714);
nor U11656 (N_11656,N_7733,N_8800);
xnor U11657 (N_11657,N_9351,N_8683);
xor U11658 (N_11658,N_9454,N_8815);
nor U11659 (N_11659,N_7801,N_7515);
nor U11660 (N_11660,N_7671,N_8172);
or U11661 (N_11661,N_7679,N_9409);
and U11662 (N_11662,N_9473,N_9794);
nand U11663 (N_11663,N_7796,N_8136);
or U11664 (N_11664,N_7666,N_8880);
nor U11665 (N_11665,N_9012,N_8984);
xor U11666 (N_11666,N_9179,N_7991);
or U11667 (N_11667,N_7696,N_7676);
nor U11668 (N_11668,N_9056,N_9300);
nor U11669 (N_11669,N_8836,N_9391);
nor U11670 (N_11670,N_9547,N_8205);
nand U11671 (N_11671,N_8419,N_9360);
or U11672 (N_11672,N_9006,N_8421);
nor U11673 (N_11673,N_8568,N_9897);
nand U11674 (N_11674,N_8109,N_8853);
or U11675 (N_11675,N_8638,N_9837);
and U11676 (N_11676,N_7606,N_9492);
nor U11677 (N_11677,N_8095,N_8029);
nand U11678 (N_11678,N_7565,N_8630);
nand U11679 (N_11679,N_8060,N_7640);
or U11680 (N_11680,N_9588,N_9490);
or U11681 (N_11681,N_9252,N_9583);
or U11682 (N_11682,N_9563,N_9001);
or U11683 (N_11683,N_7622,N_9022);
or U11684 (N_11684,N_8698,N_8867);
nor U11685 (N_11685,N_8528,N_9860);
xor U11686 (N_11686,N_8066,N_9321);
nand U11687 (N_11687,N_8557,N_7737);
xor U11688 (N_11688,N_9205,N_9226);
nand U11689 (N_11689,N_9772,N_7910);
nor U11690 (N_11690,N_7917,N_8786);
nand U11691 (N_11691,N_8679,N_7839);
nand U11692 (N_11692,N_9028,N_7726);
nand U11693 (N_11693,N_8250,N_9233);
nor U11694 (N_11694,N_8022,N_9930);
nor U11695 (N_11695,N_8830,N_9847);
and U11696 (N_11696,N_8131,N_9861);
xnor U11697 (N_11697,N_8570,N_9513);
and U11698 (N_11698,N_8872,N_9616);
or U11699 (N_11699,N_9361,N_9370);
nand U11700 (N_11700,N_8798,N_8721);
and U11701 (N_11701,N_7584,N_9550);
and U11702 (N_11702,N_9398,N_8656);
nor U11703 (N_11703,N_7638,N_9847);
xor U11704 (N_11704,N_8174,N_7552);
nor U11705 (N_11705,N_9497,N_9008);
or U11706 (N_11706,N_8311,N_9593);
xnor U11707 (N_11707,N_7741,N_8392);
nand U11708 (N_11708,N_8569,N_8496);
and U11709 (N_11709,N_9349,N_9431);
and U11710 (N_11710,N_8772,N_8793);
and U11711 (N_11711,N_9519,N_8830);
and U11712 (N_11712,N_8814,N_8962);
and U11713 (N_11713,N_8680,N_8441);
nand U11714 (N_11714,N_7731,N_7681);
nor U11715 (N_11715,N_7861,N_9536);
and U11716 (N_11716,N_8205,N_8368);
and U11717 (N_11717,N_9332,N_9579);
xnor U11718 (N_11718,N_8866,N_8475);
nor U11719 (N_11719,N_7882,N_9196);
nor U11720 (N_11720,N_9087,N_7710);
or U11721 (N_11721,N_8131,N_8574);
nor U11722 (N_11722,N_9303,N_8886);
and U11723 (N_11723,N_9315,N_8693);
and U11724 (N_11724,N_9874,N_8574);
xnor U11725 (N_11725,N_9520,N_9785);
xor U11726 (N_11726,N_9052,N_7848);
nand U11727 (N_11727,N_8076,N_9300);
nand U11728 (N_11728,N_9983,N_8187);
or U11729 (N_11729,N_8215,N_9960);
or U11730 (N_11730,N_7888,N_8029);
xor U11731 (N_11731,N_7526,N_8419);
nor U11732 (N_11732,N_7514,N_8809);
nor U11733 (N_11733,N_8541,N_8902);
or U11734 (N_11734,N_7511,N_9023);
xnor U11735 (N_11735,N_7550,N_9197);
and U11736 (N_11736,N_7857,N_8916);
nand U11737 (N_11737,N_9484,N_9311);
nor U11738 (N_11738,N_8117,N_8040);
nor U11739 (N_11739,N_9149,N_9071);
and U11740 (N_11740,N_9393,N_8375);
or U11741 (N_11741,N_9731,N_9516);
xor U11742 (N_11742,N_8840,N_9678);
xor U11743 (N_11743,N_7875,N_7655);
nand U11744 (N_11744,N_8699,N_9499);
or U11745 (N_11745,N_7768,N_8779);
and U11746 (N_11746,N_8669,N_9275);
nor U11747 (N_11747,N_9513,N_9984);
xnor U11748 (N_11748,N_9330,N_9034);
and U11749 (N_11749,N_8985,N_9896);
or U11750 (N_11750,N_9355,N_8782);
nor U11751 (N_11751,N_8845,N_9798);
xnor U11752 (N_11752,N_7784,N_7729);
nand U11753 (N_11753,N_8038,N_9331);
and U11754 (N_11754,N_7500,N_8208);
and U11755 (N_11755,N_8372,N_8717);
and U11756 (N_11756,N_9373,N_9038);
and U11757 (N_11757,N_8387,N_9970);
xnor U11758 (N_11758,N_8581,N_7882);
or U11759 (N_11759,N_8892,N_8218);
nor U11760 (N_11760,N_9939,N_7809);
nor U11761 (N_11761,N_8436,N_9404);
xor U11762 (N_11762,N_7638,N_8874);
xor U11763 (N_11763,N_9544,N_8275);
xnor U11764 (N_11764,N_8545,N_7747);
and U11765 (N_11765,N_8136,N_9016);
xnor U11766 (N_11766,N_7763,N_9538);
nor U11767 (N_11767,N_9122,N_7777);
or U11768 (N_11768,N_7961,N_9656);
and U11769 (N_11769,N_9193,N_8885);
or U11770 (N_11770,N_7532,N_8274);
xnor U11771 (N_11771,N_9565,N_9859);
nand U11772 (N_11772,N_8489,N_8257);
nor U11773 (N_11773,N_8275,N_9128);
xnor U11774 (N_11774,N_9332,N_8402);
nor U11775 (N_11775,N_7649,N_8825);
or U11776 (N_11776,N_9909,N_8538);
or U11777 (N_11777,N_7594,N_9261);
or U11778 (N_11778,N_9030,N_9200);
nand U11779 (N_11779,N_9565,N_7977);
or U11780 (N_11780,N_9007,N_9287);
nand U11781 (N_11781,N_8434,N_8990);
or U11782 (N_11782,N_9882,N_9248);
and U11783 (N_11783,N_9728,N_9518);
or U11784 (N_11784,N_9841,N_8960);
or U11785 (N_11785,N_9797,N_8207);
xnor U11786 (N_11786,N_8789,N_9481);
nor U11787 (N_11787,N_8347,N_9784);
or U11788 (N_11788,N_9788,N_7625);
and U11789 (N_11789,N_7857,N_7720);
or U11790 (N_11790,N_9083,N_9680);
nand U11791 (N_11791,N_8263,N_8535);
and U11792 (N_11792,N_9040,N_9438);
or U11793 (N_11793,N_9493,N_8427);
nor U11794 (N_11794,N_8347,N_7811);
nand U11795 (N_11795,N_9364,N_8732);
nor U11796 (N_11796,N_8208,N_8388);
or U11797 (N_11797,N_8851,N_8645);
or U11798 (N_11798,N_8651,N_8018);
and U11799 (N_11799,N_9150,N_8395);
nand U11800 (N_11800,N_8158,N_8923);
nand U11801 (N_11801,N_9118,N_7730);
nand U11802 (N_11802,N_7790,N_9794);
nand U11803 (N_11803,N_9207,N_9570);
or U11804 (N_11804,N_9556,N_9146);
nand U11805 (N_11805,N_8954,N_8317);
nand U11806 (N_11806,N_8579,N_9878);
xnor U11807 (N_11807,N_9462,N_7739);
nor U11808 (N_11808,N_9079,N_8613);
or U11809 (N_11809,N_9871,N_9613);
xor U11810 (N_11810,N_8420,N_7808);
and U11811 (N_11811,N_7951,N_8454);
xnor U11812 (N_11812,N_8021,N_9517);
nand U11813 (N_11813,N_9437,N_7908);
nand U11814 (N_11814,N_9932,N_9197);
and U11815 (N_11815,N_7772,N_8413);
and U11816 (N_11816,N_8592,N_7838);
xor U11817 (N_11817,N_7759,N_9622);
nand U11818 (N_11818,N_9697,N_8657);
and U11819 (N_11819,N_9450,N_8739);
nand U11820 (N_11820,N_7919,N_9058);
nand U11821 (N_11821,N_8563,N_7986);
and U11822 (N_11822,N_7562,N_7833);
xor U11823 (N_11823,N_8909,N_8227);
nor U11824 (N_11824,N_8317,N_8714);
nor U11825 (N_11825,N_9044,N_7940);
or U11826 (N_11826,N_8326,N_8000);
or U11827 (N_11827,N_9707,N_8400);
nand U11828 (N_11828,N_9730,N_9482);
and U11829 (N_11829,N_7572,N_9870);
nor U11830 (N_11830,N_9876,N_9769);
nor U11831 (N_11831,N_9988,N_8296);
xnor U11832 (N_11832,N_7741,N_9183);
or U11833 (N_11833,N_9315,N_9921);
nand U11834 (N_11834,N_8632,N_9307);
nor U11835 (N_11835,N_9418,N_8850);
nand U11836 (N_11836,N_8226,N_7872);
and U11837 (N_11837,N_8598,N_8051);
xnor U11838 (N_11838,N_8766,N_7507);
nand U11839 (N_11839,N_8730,N_8055);
nor U11840 (N_11840,N_8204,N_9390);
and U11841 (N_11841,N_8491,N_8673);
nand U11842 (N_11842,N_9311,N_8737);
nand U11843 (N_11843,N_8149,N_8996);
nor U11844 (N_11844,N_8395,N_7932);
nand U11845 (N_11845,N_8472,N_8854);
and U11846 (N_11846,N_9738,N_7833);
or U11847 (N_11847,N_8644,N_8308);
xor U11848 (N_11848,N_7681,N_8601);
nand U11849 (N_11849,N_9697,N_9715);
xor U11850 (N_11850,N_9429,N_9511);
and U11851 (N_11851,N_9253,N_9473);
nand U11852 (N_11852,N_9340,N_9174);
nor U11853 (N_11853,N_8565,N_9220);
nand U11854 (N_11854,N_8931,N_8282);
and U11855 (N_11855,N_8971,N_9906);
and U11856 (N_11856,N_9757,N_9213);
and U11857 (N_11857,N_8226,N_8375);
and U11858 (N_11858,N_8905,N_8897);
and U11859 (N_11859,N_9903,N_8816);
and U11860 (N_11860,N_8665,N_9139);
xor U11861 (N_11861,N_9541,N_9316);
or U11862 (N_11862,N_8241,N_8019);
nand U11863 (N_11863,N_9153,N_9338);
nor U11864 (N_11864,N_7820,N_8629);
nand U11865 (N_11865,N_9477,N_8695);
and U11866 (N_11866,N_7717,N_8236);
and U11867 (N_11867,N_8730,N_8137);
nor U11868 (N_11868,N_8246,N_8596);
or U11869 (N_11869,N_9641,N_7898);
nand U11870 (N_11870,N_9981,N_9320);
xor U11871 (N_11871,N_9171,N_9070);
xnor U11872 (N_11872,N_8694,N_8673);
or U11873 (N_11873,N_7998,N_8247);
or U11874 (N_11874,N_9496,N_8248);
xor U11875 (N_11875,N_7906,N_7716);
nor U11876 (N_11876,N_9215,N_7713);
or U11877 (N_11877,N_8146,N_8243);
xor U11878 (N_11878,N_9546,N_8887);
nor U11879 (N_11879,N_9331,N_9770);
nand U11880 (N_11880,N_9202,N_8292);
nor U11881 (N_11881,N_8387,N_8406);
xnor U11882 (N_11882,N_8639,N_9553);
or U11883 (N_11883,N_8908,N_9652);
nor U11884 (N_11884,N_8542,N_8992);
and U11885 (N_11885,N_7588,N_8947);
nand U11886 (N_11886,N_8369,N_7918);
or U11887 (N_11887,N_8881,N_7640);
nand U11888 (N_11888,N_8473,N_7803);
or U11889 (N_11889,N_9529,N_8883);
nand U11890 (N_11890,N_9478,N_8982);
nand U11891 (N_11891,N_9614,N_8936);
and U11892 (N_11892,N_7735,N_8347);
or U11893 (N_11893,N_7503,N_7788);
nor U11894 (N_11894,N_7570,N_8260);
nor U11895 (N_11895,N_9083,N_9618);
and U11896 (N_11896,N_9406,N_9211);
xor U11897 (N_11897,N_9599,N_9089);
and U11898 (N_11898,N_8298,N_7762);
nor U11899 (N_11899,N_8635,N_8290);
nor U11900 (N_11900,N_9406,N_9631);
or U11901 (N_11901,N_9977,N_9574);
xnor U11902 (N_11902,N_8823,N_7759);
nand U11903 (N_11903,N_9767,N_8153);
nor U11904 (N_11904,N_9524,N_9453);
nor U11905 (N_11905,N_7586,N_7652);
or U11906 (N_11906,N_8056,N_8263);
and U11907 (N_11907,N_9114,N_8304);
or U11908 (N_11908,N_8944,N_8797);
nor U11909 (N_11909,N_9066,N_8212);
nor U11910 (N_11910,N_7607,N_9587);
nor U11911 (N_11911,N_8137,N_8094);
nor U11912 (N_11912,N_8110,N_9981);
xnor U11913 (N_11913,N_7596,N_7734);
and U11914 (N_11914,N_7576,N_8307);
xor U11915 (N_11915,N_9546,N_7678);
xor U11916 (N_11916,N_9147,N_7636);
nand U11917 (N_11917,N_8072,N_9921);
xor U11918 (N_11918,N_8383,N_7578);
xnor U11919 (N_11919,N_8859,N_9441);
or U11920 (N_11920,N_9501,N_7550);
or U11921 (N_11921,N_8035,N_9696);
and U11922 (N_11922,N_8208,N_9256);
and U11923 (N_11923,N_8744,N_8097);
or U11924 (N_11924,N_7627,N_8522);
nand U11925 (N_11925,N_8105,N_9510);
nor U11926 (N_11926,N_7721,N_9697);
or U11927 (N_11927,N_8739,N_7816);
or U11928 (N_11928,N_7917,N_9865);
and U11929 (N_11929,N_9950,N_8341);
nor U11930 (N_11930,N_9132,N_9946);
and U11931 (N_11931,N_8368,N_7727);
nand U11932 (N_11932,N_7768,N_8519);
and U11933 (N_11933,N_9524,N_9558);
nand U11934 (N_11934,N_9585,N_8030);
or U11935 (N_11935,N_7976,N_9463);
xnor U11936 (N_11936,N_9553,N_7629);
or U11937 (N_11937,N_8595,N_7958);
or U11938 (N_11938,N_9483,N_9773);
and U11939 (N_11939,N_8837,N_8266);
nor U11940 (N_11940,N_9171,N_8429);
nand U11941 (N_11941,N_7794,N_8953);
and U11942 (N_11942,N_8251,N_8637);
or U11943 (N_11943,N_9338,N_8442);
xnor U11944 (N_11944,N_8791,N_9439);
and U11945 (N_11945,N_9110,N_8607);
or U11946 (N_11946,N_8458,N_8431);
or U11947 (N_11947,N_8331,N_9361);
xnor U11948 (N_11948,N_9165,N_9251);
xor U11949 (N_11949,N_8133,N_9274);
nand U11950 (N_11950,N_7703,N_9615);
nor U11951 (N_11951,N_9222,N_8152);
or U11952 (N_11952,N_7662,N_9467);
nor U11953 (N_11953,N_9057,N_8974);
nor U11954 (N_11954,N_7780,N_9311);
nand U11955 (N_11955,N_9050,N_8122);
xnor U11956 (N_11956,N_7604,N_9675);
and U11957 (N_11957,N_8980,N_9809);
nor U11958 (N_11958,N_9507,N_7875);
nand U11959 (N_11959,N_8725,N_8410);
and U11960 (N_11960,N_7834,N_9809);
nand U11961 (N_11961,N_8445,N_8447);
nor U11962 (N_11962,N_8295,N_7899);
nand U11963 (N_11963,N_9723,N_8179);
nor U11964 (N_11964,N_8674,N_9444);
xor U11965 (N_11965,N_9412,N_7645);
nor U11966 (N_11966,N_8970,N_9153);
nor U11967 (N_11967,N_8811,N_9877);
nand U11968 (N_11968,N_7566,N_7629);
xnor U11969 (N_11969,N_9724,N_9322);
nand U11970 (N_11970,N_7694,N_9296);
and U11971 (N_11971,N_8054,N_7770);
nand U11972 (N_11972,N_8655,N_9595);
or U11973 (N_11973,N_7851,N_8859);
xor U11974 (N_11974,N_7848,N_7951);
nor U11975 (N_11975,N_9017,N_8587);
nand U11976 (N_11976,N_9342,N_7839);
and U11977 (N_11977,N_8825,N_8696);
or U11978 (N_11978,N_8288,N_7970);
nand U11979 (N_11979,N_8564,N_7559);
or U11980 (N_11980,N_8530,N_8746);
nor U11981 (N_11981,N_8970,N_7934);
and U11982 (N_11982,N_7927,N_8866);
xor U11983 (N_11983,N_9576,N_8974);
nand U11984 (N_11984,N_8756,N_7714);
or U11985 (N_11985,N_8529,N_7694);
xnor U11986 (N_11986,N_9254,N_7512);
and U11987 (N_11987,N_8091,N_7931);
xor U11988 (N_11988,N_8125,N_8026);
and U11989 (N_11989,N_8072,N_7707);
xor U11990 (N_11990,N_9321,N_8159);
nand U11991 (N_11991,N_9803,N_8448);
or U11992 (N_11992,N_9857,N_8835);
or U11993 (N_11993,N_8192,N_7974);
or U11994 (N_11994,N_8707,N_7586);
nand U11995 (N_11995,N_8154,N_9358);
xnor U11996 (N_11996,N_9525,N_8117);
and U11997 (N_11997,N_9561,N_9483);
and U11998 (N_11998,N_8224,N_8888);
nor U11999 (N_11999,N_9770,N_9199);
or U12000 (N_12000,N_8872,N_7995);
nor U12001 (N_12001,N_9275,N_8256);
or U12002 (N_12002,N_8798,N_7516);
nand U12003 (N_12003,N_9195,N_8393);
and U12004 (N_12004,N_7900,N_9490);
and U12005 (N_12005,N_7728,N_9629);
nor U12006 (N_12006,N_7523,N_7587);
nor U12007 (N_12007,N_8286,N_9624);
or U12008 (N_12008,N_8784,N_9606);
nand U12009 (N_12009,N_9664,N_9075);
or U12010 (N_12010,N_8973,N_9593);
or U12011 (N_12011,N_8396,N_7645);
and U12012 (N_12012,N_8692,N_8723);
xnor U12013 (N_12013,N_8550,N_8307);
nor U12014 (N_12014,N_9085,N_9222);
nor U12015 (N_12015,N_8950,N_8671);
xnor U12016 (N_12016,N_8665,N_8904);
nor U12017 (N_12017,N_8515,N_9647);
xor U12018 (N_12018,N_8101,N_8280);
nand U12019 (N_12019,N_9516,N_8989);
xor U12020 (N_12020,N_8461,N_8867);
nand U12021 (N_12021,N_8829,N_8573);
xor U12022 (N_12022,N_8850,N_8790);
nor U12023 (N_12023,N_9858,N_8413);
or U12024 (N_12024,N_7727,N_9213);
or U12025 (N_12025,N_9968,N_9153);
xor U12026 (N_12026,N_8163,N_8696);
or U12027 (N_12027,N_7510,N_8202);
nor U12028 (N_12028,N_7543,N_9087);
xor U12029 (N_12029,N_8284,N_9565);
and U12030 (N_12030,N_9017,N_8295);
and U12031 (N_12031,N_9369,N_8201);
nor U12032 (N_12032,N_9678,N_9222);
xor U12033 (N_12033,N_9442,N_8317);
and U12034 (N_12034,N_8884,N_9144);
xor U12035 (N_12035,N_8071,N_9789);
nand U12036 (N_12036,N_7651,N_7874);
nor U12037 (N_12037,N_7500,N_9731);
nor U12038 (N_12038,N_9412,N_8407);
and U12039 (N_12039,N_8615,N_9779);
and U12040 (N_12040,N_9423,N_7775);
and U12041 (N_12041,N_8370,N_9590);
nor U12042 (N_12042,N_8765,N_9604);
xor U12043 (N_12043,N_8452,N_8541);
xor U12044 (N_12044,N_9373,N_7767);
and U12045 (N_12045,N_7855,N_7678);
xor U12046 (N_12046,N_9161,N_8438);
or U12047 (N_12047,N_7707,N_9207);
nor U12048 (N_12048,N_7898,N_8127);
xor U12049 (N_12049,N_8232,N_9844);
nor U12050 (N_12050,N_8273,N_8074);
and U12051 (N_12051,N_7639,N_8094);
nand U12052 (N_12052,N_8341,N_9240);
and U12053 (N_12053,N_9318,N_7784);
or U12054 (N_12054,N_9731,N_8849);
and U12055 (N_12055,N_9214,N_8435);
or U12056 (N_12056,N_8757,N_8440);
and U12057 (N_12057,N_8468,N_8929);
nor U12058 (N_12058,N_9657,N_7857);
and U12059 (N_12059,N_9749,N_7867);
xnor U12060 (N_12060,N_8712,N_9595);
xnor U12061 (N_12061,N_9564,N_8456);
xor U12062 (N_12062,N_7710,N_9233);
and U12063 (N_12063,N_9819,N_8952);
xor U12064 (N_12064,N_9046,N_8550);
and U12065 (N_12065,N_9198,N_8480);
or U12066 (N_12066,N_7740,N_8822);
or U12067 (N_12067,N_7611,N_9850);
nand U12068 (N_12068,N_8393,N_9969);
or U12069 (N_12069,N_9983,N_8266);
xor U12070 (N_12070,N_8174,N_9874);
nor U12071 (N_12071,N_9825,N_8567);
nand U12072 (N_12072,N_7992,N_9452);
nor U12073 (N_12073,N_7524,N_9881);
and U12074 (N_12074,N_7697,N_8410);
or U12075 (N_12075,N_8944,N_9957);
nand U12076 (N_12076,N_9563,N_7538);
and U12077 (N_12077,N_7665,N_9483);
nand U12078 (N_12078,N_9455,N_9894);
nand U12079 (N_12079,N_8142,N_7563);
nand U12080 (N_12080,N_8894,N_9322);
nor U12081 (N_12081,N_8497,N_9954);
nand U12082 (N_12082,N_8073,N_8142);
and U12083 (N_12083,N_8679,N_7751);
and U12084 (N_12084,N_9594,N_9357);
and U12085 (N_12085,N_9423,N_8161);
or U12086 (N_12086,N_9527,N_7593);
and U12087 (N_12087,N_8213,N_7538);
or U12088 (N_12088,N_9632,N_7749);
or U12089 (N_12089,N_9723,N_8544);
or U12090 (N_12090,N_8181,N_8480);
xor U12091 (N_12091,N_9361,N_7953);
nand U12092 (N_12092,N_9482,N_7590);
nor U12093 (N_12093,N_7986,N_9780);
nand U12094 (N_12094,N_8815,N_8686);
nor U12095 (N_12095,N_9028,N_7544);
nand U12096 (N_12096,N_7588,N_9131);
nand U12097 (N_12097,N_8580,N_8476);
or U12098 (N_12098,N_7921,N_8042);
xor U12099 (N_12099,N_8630,N_8789);
and U12100 (N_12100,N_8174,N_9185);
or U12101 (N_12101,N_8596,N_9944);
or U12102 (N_12102,N_8959,N_9910);
xnor U12103 (N_12103,N_7647,N_7569);
xor U12104 (N_12104,N_7665,N_9290);
xor U12105 (N_12105,N_7727,N_9946);
or U12106 (N_12106,N_7587,N_8539);
nor U12107 (N_12107,N_9943,N_8397);
xor U12108 (N_12108,N_9006,N_9415);
nor U12109 (N_12109,N_8027,N_8266);
nand U12110 (N_12110,N_9129,N_7609);
xor U12111 (N_12111,N_8151,N_8817);
or U12112 (N_12112,N_7597,N_9961);
or U12113 (N_12113,N_9299,N_9310);
nand U12114 (N_12114,N_9699,N_9347);
or U12115 (N_12115,N_9690,N_8558);
xor U12116 (N_12116,N_9504,N_9959);
or U12117 (N_12117,N_9083,N_9462);
xnor U12118 (N_12118,N_9172,N_8673);
nor U12119 (N_12119,N_8524,N_9252);
and U12120 (N_12120,N_9260,N_8610);
nand U12121 (N_12121,N_8367,N_8321);
nor U12122 (N_12122,N_9727,N_9393);
or U12123 (N_12123,N_7862,N_7571);
or U12124 (N_12124,N_7660,N_8659);
xnor U12125 (N_12125,N_7954,N_8483);
nor U12126 (N_12126,N_8381,N_8033);
or U12127 (N_12127,N_7656,N_8473);
xor U12128 (N_12128,N_8158,N_8732);
nand U12129 (N_12129,N_9964,N_9253);
or U12130 (N_12130,N_7532,N_7885);
xor U12131 (N_12131,N_7747,N_9239);
nor U12132 (N_12132,N_8433,N_7792);
or U12133 (N_12133,N_8731,N_9539);
xor U12134 (N_12134,N_8500,N_9537);
nor U12135 (N_12135,N_8375,N_8737);
and U12136 (N_12136,N_9390,N_7977);
xor U12137 (N_12137,N_9619,N_7618);
xor U12138 (N_12138,N_8081,N_9065);
and U12139 (N_12139,N_9777,N_8363);
and U12140 (N_12140,N_9427,N_9565);
xor U12141 (N_12141,N_9640,N_9818);
and U12142 (N_12142,N_9940,N_7968);
or U12143 (N_12143,N_8148,N_9329);
and U12144 (N_12144,N_9798,N_9461);
xor U12145 (N_12145,N_8244,N_8328);
or U12146 (N_12146,N_7655,N_8667);
and U12147 (N_12147,N_9485,N_9149);
nand U12148 (N_12148,N_9418,N_8223);
xnor U12149 (N_12149,N_9633,N_7675);
nand U12150 (N_12150,N_8231,N_7941);
nor U12151 (N_12151,N_8791,N_9462);
or U12152 (N_12152,N_9780,N_8876);
nand U12153 (N_12153,N_9012,N_8686);
nor U12154 (N_12154,N_8862,N_8831);
and U12155 (N_12155,N_8313,N_9762);
or U12156 (N_12156,N_7839,N_8380);
or U12157 (N_12157,N_7908,N_9466);
nor U12158 (N_12158,N_8324,N_9688);
or U12159 (N_12159,N_7615,N_9738);
nand U12160 (N_12160,N_8799,N_9700);
or U12161 (N_12161,N_9373,N_8265);
or U12162 (N_12162,N_9860,N_7585);
and U12163 (N_12163,N_9234,N_9697);
or U12164 (N_12164,N_9517,N_7848);
and U12165 (N_12165,N_9977,N_9244);
or U12166 (N_12166,N_7508,N_8743);
nor U12167 (N_12167,N_9292,N_7672);
nand U12168 (N_12168,N_9091,N_8404);
or U12169 (N_12169,N_9815,N_9665);
nand U12170 (N_12170,N_7922,N_7946);
xnor U12171 (N_12171,N_9628,N_9761);
xor U12172 (N_12172,N_9362,N_9670);
nand U12173 (N_12173,N_7667,N_8384);
xnor U12174 (N_12174,N_8533,N_9517);
nand U12175 (N_12175,N_9439,N_8700);
or U12176 (N_12176,N_8408,N_7631);
or U12177 (N_12177,N_8464,N_9306);
nor U12178 (N_12178,N_8833,N_9137);
nand U12179 (N_12179,N_9309,N_7580);
nand U12180 (N_12180,N_9606,N_9915);
nor U12181 (N_12181,N_8391,N_9272);
nor U12182 (N_12182,N_9641,N_8871);
nor U12183 (N_12183,N_8520,N_8765);
nand U12184 (N_12184,N_7749,N_8752);
and U12185 (N_12185,N_7547,N_9868);
nand U12186 (N_12186,N_8324,N_9054);
xor U12187 (N_12187,N_9221,N_8402);
nor U12188 (N_12188,N_9746,N_9342);
nor U12189 (N_12189,N_9788,N_7725);
and U12190 (N_12190,N_8795,N_7715);
nand U12191 (N_12191,N_8579,N_7984);
nor U12192 (N_12192,N_8073,N_9658);
or U12193 (N_12193,N_8335,N_7529);
nor U12194 (N_12194,N_8343,N_8380);
nor U12195 (N_12195,N_8071,N_8815);
nand U12196 (N_12196,N_8122,N_9942);
nor U12197 (N_12197,N_9714,N_7603);
and U12198 (N_12198,N_7997,N_8067);
nor U12199 (N_12199,N_9961,N_8248);
or U12200 (N_12200,N_8374,N_7613);
or U12201 (N_12201,N_8980,N_9395);
xnor U12202 (N_12202,N_9486,N_8282);
nand U12203 (N_12203,N_9176,N_9073);
nor U12204 (N_12204,N_9878,N_7973);
nand U12205 (N_12205,N_9708,N_8180);
or U12206 (N_12206,N_8716,N_8051);
nor U12207 (N_12207,N_8647,N_7638);
xnor U12208 (N_12208,N_8968,N_8806);
and U12209 (N_12209,N_9010,N_8826);
and U12210 (N_12210,N_8365,N_9394);
nand U12211 (N_12211,N_9021,N_8801);
nor U12212 (N_12212,N_8799,N_8944);
xor U12213 (N_12213,N_7629,N_7781);
nand U12214 (N_12214,N_9895,N_8407);
or U12215 (N_12215,N_8740,N_8460);
or U12216 (N_12216,N_8093,N_8819);
and U12217 (N_12217,N_8224,N_9872);
or U12218 (N_12218,N_8130,N_9060);
xor U12219 (N_12219,N_8128,N_7853);
xnor U12220 (N_12220,N_8631,N_9829);
and U12221 (N_12221,N_9150,N_7779);
nand U12222 (N_12222,N_9279,N_9120);
nand U12223 (N_12223,N_8768,N_9644);
xor U12224 (N_12224,N_8390,N_9789);
and U12225 (N_12225,N_9351,N_8930);
and U12226 (N_12226,N_7750,N_8035);
nand U12227 (N_12227,N_7800,N_7859);
nor U12228 (N_12228,N_8415,N_8846);
or U12229 (N_12229,N_8812,N_8132);
or U12230 (N_12230,N_9619,N_7554);
or U12231 (N_12231,N_7714,N_9708);
xor U12232 (N_12232,N_8130,N_7664);
or U12233 (N_12233,N_8636,N_8962);
nor U12234 (N_12234,N_7772,N_8679);
xnor U12235 (N_12235,N_9971,N_8380);
xnor U12236 (N_12236,N_8257,N_7774);
or U12237 (N_12237,N_7521,N_7500);
nor U12238 (N_12238,N_8348,N_9661);
xnor U12239 (N_12239,N_9248,N_8380);
nand U12240 (N_12240,N_9309,N_8380);
or U12241 (N_12241,N_7783,N_8589);
xor U12242 (N_12242,N_8450,N_8541);
nand U12243 (N_12243,N_9932,N_8294);
or U12244 (N_12244,N_8562,N_9830);
nor U12245 (N_12245,N_8525,N_8585);
and U12246 (N_12246,N_9615,N_8995);
nand U12247 (N_12247,N_8616,N_9559);
nand U12248 (N_12248,N_8886,N_9657);
xor U12249 (N_12249,N_8340,N_7540);
and U12250 (N_12250,N_8159,N_9441);
and U12251 (N_12251,N_9115,N_7650);
and U12252 (N_12252,N_8353,N_8520);
and U12253 (N_12253,N_9680,N_9880);
and U12254 (N_12254,N_8331,N_9157);
nor U12255 (N_12255,N_9930,N_8405);
and U12256 (N_12256,N_9770,N_9217);
xor U12257 (N_12257,N_9176,N_8184);
nand U12258 (N_12258,N_8442,N_7958);
nor U12259 (N_12259,N_7556,N_7838);
nand U12260 (N_12260,N_9528,N_9099);
nor U12261 (N_12261,N_7688,N_7965);
nor U12262 (N_12262,N_9911,N_9305);
and U12263 (N_12263,N_9044,N_9707);
and U12264 (N_12264,N_7830,N_8568);
or U12265 (N_12265,N_7689,N_8799);
nor U12266 (N_12266,N_8136,N_9674);
xnor U12267 (N_12267,N_7520,N_9630);
xnor U12268 (N_12268,N_8936,N_8049);
nand U12269 (N_12269,N_9159,N_9028);
and U12270 (N_12270,N_7864,N_7533);
xor U12271 (N_12271,N_9014,N_9522);
or U12272 (N_12272,N_9475,N_8690);
or U12273 (N_12273,N_8111,N_9683);
xor U12274 (N_12274,N_7829,N_9412);
or U12275 (N_12275,N_8352,N_8119);
and U12276 (N_12276,N_9441,N_8648);
or U12277 (N_12277,N_8666,N_9764);
xnor U12278 (N_12278,N_8693,N_8905);
nand U12279 (N_12279,N_9411,N_9453);
nand U12280 (N_12280,N_7657,N_9863);
and U12281 (N_12281,N_8984,N_8332);
xor U12282 (N_12282,N_9192,N_8962);
nand U12283 (N_12283,N_9866,N_9798);
or U12284 (N_12284,N_7882,N_8960);
or U12285 (N_12285,N_9329,N_9021);
xnor U12286 (N_12286,N_7536,N_8573);
nor U12287 (N_12287,N_8924,N_9288);
and U12288 (N_12288,N_8434,N_9532);
or U12289 (N_12289,N_8765,N_7845);
and U12290 (N_12290,N_8101,N_8246);
and U12291 (N_12291,N_8309,N_9378);
nand U12292 (N_12292,N_9342,N_8400);
or U12293 (N_12293,N_7967,N_9415);
xor U12294 (N_12294,N_9836,N_9288);
xnor U12295 (N_12295,N_9885,N_9878);
or U12296 (N_12296,N_9517,N_9616);
or U12297 (N_12297,N_8234,N_9434);
xnor U12298 (N_12298,N_8734,N_9063);
xor U12299 (N_12299,N_7653,N_8372);
nor U12300 (N_12300,N_9961,N_7517);
or U12301 (N_12301,N_8088,N_8408);
nand U12302 (N_12302,N_8286,N_9940);
and U12303 (N_12303,N_7822,N_8324);
xnor U12304 (N_12304,N_8353,N_9385);
nand U12305 (N_12305,N_9826,N_7604);
nor U12306 (N_12306,N_9230,N_8962);
xor U12307 (N_12307,N_9587,N_8788);
nand U12308 (N_12308,N_7717,N_9852);
and U12309 (N_12309,N_9332,N_9847);
xnor U12310 (N_12310,N_7854,N_9184);
nor U12311 (N_12311,N_7996,N_7985);
and U12312 (N_12312,N_9087,N_9333);
or U12313 (N_12313,N_7942,N_8693);
nor U12314 (N_12314,N_8753,N_7695);
xnor U12315 (N_12315,N_9093,N_8725);
and U12316 (N_12316,N_9117,N_7962);
and U12317 (N_12317,N_9340,N_7808);
or U12318 (N_12318,N_7735,N_9890);
nor U12319 (N_12319,N_9177,N_8951);
nor U12320 (N_12320,N_8536,N_9747);
or U12321 (N_12321,N_8921,N_9320);
nand U12322 (N_12322,N_8193,N_7936);
nor U12323 (N_12323,N_7604,N_9440);
xnor U12324 (N_12324,N_7667,N_8589);
xnor U12325 (N_12325,N_8941,N_8592);
and U12326 (N_12326,N_8401,N_8313);
nand U12327 (N_12327,N_9342,N_8513);
nor U12328 (N_12328,N_9876,N_9442);
xor U12329 (N_12329,N_8159,N_8883);
or U12330 (N_12330,N_7827,N_8199);
xor U12331 (N_12331,N_8955,N_8164);
and U12332 (N_12332,N_9808,N_8180);
or U12333 (N_12333,N_9383,N_8294);
nand U12334 (N_12334,N_9327,N_8684);
and U12335 (N_12335,N_7882,N_8285);
xnor U12336 (N_12336,N_8064,N_8051);
xor U12337 (N_12337,N_9884,N_8451);
xnor U12338 (N_12338,N_8125,N_8364);
xor U12339 (N_12339,N_8169,N_7699);
nand U12340 (N_12340,N_9212,N_9122);
nand U12341 (N_12341,N_8145,N_9782);
nor U12342 (N_12342,N_7690,N_9561);
nand U12343 (N_12343,N_7513,N_7563);
and U12344 (N_12344,N_9407,N_8553);
nor U12345 (N_12345,N_8437,N_9756);
and U12346 (N_12346,N_9439,N_8488);
xor U12347 (N_12347,N_8016,N_9411);
or U12348 (N_12348,N_9459,N_7754);
xnor U12349 (N_12349,N_9237,N_7880);
nand U12350 (N_12350,N_9532,N_7559);
xor U12351 (N_12351,N_9052,N_9565);
xnor U12352 (N_12352,N_9443,N_8318);
or U12353 (N_12353,N_8090,N_8752);
or U12354 (N_12354,N_8525,N_7729);
or U12355 (N_12355,N_8794,N_8491);
nand U12356 (N_12356,N_9496,N_8170);
nor U12357 (N_12357,N_9508,N_9564);
xor U12358 (N_12358,N_9350,N_9611);
nand U12359 (N_12359,N_9671,N_9984);
nor U12360 (N_12360,N_7823,N_9055);
nand U12361 (N_12361,N_9092,N_9246);
nand U12362 (N_12362,N_8217,N_8934);
or U12363 (N_12363,N_9674,N_9058);
xnor U12364 (N_12364,N_8516,N_9056);
nand U12365 (N_12365,N_8574,N_9636);
nand U12366 (N_12366,N_8965,N_8815);
nor U12367 (N_12367,N_9964,N_8457);
nor U12368 (N_12368,N_7706,N_8959);
nand U12369 (N_12369,N_8331,N_9307);
nor U12370 (N_12370,N_8523,N_9021);
nand U12371 (N_12371,N_7753,N_7918);
nor U12372 (N_12372,N_8050,N_9959);
nand U12373 (N_12373,N_9588,N_8076);
and U12374 (N_12374,N_8855,N_8674);
or U12375 (N_12375,N_8885,N_9261);
and U12376 (N_12376,N_8232,N_9202);
nor U12377 (N_12377,N_8264,N_8358);
and U12378 (N_12378,N_7546,N_8927);
nand U12379 (N_12379,N_8826,N_9690);
or U12380 (N_12380,N_8965,N_9940);
and U12381 (N_12381,N_8523,N_8929);
nand U12382 (N_12382,N_8479,N_9248);
nor U12383 (N_12383,N_9735,N_7518);
xnor U12384 (N_12384,N_8659,N_9741);
nor U12385 (N_12385,N_9872,N_8907);
and U12386 (N_12386,N_9361,N_9669);
nand U12387 (N_12387,N_8803,N_8628);
nand U12388 (N_12388,N_7826,N_8701);
nor U12389 (N_12389,N_8492,N_9278);
and U12390 (N_12390,N_7988,N_8542);
or U12391 (N_12391,N_9950,N_7770);
or U12392 (N_12392,N_9426,N_8096);
xnor U12393 (N_12393,N_8554,N_8720);
and U12394 (N_12394,N_8046,N_7979);
xnor U12395 (N_12395,N_8442,N_8154);
nor U12396 (N_12396,N_9033,N_7865);
and U12397 (N_12397,N_8603,N_7568);
nor U12398 (N_12398,N_8562,N_8673);
and U12399 (N_12399,N_7680,N_9389);
nor U12400 (N_12400,N_9057,N_7610);
nand U12401 (N_12401,N_9268,N_8749);
or U12402 (N_12402,N_9869,N_9052);
nor U12403 (N_12403,N_7871,N_9046);
nand U12404 (N_12404,N_7568,N_9244);
and U12405 (N_12405,N_8282,N_8610);
nor U12406 (N_12406,N_9619,N_7691);
nor U12407 (N_12407,N_8907,N_8841);
and U12408 (N_12408,N_9067,N_9238);
nor U12409 (N_12409,N_9359,N_9294);
or U12410 (N_12410,N_9600,N_9943);
and U12411 (N_12411,N_8658,N_8893);
nor U12412 (N_12412,N_8845,N_9546);
and U12413 (N_12413,N_7967,N_8380);
nor U12414 (N_12414,N_9469,N_8839);
xnor U12415 (N_12415,N_9393,N_8501);
or U12416 (N_12416,N_9873,N_8792);
and U12417 (N_12417,N_8805,N_7637);
xnor U12418 (N_12418,N_9501,N_8637);
nand U12419 (N_12419,N_8497,N_8021);
nor U12420 (N_12420,N_9048,N_9442);
nand U12421 (N_12421,N_7879,N_9636);
nor U12422 (N_12422,N_7543,N_9105);
nor U12423 (N_12423,N_8469,N_9595);
or U12424 (N_12424,N_8599,N_9085);
nand U12425 (N_12425,N_9483,N_7836);
or U12426 (N_12426,N_8222,N_8585);
or U12427 (N_12427,N_8900,N_8424);
or U12428 (N_12428,N_8138,N_8598);
nor U12429 (N_12429,N_9090,N_7681);
nor U12430 (N_12430,N_9434,N_8987);
nand U12431 (N_12431,N_9604,N_9385);
xor U12432 (N_12432,N_7877,N_9702);
nand U12433 (N_12433,N_7978,N_7789);
and U12434 (N_12434,N_8805,N_8677);
nand U12435 (N_12435,N_7933,N_9106);
and U12436 (N_12436,N_8779,N_9161);
and U12437 (N_12437,N_8425,N_9324);
or U12438 (N_12438,N_7647,N_7940);
or U12439 (N_12439,N_9090,N_8941);
nor U12440 (N_12440,N_8662,N_7839);
or U12441 (N_12441,N_8001,N_9047);
xor U12442 (N_12442,N_8554,N_7537);
or U12443 (N_12443,N_9954,N_8605);
nor U12444 (N_12444,N_7990,N_9253);
nand U12445 (N_12445,N_9477,N_9281);
nand U12446 (N_12446,N_8412,N_9793);
and U12447 (N_12447,N_9768,N_9951);
and U12448 (N_12448,N_8446,N_9048);
and U12449 (N_12449,N_9372,N_8984);
nand U12450 (N_12450,N_8962,N_7876);
xor U12451 (N_12451,N_9716,N_9317);
and U12452 (N_12452,N_9077,N_9275);
and U12453 (N_12453,N_9949,N_7566);
nand U12454 (N_12454,N_8911,N_8858);
nor U12455 (N_12455,N_9040,N_7899);
or U12456 (N_12456,N_9602,N_7509);
and U12457 (N_12457,N_8817,N_8130);
and U12458 (N_12458,N_7579,N_9652);
nand U12459 (N_12459,N_8161,N_9935);
xor U12460 (N_12460,N_9513,N_9916);
nand U12461 (N_12461,N_7848,N_8461);
and U12462 (N_12462,N_8463,N_9061);
nor U12463 (N_12463,N_8080,N_9068);
xnor U12464 (N_12464,N_8113,N_8349);
nor U12465 (N_12465,N_9164,N_8186);
or U12466 (N_12466,N_8133,N_9844);
xnor U12467 (N_12467,N_9106,N_8406);
or U12468 (N_12468,N_8371,N_9289);
xnor U12469 (N_12469,N_7999,N_8645);
nor U12470 (N_12470,N_8004,N_9946);
nand U12471 (N_12471,N_7770,N_8475);
nand U12472 (N_12472,N_8266,N_9348);
and U12473 (N_12473,N_9292,N_9878);
xor U12474 (N_12474,N_8673,N_9211);
or U12475 (N_12475,N_9732,N_8344);
nand U12476 (N_12476,N_9545,N_8243);
or U12477 (N_12477,N_7718,N_8326);
nor U12478 (N_12478,N_7922,N_8929);
or U12479 (N_12479,N_7638,N_8769);
and U12480 (N_12480,N_8632,N_8599);
or U12481 (N_12481,N_9922,N_8326);
or U12482 (N_12482,N_7855,N_8292);
and U12483 (N_12483,N_7863,N_8297);
nor U12484 (N_12484,N_8008,N_9912);
nand U12485 (N_12485,N_7890,N_7885);
nor U12486 (N_12486,N_7559,N_8604);
nor U12487 (N_12487,N_9199,N_7882);
and U12488 (N_12488,N_9300,N_8050);
nor U12489 (N_12489,N_7748,N_9496);
and U12490 (N_12490,N_7965,N_9400);
or U12491 (N_12491,N_9046,N_9881);
or U12492 (N_12492,N_7670,N_9389);
and U12493 (N_12493,N_7630,N_8199);
and U12494 (N_12494,N_7923,N_8730);
and U12495 (N_12495,N_7823,N_9307);
nor U12496 (N_12496,N_9975,N_8891);
xor U12497 (N_12497,N_9734,N_7724);
xnor U12498 (N_12498,N_8280,N_9818);
nor U12499 (N_12499,N_8179,N_7587);
nor U12500 (N_12500,N_10006,N_11006);
xor U12501 (N_12501,N_10385,N_11928);
and U12502 (N_12502,N_11197,N_12153);
nor U12503 (N_12503,N_10184,N_12069);
nand U12504 (N_12504,N_11272,N_11316);
nor U12505 (N_12505,N_12093,N_11719);
and U12506 (N_12506,N_11830,N_10279);
nor U12507 (N_12507,N_11969,N_10232);
and U12508 (N_12508,N_11948,N_10679);
xnor U12509 (N_12509,N_11825,N_11979);
and U12510 (N_12510,N_11766,N_10701);
nand U12511 (N_12511,N_12223,N_11417);
nor U12512 (N_12512,N_10377,N_10863);
nor U12513 (N_12513,N_11765,N_11521);
nand U12514 (N_12514,N_11322,N_11929);
nand U12515 (N_12515,N_12475,N_11294);
or U12516 (N_12516,N_11756,N_10563);
nand U12517 (N_12517,N_11542,N_10722);
xnor U12518 (N_12518,N_10606,N_10816);
nand U12519 (N_12519,N_10354,N_10877);
nor U12520 (N_12520,N_10486,N_12192);
xnor U12521 (N_12521,N_11736,N_11471);
nand U12522 (N_12522,N_11022,N_12406);
and U12523 (N_12523,N_12315,N_12477);
xor U12524 (N_12524,N_10352,N_11643);
xor U12525 (N_12525,N_10144,N_10161);
xor U12526 (N_12526,N_10862,N_12458);
nor U12527 (N_12527,N_11485,N_12374);
nor U12528 (N_12528,N_12484,N_11448);
xnor U12529 (N_12529,N_11382,N_10454);
xor U12530 (N_12530,N_11386,N_11149);
nor U12531 (N_12531,N_10704,N_11604);
or U12532 (N_12532,N_10527,N_10441);
xor U12533 (N_12533,N_11293,N_12098);
nor U12534 (N_12534,N_11458,N_11051);
or U12535 (N_12535,N_10294,N_10258);
nand U12536 (N_12536,N_12037,N_12221);
or U12537 (N_12537,N_10605,N_12411);
or U12538 (N_12538,N_11469,N_12397);
nand U12539 (N_12539,N_10781,N_11374);
xnor U12540 (N_12540,N_11039,N_10149);
and U12541 (N_12541,N_11452,N_10236);
nor U12542 (N_12542,N_10005,N_12030);
and U12543 (N_12543,N_10371,N_12470);
or U12544 (N_12544,N_10769,N_10539);
or U12545 (N_12545,N_11633,N_10755);
xor U12546 (N_12546,N_11373,N_11733);
nand U12547 (N_12547,N_11170,N_12033);
nand U12548 (N_12548,N_12287,N_12201);
xor U12549 (N_12549,N_11539,N_11284);
xnor U12550 (N_12550,N_10423,N_10641);
nand U12551 (N_12551,N_10492,N_10518);
and U12552 (N_12552,N_10947,N_12330);
or U12553 (N_12553,N_10452,N_10218);
xnor U12554 (N_12554,N_12480,N_11744);
xnor U12555 (N_12555,N_12266,N_10920);
nor U12556 (N_12556,N_10474,N_10455);
or U12557 (N_12557,N_10783,N_11481);
and U12558 (N_12558,N_11913,N_10439);
and U12559 (N_12559,N_11487,N_10536);
and U12560 (N_12560,N_12068,N_10030);
or U12561 (N_12561,N_11531,N_11171);
nand U12562 (N_12562,N_10938,N_10712);
and U12563 (N_12563,N_11876,N_10225);
nand U12564 (N_12564,N_10136,N_11501);
nand U12565 (N_12565,N_12214,N_12301);
nor U12566 (N_12566,N_11924,N_10212);
or U12567 (N_12567,N_11918,N_11499);
nor U12568 (N_12568,N_10021,N_12238);
or U12569 (N_12569,N_10747,N_12324);
or U12570 (N_12570,N_10569,N_12229);
nand U12571 (N_12571,N_12228,N_12151);
xnor U12572 (N_12572,N_11721,N_10885);
xnor U12573 (N_12573,N_10264,N_11617);
or U12574 (N_12574,N_11627,N_11999);
xor U12575 (N_12575,N_11800,N_11219);
or U12576 (N_12576,N_11804,N_10159);
or U12577 (N_12577,N_11698,N_11465);
xor U12578 (N_12578,N_10626,N_10427);
and U12579 (N_12579,N_10115,N_11693);
nand U12580 (N_12580,N_12144,N_10754);
nand U12581 (N_12581,N_10231,N_10241);
nor U12582 (N_12582,N_10465,N_11921);
or U12583 (N_12583,N_10538,N_10117);
nor U12584 (N_12584,N_10100,N_10227);
nor U12585 (N_12585,N_12158,N_10449);
xnor U12586 (N_12586,N_12461,N_11433);
nor U12587 (N_12587,N_10523,N_12465);
or U12588 (N_12588,N_12118,N_10824);
nor U12589 (N_12589,N_12125,N_11413);
xor U12590 (N_12590,N_12468,N_12169);
and U12591 (N_12591,N_10571,N_10095);
nor U12592 (N_12592,N_10444,N_11184);
and U12593 (N_12593,N_11728,N_11982);
nand U12594 (N_12594,N_12076,N_10806);
and U12595 (N_12595,N_11562,N_12402);
and U12596 (N_12596,N_11420,N_11391);
or U12597 (N_12597,N_10811,N_12172);
nand U12598 (N_12598,N_12494,N_10965);
nand U12599 (N_12599,N_10414,N_11097);
and U12600 (N_12600,N_11988,N_11571);
nor U12601 (N_12601,N_12224,N_11343);
xnor U12602 (N_12602,N_10167,N_11259);
xor U12603 (N_12603,N_10696,N_10316);
nor U12604 (N_12604,N_12352,N_11887);
xor U12605 (N_12605,N_12104,N_12450);
xor U12606 (N_12606,N_11215,N_11598);
nor U12607 (N_12607,N_12060,N_11187);
or U12608 (N_12608,N_12323,N_11032);
nor U12609 (N_12609,N_11176,N_10731);
and U12610 (N_12610,N_11218,N_12120);
and U12611 (N_12611,N_10209,N_11372);
xnor U12612 (N_12612,N_10660,N_10768);
nand U12613 (N_12613,N_10510,N_11737);
nand U12614 (N_12614,N_11415,N_11667);
or U12615 (N_12615,N_10409,N_11300);
nand U12616 (N_12616,N_10949,N_10586);
nor U12617 (N_12617,N_10958,N_10201);
or U12618 (N_12618,N_11962,N_10173);
nand U12619 (N_12619,N_11730,N_12176);
nand U12620 (N_12620,N_12325,N_11466);
nor U12621 (N_12621,N_11623,N_10331);
xnor U12622 (N_12622,N_11624,N_10237);
nand U12623 (N_12623,N_11971,N_10633);
xor U12624 (N_12624,N_10598,N_11726);
xor U12625 (N_12625,N_12463,N_11524);
or U12626 (N_12626,N_11861,N_11011);
or U12627 (N_12627,N_12380,N_12211);
nor U12628 (N_12628,N_10139,N_12428);
or U12629 (N_12629,N_11870,N_10883);
xnor U12630 (N_12630,N_12369,N_11354);
nand U12631 (N_12631,N_11670,N_11673);
nor U12632 (N_12632,N_10673,N_11664);
and U12633 (N_12633,N_11050,N_11684);
and U12634 (N_12634,N_10813,N_10695);
or U12635 (N_12635,N_10993,N_11102);
xnor U12636 (N_12636,N_10562,N_11828);
or U12637 (N_12637,N_12002,N_10537);
nor U12638 (N_12638,N_11334,N_11541);
xor U12639 (N_12639,N_11826,N_12167);
and U12640 (N_12640,N_11062,N_11056);
nor U12641 (N_12641,N_10891,N_11656);
and U12642 (N_12642,N_10016,N_10265);
nor U12643 (N_12643,N_12081,N_12162);
xor U12644 (N_12644,N_12225,N_11360);
or U12645 (N_12645,N_12471,N_11194);
xor U12646 (N_12646,N_11101,N_11907);
nand U12647 (N_12647,N_10573,N_11427);
nand U12648 (N_12648,N_11764,N_11209);
nand U12649 (N_12649,N_10150,N_12300);
nor U12650 (N_12650,N_11915,N_12283);
nor U12651 (N_12651,N_12353,N_10437);
nand U12652 (N_12652,N_10203,N_10109);
and U12653 (N_12653,N_12044,N_10770);
or U12654 (N_12654,N_10828,N_12263);
nand U12655 (N_12655,N_11064,N_11709);
xor U12656 (N_12656,N_10574,N_10336);
nor U12657 (N_12657,N_11088,N_11949);
nor U12658 (N_12658,N_12043,N_12491);
or U12659 (N_12659,N_10047,N_10353);
nor U12660 (N_12660,N_11424,N_11973);
or U12661 (N_12661,N_12213,N_10359);
and U12662 (N_12662,N_11076,N_11271);
nor U12663 (N_12663,N_10752,N_11147);
nand U12664 (N_12664,N_10915,N_11526);
nor U12665 (N_12665,N_11137,N_11378);
xnor U12666 (N_12666,N_10322,N_12483);
and U12667 (N_12667,N_11871,N_11500);
or U12668 (N_12668,N_12137,N_10189);
or U12669 (N_12669,N_11642,N_11063);
nor U12670 (N_12670,N_11312,N_12115);
or U12671 (N_12671,N_11394,N_12009);
nand U12672 (N_12672,N_10330,N_12251);
or U12673 (N_12673,N_11952,N_11460);
or U12674 (N_12674,N_10000,N_10587);
or U12675 (N_12675,N_12050,N_12379);
or U12676 (N_12676,N_10960,N_10317);
nand U12677 (N_12677,N_10007,N_11860);
and U12678 (N_12678,N_12121,N_11114);
or U12679 (N_12679,N_10106,N_11156);
and U12680 (N_12680,N_10499,N_11486);
and U12681 (N_12681,N_10799,N_10224);
xnor U12682 (N_12682,N_10299,N_12420);
or U12683 (N_12683,N_10276,N_10420);
xor U12684 (N_12684,N_10089,N_12419);
or U12685 (N_12685,N_11936,N_10325);
xor U12686 (N_12686,N_11290,N_11798);
or U12687 (N_12687,N_12499,N_11514);
xor U12688 (N_12688,N_10989,N_10063);
nor U12689 (N_12689,N_11115,N_11277);
xnor U12690 (N_12690,N_12070,N_11805);
nand U12691 (N_12691,N_10200,N_10478);
nand U12692 (N_12692,N_11264,N_11318);
xnor U12693 (N_12693,N_10942,N_10341);
xnor U12694 (N_12694,N_10533,N_10559);
or U12695 (N_12695,N_10055,N_11474);
or U12696 (N_12696,N_10254,N_11456);
xor U12697 (N_12697,N_12026,N_12331);
nand U12698 (N_12698,N_10540,N_11945);
xor U12699 (N_12699,N_10829,N_11069);
and U12700 (N_12700,N_10097,N_11302);
nor U12701 (N_12701,N_11037,N_11462);
and U12702 (N_12702,N_10937,N_11793);
or U12703 (N_12703,N_10708,N_10982);
nand U12704 (N_12704,N_11490,N_12448);
nor U12705 (N_12705,N_12286,N_11132);
nor U12706 (N_12706,N_12234,N_12431);
and U12707 (N_12707,N_11757,N_11204);
or U12708 (N_12708,N_11074,N_11620);
and U12709 (N_12709,N_11365,N_12047);
and U12710 (N_12710,N_10066,N_10335);
xnor U12711 (N_12711,N_11968,N_12433);
and U12712 (N_12712,N_12036,N_11152);
or U12713 (N_12713,N_10373,N_12342);
xnor U12714 (N_12714,N_11889,N_10864);
and U12715 (N_12715,N_11375,N_10168);
xor U12716 (N_12716,N_10363,N_11845);
nand U12717 (N_12717,N_11364,N_10865);
nor U12718 (N_12718,N_10567,N_11496);
xnor U12719 (N_12719,N_11168,N_10155);
xnor U12720 (N_12720,N_10820,N_12080);
or U12721 (N_12721,N_12393,N_12421);
or U12722 (N_12722,N_12000,N_11618);
nor U12723 (N_12723,N_12216,N_11282);
nor U12724 (N_12724,N_11724,N_12001);
nand U12725 (N_12725,N_10645,N_10302);
xor U12726 (N_12726,N_12179,N_11966);
and U12727 (N_12727,N_11153,N_11538);
xor U12728 (N_12728,N_10070,N_11444);
xor U12729 (N_12729,N_11641,N_12049);
nor U12730 (N_12730,N_12261,N_12347);
or U12731 (N_12731,N_10931,N_11864);
nand U12732 (N_12732,N_10910,N_10718);
nand U12733 (N_12733,N_10018,N_12103);
and U12734 (N_12734,N_10978,N_11634);
xor U12735 (N_12735,N_10493,N_11105);
and U12736 (N_12736,N_11447,N_10187);
nand U12737 (N_12737,N_10471,N_11042);
and U12738 (N_12738,N_10566,N_11067);
or U12739 (N_12739,N_10088,N_10948);
and U12740 (N_12740,N_12159,N_10923);
nor U12741 (N_12741,N_10514,N_10164);
nand U12742 (N_12742,N_11543,N_12269);
or U12743 (N_12743,N_10152,N_11802);
and U12744 (N_12744,N_11650,N_12016);
nor U12745 (N_12745,N_10779,N_10797);
nand U12746 (N_12746,N_11100,N_11640);
or U12747 (N_12747,N_11348,N_10616);
and U12748 (N_12748,N_10810,N_12059);
xnor U12749 (N_12749,N_11278,N_12271);
or U12750 (N_12750,N_10108,N_11545);
or U12751 (N_12751,N_11236,N_10318);
nand U12752 (N_12752,N_11903,N_12446);
nand U12753 (N_12753,N_12004,N_11154);
and U12754 (N_12754,N_11732,N_12123);
or U12755 (N_12755,N_11108,N_11925);
nor U12756 (N_12756,N_11905,N_11705);
or U12757 (N_12757,N_10214,N_11546);
nand U12758 (N_12758,N_10308,N_12456);
nor U12759 (N_12759,N_10705,N_10368);
and U12760 (N_12760,N_11116,N_12147);
xor U12761 (N_12761,N_11279,N_10686);
xor U12762 (N_12762,N_12436,N_11252);
nand U12763 (N_12763,N_11609,N_11722);
nor U12764 (N_12764,N_10422,N_11307);
nand U12765 (N_12765,N_11159,N_11972);
nand U12766 (N_12766,N_10242,N_12321);
xor U12767 (N_12767,N_10814,N_12349);
nor U12768 (N_12768,N_10303,N_12156);
xnor U12769 (N_12769,N_11916,N_10488);
and U12770 (N_12770,N_11926,N_10991);
xnor U12771 (N_12771,N_10288,N_11580);
nand U12772 (N_12772,N_10328,N_10290);
nor U12773 (N_12773,N_11213,N_10547);
nand U12774 (N_12774,N_11563,N_12275);
and U12775 (N_12775,N_11525,N_11495);
nor U12776 (N_12776,N_11164,N_10825);
nor U12777 (N_12777,N_11893,N_11119);
nor U12778 (N_12778,N_11031,N_10413);
and U12779 (N_12779,N_12074,N_11175);
or U12780 (N_12780,N_11603,N_10116);
nor U12781 (N_12781,N_11321,N_10740);
xnor U12782 (N_12782,N_11553,N_11414);
nor U12783 (N_12783,N_11345,N_12164);
and U12784 (N_12784,N_11216,N_10376);
nor U12785 (N_12785,N_11748,N_12295);
nor U12786 (N_12786,N_11699,N_12140);
nand U12787 (N_12787,N_11529,N_12362);
xor U12788 (N_12788,N_11827,N_10542);
or U12789 (N_12789,N_11353,N_11058);
nor U12790 (N_12790,N_12363,N_10917);
xor U12791 (N_12791,N_12392,N_12048);
nor U12792 (N_12792,N_10529,N_10979);
nand U12793 (N_12793,N_12398,N_12240);
xnor U12794 (N_12794,N_11549,N_11970);
and U12795 (N_12795,N_10699,N_10798);
nor U12796 (N_12796,N_12054,N_12046);
xnor U12797 (N_12797,N_10012,N_12438);
xor U12798 (N_12798,N_12249,N_12385);
or U12799 (N_12799,N_12086,N_11686);
or U12800 (N_12800,N_10326,N_11053);
xor U12801 (N_12801,N_10138,N_11400);
nor U12802 (N_12802,N_10516,N_11397);
nand U12803 (N_12803,N_10585,N_12195);
nand U12804 (N_12804,N_10684,N_12417);
xor U12805 (N_12805,N_11513,N_11834);
xor U12806 (N_12806,N_12360,N_11081);
or U12807 (N_12807,N_10871,N_10301);
or U12808 (N_12808,N_11082,N_10064);
nor U12809 (N_12809,N_10190,N_11850);
xnor U12810 (N_12810,N_11872,N_11778);
or U12811 (N_12811,N_12361,N_10596);
xor U12812 (N_12812,N_11644,N_10506);
nor U12813 (N_12813,N_10837,N_11434);
nand U12814 (N_12814,N_11848,N_10132);
xor U12815 (N_12815,N_12305,N_11174);
or U12816 (N_12816,N_10153,N_10672);
nand U12817 (N_12817,N_10742,N_11977);
or U12818 (N_12818,N_11878,N_11577);
or U12819 (N_12819,N_10804,N_11773);
or U12820 (N_12820,N_10323,N_11946);
and U12821 (N_12821,N_10940,N_11480);
nor U12822 (N_12822,N_11654,N_12052);
xor U12823 (N_12823,N_11810,N_10846);
nand U12824 (N_12824,N_12449,N_12467);
xnor U12825 (N_12825,N_10994,N_11616);
or U12826 (N_12826,N_10916,N_11281);
or U12827 (N_12827,N_10997,N_12018);
and U12828 (N_12828,N_12114,N_12190);
xnor U12829 (N_12829,N_11412,N_11750);
nand U12830 (N_12830,N_10381,N_11422);
or U12831 (N_12831,N_10784,N_11986);
nand U12832 (N_12832,N_11505,N_12490);
or U12833 (N_12833,N_11983,N_11379);
xnor U12834 (N_12834,N_11298,N_11574);
nor U12835 (N_12835,N_10908,N_12241);
or U12836 (N_12836,N_10685,N_11919);
or U12837 (N_12837,N_10522,N_11844);
nand U12838 (N_12838,N_11430,N_11110);
nand U12839 (N_12839,N_10496,N_10895);
xnor U12840 (N_12840,N_10584,N_10142);
and U12841 (N_12841,N_11285,N_10032);
nand U12842 (N_12842,N_11877,N_10850);
nor U12843 (N_12843,N_10295,N_12196);
or U12844 (N_12844,N_10560,N_10428);
xnor U12845 (N_12845,N_12028,N_10807);
or U12846 (N_12846,N_10001,N_12034);
or U12847 (N_12847,N_11221,N_12337);
and U12848 (N_12848,N_10525,N_10186);
nand U12849 (N_12849,N_10347,N_10904);
nand U12850 (N_12850,N_12375,N_11262);
nand U12851 (N_12851,N_11036,N_11183);
and U12852 (N_12852,N_10096,N_12005);
nand U12853 (N_12853,N_11342,N_12365);
and U12854 (N_12854,N_10172,N_11852);
nand U12855 (N_12855,N_10860,N_10886);
nand U12856 (N_12856,N_11685,N_10374);
nor U12857 (N_12857,N_12107,N_10730);
nand U12858 (N_12858,N_11244,N_11955);
and U12859 (N_12859,N_11791,N_10872);
xor U12860 (N_12860,N_11350,N_10221);
and U12861 (N_12861,N_11729,N_10126);
nor U12862 (N_12862,N_10130,N_11276);
xnor U12863 (N_12863,N_11033,N_10051);
nor U12864 (N_12864,N_11357,N_10213);
and U12865 (N_12865,N_10791,N_11932);
and U12866 (N_12866,N_10834,N_10313);
or U12867 (N_12867,N_11167,N_12388);
xor U12868 (N_12868,N_11220,N_10456);
nor U12869 (N_12869,N_12035,N_10630);
xor U12870 (N_12870,N_10086,N_10462);
nand U12871 (N_12871,N_12441,N_11269);
or U12872 (N_12872,N_11718,N_10059);
or U12873 (N_12873,N_11048,N_11193);
or U12874 (N_12874,N_10776,N_12181);
xor U12875 (N_12875,N_10995,N_10416);
and U12876 (N_12876,N_10083,N_10244);
or U12877 (N_12877,N_10102,N_11573);
xnor U12878 (N_12878,N_10678,N_10889);
and U12879 (N_12879,N_10350,N_11532);
nor U12880 (N_12880,N_11061,N_11892);
nor U12881 (N_12881,N_12495,N_12313);
nand U12882 (N_12882,N_11984,N_10654);
xor U12883 (N_12883,N_12279,N_11157);
nand U12884 (N_12884,N_12403,N_12289);
nand U12885 (N_12885,N_10447,N_11291);
and U12886 (N_12886,N_10892,N_11837);
nand U12887 (N_12887,N_10440,N_11613);
and U12888 (N_12888,N_12227,N_11941);
or U12889 (N_12889,N_12186,N_12101);
or U12890 (N_12890,N_10838,N_10078);
nor U12891 (N_12891,N_10387,N_11403);
nor U12892 (N_12892,N_11833,N_10952);
nand U12893 (N_12893,N_11470,N_10469);
or U12894 (N_12894,N_12299,N_12226);
nand U12895 (N_12895,N_11239,N_11383);
xnor U12896 (N_12896,N_11743,N_10135);
and U12897 (N_12897,N_11985,N_10287);
or U12898 (N_12898,N_10763,N_12237);
nand U12899 (N_12899,N_12307,N_11619);
nand U12900 (N_12900,N_11188,N_10031);
nand U12901 (N_12901,N_11572,N_10998);
xnor U12902 (N_12902,N_11150,N_11669);
xnor U12903 (N_12903,N_11402,N_11856);
nand U12904 (N_12904,N_11146,N_12222);
xor U12905 (N_12905,N_11071,N_10104);
xnor U12906 (N_12906,N_11681,N_11326);
nor U12907 (N_12907,N_11720,N_11831);
nor U12908 (N_12908,N_11865,N_10194);
nor U12909 (N_12909,N_10852,N_11052);
nor U12910 (N_12910,N_10248,N_10670);
nand U12911 (N_12911,N_11059,N_10162);
xor U12912 (N_12912,N_11843,N_10651);
xnor U12913 (N_12913,N_11004,N_12145);
nor U12914 (N_12914,N_11077,N_10577);
and U12915 (N_12915,N_11746,N_11672);
xnor U12916 (N_12916,N_10022,N_10709);
or U12917 (N_12917,N_12454,N_11320);
and U12918 (N_12918,N_11958,N_11129);
or U12919 (N_12919,N_11832,N_10627);
nand U12920 (N_12920,N_10946,N_10913);
nand U12921 (N_12921,N_11938,N_11161);
or U12922 (N_12922,N_11410,N_11803);
nor U12923 (N_12923,N_11185,N_10737);
nor U12924 (N_12924,N_11993,N_10391);
and U12925 (N_12925,N_10592,N_10234);
nand U12926 (N_12926,N_11884,N_11854);
xor U12927 (N_12927,N_12487,N_10817);
and U12928 (N_12928,N_11712,N_12110);
and U12929 (N_12929,N_10226,N_11859);
nor U12930 (N_12930,N_11628,N_11073);
xnor U12931 (N_12931,N_10042,N_11464);
xor U12932 (N_12932,N_10683,N_10690);
and U12933 (N_12933,N_10480,N_10056);
xor U12934 (N_12934,N_10246,N_12314);
nand U12935 (N_12935,N_11506,N_10068);
nor U12936 (N_12936,N_12303,N_12130);
xor U12937 (N_12937,N_10069,N_10773);
or U12938 (N_12938,N_12090,N_11917);
xnor U12939 (N_12939,N_11027,N_10141);
nor U12940 (N_12940,N_10694,N_11260);
and U12941 (N_12941,N_11639,N_11547);
nand U12942 (N_12942,N_10169,N_11190);
nor U12943 (N_12943,N_11047,N_11551);
nor U12944 (N_12944,N_12232,N_10457);
nand U12945 (N_12945,N_11449,N_11367);
and U12946 (N_12946,N_12492,N_12294);
nand U12947 (N_12947,N_12407,N_10581);
nor U12948 (N_12948,N_12209,N_12170);
and U12949 (N_12949,N_10981,N_11621);
xnor U12950 (N_12950,N_12011,N_10366);
or U12951 (N_12951,N_11177,N_12102);
nor U12952 (N_12952,N_11679,N_10125);
nand U12953 (N_12953,N_11333,N_11661);
and U12954 (N_12954,N_11181,N_10235);
nand U12955 (N_12955,N_10517,N_11675);
or U12956 (N_12956,N_10733,N_10604);
and U12957 (N_12957,N_11266,N_10925);
or U12958 (N_12958,N_11223,N_11337);
or U12959 (N_12959,N_11610,N_11035);
or U12960 (N_12960,N_11034,N_10667);
xor U12961 (N_12961,N_11891,N_11787);
nand U12962 (N_12962,N_11384,N_11411);
nor U12963 (N_12963,N_11245,N_11070);
nand U12964 (N_12964,N_11346,N_11760);
nor U12965 (N_12965,N_11380,N_12377);
xor U12966 (N_12966,N_11901,N_12437);
nand U12967 (N_12967,N_12119,N_11120);
nor U12968 (N_12968,N_12168,N_10549);
xor U12969 (N_12969,N_10782,N_11991);
xnor U12970 (N_12970,N_11680,N_12188);
nand U12971 (N_12971,N_10393,N_11428);
xnor U12972 (N_12972,N_11358,N_12346);
or U12973 (N_12973,N_11151,N_11607);
nor U12974 (N_12974,N_11920,N_11090);
or U12975 (N_12975,N_10570,N_11782);
xor U12976 (N_12976,N_12466,N_10611);
nand U12977 (N_12977,N_10181,N_11601);
nand U12978 (N_12978,N_12252,N_10340);
nand U12979 (N_12979,N_12094,N_11040);
nor U12980 (N_12980,N_12218,N_12354);
nor U12981 (N_12981,N_11359,N_10866);
and U12982 (N_12982,N_11301,N_11683);
or U12983 (N_12983,N_11224,N_12173);
and U12984 (N_12984,N_10901,N_10970);
or U12985 (N_12985,N_11015,N_10687);
xnor U12986 (N_12986,N_11385,N_11296);
and U12987 (N_12987,N_12285,N_11468);
or U12988 (N_12988,N_11752,N_10650);
nor U12989 (N_12989,N_12150,N_10835);
or U12990 (N_12990,N_11688,N_10035);
nand U12991 (N_12991,N_11657,N_10725);
or U12992 (N_12992,N_10726,N_10927);
nand U12993 (N_12993,N_11611,N_11173);
nand U12994 (N_12994,N_12200,N_11297);
nor U12995 (N_12995,N_10888,N_11370);
nand U12996 (N_12996,N_11786,N_10481);
nor U12997 (N_12997,N_10268,N_10924);
and U12998 (N_12998,N_10874,N_10384);
and U12999 (N_12999,N_10476,N_12488);
xnor U13000 (N_13000,N_10634,N_11519);
or U13001 (N_13001,N_11099,N_10280);
nor U13002 (N_13002,N_11695,N_10858);
nor U13003 (N_13003,N_12308,N_11361);
or U13004 (N_13004,N_10849,N_10568);
nand U13005 (N_13005,N_10233,N_10753);
xnor U13006 (N_13006,N_11442,N_11863);
and U13007 (N_13007,N_12250,N_11777);
or U13008 (N_13008,N_10171,N_11961);
xor U13009 (N_13009,N_11423,N_11046);
and U13010 (N_13010,N_12427,N_10692);
nand U13011 (N_13011,N_10578,N_10050);
nand U13012 (N_13012,N_10610,N_12497);
nor U13013 (N_13013,N_10121,N_12444);
nand U13014 (N_13014,N_12206,N_12442);
and U13015 (N_13015,N_10648,N_11890);
or U13016 (N_13016,N_10297,N_12412);
nand U13017 (N_13017,N_11912,N_12344);
xor U13018 (N_13018,N_10943,N_11484);
and U13019 (N_13019,N_11125,N_11597);
nand U13020 (N_13020,N_10772,N_12350);
or U13021 (N_13021,N_11774,N_10968);
or U13022 (N_13022,N_10661,N_10832);
nand U13023 (N_13023,N_11240,N_12012);
nor U13024 (N_13024,N_11242,N_11446);
or U13025 (N_13025,N_10595,N_11304);
nor U13026 (N_13026,N_12141,N_10809);
nand U13027 (N_13027,N_11569,N_11596);
or U13028 (N_13028,N_11356,N_10274);
nand U13029 (N_13029,N_10922,N_10550);
or U13030 (N_13030,N_11819,N_11237);
and U13031 (N_13031,N_10305,N_12373);
xor U13032 (N_13032,N_10113,N_12462);
nand U13033 (N_13033,N_12215,N_10756);
nand U13034 (N_13034,N_10962,N_11166);
and U13035 (N_13035,N_11274,N_12293);
nor U13036 (N_13036,N_11494,N_11024);
or U13037 (N_13037,N_10795,N_10123);
and U13038 (N_13038,N_11376,N_10878);
nor U13039 (N_13039,N_11179,N_12291);
or U13040 (N_13040,N_11112,N_11755);
nor U13041 (N_13041,N_12338,N_11857);
or U13042 (N_13042,N_12327,N_10238);
nor U13043 (N_13043,N_12255,N_10513);
nor U13044 (N_13044,N_11771,N_10624);
nor U13045 (N_13045,N_10076,N_11632);
nor U13046 (N_13046,N_10986,N_10855);
and U13047 (N_13047,N_10446,N_10620);
nor U13048 (N_13048,N_11504,N_10215);
and U13049 (N_13049,N_12399,N_12099);
nor U13050 (N_13050,N_10959,N_11253);
or U13051 (N_13051,N_10128,N_10219);
xor U13052 (N_13052,N_10875,N_10561);
nor U13053 (N_13053,N_11906,N_11707);
and U13054 (N_13054,N_10494,N_11232);
nand U13055 (N_13055,N_12268,N_10147);
and U13056 (N_13056,N_11522,N_11691);
and U13057 (N_13057,N_10579,N_11731);
or U13058 (N_13058,N_11779,N_12358);
nand U13059 (N_13059,N_12230,N_11195);
or U13060 (N_13060,N_11996,N_11959);
nor U13061 (N_13061,N_10703,N_12084);
xor U13062 (N_13062,N_11593,N_10495);
or U13063 (N_13063,N_11226,N_10751);
and U13064 (N_13064,N_11113,N_11128);
xor U13065 (N_13065,N_10170,N_10618);
and U13066 (N_13066,N_11582,N_10609);
nand U13067 (N_13067,N_10028,N_10289);
nand U13068 (N_13068,N_12022,N_12443);
nor U13069 (N_13069,N_12088,N_10912);
nand U13070 (N_13070,N_10277,N_11735);
nor U13071 (N_13071,N_12292,N_11377);
nor U13072 (N_13072,N_11653,N_11763);
and U13073 (N_13073,N_11663,N_11319);
xor U13074 (N_13074,N_12333,N_10721);
nor U13075 (N_13075,N_11587,N_11660);
nand U13076 (N_13076,N_11169,N_10029);
or U13077 (N_13077,N_11638,N_11339);
xnor U13078 (N_13078,N_11029,N_10105);
or U13079 (N_13079,N_12296,N_12381);
nor U13080 (N_13080,N_11678,N_11838);
nand U13081 (N_13081,N_11016,N_12335);
or U13082 (N_13082,N_10902,N_12257);
or U13083 (N_13083,N_10778,N_10839);
nor U13084 (N_13084,N_10075,N_11419);
or U13085 (N_13085,N_12219,N_10664);
and U13086 (N_13086,N_10674,N_10327);
nand U13087 (N_13087,N_10467,N_10211);
nand U13088 (N_13088,N_10191,N_12116);
and U13089 (N_13089,N_11794,N_10509);
xnor U13090 (N_13090,N_11436,N_11862);
nand U13091 (N_13091,N_10572,N_11923);
xor U13092 (N_13092,N_11254,N_12262);
nor U13093 (N_13093,N_10830,N_10253);
nand U13094 (N_13094,N_12259,N_12309);
and U13095 (N_13095,N_12455,N_10653);
and U13096 (N_13096,N_10929,N_11142);
or U13097 (N_13097,N_11362,N_10020);
xor U13098 (N_13098,N_11330,N_10195);
or U13099 (N_13099,N_12476,N_11835);
nor U13100 (N_13100,N_11241,N_11741);
nor U13101 (N_13101,N_11956,N_10720);
or U13102 (N_13102,N_12112,N_11355);
nand U13103 (N_13103,N_11510,N_10009);
nor U13104 (N_13104,N_12387,N_10484);
xnor U13105 (N_13105,N_12356,N_10762);
nor U13106 (N_13106,N_11409,N_10801);
nand U13107 (N_13107,N_12367,N_10790);
xor U13108 (N_13108,N_10399,N_11781);
and U13109 (N_13109,N_10372,N_11516);
nand U13110 (N_13110,N_10247,N_11965);
or U13111 (N_13111,N_10239,N_10450);
and U13112 (N_13112,N_11612,N_11231);
and U13113 (N_13113,N_11950,N_10662);
nor U13114 (N_13114,N_12415,N_12316);
nand U13115 (N_13115,N_11625,N_10081);
nand U13116 (N_13116,N_12132,N_11818);
and U13117 (N_13117,N_10329,N_12320);
and U13118 (N_13118,N_11314,N_11790);
and U13119 (N_13119,N_11690,N_12134);
nand U13120 (N_13120,N_10358,N_11021);
and U13121 (N_13121,N_12174,N_11280);
xnor U13122 (N_13122,N_10992,N_10859);
xor U13123 (N_13123,N_11842,N_11257);
xnor U13124 (N_13124,N_10143,N_10229);
or U13125 (N_13125,N_10285,N_12368);
nor U13126 (N_13126,N_10443,N_11783);
xnor U13127 (N_13127,N_11313,N_10292);
nor U13128 (N_13128,N_12235,N_11135);
nor U13129 (N_13129,N_11694,N_11987);
and U13130 (N_13130,N_10103,N_11198);
xor U13131 (N_13131,N_10048,N_10615);
or U13132 (N_13132,N_11989,N_10174);
xor U13133 (N_13133,N_12109,N_12071);
nand U13134 (N_13134,N_12473,N_12027);
nor U13135 (N_13135,N_10735,N_10575);
nor U13136 (N_13136,N_11002,N_11963);
nor U13137 (N_13137,N_12322,N_10635);
nor U13138 (N_13138,N_11398,N_11517);
or U13139 (N_13139,N_10008,N_12166);
or U13140 (N_13140,N_12231,N_12474);
xnor U13141 (N_13141,N_10383,N_12185);
xor U13142 (N_13142,N_12146,N_10342);
or U13143 (N_13143,N_11692,N_10283);
and U13144 (N_13144,N_12414,N_10556);
nand U13145 (N_13145,N_12267,N_11498);
nand U13146 (N_13146,N_11875,N_10208);
nor U13147 (N_13147,N_12359,N_10950);
nor U13148 (N_13148,N_10319,N_11138);
or U13149 (N_13149,N_12152,N_12180);
and U13150 (N_13150,N_10511,N_11700);
and U13151 (N_13151,N_10882,N_11246);
nand U13152 (N_13152,N_12478,N_12423);
nand U13153 (N_13153,N_11013,N_10154);
or U13154 (N_13154,N_12031,N_12032);
or U13155 (N_13155,N_11192,N_10463);
nand U13156 (N_13156,N_12023,N_10582);
nor U13157 (N_13157,N_12177,N_10818);
or U13158 (N_13158,N_12100,N_10543);
nand U13159 (N_13159,N_11256,N_10228);
nand U13160 (N_13160,N_10072,N_10821);
xor U13161 (N_13161,N_11584,N_10906);
or U13162 (N_13162,N_10911,N_10346);
nor U13163 (N_13163,N_11288,N_10907);
nor U13164 (N_13164,N_11205,N_10085);
nor U13165 (N_13165,N_11491,N_10802);
and U13166 (N_13166,N_11457,N_10101);
and U13167 (N_13167,N_11512,N_12372);
xnor U13168 (N_13168,N_12464,N_10652);
nor U13169 (N_13169,N_11309,N_11265);
nand U13170 (N_13170,N_11476,N_10193);
xor U13171 (N_13171,N_10442,N_10879);
nor U13172 (N_13172,N_12045,N_12284);
xor U13173 (N_13173,N_10900,N_11964);
nand U13174 (N_13174,N_11206,N_10357);
and U13175 (N_13175,N_10343,N_11225);
or U13176 (N_13176,N_10112,N_10320);
or U13177 (N_13177,N_12057,N_10430);
nor U13178 (N_13178,N_10388,N_11352);
xor U13179 (N_13179,N_11590,N_10306);
xnor U13180 (N_13180,N_11579,N_10362);
and U13181 (N_13181,N_10520,N_10857);
xnor U13182 (N_13182,N_11914,N_11199);
and U13183 (N_13183,N_10564,N_10309);
nor U13184 (N_13184,N_10739,N_10025);
or U13185 (N_13185,N_12208,N_12183);
xor U13186 (N_13186,N_10944,N_10682);
and U13187 (N_13187,N_12376,N_10099);
or U13188 (N_13188,N_11761,N_12161);
and U13189 (N_13189,N_10896,N_11874);
and U13190 (N_13190,N_11019,N_11637);
and U13191 (N_13191,N_11759,N_11769);
xor U13192 (N_13192,N_11909,N_10470);
nand U13193 (N_13193,N_10919,N_10744);
and U13194 (N_13194,N_10259,N_10786);
and U13195 (N_13195,N_11836,N_11094);
nand U13196 (N_13196,N_12078,N_10675);
or U13197 (N_13197,N_11305,N_12020);
and U13198 (N_13198,N_12435,N_11704);
nand U13199 (N_13199,N_10980,N_10870);
and U13200 (N_13200,N_10515,N_10489);
and U13201 (N_13201,N_10716,N_12019);
nor U13202 (N_13202,N_11622,N_10053);
or U13203 (N_13203,N_11528,N_10714);
and U13204 (N_13204,N_11841,N_11954);
xnor U13205 (N_13205,N_10151,N_10337);
nor U13206 (N_13206,N_12017,N_10792);
nor U13207 (N_13207,N_11868,N_11258);
xnor U13208 (N_13208,N_11751,N_12142);
nand U13209 (N_13209,N_10389,N_12332);
and U13210 (N_13210,N_12182,N_11208);
xor U13211 (N_13211,N_11186,N_11997);
nand U13212 (N_13212,N_11608,N_10148);
nor U13213 (N_13213,N_11537,N_12066);
nand U13214 (N_13214,N_11057,N_11044);
or U13215 (N_13215,N_11897,N_11003);
and U13216 (N_13216,N_10812,N_10397);
or U13217 (N_13217,N_10967,N_11025);
nor U13218 (N_13218,N_11662,N_12390);
nor U13219 (N_13219,N_10727,N_11068);
xor U13220 (N_13220,N_10324,N_10351);
nand U13221 (N_13221,N_10702,N_11723);
nor U13222 (N_13222,N_10707,N_11392);
xnor U13223 (N_13223,N_11123,N_11867);
xnor U13224 (N_13224,N_10243,N_10766);
nor U13225 (N_13225,N_11899,N_10344);
xnor U13226 (N_13226,N_10404,N_11829);
nor U13227 (N_13227,N_10251,N_10833);
xor U13228 (N_13228,N_10483,N_11515);
nand U13229 (N_13229,N_10659,N_10067);
xnor U13230 (N_13230,N_10256,N_11109);
or U13231 (N_13231,N_11631,N_11817);
nor U13232 (N_13232,N_10255,N_11472);
or U13233 (N_13233,N_10304,N_10110);
nand U13234 (N_13234,N_12382,N_12007);
and U13235 (N_13235,N_11440,N_12191);
nor U13236 (N_13236,N_10724,N_11749);
and U13237 (N_13237,N_10710,N_10897);
xor U13238 (N_13238,N_11368,N_11713);
xor U13239 (N_13239,N_11646,N_10079);
or U13240 (N_13240,N_11250,N_12053);
nand U13241 (N_13241,N_10176,N_11315);
or U13242 (N_13242,N_12148,N_11421);
nor U13243 (N_13243,N_11586,N_10939);
nand U13244 (N_13244,N_10951,N_12212);
and U13245 (N_13245,N_12010,N_11230);
and U13246 (N_13246,N_11881,N_12113);
nand U13247 (N_13247,N_10794,N_10873);
or U13248 (N_13248,N_11030,N_11933);
xnor U13249 (N_13249,N_11396,N_11085);
and U13250 (N_13250,N_11191,N_12310);
and U13251 (N_13251,N_11243,N_10405);
xor U13252 (N_13252,N_10805,N_11858);
nor U13253 (N_13253,N_10969,N_10180);
nor U13254 (N_13254,N_10269,N_12067);
or U13255 (N_13255,N_11317,N_11455);
nand U13256 (N_13256,N_11180,N_12175);
and U13257 (N_13257,N_10693,N_10003);
xnor U13258 (N_13258,N_10780,N_10044);
and U13259 (N_13259,N_12077,N_11944);
nand U13260 (N_13260,N_11942,N_11687);
nand U13261 (N_13261,N_12452,N_10531);
xnor U13262 (N_13262,N_10436,N_11715);
nand U13263 (N_13263,N_11441,N_10623);
nor U13264 (N_13264,N_10298,N_11235);
and U13265 (N_13265,N_10146,N_11247);
nand U13266 (N_13266,N_10240,N_10545);
or U13267 (N_13267,N_10039,N_10819);
nor U13268 (N_13268,N_12357,N_10761);
nor U13269 (N_13269,N_11943,N_11647);
nor U13270 (N_13270,N_10482,N_10988);
and U13271 (N_13271,N_12143,N_10458);
xor U13272 (N_13272,N_12006,N_11851);
nand U13273 (N_13273,N_11233,N_10396);
nor U13274 (N_13274,N_11306,N_10640);
xnor U13275 (N_13275,N_10521,N_11614);
or U13276 (N_13276,N_10134,N_10369);
xor U13277 (N_13277,N_10861,N_12424);
nand U13278 (N_13278,N_11822,N_11155);
nor U13279 (N_13279,N_11425,N_10196);
nor U13280 (N_13280,N_11811,N_11702);
and U13281 (N_13281,N_10411,N_11789);
nand U13282 (N_13282,N_10333,N_10854);
and U13283 (N_13283,N_12108,N_10512);
nor U13284 (N_13284,N_11014,N_10137);
nor U13285 (N_13285,N_11533,N_12451);
xor U13286 (N_13286,N_11093,N_10058);
nor U13287 (N_13287,N_11018,N_10848);
or U13288 (N_13288,N_12281,N_10477);
or U13289 (N_13289,N_12256,N_10715);
xor U13290 (N_13290,N_10614,N_10185);
and U13291 (N_13291,N_10777,N_10771);
nor U13292 (N_13292,N_10419,N_11005);
xnor U13293 (N_13293,N_10734,N_11103);
nand U13294 (N_13294,N_11045,N_11072);
and U13295 (N_13295,N_11325,N_11534);
or U13296 (N_13296,N_11308,N_11557);
or U13297 (N_13297,N_11341,N_11814);
nand U13298 (N_13298,N_10270,N_10932);
nor U13299 (N_13299,N_11570,N_11768);
or U13300 (N_13300,N_10311,N_10338);
or U13301 (N_13301,N_11816,N_11507);
and U13302 (N_13302,N_11605,N_10023);
and U13303 (N_13303,N_12260,N_10836);
and U13304 (N_13304,N_11775,N_12189);
or U13305 (N_13305,N_10551,N_10014);
and U13306 (N_13306,N_11126,N_10964);
xnor U13307 (N_13307,N_12021,N_12041);
or U13308 (N_13308,N_10757,N_11338);
xor U13309 (N_13309,N_12083,N_11130);
nor U13310 (N_13310,N_11898,N_10914);
nand U13311 (N_13311,N_10745,N_10636);
nor U13312 (N_13312,N_10356,N_10894);
nand U13313 (N_13313,N_12432,N_11331);
or U13314 (N_13314,N_10321,N_10738);
nor U13315 (N_13315,N_12418,N_10158);
or U13316 (N_13316,N_12124,N_11974);
xnor U13317 (N_13317,N_11054,N_11583);
nor U13318 (N_13318,N_11172,N_11366);
xor U13319 (N_13319,N_10037,N_10534);
nand U13320 (N_13320,N_12233,N_11710);
nor U13321 (N_13321,N_10845,N_11568);
xnor U13322 (N_13322,N_11162,N_12445);
xor U13323 (N_13323,N_10230,N_12149);
nor U13324 (N_13324,N_10985,N_10131);
xnor U13325 (N_13325,N_10729,N_10062);
and U13326 (N_13326,N_10749,N_11600);
and U13327 (N_13327,N_11292,N_10293);
and U13328 (N_13328,N_10711,N_11957);
xor U13329 (N_13329,N_10607,N_10300);
or U13330 (N_13330,N_11839,N_11886);
and U13331 (N_13331,N_10315,N_12131);
and U13332 (N_13332,N_10296,N_11238);
xnor U13333 (N_13333,N_10637,N_11855);
nor U13334 (N_13334,N_10760,N_11711);
nor U13335 (N_13335,N_10206,N_10921);
nand U13336 (N_13336,N_11770,N_11548);
xnor U13337 (N_13337,N_11535,N_10261);
and U13338 (N_13338,N_11055,N_11473);
or U13339 (N_13339,N_11588,N_11387);
nand U13340 (N_13340,N_12122,N_10956);
xnor U13341 (N_13341,N_10129,N_11453);
nor U13342 (N_13342,N_12105,N_11561);
and U13343 (N_13343,N_10400,N_11426);
xnor U13344 (N_13344,N_11163,N_10909);
or U13345 (N_13345,N_11995,N_10576);
nand U13346 (N_13346,N_12133,N_12254);
nand U13347 (N_13347,N_12091,N_10034);
nor U13348 (N_13348,N_10928,N_10593);
xnor U13349 (N_13349,N_12258,N_12247);
nand U13350 (N_13350,N_11461,N_12117);
nand U13351 (N_13351,N_11630,N_11998);
or U13352 (N_13352,N_11127,N_11332);
nor U13353 (N_13353,N_10010,N_10013);
and U13354 (N_13354,N_12097,N_10646);
nor U13355 (N_13355,N_11931,N_11286);
or U13356 (N_13356,N_10314,N_10332);
nor U13357 (N_13357,N_10491,N_11202);
or U13358 (N_13358,N_11747,N_10983);
xor U13359 (N_13359,N_11178,N_11559);
and U13360 (N_13360,N_10468,N_12242);
nor U13361 (N_13361,N_10649,N_10528);
nand U13362 (N_13362,N_11981,N_10934);
and U13363 (N_13363,N_10210,N_10166);
or U13364 (N_13364,N_10127,N_10464);
or U13365 (N_13365,N_10094,N_11930);
xor U13366 (N_13366,N_11992,N_11438);
xnor U13367 (N_13367,N_10163,N_12384);
or U13368 (N_13368,N_10608,N_10183);
and U13369 (N_13369,N_12265,N_10869);
and U13370 (N_13370,N_11846,N_12095);
xnor U13371 (N_13371,N_10665,N_10502);
nand U13372 (N_13372,N_10179,N_12129);
nand U13373 (N_13373,N_11976,N_12171);
or U13374 (N_13374,N_12429,N_10033);
and U13375 (N_13375,N_12334,N_11261);
and U13376 (N_13376,N_11910,N_11558);
nor U13377 (N_13377,N_11592,N_10061);
nor U13378 (N_13378,N_11273,N_11095);
nand U13379 (N_13379,N_10156,N_11708);
or U13380 (N_13380,N_10084,N_12024);
nor U13381 (N_13381,N_10412,N_10666);
or U13382 (N_13382,N_10591,N_10597);
nand U13383 (N_13383,N_11739,N_11010);
xnor U13384 (N_13384,N_10594,N_11122);
nand U13385 (N_13385,N_10250,N_11734);
or U13386 (N_13386,N_12386,N_10853);
and U13387 (N_13387,N_10431,N_10433);
nand U13388 (N_13388,N_10856,N_10429);
xor U13389 (N_13389,N_10827,N_10177);
and U13390 (N_13390,N_10004,N_11201);
nor U13391 (N_13391,N_10973,N_12194);
or U13392 (N_13392,N_12253,N_12348);
or U13393 (N_13393,N_12297,N_11478);
or U13394 (N_13394,N_12426,N_11994);
nand U13395 (N_13395,N_11815,N_11049);
nor U13396 (N_13396,N_11459,N_12273);
and U13397 (N_13397,N_12106,N_12136);
and U13398 (N_13398,N_10957,N_11785);
nor U13399 (N_13399,N_10697,N_11758);
and U13400 (N_13400,N_11482,N_10996);
and U13401 (N_13401,N_11823,N_11086);
and U13402 (N_13402,N_10199,N_11677);
or U13403 (N_13403,N_11437,N_11324);
or U13404 (N_13404,N_11117,N_11477);
nor U13405 (N_13405,N_11275,N_11902);
nand U13406 (N_13406,N_11454,N_10466);
and U13407 (N_13407,N_10548,N_11706);
nand U13408 (N_13408,N_11518,N_10823);
xnor U13409 (N_13409,N_10355,N_11001);
nor U13410 (N_13410,N_12457,N_11148);
or U13411 (N_13411,N_11767,N_10984);
nand U13412 (N_13412,N_11483,N_11141);
xor U13413 (N_13413,N_10407,N_10120);
nor U13414 (N_13414,N_11497,N_11078);
xnor U13415 (N_13415,N_10065,N_11849);
xor U13416 (N_13416,N_10479,N_12282);
and U13417 (N_13417,N_11489,N_11927);
nor U13418 (N_13418,N_10307,N_11578);
or U13419 (N_13419,N_11594,N_11820);
nor U13420 (N_13420,N_11560,N_10750);
and U13421 (N_13421,N_10334,N_11311);
nand U13422 (N_13422,N_10046,N_10082);
and U13423 (N_13423,N_11251,N_10800);
or U13424 (N_13424,N_11075,N_10966);
or U13425 (N_13425,N_10647,N_10600);
nand U13426 (N_13426,N_10881,N_12128);
xor U13427 (N_13427,N_10977,N_12351);
xor U13428 (N_13428,N_11492,N_10438);
and U13429 (N_13429,N_11404,N_12075);
nand U13430 (N_13430,N_11263,N_10114);
nor U13431 (N_13431,N_11576,N_12111);
and U13432 (N_13432,N_11008,N_10475);
and U13433 (N_13433,N_11463,N_12311);
nor U13434 (N_13434,N_11327,N_12204);
nor U13435 (N_13435,N_11806,N_12217);
and U13436 (N_13436,N_12096,N_11947);
xnor U13437 (N_13437,N_10974,N_10448);
or U13438 (N_13438,N_10160,N_11536);
nor U13439 (N_13439,N_10642,N_12329);
xnor U13440 (N_13440,N_10435,N_10249);
or U13441 (N_13441,N_10077,N_12413);
nand U13442 (N_13442,N_10425,N_10622);
xor U13443 (N_13443,N_10743,N_11703);
or U13444 (N_13444,N_10815,N_11797);
nor U13445 (N_13445,N_12264,N_10767);
xor U13446 (N_13446,N_10987,N_10410);
nor U13447 (N_13447,N_12339,N_11880);
or U13448 (N_13448,N_10262,N_10286);
and U13449 (N_13449,N_11121,N_12210);
nand U13450 (N_13450,N_10669,N_10868);
xor U13451 (N_13451,N_11809,N_11287);
nand U13452 (N_13452,N_10281,N_12038);
xnor U13453 (N_13453,N_10080,N_11882);
nand U13454 (N_13454,N_12178,N_11796);
and U13455 (N_13455,N_11295,N_11606);
xnor U13456 (N_13456,N_10880,N_11937);
or U13457 (N_13457,N_10691,N_12203);
xor U13458 (N_13458,N_10403,N_10524);
nor U13459 (N_13459,N_12408,N_11540);
and U13460 (N_13460,N_12198,N_11347);
or U13461 (N_13461,N_11203,N_11762);
and U13462 (N_13462,N_10460,N_10060);
nor U13463 (N_13463,N_10119,N_11740);
nand U13464 (N_13464,N_10178,N_10379);
or U13465 (N_13465,N_12025,N_11869);
nand U13466 (N_13466,N_11585,N_12065);
xnor U13467 (N_13467,N_12040,N_12139);
and U13468 (N_13468,N_11674,N_11408);
nand U13469 (N_13469,N_10017,N_10583);
nor U13470 (N_13470,N_10418,N_10899);
or U13471 (N_13471,N_10091,N_12138);
nand U13472 (N_13472,N_10680,N_12290);
or U13473 (N_13473,N_10558,N_12087);
nand U13474 (N_13474,N_11189,N_10284);
and U13475 (N_13475,N_11165,N_12447);
or U13476 (N_13476,N_11303,N_10360);
nor U13477 (N_13477,N_10043,N_11935);
and U13478 (N_13478,N_11267,N_11043);
nor U13479 (N_13479,N_10175,N_10599);
nor U13480 (N_13480,N_10546,N_10963);
and U13481 (N_13481,N_10706,N_12055);
nor U13482 (N_13482,N_10764,N_11038);
and U13483 (N_13483,N_12013,N_10619);
nand U13484 (N_13484,N_10590,N_11866);
or U13485 (N_13485,N_10398,N_10613);
xor U13486 (N_13486,N_11248,N_11648);
or U13487 (N_13487,N_12394,N_11655);
nor U13488 (N_13488,N_11416,N_12015);
and U13489 (N_13489,N_11371,N_10339);
or U13490 (N_13490,N_10133,N_11754);
nand U13491 (N_13491,N_10876,N_12482);
or U13492 (N_13492,N_10038,N_10736);
nand U13493 (N_13493,N_10748,N_11668);
or U13494 (N_13494,N_11503,N_10382);
xnor U13495 (N_13495,N_11894,N_12395);
nand U13496 (N_13496,N_11873,N_11445);
xnor U13497 (N_13497,N_10252,N_10207);
or U13498 (N_13498,N_11951,N_12459);
nand U13499 (N_13499,N_12079,N_10364);
and U13500 (N_13500,N_12343,N_12326);
nor U13501 (N_13501,N_12127,N_12008);
or U13502 (N_13502,N_11566,N_10459);
xnor U13503 (N_13503,N_10723,N_12205);
and U13504 (N_13504,N_11896,N_10758);
xnor U13505 (N_13505,N_11084,N_10093);
or U13506 (N_13506,N_11020,N_10011);
nand U13507 (N_13507,N_11530,N_11883);
and U13508 (N_13508,N_10282,N_12422);
nand U13509 (N_13509,N_11388,N_10588);
or U13510 (N_13510,N_10655,N_11544);
xor U13511 (N_13511,N_10532,N_10204);
or U13512 (N_13512,N_10741,N_11023);
xor U13513 (N_13513,N_10401,N_12460);
xnor U13514 (N_13514,N_10639,N_12400);
xnor U13515 (N_13515,N_10580,N_12014);
nand U13516 (N_13516,N_10840,N_10165);
nand U13517 (N_13517,N_11079,N_10361);
xnor U13518 (N_13518,N_10392,N_11401);
or U13519 (N_13519,N_11012,N_10107);
or U13520 (N_13520,N_11780,N_11717);
xnor U13521 (N_13521,N_11527,N_10841);
xor U13522 (N_13522,N_11399,N_10933);
and U13523 (N_13523,N_10312,N_10272);
nand U13524 (N_13524,N_11328,N_12056);
nand U13525 (N_13525,N_10267,N_10490);
and U13526 (N_13526,N_10732,N_10935);
xnor U13527 (N_13527,N_11349,N_11922);
or U13528 (N_13528,N_11133,N_10717);
xor U13529 (N_13529,N_10124,N_12193);
and U13530 (N_13530,N_11742,N_11393);
nor U13531 (N_13531,N_11807,N_10903);
nor U13532 (N_13532,N_11595,N_12304);
and U13533 (N_13533,N_11340,N_10375);
nor U13534 (N_13534,N_11211,N_10390);
nor U13535 (N_13535,N_11017,N_11299);
nand U13536 (N_13536,N_11009,N_12366);
and U13537 (N_13537,N_11953,N_11196);
nand U13538 (N_13538,N_12270,N_11666);
or U13539 (N_13539,N_11143,N_11418);
xnor U13540 (N_13540,N_12245,N_11249);
nand U13541 (N_13541,N_10098,N_10971);
nor U13542 (N_13542,N_11725,N_10157);
nand U13543 (N_13543,N_12370,N_10976);
or U13544 (N_13544,N_10402,N_12288);
nor U13545 (N_13545,N_12085,N_10554);
or U13546 (N_13546,N_11395,N_11092);
nand U13547 (N_13547,N_10918,N_10700);
nor U13548 (N_13548,N_11026,N_10898);
nor U13549 (N_13549,N_10198,N_12246);
and U13550 (N_13550,N_11990,N_12383);
nor U13551 (N_13551,N_11479,N_12336);
nor U13552 (N_13552,N_10041,N_10789);
or U13553 (N_13553,N_12391,N_10954);
xor U13554 (N_13554,N_11139,N_11772);
nor U13555 (N_13555,N_11626,N_12345);
nand U13556 (N_13556,N_10386,N_10688);
and U13557 (N_13557,N_11784,N_10544);
xor U13558 (N_13558,N_11808,N_11615);
xor U13559 (N_13559,N_10310,N_10671);
and U13560 (N_13560,N_11229,N_11885);
nor U13561 (N_13561,N_10415,N_10719);
nand U13562 (N_13562,N_12434,N_10197);
or U13563 (N_13563,N_10713,N_12061);
or U13564 (N_13564,N_12072,N_10054);
or U13565 (N_13565,N_10826,N_11060);
nor U13566 (N_13566,N_10485,N_10847);
and U13567 (N_13567,N_10526,N_12479);
or U13568 (N_13568,N_12272,N_11207);
and U13569 (N_13569,N_12341,N_10628);
nor U13570 (N_13570,N_10676,N_11799);
nor U13571 (N_13571,N_10698,N_10793);
and U13572 (N_13572,N_11888,N_12042);
or U13573 (N_13573,N_12154,N_10507);
or U13574 (N_13574,N_12003,N_11488);
or U13575 (N_13575,N_12485,N_12243);
and U13576 (N_13576,N_10071,N_11098);
or U13577 (N_13577,N_11323,N_12378);
xor U13578 (N_13578,N_11813,N_11602);
nor U13579 (N_13579,N_11879,N_10370);
xor U13580 (N_13580,N_12298,N_10785);
nand U13581 (N_13581,N_10535,N_11581);
xor U13582 (N_13582,N_10905,N_10625);
nand U13583 (N_13583,N_11227,N_12058);
xor U13584 (N_13584,N_11940,N_11555);
and U13585 (N_13585,N_10275,N_11111);
and U13586 (N_13586,N_10774,N_10519);
and U13587 (N_13587,N_11134,N_12135);
nand U13588 (N_13588,N_11671,N_10656);
or U13589 (N_13589,N_11908,N_11475);
nand U13590 (N_13590,N_11960,N_11389);
and U13591 (N_13591,N_11939,N_10216);
nor U13592 (N_13592,N_10765,N_11140);
or U13593 (N_13593,N_10851,N_11083);
xnor U13594 (N_13594,N_11824,N_11651);
xor U13595 (N_13595,N_10617,N_12073);
nor U13596 (N_13596,N_10555,N_11567);
nand U13597 (N_13597,N_10638,N_10498);
or U13598 (N_13598,N_11255,N_11096);
nor U13599 (N_13599,N_11659,N_11738);
or U13600 (N_13600,N_10557,N_11645);
and U13601 (N_13601,N_10990,N_12306);
and U13602 (N_13602,N_10953,N_10999);
and U13603 (N_13603,N_10394,N_11118);
or U13604 (N_13604,N_10887,N_11511);
nor U13605 (N_13605,N_11066,N_11552);
xor U13606 (N_13606,N_10844,N_11911);
nand U13607 (N_13607,N_12364,N_12092);
and U13608 (N_13608,N_11520,N_11565);
xnor U13609 (N_13609,N_10348,N_12029);
or U13610 (N_13610,N_10291,N_10621);
or U13611 (N_13611,N_11310,N_12496);
nor U13612 (N_13612,N_10842,N_11406);
nand U13613 (N_13613,N_10257,N_10278);
nand U13614 (N_13614,N_10893,N_11716);
xnor U13615 (N_13615,N_12277,N_12389);
nor U13616 (N_13616,N_11270,N_11407);
or U13617 (N_13617,N_11801,N_12302);
nand U13618 (N_13618,N_10271,N_12425);
and U13619 (N_13619,N_11556,N_11980);
xor U13620 (N_13620,N_11493,N_10222);
or U13621 (N_13621,N_10508,N_11158);
and U13622 (N_13622,N_10867,N_12248);
xor U13623 (N_13623,N_12280,N_10349);
or U13624 (N_13624,N_12244,N_11283);
nor U13625 (N_13625,N_11234,N_10808);
nand U13626 (N_13626,N_11676,N_10245);
nand U13627 (N_13627,N_10955,N_11714);
and U13628 (N_13628,N_10552,N_12089);
nand U13629 (N_13629,N_10260,N_11701);
and U13630 (N_13630,N_10263,N_10453);
and U13631 (N_13631,N_11900,N_11124);
or U13632 (N_13632,N_11599,N_10434);
xnor U13633 (N_13633,N_10505,N_12199);
and U13634 (N_13634,N_10380,N_10202);
and U13635 (N_13635,N_11222,N_10643);
xnor U13636 (N_13636,N_12202,N_11363);
nor U13637 (N_13637,N_11144,N_10002);
and U13638 (N_13638,N_11131,N_11467);
xnor U13639 (N_13639,N_12317,N_11217);
or U13640 (N_13640,N_11934,N_10501);
nand U13641 (N_13641,N_10217,N_10073);
and U13642 (N_13642,N_10445,N_11652);
and U13643 (N_13643,N_10831,N_11000);
xor U13644 (N_13644,N_12051,N_10426);
nand U13645 (N_13645,N_11649,N_10188);
nor U13646 (N_13646,N_12236,N_10367);
or U13647 (N_13647,N_10796,N_10972);
nor U13648 (N_13648,N_12416,N_10602);
or U13649 (N_13649,N_10111,N_12207);
or U13650 (N_13650,N_10019,N_11443);
xnor U13651 (N_13651,N_11214,N_12157);
xor U13652 (N_13652,N_10192,N_11432);
nand U13653 (N_13653,N_10681,N_11136);
nor U13654 (N_13654,N_10658,N_10182);
nor U13655 (N_13655,N_10472,N_12276);
and U13656 (N_13656,N_10451,N_10432);
nor U13657 (N_13657,N_10629,N_12155);
nand U13658 (N_13658,N_10677,N_10026);
and U13659 (N_13659,N_10365,N_12063);
xnor U13660 (N_13660,N_12312,N_10589);
nor U13661 (N_13661,N_10473,N_10087);
or U13662 (N_13662,N_11212,N_10632);
and U13663 (N_13663,N_11665,N_11753);
nand U13664 (N_13664,N_10612,N_10395);
or U13665 (N_13665,N_10890,N_11429);
and U13666 (N_13666,N_11853,N_11792);
nor U13667 (N_13667,N_11041,N_11847);
and U13668 (N_13668,N_10421,N_11289);
nand U13669 (N_13669,N_11636,N_11795);
xnor U13670 (N_13670,N_10631,N_10530);
and U13671 (N_13671,N_11696,N_12371);
or U13672 (N_13672,N_10057,N_11788);
and U13673 (N_13673,N_10036,N_10553);
or U13674 (N_13674,N_11591,N_10689);
xor U13675 (N_13675,N_12184,N_10926);
or U13676 (N_13676,N_12481,N_11840);
and U13677 (N_13677,N_11007,N_11697);
nand U13678 (N_13678,N_12163,N_10417);
nand U13679 (N_13679,N_11369,N_11351);
and U13680 (N_13680,N_10503,N_10266);
and U13681 (N_13681,N_10145,N_11435);
or U13682 (N_13682,N_11091,N_11727);
nand U13683 (N_13683,N_12440,N_12082);
xnor U13684 (N_13684,N_12396,N_11336);
nand U13685 (N_13685,N_11089,N_12355);
and U13686 (N_13686,N_11978,N_10122);
nor U13687 (N_13687,N_10015,N_10930);
and U13688 (N_13688,N_11106,N_12126);
xor U13689 (N_13689,N_10788,N_11080);
xnor U13690 (N_13690,N_10504,N_11268);
or U13691 (N_13691,N_12220,N_12274);
xnor U13692 (N_13692,N_11508,N_10092);
nor U13693 (N_13693,N_11658,N_10140);
and U13694 (N_13694,N_10603,N_10223);
xor U13695 (N_13695,N_11589,N_11967);
nand U13696 (N_13696,N_12062,N_11104);
and U13697 (N_13697,N_10843,N_10027);
nand U13698 (N_13698,N_11523,N_11228);
nand U13699 (N_13699,N_10775,N_10541);
xnor U13700 (N_13700,N_10803,N_11564);
nand U13701 (N_13701,N_10406,N_12430);
nor U13702 (N_13702,N_10975,N_11344);
nand U13703 (N_13703,N_10728,N_10787);
and U13704 (N_13704,N_10487,N_10378);
or U13705 (N_13705,N_10045,N_11381);
or U13706 (N_13706,N_12489,N_12409);
nand U13707 (N_13707,N_11210,N_11895);
or U13708 (N_13708,N_11812,N_11550);
xnor U13709 (N_13709,N_10668,N_12472);
and U13710 (N_13710,N_10024,N_10049);
nor U13711 (N_13711,N_11904,N_11145);
xnor U13712 (N_13712,N_12318,N_10657);
and U13713 (N_13713,N_10565,N_10500);
xor U13714 (N_13714,N_11065,N_12160);
nor U13715 (N_13715,N_10961,N_11745);
and U13716 (N_13716,N_11689,N_10408);
nand U13717 (N_13717,N_11107,N_10644);
nand U13718 (N_13718,N_12469,N_12328);
and U13719 (N_13719,N_11439,N_12404);
or U13720 (N_13720,N_12453,N_10461);
nand U13721 (N_13721,N_12239,N_10220);
nand U13722 (N_13722,N_11682,N_12405);
xnor U13723 (N_13723,N_11329,N_10273);
nor U13724 (N_13724,N_12064,N_10074);
xor U13725 (N_13725,N_12493,N_11405);
xnor U13726 (N_13726,N_11629,N_11028);
nor U13727 (N_13727,N_11575,N_10936);
or U13728 (N_13728,N_11390,N_11451);
or U13729 (N_13729,N_12187,N_12340);
nand U13730 (N_13730,N_10601,N_11554);
xor U13731 (N_13731,N_12401,N_12278);
nor U13732 (N_13732,N_10090,N_11087);
nand U13733 (N_13733,N_12439,N_12319);
or U13734 (N_13734,N_11776,N_10822);
or U13735 (N_13735,N_10118,N_11635);
or U13736 (N_13736,N_11975,N_11160);
and U13737 (N_13737,N_11335,N_11182);
nand U13738 (N_13738,N_12165,N_11200);
nand U13739 (N_13739,N_10205,N_10052);
or U13740 (N_13740,N_12410,N_10941);
xor U13741 (N_13741,N_12039,N_10759);
or U13742 (N_13742,N_10945,N_12197);
or U13743 (N_13743,N_10424,N_11431);
and U13744 (N_13744,N_12486,N_10497);
or U13745 (N_13745,N_10884,N_11502);
nor U13746 (N_13746,N_11509,N_10040);
xnor U13747 (N_13747,N_10345,N_11821);
nor U13748 (N_13748,N_10663,N_11450);
nor U13749 (N_13749,N_10746,N_12498);
or U13750 (N_13750,N_12260,N_11028);
nand U13751 (N_13751,N_10244,N_10088);
and U13752 (N_13752,N_11332,N_10759);
nor U13753 (N_13753,N_12183,N_11423);
and U13754 (N_13754,N_11009,N_11419);
xor U13755 (N_13755,N_11457,N_11741);
or U13756 (N_13756,N_10001,N_11278);
nor U13757 (N_13757,N_11931,N_11121);
xnor U13758 (N_13758,N_12112,N_11144);
nand U13759 (N_13759,N_10717,N_12451);
and U13760 (N_13760,N_12375,N_10663);
nand U13761 (N_13761,N_12380,N_12474);
or U13762 (N_13762,N_11722,N_12394);
or U13763 (N_13763,N_11058,N_12051);
and U13764 (N_13764,N_11695,N_10210);
nand U13765 (N_13765,N_12474,N_12156);
and U13766 (N_13766,N_11771,N_11248);
nand U13767 (N_13767,N_10306,N_10832);
nand U13768 (N_13768,N_11121,N_10307);
or U13769 (N_13769,N_10575,N_10422);
nor U13770 (N_13770,N_11151,N_10416);
or U13771 (N_13771,N_12455,N_11977);
and U13772 (N_13772,N_10658,N_11724);
nor U13773 (N_13773,N_10375,N_11632);
or U13774 (N_13774,N_11621,N_12225);
and U13775 (N_13775,N_10223,N_10328);
or U13776 (N_13776,N_10986,N_11908);
xnor U13777 (N_13777,N_11933,N_11447);
xnor U13778 (N_13778,N_11525,N_10762);
xor U13779 (N_13779,N_10690,N_10513);
nor U13780 (N_13780,N_11201,N_12471);
xor U13781 (N_13781,N_11269,N_11118);
and U13782 (N_13782,N_10079,N_11529);
or U13783 (N_13783,N_11437,N_10278);
nor U13784 (N_13784,N_11665,N_11198);
xor U13785 (N_13785,N_11267,N_10489);
xor U13786 (N_13786,N_11554,N_11913);
xor U13787 (N_13787,N_10844,N_11942);
xnor U13788 (N_13788,N_10529,N_10401);
or U13789 (N_13789,N_11861,N_10287);
or U13790 (N_13790,N_11818,N_10659);
nand U13791 (N_13791,N_11984,N_10824);
and U13792 (N_13792,N_10408,N_11378);
or U13793 (N_13793,N_10060,N_11469);
and U13794 (N_13794,N_11173,N_10823);
xor U13795 (N_13795,N_10398,N_11968);
and U13796 (N_13796,N_12194,N_10519);
and U13797 (N_13797,N_10708,N_10477);
and U13798 (N_13798,N_12010,N_12213);
or U13799 (N_13799,N_10695,N_12340);
nor U13800 (N_13800,N_10407,N_10539);
and U13801 (N_13801,N_12024,N_11355);
and U13802 (N_13802,N_12316,N_11312);
xor U13803 (N_13803,N_10896,N_10572);
or U13804 (N_13804,N_12302,N_11082);
nor U13805 (N_13805,N_10144,N_11337);
nor U13806 (N_13806,N_10885,N_10466);
xnor U13807 (N_13807,N_11581,N_10286);
or U13808 (N_13808,N_11621,N_12330);
nor U13809 (N_13809,N_11165,N_10973);
xnor U13810 (N_13810,N_10014,N_11053);
nor U13811 (N_13811,N_10356,N_12273);
or U13812 (N_13812,N_12114,N_12189);
nand U13813 (N_13813,N_11014,N_11270);
xnor U13814 (N_13814,N_11926,N_11421);
xor U13815 (N_13815,N_12035,N_10674);
or U13816 (N_13816,N_10171,N_10889);
xnor U13817 (N_13817,N_10631,N_10932);
xor U13818 (N_13818,N_11672,N_11285);
or U13819 (N_13819,N_12069,N_10647);
and U13820 (N_13820,N_11358,N_10651);
xor U13821 (N_13821,N_10921,N_11491);
xor U13822 (N_13822,N_10494,N_11299);
nand U13823 (N_13823,N_10179,N_10994);
nand U13824 (N_13824,N_11909,N_10653);
or U13825 (N_13825,N_10327,N_10562);
nor U13826 (N_13826,N_10234,N_12103);
or U13827 (N_13827,N_10590,N_12295);
nand U13828 (N_13828,N_12122,N_11110);
nor U13829 (N_13829,N_10586,N_11939);
nor U13830 (N_13830,N_10877,N_10774);
and U13831 (N_13831,N_10982,N_11386);
nor U13832 (N_13832,N_10737,N_10573);
nand U13833 (N_13833,N_11796,N_12209);
and U13834 (N_13834,N_11201,N_11620);
and U13835 (N_13835,N_12103,N_10176);
nor U13836 (N_13836,N_11762,N_10913);
xor U13837 (N_13837,N_11308,N_11233);
and U13838 (N_13838,N_12434,N_12281);
and U13839 (N_13839,N_11764,N_11422);
or U13840 (N_13840,N_11536,N_11947);
nand U13841 (N_13841,N_11747,N_11405);
or U13842 (N_13842,N_10426,N_11313);
xor U13843 (N_13843,N_11809,N_11333);
and U13844 (N_13844,N_10421,N_10856);
nor U13845 (N_13845,N_11157,N_10457);
and U13846 (N_13846,N_11802,N_10472);
or U13847 (N_13847,N_10673,N_12271);
nor U13848 (N_13848,N_12238,N_10638);
and U13849 (N_13849,N_11760,N_11119);
or U13850 (N_13850,N_12422,N_10376);
and U13851 (N_13851,N_10006,N_11615);
and U13852 (N_13852,N_11670,N_12211);
or U13853 (N_13853,N_10621,N_11397);
nand U13854 (N_13854,N_11334,N_11212);
nand U13855 (N_13855,N_10170,N_11988);
xnor U13856 (N_13856,N_10942,N_10436);
nand U13857 (N_13857,N_11566,N_12383);
or U13858 (N_13858,N_11679,N_10861);
and U13859 (N_13859,N_11666,N_10418);
xor U13860 (N_13860,N_10689,N_12429);
xor U13861 (N_13861,N_12195,N_11936);
nand U13862 (N_13862,N_10656,N_11776);
nand U13863 (N_13863,N_10454,N_12066);
and U13864 (N_13864,N_10514,N_11264);
or U13865 (N_13865,N_11139,N_11695);
and U13866 (N_13866,N_11184,N_11106);
xor U13867 (N_13867,N_12100,N_11140);
and U13868 (N_13868,N_10213,N_10543);
xnor U13869 (N_13869,N_11523,N_12334);
or U13870 (N_13870,N_11388,N_10887);
and U13871 (N_13871,N_11654,N_10983);
or U13872 (N_13872,N_11274,N_10094);
nand U13873 (N_13873,N_10047,N_10858);
nor U13874 (N_13874,N_10279,N_12102);
xor U13875 (N_13875,N_10716,N_11516);
nand U13876 (N_13876,N_10977,N_11054);
nand U13877 (N_13877,N_11442,N_12419);
or U13878 (N_13878,N_10274,N_10661);
or U13879 (N_13879,N_12305,N_11784);
nand U13880 (N_13880,N_11855,N_10962);
and U13881 (N_13881,N_10372,N_12049);
xnor U13882 (N_13882,N_11440,N_12102);
nand U13883 (N_13883,N_12488,N_10826);
nor U13884 (N_13884,N_10524,N_10013);
nor U13885 (N_13885,N_11421,N_10740);
nor U13886 (N_13886,N_10414,N_10524);
nand U13887 (N_13887,N_10038,N_11499);
xor U13888 (N_13888,N_10353,N_11664);
nor U13889 (N_13889,N_11166,N_11314);
nor U13890 (N_13890,N_12086,N_10440);
nor U13891 (N_13891,N_10821,N_12465);
xnor U13892 (N_13892,N_11775,N_11661);
nand U13893 (N_13893,N_10982,N_10487);
or U13894 (N_13894,N_11546,N_10110);
nand U13895 (N_13895,N_11066,N_12339);
or U13896 (N_13896,N_11731,N_10477);
or U13897 (N_13897,N_10485,N_10331);
nand U13898 (N_13898,N_10023,N_12419);
nand U13899 (N_13899,N_12057,N_10102);
xnor U13900 (N_13900,N_11576,N_10085);
nor U13901 (N_13901,N_12061,N_12211);
nand U13902 (N_13902,N_11449,N_11365);
and U13903 (N_13903,N_12481,N_12112);
nor U13904 (N_13904,N_11231,N_11688);
and U13905 (N_13905,N_10137,N_10221);
xor U13906 (N_13906,N_11520,N_11203);
nor U13907 (N_13907,N_10447,N_10441);
and U13908 (N_13908,N_10688,N_10571);
and U13909 (N_13909,N_12182,N_12195);
nor U13910 (N_13910,N_12007,N_10886);
or U13911 (N_13911,N_12139,N_12180);
nor U13912 (N_13912,N_10754,N_11023);
or U13913 (N_13913,N_12433,N_10764);
xor U13914 (N_13914,N_10476,N_10038);
or U13915 (N_13915,N_11144,N_11968);
xnor U13916 (N_13916,N_12295,N_11911);
nand U13917 (N_13917,N_12454,N_10718);
nor U13918 (N_13918,N_11826,N_10720);
and U13919 (N_13919,N_11690,N_10753);
or U13920 (N_13920,N_11972,N_12475);
nor U13921 (N_13921,N_12423,N_10644);
nor U13922 (N_13922,N_10566,N_10170);
nand U13923 (N_13923,N_11289,N_11960);
nand U13924 (N_13924,N_10001,N_10085);
nor U13925 (N_13925,N_10557,N_12305);
xnor U13926 (N_13926,N_12479,N_11299);
nand U13927 (N_13927,N_10072,N_12272);
nand U13928 (N_13928,N_11487,N_11678);
nor U13929 (N_13929,N_10523,N_11514);
nand U13930 (N_13930,N_11956,N_10698);
or U13931 (N_13931,N_10695,N_10610);
or U13932 (N_13932,N_11467,N_10410);
nor U13933 (N_13933,N_10987,N_10495);
nand U13934 (N_13934,N_10276,N_11205);
or U13935 (N_13935,N_12384,N_10740);
xnor U13936 (N_13936,N_11816,N_10814);
nand U13937 (N_13937,N_10033,N_12316);
nor U13938 (N_13938,N_11081,N_11413);
or U13939 (N_13939,N_12099,N_11700);
nand U13940 (N_13940,N_11001,N_11527);
and U13941 (N_13941,N_11774,N_11403);
nand U13942 (N_13942,N_12047,N_10115);
nor U13943 (N_13943,N_11763,N_12148);
and U13944 (N_13944,N_10416,N_10024);
nor U13945 (N_13945,N_10864,N_10984);
nand U13946 (N_13946,N_10514,N_11992);
nand U13947 (N_13947,N_11301,N_12225);
or U13948 (N_13948,N_11614,N_11242);
or U13949 (N_13949,N_10388,N_10930);
xnor U13950 (N_13950,N_11283,N_10285);
and U13951 (N_13951,N_10863,N_10770);
nand U13952 (N_13952,N_12163,N_12216);
nand U13953 (N_13953,N_12316,N_12398);
or U13954 (N_13954,N_11434,N_10438);
or U13955 (N_13955,N_10988,N_10771);
nor U13956 (N_13956,N_11373,N_11959);
nand U13957 (N_13957,N_12490,N_10262);
nor U13958 (N_13958,N_10321,N_10375);
or U13959 (N_13959,N_11810,N_11980);
xnor U13960 (N_13960,N_10671,N_12074);
xnor U13961 (N_13961,N_10431,N_10661);
and U13962 (N_13962,N_11898,N_11553);
or U13963 (N_13963,N_10197,N_11401);
nor U13964 (N_13964,N_12332,N_11234);
nor U13965 (N_13965,N_12207,N_12304);
nand U13966 (N_13966,N_10490,N_10337);
nor U13967 (N_13967,N_10724,N_10039);
xnor U13968 (N_13968,N_10378,N_11113);
nor U13969 (N_13969,N_11255,N_10594);
nor U13970 (N_13970,N_11281,N_12102);
or U13971 (N_13971,N_10079,N_11058);
or U13972 (N_13972,N_11217,N_10752);
or U13973 (N_13973,N_10144,N_10592);
or U13974 (N_13974,N_11059,N_11789);
xnor U13975 (N_13975,N_12368,N_10611);
nand U13976 (N_13976,N_11054,N_12030);
nor U13977 (N_13977,N_10860,N_12207);
and U13978 (N_13978,N_10446,N_10570);
xor U13979 (N_13979,N_10659,N_11097);
and U13980 (N_13980,N_11526,N_11343);
xnor U13981 (N_13981,N_10758,N_11844);
nand U13982 (N_13982,N_10818,N_11848);
nand U13983 (N_13983,N_10480,N_10339);
nor U13984 (N_13984,N_10049,N_10146);
and U13985 (N_13985,N_10611,N_11406);
and U13986 (N_13986,N_12056,N_11340);
nor U13987 (N_13987,N_11151,N_12340);
nand U13988 (N_13988,N_11054,N_11670);
and U13989 (N_13989,N_12001,N_12246);
and U13990 (N_13990,N_10075,N_10347);
or U13991 (N_13991,N_11524,N_11559);
nand U13992 (N_13992,N_11706,N_11177);
nor U13993 (N_13993,N_10785,N_11568);
nor U13994 (N_13994,N_11278,N_10137);
or U13995 (N_13995,N_11902,N_11915);
or U13996 (N_13996,N_11873,N_12402);
or U13997 (N_13997,N_12296,N_10366);
or U13998 (N_13998,N_11086,N_10819);
nor U13999 (N_13999,N_11575,N_11432);
or U14000 (N_14000,N_10820,N_11466);
nand U14001 (N_14001,N_11929,N_11481);
or U14002 (N_14002,N_11600,N_11374);
xor U14003 (N_14003,N_12329,N_11761);
xor U14004 (N_14004,N_10129,N_10042);
nand U14005 (N_14005,N_11997,N_11238);
nor U14006 (N_14006,N_10284,N_11154);
nand U14007 (N_14007,N_11004,N_11737);
nor U14008 (N_14008,N_10394,N_10970);
and U14009 (N_14009,N_11685,N_10795);
and U14010 (N_14010,N_12220,N_11471);
nor U14011 (N_14011,N_10882,N_11638);
nor U14012 (N_14012,N_10069,N_10128);
nor U14013 (N_14013,N_11306,N_12489);
nand U14014 (N_14014,N_12421,N_10926);
or U14015 (N_14015,N_12097,N_11275);
xnor U14016 (N_14016,N_12065,N_11606);
and U14017 (N_14017,N_11201,N_11644);
nand U14018 (N_14018,N_11007,N_12286);
xor U14019 (N_14019,N_11301,N_10802);
nand U14020 (N_14020,N_10058,N_11014);
nor U14021 (N_14021,N_10517,N_10006);
xnor U14022 (N_14022,N_10328,N_11992);
xnor U14023 (N_14023,N_11264,N_11584);
nor U14024 (N_14024,N_11095,N_12355);
or U14025 (N_14025,N_12228,N_10228);
nand U14026 (N_14026,N_11386,N_11749);
and U14027 (N_14027,N_12034,N_12275);
xor U14028 (N_14028,N_12085,N_11289);
nor U14029 (N_14029,N_10876,N_10140);
nand U14030 (N_14030,N_11942,N_11395);
nor U14031 (N_14031,N_11554,N_11774);
nor U14032 (N_14032,N_12015,N_10609);
and U14033 (N_14033,N_10417,N_10496);
or U14034 (N_14034,N_10487,N_10207);
nor U14035 (N_14035,N_10727,N_10605);
xor U14036 (N_14036,N_11828,N_12161);
and U14037 (N_14037,N_10401,N_11235);
and U14038 (N_14038,N_12433,N_12196);
nand U14039 (N_14039,N_12106,N_11121);
xnor U14040 (N_14040,N_10215,N_11665);
nand U14041 (N_14041,N_10964,N_10211);
nor U14042 (N_14042,N_11079,N_12186);
nor U14043 (N_14043,N_10316,N_10774);
or U14044 (N_14044,N_10338,N_10042);
and U14045 (N_14045,N_10052,N_10778);
and U14046 (N_14046,N_10838,N_11270);
xor U14047 (N_14047,N_10068,N_11839);
or U14048 (N_14048,N_10822,N_10684);
and U14049 (N_14049,N_12245,N_11996);
or U14050 (N_14050,N_12338,N_10072);
and U14051 (N_14051,N_11541,N_10090);
and U14052 (N_14052,N_10809,N_10280);
and U14053 (N_14053,N_10946,N_11257);
or U14054 (N_14054,N_10313,N_11748);
nor U14055 (N_14055,N_11219,N_11404);
nor U14056 (N_14056,N_11113,N_11048);
xor U14057 (N_14057,N_11371,N_11340);
or U14058 (N_14058,N_10053,N_10241);
and U14059 (N_14059,N_12085,N_11753);
nand U14060 (N_14060,N_12482,N_10923);
xnor U14061 (N_14061,N_10634,N_11706);
xor U14062 (N_14062,N_11556,N_11564);
nor U14063 (N_14063,N_11299,N_10295);
nor U14064 (N_14064,N_12418,N_10152);
and U14065 (N_14065,N_11391,N_12042);
xor U14066 (N_14066,N_12172,N_12278);
nor U14067 (N_14067,N_10365,N_10931);
and U14068 (N_14068,N_10147,N_11421);
xor U14069 (N_14069,N_12297,N_11973);
nand U14070 (N_14070,N_10976,N_10896);
nor U14071 (N_14071,N_12242,N_10907);
or U14072 (N_14072,N_10647,N_11660);
and U14073 (N_14073,N_12227,N_12247);
and U14074 (N_14074,N_10423,N_11157);
or U14075 (N_14075,N_11901,N_11310);
nand U14076 (N_14076,N_10991,N_11376);
or U14077 (N_14077,N_10326,N_11224);
nand U14078 (N_14078,N_11602,N_10600);
and U14079 (N_14079,N_10137,N_11857);
xor U14080 (N_14080,N_12225,N_11357);
nand U14081 (N_14081,N_12253,N_12119);
nor U14082 (N_14082,N_11252,N_12421);
or U14083 (N_14083,N_11424,N_11198);
nor U14084 (N_14084,N_11867,N_11225);
or U14085 (N_14085,N_11847,N_10880);
nand U14086 (N_14086,N_12121,N_12324);
and U14087 (N_14087,N_11679,N_11446);
nor U14088 (N_14088,N_11959,N_12104);
nor U14089 (N_14089,N_12204,N_12234);
or U14090 (N_14090,N_11125,N_10572);
xnor U14091 (N_14091,N_10292,N_11995);
or U14092 (N_14092,N_11102,N_10889);
or U14093 (N_14093,N_10717,N_10829);
or U14094 (N_14094,N_12271,N_11128);
nor U14095 (N_14095,N_11231,N_10437);
and U14096 (N_14096,N_10683,N_11647);
nand U14097 (N_14097,N_11598,N_12232);
xor U14098 (N_14098,N_10368,N_12271);
xor U14099 (N_14099,N_10599,N_10844);
nor U14100 (N_14100,N_11779,N_11405);
and U14101 (N_14101,N_10966,N_11590);
and U14102 (N_14102,N_11921,N_11240);
and U14103 (N_14103,N_12027,N_11767);
xor U14104 (N_14104,N_10554,N_11246);
nor U14105 (N_14105,N_11665,N_11329);
and U14106 (N_14106,N_10039,N_12240);
and U14107 (N_14107,N_10305,N_10809);
and U14108 (N_14108,N_11377,N_10870);
and U14109 (N_14109,N_10921,N_10295);
xor U14110 (N_14110,N_12445,N_12185);
and U14111 (N_14111,N_12184,N_11192);
or U14112 (N_14112,N_10153,N_10322);
nor U14113 (N_14113,N_11679,N_10297);
xnor U14114 (N_14114,N_10380,N_11736);
or U14115 (N_14115,N_10134,N_10982);
nand U14116 (N_14116,N_10581,N_10358);
xor U14117 (N_14117,N_11624,N_11774);
nor U14118 (N_14118,N_10124,N_11203);
xnor U14119 (N_14119,N_11693,N_10597);
nor U14120 (N_14120,N_12476,N_12400);
and U14121 (N_14121,N_10504,N_11064);
or U14122 (N_14122,N_11241,N_11990);
and U14123 (N_14123,N_11232,N_10692);
nor U14124 (N_14124,N_12242,N_12436);
or U14125 (N_14125,N_10653,N_12015);
nor U14126 (N_14126,N_10204,N_10497);
nand U14127 (N_14127,N_10304,N_11831);
nor U14128 (N_14128,N_10818,N_12279);
xor U14129 (N_14129,N_11556,N_11756);
nand U14130 (N_14130,N_10761,N_11067);
nand U14131 (N_14131,N_11842,N_12303);
nand U14132 (N_14132,N_10573,N_10316);
nand U14133 (N_14133,N_10819,N_11823);
and U14134 (N_14134,N_10593,N_12232);
nor U14135 (N_14135,N_12080,N_12166);
or U14136 (N_14136,N_12431,N_11348);
or U14137 (N_14137,N_11703,N_10888);
nand U14138 (N_14138,N_12041,N_10841);
or U14139 (N_14139,N_10702,N_10973);
and U14140 (N_14140,N_12116,N_10022);
xnor U14141 (N_14141,N_10025,N_11145);
or U14142 (N_14142,N_11964,N_10940);
nor U14143 (N_14143,N_10750,N_11503);
nor U14144 (N_14144,N_10186,N_11584);
nand U14145 (N_14145,N_11569,N_11865);
or U14146 (N_14146,N_11049,N_11485);
nor U14147 (N_14147,N_10220,N_11984);
xnor U14148 (N_14148,N_10750,N_11628);
or U14149 (N_14149,N_10597,N_11993);
and U14150 (N_14150,N_12401,N_10771);
or U14151 (N_14151,N_11090,N_10845);
nor U14152 (N_14152,N_11320,N_11109);
xor U14153 (N_14153,N_12489,N_12490);
or U14154 (N_14154,N_10844,N_11189);
and U14155 (N_14155,N_12357,N_11240);
xnor U14156 (N_14156,N_11939,N_10603);
and U14157 (N_14157,N_11938,N_10427);
nand U14158 (N_14158,N_10990,N_11286);
nand U14159 (N_14159,N_12095,N_11673);
nand U14160 (N_14160,N_10829,N_10540);
and U14161 (N_14161,N_12162,N_10646);
or U14162 (N_14162,N_10878,N_10652);
and U14163 (N_14163,N_12177,N_10192);
nor U14164 (N_14164,N_11787,N_10371);
nor U14165 (N_14165,N_12195,N_11915);
or U14166 (N_14166,N_10778,N_11231);
and U14167 (N_14167,N_10734,N_11427);
and U14168 (N_14168,N_10116,N_11663);
nor U14169 (N_14169,N_10461,N_12226);
nand U14170 (N_14170,N_11155,N_10675);
or U14171 (N_14171,N_11485,N_12343);
nand U14172 (N_14172,N_12214,N_12392);
xor U14173 (N_14173,N_11891,N_11836);
nand U14174 (N_14174,N_11722,N_12262);
and U14175 (N_14175,N_10798,N_11161);
nor U14176 (N_14176,N_10606,N_10798);
xor U14177 (N_14177,N_10429,N_11584);
xnor U14178 (N_14178,N_11048,N_11919);
and U14179 (N_14179,N_10105,N_10836);
nor U14180 (N_14180,N_10640,N_12337);
and U14181 (N_14181,N_10614,N_10523);
nand U14182 (N_14182,N_10059,N_10072);
nor U14183 (N_14183,N_10161,N_11361);
nor U14184 (N_14184,N_11510,N_12110);
or U14185 (N_14185,N_11438,N_11281);
nor U14186 (N_14186,N_12109,N_11870);
xnor U14187 (N_14187,N_11777,N_10034);
xnor U14188 (N_14188,N_10856,N_11970);
nand U14189 (N_14189,N_10933,N_11431);
nor U14190 (N_14190,N_10691,N_11202);
and U14191 (N_14191,N_10951,N_10506);
and U14192 (N_14192,N_11000,N_11117);
nand U14193 (N_14193,N_11210,N_11419);
and U14194 (N_14194,N_12381,N_10237);
and U14195 (N_14195,N_11133,N_12383);
nor U14196 (N_14196,N_11237,N_10686);
and U14197 (N_14197,N_11194,N_10899);
xor U14198 (N_14198,N_11953,N_12293);
xor U14199 (N_14199,N_11855,N_12392);
xnor U14200 (N_14200,N_10835,N_11414);
xor U14201 (N_14201,N_12179,N_11351);
nor U14202 (N_14202,N_11217,N_11611);
and U14203 (N_14203,N_11946,N_11574);
nor U14204 (N_14204,N_11816,N_12141);
or U14205 (N_14205,N_12461,N_10879);
nor U14206 (N_14206,N_10694,N_10227);
or U14207 (N_14207,N_11566,N_11573);
xnor U14208 (N_14208,N_12103,N_10295);
and U14209 (N_14209,N_11934,N_12177);
nor U14210 (N_14210,N_11987,N_10000);
nor U14211 (N_14211,N_10916,N_11205);
and U14212 (N_14212,N_10783,N_10337);
xor U14213 (N_14213,N_12241,N_10549);
xnor U14214 (N_14214,N_11987,N_10626);
xnor U14215 (N_14215,N_11368,N_10249);
or U14216 (N_14216,N_10202,N_12353);
xnor U14217 (N_14217,N_11007,N_11943);
and U14218 (N_14218,N_10625,N_10544);
nand U14219 (N_14219,N_11028,N_10804);
nand U14220 (N_14220,N_11143,N_11367);
or U14221 (N_14221,N_11739,N_12390);
xor U14222 (N_14222,N_11154,N_11054);
or U14223 (N_14223,N_12475,N_10928);
and U14224 (N_14224,N_12331,N_10940);
and U14225 (N_14225,N_10865,N_12353);
xor U14226 (N_14226,N_10534,N_10244);
or U14227 (N_14227,N_10378,N_11581);
xnor U14228 (N_14228,N_11175,N_11431);
and U14229 (N_14229,N_11621,N_10204);
nand U14230 (N_14230,N_12443,N_12442);
xnor U14231 (N_14231,N_11584,N_11306);
and U14232 (N_14232,N_10107,N_11045);
nor U14233 (N_14233,N_10411,N_10821);
nand U14234 (N_14234,N_10988,N_11757);
xnor U14235 (N_14235,N_11919,N_12239);
xnor U14236 (N_14236,N_11742,N_11147);
nand U14237 (N_14237,N_10697,N_10864);
and U14238 (N_14238,N_10245,N_10111);
and U14239 (N_14239,N_10153,N_10928);
nor U14240 (N_14240,N_10087,N_10185);
xor U14241 (N_14241,N_10085,N_11007);
and U14242 (N_14242,N_10871,N_12108);
or U14243 (N_14243,N_12482,N_10569);
or U14244 (N_14244,N_10574,N_12280);
nand U14245 (N_14245,N_11548,N_12127);
xnor U14246 (N_14246,N_12267,N_12178);
or U14247 (N_14247,N_10403,N_10584);
or U14248 (N_14248,N_10667,N_10600);
xnor U14249 (N_14249,N_10250,N_11348);
and U14250 (N_14250,N_10856,N_12024);
and U14251 (N_14251,N_12001,N_11739);
or U14252 (N_14252,N_10834,N_12366);
nor U14253 (N_14253,N_12460,N_10168);
nor U14254 (N_14254,N_11720,N_10937);
or U14255 (N_14255,N_10230,N_12448);
nand U14256 (N_14256,N_11069,N_12438);
or U14257 (N_14257,N_12340,N_12038);
nor U14258 (N_14258,N_10593,N_10133);
nor U14259 (N_14259,N_10533,N_11987);
nor U14260 (N_14260,N_11451,N_11138);
nor U14261 (N_14261,N_12419,N_11173);
nor U14262 (N_14262,N_10280,N_10889);
or U14263 (N_14263,N_11814,N_10934);
xnor U14264 (N_14264,N_11797,N_11178);
nor U14265 (N_14265,N_10048,N_10898);
or U14266 (N_14266,N_12312,N_12452);
nor U14267 (N_14267,N_10967,N_10866);
or U14268 (N_14268,N_10597,N_11076);
and U14269 (N_14269,N_11687,N_10559);
and U14270 (N_14270,N_12346,N_10248);
nand U14271 (N_14271,N_11541,N_11726);
nand U14272 (N_14272,N_10355,N_12411);
nor U14273 (N_14273,N_10234,N_11503);
nand U14274 (N_14274,N_10197,N_10012);
nor U14275 (N_14275,N_10924,N_10281);
or U14276 (N_14276,N_10847,N_10003);
xor U14277 (N_14277,N_10264,N_11456);
and U14278 (N_14278,N_10775,N_10716);
or U14279 (N_14279,N_11614,N_10606);
or U14280 (N_14280,N_12256,N_11783);
nand U14281 (N_14281,N_11311,N_11385);
nor U14282 (N_14282,N_11831,N_12478);
nor U14283 (N_14283,N_11015,N_11273);
nand U14284 (N_14284,N_11702,N_11312);
and U14285 (N_14285,N_10625,N_10828);
nor U14286 (N_14286,N_11228,N_11437);
nor U14287 (N_14287,N_10957,N_12497);
and U14288 (N_14288,N_11700,N_11692);
or U14289 (N_14289,N_10529,N_12422);
or U14290 (N_14290,N_12204,N_11424);
xor U14291 (N_14291,N_11816,N_10119);
xor U14292 (N_14292,N_11489,N_10168);
xnor U14293 (N_14293,N_12281,N_10726);
or U14294 (N_14294,N_10420,N_10853);
nand U14295 (N_14295,N_11065,N_11947);
xor U14296 (N_14296,N_10051,N_11583);
or U14297 (N_14297,N_10260,N_10181);
nor U14298 (N_14298,N_10804,N_10937);
xnor U14299 (N_14299,N_10806,N_11479);
or U14300 (N_14300,N_10437,N_11052);
or U14301 (N_14301,N_12127,N_11299);
nor U14302 (N_14302,N_11858,N_12033);
xnor U14303 (N_14303,N_10949,N_11236);
and U14304 (N_14304,N_11866,N_12348);
nor U14305 (N_14305,N_11307,N_12060);
nand U14306 (N_14306,N_10996,N_10991);
and U14307 (N_14307,N_10564,N_11377);
and U14308 (N_14308,N_11997,N_10951);
xor U14309 (N_14309,N_10107,N_12362);
or U14310 (N_14310,N_10319,N_11374);
nor U14311 (N_14311,N_10123,N_11652);
and U14312 (N_14312,N_11043,N_11131);
and U14313 (N_14313,N_10787,N_11513);
xor U14314 (N_14314,N_11400,N_12278);
nand U14315 (N_14315,N_11580,N_10154);
nand U14316 (N_14316,N_12467,N_11736);
and U14317 (N_14317,N_10118,N_11927);
and U14318 (N_14318,N_10734,N_12406);
nor U14319 (N_14319,N_12088,N_12251);
or U14320 (N_14320,N_11180,N_11103);
xnor U14321 (N_14321,N_10145,N_11193);
nand U14322 (N_14322,N_10330,N_11128);
or U14323 (N_14323,N_10554,N_10142);
xnor U14324 (N_14324,N_11281,N_10881);
and U14325 (N_14325,N_10483,N_12494);
nor U14326 (N_14326,N_12395,N_10544);
and U14327 (N_14327,N_10186,N_11450);
nand U14328 (N_14328,N_10777,N_11809);
xnor U14329 (N_14329,N_12152,N_10032);
xnor U14330 (N_14330,N_10466,N_11063);
xor U14331 (N_14331,N_11587,N_11392);
and U14332 (N_14332,N_12056,N_10229);
nand U14333 (N_14333,N_10073,N_12064);
xor U14334 (N_14334,N_11032,N_10751);
xnor U14335 (N_14335,N_10973,N_11388);
nor U14336 (N_14336,N_12011,N_10468);
and U14337 (N_14337,N_11135,N_10407);
nor U14338 (N_14338,N_11390,N_11840);
nor U14339 (N_14339,N_11662,N_10545);
or U14340 (N_14340,N_11186,N_10817);
or U14341 (N_14341,N_10039,N_10193);
nor U14342 (N_14342,N_10892,N_11563);
nor U14343 (N_14343,N_11509,N_10237);
and U14344 (N_14344,N_11619,N_11621);
nor U14345 (N_14345,N_12168,N_11971);
nor U14346 (N_14346,N_11291,N_12333);
nor U14347 (N_14347,N_12343,N_12211);
nand U14348 (N_14348,N_12026,N_10603);
nand U14349 (N_14349,N_12113,N_11581);
nor U14350 (N_14350,N_12113,N_10246);
xnor U14351 (N_14351,N_11700,N_12445);
or U14352 (N_14352,N_10448,N_10008);
nor U14353 (N_14353,N_10594,N_11908);
xor U14354 (N_14354,N_10457,N_12075);
xnor U14355 (N_14355,N_12258,N_11145);
and U14356 (N_14356,N_12220,N_10476);
xnor U14357 (N_14357,N_12141,N_11568);
nor U14358 (N_14358,N_11917,N_11620);
and U14359 (N_14359,N_11982,N_10864);
xor U14360 (N_14360,N_11151,N_11339);
or U14361 (N_14361,N_10541,N_11531);
and U14362 (N_14362,N_10258,N_12107);
xnor U14363 (N_14363,N_11050,N_12434);
and U14364 (N_14364,N_11190,N_10988);
nor U14365 (N_14365,N_11512,N_10896);
xor U14366 (N_14366,N_10566,N_11767);
or U14367 (N_14367,N_12076,N_10946);
or U14368 (N_14368,N_12286,N_11494);
nor U14369 (N_14369,N_10339,N_10250);
and U14370 (N_14370,N_12012,N_10072);
or U14371 (N_14371,N_11790,N_11337);
or U14372 (N_14372,N_12415,N_10822);
nor U14373 (N_14373,N_11781,N_10241);
xor U14374 (N_14374,N_11480,N_12451);
xor U14375 (N_14375,N_10177,N_11310);
nor U14376 (N_14376,N_10037,N_11122);
or U14377 (N_14377,N_10630,N_12427);
xnor U14378 (N_14378,N_11986,N_11660);
or U14379 (N_14379,N_10708,N_11269);
xnor U14380 (N_14380,N_12414,N_10226);
and U14381 (N_14381,N_10464,N_11242);
nor U14382 (N_14382,N_10062,N_11190);
nand U14383 (N_14383,N_10863,N_10514);
nand U14384 (N_14384,N_12017,N_11890);
nor U14385 (N_14385,N_11174,N_11335);
xnor U14386 (N_14386,N_10728,N_10257);
nor U14387 (N_14387,N_10979,N_10128);
nor U14388 (N_14388,N_10185,N_10633);
xnor U14389 (N_14389,N_11141,N_12173);
nor U14390 (N_14390,N_10556,N_10204);
nand U14391 (N_14391,N_10895,N_12110);
xnor U14392 (N_14392,N_12159,N_12392);
nor U14393 (N_14393,N_10450,N_11366);
or U14394 (N_14394,N_12307,N_11631);
or U14395 (N_14395,N_11135,N_10108);
and U14396 (N_14396,N_11860,N_10519);
or U14397 (N_14397,N_12474,N_11509);
nand U14398 (N_14398,N_12005,N_10601);
or U14399 (N_14399,N_12181,N_12131);
nand U14400 (N_14400,N_11060,N_12170);
and U14401 (N_14401,N_12183,N_11937);
or U14402 (N_14402,N_12188,N_10624);
nor U14403 (N_14403,N_11491,N_11377);
xnor U14404 (N_14404,N_11287,N_11415);
nor U14405 (N_14405,N_11687,N_11123);
nor U14406 (N_14406,N_10114,N_12351);
xor U14407 (N_14407,N_10917,N_11325);
xor U14408 (N_14408,N_11384,N_10608);
or U14409 (N_14409,N_10634,N_11748);
or U14410 (N_14410,N_10066,N_12431);
nor U14411 (N_14411,N_11561,N_12422);
or U14412 (N_14412,N_10110,N_11647);
and U14413 (N_14413,N_10230,N_10556);
or U14414 (N_14414,N_12334,N_12022);
or U14415 (N_14415,N_10495,N_12117);
nand U14416 (N_14416,N_11174,N_11678);
and U14417 (N_14417,N_11130,N_10052);
and U14418 (N_14418,N_11682,N_10769);
nor U14419 (N_14419,N_12436,N_10666);
xnor U14420 (N_14420,N_10178,N_11034);
nand U14421 (N_14421,N_12458,N_11289);
nor U14422 (N_14422,N_10102,N_11682);
nor U14423 (N_14423,N_11420,N_10081);
xor U14424 (N_14424,N_10610,N_10214);
xor U14425 (N_14425,N_12335,N_10664);
xnor U14426 (N_14426,N_12330,N_10949);
xnor U14427 (N_14427,N_10394,N_10629);
or U14428 (N_14428,N_12097,N_10427);
xnor U14429 (N_14429,N_10311,N_11869);
nor U14430 (N_14430,N_10135,N_11969);
xnor U14431 (N_14431,N_10131,N_11225);
xnor U14432 (N_14432,N_11083,N_11284);
and U14433 (N_14433,N_10635,N_11024);
nand U14434 (N_14434,N_11027,N_12004);
nor U14435 (N_14435,N_11505,N_11878);
and U14436 (N_14436,N_12396,N_10459);
xor U14437 (N_14437,N_12456,N_10797);
xnor U14438 (N_14438,N_10822,N_11381);
nand U14439 (N_14439,N_12208,N_10252);
and U14440 (N_14440,N_11189,N_11659);
nor U14441 (N_14441,N_11425,N_10572);
or U14442 (N_14442,N_12445,N_12124);
nand U14443 (N_14443,N_11306,N_11174);
and U14444 (N_14444,N_11557,N_11894);
and U14445 (N_14445,N_12463,N_10041);
nor U14446 (N_14446,N_10038,N_10848);
or U14447 (N_14447,N_12083,N_10583);
nand U14448 (N_14448,N_11823,N_11794);
or U14449 (N_14449,N_10894,N_11583);
nor U14450 (N_14450,N_10786,N_11903);
or U14451 (N_14451,N_10964,N_10773);
or U14452 (N_14452,N_10679,N_11451);
and U14453 (N_14453,N_11960,N_10010);
xnor U14454 (N_14454,N_11208,N_11362);
and U14455 (N_14455,N_11466,N_11163);
xor U14456 (N_14456,N_10047,N_12421);
nor U14457 (N_14457,N_10069,N_10871);
or U14458 (N_14458,N_12217,N_10410);
nor U14459 (N_14459,N_11008,N_10790);
nor U14460 (N_14460,N_11229,N_11497);
nand U14461 (N_14461,N_11098,N_11175);
nand U14462 (N_14462,N_10038,N_10831);
and U14463 (N_14463,N_12212,N_10598);
nor U14464 (N_14464,N_10637,N_12256);
xnor U14465 (N_14465,N_10596,N_10888);
nor U14466 (N_14466,N_11838,N_12103);
nor U14467 (N_14467,N_11110,N_11727);
or U14468 (N_14468,N_10294,N_10350);
nand U14469 (N_14469,N_10789,N_12116);
and U14470 (N_14470,N_11309,N_11386);
and U14471 (N_14471,N_10014,N_10900);
nor U14472 (N_14472,N_10983,N_12147);
and U14473 (N_14473,N_11962,N_10828);
or U14474 (N_14474,N_11072,N_11800);
and U14475 (N_14475,N_11791,N_11320);
and U14476 (N_14476,N_10283,N_12364);
or U14477 (N_14477,N_12437,N_10004);
nand U14478 (N_14478,N_11732,N_11315);
and U14479 (N_14479,N_12395,N_10043);
xnor U14480 (N_14480,N_10131,N_11391);
xor U14481 (N_14481,N_11049,N_11678);
nand U14482 (N_14482,N_10139,N_11124);
nand U14483 (N_14483,N_12018,N_10468);
or U14484 (N_14484,N_10896,N_10101);
nand U14485 (N_14485,N_11582,N_10286);
or U14486 (N_14486,N_10840,N_10243);
xnor U14487 (N_14487,N_11601,N_12346);
or U14488 (N_14488,N_11563,N_12497);
xor U14489 (N_14489,N_11679,N_10996);
or U14490 (N_14490,N_11468,N_10342);
or U14491 (N_14491,N_11887,N_11536);
nor U14492 (N_14492,N_12210,N_11062);
and U14493 (N_14493,N_10650,N_12349);
nor U14494 (N_14494,N_11705,N_11269);
nand U14495 (N_14495,N_12184,N_11055);
and U14496 (N_14496,N_11278,N_11419);
xor U14497 (N_14497,N_11997,N_10000);
nand U14498 (N_14498,N_12268,N_10705);
nand U14499 (N_14499,N_11863,N_11808);
nor U14500 (N_14500,N_11718,N_12368);
and U14501 (N_14501,N_11486,N_12046);
or U14502 (N_14502,N_11903,N_10913);
nor U14503 (N_14503,N_10895,N_10947);
or U14504 (N_14504,N_12450,N_11299);
or U14505 (N_14505,N_12429,N_11727);
xnor U14506 (N_14506,N_10885,N_10380);
xnor U14507 (N_14507,N_10894,N_10329);
nand U14508 (N_14508,N_11456,N_12404);
nor U14509 (N_14509,N_11961,N_11380);
or U14510 (N_14510,N_10605,N_10595);
or U14511 (N_14511,N_11639,N_10463);
nand U14512 (N_14512,N_11931,N_10806);
or U14513 (N_14513,N_12478,N_11947);
and U14514 (N_14514,N_11948,N_10012);
nand U14515 (N_14515,N_10024,N_10244);
nand U14516 (N_14516,N_10595,N_12408);
nand U14517 (N_14517,N_11991,N_10233);
nand U14518 (N_14518,N_11953,N_10187);
xor U14519 (N_14519,N_11431,N_12396);
or U14520 (N_14520,N_11723,N_12241);
and U14521 (N_14521,N_12424,N_11732);
nand U14522 (N_14522,N_11187,N_11471);
or U14523 (N_14523,N_12331,N_11044);
and U14524 (N_14524,N_12388,N_10297);
nand U14525 (N_14525,N_11343,N_11906);
nor U14526 (N_14526,N_11540,N_11126);
and U14527 (N_14527,N_10575,N_10751);
and U14528 (N_14528,N_11042,N_12499);
xor U14529 (N_14529,N_11841,N_11117);
nand U14530 (N_14530,N_11078,N_10668);
and U14531 (N_14531,N_11498,N_12116);
xor U14532 (N_14532,N_12319,N_11663);
nor U14533 (N_14533,N_12478,N_10119);
nor U14534 (N_14534,N_11703,N_11440);
nor U14535 (N_14535,N_11751,N_10875);
and U14536 (N_14536,N_12169,N_11616);
nand U14537 (N_14537,N_12295,N_10990);
or U14538 (N_14538,N_10643,N_10901);
and U14539 (N_14539,N_10104,N_10895);
xnor U14540 (N_14540,N_11226,N_11168);
xor U14541 (N_14541,N_11343,N_11478);
xor U14542 (N_14542,N_12034,N_12308);
and U14543 (N_14543,N_10831,N_11165);
and U14544 (N_14544,N_10905,N_12472);
and U14545 (N_14545,N_11367,N_10037);
xor U14546 (N_14546,N_10445,N_10734);
and U14547 (N_14547,N_12202,N_12490);
nor U14548 (N_14548,N_10241,N_10140);
nand U14549 (N_14549,N_10444,N_11542);
xor U14550 (N_14550,N_11900,N_11227);
xor U14551 (N_14551,N_11564,N_11861);
nor U14552 (N_14552,N_11443,N_11168);
nand U14553 (N_14553,N_11046,N_10114);
xor U14554 (N_14554,N_10032,N_11157);
nor U14555 (N_14555,N_11778,N_11484);
or U14556 (N_14556,N_12047,N_11345);
or U14557 (N_14557,N_11534,N_11093);
and U14558 (N_14558,N_11681,N_10259);
and U14559 (N_14559,N_10369,N_11020);
or U14560 (N_14560,N_11161,N_11796);
xnor U14561 (N_14561,N_12379,N_12352);
or U14562 (N_14562,N_10641,N_11324);
nand U14563 (N_14563,N_10354,N_10742);
xnor U14564 (N_14564,N_11212,N_12394);
or U14565 (N_14565,N_10417,N_10666);
or U14566 (N_14566,N_10239,N_10844);
and U14567 (N_14567,N_12499,N_11602);
or U14568 (N_14568,N_11316,N_11121);
and U14569 (N_14569,N_10269,N_12096);
or U14570 (N_14570,N_10210,N_10818);
and U14571 (N_14571,N_11201,N_10475);
and U14572 (N_14572,N_10783,N_10015);
or U14573 (N_14573,N_10190,N_11823);
and U14574 (N_14574,N_11116,N_10699);
or U14575 (N_14575,N_12055,N_12369);
xnor U14576 (N_14576,N_10260,N_11659);
xor U14577 (N_14577,N_12153,N_11153);
and U14578 (N_14578,N_10427,N_12022);
and U14579 (N_14579,N_12070,N_11383);
nor U14580 (N_14580,N_10393,N_11970);
nor U14581 (N_14581,N_11908,N_10945);
and U14582 (N_14582,N_10138,N_11429);
or U14583 (N_14583,N_10672,N_11453);
or U14584 (N_14584,N_10680,N_10543);
xnor U14585 (N_14585,N_11982,N_10607);
nor U14586 (N_14586,N_10232,N_12376);
xnor U14587 (N_14587,N_11128,N_11994);
nand U14588 (N_14588,N_11443,N_11254);
nand U14589 (N_14589,N_12233,N_11063);
and U14590 (N_14590,N_12035,N_10720);
xor U14591 (N_14591,N_10629,N_10391);
and U14592 (N_14592,N_10309,N_11504);
nand U14593 (N_14593,N_10911,N_12089);
and U14594 (N_14594,N_11904,N_11822);
and U14595 (N_14595,N_10031,N_11258);
nor U14596 (N_14596,N_11374,N_11225);
and U14597 (N_14597,N_10125,N_10334);
nand U14598 (N_14598,N_11736,N_11799);
or U14599 (N_14599,N_11833,N_11856);
or U14600 (N_14600,N_11279,N_10436);
nor U14601 (N_14601,N_12055,N_11021);
or U14602 (N_14602,N_10986,N_12011);
or U14603 (N_14603,N_10587,N_10366);
xnor U14604 (N_14604,N_10545,N_11747);
and U14605 (N_14605,N_11377,N_11386);
or U14606 (N_14606,N_11135,N_10167);
nand U14607 (N_14607,N_12495,N_10755);
or U14608 (N_14608,N_10276,N_10249);
and U14609 (N_14609,N_10950,N_10750);
or U14610 (N_14610,N_12293,N_11552);
or U14611 (N_14611,N_11109,N_10630);
and U14612 (N_14612,N_10257,N_12354);
xor U14613 (N_14613,N_11383,N_12138);
nand U14614 (N_14614,N_10765,N_10968);
nor U14615 (N_14615,N_10521,N_12103);
nand U14616 (N_14616,N_12220,N_12375);
nand U14617 (N_14617,N_11975,N_10822);
nor U14618 (N_14618,N_10207,N_11590);
nor U14619 (N_14619,N_12357,N_11873);
nor U14620 (N_14620,N_10073,N_11240);
or U14621 (N_14621,N_12264,N_11855);
xnor U14622 (N_14622,N_11383,N_10292);
or U14623 (N_14623,N_11735,N_12061);
and U14624 (N_14624,N_12177,N_12268);
and U14625 (N_14625,N_12350,N_12046);
or U14626 (N_14626,N_11023,N_11866);
nand U14627 (N_14627,N_12272,N_12166);
xnor U14628 (N_14628,N_11265,N_10706);
and U14629 (N_14629,N_11432,N_10269);
xor U14630 (N_14630,N_11865,N_10772);
nor U14631 (N_14631,N_10180,N_11584);
or U14632 (N_14632,N_12081,N_11149);
or U14633 (N_14633,N_10588,N_11794);
nor U14634 (N_14634,N_12110,N_10072);
or U14635 (N_14635,N_11008,N_10981);
or U14636 (N_14636,N_11722,N_11329);
and U14637 (N_14637,N_11719,N_11287);
nor U14638 (N_14638,N_11159,N_12030);
or U14639 (N_14639,N_10753,N_10689);
or U14640 (N_14640,N_11358,N_12356);
or U14641 (N_14641,N_12197,N_11813);
and U14642 (N_14642,N_10893,N_10296);
xnor U14643 (N_14643,N_10003,N_12272);
nor U14644 (N_14644,N_11794,N_11425);
nand U14645 (N_14645,N_10157,N_11413);
nand U14646 (N_14646,N_11228,N_12020);
xor U14647 (N_14647,N_10599,N_12065);
nor U14648 (N_14648,N_10176,N_12409);
and U14649 (N_14649,N_11763,N_12085);
xor U14650 (N_14650,N_11020,N_10728);
or U14651 (N_14651,N_10911,N_11511);
nand U14652 (N_14652,N_12080,N_10310);
xor U14653 (N_14653,N_11862,N_11087);
and U14654 (N_14654,N_12405,N_10407);
or U14655 (N_14655,N_10097,N_10943);
xnor U14656 (N_14656,N_11271,N_10755);
nor U14657 (N_14657,N_11741,N_10296);
xor U14658 (N_14658,N_12183,N_11294);
or U14659 (N_14659,N_10696,N_11829);
nor U14660 (N_14660,N_11437,N_12123);
or U14661 (N_14661,N_11349,N_11840);
xnor U14662 (N_14662,N_12260,N_11196);
or U14663 (N_14663,N_10200,N_11084);
nand U14664 (N_14664,N_11297,N_11734);
nor U14665 (N_14665,N_10564,N_11298);
xnor U14666 (N_14666,N_10757,N_10939);
nand U14667 (N_14667,N_11906,N_11862);
xnor U14668 (N_14668,N_11853,N_10136);
and U14669 (N_14669,N_10824,N_10183);
nor U14670 (N_14670,N_10090,N_11859);
and U14671 (N_14671,N_12069,N_11338);
nand U14672 (N_14672,N_10262,N_12499);
and U14673 (N_14673,N_12151,N_10842);
nor U14674 (N_14674,N_10929,N_10800);
and U14675 (N_14675,N_10777,N_11450);
and U14676 (N_14676,N_11897,N_11811);
and U14677 (N_14677,N_11668,N_10941);
nand U14678 (N_14678,N_11203,N_11143);
nand U14679 (N_14679,N_12359,N_11566);
and U14680 (N_14680,N_11934,N_12367);
xnor U14681 (N_14681,N_10638,N_10043);
or U14682 (N_14682,N_10135,N_12473);
and U14683 (N_14683,N_12007,N_10998);
xnor U14684 (N_14684,N_10367,N_10928);
and U14685 (N_14685,N_12382,N_11453);
or U14686 (N_14686,N_10290,N_10452);
nand U14687 (N_14687,N_11571,N_10802);
or U14688 (N_14688,N_11642,N_11148);
nor U14689 (N_14689,N_11069,N_11607);
xnor U14690 (N_14690,N_12399,N_11560);
nor U14691 (N_14691,N_10999,N_11422);
xnor U14692 (N_14692,N_10801,N_12019);
nor U14693 (N_14693,N_11819,N_11288);
nand U14694 (N_14694,N_11078,N_11872);
xnor U14695 (N_14695,N_11828,N_10008);
or U14696 (N_14696,N_10486,N_11398);
or U14697 (N_14697,N_10410,N_11113);
xor U14698 (N_14698,N_11097,N_12226);
xnor U14699 (N_14699,N_10233,N_11825);
nor U14700 (N_14700,N_10129,N_11342);
and U14701 (N_14701,N_10969,N_10908);
nand U14702 (N_14702,N_11464,N_11088);
xnor U14703 (N_14703,N_12107,N_10244);
or U14704 (N_14704,N_10554,N_10567);
xor U14705 (N_14705,N_12096,N_10726);
or U14706 (N_14706,N_11462,N_11351);
nand U14707 (N_14707,N_11960,N_10156);
or U14708 (N_14708,N_11727,N_11193);
nor U14709 (N_14709,N_10405,N_10137);
nor U14710 (N_14710,N_11650,N_10250);
nor U14711 (N_14711,N_12494,N_11079);
and U14712 (N_14712,N_11442,N_10677);
nand U14713 (N_14713,N_11354,N_11626);
xor U14714 (N_14714,N_11933,N_10628);
xor U14715 (N_14715,N_10956,N_10663);
nor U14716 (N_14716,N_10660,N_11150);
xnor U14717 (N_14717,N_11123,N_10201);
or U14718 (N_14718,N_10248,N_10379);
or U14719 (N_14719,N_10993,N_12155);
and U14720 (N_14720,N_11390,N_11578);
xnor U14721 (N_14721,N_10780,N_10213);
nand U14722 (N_14722,N_11384,N_11225);
xnor U14723 (N_14723,N_10194,N_11749);
nor U14724 (N_14724,N_11223,N_12447);
xnor U14725 (N_14725,N_11238,N_10684);
or U14726 (N_14726,N_10137,N_11503);
xnor U14727 (N_14727,N_11953,N_12317);
and U14728 (N_14728,N_10240,N_10615);
and U14729 (N_14729,N_11815,N_11764);
and U14730 (N_14730,N_12039,N_11099);
xnor U14731 (N_14731,N_11984,N_11640);
nor U14732 (N_14732,N_10183,N_10026);
nor U14733 (N_14733,N_12450,N_10137);
and U14734 (N_14734,N_10618,N_11340);
xor U14735 (N_14735,N_10045,N_10962);
or U14736 (N_14736,N_11247,N_11803);
nand U14737 (N_14737,N_10882,N_12272);
and U14738 (N_14738,N_10215,N_10778);
and U14739 (N_14739,N_10548,N_12374);
nor U14740 (N_14740,N_10195,N_11575);
or U14741 (N_14741,N_12327,N_11455);
and U14742 (N_14742,N_10004,N_12005);
and U14743 (N_14743,N_10171,N_12057);
nand U14744 (N_14744,N_11669,N_10065);
or U14745 (N_14745,N_10898,N_10469);
nor U14746 (N_14746,N_10871,N_11622);
nor U14747 (N_14747,N_12037,N_10317);
or U14748 (N_14748,N_11843,N_12279);
xor U14749 (N_14749,N_11405,N_10899);
xnor U14750 (N_14750,N_10834,N_12482);
xor U14751 (N_14751,N_11668,N_10932);
xor U14752 (N_14752,N_10439,N_12039);
and U14753 (N_14753,N_11907,N_11048);
or U14754 (N_14754,N_11658,N_11068);
xnor U14755 (N_14755,N_11370,N_11815);
xor U14756 (N_14756,N_11792,N_10746);
or U14757 (N_14757,N_11798,N_10246);
nor U14758 (N_14758,N_10777,N_11750);
nand U14759 (N_14759,N_10672,N_12015);
xor U14760 (N_14760,N_10892,N_10432);
xor U14761 (N_14761,N_11787,N_12147);
and U14762 (N_14762,N_10182,N_12464);
nor U14763 (N_14763,N_10198,N_12460);
and U14764 (N_14764,N_10789,N_10819);
and U14765 (N_14765,N_11155,N_11860);
and U14766 (N_14766,N_11729,N_12123);
nand U14767 (N_14767,N_11194,N_10285);
and U14768 (N_14768,N_10090,N_10275);
xnor U14769 (N_14769,N_10080,N_10677);
xnor U14770 (N_14770,N_11689,N_10728);
or U14771 (N_14771,N_11467,N_11799);
and U14772 (N_14772,N_11725,N_10806);
nor U14773 (N_14773,N_12205,N_11700);
nand U14774 (N_14774,N_10817,N_10146);
nor U14775 (N_14775,N_10379,N_12324);
and U14776 (N_14776,N_11520,N_12480);
or U14777 (N_14777,N_10852,N_10268);
or U14778 (N_14778,N_10926,N_11653);
and U14779 (N_14779,N_10205,N_12439);
nor U14780 (N_14780,N_12165,N_10800);
or U14781 (N_14781,N_10848,N_10333);
or U14782 (N_14782,N_10559,N_11433);
nand U14783 (N_14783,N_12289,N_12311);
nand U14784 (N_14784,N_10857,N_12090);
or U14785 (N_14785,N_11635,N_11715);
or U14786 (N_14786,N_10032,N_10014);
xnor U14787 (N_14787,N_10952,N_12169);
xor U14788 (N_14788,N_12378,N_10562);
and U14789 (N_14789,N_12215,N_11652);
nand U14790 (N_14790,N_10900,N_11256);
and U14791 (N_14791,N_10003,N_10985);
xnor U14792 (N_14792,N_10488,N_11664);
nor U14793 (N_14793,N_11894,N_11223);
or U14794 (N_14794,N_11393,N_11093);
xor U14795 (N_14795,N_11595,N_10811);
xnor U14796 (N_14796,N_10747,N_10716);
xnor U14797 (N_14797,N_11243,N_10462);
nor U14798 (N_14798,N_10978,N_10592);
or U14799 (N_14799,N_10941,N_11034);
xor U14800 (N_14800,N_12424,N_10769);
nor U14801 (N_14801,N_11974,N_11883);
and U14802 (N_14802,N_10906,N_10047);
nand U14803 (N_14803,N_11616,N_11843);
nand U14804 (N_14804,N_10753,N_12182);
nor U14805 (N_14805,N_11639,N_11233);
nand U14806 (N_14806,N_11805,N_10261);
xnor U14807 (N_14807,N_11122,N_10588);
nand U14808 (N_14808,N_10659,N_10435);
nand U14809 (N_14809,N_10402,N_10340);
nand U14810 (N_14810,N_10044,N_11858);
xor U14811 (N_14811,N_11106,N_12271);
and U14812 (N_14812,N_10830,N_10535);
and U14813 (N_14813,N_10568,N_10987);
and U14814 (N_14814,N_10065,N_11633);
and U14815 (N_14815,N_10723,N_12324);
or U14816 (N_14816,N_10179,N_10050);
nor U14817 (N_14817,N_12488,N_11652);
and U14818 (N_14818,N_12126,N_11928);
xnor U14819 (N_14819,N_11323,N_11862);
and U14820 (N_14820,N_11249,N_10091);
and U14821 (N_14821,N_11263,N_10050);
and U14822 (N_14822,N_12428,N_10535);
or U14823 (N_14823,N_12067,N_10345);
xnor U14824 (N_14824,N_10816,N_11995);
xnor U14825 (N_14825,N_11217,N_12487);
or U14826 (N_14826,N_10414,N_12342);
and U14827 (N_14827,N_11717,N_10514);
nand U14828 (N_14828,N_11072,N_10863);
and U14829 (N_14829,N_12138,N_11006);
xnor U14830 (N_14830,N_11444,N_11157);
and U14831 (N_14831,N_10039,N_11373);
xor U14832 (N_14832,N_10375,N_11390);
nor U14833 (N_14833,N_11896,N_11755);
nor U14834 (N_14834,N_10579,N_12309);
and U14835 (N_14835,N_10721,N_12122);
or U14836 (N_14836,N_10034,N_10897);
nand U14837 (N_14837,N_11797,N_10859);
xor U14838 (N_14838,N_10544,N_12213);
nor U14839 (N_14839,N_11665,N_10077);
xnor U14840 (N_14840,N_11176,N_10922);
or U14841 (N_14841,N_10832,N_10525);
nor U14842 (N_14842,N_10236,N_10944);
or U14843 (N_14843,N_11959,N_10856);
and U14844 (N_14844,N_12347,N_11663);
or U14845 (N_14845,N_11097,N_11266);
xor U14846 (N_14846,N_11411,N_10194);
or U14847 (N_14847,N_12401,N_10627);
nand U14848 (N_14848,N_11457,N_12284);
or U14849 (N_14849,N_12286,N_12186);
nand U14850 (N_14850,N_11324,N_11166);
xor U14851 (N_14851,N_10564,N_12228);
xnor U14852 (N_14852,N_10309,N_11697);
or U14853 (N_14853,N_11767,N_12391);
xnor U14854 (N_14854,N_10842,N_11323);
nand U14855 (N_14855,N_11341,N_10590);
nor U14856 (N_14856,N_11254,N_11412);
nor U14857 (N_14857,N_10387,N_11070);
xnor U14858 (N_14858,N_11465,N_11708);
or U14859 (N_14859,N_11406,N_12351);
or U14860 (N_14860,N_11293,N_10151);
xor U14861 (N_14861,N_11170,N_12389);
and U14862 (N_14862,N_11673,N_10687);
or U14863 (N_14863,N_11042,N_11795);
nor U14864 (N_14864,N_12459,N_10943);
nor U14865 (N_14865,N_10488,N_11897);
nand U14866 (N_14866,N_12276,N_11578);
nor U14867 (N_14867,N_11820,N_12250);
nor U14868 (N_14868,N_10067,N_11782);
or U14869 (N_14869,N_11228,N_10409);
or U14870 (N_14870,N_10505,N_11101);
and U14871 (N_14871,N_11446,N_10987);
or U14872 (N_14872,N_11045,N_11673);
xor U14873 (N_14873,N_10733,N_10857);
and U14874 (N_14874,N_10153,N_11754);
xnor U14875 (N_14875,N_10834,N_12134);
nor U14876 (N_14876,N_12207,N_10710);
and U14877 (N_14877,N_10403,N_11704);
nor U14878 (N_14878,N_11715,N_12437);
nor U14879 (N_14879,N_12459,N_10893);
xnor U14880 (N_14880,N_10039,N_11827);
or U14881 (N_14881,N_12370,N_11409);
or U14882 (N_14882,N_10366,N_11253);
or U14883 (N_14883,N_11251,N_10590);
or U14884 (N_14884,N_12499,N_11779);
xnor U14885 (N_14885,N_10315,N_11105);
or U14886 (N_14886,N_10676,N_12423);
or U14887 (N_14887,N_11568,N_10120);
xnor U14888 (N_14888,N_11546,N_11108);
xnor U14889 (N_14889,N_11082,N_12439);
nor U14890 (N_14890,N_10065,N_12480);
xnor U14891 (N_14891,N_10642,N_11552);
xnor U14892 (N_14892,N_12390,N_10489);
nand U14893 (N_14893,N_10830,N_11779);
and U14894 (N_14894,N_10580,N_11059);
xor U14895 (N_14895,N_10841,N_12034);
or U14896 (N_14896,N_12227,N_11416);
nor U14897 (N_14897,N_10950,N_11530);
and U14898 (N_14898,N_10621,N_10981);
xor U14899 (N_14899,N_11235,N_10472);
nor U14900 (N_14900,N_11308,N_10681);
nor U14901 (N_14901,N_10614,N_10534);
nor U14902 (N_14902,N_11926,N_11647);
and U14903 (N_14903,N_10241,N_11976);
or U14904 (N_14904,N_10756,N_10285);
or U14905 (N_14905,N_10255,N_10659);
nand U14906 (N_14906,N_12198,N_10697);
xnor U14907 (N_14907,N_10063,N_11892);
or U14908 (N_14908,N_11050,N_10409);
xnor U14909 (N_14909,N_11339,N_11221);
nand U14910 (N_14910,N_10280,N_10066);
or U14911 (N_14911,N_11646,N_11547);
or U14912 (N_14912,N_11392,N_10338);
nor U14913 (N_14913,N_11746,N_12438);
xnor U14914 (N_14914,N_12304,N_10789);
xnor U14915 (N_14915,N_10678,N_10199);
xnor U14916 (N_14916,N_10017,N_12421);
and U14917 (N_14917,N_11837,N_10037);
and U14918 (N_14918,N_10805,N_11269);
nand U14919 (N_14919,N_10305,N_10745);
nand U14920 (N_14920,N_11675,N_11778);
nand U14921 (N_14921,N_10171,N_11891);
nor U14922 (N_14922,N_10675,N_11367);
or U14923 (N_14923,N_10625,N_12229);
xor U14924 (N_14924,N_12336,N_12189);
or U14925 (N_14925,N_11539,N_12499);
or U14926 (N_14926,N_11554,N_12355);
nand U14927 (N_14927,N_12311,N_11719);
xnor U14928 (N_14928,N_11003,N_10086);
or U14929 (N_14929,N_12140,N_12458);
or U14930 (N_14930,N_12412,N_10004);
and U14931 (N_14931,N_11942,N_11352);
nor U14932 (N_14932,N_11171,N_11508);
xor U14933 (N_14933,N_10478,N_11812);
or U14934 (N_14934,N_10439,N_10070);
xnor U14935 (N_14935,N_11424,N_11330);
and U14936 (N_14936,N_11513,N_11341);
nor U14937 (N_14937,N_11219,N_10996);
xnor U14938 (N_14938,N_11866,N_11256);
and U14939 (N_14939,N_10575,N_10297);
nand U14940 (N_14940,N_10296,N_10086);
or U14941 (N_14941,N_10759,N_11275);
nor U14942 (N_14942,N_10211,N_11264);
xnor U14943 (N_14943,N_11623,N_12014);
nor U14944 (N_14944,N_10934,N_12448);
and U14945 (N_14945,N_10330,N_10156);
or U14946 (N_14946,N_10177,N_12449);
or U14947 (N_14947,N_10707,N_11755);
nand U14948 (N_14948,N_11666,N_11910);
xor U14949 (N_14949,N_11466,N_12052);
or U14950 (N_14950,N_10592,N_12430);
xor U14951 (N_14951,N_10634,N_10576);
nand U14952 (N_14952,N_10913,N_11642);
or U14953 (N_14953,N_10596,N_11654);
or U14954 (N_14954,N_10933,N_10787);
xnor U14955 (N_14955,N_10593,N_11315);
xor U14956 (N_14956,N_11435,N_11207);
xor U14957 (N_14957,N_11732,N_11077);
or U14958 (N_14958,N_12360,N_11619);
xnor U14959 (N_14959,N_11998,N_12047);
nand U14960 (N_14960,N_11037,N_11761);
xnor U14961 (N_14961,N_11257,N_11662);
and U14962 (N_14962,N_10176,N_10140);
and U14963 (N_14963,N_12232,N_10778);
nor U14964 (N_14964,N_10038,N_10620);
and U14965 (N_14965,N_10750,N_11650);
or U14966 (N_14966,N_11985,N_11698);
nand U14967 (N_14967,N_10588,N_10276);
xor U14968 (N_14968,N_11907,N_10486);
or U14969 (N_14969,N_10146,N_12135);
or U14970 (N_14970,N_10691,N_10821);
or U14971 (N_14971,N_10969,N_12335);
nand U14972 (N_14972,N_10222,N_11368);
or U14973 (N_14973,N_10276,N_11310);
or U14974 (N_14974,N_12458,N_11004);
and U14975 (N_14975,N_11382,N_10914);
or U14976 (N_14976,N_11198,N_11631);
and U14977 (N_14977,N_11837,N_11277);
xnor U14978 (N_14978,N_11592,N_12247);
nor U14979 (N_14979,N_10060,N_11607);
or U14980 (N_14980,N_10105,N_10700);
or U14981 (N_14981,N_11000,N_11545);
nor U14982 (N_14982,N_11698,N_10597);
and U14983 (N_14983,N_10570,N_11980);
nand U14984 (N_14984,N_11475,N_11582);
nand U14985 (N_14985,N_11598,N_10782);
nor U14986 (N_14986,N_12417,N_10132);
nand U14987 (N_14987,N_12257,N_10976);
nand U14988 (N_14988,N_11154,N_11370);
or U14989 (N_14989,N_11957,N_11099);
nand U14990 (N_14990,N_11492,N_10147);
xor U14991 (N_14991,N_12461,N_12493);
and U14992 (N_14992,N_10725,N_11674);
and U14993 (N_14993,N_12429,N_10662);
or U14994 (N_14994,N_11067,N_12202);
nand U14995 (N_14995,N_10203,N_11336);
and U14996 (N_14996,N_11810,N_10210);
xor U14997 (N_14997,N_10012,N_11593);
and U14998 (N_14998,N_12406,N_10385);
and U14999 (N_14999,N_10826,N_12045);
or U15000 (N_15000,N_14891,N_12518);
and U15001 (N_15001,N_14825,N_13397);
and U15002 (N_15002,N_13529,N_14782);
xor U15003 (N_15003,N_14513,N_14717);
xnor U15004 (N_15004,N_12529,N_13146);
xnor U15005 (N_15005,N_14029,N_13619);
xnor U15006 (N_15006,N_12698,N_12702);
or U15007 (N_15007,N_14224,N_14548);
nor U15008 (N_15008,N_14003,N_12586);
nor U15009 (N_15009,N_14150,N_13066);
nand U15010 (N_15010,N_13392,N_13271);
nor U15011 (N_15011,N_13368,N_14960);
xnor U15012 (N_15012,N_13039,N_14039);
and U15013 (N_15013,N_14893,N_13701);
nand U15014 (N_15014,N_14794,N_14523);
nor U15015 (N_15015,N_13280,N_13053);
nor U15016 (N_15016,N_13449,N_14242);
and U15017 (N_15017,N_14652,N_13434);
nand U15018 (N_15018,N_14524,N_13415);
nor U15019 (N_15019,N_14184,N_13616);
or U15020 (N_15020,N_14379,N_14958);
and U15021 (N_15021,N_12973,N_12956);
nor U15022 (N_15022,N_13906,N_12836);
and U15023 (N_15023,N_12990,N_13017);
or U15024 (N_15024,N_12631,N_12553);
nand U15025 (N_15025,N_14102,N_14462);
and U15026 (N_15026,N_14816,N_14533);
or U15027 (N_15027,N_14896,N_13383);
xor U15028 (N_15028,N_14270,N_14147);
nor U15029 (N_15029,N_12985,N_13268);
xor U15030 (N_15030,N_14457,N_12515);
nand U15031 (N_15031,N_13834,N_13676);
xnor U15032 (N_15032,N_14736,N_13174);
or U15033 (N_15033,N_12654,N_13236);
xor U15034 (N_15034,N_13102,N_12732);
nand U15035 (N_15035,N_14112,N_13260);
and U15036 (N_15036,N_14752,N_13806);
nor U15037 (N_15037,N_14624,N_12886);
xnor U15038 (N_15038,N_14635,N_13962);
and U15039 (N_15039,N_13876,N_14632);
xor U15040 (N_15040,N_12940,N_13028);
or U15041 (N_15041,N_14257,N_12652);
nand U15042 (N_15042,N_14655,N_14601);
nand U15043 (N_15043,N_13703,N_14053);
and U15044 (N_15044,N_13391,N_13508);
nand U15045 (N_15045,N_13851,N_14784);
xnor U15046 (N_15046,N_14827,N_13231);
and U15047 (N_15047,N_13126,N_14708);
nand U15048 (N_15048,N_13172,N_13615);
xor U15049 (N_15049,N_13599,N_12582);
nand U15050 (N_15050,N_14515,N_14249);
or U15051 (N_15051,N_12658,N_13071);
and U15052 (N_15052,N_13119,N_14895);
or U15053 (N_15053,N_12934,N_13805);
and U15054 (N_15054,N_12954,N_12630);
nor U15055 (N_15055,N_14351,N_13495);
nor U15056 (N_15056,N_13474,N_14144);
and U15057 (N_15057,N_14110,N_12651);
nand U15058 (N_15058,N_12982,N_13341);
nand U15059 (N_15059,N_14553,N_13413);
and U15060 (N_15060,N_13734,N_13334);
xor U15061 (N_15061,N_13914,N_13904);
and U15062 (N_15062,N_13414,N_13762);
or U15063 (N_15063,N_13234,N_13627);
nor U15064 (N_15064,N_13848,N_12864);
nor U15065 (N_15065,N_14436,N_14483);
or U15066 (N_15066,N_12599,N_13836);
and U15067 (N_15067,N_13041,N_13117);
nand U15068 (N_15068,N_13357,N_13927);
xnor U15069 (N_15069,N_12689,N_12547);
and U15070 (N_15070,N_13749,N_13583);
and U15071 (N_15071,N_13592,N_13249);
nand U15072 (N_15072,N_14921,N_14686);
xnor U15073 (N_15073,N_12841,N_14608);
and U15074 (N_15074,N_14231,N_13623);
or U15075 (N_15075,N_13165,N_14022);
or U15076 (N_15076,N_14616,N_13277);
or U15077 (N_15077,N_14016,N_14550);
and U15078 (N_15078,N_13575,N_13767);
xnor U15079 (N_15079,N_14063,N_14567);
nor U15080 (N_15080,N_14541,N_13170);
and U15081 (N_15081,N_14157,N_14341);
nand U15082 (N_15082,N_13689,N_13861);
nor U15083 (N_15083,N_14335,N_14946);
xor U15084 (N_15084,N_12895,N_14968);
and U15085 (N_15085,N_13006,N_13540);
nor U15086 (N_15086,N_12613,N_13664);
and U15087 (N_15087,N_13224,N_12949);
nor U15088 (N_15088,N_13284,N_13443);
and U15089 (N_15089,N_14178,N_13079);
nand U15090 (N_15090,N_14589,N_13845);
or U15091 (N_15091,N_14132,N_13240);
nor U15092 (N_15092,N_12984,N_14729);
nor U15093 (N_15093,N_13296,N_12745);
and U15094 (N_15094,N_13156,N_13572);
xor U15095 (N_15095,N_12980,N_14767);
and U15096 (N_15096,N_14870,N_14631);
nor U15097 (N_15097,N_13469,N_14555);
or U15098 (N_15098,N_12693,N_13010);
xnor U15099 (N_15099,N_12675,N_14491);
xnor U15100 (N_15100,N_12873,N_12624);
and U15101 (N_15101,N_12533,N_13747);
nor U15102 (N_15102,N_12541,N_14644);
xnor U15103 (N_15103,N_14252,N_13486);
or U15104 (N_15104,N_13441,N_14780);
xnor U15105 (N_15105,N_14793,N_14975);
nor U15106 (N_15106,N_14439,N_14807);
nor U15107 (N_15107,N_13931,N_12998);
xnor U15108 (N_15108,N_14050,N_12816);
and U15109 (N_15109,N_13150,N_12749);
and U15110 (N_15110,N_13223,N_13919);
xnor U15111 (N_15111,N_13106,N_12712);
nand U15112 (N_15112,N_13728,N_14255);
and U15113 (N_15113,N_13332,N_13645);
nand U15114 (N_15114,N_14872,N_12629);
nand U15115 (N_15115,N_13807,N_14206);
or U15116 (N_15116,N_14540,N_14714);
and U15117 (N_15117,N_13889,N_12728);
and U15118 (N_15118,N_14750,N_14187);
or U15119 (N_15119,N_14017,N_14596);
nand U15120 (N_15120,N_13633,N_14938);
nor U15121 (N_15121,N_14098,N_13109);
and U15122 (N_15122,N_13325,N_13941);
nor U15123 (N_15123,N_13754,N_13976);
and U15124 (N_15124,N_13909,N_14575);
and U15125 (N_15125,N_13573,N_13359);
and U15126 (N_15126,N_13131,N_13228);
xnor U15127 (N_15127,N_14398,N_13366);
and U15128 (N_15128,N_13644,N_14674);
and U15129 (N_15129,N_14700,N_13499);
and U15130 (N_15130,N_13925,N_14223);
xnor U15131 (N_15131,N_14311,N_13061);
nand U15132 (N_15132,N_13120,N_13207);
nand U15133 (N_15133,N_13995,N_13149);
or U15134 (N_15134,N_14478,N_13245);
xnor U15135 (N_15135,N_12759,N_13830);
and U15136 (N_15136,N_12594,N_13542);
nor U15137 (N_15137,N_13446,N_13381);
nor U15138 (N_15138,N_12707,N_13569);
nand U15139 (N_15139,N_14226,N_13517);
nand U15140 (N_15140,N_14662,N_12771);
and U15141 (N_15141,N_12604,N_14578);
nand U15142 (N_15142,N_13980,N_13233);
xor U15143 (N_15143,N_14072,N_12569);
xnor U15144 (N_15144,N_14585,N_13140);
nor U15145 (N_15145,N_14289,N_14582);
and U15146 (N_15146,N_14977,N_13211);
nor U15147 (N_15147,N_13698,N_14762);
and U15148 (N_15148,N_14395,N_14389);
nand U15149 (N_15149,N_14306,N_14120);
xnor U15150 (N_15150,N_13872,N_13226);
and U15151 (N_15151,N_13369,N_12825);
and U15152 (N_15152,N_14724,N_13626);
nand U15153 (N_15153,N_13266,N_12963);
nor U15154 (N_15154,N_13541,N_14962);
nand U15155 (N_15155,N_14472,N_14739);
or U15156 (N_15156,N_14667,N_13073);
and U15157 (N_15157,N_13304,N_13781);
nor U15158 (N_15158,N_13099,N_12791);
or U15159 (N_15159,N_12930,N_12952);
or U15160 (N_15160,N_13076,N_13206);
or U15161 (N_15161,N_12860,N_12892);
nand U15162 (N_15162,N_14416,N_14365);
nor U15163 (N_15163,N_13029,N_14012);
xor U15164 (N_15164,N_14262,N_12716);
and U15165 (N_15165,N_13780,N_13898);
xor U15166 (N_15166,N_13450,N_14054);
nor U15167 (N_15167,N_13351,N_13046);
nor U15168 (N_15168,N_13487,N_14526);
and U15169 (N_15169,N_14275,N_13994);
xnor U15170 (N_15170,N_14103,N_14878);
or U15171 (N_15171,N_13072,N_12968);
or U15172 (N_15172,N_14285,N_13860);
nor U15173 (N_15173,N_13605,N_14598);
nand U15174 (N_15174,N_13204,N_14430);
xnor U15175 (N_15175,N_14067,N_14511);
nor U15176 (N_15176,N_13763,N_14517);
and U15177 (N_15177,N_12750,N_14431);
nor U15178 (N_15178,N_14479,N_14902);
or U15179 (N_15179,N_14497,N_14857);
nand U15180 (N_15180,N_12876,N_13320);
or U15181 (N_15181,N_14682,N_13850);
and U15182 (N_15182,N_13247,N_13577);
nor U15183 (N_15183,N_12919,N_13180);
xnor U15184 (N_15184,N_12875,N_14786);
xnor U15185 (N_15185,N_14888,N_14591);
xor U15186 (N_15186,N_14373,N_13404);
or U15187 (N_15187,N_13500,N_13510);
nor U15188 (N_15188,N_12822,N_13534);
xnor U15189 (N_15189,N_14864,N_12986);
and U15190 (N_15190,N_12953,N_13839);
or U15191 (N_15191,N_14688,N_14507);
nor U15192 (N_15192,N_14485,N_14279);
nor U15193 (N_15193,N_14444,N_13853);
or U15194 (N_15194,N_13974,N_14121);
nand U15195 (N_15195,N_14159,N_13518);
nand U15196 (N_15196,N_14399,N_14097);
and U15197 (N_15197,N_13330,N_12598);
or U15198 (N_15198,N_14111,N_13936);
xor U15199 (N_15199,N_14302,N_14445);
nor U15200 (N_15200,N_14592,N_13103);
xor U15201 (N_15201,N_12969,N_14455);
nor U15202 (N_15202,N_14496,N_13602);
and U15203 (N_15203,N_13630,N_14031);
xnor U15204 (N_15204,N_14980,N_14355);
xor U15205 (N_15205,N_14613,N_13164);
nor U15206 (N_15206,N_13917,N_14030);
nand U15207 (N_15207,N_14402,N_14267);
nand U15208 (N_15208,N_12787,N_13586);
nand U15209 (N_15209,N_13580,N_13353);
nand U15210 (N_15210,N_14787,N_12572);
or U15211 (N_15211,N_14703,N_14331);
xor U15212 (N_15212,N_12931,N_13018);
nor U15213 (N_15213,N_13888,N_14074);
or U15214 (N_15214,N_14238,N_14182);
or U15215 (N_15215,N_12843,N_14308);
nor U15216 (N_15216,N_12577,N_14475);
and U15217 (N_15217,N_13873,N_13560);
or U15218 (N_15218,N_14099,N_12850);
nor U15219 (N_15219,N_13212,N_12877);
or U15220 (N_15220,N_13826,N_14435);
or U15221 (N_15221,N_13915,N_14446);
and U15222 (N_15222,N_13827,N_13321);
or U15223 (N_15223,N_14059,N_12726);
or U15224 (N_15224,N_14846,N_13455);
xnor U15225 (N_15225,N_14163,N_13355);
and U15226 (N_15226,N_14656,N_12605);
nor U15227 (N_15227,N_13907,N_12844);
xor U15228 (N_15228,N_14153,N_13646);
and U15229 (N_15229,N_14188,N_13857);
nand U15230 (N_15230,N_12817,N_12643);
nor U15231 (N_15231,N_12751,N_13312);
nand U15232 (N_15232,N_13399,N_12508);
nor U15233 (N_15233,N_14149,N_12758);
and U15234 (N_15234,N_14284,N_13802);
nor U15235 (N_15235,N_13891,N_14010);
or U15236 (N_15236,N_14551,N_14327);
nor U15237 (N_15237,N_14698,N_14769);
xnor U15238 (N_15238,N_12829,N_13821);
nor U15239 (N_15239,N_14143,N_13407);
nand U15240 (N_15240,N_12893,N_14917);
or U15241 (N_15241,N_14114,N_12616);
nand U15242 (N_15242,N_13971,N_14338);
nand U15243 (N_15243,N_12609,N_14384);
nand U15244 (N_15244,N_12555,N_13622);
or U15245 (N_15245,N_12708,N_13112);
xnor U15246 (N_15246,N_13253,N_14244);
nand U15247 (N_15247,N_13856,N_12789);
nand U15248 (N_15248,N_14773,N_12858);
and U15249 (N_15249,N_13568,N_14577);
or U15250 (N_15250,N_14826,N_14198);
nand U15251 (N_15251,N_14563,N_12857);
and U15252 (N_15252,N_14790,N_14746);
nor U15253 (N_15253,N_12951,N_14874);
xor U15254 (N_15254,N_12838,N_13267);
xor U15255 (N_15255,N_14428,N_14981);
or U15256 (N_15256,N_12746,N_13611);
or U15257 (N_15257,N_14948,N_14957);
or U15258 (N_15258,N_12792,N_13905);
and U15259 (N_15259,N_13513,N_14650);
nand U15260 (N_15260,N_13973,N_13711);
or U15261 (N_15261,N_14680,N_12946);
nor U15262 (N_15262,N_14026,N_14564);
and U15263 (N_15263,N_13649,N_13547);
nor U15264 (N_15264,N_14926,N_13471);
nand U15265 (N_15265,N_12706,N_14875);
xor U15266 (N_15266,N_13181,N_14015);
or U15267 (N_15267,N_14869,N_13757);
nand U15268 (N_15268,N_14818,N_14276);
or U15269 (N_15269,N_14057,N_14712);
nor U15270 (N_15270,N_13273,N_13512);
or U15271 (N_15271,N_12589,N_14303);
nand U15272 (N_15272,N_12863,N_13804);
and U15273 (N_15273,N_14629,N_12507);
or U15274 (N_15274,N_14751,N_14309);
xor U15275 (N_15275,N_13666,N_13101);
nand U15276 (N_15276,N_14393,N_12575);
nor U15277 (N_15277,N_14861,N_13854);
nor U15278 (N_15278,N_13721,N_13171);
nor U15279 (N_15279,N_14219,N_14670);
xor U15280 (N_15280,N_12635,N_13582);
nor U15281 (N_15281,N_14673,N_12981);
xor U15282 (N_15282,N_13688,N_14953);
or U15283 (N_15283,N_13758,N_14810);
or U15284 (N_15284,N_14142,N_13459);
or U15285 (N_15285,N_13186,N_13288);
xnor U15286 (N_15286,N_12724,N_12775);
nor U15287 (N_15287,N_13022,N_12818);
nor U15288 (N_15288,N_14944,N_13343);
nand U15289 (N_15289,N_13870,N_14477);
nor U15290 (N_15290,N_14868,N_13691);
nand U15291 (N_15291,N_13261,N_12692);
or U15292 (N_15292,N_13539,N_12853);
nor U15293 (N_15293,N_13981,N_12512);
or U15294 (N_15294,N_13335,N_13048);
nand U15295 (N_15295,N_12747,N_12677);
and U15296 (N_15296,N_14612,N_13057);
nand U15297 (N_15297,N_13803,N_14676);
nand U15298 (N_15298,N_12719,N_14900);
xnor U15299 (N_15299,N_14155,N_13151);
xnor U15300 (N_15300,N_13667,N_14630);
or U15301 (N_15301,N_14521,N_14593);
nand U15302 (N_15302,N_12754,N_13902);
nand U15303 (N_15303,N_13983,N_14177);
xnor U15304 (N_15304,N_14576,N_13173);
nor U15305 (N_15305,N_13571,N_14572);
nor U15306 (N_15306,N_13935,N_14065);
nand U15307 (N_15307,N_14903,N_14726);
nand U15308 (N_15308,N_13822,N_13933);
xor U15309 (N_15309,N_13525,N_12686);
nor U15310 (N_15310,N_14509,N_12717);
and U15311 (N_15311,N_13141,N_13522);
nand U15312 (N_15312,N_14976,N_12606);
xnor U15313 (N_15313,N_12567,N_14222);
or U15314 (N_15314,N_14469,N_14693);
and U15315 (N_15315,N_14738,N_13593);
or U15316 (N_15316,N_13669,N_12861);
and U15317 (N_15317,N_13093,N_13373);
nor U15318 (N_15318,N_14210,N_13384);
xor U15319 (N_15319,N_14452,N_12912);
xor U15320 (N_15320,N_13563,N_14518);
and U15321 (N_15321,N_13910,N_12849);
xnor U15322 (N_15322,N_14245,N_14218);
nor U15323 (N_15323,N_13968,N_14374);
xor U15324 (N_15324,N_13685,N_14089);
xnor U15325 (N_15325,N_14552,N_13238);
and U15326 (N_15326,N_13454,N_14606);
or U15327 (N_15327,N_14221,N_12997);
nor U15328 (N_15328,N_13793,N_14328);
or U15329 (N_15329,N_13085,N_12942);
xnor U15330 (N_15330,N_13221,N_13144);
nand U15331 (N_15331,N_14522,N_13027);
or U15332 (N_15332,N_12902,N_14332);
and U15333 (N_15333,N_13175,N_13531);
xnor U15334 (N_15334,N_12568,N_14898);
nor U15335 (N_15335,N_13641,N_13768);
or U15336 (N_15336,N_14002,N_14964);
nand U15337 (N_15337,N_12960,N_14979);
or U15338 (N_15338,N_13059,N_14091);
or U15339 (N_15339,N_12500,N_13423);
nor U15340 (N_15340,N_12640,N_12506);
and U15341 (N_15341,N_12774,N_13394);
nor U15342 (N_15342,N_13695,N_14843);
nor U15343 (N_15343,N_13969,N_13421);
nor U15344 (N_15344,N_13254,N_14080);
xnor U15345 (N_15345,N_14607,N_14663);
or U15346 (N_15346,N_13672,N_14025);
or U15347 (N_15347,N_12896,N_13752);
and U15348 (N_15348,N_13772,N_13301);
or U15349 (N_15349,N_14645,N_13289);
xnor U15350 (N_15350,N_14194,N_14354);
or U15351 (N_15351,N_13647,N_13938);
nand U15352 (N_15352,N_14183,N_14077);
or U15353 (N_15353,N_14251,N_13723);
or U15354 (N_15354,N_13852,N_13246);
nand U15355 (N_15355,N_13589,N_14538);
and U15356 (N_15356,N_14137,N_14036);
xor U15357 (N_15357,N_14201,N_13045);
xnor U15358 (N_15358,N_13142,N_12559);
nand U15359 (N_15359,N_13635,N_13725);
or U15360 (N_15360,N_14855,N_13411);
and U15361 (N_15361,N_12536,N_14488);
nor U15362 (N_15362,N_14919,N_12557);
and U15363 (N_15363,N_13782,N_12727);
nand U15364 (N_15364,N_13581,N_14618);
and U15365 (N_15365,N_13811,N_13696);
and U15366 (N_15366,N_12859,N_14704);
and U15367 (N_15367,N_13502,N_14837);
and U15368 (N_15368,N_12827,N_14281);
and U15369 (N_15369,N_14815,N_13978);
or U15370 (N_15370,N_13730,N_13303);
or U15371 (N_15371,N_13086,N_13556);
nor U15372 (N_15372,N_12539,N_14557);
or U15373 (N_15373,N_12521,N_13435);
and U15374 (N_15374,N_13333,N_13614);
or U15375 (N_15375,N_12538,N_14623);
or U15376 (N_15376,N_14007,N_13796);
and U15377 (N_15377,N_13713,N_12554);
and U15378 (N_15378,N_14191,N_14679);
nand U15379 (N_15379,N_12691,N_13433);
nor U15380 (N_15380,N_13208,N_12979);
xnor U15381 (N_15381,N_14918,N_13197);
xnor U15382 (N_15382,N_14162,N_13179);
nand U15383 (N_15383,N_12528,N_13727);
nor U15384 (N_15384,N_13682,N_13470);
nor U15385 (N_15385,N_14772,N_14675);
and U15386 (N_15386,N_12803,N_14368);
nand U15387 (N_15387,N_14971,N_13339);
nand U15388 (N_15388,N_14443,N_14106);
nor U15389 (N_15389,N_12842,N_12779);
or U15390 (N_15390,N_13153,N_14290);
xor U15391 (N_15391,N_13004,N_13432);
and U15392 (N_15392,N_12770,N_14505);
and U15393 (N_15393,N_14427,N_14955);
nand U15394 (N_15394,N_13760,N_13417);
nand U15395 (N_15395,N_14997,N_13008);
nand U15396 (N_15396,N_12773,N_14310);
or U15397 (N_15397,N_14535,N_13604);
and U15398 (N_15398,N_13504,N_13143);
nand U15399 (N_15399,N_14824,N_14292);
and U15400 (N_15400,N_13610,N_13298);
or U15401 (N_15401,N_13188,N_14580);
xnor U15402 (N_15402,N_14045,N_14766);
xor U15403 (N_15403,N_13503,N_14135);
or U15404 (N_15404,N_14940,N_13490);
nor U15405 (N_15405,N_14021,N_13920);
and U15406 (N_15406,N_13396,N_14614);
and U15407 (N_15407,N_14910,N_13452);
xor U15408 (N_15408,N_14009,N_14569);
xor U15409 (N_15409,N_13609,N_14419);
or U15410 (N_15410,N_14889,N_14125);
nor U15411 (N_15411,N_12757,N_13951);
xor U15412 (N_15412,N_12656,N_14081);
xnor U15413 (N_15413,N_13596,N_14839);
xor U15414 (N_15414,N_12871,N_14634);
and U15415 (N_15415,N_14972,N_13833);
nor U15416 (N_15416,N_12748,N_14378);
nand U15417 (N_15417,N_12525,N_13631);
or U15418 (N_15418,N_14988,N_13629);
xnor U15419 (N_15419,N_14295,N_14096);
nor U15420 (N_15420,N_12905,N_14247);
or U15421 (N_15421,N_14024,N_12617);
or U15422 (N_15422,N_12709,N_12994);
nor U15423 (N_15423,N_14808,N_12962);
nand U15424 (N_15424,N_13402,N_13838);
or U15425 (N_15425,N_14792,N_13892);
nand U15426 (N_15426,N_13603,N_12904);
xnor U15427 (N_15427,N_13511,N_14494);
nand U15428 (N_15428,N_13939,N_13986);
xnor U15429 (N_15429,N_14265,N_13007);
or U15430 (N_15430,N_13350,N_13679);
or U15431 (N_15431,N_13779,N_14118);
or U15432 (N_15432,N_14042,N_14851);
xnor U15433 (N_15433,N_14728,N_13177);
xor U15434 (N_15434,N_14300,N_12882);
or U15435 (N_15435,N_12696,N_12657);
and U15436 (N_15436,N_14361,N_14881);
or U15437 (N_15437,N_14761,N_14266);
and U15438 (N_15438,N_13192,N_13044);
nor U15439 (N_15439,N_13792,N_12808);
nand U15440 (N_15440,N_13913,N_12522);
nor U15441 (N_15441,N_13315,N_12958);
xnor U15442 (N_15442,N_12523,N_14146);
nor U15443 (N_15443,N_13795,N_14508);
and U15444 (N_15444,N_13726,N_12936);
and U15445 (N_15445,N_13160,N_13408);
nand U15446 (N_15446,N_14196,N_13998);
nor U15447 (N_15447,N_14038,N_14033);
xor U15448 (N_15448,N_13567,N_14941);
and U15449 (N_15449,N_13673,N_13750);
nor U15450 (N_15450,N_13942,N_13736);
or U15451 (N_15451,N_13544,N_14537);
and U15452 (N_15452,N_14706,N_14858);
xnor U15453 (N_15453,N_12637,N_14967);
or U15454 (N_15454,N_12744,N_13447);
xor U15455 (N_15455,N_12831,N_13038);
and U15456 (N_15456,N_14417,N_13965);
and U15457 (N_15457,N_13482,N_12510);
xnor U15458 (N_15458,N_13809,N_13922);
xor U15459 (N_15459,N_14418,N_14415);
nand U15460 (N_15460,N_14713,N_14109);
or U15461 (N_15461,N_13466,N_14811);
nor U15462 (N_15462,N_13576,N_13895);
xnor U15463 (N_15463,N_12741,N_14768);
xor U15464 (N_15464,N_13241,N_12502);
or U15465 (N_15465,N_12671,N_13020);
nor U15466 (N_15466,N_14646,N_12537);
or U15467 (N_15467,N_14179,N_14775);
nand U15468 (N_15468,N_13775,N_13125);
nor U15469 (N_15469,N_14214,N_12763);
and U15470 (N_15470,N_13114,N_14156);
and U15471 (N_15471,N_14558,N_14107);
nand U15472 (N_15472,N_12846,N_13379);
nand U15473 (N_15473,N_13054,N_13637);
xnor U15474 (N_15474,N_13710,N_14689);
nand U15475 (N_15475,N_12782,N_13157);
nor U15476 (N_15476,N_14885,N_14441);
or U15477 (N_15477,N_13347,N_12784);
xnor U15478 (N_15478,N_12901,N_14539);
nor U15479 (N_15479,N_14754,N_14930);
nor U15480 (N_15480,N_14573,N_14165);
and U15481 (N_15481,N_14731,N_13444);
nor U15482 (N_15482,N_12649,N_13702);
xnor U15483 (N_15483,N_13650,N_13538);
nor U15484 (N_15484,N_14833,N_14649);
nor U15485 (N_15485,N_12802,N_13185);
nor U15486 (N_15486,N_13476,N_14315);
nand U15487 (N_15487,N_12993,N_12591);
xnor U15488 (N_15488,N_13235,N_13047);
and U15489 (N_15489,N_14641,N_12628);
and U15490 (N_15490,N_14264,N_14943);
nor U15491 (N_15491,N_13816,N_13243);
nand U15492 (N_15492,N_14041,N_14161);
nand U15493 (N_15493,N_13064,N_13662);
and U15494 (N_15494,N_14745,N_14407);
nor U15495 (N_15495,N_14531,N_14055);
and U15496 (N_15496,N_14248,N_12738);
and U15497 (N_15497,N_12534,N_13201);
nor U15498 (N_15498,N_12928,N_14383);
xor U15499 (N_15499,N_12627,N_14805);
or U15500 (N_15500,N_13712,N_12926);
nand U15501 (N_15501,N_14923,N_13523);
nand U15502 (N_15502,N_14892,N_14282);
xnor U15503 (N_15503,N_13098,N_14806);
or U15504 (N_15504,N_13743,N_13481);
or U15505 (N_15505,N_13422,N_13875);
nand U15506 (N_15506,N_12564,N_13265);
or U15507 (N_15507,N_14721,N_13928);
nor U15508 (N_15508,N_14071,N_13262);
or U15509 (N_15509,N_12639,N_13776);
and U15510 (N_15510,N_13944,N_14758);
nor U15511 (N_15511,N_14287,N_12739);
or U15512 (N_15512,N_14486,N_13708);
and U15513 (N_15513,N_12597,N_14659);
nand U15514 (N_15514,N_13274,N_13216);
nand U15515 (N_15515,N_13532,N_13055);
nand U15516 (N_15516,N_14447,N_12948);
or U15517 (N_15517,N_13570,N_13338);
and U15518 (N_15518,N_12711,N_14740);
or U15519 (N_15519,N_12669,N_13349);
or U15520 (N_15520,N_12959,N_14908);
xnor U15521 (N_15521,N_13348,N_13770);
or U15522 (N_15522,N_12543,N_13656);
nand U15523 (N_15523,N_12713,N_14438);
or U15524 (N_15524,N_14587,N_13787);
xor U15525 (N_15525,N_13410,N_13084);
and U15526 (N_15526,N_13864,N_14711);
nor U15527 (N_15527,N_14985,N_12673);
and U15528 (N_15528,N_14732,N_13279);
and U15529 (N_15529,N_13395,N_13195);
and U15530 (N_15530,N_12937,N_13345);
and U15531 (N_15531,N_14990,N_14253);
and U15532 (N_15532,N_14233,N_14989);
nand U15533 (N_15533,N_13001,N_13880);
or U15534 (N_15534,N_13270,N_14359);
nand U15535 (N_15535,N_13960,N_13285);
or U15536 (N_15536,N_14661,N_14449);
xnor U15537 (N_15537,N_12524,N_12911);
and U15538 (N_15538,N_12851,N_14747);
nor U15539 (N_15539,N_13091,N_12513);
or U15540 (N_15540,N_13884,N_13217);
nand U15541 (N_15541,N_12687,N_12618);
xnor U15542 (N_15542,N_14131,N_13595);
nor U15543 (N_15543,N_14757,N_13999);
nand U15544 (N_15544,N_14894,N_14829);
nor U15545 (N_15545,N_13478,N_14241);
nor U15546 (N_15546,N_14776,N_14742);
xnor U15547 (N_15547,N_13483,N_14709);
nand U15548 (N_15548,N_14566,N_13317);
or U15549 (N_15549,N_12879,N_14258);
and U15550 (N_15550,N_14883,N_14696);
nand U15551 (N_15551,N_13565,N_13600);
and U15552 (N_15552,N_13731,N_13494);
nand U15553 (N_15553,N_12920,N_14489);
and U15554 (N_15554,N_14356,N_13081);
nor U15555 (N_15555,N_13882,N_13566);
or U15556 (N_15556,N_14404,N_14410);
nor U15557 (N_15557,N_14138,N_14340);
xnor U15558 (N_15558,N_14463,N_13653);
xor U15559 (N_15559,N_14350,N_14216);
and U15560 (N_15560,N_12505,N_12663);
xor U15561 (N_15561,N_13309,N_14464);
or U15562 (N_15562,N_14154,N_13943);
xnor U15563 (N_15563,N_13219,N_13137);
xnor U15564 (N_15564,N_14545,N_13606);
and U15565 (N_15565,N_13451,N_12558);
xor U15566 (N_15566,N_12955,N_12610);
and U15567 (N_15567,N_14687,N_14334);
and U15568 (N_15568,N_14301,N_13252);
xor U15569 (N_15569,N_14049,N_12588);
and U15570 (N_15570,N_13766,N_14602);
and U15571 (N_15571,N_13670,N_14396);
and U15572 (N_15572,N_13977,N_14996);
nor U15573 (N_15573,N_13774,N_12753);
xnor U15574 (N_15574,N_13448,N_14158);
nand U15575 (N_15575,N_14305,N_14493);
nand U15576 (N_15576,N_13344,N_14856);
nor U15577 (N_15577,N_12516,N_13945);
and U15578 (N_15578,N_13671,N_13364);
or U15579 (N_15579,N_14619,N_14073);
or U15580 (N_15580,N_12805,N_12603);
or U15581 (N_15581,N_14819,N_12647);
and U15582 (N_15582,N_13390,N_14064);
and U15583 (N_15583,N_14669,N_13899);
nand U15584 (N_15584,N_14809,N_14638);
nand U15585 (N_15585,N_12809,N_13092);
nand U15586 (N_15586,N_12607,N_12927);
or U15587 (N_15587,N_14454,N_12813);
and U15588 (N_15588,N_12593,N_14835);
or U15589 (N_15589,N_12576,N_14841);
and U15590 (N_15590,N_14105,N_12910);
xnor U15591 (N_15591,N_13755,N_12974);
nor U15592 (N_15592,N_12565,N_13578);
nor U15593 (N_15593,N_12560,N_13618);
and U15594 (N_15594,N_12971,N_13958);
and U15595 (N_15595,N_13955,N_13037);
xnor U15596 (N_15596,N_14886,N_14859);
nand U15597 (N_15597,N_14199,N_14705);
and U15598 (N_15598,N_14476,N_12801);
nand U15599 (N_15599,N_14370,N_14764);
nor U15600 (N_15600,N_14160,N_13842);
xor U15601 (N_15601,N_14195,N_14040);
and U15602 (N_15602,N_13431,N_12913);
or U15603 (N_15603,N_13406,N_12583);
or U15604 (N_15604,N_14876,N_13632);
nand U15605 (N_15605,N_12788,N_13621);
and U15606 (N_15606,N_13657,N_13966);
nor U15607 (N_15607,N_13658,N_13783);
nand U15608 (N_15608,N_13916,N_14048);
xor U15609 (N_15609,N_13484,N_12966);
and U15610 (N_15610,N_13700,N_14286);
nand U15611 (N_15611,N_13520,N_14554);
nor U15612 (N_15612,N_13733,N_12991);
nor U15613 (N_15613,N_14205,N_13276);
xnor U15614 (N_15614,N_14200,N_13050);
xor U15615 (N_15615,N_12736,N_14474);
xnor U15616 (N_15616,N_13202,N_14207);
or U15617 (N_15617,N_14128,N_12799);
nor U15618 (N_15618,N_13900,N_13002);
or U15619 (N_15619,N_14375,N_13901);
xor U15620 (N_15620,N_14405,N_13724);
and U15621 (N_15621,N_14083,N_14615);
nor U15622 (N_15622,N_14408,N_14934);
nand U15623 (N_15623,N_14753,N_14610);
nand U15624 (N_15624,N_14314,N_13340);
xnor U15625 (N_15625,N_12950,N_14528);
xnor U15626 (N_15626,N_13051,N_12562);
xor U15627 (N_15627,N_13374,N_13964);
and U15628 (N_15628,N_13294,N_14707);
nor U15629 (N_15629,N_14423,N_13293);
xnor U15630 (N_15630,N_13549,N_12790);
nand U15631 (N_15631,N_13498,N_12566);
nand U15632 (N_15632,N_12570,N_12992);
or U15633 (N_15633,N_14579,N_12581);
or U15634 (N_15634,N_14392,N_13387);
and U15635 (N_15635,N_14914,N_13264);
xor U15636 (N_15636,N_14230,N_13947);
nand U15637 (N_15637,N_14371,N_14832);
and U15638 (N_15638,N_13720,N_14969);
nor U15639 (N_15639,N_13718,N_12661);
or U15640 (N_15640,N_14970,N_13352);
nor U15641 (N_15641,N_13832,N_14326);
nand U15642 (N_15642,N_13810,N_14799);
nor U15643 (N_15643,N_13196,N_13970);
and U15644 (N_15644,N_13295,N_12819);
and U15645 (N_15645,N_14913,N_13021);
nand U15646 (N_15646,N_13287,N_14298);
or U15647 (N_15647,N_13528,N_13985);
or U15648 (N_15648,N_14259,N_14113);
xnor U15649 (N_15649,N_13378,N_14492);
or U15650 (N_15650,N_13859,N_12550);
nor U15651 (N_15651,N_13198,N_13162);
or U15652 (N_15652,N_13166,N_13744);
xor U15653 (N_15653,N_14394,N_13220);
nor U15654 (N_15654,N_14774,N_14277);
or U15655 (N_15655,N_13199,N_14167);
xnor U15656 (N_15656,N_14145,N_14571);
xor U15657 (N_15657,N_14240,N_13612);
nand U15658 (N_15658,N_12826,N_13784);
nor U15659 (N_15659,N_14671,N_14544);
nor U15660 (N_15660,N_12929,N_14838);
or U15661 (N_15661,N_14192,N_13479);
nor U15662 (N_15662,N_14090,N_13745);
or U15663 (N_15663,N_14380,N_14372);
or U15664 (N_15664,N_13699,N_13427);
nand U15665 (N_15665,N_13598,N_14681);
nor U15666 (N_15666,N_13203,N_14465);
or U15667 (N_15667,N_14261,N_14343);
and U15668 (N_15668,N_14744,N_13588);
and U15669 (N_15669,N_13176,N_13472);
or U15670 (N_15670,N_14453,N_14237);
xor U15671 (N_15671,N_12718,N_12530);
or U15672 (N_15672,N_14060,N_13453);
xnor U15673 (N_15673,N_14723,N_14748);
nor U15674 (N_15674,N_13751,N_14949);
and U15675 (N_15675,N_12899,N_14250);
xnor U15676 (N_15676,N_13154,N_13526);
nand U15677 (N_15677,N_13855,N_14100);
nand U15678 (N_15678,N_13089,N_14694);
or U15679 (N_15679,N_13460,N_13136);
or U15680 (N_15680,N_12725,N_13405);
or U15681 (N_15681,N_13428,N_14877);
xnor U15682 (N_15682,N_12587,N_13040);
nand U15683 (N_15683,N_14741,N_12845);
nand U15684 (N_15684,N_12909,N_12764);
nand U15685 (N_15685,N_13465,N_14202);
nand U15686 (N_15686,N_13439,N_13639);
and U15687 (N_15687,N_13817,N_13785);
and U15688 (N_15688,N_14801,N_13675);
nor U15689 (N_15689,N_14280,N_14299);
nand U15690 (N_15690,N_14658,N_13831);
xor U15691 (N_15691,N_14358,N_14490);
nand U15692 (N_15692,N_14672,N_14570);
or U15693 (N_15693,N_14369,N_14499);
xnor U15694 (N_15694,N_14078,N_14307);
and U15695 (N_15695,N_14095,N_14637);
and U15696 (N_15696,N_14330,N_12804);
and U15697 (N_15697,N_13704,N_14366);
nor U15698 (N_15698,N_13654,N_12595);
or U15699 (N_15699,N_13954,N_14848);
or U15700 (N_15700,N_12869,N_13987);
or U15701 (N_15701,N_13677,N_14434);
nand U15702 (N_15702,N_14804,N_14058);
and U15703 (N_15703,N_12674,N_14180);
and U15704 (N_15704,N_12768,N_14734);
xor U15705 (N_15705,N_14916,N_12975);
xor U15706 (N_15706,N_14339,N_13553);
or U15707 (N_15707,N_12682,N_12815);
nand U15708 (N_15708,N_14425,N_14397);
xnor U15709 (N_15709,N_12579,N_12761);
and U15710 (N_15710,N_14000,N_14722);
and U15711 (N_15711,N_14845,N_13659);
or U15712 (N_15712,N_14412,N_14117);
xnor U15713 (N_15713,N_12650,N_13232);
or U15714 (N_15714,N_14909,N_14684);
xnor U15715 (N_15715,N_14133,N_14062);
or U15716 (N_15716,N_12752,N_12794);
nor U15717 (N_15717,N_13155,N_14512);
or U15718 (N_15718,N_13409,N_13087);
and U15719 (N_15719,N_14690,N_14501);
or U15720 (N_15720,N_12812,N_13108);
xnor U15721 (N_15721,N_12546,N_13372);
nand U15722 (N_15722,N_14387,N_13272);
and U15723 (N_15723,N_12964,N_12737);
or U15724 (N_15724,N_14935,N_14924);
xor U15725 (N_15725,N_14329,N_12972);
and U15726 (N_15726,N_14730,N_12820);
xor U15727 (N_15727,N_14424,N_14814);
and U15728 (N_15728,N_12967,N_14516);
nand U15729 (N_15729,N_13305,N_14429);
nand U15730 (N_15730,N_14657,N_14963);
or U15731 (N_15731,N_14193,N_13138);
nand U15732 (N_15732,N_13013,N_14088);
nor U15733 (N_15733,N_14834,N_12642);
nand U15734 (N_15734,N_13400,N_12957);
nor U15735 (N_15735,N_13376,N_14254);
xnor U15736 (N_15736,N_12903,N_12700);
xor U15737 (N_15737,N_12561,N_13742);
nor U15738 (N_15738,N_13382,N_13881);
nor U15739 (N_15739,N_14920,N_13819);
xor U15740 (N_15740,N_13291,N_13132);
xnor U15741 (N_15741,N_13095,N_12965);
nand U15742 (N_15742,N_12735,N_14879);
or U15743 (N_15743,N_13769,N_13300);
or U15744 (N_15744,N_12855,N_13869);
or U15745 (N_15745,N_14595,N_13678);
or U15746 (N_15746,N_13227,N_13501);
and U15747 (N_15747,N_12793,N_13505);
xnor U15748 (N_15748,N_12780,N_13923);
nor U15749 (N_15749,N_14268,N_12527);
nand U15750 (N_15750,N_13297,N_12573);
xnor U15751 (N_15751,N_14974,N_13133);
nor U15752 (N_15752,N_14333,N_13858);
nand U15753 (N_15753,N_14318,N_14905);
xor U15754 (N_15754,N_12989,N_12596);
nor U15755 (N_15755,N_14043,N_12695);
nand U15756 (N_15756,N_14070,N_13709);
or U15757 (N_15757,N_14556,N_13467);
xnor U15758 (N_15758,N_14450,N_13961);
and U15759 (N_15759,N_13191,N_12722);
or U15760 (N_15760,N_14460,N_12796);
nor U15761 (N_15761,N_14319,N_14260);
and U15762 (N_15762,N_13584,N_13485);
nand U15763 (N_15763,N_13370,N_14547);
nand U15764 (N_15764,N_14765,N_14484);
nor U15765 (N_15765,N_13648,N_14386);
nand U15766 (N_15766,N_13167,N_13557);
or U15767 (N_15767,N_14785,N_12590);
nor U15768 (N_15768,N_13844,N_13292);
nor U15769 (N_15769,N_13473,N_12943);
or U15770 (N_15770,N_13283,N_13105);
nand U15771 (N_15771,N_13843,N_13740);
nand U15772 (N_15772,N_14844,N_13107);
nor U15773 (N_15773,N_13846,N_13823);
nand U15774 (N_15774,N_13075,N_12891);
or U15775 (N_15775,N_13316,N_13375);
nor U15776 (N_15776,N_14904,N_13222);
nor U15777 (N_15777,N_14936,N_12797);
nand U15778 (N_15778,N_12821,N_14409);
nor U15779 (N_15779,N_14376,N_12666);
nor U15780 (N_15780,N_13477,N_13997);
nor U15781 (N_15781,N_14568,N_13777);
and U15782 (N_15782,N_13496,N_14823);
xor U15783 (N_15783,N_12623,N_14562);
nand U15784 (N_15784,N_14421,N_14413);
xnor U15785 (N_15785,N_13060,N_14939);
nor U15786 (N_15786,N_14175,N_13242);
and U15787 (N_15787,N_14866,N_13737);
or U15788 (N_15788,N_13791,N_13634);
xnor U15789 (N_15789,N_14189,N_14973);
nor U15790 (N_15790,N_13812,N_12921);
and U15791 (N_15791,N_13210,N_13328);
nand U15792 (N_15792,N_14164,N_13134);
nor U15793 (N_15793,N_14082,N_13705);
nand U15794 (N_15794,N_14867,N_12885);
nor U15795 (N_15795,N_12872,N_13594);
xnor U15796 (N_15796,N_12918,N_14791);
xor U15797 (N_15797,N_12641,N_14344);
nand U15798 (N_15798,N_13070,N_12832);
or U15799 (N_15799,N_13310,N_14174);
nand U15800 (N_15800,N_12511,N_13275);
nor U15801 (N_15801,N_14220,N_14947);
and U15802 (N_15802,N_13607,N_13278);
or U15803 (N_15803,N_14203,N_13128);
and U15804 (N_15804,N_14559,N_14648);
and U15805 (N_15805,N_14588,N_14468);
and U15806 (N_15806,N_12833,N_13365);
nor U15807 (N_15807,N_13948,N_14725);
nand U15808 (N_15808,N_14448,N_13597);
nor U15809 (N_15809,N_12767,N_14217);
or U15810 (N_15810,N_14119,N_13182);
xnor U15811 (N_15811,N_12944,N_12795);
or U15812 (N_15812,N_14850,N_12517);
and U15813 (N_15813,N_13952,N_14246);
nand U15814 (N_15814,N_12880,N_14459);
and U15815 (N_15815,N_13256,N_14437);
nand U15816 (N_15816,N_13282,N_14697);
and U15817 (N_15817,N_13458,N_13302);
nor U15818 (N_15818,N_14288,N_13660);
nand U15819 (N_15819,N_13601,N_14005);
and U15820 (N_15820,N_14779,N_13530);
or U15821 (N_15821,N_12644,N_13535);
nand U15822 (N_15822,N_14597,N_13281);
nand U15823 (N_15823,N_13214,N_14228);
and U15824 (N_15824,N_14993,N_12874);
and U15825 (N_15825,N_13014,N_13169);
nand U15826 (N_15826,N_13329,N_13874);
nand U15827 (N_15827,N_13356,N_14911);
nor U15828 (N_15828,N_13323,N_14293);
nor U15829 (N_15829,N_13094,N_13789);
or U15830 (N_15830,N_12783,N_13558);
xnor U15831 (N_15831,N_12645,N_12592);
nand U15832 (N_15832,N_12634,N_14400);
and U15833 (N_15833,N_14865,N_14660);
and U15834 (N_15834,N_14899,N_14828);
xor U15835 (N_15835,N_12848,N_13438);
or U15836 (N_15836,N_14470,N_13313);
and U15837 (N_15837,N_13468,N_13932);
or U15838 (N_15838,N_12924,N_12626);
nand U15839 (N_15839,N_13122,N_13684);
and U15840 (N_15840,N_14362,N_13401);
xor U15841 (N_15841,N_13908,N_14076);
nand U15842 (N_15842,N_13878,N_13849);
and U15843 (N_15843,N_13464,N_12781);
nand U15844 (N_15844,N_13011,N_13097);
nand U15845 (N_15845,N_13536,N_12531);
or U15846 (N_15846,N_13687,N_14942);
xnor U15847 (N_15847,N_13436,N_12684);
or U15848 (N_15848,N_13111,N_13113);
and U15849 (N_15849,N_14345,N_13327);
or U15850 (N_15850,N_12814,N_13871);
and U15851 (N_15851,N_13665,N_12835);
nand U15852 (N_15852,N_14403,N_14915);
and U15853 (N_15853,N_14506,N_12978);
nand U15854 (N_15854,N_14534,N_13118);
and U15855 (N_15855,N_14783,N_13440);
or U15856 (N_15856,N_14560,N_14337);
or U15857 (N_15857,N_12601,N_12667);
nor U15858 (N_15858,N_12668,N_12828);
and U15859 (N_15859,N_13110,N_14391);
nor U15860 (N_15860,N_14611,N_13564);
xnor U15861 (N_15861,N_13554,N_14461);
and U15862 (N_15862,N_14027,N_12823);
and U15863 (N_15863,N_13524,N_13342);
or U15864 (N_15864,N_14796,N_14605);
and U15865 (N_15865,N_14627,N_14134);
nor U15866 (N_15866,N_12995,N_13979);
and U15867 (N_15867,N_14294,N_14466);
nor U15868 (N_15868,N_14927,N_12888);
or U15869 (N_15869,N_12548,N_13761);
or U15870 (N_15870,N_14347,N_12683);
xnor U15871 (N_15871,N_13189,N_13988);
xnor U15872 (N_15872,N_13940,N_13259);
xor U15873 (N_15873,N_13418,N_14932);
nor U15874 (N_15874,N_13879,N_13587);
nor U15875 (N_15875,N_14702,N_14390);
xnor U15876 (N_15876,N_14862,N_14532);
nor U15877 (N_15877,N_13158,N_13358);
nor U15878 (N_15878,N_13716,N_13579);
xor U15879 (N_15879,N_13425,N_13608);
nor U15880 (N_15880,N_14520,N_13403);
or U15881 (N_15881,N_12509,N_12660);
xor U15882 (N_15882,N_14273,N_13778);
nor U15883 (N_15883,N_12535,N_12760);
nor U15884 (N_15884,N_14422,N_13385);
nand U15885 (N_15885,N_13957,N_13121);
or U15886 (N_15886,N_14795,N_14830);
nand U15887 (N_15887,N_14549,N_14061);
xor U15888 (N_15888,N_13035,N_13866);
nand U15889 (N_15889,N_14514,N_14176);
nor U15890 (N_15890,N_12865,N_14227);
and U15891 (N_15891,N_12514,N_14536);
xor U15892 (N_15892,N_13865,N_12659);
and U15893 (N_15893,N_14956,N_12542);
and U15894 (N_15894,N_14737,N_14749);
xnor U15895 (N_15895,N_14984,N_13559);
xor U15896 (N_15896,N_12678,N_13729);
nor U15897 (N_15897,N_13025,N_14603);
or U15898 (N_15898,N_12916,N_13516);
nor U15899 (N_15899,N_13424,N_14952);
and U15900 (N_15900,N_13354,N_14743);
and U15901 (N_15901,N_13837,N_13286);
nor U15902 (N_15902,N_14890,N_13062);
nand U15903 (N_15903,N_14701,N_13642);
nand U15904 (N_15904,N_14929,N_13462);
xnor U15905 (N_15905,N_14880,N_12765);
xor U15906 (N_15906,N_14243,N_12670);
xor U15907 (N_15907,N_13096,N_13042);
and U15908 (N_15908,N_13640,N_14001);
or U15909 (N_15909,N_12908,N_12632);
and U15910 (N_15910,N_13032,N_14023);
nand U15911 (N_15911,N_14456,N_12935);
nor U15912 (N_15912,N_14840,N_14668);
nor U15913 (N_15913,N_12615,N_13115);
xor U15914 (N_15914,N_13717,N_14092);
or U15915 (N_15915,N_14151,N_14104);
xnor U15916 (N_15916,N_14381,N_13692);
or U15917 (N_15917,N_12854,N_12633);
and U15918 (N_15918,N_14781,N_14360);
and U15919 (N_15919,N_12612,N_13697);
xor U15920 (N_15920,N_14803,N_13248);
nor U15921 (N_15921,N_13065,N_14653);
nand U15922 (N_15922,N_14066,N_13628);
nor U15923 (N_15923,N_14912,N_14313);
nor U15924 (N_15924,N_14433,N_13975);
and U15925 (N_15925,N_14755,N_12743);
and U15926 (N_15926,N_13290,N_13552);
nor U15927 (N_15927,N_14978,N_13123);
or U15928 (N_15928,N_13147,N_12580);
nand U15929 (N_15929,N_13056,N_13183);
or U15930 (N_15930,N_12914,N_14004);
and U15931 (N_15931,N_14854,N_14503);
or U15932 (N_15932,N_13840,N_13367);
or U15933 (N_15933,N_14642,N_13847);
xor U15934 (N_15934,N_14543,N_14604);
and U15935 (N_15935,N_13159,N_12881);
nand U15936 (N_15936,N_14831,N_12520);
nor U15937 (N_15937,N_13690,N_13863);
or U15938 (N_15938,N_13956,N_13896);
nor U15939 (N_15939,N_14108,N_13336);
nor U15940 (N_15940,N_14442,N_13707);
xor U15941 (N_15941,N_12545,N_12697);
nor U15942 (N_15942,N_13661,N_14116);
xnor U15943 (N_15943,N_12766,N_13319);
or U15944 (N_15944,N_14052,N_13613);
xnor U15945 (N_15945,N_14849,N_14209);
xor U15946 (N_15946,N_14519,N_14323);
and U15947 (N_15947,N_13521,N_14342);
or U15948 (N_15948,N_14763,N_14720);
or U15949 (N_15949,N_14777,N_14140);
or U15950 (N_15950,N_12866,N_12600);
or U15951 (N_15951,N_13230,N_13429);
nand U15952 (N_15952,N_12731,N_12999);
xnor U15953 (N_15953,N_14211,N_14590);
xor U15954 (N_15954,N_13655,N_13543);
or U15955 (N_15955,N_12983,N_12621);
or U15956 (N_15956,N_12614,N_12694);
xnor U15957 (N_15957,N_13306,N_14788);
or U15958 (N_15958,N_13000,N_12563);
nand U15959 (N_15959,N_13813,N_13225);
xnor U15960 (N_15960,N_14316,N_13926);
and U15961 (N_15961,N_13497,N_13990);
nor U15962 (N_15962,N_13625,N_14651);
xor U15963 (N_15963,N_14481,N_12778);
nand U15964 (N_15964,N_12699,N_14086);
or U15965 (N_15965,N_14759,N_14527);
or U15966 (N_15966,N_14710,N_14691);
nand U15967 (N_15967,N_12830,N_13862);
xnor U15968 (N_15968,N_14925,N_14229);
or U15969 (N_15969,N_13326,N_13893);
nand U15970 (N_15970,N_13036,N_13732);
xor U15971 (N_15971,N_14234,N_13049);
nor U15972 (N_15972,N_13318,N_13937);
or U15973 (N_15973,N_13026,N_13250);
nor U15974 (N_15974,N_13590,N_13897);
nor U15975 (N_15975,N_14992,N_14044);
nand U15976 (N_15976,N_14817,N_12811);
nand U15977 (N_15977,N_13068,N_14297);
and U15978 (N_15978,N_13324,N_13239);
xor U15979 (N_15979,N_12544,N_12636);
nand U15980 (N_15980,N_13489,N_13322);
nor U15981 (N_15981,N_13083,N_14599);
xnor U15982 (N_15982,N_14860,N_13033);
and U15983 (N_15983,N_12503,N_14451);
nor U15984 (N_15984,N_13088,N_14987);
nand U15985 (N_15985,N_13377,N_14873);
nand U15986 (N_15986,N_14677,N_12740);
or U15987 (N_15987,N_14812,N_13993);
xnor U15988 (N_15988,N_12685,N_14482);
nor U15989 (N_15989,N_14037,N_12939);
and U15990 (N_15990,N_14594,N_13104);
nor U15991 (N_15991,N_14715,N_13263);
nor U15992 (N_15992,N_12887,N_14625);
nor U15993 (N_15993,N_14126,N_13546);
nor U15994 (N_15994,N_13005,N_13918);
xnor U15995 (N_15995,N_14085,N_14148);
or U15996 (N_15996,N_12742,N_14583);
nor U15997 (N_15997,N_13674,N_14821);
or U15998 (N_15998,N_14168,N_13461);
nor U15999 (N_15999,N_14028,N_13638);
or U16000 (N_16000,N_13548,N_14542);
nor U16001 (N_16001,N_13492,N_14263);
nand U16002 (N_16002,N_14232,N_13533);
nor U16003 (N_16003,N_14500,N_13934);
and U16004 (N_16004,N_13984,N_14778);
nand U16005 (N_16005,N_14954,N_13412);
nor U16006 (N_16006,N_13218,N_12807);
xnor U16007 (N_16007,N_13215,N_12703);
xnor U16008 (N_16008,N_14406,N_12769);
or U16009 (N_16009,N_14678,N_13591);
nand U16010 (N_16010,N_14171,N_13788);
xor U16011 (N_16011,N_14212,N_12837);
nor U16012 (N_16012,N_13867,N_13735);
xor U16013 (N_16013,N_13361,N_13034);
nor U16014 (N_16014,N_14186,N_14411);
or U16015 (N_16015,N_12705,N_13251);
and U16016 (N_16016,N_14215,N_13989);
nor U16017 (N_16017,N_13746,N_12704);
and U16018 (N_16018,N_14364,N_12839);
xnor U16019 (N_16019,N_12756,N_14385);
nor U16020 (N_16020,N_13959,N_13178);
nand U16021 (N_16021,N_14665,N_14166);
or U16022 (N_16022,N_14622,N_13643);
and U16023 (N_16023,N_14087,N_13184);
nor U16024 (N_16024,N_14931,N_14414);
xor U16025 (N_16025,N_13636,N_13024);
xnor U16026 (N_16026,N_14236,N_14008);
xnor U16027 (N_16027,N_14628,N_14320);
xor U16028 (N_16028,N_14666,N_13130);
nand U16029 (N_16029,N_13877,N_13756);
nor U16030 (N_16030,N_14820,N_13972);
nor U16031 (N_16031,N_14278,N_14173);
nor U16032 (N_16032,N_12676,N_14181);
nor U16033 (N_16033,N_14139,N_12970);
xnor U16034 (N_16034,N_14863,N_12987);
and U16035 (N_16035,N_14056,N_12611);
or U16036 (N_16036,N_12608,N_13031);
nor U16037 (N_16037,N_13620,N_13714);
or U16038 (N_16038,N_14352,N_13363);
xnor U16039 (N_16039,N_14324,N_13652);
xnor U16040 (N_16040,N_14169,N_14882);
or U16041 (N_16041,N_13886,N_13924);
nor U16042 (N_16042,N_12662,N_14639);
nor U16043 (N_16043,N_13311,N_14432);
or U16044 (N_16044,N_13828,N_13753);
nor U16045 (N_16045,N_13480,N_13012);
and U16046 (N_16046,N_13237,N_12977);
nand U16047 (N_16047,N_12715,N_14336);
and U16048 (N_16048,N_14011,N_13016);
or U16049 (N_16049,N_12729,N_13739);
or U16050 (N_16050,N_12867,N_14727);
or U16051 (N_16051,N_13801,N_12786);
nor U16052 (N_16052,N_13765,N_13624);
and U16053 (N_16053,N_14136,N_12578);
or U16054 (N_16054,N_13127,N_14208);
xnor U16055 (N_16055,N_12941,N_14760);
or U16056 (N_16056,N_13426,N_14321);
xor U16057 (N_16057,N_13894,N_12755);
nor U16058 (N_16058,N_13950,N_14274);
and U16059 (N_16059,N_13229,N_12664);
xnor U16060 (N_16060,N_12961,N_14897);
or U16061 (N_16061,N_13129,N_13835);
nor U16062 (N_16062,N_13269,N_13991);
nor U16063 (N_16063,N_13885,N_14349);
nand U16064 (N_16064,N_14152,N_12890);
nor U16065 (N_16065,N_14718,N_13074);
nand U16066 (N_16066,N_14296,N_13463);
or U16067 (N_16067,N_13437,N_14141);
and U16068 (N_16068,N_14020,N_14884);
xnor U16069 (N_16069,N_12584,N_12720);
or U16070 (N_16070,N_12868,N_13930);
nand U16071 (N_16071,N_14561,N_14621);
and U16072 (N_16072,N_13929,N_13818);
nand U16073 (N_16073,N_12551,N_14235);
nand U16074 (N_16074,N_14525,N_12585);
and U16075 (N_16075,N_12714,N_14019);
or U16076 (N_16076,N_13080,N_14999);
nor U16077 (N_16077,N_14283,N_14357);
nand U16078 (N_16078,N_13393,N_14922);
or U16079 (N_16079,N_14654,N_14353);
nor U16080 (N_16080,N_14322,N_14797);
nand U16081 (N_16081,N_12532,N_13963);
xnor U16082 (N_16082,N_14617,N_14586);
nor U16083 (N_16083,N_12540,N_14719);
and U16084 (N_16084,N_14907,N_14115);
xnor U16085 (N_16085,N_12619,N_14312);
or U16086 (N_16086,N_14122,N_12889);
xnor U16087 (N_16087,N_14269,N_12938);
or U16088 (N_16088,N_14965,N_13100);
nor U16089 (N_16089,N_14529,N_14847);
nor U16090 (N_16090,N_12884,N_14471);
nor U16091 (N_16091,N_13514,N_13190);
xor U16092 (N_16092,N_14051,N_13890);
nand U16093 (N_16093,N_12945,N_12894);
and U16094 (N_16094,N_13764,N_14170);
xor U16095 (N_16095,N_12917,N_14871);
nor U16096 (N_16096,N_13063,N_12856);
nor U16097 (N_16097,N_13799,N_13090);
or U16098 (N_16098,N_13255,N_12907);
or U16099 (N_16099,N_13148,N_13883);
xor U16100 (N_16100,N_14124,N_13398);
and U16101 (N_16101,N_12638,N_14565);
xor U16102 (N_16102,N_13808,N_14046);
nor U16103 (N_16103,N_14272,N_12653);
nor U16104 (N_16104,N_14950,N_13617);
or U16105 (N_16105,N_13337,N_13738);
nor U16106 (N_16106,N_13759,N_14069);
nor U16107 (N_16107,N_14504,N_12996);
nor U16108 (N_16108,N_13386,N_14695);
nand U16109 (N_16109,N_12648,N_14995);
nor U16110 (N_16110,N_14546,N_13200);
and U16111 (N_16111,N_14426,N_14271);
and U16112 (N_16112,N_14190,N_14346);
or U16113 (N_16113,N_13771,N_13015);
or U16114 (N_16114,N_12772,N_12798);
nor U16115 (N_16115,N_14959,N_12602);
or U16116 (N_16116,N_14928,N_13953);
nand U16117 (N_16117,N_14735,N_13992);
and U16118 (N_16118,N_14480,N_12655);
or U16119 (N_16119,N_14800,N_14388);
nand U16120 (N_16120,N_13456,N_14813);
or U16121 (N_16121,N_13445,N_12681);
or U16122 (N_16122,N_14094,N_13912);
or U16123 (N_16123,N_13205,N_14467);
or U16124 (N_16124,N_14685,N_14013);
and U16125 (N_16125,N_13574,N_13800);
and U16126 (N_16126,N_14647,N_13163);
nor U16127 (N_16127,N_13213,N_12870);
nor U16128 (N_16128,N_14966,N_13527);
xor U16129 (N_16129,N_14377,N_13887);
nor U16130 (N_16130,N_14325,N_14756);
or U16131 (N_16131,N_14798,N_14034);
nor U16132 (N_16132,N_13519,N_12730);
or U16133 (N_16133,N_14498,N_13681);
and U16134 (N_16134,N_13561,N_12646);
or U16135 (N_16135,N_13825,N_12690);
or U16136 (N_16136,N_12883,N_14626);
nand U16137 (N_16137,N_13946,N_14998);
or U16138 (N_16138,N_14317,N_12785);
nor U16139 (N_16139,N_12922,N_14901);
xnor U16140 (N_16140,N_13982,N_14006);
nor U16141 (N_16141,N_13388,N_14664);
xnor U16142 (N_16142,N_14018,N_13124);
nand U16143 (N_16143,N_12622,N_12834);
and U16144 (N_16144,N_13069,N_13331);
xor U16145 (N_16145,N_13430,N_13488);
xor U16146 (N_16146,N_14982,N_14986);
nand U16147 (N_16147,N_14256,N_13077);
xor U16148 (N_16148,N_12840,N_14458);
nand U16149 (N_16149,N_13562,N_13491);
and U16150 (N_16150,N_14692,N_13797);
or U16151 (N_16151,N_13019,N_14733);
xor U16152 (N_16152,N_13903,N_12519);
and U16153 (N_16153,N_14574,N_13814);
and U16154 (N_16154,N_13493,N_14906);
nor U16155 (N_16155,N_13507,N_13545);
nand U16156 (N_16156,N_13537,N_13161);
xnor U16157 (N_16157,N_14348,N_14093);
or U16158 (N_16158,N_13815,N_12988);
xor U16159 (N_16159,N_13686,N_13715);
or U16160 (N_16160,N_13996,N_12680);
nand U16161 (N_16161,N_13009,N_13550);
nand U16162 (N_16162,N_13362,N_12620);
and U16163 (N_16163,N_13209,N_13515);
nand U16164 (N_16164,N_12897,N_14937);
nand U16165 (N_16165,N_12734,N_14852);
xor U16166 (N_16166,N_14047,N_13360);
or U16167 (N_16167,N_14530,N_13829);
xor U16168 (N_16168,N_14510,N_14716);
xnor U16169 (N_16169,N_12526,N_14581);
xor U16170 (N_16170,N_14225,N_13145);
xnor U16171 (N_16171,N_14014,N_12933);
and U16172 (N_16172,N_13506,N_13078);
nand U16173 (N_16173,N_13194,N_12625);
and U16174 (N_16174,N_14130,N_12688);
xor U16175 (N_16175,N_13258,N_13680);
xor U16176 (N_16176,N_13824,N_13585);
and U16177 (N_16177,N_13082,N_14609);
or U16178 (N_16178,N_14643,N_12915);
and U16179 (N_16179,N_13380,N_14079);
and U16180 (N_16180,N_14771,N_14887);
nor U16181 (N_16181,N_13921,N_12733);
nand U16182 (N_16182,N_14495,N_13043);
xnor U16183 (N_16183,N_13052,N_12777);
or U16184 (N_16184,N_12501,N_13794);
xor U16185 (N_16185,N_14487,N_12900);
nand U16186 (N_16186,N_12723,N_14440);
xnor U16187 (N_16187,N_12552,N_13693);
or U16188 (N_16188,N_13257,N_13841);
or U16189 (N_16189,N_14502,N_13719);
and U16190 (N_16190,N_13555,N_14127);
nor U16191 (N_16191,N_13139,N_13820);
or U16192 (N_16192,N_14291,N_12806);
nand U16193 (N_16193,N_13706,N_14123);
nor U16194 (N_16194,N_12549,N_13741);
nand U16195 (N_16195,N_14945,N_13949);
xnor U16196 (N_16196,N_13786,N_13773);
and U16197 (N_16197,N_13694,N_14204);
and U16198 (N_16198,N_12862,N_14401);
xnor U16199 (N_16199,N_14213,N_12925);
or U16200 (N_16200,N_14239,N_13722);
nor U16201 (N_16201,N_12762,N_13187);
nand U16202 (N_16202,N_14600,N_13152);
or U16203 (N_16203,N_13967,N_14991);
and U16204 (N_16204,N_13308,N_13798);
xor U16205 (N_16205,N_14842,N_13307);
and U16206 (N_16206,N_12947,N_12810);
nor U16207 (N_16207,N_13244,N_13663);
xor U16208 (N_16208,N_14367,N_14197);
or U16209 (N_16209,N_14363,N_12665);
and U16210 (N_16210,N_13651,N_14068);
and U16211 (N_16211,N_14822,N_13683);
nand U16212 (N_16212,N_12923,N_12824);
nor U16213 (N_16213,N_12721,N_13003);
and U16214 (N_16214,N_12847,N_14683);
nor U16215 (N_16215,N_13067,N_12504);
or U16216 (N_16216,N_14961,N_13475);
xnor U16217 (N_16217,N_14640,N_14101);
nor U16218 (N_16218,N_14129,N_13346);
xor U16219 (N_16219,N_13668,N_13168);
nand U16220 (N_16220,N_14473,N_12710);
xnor U16221 (N_16221,N_13299,N_14636);
nor U16222 (N_16222,N_12556,N_13868);
and U16223 (N_16223,N_12800,N_13748);
nand U16224 (N_16224,N_13193,N_14770);
nand U16225 (N_16225,N_14185,N_14084);
nand U16226 (N_16226,N_13023,N_13116);
nor U16227 (N_16227,N_13416,N_14789);
nand U16228 (N_16228,N_14994,N_12878);
nand U16229 (N_16229,N_12776,N_14620);
xnor U16230 (N_16230,N_13314,N_14951);
or U16231 (N_16231,N_14075,N_13509);
xnor U16232 (N_16232,N_14035,N_14699);
or U16233 (N_16233,N_14382,N_14032);
and U16234 (N_16234,N_14584,N_13420);
nand U16235 (N_16235,N_13911,N_12672);
nor U16236 (N_16236,N_14853,N_13790);
and U16237 (N_16237,N_14933,N_13058);
and U16238 (N_16238,N_14304,N_13389);
nor U16239 (N_16239,N_13419,N_14836);
nand U16240 (N_16240,N_14983,N_12976);
nor U16241 (N_16241,N_14802,N_12574);
nand U16242 (N_16242,N_13371,N_14172);
xnor U16243 (N_16243,N_12906,N_12932);
nor U16244 (N_16244,N_12852,N_14420);
nor U16245 (N_16245,N_13442,N_13551);
or U16246 (N_16246,N_13135,N_14633);
xor U16247 (N_16247,N_12898,N_12571);
or U16248 (N_16248,N_12679,N_12701);
nor U16249 (N_16249,N_13030,N_13457);
or U16250 (N_16250,N_12622,N_13779);
or U16251 (N_16251,N_13202,N_14455);
or U16252 (N_16252,N_13308,N_13006);
nand U16253 (N_16253,N_13959,N_14738);
and U16254 (N_16254,N_12837,N_14925);
or U16255 (N_16255,N_13883,N_13691);
or U16256 (N_16256,N_13013,N_13724);
nor U16257 (N_16257,N_13084,N_12980);
nand U16258 (N_16258,N_14839,N_13795);
nor U16259 (N_16259,N_12758,N_14513);
and U16260 (N_16260,N_13755,N_13184);
or U16261 (N_16261,N_13154,N_12632);
or U16262 (N_16262,N_14486,N_14868);
or U16263 (N_16263,N_12683,N_14094);
nor U16264 (N_16264,N_13844,N_14045);
nand U16265 (N_16265,N_13192,N_14579);
and U16266 (N_16266,N_13670,N_12997);
or U16267 (N_16267,N_14387,N_14019);
or U16268 (N_16268,N_13487,N_13579);
xnor U16269 (N_16269,N_14585,N_13411);
or U16270 (N_16270,N_13783,N_13210);
xnor U16271 (N_16271,N_13039,N_14036);
or U16272 (N_16272,N_13147,N_12677);
or U16273 (N_16273,N_13906,N_13009);
xor U16274 (N_16274,N_14272,N_14579);
nor U16275 (N_16275,N_12950,N_14019);
or U16276 (N_16276,N_14672,N_13291);
or U16277 (N_16277,N_14792,N_14703);
or U16278 (N_16278,N_13045,N_13854);
nand U16279 (N_16279,N_14718,N_14140);
xor U16280 (N_16280,N_12903,N_13794);
nor U16281 (N_16281,N_12764,N_14826);
nor U16282 (N_16282,N_13304,N_14823);
or U16283 (N_16283,N_14997,N_14036);
and U16284 (N_16284,N_13129,N_14012);
nand U16285 (N_16285,N_14274,N_13476);
or U16286 (N_16286,N_14608,N_13444);
xnor U16287 (N_16287,N_13847,N_12579);
xor U16288 (N_16288,N_13197,N_14101);
xnor U16289 (N_16289,N_14409,N_14328);
xor U16290 (N_16290,N_13837,N_14787);
nand U16291 (N_16291,N_13962,N_14831);
nand U16292 (N_16292,N_14264,N_13339);
nor U16293 (N_16293,N_14362,N_13580);
nand U16294 (N_16294,N_12588,N_14291);
or U16295 (N_16295,N_13012,N_12558);
nand U16296 (N_16296,N_13760,N_12740);
xnor U16297 (N_16297,N_12871,N_14238);
nand U16298 (N_16298,N_13249,N_14094);
xor U16299 (N_16299,N_14173,N_12590);
nor U16300 (N_16300,N_13186,N_14812);
or U16301 (N_16301,N_12889,N_14191);
nand U16302 (N_16302,N_14493,N_13117);
nor U16303 (N_16303,N_14071,N_14361);
xnor U16304 (N_16304,N_13937,N_13216);
or U16305 (N_16305,N_14006,N_14790);
and U16306 (N_16306,N_13608,N_13333);
nand U16307 (N_16307,N_14312,N_13684);
nand U16308 (N_16308,N_13673,N_13487);
and U16309 (N_16309,N_14007,N_13289);
and U16310 (N_16310,N_13355,N_13268);
or U16311 (N_16311,N_14602,N_13708);
xnor U16312 (N_16312,N_14015,N_13637);
nor U16313 (N_16313,N_14337,N_14794);
xor U16314 (N_16314,N_14287,N_14380);
and U16315 (N_16315,N_13036,N_12870);
and U16316 (N_16316,N_13022,N_12551);
or U16317 (N_16317,N_13547,N_13511);
nand U16318 (N_16318,N_13718,N_13283);
xnor U16319 (N_16319,N_14327,N_12939);
nand U16320 (N_16320,N_14435,N_13688);
nand U16321 (N_16321,N_12759,N_13393);
or U16322 (N_16322,N_13943,N_14475);
and U16323 (N_16323,N_12836,N_12903);
or U16324 (N_16324,N_14584,N_13728);
xnor U16325 (N_16325,N_12981,N_13574);
or U16326 (N_16326,N_13923,N_14803);
nand U16327 (N_16327,N_14344,N_14661);
xnor U16328 (N_16328,N_13651,N_14375);
and U16329 (N_16329,N_13824,N_12956);
and U16330 (N_16330,N_14008,N_13284);
or U16331 (N_16331,N_14982,N_14084);
or U16332 (N_16332,N_14793,N_14485);
xor U16333 (N_16333,N_12931,N_14032);
and U16334 (N_16334,N_14178,N_12797);
nor U16335 (N_16335,N_14932,N_14853);
nand U16336 (N_16336,N_14693,N_14277);
nor U16337 (N_16337,N_14556,N_13861);
nor U16338 (N_16338,N_14738,N_12759);
nor U16339 (N_16339,N_14376,N_14959);
nor U16340 (N_16340,N_14706,N_13508);
nand U16341 (N_16341,N_14654,N_12523);
nand U16342 (N_16342,N_12507,N_14843);
nand U16343 (N_16343,N_14419,N_13254);
xnor U16344 (N_16344,N_13386,N_13563);
and U16345 (N_16345,N_13862,N_13731);
nor U16346 (N_16346,N_14628,N_14428);
nor U16347 (N_16347,N_12734,N_13326);
xnor U16348 (N_16348,N_13614,N_13737);
nor U16349 (N_16349,N_13157,N_14396);
or U16350 (N_16350,N_14217,N_14590);
nand U16351 (N_16351,N_12786,N_13811);
xnor U16352 (N_16352,N_14287,N_14089);
or U16353 (N_16353,N_14761,N_12979);
and U16354 (N_16354,N_14072,N_13509);
nand U16355 (N_16355,N_13846,N_14804);
or U16356 (N_16356,N_13759,N_14139);
or U16357 (N_16357,N_12565,N_13162);
and U16358 (N_16358,N_12841,N_13336);
and U16359 (N_16359,N_13299,N_12829);
and U16360 (N_16360,N_14199,N_14638);
nor U16361 (N_16361,N_14355,N_14787);
nand U16362 (N_16362,N_13214,N_14003);
nand U16363 (N_16363,N_14318,N_13415);
xor U16364 (N_16364,N_13833,N_14335);
nor U16365 (N_16365,N_13133,N_12913);
or U16366 (N_16366,N_14324,N_13401);
xor U16367 (N_16367,N_13040,N_12596);
xor U16368 (N_16368,N_14342,N_12619);
nor U16369 (N_16369,N_14498,N_13724);
or U16370 (N_16370,N_14340,N_13726);
nor U16371 (N_16371,N_14885,N_13880);
xnor U16372 (N_16372,N_13098,N_13319);
nor U16373 (N_16373,N_12534,N_13969);
xor U16374 (N_16374,N_14237,N_12923);
xor U16375 (N_16375,N_12999,N_13412);
and U16376 (N_16376,N_12827,N_14889);
nand U16377 (N_16377,N_14100,N_13745);
nand U16378 (N_16378,N_14728,N_14094);
nor U16379 (N_16379,N_12695,N_14631);
xor U16380 (N_16380,N_13152,N_14472);
nand U16381 (N_16381,N_13535,N_13265);
and U16382 (N_16382,N_13173,N_13572);
or U16383 (N_16383,N_13153,N_14627);
nand U16384 (N_16384,N_13530,N_14166);
xor U16385 (N_16385,N_14893,N_14417);
nor U16386 (N_16386,N_13009,N_14880);
xor U16387 (N_16387,N_13797,N_14868);
nor U16388 (N_16388,N_13456,N_13486);
or U16389 (N_16389,N_13721,N_14652);
xor U16390 (N_16390,N_12950,N_13920);
nand U16391 (N_16391,N_14268,N_14816);
xnor U16392 (N_16392,N_12552,N_12874);
nand U16393 (N_16393,N_14958,N_13644);
or U16394 (N_16394,N_14876,N_14892);
nand U16395 (N_16395,N_13213,N_13980);
nor U16396 (N_16396,N_13016,N_13513);
and U16397 (N_16397,N_13683,N_13701);
and U16398 (N_16398,N_12787,N_13891);
nand U16399 (N_16399,N_14122,N_12877);
nand U16400 (N_16400,N_12862,N_13575);
nand U16401 (N_16401,N_12762,N_13389);
nand U16402 (N_16402,N_13469,N_13058);
nand U16403 (N_16403,N_14229,N_13809);
nand U16404 (N_16404,N_14847,N_13031);
and U16405 (N_16405,N_14514,N_13167);
and U16406 (N_16406,N_13076,N_13665);
and U16407 (N_16407,N_13677,N_13290);
or U16408 (N_16408,N_14155,N_14775);
and U16409 (N_16409,N_14468,N_14699);
and U16410 (N_16410,N_13669,N_13087);
nor U16411 (N_16411,N_13660,N_13028);
nor U16412 (N_16412,N_12864,N_12874);
or U16413 (N_16413,N_12697,N_14939);
or U16414 (N_16414,N_12975,N_12740);
xnor U16415 (N_16415,N_12563,N_13290);
and U16416 (N_16416,N_14993,N_14839);
nand U16417 (N_16417,N_14113,N_13307);
nor U16418 (N_16418,N_13355,N_13920);
nor U16419 (N_16419,N_14934,N_14132);
xnor U16420 (N_16420,N_14415,N_12545);
nor U16421 (N_16421,N_14329,N_14693);
and U16422 (N_16422,N_13340,N_14176);
nor U16423 (N_16423,N_13844,N_13842);
nor U16424 (N_16424,N_13768,N_13898);
nor U16425 (N_16425,N_13232,N_14840);
nor U16426 (N_16426,N_14044,N_13337);
or U16427 (N_16427,N_14500,N_14411);
xnor U16428 (N_16428,N_13134,N_14241);
nand U16429 (N_16429,N_14282,N_12862);
nand U16430 (N_16430,N_13344,N_14133);
and U16431 (N_16431,N_14094,N_13305);
or U16432 (N_16432,N_14484,N_12666);
nand U16433 (N_16433,N_14712,N_13701);
and U16434 (N_16434,N_13272,N_12918);
and U16435 (N_16435,N_14279,N_13548);
nor U16436 (N_16436,N_14307,N_13689);
xnor U16437 (N_16437,N_12725,N_13852);
or U16438 (N_16438,N_13108,N_14461);
xor U16439 (N_16439,N_13694,N_13501);
or U16440 (N_16440,N_14055,N_12995);
and U16441 (N_16441,N_14359,N_12965);
or U16442 (N_16442,N_14555,N_14968);
nor U16443 (N_16443,N_13573,N_13968);
nand U16444 (N_16444,N_13047,N_13213);
or U16445 (N_16445,N_14733,N_13416);
xnor U16446 (N_16446,N_14551,N_13105);
or U16447 (N_16447,N_14962,N_13942);
or U16448 (N_16448,N_13468,N_13941);
nor U16449 (N_16449,N_12777,N_13081);
xor U16450 (N_16450,N_12596,N_13521);
and U16451 (N_16451,N_13261,N_13063);
and U16452 (N_16452,N_14113,N_13305);
or U16453 (N_16453,N_13833,N_14672);
nor U16454 (N_16454,N_14120,N_14578);
or U16455 (N_16455,N_13671,N_14167);
nand U16456 (N_16456,N_14732,N_13789);
xor U16457 (N_16457,N_12798,N_14248);
and U16458 (N_16458,N_13320,N_13444);
xnor U16459 (N_16459,N_13450,N_12613);
or U16460 (N_16460,N_14463,N_14810);
or U16461 (N_16461,N_13222,N_14679);
and U16462 (N_16462,N_14227,N_13764);
xor U16463 (N_16463,N_13210,N_12940);
xnor U16464 (N_16464,N_13205,N_13908);
nor U16465 (N_16465,N_12853,N_14069);
nor U16466 (N_16466,N_14284,N_14635);
or U16467 (N_16467,N_12640,N_12701);
xor U16468 (N_16468,N_12529,N_14566);
nand U16469 (N_16469,N_13460,N_14605);
and U16470 (N_16470,N_13203,N_13099);
xnor U16471 (N_16471,N_14890,N_14847);
and U16472 (N_16472,N_14235,N_14336);
or U16473 (N_16473,N_13453,N_13710);
xor U16474 (N_16474,N_14575,N_12995);
nor U16475 (N_16475,N_12798,N_13223);
and U16476 (N_16476,N_13725,N_12571);
or U16477 (N_16477,N_14914,N_13274);
and U16478 (N_16478,N_14789,N_14781);
xnor U16479 (N_16479,N_13969,N_13268);
nand U16480 (N_16480,N_13247,N_12824);
or U16481 (N_16481,N_13310,N_14974);
nor U16482 (N_16482,N_13811,N_12575);
xnor U16483 (N_16483,N_14841,N_13995);
nor U16484 (N_16484,N_12692,N_13048);
or U16485 (N_16485,N_14208,N_13514);
and U16486 (N_16486,N_12798,N_14226);
nand U16487 (N_16487,N_14598,N_13768);
xor U16488 (N_16488,N_14636,N_12740);
xnor U16489 (N_16489,N_12981,N_13395);
nor U16490 (N_16490,N_14379,N_12866);
nor U16491 (N_16491,N_14385,N_14989);
nand U16492 (N_16492,N_14851,N_14881);
and U16493 (N_16493,N_14713,N_12962);
nand U16494 (N_16494,N_12570,N_13614);
xnor U16495 (N_16495,N_14852,N_12778);
or U16496 (N_16496,N_13387,N_12899);
xnor U16497 (N_16497,N_12734,N_14586);
or U16498 (N_16498,N_14368,N_13878);
or U16499 (N_16499,N_13072,N_14186);
xnor U16500 (N_16500,N_13294,N_14939);
xnor U16501 (N_16501,N_14944,N_13803);
or U16502 (N_16502,N_13586,N_14428);
and U16503 (N_16503,N_12889,N_14515);
and U16504 (N_16504,N_12900,N_14513);
xor U16505 (N_16505,N_14258,N_13600);
xnor U16506 (N_16506,N_14508,N_14899);
nand U16507 (N_16507,N_12796,N_13823);
and U16508 (N_16508,N_14574,N_14339);
nand U16509 (N_16509,N_14940,N_14275);
nand U16510 (N_16510,N_13205,N_14087);
and U16511 (N_16511,N_13693,N_13636);
or U16512 (N_16512,N_13740,N_14703);
nor U16513 (N_16513,N_13464,N_13013);
nor U16514 (N_16514,N_12660,N_12868);
xor U16515 (N_16515,N_14120,N_12644);
nor U16516 (N_16516,N_12827,N_13267);
nor U16517 (N_16517,N_14070,N_13624);
xor U16518 (N_16518,N_12621,N_14038);
nor U16519 (N_16519,N_14262,N_14698);
nor U16520 (N_16520,N_13956,N_14589);
nand U16521 (N_16521,N_12709,N_13013);
nor U16522 (N_16522,N_13546,N_13133);
and U16523 (N_16523,N_13582,N_12519);
and U16524 (N_16524,N_13313,N_12571);
xnor U16525 (N_16525,N_14558,N_14505);
and U16526 (N_16526,N_13470,N_13424);
or U16527 (N_16527,N_13271,N_12697);
and U16528 (N_16528,N_13404,N_14687);
or U16529 (N_16529,N_13005,N_13616);
or U16530 (N_16530,N_13778,N_13676);
and U16531 (N_16531,N_14408,N_14278);
nand U16532 (N_16532,N_13426,N_14729);
and U16533 (N_16533,N_12712,N_13263);
nand U16534 (N_16534,N_14827,N_12652);
or U16535 (N_16535,N_13513,N_12623);
nor U16536 (N_16536,N_13408,N_14095);
and U16537 (N_16537,N_13850,N_13218);
nand U16538 (N_16538,N_14105,N_13051);
and U16539 (N_16539,N_14751,N_14585);
and U16540 (N_16540,N_12583,N_13208);
and U16541 (N_16541,N_13835,N_14722);
and U16542 (N_16542,N_14696,N_13815);
nor U16543 (N_16543,N_14209,N_13872);
nor U16544 (N_16544,N_14527,N_13307);
nand U16545 (N_16545,N_14411,N_12765);
nor U16546 (N_16546,N_12674,N_13834);
or U16547 (N_16547,N_12958,N_14708);
xnor U16548 (N_16548,N_14342,N_14360);
nor U16549 (N_16549,N_13187,N_14847);
and U16550 (N_16550,N_14465,N_14730);
xnor U16551 (N_16551,N_13040,N_14072);
nor U16552 (N_16552,N_14379,N_12749);
nor U16553 (N_16553,N_13523,N_14233);
xnor U16554 (N_16554,N_14132,N_12728);
nor U16555 (N_16555,N_13169,N_13912);
xor U16556 (N_16556,N_14432,N_14545);
or U16557 (N_16557,N_14021,N_13989);
and U16558 (N_16558,N_13940,N_13222);
nand U16559 (N_16559,N_13492,N_14462);
nor U16560 (N_16560,N_12780,N_14893);
nor U16561 (N_16561,N_13694,N_14822);
xnor U16562 (N_16562,N_14951,N_12949);
nand U16563 (N_16563,N_14659,N_12739);
or U16564 (N_16564,N_12790,N_14766);
nor U16565 (N_16565,N_12516,N_14851);
nor U16566 (N_16566,N_14873,N_13289);
or U16567 (N_16567,N_14587,N_13803);
nand U16568 (N_16568,N_13265,N_14385);
and U16569 (N_16569,N_13037,N_13491);
nand U16570 (N_16570,N_13512,N_14371);
xnor U16571 (N_16571,N_14710,N_13969);
nand U16572 (N_16572,N_14430,N_12704);
or U16573 (N_16573,N_13377,N_13660);
or U16574 (N_16574,N_14144,N_12572);
nand U16575 (N_16575,N_14193,N_13786);
nor U16576 (N_16576,N_13216,N_14081);
and U16577 (N_16577,N_13223,N_12778);
or U16578 (N_16578,N_13941,N_14163);
nand U16579 (N_16579,N_14388,N_14167);
nand U16580 (N_16580,N_12945,N_12639);
nand U16581 (N_16581,N_14116,N_14422);
or U16582 (N_16582,N_14485,N_14767);
nand U16583 (N_16583,N_14916,N_12632);
nand U16584 (N_16584,N_14564,N_14856);
nand U16585 (N_16585,N_14305,N_13388);
and U16586 (N_16586,N_13231,N_12914);
xnor U16587 (N_16587,N_14020,N_14587);
xnor U16588 (N_16588,N_13448,N_13055);
nand U16589 (N_16589,N_13157,N_14586);
nand U16590 (N_16590,N_13783,N_12728);
xor U16591 (N_16591,N_13415,N_14424);
xnor U16592 (N_16592,N_14405,N_14684);
nor U16593 (N_16593,N_14530,N_13605);
nor U16594 (N_16594,N_14303,N_12716);
and U16595 (N_16595,N_12725,N_13128);
xnor U16596 (N_16596,N_14395,N_12830);
xnor U16597 (N_16597,N_12972,N_14970);
nor U16598 (N_16598,N_14922,N_13215);
xor U16599 (N_16599,N_14942,N_14520);
nor U16600 (N_16600,N_14023,N_14565);
and U16601 (N_16601,N_14301,N_13813);
nand U16602 (N_16602,N_13637,N_14124);
or U16603 (N_16603,N_12638,N_13074);
nor U16604 (N_16604,N_14065,N_13778);
xnor U16605 (N_16605,N_12626,N_14698);
nand U16606 (N_16606,N_13685,N_13652);
nor U16607 (N_16607,N_13157,N_13321);
nor U16608 (N_16608,N_14555,N_14662);
nor U16609 (N_16609,N_14264,N_12925);
or U16610 (N_16610,N_14812,N_13748);
nand U16611 (N_16611,N_14016,N_13481);
nand U16612 (N_16612,N_14637,N_14701);
nand U16613 (N_16613,N_12764,N_14400);
nand U16614 (N_16614,N_14616,N_13199);
nand U16615 (N_16615,N_13505,N_13391);
nand U16616 (N_16616,N_12726,N_14425);
nor U16617 (N_16617,N_14399,N_13795);
nor U16618 (N_16618,N_13261,N_13946);
nor U16619 (N_16619,N_13965,N_13710);
and U16620 (N_16620,N_14621,N_14435);
and U16621 (N_16621,N_13324,N_13473);
or U16622 (N_16622,N_13009,N_14638);
xor U16623 (N_16623,N_13029,N_13361);
xnor U16624 (N_16624,N_12519,N_14150);
nand U16625 (N_16625,N_13523,N_13059);
nand U16626 (N_16626,N_12714,N_13184);
and U16627 (N_16627,N_14016,N_12535);
nor U16628 (N_16628,N_14471,N_14864);
or U16629 (N_16629,N_14790,N_13518);
or U16630 (N_16630,N_14390,N_14597);
xnor U16631 (N_16631,N_12724,N_14452);
nor U16632 (N_16632,N_13643,N_12806);
xor U16633 (N_16633,N_14160,N_14642);
nor U16634 (N_16634,N_14104,N_14991);
xnor U16635 (N_16635,N_13407,N_13971);
or U16636 (N_16636,N_14250,N_14070);
nor U16637 (N_16637,N_14422,N_12865);
xor U16638 (N_16638,N_12910,N_13333);
and U16639 (N_16639,N_12971,N_14192);
or U16640 (N_16640,N_14794,N_14290);
xor U16641 (N_16641,N_14416,N_13119);
or U16642 (N_16642,N_12641,N_13759);
or U16643 (N_16643,N_14887,N_13322);
or U16644 (N_16644,N_13070,N_14583);
nor U16645 (N_16645,N_13526,N_12876);
nor U16646 (N_16646,N_14167,N_14504);
and U16647 (N_16647,N_14072,N_13087);
nor U16648 (N_16648,N_13861,N_14105);
and U16649 (N_16649,N_14954,N_12882);
or U16650 (N_16650,N_12786,N_14542);
and U16651 (N_16651,N_14121,N_13973);
nand U16652 (N_16652,N_13525,N_13220);
nand U16653 (N_16653,N_13309,N_14859);
and U16654 (N_16654,N_12813,N_13418);
xor U16655 (N_16655,N_13543,N_14417);
xnor U16656 (N_16656,N_14398,N_12834);
and U16657 (N_16657,N_13631,N_14017);
and U16658 (N_16658,N_14593,N_12969);
nand U16659 (N_16659,N_14085,N_14909);
and U16660 (N_16660,N_14700,N_14485);
or U16661 (N_16661,N_12877,N_14544);
or U16662 (N_16662,N_12758,N_14307);
and U16663 (N_16663,N_13768,N_12551);
or U16664 (N_16664,N_13492,N_12782);
or U16665 (N_16665,N_13714,N_14163);
and U16666 (N_16666,N_14793,N_14735);
and U16667 (N_16667,N_13896,N_13441);
nor U16668 (N_16668,N_13674,N_12532);
and U16669 (N_16669,N_14445,N_14990);
xnor U16670 (N_16670,N_14651,N_13526);
nand U16671 (N_16671,N_14902,N_12625);
nor U16672 (N_16672,N_14518,N_14761);
xnor U16673 (N_16673,N_14013,N_13554);
nand U16674 (N_16674,N_14922,N_13204);
and U16675 (N_16675,N_14446,N_14116);
nand U16676 (N_16676,N_13652,N_14796);
nand U16677 (N_16677,N_14467,N_13472);
or U16678 (N_16678,N_13362,N_13173);
nor U16679 (N_16679,N_13666,N_13815);
or U16680 (N_16680,N_14796,N_14007);
xnor U16681 (N_16681,N_13146,N_13836);
xor U16682 (N_16682,N_13072,N_14498);
and U16683 (N_16683,N_13004,N_14311);
xor U16684 (N_16684,N_13429,N_14413);
and U16685 (N_16685,N_13448,N_14783);
xnor U16686 (N_16686,N_13042,N_14100);
and U16687 (N_16687,N_13041,N_12683);
or U16688 (N_16688,N_14502,N_13683);
or U16689 (N_16689,N_14937,N_12895);
nor U16690 (N_16690,N_13176,N_13687);
nand U16691 (N_16691,N_12929,N_13808);
or U16692 (N_16692,N_13652,N_14140);
nand U16693 (N_16693,N_14278,N_14672);
nor U16694 (N_16694,N_12958,N_13847);
nand U16695 (N_16695,N_12905,N_14781);
nor U16696 (N_16696,N_13231,N_13391);
or U16697 (N_16697,N_14339,N_13732);
and U16698 (N_16698,N_13290,N_14847);
xor U16699 (N_16699,N_14755,N_13850);
or U16700 (N_16700,N_13859,N_12592);
or U16701 (N_16701,N_14567,N_14017);
and U16702 (N_16702,N_13610,N_14510);
nand U16703 (N_16703,N_14448,N_14843);
and U16704 (N_16704,N_13401,N_12574);
nor U16705 (N_16705,N_14069,N_12946);
xor U16706 (N_16706,N_14474,N_13895);
nand U16707 (N_16707,N_13119,N_14509);
nand U16708 (N_16708,N_14745,N_12737);
nor U16709 (N_16709,N_14321,N_12875);
or U16710 (N_16710,N_13575,N_13285);
or U16711 (N_16711,N_14822,N_13252);
xor U16712 (N_16712,N_13396,N_12625);
nor U16713 (N_16713,N_13952,N_14537);
nand U16714 (N_16714,N_14469,N_13731);
or U16715 (N_16715,N_14636,N_13734);
and U16716 (N_16716,N_14471,N_14700);
or U16717 (N_16717,N_14699,N_14864);
and U16718 (N_16718,N_14413,N_13479);
nand U16719 (N_16719,N_14404,N_13173);
xnor U16720 (N_16720,N_14821,N_14370);
and U16721 (N_16721,N_13744,N_14476);
or U16722 (N_16722,N_14528,N_13049);
nor U16723 (N_16723,N_14711,N_14381);
nand U16724 (N_16724,N_13713,N_12676);
xor U16725 (N_16725,N_14687,N_13130);
xnor U16726 (N_16726,N_12699,N_12655);
xor U16727 (N_16727,N_13998,N_14582);
nor U16728 (N_16728,N_14349,N_14733);
or U16729 (N_16729,N_14698,N_13826);
xor U16730 (N_16730,N_12860,N_13282);
or U16731 (N_16731,N_13725,N_13747);
nand U16732 (N_16732,N_13552,N_14155);
xnor U16733 (N_16733,N_14323,N_14439);
nand U16734 (N_16734,N_12646,N_13195);
and U16735 (N_16735,N_14274,N_13211);
nor U16736 (N_16736,N_13250,N_13949);
xor U16737 (N_16737,N_14617,N_13932);
nand U16738 (N_16738,N_13129,N_13802);
nor U16739 (N_16739,N_12876,N_14787);
or U16740 (N_16740,N_14383,N_12995);
xor U16741 (N_16741,N_14887,N_13189);
xnor U16742 (N_16742,N_14922,N_14643);
or U16743 (N_16743,N_13476,N_13180);
nor U16744 (N_16744,N_14637,N_13399);
and U16745 (N_16745,N_14379,N_12767);
nor U16746 (N_16746,N_13954,N_13923);
and U16747 (N_16747,N_13018,N_14099);
xor U16748 (N_16748,N_14942,N_13832);
nand U16749 (N_16749,N_14453,N_12793);
xor U16750 (N_16750,N_14331,N_13072);
xnor U16751 (N_16751,N_14329,N_12516);
nand U16752 (N_16752,N_14174,N_14242);
and U16753 (N_16753,N_14498,N_14679);
or U16754 (N_16754,N_14445,N_14151);
and U16755 (N_16755,N_14401,N_14627);
xnor U16756 (N_16756,N_14496,N_13881);
or U16757 (N_16757,N_14390,N_12582);
nand U16758 (N_16758,N_13752,N_13443);
or U16759 (N_16759,N_14026,N_12761);
xor U16760 (N_16760,N_13463,N_14561);
nand U16761 (N_16761,N_13746,N_13160);
and U16762 (N_16762,N_14672,N_13852);
and U16763 (N_16763,N_14275,N_13581);
xnor U16764 (N_16764,N_13711,N_13807);
and U16765 (N_16765,N_14903,N_14832);
xnor U16766 (N_16766,N_14712,N_13970);
or U16767 (N_16767,N_12802,N_13840);
or U16768 (N_16768,N_12675,N_14931);
xnor U16769 (N_16769,N_13762,N_14339);
xnor U16770 (N_16770,N_12606,N_14471);
and U16771 (N_16771,N_12799,N_12657);
and U16772 (N_16772,N_14989,N_12998);
xnor U16773 (N_16773,N_12767,N_12763);
and U16774 (N_16774,N_14070,N_13857);
nor U16775 (N_16775,N_14898,N_13805);
nand U16776 (N_16776,N_14100,N_14460);
xor U16777 (N_16777,N_13348,N_14452);
nand U16778 (N_16778,N_13192,N_12864);
xnor U16779 (N_16779,N_12761,N_13437);
or U16780 (N_16780,N_13260,N_13221);
or U16781 (N_16781,N_13827,N_13993);
xnor U16782 (N_16782,N_13405,N_12829);
or U16783 (N_16783,N_14086,N_14965);
nand U16784 (N_16784,N_13736,N_13933);
and U16785 (N_16785,N_13166,N_14680);
nor U16786 (N_16786,N_13430,N_12665);
xnor U16787 (N_16787,N_12522,N_12934);
and U16788 (N_16788,N_12602,N_13146);
nor U16789 (N_16789,N_14436,N_12531);
or U16790 (N_16790,N_13533,N_13934);
and U16791 (N_16791,N_14368,N_12829);
and U16792 (N_16792,N_14262,N_13236);
xnor U16793 (N_16793,N_14759,N_12733);
or U16794 (N_16794,N_12670,N_13042);
nor U16795 (N_16795,N_14180,N_14126);
or U16796 (N_16796,N_14999,N_13116);
nor U16797 (N_16797,N_13603,N_12681);
xnor U16798 (N_16798,N_14466,N_12670);
or U16799 (N_16799,N_12751,N_12921);
or U16800 (N_16800,N_13764,N_14071);
or U16801 (N_16801,N_12631,N_13850);
nor U16802 (N_16802,N_13993,N_14256);
or U16803 (N_16803,N_13842,N_13393);
or U16804 (N_16804,N_13380,N_13077);
and U16805 (N_16805,N_13747,N_12928);
and U16806 (N_16806,N_13661,N_13194);
and U16807 (N_16807,N_13208,N_13335);
and U16808 (N_16808,N_14491,N_14555);
and U16809 (N_16809,N_13579,N_13153);
or U16810 (N_16810,N_14628,N_14079);
nor U16811 (N_16811,N_14323,N_14749);
or U16812 (N_16812,N_14328,N_14602);
or U16813 (N_16813,N_12717,N_14861);
nand U16814 (N_16814,N_13768,N_14414);
or U16815 (N_16815,N_12784,N_13977);
xnor U16816 (N_16816,N_14519,N_14244);
nand U16817 (N_16817,N_13659,N_14053);
xnor U16818 (N_16818,N_13068,N_14474);
or U16819 (N_16819,N_13688,N_14050);
and U16820 (N_16820,N_14547,N_12517);
xnor U16821 (N_16821,N_13348,N_13007);
or U16822 (N_16822,N_13662,N_13334);
and U16823 (N_16823,N_13193,N_14317);
xnor U16824 (N_16824,N_14341,N_12608);
xor U16825 (N_16825,N_13491,N_12737);
xnor U16826 (N_16826,N_14731,N_14577);
xnor U16827 (N_16827,N_14664,N_12729);
xnor U16828 (N_16828,N_13264,N_12930);
and U16829 (N_16829,N_13171,N_13388);
xnor U16830 (N_16830,N_14329,N_14948);
or U16831 (N_16831,N_13293,N_14019);
nand U16832 (N_16832,N_12880,N_14338);
and U16833 (N_16833,N_14797,N_13525);
nand U16834 (N_16834,N_14467,N_13314);
nand U16835 (N_16835,N_12607,N_13840);
or U16836 (N_16836,N_12746,N_12857);
or U16837 (N_16837,N_13579,N_14270);
or U16838 (N_16838,N_13089,N_13590);
xor U16839 (N_16839,N_12957,N_14542);
xnor U16840 (N_16840,N_14121,N_14389);
nor U16841 (N_16841,N_14821,N_14752);
and U16842 (N_16842,N_13142,N_14099);
xor U16843 (N_16843,N_12548,N_12972);
nand U16844 (N_16844,N_14490,N_14763);
nor U16845 (N_16845,N_12857,N_13048);
and U16846 (N_16846,N_14705,N_14729);
xnor U16847 (N_16847,N_14582,N_14981);
nand U16848 (N_16848,N_14704,N_13563);
nor U16849 (N_16849,N_14648,N_14966);
xnor U16850 (N_16850,N_13604,N_13325);
or U16851 (N_16851,N_12608,N_12731);
nand U16852 (N_16852,N_13037,N_13611);
xnor U16853 (N_16853,N_14982,N_13086);
xnor U16854 (N_16854,N_14418,N_13533);
and U16855 (N_16855,N_12614,N_13666);
nor U16856 (N_16856,N_13966,N_14651);
and U16857 (N_16857,N_13685,N_13407);
nor U16858 (N_16858,N_13695,N_14260);
nor U16859 (N_16859,N_12580,N_12823);
nor U16860 (N_16860,N_14842,N_13225);
nand U16861 (N_16861,N_13153,N_12661);
nand U16862 (N_16862,N_14451,N_13978);
and U16863 (N_16863,N_14612,N_12886);
xor U16864 (N_16864,N_13299,N_12543);
nor U16865 (N_16865,N_13765,N_12739);
nand U16866 (N_16866,N_14693,N_14169);
nand U16867 (N_16867,N_14172,N_14102);
nand U16868 (N_16868,N_14208,N_14953);
or U16869 (N_16869,N_12545,N_13184);
nor U16870 (N_16870,N_14250,N_13693);
and U16871 (N_16871,N_13690,N_13267);
nand U16872 (N_16872,N_14344,N_14625);
or U16873 (N_16873,N_13389,N_14009);
xor U16874 (N_16874,N_13206,N_12637);
xnor U16875 (N_16875,N_14149,N_14173);
nor U16876 (N_16876,N_12723,N_14694);
and U16877 (N_16877,N_14879,N_14583);
and U16878 (N_16878,N_12550,N_13062);
and U16879 (N_16879,N_14351,N_12558);
or U16880 (N_16880,N_14186,N_13222);
xnor U16881 (N_16881,N_13877,N_14466);
xnor U16882 (N_16882,N_14412,N_13235);
or U16883 (N_16883,N_13351,N_13651);
xor U16884 (N_16884,N_13593,N_13795);
nand U16885 (N_16885,N_12774,N_14436);
nand U16886 (N_16886,N_12826,N_12688);
nand U16887 (N_16887,N_13470,N_14117);
nor U16888 (N_16888,N_14405,N_14120);
or U16889 (N_16889,N_14795,N_14494);
xor U16890 (N_16890,N_14369,N_14228);
xor U16891 (N_16891,N_14721,N_14344);
nor U16892 (N_16892,N_13734,N_14653);
and U16893 (N_16893,N_13308,N_14577);
nand U16894 (N_16894,N_12952,N_14772);
xnor U16895 (N_16895,N_14739,N_14192);
xnor U16896 (N_16896,N_14372,N_14475);
or U16897 (N_16897,N_12763,N_14789);
nor U16898 (N_16898,N_13164,N_13813);
nor U16899 (N_16899,N_14164,N_12947);
or U16900 (N_16900,N_13181,N_13824);
nor U16901 (N_16901,N_14112,N_14647);
nor U16902 (N_16902,N_14413,N_14480);
and U16903 (N_16903,N_13809,N_13762);
xor U16904 (N_16904,N_14111,N_12754);
or U16905 (N_16905,N_14349,N_13966);
and U16906 (N_16906,N_12739,N_14616);
nand U16907 (N_16907,N_13376,N_13047);
xnor U16908 (N_16908,N_13566,N_12645);
nand U16909 (N_16909,N_13464,N_13511);
and U16910 (N_16910,N_14662,N_12995);
xnor U16911 (N_16911,N_14388,N_12650);
or U16912 (N_16912,N_13972,N_12745);
and U16913 (N_16913,N_13060,N_12911);
nor U16914 (N_16914,N_12539,N_14250);
and U16915 (N_16915,N_14665,N_12849);
xor U16916 (N_16916,N_14724,N_13187);
and U16917 (N_16917,N_14637,N_14476);
and U16918 (N_16918,N_13350,N_13382);
and U16919 (N_16919,N_14752,N_13445);
nand U16920 (N_16920,N_12621,N_12931);
and U16921 (N_16921,N_13718,N_12977);
nand U16922 (N_16922,N_12699,N_12507);
xnor U16923 (N_16923,N_14637,N_14323);
or U16924 (N_16924,N_12583,N_14011);
nand U16925 (N_16925,N_12735,N_14236);
xnor U16926 (N_16926,N_13089,N_14584);
or U16927 (N_16927,N_13926,N_14176);
nand U16928 (N_16928,N_14536,N_14834);
and U16929 (N_16929,N_13340,N_12711);
and U16930 (N_16930,N_13981,N_13999);
xor U16931 (N_16931,N_12807,N_14399);
nor U16932 (N_16932,N_12724,N_13276);
nand U16933 (N_16933,N_14584,N_12887);
or U16934 (N_16934,N_13647,N_13023);
nor U16935 (N_16935,N_13230,N_13667);
or U16936 (N_16936,N_12535,N_14619);
nand U16937 (N_16937,N_13764,N_12923);
or U16938 (N_16938,N_13712,N_12772);
xnor U16939 (N_16939,N_13213,N_13359);
or U16940 (N_16940,N_14886,N_13730);
xnor U16941 (N_16941,N_14440,N_13301);
nor U16942 (N_16942,N_12692,N_13804);
and U16943 (N_16943,N_14510,N_12855);
nor U16944 (N_16944,N_14564,N_14109);
nand U16945 (N_16945,N_12793,N_12686);
and U16946 (N_16946,N_13707,N_12911);
xor U16947 (N_16947,N_12772,N_13907);
or U16948 (N_16948,N_14386,N_13165);
nand U16949 (N_16949,N_14857,N_13951);
and U16950 (N_16950,N_14455,N_13707);
nor U16951 (N_16951,N_13598,N_12922);
nor U16952 (N_16952,N_13946,N_14565);
nor U16953 (N_16953,N_14456,N_14659);
nand U16954 (N_16954,N_14574,N_14005);
nand U16955 (N_16955,N_13398,N_14623);
or U16956 (N_16956,N_14170,N_14945);
nor U16957 (N_16957,N_14455,N_14308);
xnor U16958 (N_16958,N_14385,N_14748);
nand U16959 (N_16959,N_14715,N_13489);
or U16960 (N_16960,N_12545,N_12722);
or U16961 (N_16961,N_14166,N_14295);
nor U16962 (N_16962,N_14089,N_12979);
xor U16963 (N_16963,N_14714,N_12914);
xor U16964 (N_16964,N_14929,N_14785);
xor U16965 (N_16965,N_14553,N_14120);
or U16966 (N_16966,N_13111,N_14018);
nor U16967 (N_16967,N_14636,N_12958);
nor U16968 (N_16968,N_13905,N_13692);
or U16969 (N_16969,N_12590,N_12901);
nand U16970 (N_16970,N_14535,N_14171);
or U16971 (N_16971,N_14151,N_13340);
xor U16972 (N_16972,N_13305,N_13251);
and U16973 (N_16973,N_13861,N_12846);
xnor U16974 (N_16974,N_12606,N_13969);
nor U16975 (N_16975,N_13243,N_14340);
xor U16976 (N_16976,N_14189,N_12780);
nor U16977 (N_16977,N_14838,N_14166);
and U16978 (N_16978,N_14101,N_14982);
and U16979 (N_16979,N_13117,N_13483);
nand U16980 (N_16980,N_14082,N_12776);
nand U16981 (N_16981,N_13807,N_14532);
and U16982 (N_16982,N_13807,N_12605);
and U16983 (N_16983,N_12645,N_13447);
or U16984 (N_16984,N_14693,N_14171);
or U16985 (N_16985,N_13863,N_14205);
and U16986 (N_16986,N_13611,N_14134);
xor U16987 (N_16987,N_14580,N_14524);
xnor U16988 (N_16988,N_14275,N_14258);
nand U16989 (N_16989,N_12851,N_13137);
xnor U16990 (N_16990,N_14222,N_14215);
nor U16991 (N_16991,N_13195,N_14995);
xor U16992 (N_16992,N_13407,N_14815);
nand U16993 (N_16993,N_12807,N_13879);
or U16994 (N_16994,N_12833,N_13773);
xnor U16995 (N_16995,N_14143,N_12966);
nand U16996 (N_16996,N_13897,N_14755);
or U16997 (N_16997,N_13191,N_14776);
or U16998 (N_16998,N_14451,N_14639);
or U16999 (N_16999,N_12532,N_13811);
or U17000 (N_17000,N_14761,N_13598);
and U17001 (N_17001,N_13304,N_12809);
and U17002 (N_17002,N_13607,N_14204);
nand U17003 (N_17003,N_13629,N_14863);
xnor U17004 (N_17004,N_14403,N_12988);
nand U17005 (N_17005,N_14798,N_14846);
xnor U17006 (N_17006,N_14466,N_13388);
and U17007 (N_17007,N_14178,N_13026);
nand U17008 (N_17008,N_13704,N_13538);
or U17009 (N_17009,N_14628,N_13445);
xnor U17010 (N_17010,N_12733,N_14252);
and U17011 (N_17011,N_12688,N_14579);
and U17012 (N_17012,N_13381,N_14737);
or U17013 (N_17013,N_13613,N_12587);
or U17014 (N_17014,N_13780,N_13766);
and U17015 (N_17015,N_13216,N_14118);
nand U17016 (N_17016,N_13069,N_13937);
and U17017 (N_17017,N_14442,N_14329);
and U17018 (N_17018,N_13558,N_14029);
nor U17019 (N_17019,N_13323,N_12545);
or U17020 (N_17020,N_14832,N_14270);
or U17021 (N_17021,N_13223,N_13996);
or U17022 (N_17022,N_13609,N_13912);
nor U17023 (N_17023,N_13344,N_12786);
and U17024 (N_17024,N_13572,N_14801);
nor U17025 (N_17025,N_13247,N_14458);
nand U17026 (N_17026,N_14590,N_13414);
nand U17027 (N_17027,N_14315,N_14098);
xor U17028 (N_17028,N_12829,N_14033);
and U17029 (N_17029,N_13888,N_13900);
nor U17030 (N_17030,N_13185,N_13551);
nand U17031 (N_17031,N_14577,N_14427);
nand U17032 (N_17032,N_14517,N_12876);
or U17033 (N_17033,N_13308,N_14549);
xor U17034 (N_17034,N_14098,N_14947);
nor U17035 (N_17035,N_13296,N_12515);
nand U17036 (N_17036,N_14206,N_13131);
and U17037 (N_17037,N_12856,N_13372);
or U17038 (N_17038,N_13676,N_13225);
or U17039 (N_17039,N_14546,N_12560);
nor U17040 (N_17040,N_14047,N_13426);
nor U17041 (N_17041,N_12854,N_14524);
or U17042 (N_17042,N_14519,N_13217);
nor U17043 (N_17043,N_14860,N_13516);
or U17044 (N_17044,N_14436,N_12711);
nand U17045 (N_17045,N_14489,N_12688);
and U17046 (N_17046,N_13969,N_14976);
or U17047 (N_17047,N_12607,N_14863);
nand U17048 (N_17048,N_13087,N_12623);
and U17049 (N_17049,N_14952,N_13556);
and U17050 (N_17050,N_12758,N_14643);
nand U17051 (N_17051,N_12984,N_13940);
xor U17052 (N_17052,N_13597,N_12527);
xor U17053 (N_17053,N_13706,N_13251);
nand U17054 (N_17054,N_13120,N_13539);
nand U17055 (N_17055,N_14164,N_14347);
or U17056 (N_17056,N_14883,N_14386);
and U17057 (N_17057,N_14768,N_12857);
and U17058 (N_17058,N_13355,N_14382);
nor U17059 (N_17059,N_13603,N_13137);
xnor U17060 (N_17060,N_14176,N_12831);
or U17061 (N_17061,N_14514,N_14256);
or U17062 (N_17062,N_13399,N_14420);
or U17063 (N_17063,N_12685,N_14878);
or U17064 (N_17064,N_13155,N_13034);
nand U17065 (N_17065,N_14537,N_13053);
xnor U17066 (N_17066,N_13688,N_14946);
or U17067 (N_17067,N_13738,N_13520);
and U17068 (N_17068,N_13338,N_13372);
or U17069 (N_17069,N_14458,N_14000);
xnor U17070 (N_17070,N_14550,N_12800);
nor U17071 (N_17071,N_12924,N_13168);
nand U17072 (N_17072,N_13677,N_14863);
xnor U17073 (N_17073,N_13423,N_13288);
nand U17074 (N_17074,N_13456,N_12920);
nand U17075 (N_17075,N_14611,N_13179);
or U17076 (N_17076,N_14837,N_14116);
nand U17077 (N_17077,N_13957,N_13404);
or U17078 (N_17078,N_14819,N_13889);
or U17079 (N_17079,N_13833,N_14061);
or U17080 (N_17080,N_14757,N_13693);
nor U17081 (N_17081,N_14531,N_14956);
nand U17082 (N_17082,N_12674,N_14636);
and U17083 (N_17083,N_12802,N_14213);
nor U17084 (N_17084,N_13974,N_13236);
nor U17085 (N_17085,N_12525,N_14558);
or U17086 (N_17086,N_13222,N_13468);
nor U17087 (N_17087,N_13539,N_12615);
or U17088 (N_17088,N_13191,N_12904);
and U17089 (N_17089,N_14407,N_13390);
and U17090 (N_17090,N_14530,N_12958);
xnor U17091 (N_17091,N_14416,N_13521);
nor U17092 (N_17092,N_14512,N_13232);
xnor U17093 (N_17093,N_12640,N_13391);
nand U17094 (N_17094,N_13629,N_14749);
or U17095 (N_17095,N_13317,N_13973);
nor U17096 (N_17096,N_14959,N_14371);
and U17097 (N_17097,N_13862,N_13361);
nand U17098 (N_17098,N_13931,N_13340);
nor U17099 (N_17099,N_13639,N_12986);
xnor U17100 (N_17100,N_14053,N_13490);
nor U17101 (N_17101,N_14913,N_12710);
nand U17102 (N_17102,N_14569,N_12655);
or U17103 (N_17103,N_12838,N_14181);
nand U17104 (N_17104,N_14253,N_14934);
or U17105 (N_17105,N_12868,N_13331);
nand U17106 (N_17106,N_14395,N_13506);
xor U17107 (N_17107,N_12739,N_14576);
and U17108 (N_17108,N_14115,N_14722);
xnor U17109 (N_17109,N_13289,N_13355);
nor U17110 (N_17110,N_13819,N_13686);
nor U17111 (N_17111,N_14408,N_13761);
and U17112 (N_17112,N_14758,N_12745);
and U17113 (N_17113,N_14960,N_13454);
xor U17114 (N_17114,N_13964,N_13311);
nand U17115 (N_17115,N_14685,N_14281);
and U17116 (N_17116,N_13283,N_14550);
xnor U17117 (N_17117,N_13922,N_14708);
or U17118 (N_17118,N_14265,N_13461);
nand U17119 (N_17119,N_14429,N_14270);
nor U17120 (N_17120,N_14154,N_12968);
nor U17121 (N_17121,N_14511,N_13606);
or U17122 (N_17122,N_12603,N_13373);
or U17123 (N_17123,N_13122,N_13539);
xor U17124 (N_17124,N_13778,N_12727);
and U17125 (N_17125,N_12619,N_14954);
and U17126 (N_17126,N_14932,N_14628);
nand U17127 (N_17127,N_13337,N_14901);
and U17128 (N_17128,N_12787,N_14188);
xnor U17129 (N_17129,N_14693,N_12953);
nand U17130 (N_17130,N_12940,N_12971);
nand U17131 (N_17131,N_13613,N_14383);
xor U17132 (N_17132,N_12973,N_14468);
nor U17133 (N_17133,N_14928,N_13678);
or U17134 (N_17134,N_14896,N_13868);
xnor U17135 (N_17135,N_12822,N_13565);
nor U17136 (N_17136,N_12878,N_12941);
nor U17137 (N_17137,N_13307,N_14405);
xor U17138 (N_17138,N_13040,N_14012);
xnor U17139 (N_17139,N_14137,N_13621);
nand U17140 (N_17140,N_14072,N_13687);
xnor U17141 (N_17141,N_12695,N_14131);
or U17142 (N_17142,N_13702,N_14107);
or U17143 (N_17143,N_13220,N_13694);
or U17144 (N_17144,N_13675,N_13321);
and U17145 (N_17145,N_14051,N_14724);
nor U17146 (N_17146,N_12892,N_12765);
nand U17147 (N_17147,N_12983,N_13042);
xor U17148 (N_17148,N_13104,N_12652);
nor U17149 (N_17149,N_14534,N_13665);
or U17150 (N_17150,N_13982,N_14792);
or U17151 (N_17151,N_13941,N_14502);
and U17152 (N_17152,N_13275,N_14658);
or U17153 (N_17153,N_14738,N_14466);
nor U17154 (N_17154,N_13118,N_13621);
or U17155 (N_17155,N_12881,N_14288);
and U17156 (N_17156,N_12881,N_13970);
nor U17157 (N_17157,N_12650,N_14409);
nand U17158 (N_17158,N_13533,N_13765);
or U17159 (N_17159,N_13107,N_14234);
xnor U17160 (N_17160,N_13088,N_13062);
nor U17161 (N_17161,N_13875,N_14332);
xnor U17162 (N_17162,N_14463,N_14588);
nor U17163 (N_17163,N_12841,N_14339);
and U17164 (N_17164,N_13598,N_14240);
nand U17165 (N_17165,N_12787,N_14849);
xor U17166 (N_17166,N_12882,N_14432);
and U17167 (N_17167,N_13097,N_14857);
and U17168 (N_17168,N_12890,N_14023);
nand U17169 (N_17169,N_13826,N_12812);
nand U17170 (N_17170,N_14989,N_13262);
and U17171 (N_17171,N_13689,N_13746);
nor U17172 (N_17172,N_14384,N_13450);
and U17173 (N_17173,N_12762,N_14329);
and U17174 (N_17174,N_13432,N_12935);
or U17175 (N_17175,N_13368,N_14355);
xor U17176 (N_17176,N_12625,N_14832);
and U17177 (N_17177,N_14629,N_13565);
nor U17178 (N_17178,N_14893,N_13363);
nand U17179 (N_17179,N_13569,N_14273);
or U17180 (N_17180,N_14505,N_13085);
nor U17181 (N_17181,N_13751,N_14036);
nand U17182 (N_17182,N_14859,N_14441);
xor U17183 (N_17183,N_13312,N_14677);
nor U17184 (N_17184,N_12697,N_12999);
xor U17185 (N_17185,N_14072,N_14069);
and U17186 (N_17186,N_14294,N_13713);
xnor U17187 (N_17187,N_13186,N_14130);
xnor U17188 (N_17188,N_13174,N_12676);
nor U17189 (N_17189,N_14028,N_14088);
or U17190 (N_17190,N_14459,N_13773);
xnor U17191 (N_17191,N_12558,N_12726);
or U17192 (N_17192,N_13374,N_12679);
nor U17193 (N_17193,N_12949,N_14484);
xor U17194 (N_17194,N_14232,N_13014);
xnor U17195 (N_17195,N_13285,N_13266);
nor U17196 (N_17196,N_14586,N_13180);
nor U17197 (N_17197,N_13422,N_13552);
xor U17198 (N_17198,N_12847,N_13492);
nor U17199 (N_17199,N_14071,N_13771);
or U17200 (N_17200,N_14631,N_13763);
nor U17201 (N_17201,N_13877,N_13907);
and U17202 (N_17202,N_13862,N_12783);
nand U17203 (N_17203,N_14528,N_13254);
and U17204 (N_17204,N_14949,N_12542);
or U17205 (N_17205,N_13027,N_12810);
or U17206 (N_17206,N_12637,N_14818);
nor U17207 (N_17207,N_13456,N_14065);
or U17208 (N_17208,N_14920,N_13135);
nand U17209 (N_17209,N_14498,N_14011);
nor U17210 (N_17210,N_13252,N_13892);
and U17211 (N_17211,N_14012,N_14441);
xor U17212 (N_17212,N_13870,N_13522);
or U17213 (N_17213,N_14525,N_13476);
nor U17214 (N_17214,N_13151,N_13331);
or U17215 (N_17215,N_13906,N_13535);
and U17216 (N_17216,N_12839,N_13055);
and U17217 (N_17217,N_14164,N_14079);
and U17218 (N_17218,N_13460,N_14168);
nor U17219 (N_17219,N_14963,N_12912);
xnor U17220 (N_17220,N_14029,N_12596);
nand U17221 (N_17221,N_13643,N_14611);
xor U17222 (N_17222,N_13039,N_13499);
nor U17223 (N_17223,N_14044,N_14375);
and U17224 (N_17224,N_12912,N_13492);
xor U17225 (N_17225,N_14655,N_13449);
nor U17226 (N_17226,N_13252,N_13482);
nand U17227 (N_17227,N_14033,N_14556);
nand U17228 (N_17228,N_12798,N_13342);
and U17229 (N_17229,N_13844,N_12782);
and U17230 (N_17230,N_14447,N_13803);
and U17231 (N_17231,N_12783,N_13505);
or U17232 (N_17232,N_12640,N_13958);
xnor U17233 (N_17233,N_12514,N_13756);
nand U17234 (N_17234,N_13856,N_12567);
or U17235 (N_17235,N_14511,N_14526);
xor U17236 (N_17236,N_13677,N_13992);
xor U17237 (N_17237,N_13560,N_13037);
nand U17238 (N_17238,N_14951,N_14434);
nand U17239 (N_17239,N_14962,N_13812);
nand U17240 (N_17240,N_13712,N_13674);
nor U17241 (N_17241,N_14588,N_14608);
and U17242 (N_17242,N_14435,N_14320);
xor U17243 (N_17243,N_12737,N_13195);
and U17244 (N_17244,N_13867,N_13750);
or U17245 (N_17245,N_13738,N_14264);
and U17246 (N_17246,N_14516,N_14517);
nor U17247 (N_17247,N_13069,N_14746);
xnor U17248 (N_17248,N_14380,N_13455);
or U17249 (N_17249,N_13706,N_13608);
nor U17250 (N_17250,N_12847,N_14092);
nand U17251 (N_17251,N_14567,N_14298);
xnor U17252 (N_17252,N_14778,N_13096);
nor U17253 (N_17253,N_12504,N_14492);
nor U17254 (N_17254,N_13463,N_12844);
xor U17255 (N_17255,N_13391,N_12959);
or U17256 (N_17256,N_13634,N_13057);
nor U17257 (N_17257,N_14693,N_13406);
nor U17258 (N_17258,N_14337,N_14345);
or U17259 (N_17259,N_13795,N_14934);
and U17260 (N_17260,N_14575,N_14688);
nor U17261 (N_17261,N_14290,N_13330);
nor U17262 (N_17262,N_13934,N_13257);
and U17263 (N_17263,N_14806,N_14047);
or U17264 (N_17264,N_13319,N_13374);
xnor U17265 (N_17265,N_14583,N_14923);
nand U17266 (N_17266,N_12817,N_12733);
nand U17267 (N_17267,N_12767,N_13538);
nand U17268 (N_17268,N_12697,N_12526);
xor U17269 (N_17269,N_13651,N_14849);
xor U17270 (N_17270,N_12768,N_14199);
xnor U17271 (N_17271,N_14523,N_12895);
xnor U17272 (N_17272,N_13893,N_14590);
and U17273 (N_17273,N_12555,N_14089);
xnor U17274 (N_17274,N_14527,N_13695);
nand U17275 (N_17275,N_13506,N_13308);
xor U17276 (N_17276,N_12572,N_12898);
nand U17277 (N_17277,N_14313,N_14423);
nand U17278 (N_17278,N_12677,N_13656);
nand U17279 (N_17279,N_13553,N_14207);
and U17280 (N_17280,N_12957,N_14568);
and U17281 (N_17281,N_14981,N_14473);
and U17282 (N_17282,N_12765,N_13328);
or U17283 (N_17283,N_14844,N_13610);
nor U17284 (N_17284,N_14706,N_13806);
and U17285 (N_17285,N_12988,N_14422);
and U17286 (N_17286,N_14743,N_13353);
xnor U17287 (N_17287,N_14904,N_13926);
xor U17288 (N_17288,N_13202,N_13065);
and U17289 (N_17289,N_14760,N_12512);
or U17290 (N_17290,N_12664,N_13271);
nand U17291 (N_17291,N_12588,N_13864);
or U17292 (N_17292,N_14125,N_13708);
xor U17293 (N_17293,N_12687,N_12799);
nor U17294 (N_17294,N_13037,N_14549);
or U17295 (N_17295,N_13626,N_14109);
and U17296 (N_17296,N_13394,N_13617);
and U17297 (N_17297,N_14448,N_14101);
xor U17298 (N_17298,N_13247,N_14757);
xnor U17299 (N_17299,N_13753,N_13253);
or U17300 (N_17300,N_14704,N_13069);
xor U17301 (N_17301,N_12548,N_12542);
nor U17302 (N_17302,N_13269,N_13514);
nor U17303 (N_17303,N_13702,N_12771);
or U17304 (N_17304,N_13852,N_13208);
nor U17305 (N_17305,N_13623,N_14504);
nor U17306 (N_17306,N_13757,N_14973);
and U17307 (N_17307,N_14099,N_13615);
or U17308 (N_17308,N_12679,N_14269);
nor U17309 (N_17309,N_14275,N_14572);
xnor U17310 (N_17310,N_14747,N_13710);
and U17311 (N_17311,N_14919,N_13586);
or U17312 (N_17312,N_12631,N_14152);
nor U17313 (N_17313,N_13517,N_12872);
nor U17314 (N_17314,N_14615,N_12779);
xnor U17315 (N_17315,N_12844,N_14829);
xor U17316 (N_17316,N_14607,N_14303);
or U17317 (N_17317,N_14070,N_12628);
and U17318 (N_17318,N_14142,N_13049);
or U17319 (N_17319,N_14019,N_13031);
and U17320 (N_17320,N_14459,N_14377);
xnor U17321 (N_17321,N_14509,N_12815);
or U17322 (N_17322,N_13303,N_14401);
nor U17323 (N_17323,N_14404,N_13141);
and U17324 (N_17324,N_13611,N_14530);
and U17325 (N_17325,N_14104,N_14186);
or U17326 (N_17326,N_14648,N_12563);
xor U17327 (N_17327,N_13965,N_14564);
and U17328 (N_17328,N_14398,N_13915);
nor U17329 (N_17329,N_13555,N_13855);
nor U17330 (N_17330,N_13452,N_13464);
or U17331 (N_17331,N_13234,N_14823);
and U17332 (N_17332,N_13054,N_13456);
nor U17333 (N_17333,N_14569,N_14437);
and U17334 (N_17334,N_13089,N_14846);
or U17335 (N_17335,N_12909,N_14138);
xnor U17336 (N_17336,N_13120,N_13607);
xor U17337 (N_17337,N_13293,N_14457);
or U17338 (N_17338,N_14632,N_14899);
or U17339 (N_17339,N_14019,N_13241);
xnor U17340 (N_17340,N_12717,N_14177);
or U17341 (N_17341,N_13246,N_12739);
nor U17342 (N_17342,N_13177,N_14915);
nand U17343 (N_17343,N_13739,N_14658);
xnor U17344 (N_17344,N_12732,N_14912);
nor U17345 (N_17345,N_14774,N_14994);
and U17346 (N_17346,N_14974,N_14411);
and U17347 (N_17347,N_12695,N_13743);
nand U17348 (N_17348,N_13067,N_13589);
nand U17349 (N_17349,N_14562,N_14172);
and U17350 (N_17350,N_13451,N_13687);
xor U17351 (N_17351,N_14773,N_14631);
or U17352 (N_17352,N_13912,N_12802);
xor U17353 (N_17353,N_13312,N_12871);
nor U17354 (N_17354,N_13153,N_13986);
nand U17355 (N_17355,N_13489,N_14013);
xnor U17356 (N_17356,N_14784,N_13595);
nor U17357 (N_17357,N_13245,N_14319);
xor U17358 (N_17358,N_13358,N_13089);
nand U17359 (N_17359,N_13242,N_13295);
nor U17360 (N_17360,N_14480,N_13233);
and U17361 (N_17361,N_13822,N_13214);
nand U17362 (N_17362,N_14134,N_13527);
nand U17363 (N_17363,N_13261,N_13501);
nand U17364 (N_17364,N_13289,N_13551);
xor U17365 (N_17365,N_14396,N_13885);
nand U17366 (N_17366,N_13360,N_13236);
and U17367 (N_17367,N_12515,N_14663);
nand U17368 (N_17368,N_14582,N_14337);
or U17369 (N_17369,N_13359,N_14987);
xor U17370 (N_17370,N_12975,N_14817);
xor U17371 (N_17371,N_14186,N_14316);
nand U17372 (N_17372,N_13966,N_12510);
or U17373 (N_17373,N_12961,N_14493);
nand U17374 (N_17374,N_14017,N_14292);
or U17375 (N_17375,N_14843,N_13012);
xor U17376 (N_17376,N_12718,N_13581);
nand U17377 (N_17377,N_13579,N_13697);
or U17378 (N_17378,N_13025,N_14429);
and U17379 (N_17379,N_12965,N_13488);
and U17380 (N_17380,N_14879,N_13313);
xnor U17381 (N_17381,N_12853,N_14665);
xor U17382 (N_17382,N_12973,N_13196);
nor U17383 (N_17383,N_14025,N_14018);
and U17384 (N_17384,N_12779,N_14866);
and U17385 (N_17385,N_13380,N_13397);
and U17386 (N_17386,N_14618,N_13497);
nand U17387 (N_17387,N_13356,N_14557);
and U17388 (N_17388,N_14234,N_13063);
nand U17389 (N_17389,N_14203,N_12807);
nor U17390 (N_17390,N_13104,N_12733);
or U17391 (N_17391,N_14211,N_12983);
and U17392 (N_17392,N_14274,N_13304);
xnor U17393 (N_17393,N_13956,N_14534);
xor U17394 (N_17394,N_12958,N_13571);
and U17395 (N_17395,N_14693,N_13380);
xnor U17396 (N_17396,N_12656,N_14505);
xor U17397 (N_17397,N_13121,N_12673);
and U17398 (N_17398,N_13728,N_14284);
or U17399 (N_17399,N_13321,N_14412);
xor U17400 (N_17400,N_12597,N_12724);
nor U17401 (N_17401,N_12580,N_12627);
and U17402 (N_17402,N_12610,N_13339);
xnor U17403 (N_17403,N_13675,N_14646);
xnor U17404 (N_17404,N_13715,N_14135);
nand U17405 (N_17405,N_13152,N_14684);
nor U17406 (N_17406,N_14715,N_12500);
xnor U17407 (N_17407,N_13445,N_13157);
or U17408 (N_17408,N_14336,N_12912);
or U17409 (N_17409,N_14539,N_14803);
nand U17410 (N_17410,N_14556,N_14500);
and U17411 (N_17411,N_12966,N_13145);
nor U17412 (N_17412,N_13327,N_13377);
or U17413 (N_17413,N_14100,N_13763);
nand U17414 (N_17414,N_13769,N_14149);
and U17415 (N_17415,N_13677,N_14036);
and U17416 (N_17416,N_13493,N_14359);
nand U17417 (N_17417,N_14410,N_12959);
nand U17418 (N_17418,N_14574,N_13620);
xnor U17419 (N_17419,N_13359,N_13773);
nand U17420 (N_17420,N_14907,N_14287);
or U17421 (N_17421,N_14043,N_14347);
and U17422 (N_17422,N_14175,N_14931);
xor U17423 (N_17423,N_12864,N_13225);
nand U17424 (N_17424,N_13888,N_14583);
nand U17425 (N_17425,N_12663,N_13090);
xor U17426 (N_17426,N_14506,N_13625);
nand U17427 (N_17427,N_13253,N_12966);
xor U17428 (N_17428,N_14093,N_13817);
xnor U17429 (N_17429,N_14122,N_14896);
xnor U17430 (N_17430,N_12994,N_12535);
nand U17431 (N_17431,N_14878,N_14252);
nor U17432 (N_17432,N_14078,N_14464);
xnor U17433 (N_17433,N_13190,N_14236);
nand U17434 (N_17434,N_12770,N_13702);
xor U17435 (N_17435,N_14040,N_13956);
and U17436 (N_17436,N_13649,N_14079);
xnor U17437 (N_17437,N_13737,N_12809);
or U17438 (N_17438,N_12920,N_12659);
nand U17439 (N_17439,N_14142,N_14490);
nor U17440 (N_17440,N_14831,N_14423);
nand U17441 (N_17441,N_14512,N_12832);
or U17442 (N_17442,N_12902,N_14775);
xor U17443 (N_17443,N_13759,N_14636);
or U17444 (N_17444,N_13868,N_13723);
nand U17445 (N_17445,N_13143,N_13874);
and U17446 (N_17446,N_13505,N_14189);
nor U17447 (N_17447,N_14510,N_13645);
nor U17448 (N_17448,N_13527,N_14008);
and U17449 (N_17449,N_14487,N_14038);
or U17450 (N_17450,N_14912,N_14463);
xor U17451 (N_17451,N_14878,N_14677);
xor U17452 (N_17452,N_14140,N_14629);
nor U17453 (N_17453,N_14786,N_14230);
xnor U17454 (N_17454,N_13547,N_14131);
and U17455 (N_17455,N_14575,N_14296);
nand U17456 (N_17456,N_14585,N_14503);
nor U17457 (N_17457,N_14513,N_13735);
xor U17458 (N_17458,N_14250,N_13433);
or U17459 (N_17459,N_14546,N_13580);
or U17460 (N_17460,N_14307,N_12510);
nor U17461 (N_17461,N_14213,N_13327);
xnor U17462 (N_17462,N_13746,N_13811);
nor U17463 (N_17463,N_14983,N_13392);
xor U17464 (N_17464,N_13484,N_13791);
xor U17465 (N_17465,N_14928,N_14124);
xnor U17466 (N_17466,N_13020,N_14290);
and U17467 (N_17467,N_14724,N_14524);
or U17468 (N_17468,N_12540,N_13020);
or U17469 (N_17469,N_14139,N_13982);
and U17470 (N_17470,N_13511,N_14206);
or U17471 (N_17471,N_12531,N_13562);
xnor U17472 (N_17472,N_13964,N_14815);
nor U17473 (N_17473,N_13221,N_12707);
nand U17474 (N_17474,N_13819,N_13280);
nor U17475 (N_17475,N_13903,N_13046);
xnor U17476 (N_17476,N_13977,N_12525);
nor U17477 (N_17477,N_13607,N_12506);
nor U17478 (N_17478,N_12861,N_14391);
nand U17479 (N_17479,N_13600,N_12608);
nand U17480 (N_17480,N_13607,N_13229);
nand U17481 (N_17481,N_14807,N_14205);
xor U17482 (N_17482,N_13054,N_13689);
or U17483 (N_17483,N_13721,N_13740);
xnor U17484 (N_17484,N_14967,N_14179);
or U17485 (N_17485,N_14602,N_14542);
xor U17486 (N_17486,N_14530,N_14051);
nor U17487 (N_17487,N_13986,N_12939);
xor U17488 (N_17488,N_12916,N_12628);
nor U17489 (N_17489,N_13471,N_14512);
and U17490 (N_17490,N_12524,N_13953);
and U17491 (N_17491,N_13759,N_12686);
nor U17492 (N_17492,N_13320,N_13684);
and U17493 (N_17493,N_14457,N_14534);
xor U17494 (N_17494,N_14268,N_14076);
or U17495 (N_17495,N_14690,N_13815);
nand U17496 (N_17496,N_14869,N_14448);
xnor U17497 (N_17497,N_14784,N_13522);
or U17498 (N_17498,N_14253,N_14867);
nor U17499 (N_17499,N_13607,N_14702);
or U17500 (N_17500,N_16540,N_17427);
xnor U17501 (N_17501,N_16053,N_15623);
or U17502 (N_17502,N_15632,N_16311);
or U17503 (N_17503,N_16713,N_17183);
xnor U17504 (N_17504,N_16964,N_17310);
and U17505 (N_17505,N_15870,N_16161);
and U17506 (N_17506,N_16878,N_17385);
nor U17507 (N_17507,N_15101,N_15295);
nor U17508 (N_17508,N_16467,N_17271);
and U17509 (N_17509,N_17285,N_16308);
or U17510 (N_17510,N_17395,N_16668);
nor U17511 (N_17511,N_15279,N_16427);
and U17512 (N_17512,N_15495,N_15529);
or U17513 (N_17513,N_17269,N_15386);
nor U17514 (N_17514,N_17371,N_17067);
and U17515 (N_17515,N_16814,N_15949);
nor U17516 (N_17516,N_15210,N_17139);
nor U17517 (N_17517,N_15263,N_17042);
xor U17518 (N_17518,N_15687,N_16709);
xnor U17519 (N_17519,N_15734,N_15683);
nor U17520 (N_17520,N_16685,N_17039);
nor U17521 (N_17521,N_16682,N_16835);
xnor U17522 (N_17522,N_17128,N_16841);
nor U17523 (N_17523,N_16379,N_15666);
xnor U17524 (N_17524,N_17445,N_16784);
nor U17525 (N_17525,N_15964,N_15222);
nor U17526 (N_17526,N_16465,N_15858);
nand U17527 (N_17527,N_16799,N_16075);
nand U17528 (N_17528,N_16808,N_17469);
and U17529 (N_17529,N_15188,N_15331);
and U17530 (N_17530,N_15301,N_15780);
or U17531 (N_17531,N_16629,N_16758);
or U17532 (N_17532,N_16168,N_16130);
and U17533 (N_17533,N_17244,N_15759);
nand U17534 (N_17534,N_16309,N_16282);
nor U17535 (N_17535,N_17216,N_16577);
nand U17536 (N_17536,N_17376,N_17169);
nor U17537 (N_17537,N_16442,N_17024);
nand U17538 (N_17538,N_15934,N_17232);
xnor U17539 (N_17539,N_15347,N_17446);
nor U17540 (N_17540,N_17300,N_15288);
and U17541 (N_17541,N_17463,N_16129);
nor U17542 (N_17542,N_16355,N_16400);
nand U17543 (N_17543,N_16232,N_17093);
xnor U17544 (N_17544,N_15690,N_15004);
nand U17545 (N_17545,N_17360,N_17147);
xnor U17546 (N_17546,N_16572,N_15483);
nor U17547 (N_17547,N_15901,N_16312);
and U17548 (N_17548,N_16584,N_16836);
nand U17549 (N_17549,N_16972,N_17281);
and U17550 (N_17550,N_17037,N_15570);
xnor U17551 (N_17551,N_15430,N_17006);
nand U17552 (N_17552,N_16693,N_17411);
nor U17553 (N_17553,N_16704,N_16343);
nand U17554 (N_17554,N_15883,N_15259);
xor U17555 (N_17555,N_17292,N_17423);
nand U17556 (N_17556,N_16965,N_15557);
nor U17557 (N_17557,N_16051,N_17210);
nand U17558 (N_17558,N_15087,N_16000);
xor U17559 (N_17559,N_16422,N_15456);
nor U17560 (N_17560,N_15420,N_15232);
and U17561 (N_17561,N_15899,N_17062);
or U17562 (N_17562,N_16599,N_15152);
nor U17563 (N_17563,N_16405,N_16617);
nor U17564 (N_17564,N_16973,N_17303);
nand U17565 (N_17565,N_15991,N_17441);
xor U17566 (N_17566,N_16804,N_15798);
and U17567 (N_17567,N_17286,N_15428);
nor U17568 (N_17568,N_17461,N_16790);
or U17569 (N_17569,N_17263,N_15103);
and U17570 (N_17570,N_16194,N_17342);
or U17571 (N_17571,N_15205,N_17105);
nor U17572 (N_17572,N_15956,N_16080);
nand U17573 (N_17573,N_15241,N_15064);
nand U17574 (N_17574,N_15202,N_17011);
xnor U17575 (N_17575,N_15578,N_16543);
or U17576 (N_17576,N_16618,N_15732);
or U17577 (N_17577,N_16328,N_15487);
nand U17578 (N_17578,N_16372,N_16241);
nand U17579 (N_17579,N_15406,N_16297);
nor U17580 (N_17580,N_15309,N_15647);
nor U17581 (N_17581,N_16208,N_15182);
nand U17582 (N_17582,N_17266,N_17204);
or U17583 (N_17583,N_15165,N_15784);
nand U17584 (N_17584,N_17273,N_15958);
xor U17585 (N_17585,N_15393,N_16712);
and U17586 (N_17586,N_16528,N_16513);
or U17587 (N_17587,N_15818,N_15266);
xor U17588 (N_17588,N_16361,N_16498);
nand U17589 (N_17589,N_15919,N_15204);
and U17590 (N_17590,N_15707,N_15906);
nand U17591 (N_17591,N_17237,N_16408);
or U17592 (N_17592,N_16320,N_16741);
xor U17593 (N_17593,N_17056,N_15514);
and U17594 (N_17594,N_15536,N_15215);
nand U17595 (N_17595,N_16619,N_17077);
or U17596 (N_17596,N_16413,N_16564);
xnor U17597 (N_17597,N_16674,N_17151);
or U17598 (N_17598,N_17476,N_16763);
xor U17599 (N_17599,N_16461,N_16411);
or U17600 (N_17600,N_17185,N_15832);
xnor U17601 (N_17601,N_16363,N_17127);
or U17602 (N_17602,N_17311,N_16247);
xor U17603 (N_17603,N_16727,N_17268);
xor U17604 (N_17604,N_17061,N_15334);
nand U17605 (N_17605,N_17161,N_16217);
nor U17606 (N_17606,N_15493,N_15148);
nand U17607 (N_17607,N_16444,N_15414);
nor U17608 (N_17608,N_15836,N_17434);
nand U17609 (N_17609,N_15859,N_15564);
xor U17610 (N_17610,N_16938,N_15867);
xor U17611 (N_17611,N_16658,N_16313);
or U17612 (N_17612,N_15950,N_17012);
nand U17613 (N_17613,N_15752,N_15700);
nand U17614 (N_17614,N_16095,N_15123);
or U17615 (N_17615,N_16531,N_16567);
or U17616 (N_17616,N_16863,N_15348);
or U17617 (N_17617,N_17467,N_16470);
nor U17618 (N_17618,N_15314,N_15865);
nand U17619 (N_17619,N_15474,N_16048);
or U17620 (N_17620,N_16544,N_16036);
and U17621 (N_17621,N_17015,N_16904);
nand U17622 (N_17622,N_15960,N_16056);
or U17623 (N_17623,N_17138,N_16817);
xor U17624 (N_17624,N_15247,N_16061);
or U17625 (N_17625,N_15629,N_15109);
or U17626 (N_17626,N_16010,N_15203);
or U17627 (N_17627,N_16471,N_15404);
nor U17628 (N_17628,N_15371,N_16779);
nand U17629 (N_17629,N_16673,N_15643);
nand U17630 (N_17630,N_16201,N_17223);
nand U17631 (N_17631,N_15691,N_16446);
nand U17632 (N_17632,N_16337,N_16725);
and U17633 (N_17633,N_15135,N_16123);
xnor U17634 (N_17634,N_17453,N_15881);
nand U17635 (N_17635,N_15485,N_16918);
or U17636 (N_17636,N_16474,N_17486);
nand U17637 (N_17637,N_16516,N_17364);
nand U17638 (N_17638,N_15405,N_16407);
xnor U17639 (N_17639,N_16719,N_16738);
nor U17640 (N_17640,N_15876,N_15142);
and U17641 (N_17641,N_16750,N_17014);
nand U17642 (N_17642,N_17245,N_15472);
nor U17643 (N_17643,N_16033,N_15282);
or U17644 (N_17644,N_15534,N_16081);
or U17645 (N_17645,N_15201,N_15885);
xor U17646 (N_17646,N_16218,N_15720);
and U17647 (N_17647,N_16460,N_16625);
nand U17648 (N_17648,N_16563,N_17178);
xor U17649 (N_17649,N_16885,N_16557);
or U17650 (N_17650,N_17170,N_15340);
nor U17651 (N_17651,N_16574,N_16267);
nand U17652 (N_17652,N_15378,N_16714);
and U17653 (N_17653,N_15300,N_15754);
nor U17654 (N_17654,N_16200,N_15333);
nor U17655 (N_17655,N_15829,N_15104);
nand U17656 (N_17656,N_15339,N_15312);
or U17657 (N_17657,N_15594,N_15655);
nand U17658 (N_17658,N_16014,N_16979);
nand U17659 (N_17659,N_16266,N_17343);
xnor U17660 (N_17660,N_17470,N_16233);
nor U17661 (N_17661,N_15048,N_16649);
nor U17662 (N_17662,N_16550,N_16889);
xnor U17663 (N_17663,N_15413,N_15494);
nand U17664 (N_17664,N_17158,N_15637);
xor U17665 (N_17665,N_15617,N_16441);
xnor U17666 (N_17666,N_16590,N_16924);
or U17667 (N_17667,N_17073,N_15726);
and U17668 (N_17668,N_16490,N_16862);
xor U17669 (N_17669,N_15242,N_17316);
nor U17670 (N_17670,N_16187,N_16410);
nand U17671 (N_17671,N_16667,N_16302);
xnor U17672 (N_17672,N_16868,N_16803);
and U17673 (N_17673,N_16899,N_15531);
and U17674 (N_17674,N_17451,N_15091);
nand U17675 (N_17675,N_16393,N_17396);
nor U17676 (N_17676,N_15681,N_15149);
or U17677 (N_17677,N_17233,N_17134);
nand U17678 (N_17678,N_16115,N_15625);
nand U17679 (N_17679,N_16724,N_15774);
and U17680 (N_17680,N_17112,N_15575);
xnor U17681 (N_17681,N_15517,N_17497);
xnor U17682 (N_17682,N_16068,N_16364);
xnor U17683 (N_17683,N_15025,N_15238);
nor U17684 (N_17684,N_16083,N_16270);
xor U17685 (N_17685,N_15808,N_16542);
or U17686 (N_17686,N_17317,N_15668);
nand U17687 (N_17687,N_16031,N_17277);
nand U17688 (N_17688,N_15698,N_16155);
nand U17689 (N_17689,N_16767,N_15030);
nor U17690 (N_17690,N_16416,N_15999);
nor U17691 (N_17691,N_17013,N_16958);
and U17692 (N_17692,N_15069,N_16594);
xnor U17693 (N_17693,N_16978,N_15284);
or U17694 (N_17694,N_17438,N_17101);
xor U17695 (N_17695,N_16634,N_15506);
and U17696 (N_17696,N_16406,N_16537);
or U17697 (N_17697,N_16770,N_15535);
or U17698 (N_17698,N_17338,N_17094);
xor U17699 (N_17699,N_17033,N_16913);
and U17700 (N_17700,N_17257,N_17184);
nor U17701 (N_17701,N_16828,N_15450);
nand U17702 (N_17702,N_16394,N_17293);
and U17703 (N_17703,N_16026,N_16527);
nand U17704 (N_17704,N_17003,N_17179);
nor U17705 (N_17705,N_16339,N_17265);
nand U17706 (N_17706,N_15080,N_15872);
and U17707 (N_17707,N_15552,N_15195);
nor U17708 (N_17708,N_16316,N_17361);
nand U17709 (N_17709,N_17095,N_16521);
xnor U17710 (N_17710,N_15296,N_16191);
nand U17711 (N_17711,N_15143,N_16151);
or U17712 (N_17712,N_15515,N_15137);
nand U17713 (N_17713,N_16887,N_17374);
nor U17714 (N_17714,N_15001,N_17074);
nand U17715 (N_17715,N_15595,N_16532);
nor U17716 (N_17716,N_16482,N_15054);
nand U17717 (N_17717,N_17096,N_15212);
nor U17718 (N_17718,N_15443,N_17189);
and U17719 (N_17719,N_15528,N_15914);
nor U17720 (N_17720,N_16073,N_15351);
nand U17721 (N_17721,N_16699,N_16861);
or U17722 (N_17722,N_15937,N_15267);
or U17723 (N_17723,N_17063,N_16472);
nand U17724 (N_17724,N_16352,N_15678);
nand U17725 (N_17725,N_15381,N_15504);
nand U17726 (N_17726,N_15455,N_16568);
nor U17727 (N_17727,N_16088,N_17358);
and U17728 (N_17728,N_16058,N_15036);
nor U17729 (N_17729,N_15830,N_17218);
nor U17730 (N_17730,N_16167,N_15174);
nand U17731 (N_17731,N_15566,N_15002);
xnor U17732 (N_17732,N_15370,N_17004);
or U17733 (N_17733,N_16966,N_15421);
xnor U17734 (N_17734,N_15875,N_15618);
or U17735 (N_17735,N_16469,N_15724);
nand U17736 (N_17736,N_17082,N_17455);
xnor U17737 (N_17737,N_17367,N_15245);
nand U17738 (N_17738,N_16850,N_15947);
xor U17739 (N_17739,N_16110,N_17492);
nor U17740 (N_17740,N_17304,N_16310);
or U17741 (N_17741,N_17282,N_17239);
nor U17742 (N_17742,N_15927,N_17443);
xnor U17743 (N_17743,N_15304,N_16137);
nor U17744 (N_17744,N_16221,N_15907);
nand U17745 (N_17745,N_16744,N_16571);
or U17746 (N_17746,N_15866,N_16066);
nand U17747 (N_17747,N_16702,N_15993);
and U17748 (N_17748,N_16409,N_15039);
nand U17749 (N_17749,N_16373,N_15753);
nand U17750 (N_17750,N_16246,N_16852);
or U17751 (N_17751,N_15074,N_16652);
xor U17752 (N_17752,N_15649,N_15772);
nand U17753 (N_17753,N_17435,N_15962);
nor U17754 (N_17754,N_15837,N_16365);
xnor U17755 (N_17755,N_16140,N_17318);
and U17756 (N_17756,N_16994,N_15596);
nor U17757 (N_17757,N_16317,N_16632);
and U17758 (N_17758,N_15028,N_16288);
nand U17759 (N_17759,N_17323,N_17329);
or U17760 (N_17760,N_16038,N_16788);
xor U17761 (N_17761,N_17224,N_15363);
and U17762 (N_17762,N_15874,N_15000);
and U17763 (N_17763,N_15930,N_17088);
xnor U17764 (N_17764,N_16358,N_16975);
or U17765 (N_17765,N_16906,N_15856);
xnor U17766 (N_17766,N_15599,N_15912);
nand U17767 (N_17767,N_17291,N_15654);
xor U17768 (N_17768,N_15898,N_17118);
and U17769 (N_17769,N_17089,N_15728);
and U17770 (N_17770,N_15664,N_17044);
nor U17771 (N_17771,N_15822,N_15415);
nand U17772 (N_17772,N_15955,N_15845);
nor U17773 (N_17773,N_15692,N_15446);
or U17774 (N_17774,N_16262,N_16367);
nor U17775 (N_17775,N_17366,N_16616);
or U17776 (N_17776,N_16236,N_17188);
xnor U17777 (N_17777,N_16002,N_15640);
and U17778 (N_17778,N_16807,N_15977);
xor U17779 (N_17779,N_15886,N_16043);
xnor U17780 (N_17780,N_15737,N_16959);
and U17781 (N_17781,N_16555,N_17187);
or U17782 (N_17782,N_16020,N_17227);
and U17783 (N_17783,N_16473,N_16136);
and U17784 (N_17784,N_15055,N_15926);
and U17785 (N_17785,N_15592,N_17120);
and U17786 (N_17786,N_16145,N_15522);
xor U17787 (N_17787,N_16186,N_15855);
or U17788 (N_17788,N_16024,N_15718);
xnor U17789 (N_17789,N_15878,N_16596);
nor U17790 (N_17790,N_17252,N_17036);
or U17791 (N_17791,N_16074,N_15258);
xnor U17792 (N_17792,N_17234,N_15584);
xnor U17793 (N_17793,N_16941,N_16103);
xnor U17794 (N_17794,N_16091,N_15577);
and U17795 (N_17795,N_17045,N_17307);
nor U17796 (N_17796,N_15639,N_16812);
nand U17797 (N_17797,N_15569,N_16660);
nand U17798 (N_17798,N_15892,N_15703);
xnor U17799 (N_17799,N_15398,N_16425);
xnor U17800 (N_17800,N_15359,N_16280);
nand U17801 (N_17801,N_15470,N_15722);
or U17802 (N_17802,N_15375,N_16293);
nand U17803 (N_17803,N_15604,N_15269);
nor U17804 (N_17804,N_16937,N_15748);
and U17805 (N_17805,N_16172,N_16718);
nand U17806 (N_17806,N_15255,N_16120);
or U17807 (N_17807,N_16534,N_15889);
nor U17808 (N_17808,N_17428,N_15003);
or U17809 (N_17809,N_15920,N_15423);
or U17810 (N_17810,N_15904,N_16838);
nor U17811 (N_17811,N_16131,N_17340);
or U17812 (N_17812,N_16902,N_16475);
nor U17813 (N_17813,N_15453,N_15527);
nand U17814 (N_17814,N_15083,N_16418);
and U17815 (N_17815,N_16250,N_15477);
nand U17816 (N_17816,N_15257,N_15646);
nor U17817 (N_17817,N_16391,N_16341);
and U17818 (N_17818,N_16251,N_17473);
and U17819 (N_17819,N_16240,N_16820);
nor U17820 (N_17820,N_15662,N_16797);
nor U17821 (N_17821,N_15841,N_15262);
nand U17822 (N_17822,N_15075,N_16585);
nand U17823 (N_17823,N_15988,N_15384);
or U17824 (N_17824,N_17334,N_15923);
nor U17825 (N_17825,N_16794,N_16968);
and U17826 (N_17826,N_16381,N_15176);
nor U17827 (N_17827,N_15864,N_17295);
nor U17828 (N_17828,N_15153,N_16831);
or U17829 (N_17829,N_15161,N_16069);
xnor U17830 (N_17830,N_16519,N_17313);
nand U17831 (N_17831,N_16064,N_17000);
nor U17832 (N_17832,N_15175,N_16922);
and U17833 (N_17833,N_16325,N_16440);
nor U17834 (N_17834,N_17081,N_17274);
nand U17835 (N_17835,N_16775,N_15224);
nand U17836 (N_17836,N_16686,N_15067);
nor U17837 (N_17837,N_15173,N_15727);
xnor U17838 (N_17838,N_15987,N_16283);
and U17839 (N_17839,N_15439,N_16466);
or U17840 (N_17840,N_15248,N_15317);
or U17841 (N_17841,N_15660,N_17259);
nor U17842 (N_17842,N_15518,N_16896);
xnor U17843 (N_17843,N_16327,N_15685);
or U17844 (N_17844,N_16787,N_15234);
nand U17845 (N_17845,N_16322,N_15658);
and U17846 (N_17846,N_17436,N_16171);
or U17847 (N_17847,N_15441,N_16121);
and U17848 (N_17848,N_17191,N_15082);
nor U17849 (N_17849,N_15589,N_16087);
nor U17850 (N_17850,N_16695,N_16829);
or U17851 (N_17851,N_15277,N_17154);
nand U17852 (N_17852,N_15825,N_17162);
and U17853 (N_17853,N_17009,N_16908);
or U17854 (N_17854,N_17007,N_17198);
xor U17855 (N_17855,N_17071,N_16864);
and U17856 (N_17856,N_16759,N_15032);
and U17857 (N_17857,N_17035,N_15221);
and U17858 (N_17858,N_16261,N_16108);
and U17859 (N_17859,N_16910,N_15574);
and U17860 (N_17860,N_15719,N_17489);
or U17861 (N_17861,N_17382,N_15873);
or U17862 (N_17862,N_16291,N_15146);
or U17863 (N_17863,N_15613,N_15337);
or U17864 (N_17864,N_16396,N_16911);
xnor U17865 (N_17865,N_15403,N_17222);
xor U17866 (N_17866,N_17401,N_17080);
xor U17867 (N_17867,N_15389,N_17116);
and U17868 (N_17868,N_15480,N_15417);
or U17869 (N_17869,N_16326,N_16220);
nand U17870 (N_17870,N_16376,N_16936);
or U17871 (N_17871,N_16886,N_16215);
nor U17872 (N_17872,N_16678,N_16598);
xnor U17873 (N_17873,N_16454,N_17275);
nor U17874 (N_17874,N_15969,N_16017);
nor U17875 (N_17875,N_16622,N_15560);
and U17876 (N_17876,N_15893,N_16492);
or U17877 (N_17877,N_15014,N_15133);
and U17878 (N_17878,N_15396,N_16749);
or U17879 (N_17879,N_15448,N_16610);
nor U17880 (N_17880,N_15931,N_16995);
nand U17881 (N_17881,N_15971,N_17168);
and U17882 (N_17882,N_16299,N_17022);
nor U17883 (N_17883,N_16672,N_15547);
and U17884 (N_17884,N_17214,N_17440);
or U17885 (N_17885,N_16971,N_15435);
or U17886 (N_17886,N_15635,N_15656);
nor U17887 (N_17887,N_17398,N_16076);
and U17888 (N_17888,N_16970,N_15313);
xnor U17889 (N_17889,N_16743,N_15023);
nand U17890 (N_17890,N_16640,N_17498);
nor U17891 (N_17891,N_15896,N_16207);
and U17892 (N_17892,N_16984,N_17250);
or U17893 (N_17893,N_16637,N_15796);
nand U17894 (N_17894,N_16209,N_16184);
and U17895 (N_17895,N_17215,N_17171);
nand U17896 (N_17896,N_15997,N_15925);
nand U17897 (N_17897,N_17328,N_15177);
or U17898 (N_17898,N_15965,N_15125);
xor U17899 (N_17899,N_17392,N_15641);
nor U17900 (N_17900,N_17391,N_15422);
nand U17901 (N_17901,N_16047,N_15121);
nor U17902 (N_17902,N_17219,N_16524);
nor U17903 (N_17903,N_15828,N_16847);
nor U17904 (N_17904,N_16401,N_15373);
and U17905 (N_17905,N_16188,N_15605);
and U17906 (N_17906,N_15332,N_15492);
xnor U17907 (N_17907,N_16070,N_15061);
nor U17908 (N_17908,N_17241,N_15326);
xnor U17909 (N_17909,N_15017,N_15290);
and U17910 (N_17910,N_17430,N_17065);
and U17911 (N_17911,N_17249,N_16855);
nand U17912 (N_17912,N_15489,N_16062);
nor U17913 (N_17913,N_17331,N_16204);
and U17914 (N_17914,N_16424,N_16426);
nand U17915 (N_17915,N_15085,N_17019);
xnor U17916 (N_17916,N_15622,N_17246);
xor U17917 (N_17917,N_15524,N_17194);
xor U17918 (N_17918,N_15717,N_15814);
nor U17919 (N_17919,N_17356,N_16340);
nand U17920 (N_17920,N_16044,N_15844);
nand U17921 (N_17921,N_16366,N_15807);
xor U17922 (N_17922,N_16905,N_15994);
or U17923 (N_17923,N_15941,N_15766);
or U17924 (N_17924,N_15488,N_17055);
and U17925 (N_17925,N_17308,N_16771);
nor U17926 (N_17926,N_15037,N_16300);
xor U17927 (N_17927,N_16153,N_16977);
nor U17928 (N_17928,N_15338,N_16591);
xnor U17929 (N_17929,N_16830,N_16554);
xor U17930 (N_17930,N_16211,N_15432);
xor U17931 (N_17931,N_15760,N_15795);
nand U17932 (N_17932,N_16792,N_16739);
nand U17933 (N_17933,N_15022,N_16547);
and U17934 (N_17934,N_16037,N_17341);
and U17935 (N_17935,N_15358,N_15129);
xor U17936 (N_17936,N_17196,N_17190);
nor U17937 (N_17937,N_16898,N_16751);
nor U17938 (N_17938,N_16601,N_15507);
and U17939 (N_17939,N_16754,N_15132);
nand U17940 (N_17940,N_15088,N_15741);
xor U17941 (N_17941,N_15653,N_16375);
xnor U17942 (N_17942,N_16633,N_15297);
xnor U17943 (N_17943,N_16294,N_15005);
or U17944 (N_17944,N_15226,N_16258);
nor U17945 (N_17945,N_15180,N_15018);
or U17946 (N_17946,N_15471,N_15362);
nand U17947 (N_17947,N_16114,N_16330);
nor U17948 (N_17948,N_17348,N_16730);
nand U17949 (N_17949,N_15696,N_17163);
nand U17950 (N_17950,N_16356,N_15330);
or U17951 (N_17951,N_16022,N_15982);
xnor U17952 (N_17952,N_15544,N_16737);
nor U17953 (N_17953,N_17412,N_16272);
and U17954 (N_17954,N_17459,N_16234);
and U17955 (N_17955,N_16152,N_16996);
and U17956 (N_17956,N_16007,N_15100);
or U17957 (N_17957,N_17264,N_17439);
nor U17958 (N_17958,N_15973,N_16881);
or U17959 (N_17959,N_17468,N_15163);
or U17960 (N_17960,N_16404,N_16459);
nand U17961 (N_17961,N_16450,N_16092);
nor U17962 (N_17962,N_16742,N_16696);
xor U17963 (N_17963,N_15164,N_16222);
nand U17964 (N_17964,N_15512,N_17475);
or U17965 (N_17965,N_16548,N_17251);
nand U17966 (N_17966,N_15626,N_16858);
nand U17967 (N_17967,N_15848,N_15790);
xor U17968 (N_17968,N_17261,N_16089);
nor U17969 (N_17969,N_17491,N_15612);
nand U17970 (N_17970,N_17287,N_16694);
nor U17971 (N_17971,N_16657,N_16785);
nand U17972 (N_17972,N_16882,N_15058);
or U17973 (N_17973,N_16957,N_17109);
nand U17974 (N_17974,N_15213,N_15736);
and U17975 (N_17975,N_15981,N_16414);
nor U17976 (N_17976,N_16735,N_16039);
xnor U17977 (N_17977,N_15293,N_15156);
nor U17978 (N_17978,N_16117,N_15105);
and U17979 (N_17979,N_16745,N_17351);
nand U17980 (N_17980,N_15963,N_15523);
and U17981 (N_17981,N_16688,N_17289);
or U17982 (N_17982,N_16052,N_15851);
and U17983 (N_17983,N_15767,N_17148);
or U17984 (N_17984,N_16538,N_15498);
or U17985 (N_17985,N_15775,N_15995);
xnor U17986 (N_17986,N_15281,N_15272);
xnor U17987 (N_17987,N_16254,N_15520);
xnor U17988 (N_17988,N_17408,N_16273);
nand U17989 (N_17989,N_17280,N_16848);
nor U17990 (N_17990,N_15568,N_15806);
or U17991 (N_17991,N_16940,N_15335);
nand U17992 (N_17992,N_17452,N_15631);
nor U17993 (N_17993,N_15240,N_16578);
xor U17994 (N_17994,N_17296,N_15648);
or U17995 (N_17995,N_17302,N_16684);
nor U17996 (N_17996,N_16212,N_16664);
and U17997 (N_17997,N_15782,N_15833);
or U17998 (N_17998,N_15343,N_17336);
and U17999 (N_17999,N_15169,N_15299);
and U18000 (N_18000,N_15412,N_16183);
or U18001 (N_18001,N_15739,N_17290);
and U18002 (N_18002,N_17235,N_15645);
xnor U18003 (N_18003,N_15509,N_17032);
nand U18004 (N_18004,N_16205,N_15989);
xnor U18005 (N_18005,N_16810,N_15440);
and U18006 (N_18006,N_16565,N_16728);
and U18007 (N_18007,N_16740,N_15597);
xnor U18008 (N_18008,N_16986,N_17381);
or U18009 (N_18009,N_17378,N_15644);
nor U18010 (N_18010,N_17064,N_16976);
and U18011 (N_18011,N_16001,N_15862);
xor U18012 (N_18012,N_15765,N_16468);
or U18013 (N_18013,N_16439,N_17260);
or U18014 (N_18014,N_15467,N_15650);
or U18015 (N_18015,N_15743,N_17217);
nor U18016 (N_18016,N_17375,N_16569);
nor U18017 (N_18017,N_17104,N_17448);
or U18018 (N_18018,N_17107,N_17069);
xor U18019 (N_18019,N_16100,N_15713);
nand U18020 (N_18020,N_16801,N_16903);
xnor U18021 (N_18021,N_17403,N_15217);
and U18022 (N_18022,N_15549,N_16398);
nor U18023 (N_18023,N_15824,N_17200);
or U18024 (N_18024,N_16333,N_17373);
or U18025 (N_18025,N_17369,N_17058);
or U18026 (N_18026,N_16150,N_16562);
and U18027 (N_18027,N_15095,N_15449);
nor U18028 (N_18028,N_17460,N_16748);
nor U18029 (N_18029,N_15364,N_15126);
xor U18030 (N_18030,N_17420,N_16195);
and U18031 (N_18031,N_17208,N_16897);
and U18032 (N_18032,N_16230,N_16845);
and U18033 (N_18033,N_16974,N_16556);
xor U18034 (N_18034,N_15801,N_16782);
or U18035 (N_18035,N_17267,N_17103);
nand U18036 (N_18036,N_17149,N_16213);
and U18037 (N_18037,N_15157,N_17315);
xor U18038 (N_18038,N_15196,N_16259);
nand U18039 (N_18039,N_17068,N_17368);
nand U18040 (N_18040,N_15260,N_16950);
and U18041 (N_18041,N_15840,N_16216);
nor U18042 (N_18042,N_15992,N_15852);
and U18043 (N_18043,N_15352,N_16869);
nor U18044 (N_18044,N_15699,N_15096);
nand U18045 (N_18045,N_15688,N_15099);
xor U18046 (N_18046,N_16900,N_17027);
nand U18047 (N_18047,N_16588,N_17099);
and U18048 (N_18048,N_15278,N_15261);
nor U18049 (N_18049,N_15571,N_15586);
nor U18050 (N_18050,N_16552,N_15218);
nand U18051 (N_18051,N_16654,N_15410);
or U18052 (N_18052,N_17270,N_16265);
xnor U18053 (N_18053,N_17180,N_16529);
and U18054 (N_18054,N_15167,N_15070);
nand U18055 (N_18055,N_15322,N_16774);
and U18056 (N_18056,N_15860,N_16156);
nand U18057 (N_18057,N_15868,N_16060);
or U18058 (N_18058,N_15327,N_15539);
nor U18059 (N_18059,N_16301,N_16304);
and U18060 (N_18060,N_16387,N_15056);
xor U18061 (N_18061,N_16520,N_16920);
xor U18062 (N_18062,N_15463,N_15820);
or U18063 (N_18063,N_16860,N_16226);
or U18064 (N_18064,N_16483,N_15682);
nor U18065 (N_18065,N_16447,N_16597);
and U18066 (N_18066,N_15540,N_16493);
and U18067 (N_18067,N_16278,N_16138);
or U18068 (N_18068,N_16582,N_16306);
nand U18069 (N_18069,N_16045,N_15053);
xnor U18070 (N_18070,N_16099,N_16223);
and U18071 (N_18071,N_16698,N_16357);
nor U18072 (N_18072,N_17462,N_16178);
nor U18073 (N_18073,N_16536,N_15078);
or U18074 (N_18074,N_15183,N_16244);
and U18075 (N_18075,N_17110,N_15651);
or U18076 (N_18076,N_17236,N_16675);
and U18077 (N_18077,N_17247,N_17383);
nor U18078 (N_18078,N_16545,N_15590);
or U18079 (N_18079,N_16636,N_15679);
nand U18080 (N_18080,N_16822,N_16919);
nand U18081 (N_18081,N_16023,N_16821);
nand U18082 (N_18082,N_15433,N_15452);
nand U18083 (N_18083,N_16501,N_16951);
nand U18084 (N_18084,N_15538,N_16050);
nor U18085 (N_18085,N_16587,N_16101);
nor U18086 (N_18086,N_16586,N_15086);
nor U18087 (N_18087,N_17076,N_16846);
xnor U18088 (N_18088,N_17098,N_15178);
xnor U18089 (N_18089,N_17226,N_15044);
xor U18090 (N_18090,N_17075,N_16457);
or U18091 (N_18091,N_17314,N_17156);
or U18092 (N_18092,N_16746,N_15211);
nand U18093 (N_18093,N_16006,N_16494);
xor U18094 (N_18094,N_17283,N_17206);
and U18095 (N_18095,N_15073,N_17294);
xnor U18096 (N_18096,N_17397,N_16260);
xnor U18097 (N_18097,N_15744,N_17301);
nand U18098 (N_18098,N_15891,N_15111);
and U18099 (N_18099,N_15551,N_16224);
nand U18100 (N_18100,N_16627,N_15819);
and U18101 (N_18101,N_15380,N_15979);
xnor U18102 (N_18102,N_15140,N_15438);
or U18103 (N_18103,N_15031,N_15854);
nor U18104 (N_18104,N_16934,N_16096);
xor U18105 (N_18105,N_17352,N_16535);
and U18106 (N_18106,N_16456,N_15320);
nand U18107 (N_18107,N_16126,N_16561);
nor U18108 (N_18108,N_15811,N_17197);
or U18109 (N_18109,N_16268,N_16202);
or U18110 (N_18110,N_16013,N_15120);
and U18111 (N_18111,N_15235,N_16849);
or U18112 (N_18112,N_16755,N_17157);
xor U18113 (N_18113,N_16691,N_16546);
xnor U18114 (N_18114,N_16390,N_15329);
xor U18115 (N_18115,N_15230,N_15857);
nor U18116 (N_18116,N_17049,N_16018);
xnor U18117 (N_18117,N_15444,N_16815);
and U18118 (N_18118,N_15179,N_17025);
nor U18119 (N_18119,N_16912,N_17407);
nand U18120 (N_18120,N_17425,N_15013);
nor U18121 (N_18121,N_15611,N_17057);
nand U18122 (N_18122,N_16963,N_16179);
and U18123 (N_18123,N_16690,N_16960);
or U18124 (N_18124,N_15735,N_16107);
nor U18125 (N_18125,N_15015,N_16789);
nor U18126 (N_18126,N_15581,N_15199);
xor U18127 (N_18127,N_15786,N_15006);
nor U18128 (N_18128,N_15704,N_15318);
or U18129 (N_18129,N_16383,N_15117);
and U18130 (N_18130,N_16478,N_15697);
or U18131 (N_18131,N_16500,N_15545);
nor U18132 (N_18132,N_16488,N_15853);
nor U18133 (N_18133,N_16443,N_17386);
nor U18134 (N_18134,N_16182,N_15062);
nand U18135 (N_18135,N_17487,N_16392);
or U18136 (N_18136,N_15081,N_16507);
or U18137 (N_18137,N_16436,N_17332);
and U18138 (N_18138,N_15516,N_16421);
nor U18139 (N_18139,N_15621,N_15311);
nor U18140 (N_18140,N_16321,N_16229);
xnor U18141 (N_18141,N_16796,N_16480);
nor U18142 (N_18142,N_17370,N_16621);
xnor U18143 (N_18143,N_15310,N_15116);
nand U18144 (N_18144,N_15057,N_16783);
nand U18145 (N_18145,N_16197,N_16289);
nand U18146 (N_18146,N_15940,N_16723);
nand U18147 (N_18147,N_17354,N_16263);
nand U18148 (N_18148,N_16999,N_17464);
xnor U18149 (N_18149,N_16781,N_16559);
or U18150 (N_18150,N_16916,N_16517);
and U18151 (N_18151,N_15084,N_15465);
xor U18152 (N_18152,N_16635,N_16124);
or U18153 (N_18153,N_16997,N_15409);
nor U18154 (N_18154,N_15253,N_15065);
and U18155 (N_18155,N_16496,N_15319);
and U18156 (N_18156,N_16515,N_16235);
nor U18157 (N_18157,N_15461,N_15150);
xor U18158 (N_18158,N_15887,N_15835);
or U18159 (N_18159,N_17330,N_16747);
nor U18160 (N_18160,N_17066,N_15591);
and U18161 (N_18161,N_15770,N_15888);
and U18162 (N_18162,N_17031,N_15063);
nor U18163 (N_18163,N_17499,N_15124);
nand U18164 (N_18164,N_17070,N_16765);
nor U18165 (N_18165,N_15010,N_15812);
nand U18166 (N_18166,N_16206,N_15115);
nor U18167 (N_18167,N_15502,N_16174);
and U18168 (N_18168,N_15251,N_15108);
nor U18169 (N_18169,N_16015,N_16112);
or U18170 (N_18170,N_16707,N_16651);
nand U18171 (N_18171,N_15946,N_16351);
and U18172 (N_18172,N_16700,N_15986);
xor U18173 (N_18173,N_16666,N_16295);
xnor U18174 (N_18174,N_15271,N_16917);
nand U18175 (N_18175,N_15667,N_17297);
nor U18176 (N_18176,N_17333,N_16476);
or U18177 (N_18177,N_15607,N_17404);
nor U18178 (N_18178,N_17142,N_15090);
nand U18179 (N_18179,N_16093,N_17141);
xnor U18180 (N_18180,N_16484,N_16716);
nor U18181 (N_18181,N_15968,N_16539);
xnor U18182 (N_18182,N_16380,N_16290);
nor U18183 (N_18183,N_16005,N_15712);
nor U18184 (N_18184,N_17078,N_15499);
nand U18185 (N_18185,N_16296,N_17001);
and U18186 (N_18186,N_17402,N_16181);
nor U18187 (N_18187,N_15936,N_15503);
nand U18188 (N_18188,N_15670,N_16834);
xor U18189 (N_18189,N_15387,N_16382);
and U18190 (N_18190,N_15763,N_16883);
nor U18191 (N_18191,N_17152,N_17419);
xor U18192 (N_18192,N_16687,N_15777);
and U18193 (N_18193,N_15399,N_15229);
nand U18194 (N_18194,N_15029,N_17153);
nor U18195 (N_18195,N_16102,N_16944);
and U18196 (N_18196,N_15089,N_16602);
xor U18197 (N_18197,N_16346,N_17091);
and U18198 (N_18198,N_15530,N_16566);
or U18199 (N_18199,N_16776,N_15424);
and U18200 (N_18200,N_17450,N_16228);
nand U18201 (N_18201,N_16189,N_15019);
nand U18202 (N_18202,N_15587,N_16573);
or U18203 (N_18203,N_15171,N_16029);
or U18204 (N_18204,N_17380,N_17482);
or U18205 (N_18205,N_16487,N_15007);
xor U18206 (N_18206,N_17060,N_15911);
nand U18207 (N_18207,N_17195,N_16990);
or U18208 (N_18208,N_15961,N_15792);
nor U18209 (N_18209,N_17113,N_17084);
or U18210 (N_18210,N_15496,N_16777);
nor U18211 (N_18211,N_17123,N_17051);
and U18212 (N_18212,N_16034,N_16530);
or U18213 (N_18213,N_17344,N_15944);
xnor U18214 (N_18214,N_16106,N_16332);
and U18215 (N_18215,N_15127,N_15458);
nand U18216 (N_18216,N_17355,N_16987);
or U18217 (N_18217,N_15418,N_16437);
nand U18218 (N_18218,N_16872,N_16626);
xor U18219 (N_18219,N_15804,N_16242);
nand U18220 (N_18220,N_15379,N_17258);
xor U18221 (N_18221,N_17388,N_15368);
xnor U18222 (N_18222,N_15779,N_16276);
nand U18223 (N_18223,N_15863,N_16353);
and U18224 (N_18224,N_16607,N_16429);
xnor U18225 (N_18225,N_17406,N_16415);
xor U18226 (N_18226,N_16592,N_15943);
and U18227 (N_18227,N_15815,N_16928);
xor U18228 (N_18228,N_16495,N_16134);
and U18229 (N_18229,N_15902,N_15092);
nand U18230 (N_18230,N_15360,N_16873);
nand U18231 (N_18231,N_15638,N_15813);
and U18232 (N_18232,N_16505,N_17199);
or U18233 (N_18233,N_16347,N_15600);
or U18234 (N_18234,N_16395,N_15395);
and U18235 (N_18235,N_15939,N_17421);
xnor U18236 (N_18236,N_16842,N_17238);
nor U18237 (N_18237,N_15361,N_17026);
or U18238 (N_18238,N_15285,N_17496);
or U18239 (N_18239,N_16624,N_17335);
xnor U18240 (N_18240,N_15526,N_15394);
or U18241 (N_18241,N_17115,N_16298);
and U18242 (N_18242,N_17203,N_16004);
or U18243 (N_18243,N_15723,N_15476);
nor U18244 (N_18244,N_17494,N_15071);
or U18245 (N_18245,N_16638,N_17248);
or U18246 (N_18246,N_16576,N_16122);
nor U18247 (N_18247,N_17363,N_17490);
xor U18248 (N_18248,N_16097,N_16870);
xor U18249 (N_18249,N_16430,N_16256);
nor U18250 (N_18250,N_16533,N_16720);
nand U18251 (N_18251,N_17484,N_15580);
or U18252 (N_18252,N_16027,N_16336);
or U18253 (N_18253,N_16955,N_15021);
and U18254 (N_18254,N_15189,N_15068);
or U18255 (N_18255,N_17155,N_16643);
nand U18256 (N_18256,N_17087,N_16818);
and U18257 (N_18257,N_16953,N_16198);
and U18258 (N_18258,N_15482,N_15365);
xor U18259 (N_18259,N_16604,N_16549);
and U18260 (N_18260,N_16871,N_16992);
nand U18261 (N_18261,N_16823,N_15838);
nand U18262 (N_18262,N_17160,N_15711);
or U18263 (N_18263,N_17029,N_15565);
xnor U18264 (N_18264,N_17050,N_16455);
nor U18265 (N_18265,N_15628,N_16653);
or U18266 (N_18266,N_16084,N_17415);
or U18267 (N_18267,N_15454,N_15040);
nand U18268 (N_18268,N_16703,N_15733);
xor U18269 (N_18269,N_16662,N_16499);
and U18270 (N_18270,N_15491,N_15976);
or U18271 (N_18271,N_16943,N_16119);
nor U18272 (N_18272,N_17023,N_16163);
nand U18273 (N_18273,N_15823,N_17117);
xnor U18274 (N_18274,N_15579,N_15952);
nand U18275 (N_18275,N_16932,N_16190);
nand U18276 (N_18276,N_17030,N_15525);
nor U18277 (N_18277,N_15097,N_17319);
or U18278 (N_18278,N_17166,N_15077);
or U18279 (N_18279,N_17140,N_16608);
or U18280 (N_18280,N_16063,N_16362);
nor U18281 (N_18281,N_15805,N_15505);
or U18282 (N_18282,N_16142,N_17132);
nand U18283 (N_18283,N_15328,N_16125);
or U18284 (N_18284,N_17020,N_17175);
xnor U18285 (N_18285,N_16285,N_16154);
nor U18286 (N_18286,N_15350,N_16711);
or U18287 (N_18287,N_17253,N_16676);
and U18288 (N_18288,N_15910,N_17040);
or U18289 (N_18289,N_16319,N_15342);
and U18290 (N_18290,N_17346,N_16342);
and U18291 (N_18291,N_17177,N_16766);
and U18292 (N_18292,N_15978,N_17357);
or U18293 (N_18293,N_16504,N_17131);
nor U18294 (N_18294,N_15237,N_16722);
nand U18295 (N_18295,N_17465,N_16508);
and U18296 (N_18296,N_16463,N_16359);
and U18297 (N_18297,N_15900,N_16923);
and U18298 (N_18298,N_16772,N_17086);
and U18299 (N_18299,N_17324,N_16931);
nor U18300 (N_18300,N_15572,N_15147);
or U18301 (N_18301,N_17298,N_16570);
nor U18302 (N_18302,N_16648,N_17306);
and U18303 (N_18303,N_15513,N_15563);
nand U18304 (N_18304,N_16082,N_15555);
nand U18305 (N_18305,N_15110,N_15325);
xnor U18306 (N_18306,N_17256,N_15401);
nor U18307 (N_18307,N_15186,N_17016);
and U18308 (N_18308,N_16314,N_15139);
or U18309 (N_18309,N_16225,N_16041);
nor U18310 (N_18310,N_15608,N_16128);
and U18311 (N_18311,N_16199,N_15008);
nand U18312 (N_18312,N_15842,N_15602);
or U18313 (N_18313,N_16378,N_16967);
nand U18314 (N_18314,N_15787,N_16162);
and U18315 (N_18315,N_17090,N_16884);
and U18316 (N_18316,N_16580,N_15929);
or U18317 (N_18317,N_16945,N_15141);
xnor U18318 (N_18318,N_16933,N_16274);
nand U18319 (N_18319,N_15066,N_17174);
nor U18320 (N_18320,N_16435,N_16445);
or U18321 (N_18321,N_16837,N_15709);
or U18322 (N_18322,N_16428,N_16780);
and U18323 (N_18323,N_15219,N_15680);
or U18324 (N_18324,N_16892,N_15957);
nor U18325 (N_18325,N_17365,N_16891);
nand U18326 (N_18326,N_15742,N_17119);
or U18327 (N_18327,N_16708,N_16930);
and U18328 (N_18328,N_17221,N_16277);
xnor U18329 (N_18329,N_15882,N_16176);
nor U18330 (N_18330,N_16595,N_15603);
and U18331 (N_18331,N_17272,N_15975);
xor U18332 (N_18332,N_15794,N_16497);
nor U18333 (N_18333,N_16839,N_17159);
nor U18334 (N_18334,N_16417,N_17326);
or U18335 (N_18335,N_15402,N_15598);
and U18336 (N_18336,N_16907,N_16706);
or U18337 (N_18337,N_16512,N_16795);
xnor U18338 (N_18338,N_15663,N_16433);
nand U18339 (N_18339,N_15546,N_15307);
and U18340 (N_18340,N_15797,N_16214);
xnor U18341 (N_18341,N_17146,N_16993);
nor U18342 (N_18342,N_16451,N_17047);
nand U18343 (N_18343,N_16721,N_15052);
and U18344 (N_18344,N_16935,N_16284);
or U18345 (N_18345,N_15671,N_16249);
xor U18346 (N_18346,N_17092,N_17254);
nor U18347 (N_18347,N_16028,N_16021);
and U18348 (N_18348,N_16292,N_17347);
nor U18349 (N_18349,N_17433,N_17394);
or U18350 (N_18350,N_16196,N_17137);
or U18351 (N_18351,N_16514,N_16553);
nand U18352 (N_18352,N_16980,N_15562);
nand U18353 (N_18353,N_16303,N_15935);
xor U18354 (N_18354,N_17410,N_16773);
nor U18355 (N_18355,N_16386,N_16630);
xnor U18356 (N_18356,N_15354,N_15138);
nor U18357 (N_18357,N_16692,N_16477);
nor U18358 (N_18358,N_15469,N_16669);
and U18359 (N_18359,N_15416,N_15706);
nor U18360 (N_18360,N_16344,N_15154);
or U18361 (N_18361,N_15249,N_15252);
nor U18362 (N_18362,N_16434,N_15559);
xnor U18363 (N_18363,N_15198,N_16350);
nand U18364 (N_18364,N_16894,N_15916);
or U18365 (N_18365,N_16949,N_17312);
xor U18366 (N_18366,N_16243,N_15431);
xnor U18367 (N_18367,N_16318,N_15291);
xnor U18368 (N_18368,N_17414,N_16644);
nand U18369 (N_18369,N_17456,N_16661);
nand U18370 (N_18370,N_15756,N_15118);
nor U18371 (N_18371,N_15834,N_15305);
nand U18372 (N_18372,N_17181,N_17437);
or U18373 (N_18373,N_15582,N_15392);
and U18374 (N_18374,N_15377,N_15383);
nor U18375 (N_18375,N_16431,N_17002);
and U18376 (N_18376,N_16286,N_15909);
nor U18377 (N_18377,N_15903,N_16030);
nand U18378 (N_18378,N_16059,N_15367);
or U18379 (N_18379,N_16948,N_15627);
xor U18380 (N_18380,N_15793,N_17209);
xnor U18381 (N_18381,N_15928,N_15548);
nand U18382 (N_18382,N_15849,N_15033);
nand U18383 (N_18383,N_16879,N_15273);
nor U18384 (N_18384,N_17485,N_15847);
nand U18385 (N_18385,N_15481,N_16423);
and U18386 (N_18386,N_15466,N_17240);
or U18387 (N_18387,N_17413,N_15274);
nor U18388 (N_18388,N_17483,N_16219);
or U18389 (N_18389,N_17213,N_15382);
nor U18390 (N_18390,N_17097,N_16893);
or U18391 (N_18391,N_16939,N_17173);
xor U18392 (N_18392,N_17349,N_15208);
nor U18393 (N_18393,N_16193,N_15537);
xor U18394 (N_18394,N_16833,N_15781);
nor U18395 (N_18395,N_15731,N_17192);
nand U18396 (N_18396,N_15475,N_15614);
and U18397 (N_18397,N_15192,N_15193);
nor U18398 (N_18398,N_17010,N_16981);
xor U18399 (N_18399,N_16927,N_16732);
xnor U18400 (N_18400,N_16334,N_15918);
nand U18401 (N_18401,N_16628,N_15803);
or U18402 (N_18402,N_15740,N_16384);
or U18403 (N_18403,N_17477,N_15897);
and U18404 (N_18404,N_16526,N_15145);
nand U18405 (N_18405,N_15676,N_17176);
or U18406 (N_18406,N_16111,N_16025);
or U18407 (N_18407,N_17130,N_16854);
or U18408 (N_18408,N_15376,N_17481);
and U18409 (N_18409,N_15355,N_15214);
nand U18410 (N_18410,N_17262,N_15462);
nor U18411 (N_18411,N_15194,N_15486);
nand U18412 (N_18412,N_15672,N_16146);
nand U18413 (N_18413,N_16511,N_16593);
and U18414 (N_18414,N_15757,N_16046);
nand U18415 (N_18415,N_16844,N_16982);
nand U18416 (N_18416,N_16159,N_17320);
nand U18417 (N_18417,N_17493,N_16715);
nand U18418 (N_18418,N_17384,N_15184);
and U18419 (N_18419,N_15162,N_16094);
xor U18420 (N_18420,N_15776,N_16180);
or U18421 (N_18421,N_17136,N_16113);
nor U18422 (N_18422,N_15051,N_17379);
nor U18423 (N_18423,N_16752,N_15665);
or U18424 (N_18424,N_15344,N_16147);
or U18425 (N_18425,N_16679,N_17125);
xor U18426 (N_18426,N_16412,N_15967);
and U18427 (N_18427,N_15447,N_15231);
or U18428 (N_18428,N_15478,N_17424);
and U18429 (N_18429,N_16403,N_17230);
and U18430 (N_18430,N_15924,N_16502);
nand U18431 (N_18431,N_17122,N_15519);
xnor U18432 (N_18432,N_16255,N_15561);
xnor U18433 (N_18433,N_16756,N_16098);
or U18434 (N_18434,N_17133,N_15745);
or U18435 (N_18435,N_15556,N_16257);
xnor U18436 (N_18436,N_17079,N_16040);
nor U18437 (N_18437,N_15725,N_17005);
xor U18438 (N_18438,N_16581,N_15185);
or U18439 (N_18439,N_15270,N_16670);
xor U18440 (N_18440,N_15197,N_15011);
xnor U18441 (N_18441,N_16166,N_16231);
nor U18442 (N_18442,N_16778,N_17458);
nand U18443 (N_18443,N_16614,N_15323);
xor U18444 (N_18444,N_15541,N_17182);
nor U18445 (N_18445,N_15619,N_16518);
xnor U18446 (N_18446,N_15542,N_16677);
and U18447 (N_18447,N_16843,N_15324);
or U18448 (N_18448,N_16177,N_15460);
nor U18449 (N_18449,N_16486,N_15953);
xor U18450 (N_18450,N_15714,N_16683);
or U18451 (N_18451,N_15788,N_16315);
or U18452 (N_18452,N_17172,N_16067);
and U18453 (N_18453,N_17021,N_15216);
nor U18454 (N_18454,N_16736,N_15349);
xor U18455 (N_18455,N_16901,N_16397);
nand U18456 (N_18456,N_16385,N_17018);
and U18457 (N_18457,N_15400,N_17488);
or U18458 (N_18458,N_15298,N_16071);
or U18459 (N_18459,N_16307,N_15407);
nand U18460 (N_18460,N_15620,N_16645);
nand U18461 (N_18461,N_15035,N_15034);
nor U18462 (N_18462,N_16135,N_17043);
or U18463 (N_18463,N_15588,N_15747);
nor U18464 (N_18464,N_15716,N_15050);
and U18465 (N_18465,N_17322,N_16078);
nand U18466 (N_18466,N_15783,N_16985);
nor U18467 (N_18467,N_16275,N_16811);
nor U18468 (N_18468,N_16612,N_15106);
and U18469 (N_18469,N_17255,N_15302);
or U18470 (N_18470,N_15948,N_15128);
nor U18471 (N_18471,N_16641,N_17106);
xor U18472 (N_18472,N_17231,N_16133);
and U18473 (N_18473,N_15996,N_16615);
xnor U18474 (N_18474,N_17416,N_16185);
and U18475 (N_18475,N_15113,N_16825);
and U18476 (N_18476,N_15292,N_17444);
and U18477 (N_18477,N_17472,N_17288);
xor U18478 (N_18478,N_17309,N_15356);
nand U18479 (N_18479,N_15768,N_15501);
nand U18480 (N_18480,N_15321,N_15894);
nor U18481 (N_18481,N_17144,N_15294);
or U18482 (N_18482,N_16793,N_16926);
and U18483 (N_18483,N_16149,N_15749);
or U18484 (N_18484,N_16248,N_17321);
nand U18485 (N_18485,N_17389,N_16169);
and U18486 (N_18486,N_16867,N_17201);
and U18487 (N_18487,N_15593,N_17442);
xor U18488 (N_18488,N_16012,N_16655);
or U18489 (N_18489,N_17202,N_16323);
xnor U18490 (N_18490,N_17028,N_17145);
and U18491 (N_18491,N_17059,N_15985);
nor U18492 (N_18492,N_16009,N_16832);
nor U18493 (N_18493,N_15677,N_16157);
xor U18494 (N_18494,N_16305,N_15913);
or U18495 (N_18495,N_15701,N_16876);
xnor U18496 (N_18496,N_17393,N_16647);
nor U18497 (N_18497,N_15606,N_16819);
and U18498 (N_18498,N_16541,N_16368);
or U18499 (N_18499,N_16909,N_15047);
nand U18500 (N_18500,N_16338,N_16388);
and U18501 (N_18501,N_17279,N_16761);
nor U18502 (N_18502,N_17418,N_17164);
nand U18503 (N_18503,N_15810,N_15411);
xor U18504 (N_18504,N_16464,N_16956);
nor U18505 (N_18505,N_15686,N_17205);
nand U18506 (N_18506,N_16760,N_16271);
and U18507 (N_18507,N_16479,N_15027);
and U18508 (N_18508,N_16613,N_15112);
or U18509 (N_18509,N_16798,N_15079);
xnor U18510 (N_18510,N_16729,N_15970);
or U18511 (N_18511,N_17276,N_15445);
and U18512 (N_18512,N_16104,N_15785);
nand U18513 (N_18513,N_15130,N_15223);
nor U18514 (N_18514,N_15426,N_16160);
and U18515 (N_18515,N_16857,N_16791);
xor U18516 (N_18516,N_15256,N_16853);
nor U18517 (N_18517,N_16164,N_15689);
nor U18518 (N_18518,N_15778,N_15246);
xor U18519 (N_18519,N_15346,N_15397);
and U18520 (N_18520,N_15303,N_15933);
or U18521 (N_18521,N_16620,N_16008);
nand U18522 (N_18522,N_16609,N_15922);
xnor U18523 (N_18523,N_16840,N_16143);
nand U18524 (N_18524,N_17479,N_16827);
xor U18525 (N_18525,N_17207,N_17405);
nor U18526 (N_18526,N_17046,N_15661);
xnor U18527 (N_18527,N_17072,N_15038);
or U18528 (N_18528,N_17339,N_15227);
or U18529 (N_18529,N_17212,N_17474);
xnor U18530 (N_18530,N_16105,N_16032);
or U18531 (N_18531,N_17377,N_17432);
nand U18532 (N_18532,N_15490,N_16086);
and U18533 (N_18533,N_16462,N_15809);
xor U18534 (N_18534,N_17471,N_15160);
and U18535 (N_18535,N_16946,N_16491);
xor U18536 (N_18536,N_17495,N_16419);
xnor U18537 (N_18537,N_15984,N_16786);
and U18538 (N_18538,N_15624,N_15390);
xor U18539 (N_18539,N_15895,N_17034);
xor U18540 (N_18540,N_15306,N_17111);
or U18541 (N_18541,N_17167,N_15353);
nand U18542 (N_18542,N_16239,N_16954);
and U18543 (N_18543,N_16245,N_15045);
or U18544 (N_18544,N_15959,N_16646);
nand U18545 (N_18545,N_15729,N_15473);
and U18546 (N_18546,N_17008,N_15437);
or U18547 (N_18547,N_15041,N_15369);
and U18548 (N_18548,N_16851,N_16681);
or U18549 (N_18549,N_16551,N_16589);
nor U18550 (N_18550,N_15758,N_15094);
nand U18551 (N_18551,N_16809,N_16116);
nor U18552 (N_18552,N_15012,N_17228);
and U18553 (N_18553,N_15275,N_16757);
or U18554 (N_18554,N_16623,N_15236);
nor U18555 (N_18555,N_17124,N_15746);
nor U18556 (N_18556,N_15694,N_15385);
xor U18557 (N_18557,N_17102,N_16170);
nand U18558 (N_18558,N_15122,N_17150);
nand U18559 (N_18559,N_15107,N_15436);
nand U18560 (N_18560,N_16605,N_17041);
or U18561 (N_18561,N_15016,N_17480);
or U18562 (N_18562,N_16227,N_17372);
nor U18563 (N_18563,N_15191,N_16710);
xnor U18564 (N_18564,N_16989,N_16663);
nand U18565 (N_18565,N_15576,N_16237);
and U18566 (N_18566,N_15497,N_15059);
xor U18567 (N_18567,N_15585,N_16642);
and U18568 (N_18568,N_16731,N_17054);
nand U18569 (N_18569,N_15336,N_15773);
xnor U18570 (N_18570,N_15060,N_16345);
nor U18571 (N_18571,N_16991,N_16665);
nand U18572 (N_18572,N_15610,N_15869);
or U18573 (N_18573,N_15826,N_16506);
nor U18574 (N_18574,N_15880,N_16485);
and U18575 (N_18575,N_15046,N_15980);
nand U18576 (N_18576,N_15158,N_16874);
nand U18577 (N_18577,N_15419,N_16118);
or U18578 (N_18578,N_16509,N_16335);
nand U18579 (N_18579,N_16631,N_17447);
or U18580 (N_18580,N_16988,N_15974);
nand U18581 (N_18581,N_15114,N_16753);
nor U18582 (N_18582,N_16354,N_16525);
and U18583 (N_18583,N_16055,N_16370);
nand U18584 (N_18584,N_16701,N_15510);
nor U18585 (N_18585,N_15408,N_15945);
xnor U18586 (N_18586,N_15429,N_17053);
xor U18587 (N_18587,N_16377,N_15442);
or U18588 (N_18588,N_15457,N_17431);
xor U18589 (N_18589,N_17211,N_15020);
and U18590 (N_18590,N_17052,N_15669);
nand U18591 (N_18591,N_15233,N_15228);
nand U18592 (N_18592,N_16264,N_15043);
and U18593 (N_18593,N_15730,N_15239);
xnor U18594 (N_18594,N_16035,N_15675);
nor U18595 (N_18595,N_16481,N_15642);
nor U18596 (N_18596,N_16697,N_16090);
xnor U18597 (N_18597,N_15634,N_15464);
xor U18598 (N_18598,N_16360,N_15616);
nand U18599 (N_18599,N_15511,N_16875);
and U18600 (N_18600,N_17399,N_15573);
xor U18601 (N_18601,N_15268,N_16583);
nor U18602 (N_18602,N_16800,N_15009);
nor U18603 (N_18603,N_16816,N_17193);
xor U18604 (N_18604,N_16016,N_15693);
nor U18605 (N_18605,N_16003,N_16921);
or U18606 (N_18606,N_15190,N_16165);
nor U18607 (N_18607,N_15802,N_15877);
and U18608 (N_18608,N_16603,N_15209);
xor U18609 (N_18609,N_15799,N_15508);
and U18610 (N_18610,N_16077,N_17359);
or U18611 (N_18611,N_16139,N_17243);
nor U18612 (N_18612,N_15789,N_17229);
nand U18613 (N_18613,N_15243,N_15702);
nand U18614 (N_18614,N_16947,N_16998);
xor U18615 (N_18615,N_15425,N_16961);
nor U18616 (N_18616,N_15316,N_16175);
or U18617 (N_18617,N_17454,N_16865);
or U18618 (N_18618,N_16331,N_17362);
xor U18619 (N_18619,N_15072,N_15042);
nand U18620 (N_18620,N_16962,N_15990);
nor U18621 (N_18621,N_15289,N_16085);
xor U18622 (N_18622,N_15791,N_15884);
nor U18623 (N_18623,N_16768,N_15181);
or U18624 (N_18624,N_15673,N_17165);
nand U18625 (N_18625,N_15264,N_15771);
xor U18626 (N_18626,N_16389,N_16769);
or U18627 (N_18627,N_15172,N_16762);
nand U18628 (N_18628,N_16826,N_16510);
or U18629 (N_18629,N_17327,N_15170);
xnor U18630 (N_18630,N_16011,N_16877);
or U18631 (N_18631,N_15543,N_16019);
xnor U18632 (N_18632,N_15554,N_17135);
xor U18633 (N_18633,N_15715,N_16203);
nor U18634 (N_18634,N_16438,N_16065);
nand U18635 (N_18635,N_17186,N_17085);
or U18636 (N_18636,N_15168,N_15366);
and U18637 (N_18637,N_15388,N_15932);
nor U18638 (N_18638,N_16173,N_15372);
and U18639 (N_18639,N_15583,N_17100);
nand U18640 (N_18640,N_17038,N_15200);
nor U18641 (N_18641,N_17121,N_16279);
or U18642 (N_18642,N_15225,N_17114);
and U18643 (N_18643,N_15315,N_17350);
or U18644 (N_18644,N_16369,N_17353);
nor U18645 (N_18645,N_17429,N_15890);
and U18646 (N_18646,N_16560,N_17466);
or U18647 (N_18647,N_16806,N_16606);
nand U18648 (N_18648,N_16348,N_15954);
or U18649 (N_18649,N_15850,N_16523);
or U18650 (N_18650,N_15827,N_15738);
xor U18651 (N_18651,N_15533,N_15254);
nor U18652 (N_18652,N_15550,N_17017);
nand U18653 (N_18653,N_16054,N_16680);
and U18654 (N_18654,N_16983,N_15761);
or U18655 (N_18655,N_15966,N_17126);
xor U18656 (N_18656,N_15026,N_15357);
and U18657 (N_18657,N_15831,N_15558);
and U18658 (N_18658,N_17478,N_17284);
or U18659 (N_18659,N_16859,N_15166);
xnor U18660 (N_18660,N_15695,N_15972);
or U18661 (N_18661,N_15615,N_16127);
and U18662 (N_18662,N_15532,N_16895);
nor U18663 (N_18663,N_16734,N_17417);
nor U18664 (N_18664,N_16503,N_16452);
and U18665 (N_18665,N_15871,N_15308);
or U18666 (N_18666,N_15093,N_16880);
xnor U18667 (N_18667,N_15207,N_17305);
xor U18668 (N_18668,N_16802,N_17083);
or U18669 (N_18669,N_15119,N_15762);
xnor U18670 (N_18670,N_15636,N_16914);
or U18671 (N_18671,N_16399,N_16324);
nor U18672 (N_18672,N_16659,N_16269);
and U18673 (N_18673,N_16866,N_15908);
or U18674 (N_18674,N_16079,N_15024);
and U18675 (N_18675,N_15287,N_15286);
nand U18676 (N_18676,N_15341,N_15151);
xor U18677 (N_18677,N_16888,N_16600);
or U18678 (N_18678,N_16915,N_15244);
nor U18679 (N_18679,N_17143,N_15155);
or U18680 (N_18680,N_15839,N_17457);
xor U18681 (N_18681,N_16522,N_16650);
or U18682 (N_18682,N_16252,N_15136);
or U18683 (N_18683,N_16210,N_15102);
nand U18684 (N_18684,N_15459,N_15220);
or U18685 (N_18685,N_15134,N_15265);
nor U18686 (N_18686,N_16042,N_15280);
xor U18687 (N_18687,N_15821,N_15708);
nor U18688 (N_18688,N_16689,N_15710);
nor U18689 (N_18689,N_15659,N_16925);
xnor U18690 (N_18690,N_16856,N_16432);
nor U18691 (N_18691,N_16374,N_16158);
nor U18692 (N_18692,N_17337,N_15921);
nor U18693 (N_18693,N_16969,N_15817);
xor U18694 (N_18694,N_15276,N_15427);
nand U18695 (N_18695,N_17390,N_15468);
and U18696 (N_18696,N_15938,N_15942);
nand U18697 (N_18697,N_16402,N_15684);
nand U18698 (N_18698,N_16371,N_17409);
and U18699 (N_18699,N_15609,N_16611);
nand U18700 (N_18700,N_15076,N_15451);
or U18701 (N_18701,N_15917,N_16813);
or U18702 (N_18702,N_16281,N_15049);
nor U18703 (N_18703,N_15915,N_17325);
and U18704 (N_18704,N_17048,N_15098);
or U18705 (N_18705,N_15800,N_15764);
nand U18706 (N_18706,N_16144,N_16132);
or U18707 (N_18707,N_16458,N_15846);
xor U18708 (N_18708,N_16733,N_15951);
nand U18709 (N_18709,N_16656,N_17422);
nand U18710 (N_18710,N_17387,N_16287);
or U18711 (N_18711,N_16890,N_17225);
or U18712 (N_18712,N_15674,N_16639);
and U18713 (N_18713,N_16824,N_15755);
or U18714 (N_18714,N_15630,N_15657);
xnor U18715 (N_18715,N_16805,N_17400);
nor U18716 (N_18716,N_15721,N_15144);
nor U18717 (N_18717,N_16705,N_16057);
nor U18718 (N_18718,N_15769,N_16449);
or U18719 (N_18719,N_15187,N_15434);
nor U18720 (N_18720,N_15601,N_17345);
xor U18721 (N_18721,N_16192,N_15553);
or U18722 (N_18722,N_16141,N_16109);
and U18723 (N_18723,N_15816,N_15479);
nand U18724 (N_18724,N_16349,N_15250);
nand U18725 (N_18725,N_17299,N_15131);
nand U18726 (N_18726,N_15652,N_17129);
nor U18727 (N_18727,N_16238,N_16253);
xor U18728 (N_18728,N_15843,N_16558);
xnor U18729 (N_18729,N_16952,N_15998);
and U18730 (N_18730,N_15374,N_17449);
or U18731 (N_18731,N_17108,N_16726);
or U18732 (N_18732,N_16717,N_16575);
nor U18733 (N_18733,N_15983,N_17220);
xor U18734 (N_18734,N_15750,N_15633);
nor U18735 (N_18735,N_15484,N_16329);
and U18736 (N_18736,N_15861,N_15206);
nand U18737 (N_18737,N_15521,N_16072);
xor U18738 (N_18738,N_16049,N_16148);
xnor U18739 (N_18739,N_16489,N_17278);
and U18740 (N_18740,N_15500,N_15751);
or U18741 (N_18741,N_16929,N_15159);
nor U18742 (N_18742,N_15905,N_15879);
nor U18743 (N_18743,N_16448,N_16942);
nor U18744 (N_18744,N_15283,N_16764);
or U18745 (N_18745,N_17426,N_16453);
xor U18746 (N_18746,N_16579,N_15705);
nor U18747 (N_18747,N_17242,N_16420);
or U18748 (N_18748,N_15345,N_16671);
nor U18749 (N_18749,N_15567,N_15391);
or U18750 (N_18750,N_17113,N_15812);
nand U18751 (N_18751,N_16993,N_15685);
nand U18752 (N_18752,N_17425,N_15964);
nand U18753 (N_18753,N_16442,N_15793);
or U18754 (N_18754,N_16751,N_16285);
nand U18755 (N_18755,N_17019,N_17455);
xor U18756 (N_18756,N_16579,N_16886);
or U18757 (N_18757,N_16899,N_15669);
nand U18758 (N_18758,N_16571,N_16605);
xor U18759 (N_18759,N_16708,N_16095);
and U18760 (N_18760,N_17464,N_16692);
and U18761 (N_18761,N_15280,N_15539);
nor U18762 (N_18762,N_16913,N_17156);
and U18763 (N_18763,N_15428,N_15864);
nand U18764 (N_18764,N_15711,N_15316);
and U18765 (N_18765,N_17205,N_16984);
nand U18766 (N_18766,N_16989,N_16243);
or U18767 (N_18767,N_17482,N_16837);
nand U18768 (N_18768,N_15090,N_16949);
xnor U18769 (N_18769,N_16218,N_16882);
or U18770 (N_18770,N_15115,N_15779);
and U18771 (N_18771,N_16570,N_16763);
nand U18772 (N_18772,N_16924,N_17078);
nand U18773 (N_18773,N_15616,N_15144);
or U18774 (N_18774,N_15973,N_16467);
nand U18775 (N_18775,N_16481,N_17021);
nor U18776 (N_18776,N_16861,N_15512);
nor U18777 (N_18777,N_17390,N_15469);
xnor U18778 (N_18778,N_17431,N_16198);
xor U18779 (N_18779,N_16280,N_16220);
and U18780 (N_18780,N_16266,N_16612);
and U18781 (N_18781,N_16428,N_15375);
nor U18782 (N_18782,N_15569,N_15050);
and U18783 (N_18783,N_15747,N_16898);
nor U18784 (N_18784,N_15268,N_16175);
or U18785 (N_18785,N_17181,N_17494);
xor U18786 (N_18786,N_17058,N_17142);
nor U18787 (N_18787,N_15706,N_16715);
xnor U18788 (N_18788,N_16887,N_15461);
nand U18789 (N_18789,N_15205,N_16290);
nor U18790 (N_18790,N_16528,N_15838);
nand U18791 (N_18791,N_16036,N_15009);
or U18792 (N_18792,N_15817,N_15370);
or U18793 (N_18793,N_16032,N_17328);
and U18794 (N_18794,N_16234,N_17107);
and U18795 (N_18795,N_17055,N_17454);
xnor U18796 (N_18796,N_15721,N_16725);
or U18797 (N_18797,N_16782,N_16086);
nand U18798 (N_18798,N_17393,N_15172);
nor U18799 (N_18799,N_17043,N_15742);
nor U18800 (N_18800,N_16266,N_17237);
and U18801 (N_18801,N_16742,N_16039);
nor U18802 (N_18802,N_17023,N_16698);
xnor U18803 (N_18803,N_15599,N_15066);
nand U18804 (N_18804,N_16764,N_16156);
nand U18805 (N_18805,N_16015,N_16795);
xnor U18806 (N_18806,N_16143,N_16899);
nor U18807 (N_18807,N_15006,N_16037);
xnor U18808 (N_18808,N_15116,N_16186);
nor U18809 (N_18809,N_16847,N_16525);
nand U18810 (N_18810,N_15940,N_15740);
xnor U18811 (N_18811,N_15538,N_17170);
nor U18812 (N_18812,N_16560,N_16962);
and U18813 (N_18813,N_17472,N_15950);
or U18814 (N_18814,N_16911,N_15727);
nor U18815 (N_18815,N_17141,N_15250);
and U18816 (N_18816,N_17441,N_17313);
or U18817 (N_18817,N_16327,N_15785);
xor U18818 (N_18818,N_16462,N_17392);
nor U18819 (N_18819,N_16238,N_16465);
or U18820 (N_18820,N_16571,N_15371);
or U18821 (N_18821,N_16742,N_15864);
or U18822 (N_18822,N_17365,N_17217);
xnor U18823 (N_18823,N_15954,N_16804);
and U18824 (N_18824,N_17189,N_16135);
xnor U18825 (N_18825,N_15607,N_16430);
nand U18826 (N_18826,N_15712,N_16943);
nor U18827 (N_18827,N_16093,N_15625);
or U18828 (N_18828,N_15732,N_15266);
nand U18829 (N_18829,N_15192,N_15033);
and U18830 (N_18830,N_16181,N_17212);
xor U18831 (N_18831,N_16745,N_16844);
nor U18832 (N_18832,N_16909,N_16521);
nor U18833 (N_18833,N_15295,N_15241);
and U18834 (N_18834,N_16816,N_15751);
or U18835 (N_18835,N_17146,N_16646);
or U18836 (N_18836,N_15693,N_16645);
xnor U18837 (N_18837,N_15904,N_15848);
nor U18838 (N_18838,N_17248,N_17022);
xnor U18839 (N_18839,N_15433,N_17375);
nor U18840 (N_18840,N_16147,N_15311);
and U18841 (N_18841,N_17056,N_16466);
and U18842 (N_18842,N_15199,N_15261);
or U18843 (N_18843,N_16548,N_16857);
nor U18844 (N_18844,N_15419,N_16729);
xor U18845 (N_18845,N_16540,N_15698);
nand U18846 (N_18846,N_16943,N_15617);
xnor U18847 (N_18847,N_15688,N_16808);
nand U18848 (N_18848,N_16741,N_16582);
or U18849 (N_18849,N_15551,N_16537);
nor U18850 (N_18850,N_15192,N_17124);
nor U18851 (N_18851,N_17107,N_15140);
nand U18852 (N_18852,N_16406,N_16235);
or U18853 (N_18853,N_17363,N_17447);
nand U18854 (N_18854,N_15209,N_15675);
xnor U18855 (N_18855,N_16275,N_15576);
or U18856 (N_18856,N_16970,N_15401);
nand U18857 (N_18857,N_16728,N_17462);
nor U18858 (N_18858,N_17346,N_17009);
or U18859 (N_18859,N_15649,N_16985);
nor U18860 (N_18860,N_16308,N_17376);
nor U18861 (N_18861,N_17458,N_16766);
nand U18862 (N_18862,N_15604,N_16182);
xor U18863 (N_18863,N_16691,N_15404);
or U18864 (N_18864,N_17062,N_16093);
nand U18865 (N_18865,N_15833,N_15396);
nor U18866 (N_18866,N_16791,N_16945);
nand U18867 (N_18867,N_15760,N_15899);
or U18868 (N_18868,N_15721,N_16517);
nor U18869 (N_18869,N_15360,N_16573);
or U18870 (N_18870,N_15197,N_16662);
nor U18871 (N_18871,N_15640,N_15566);
and U18872 (N_18872,N_16498,N_16040);
or U18873 (N_18873,N_15375,N_15346);
and U18874 (N_18874,N_15351,N_15034);
nand U18875 (N_18875,N_17064,N_16777);
or U18876 (N_18876,N_15056,N_16953);
nor U18877 (N_18877,N_16115,N_15165);
nand U18878 (N_18878,N_16614,N_16849);
xor U18879 (N_18879,N_17290,N_16746);
nand U18880 (N_18880,N_15972,N_17378);
nor U18881 (N_18881,N_15833,N_16790);
nand U18882 (N_18882,N_16148,N_15098);
and U18883 (N_18883,N_15745,N_16167);
and U18884 (N_18884,N_15150,N_16576);
and U18885 (N_18885,N_16110,N_15641);
or U18886 (N_18886,N_17381,N_15298);
nor U18887 (N_18887,N_15300,N_15837);
nor U18888 (N_18888,N_15591,N_16471);
xnor U18889 (N_18889,N_16296,N_15627);
or U18890 (N_18890,N_15870,N_16446);
xnor U18891 (N_18891,N_15487,N_16962);
and U18892 (N_18892,N_16842,N_16093);
and U18893 (N_18893,N_16402,N_16217);
nand U18894 (N_18894,N_16510,N_15688);
and U18895 (N_18895,N_15679,N_15838);
nand U18896 (N_18896,N_15603,N_16529);
xnor U18897 (N_18897,N_16086,N_15918);
xor U18898 (N_18898,N_16135,N_15130);
and U18899 (N_18899,N_15448,N_16185);
nand U18900 (N_18900,N_15594,N_15707);
or U18901 (N_18901,N_16205,N_17290);
nand U18902 (N_18902,N_16378,N_16035);
nor U18903 (N_18903,N_15255,N_15000);
and U18904 (N_18904,N_16677,N_15234);
nor U18905 (N_18905,N_16529,N_16794);
nand U18906 (N_18906,N_16589,N_15200);
nor U18907 (N_18907,N_16273,N_15680);
nor U18908 (N_18908,N_16310,N_15374);
nor U18909 (N_18909,N_16280,N_17204);
or U18910 (N_18910,N_16696,N_16069);
and U18911 (N_18911,N_15547,N_17235);
xor U18912 (N_18912,N_15795,N_15932);
and U18913 (N_18913,N_16484,N_15517);
nand U18914 (N_18914,N_15551,N_15119);
and U18915 (N_18915,N_16308,N_15684);
and U18916 (N_18916,N_15232,N_17124);
nor U18917 (N_18917,N_15617,N_15878);
nand U18918 (N_18918,N_15495,N_16169);
nor U18919 (N_18919,N_15779,N_15553);
xnor U18920 (N_18920,N_15384,N_15373);
nand U18921 (N_18921,N_15352,N_15536);
xnor U18922 (N_18922,N_15859,N_16721);
and U18923 (N_18923,N_15711,N_15293);
or U18924 (N_18924,N_15369,N_15012);
nor U18925 (N_18925,N_16350,N_15825);
or U18926 (N_18926,N_15814,N_15899);
or U18927 (N_18927,N_17064,N_15919);
and U18928 (N_18928,N_16662,N_17484);
or U18929 (N_18929,N_15855,N_15754);
and U18930 (N_18930,N_16518,N_15265);
nand U18931 (N_18931,N_16414,N_16952);
nand U18932 (N_18932,N_16379,N_16314);
and U18933 (N_18933,N_16895,N_15844);
nand U18934 (N_18934,N_16934,N_17369);
and U18935 (N_18935,N_17003,N_17105);
nor U18936 (N_18936,N_17030,N_16902);
or U18937 (N_18937,N_16584,N_17061);
nand U18938 (N_18938,N_16511,N_15188);
nor U18939 (N_18939,N_15083,N_15993);
or U18940 (N_18940,N_17069,N_15070);
or U18941 (N_18941,N_16093,N_16084);
nand U18942 (N_18942,N_15967,N_15891);
xnor U18943 (N_18943,N_17043,N_15952);
or U18944 (N_18944,N_16721,N_15254);
nand U18945 (N_18945,N_16423,N_17454);
xor U18946 (N_18946,N_15798,N_15578);
and U18947 (N_18947,N_16902,N_15746);
nor U18948 (N_18948,N_16956,N_15545);
xor U18949 (N_18949,N_17184,N_15332);
or U18950 (N_18950,N_15988,N_16850);
nand U18951 (N_18951,N_17318,N_17482);
or U18952 (N_18952,N_16336,N_16016);
xnor U18953 (N_18953,N_16929,N_15846);
nand U18954 (N_18954,N_15438,N_15183);
nand U18955 (N_18955,N_15108,N_17468);
nor U18956 (N_18956,N_15488,N_16405);
or U18957 (N_18957,N_16239,N_15329);
xor U18958 (N_18958,N_16717,N_16108);
and U18959 (N_18959,N_15378,N_15683);
nand U18960 (N_18960,N_17346,N_17188);
and U18961 (N_18961,N_16583,N_16635);
or U18962 (N_18962,N_16868,N_16110);
nand U18963 (N_18963,N_15298,N_16209);
and U18964 (N_18964,N_16091,N_17017);
nor U18965 (N_18965,N_16742,N_15644);
nand U18966 (N_18966,N_17207,N_16524);
nand U18967 (N_18967,N_16821,N_16957);
xnor U18968 (N_18968,N_15553,N_15633);
and U18969 (N_18969,N_15665,N_15593);
and U18970 (N_18970,N_16860,N_16648);
xor U18971 (N_18971,N_17273,N_15489);
nor U18972 (N_18972,N_17332,N_16895);
nor U18973 (N_18973,N_16718,N_15851);
and U18974 (N_18974,N_17349,N_16498);
and U18975 (N_18975,N_15622,N_17070);
nor U18976 (N_18976,N_15976,N_16069);
or U18977 (N_18977,N_16924,N_16077);
nand U18978 (N_18978,N_15194,N_16684);
or U18979 (N_18979,N_17315,N_16570);
or U18980 (N_18980,N_17346,N_16037);
nand U18981 (N_18981,N_15767,N_15251);
nand U18982 (N_18982,N_16770,N_15325);
xor U18983 (N_18983,N_16443,N_16123);
and U18984 (N_18984,N_16360,N_17365);
nor U18985 (N_18985,N_16399,N_15118);
nand U18986 (N_18986,N_17103,N_15603);
nor U18987 (N_18987,N_16807,N_17310);
or U18988 (N_18988,N_17345,N_17204);
and U18989 (N_18989,N_16900,N_15866);
and U18990 (N_18990,N_15218,N_15948);
nor U18991 (N_18991,N_15240,N_17059);
and U18992 (N_18992,N_16777,N_15076);
nand U18993 (N_18993,N_17381,N_17177);
nand U18994 (N_18994,N_15385,N_16448);
nor U18995 (N_18995,N_15158,N_16696);
nand U18996 (N_18996,N_16775,N_15350);
nor U18997 (N_18997,N_15679,N_17145);
xor U18998 (N_18998,N_16905,N_16901);
xnor U18999 (N_18999,N_15927,N_15349);
and U19000 (N_19000,N_17221,N_15605);
xnor U19001 (N_19001,N_16408,N_16499);
xor U19002 (N_19002,N_16535,N_16828);
or U19003 (N_19003,N_15893,N_16382);
or U19004 (N_19004,N_15672,N_15950);
xor U19005 (N_19005,N_16987,N_15140);
or U19006 (N_19006,N_15164,N_16530);
nand U19007 (N_19007,N_15858,N_17388);
xnor U19008 (N_19008,N_16981,N_15255);
or U19009 (N_19009,N_17070,N_16322);
nor U19010 (N_19010,N_15611,N_15955);
or U19011 (N_19011,N_17058,N_15309);
xnor U19012 (N_19012,N_15957,N_17118);
nand U19013 (N_19013,N_16681,N_16722);
nor U19014 (N_19014,N_15751,N_16218);
nand U19015 (N_19015,N_16985,N_15837);
xnor U19016 (N_19016,N_15273,N_15582);
nand U19017 (N_19017,N_15788,N_16978);
xnor U19018 (N_19018,N_15508,N_15590);
and U19019 (N_19019,N_15786,N_16718);
nor U19020 (N_19020,N_15304,N_15757);
nor U19021 (N_19021,N_15041,N_17469);
or U19022 (N_19022,N_16045,N_16217);
xnor U19023 (N_19023,N_15368,N_16100);
and U19024 (N_19024,N_16851,N_15263);
xnor U19025 (N_19025,N_17117,N_16319);
or U19026 (N_19026,N_15401,N_15624);
nor U19027 (N_19027,N_16309,N_16004);
nor U19028 (N_19028,N_16542,N_15802);
or U19029 (N_19029,N_15765,N_15111);
nand U19030 (N_19030,N_15711,N_15897);
xnor U19031 (N_19031,N_17242,N_16780);
nor U19032 (N_19032,N_16667,N_16572);
nor U19033 (N_19033,N_16522,N_17421);
nand U19034 (N_19034,N_17492,N_15355);
nand U19035 (N_19035,N_16006,N_16179);
nand U19036 (N_19036,N_15196,N_16875);
nand U19037 (N_19037,N_15198,N_17493);
nand U19038 (N_19038,N_17423,N_15933);
and U19039 (N_19039,N_16817,N_15943);
nor U19040 (N_19040,N_15679,N_15676);
nor U19041 (N_19041,N_17157,N_16429);
or U19042 (N_19042,N_15012,N_16813);
and U19043 (N_19043,N_16473,N_15507);
nor U19044 (N_19044,N_15696,N_17411);
xor U19045 (N_19045,N_15882,N_16507);
nor U19046 (N_19046,N_15501,N_16041);
xnor U19047 (N_19047,N_17366,N_16986);
nor U19048 (N_19048,N_16636,N_16164);
xnor U19049 (N_19049,N_15647,N_16439);
and U19050 (N_19050,N_15120,N_16750);
nand U19051 (N_19051,N_16032,N_15179);
xnor U19052 (N_19052,N_16928,N_17260);
and U19053 (N_19053,N_17344,N_15805);
or U19054 (N_19054,N_16208,N_16408);
or U19055 (N_19055,N_16104,N_15362);
xnor U19056 (N_19056,N_17043,N_15939);
and U19057 (N_19057,N_17300,N_17249);
nor U19058 (N_19058,N_15958,N_16998);
xnor U19059 (N_19059,N_15276,N_15447);
and U19060 (N_19060,N_16892,N_15436);
nand U19061 (N_19061,N_16596,N_16538);
nand U19062 (N_19062,N_15334,N_15288);
nor U19063 (N_19063,N_17468,N_15596);
or U19064 (N_19064,N_15009,N_15965);
xor U19065 (N_19065,N_16777,N_15924);
xnor U19066 (N_19066,N_16038,N_15773);
nor U19067 (N_19067,N_15291,N_15487);
xnor U19068 (N_19068,N_15156,N_16544);
xnor U19069 (N_19069,N_17085,N_16782);
and U19070 (N_19070,N_15333,N_15557);
or U19071 (N_19071,N_17247,N_17032);
nor U19072 (N_19072,N_17018,N_16452);
nand U19073 (N_19073,N_15717,N_15943);
xnor U19074 (N_19074,N_16931,N_15956);
and U19075 (N_19075,N_16238,N_17135);
nand U19076 (N_19076,N_16793,N_17067);
or U19077 (N_19077,N_17121,N_16475);
or U19078 (N_19078,N_17227,N_15944);
or U19079 (N_19079,N_15902,N_16617);
or U19080 (N_19080,N_16745,N_15688);
nor U19081 (N_19081,N_15973,N_15366);
nand U19082 (N_19082,N_15473,N_16032);
nor U19083 (N_19083,N_15953,N_17134);
and U19084 (N_19084,N_15673,N_15624);
nor U19085 (N_19085,N_16216,N_16351);
xor U19086 (N_19086,N_15002,N_16032);
and U19087 (N_19087,N_16403,N_16855);
nand U19088 (N_19088,N_16443,N_15529);
and U19089 (N_19089,N_16613,N_16697);
nand U19090 (N_19090,N_17095,N_16292);
nand U19091 (N_19091,N_15844,N_17064);
or U19092 (N_19092,N_15184,N_17278);
nand U19093 (N_19093,N_16393,N_16454);
nand U19094 (N_19094,N_15091,N_16131);
or U19095 (N_19095,N_16281,N_15014);
or U19096 (N_19096,N_15820,N_16988);
xnor U19097 (N_19097,N_17112,N_16430);
or U19098 (N_19098,N_17204,N_17297);
xnor U19099 (N_19099,N_15463,N_17460);
or U19100 (N_19100,N_15778,N_17054);
and U19101 (N_19101,N_15323,N_17077);
or U19102 (N_19102,N_17393,N_15309);
nor U19103 (N_19103,N_15533,N_17236);
xnor U19104 (N_19104,N_16172,N_17061);
nand U19105 (N_19105,N_16582,N_15738);
xor U19106 (N_19106,N_17095,N_16320);
nor U19107 (N_19107,N_16097,N_15305);
nor U19108 (N_19108,N_16562,N_17010);
nand U19109 (N_19109,N_15372,N_16216);
nand U19110 (N_19110,N_17231,N_16209);
nor U19111 (N_19111,N_16848,N_16681);
or U19112 (N_19112,N_16532,N_16577);
nor U19113 (N_19113,N_15415,N_16801);
xnor U19114 (N_19114,N_15164,N_15968);
or U19115 (N_19115,N_16659,N_16538);
nand U19116 (N_19116,N_16441,N_16921);
or U19117 (N_19117,N_16298,N_15945);
xnor U19118 (N_19118,N_16574,N_16470);
or U19119 (N_19119,N_17193,N_16457);
nor U19120 (N_19120,N_15398,N_15925);
and U19121 (N_19121,N_15814,N_16298);
xor U19122 (N_19122,N_16540,N_17493);
nand U19123 (N_19123,N_16415,N_15681);
and U19124 (N_19124,N_15015,N_17301);
and U19125 (N_19125,N_17238,N_15590);
or U19126 (N_19126,N_16741,N_17313);
nand U19127 (N_19127,N_16464,N_15509);
nor U19128 (N_19128,N_16971,N_17064);
nand U19129 (N_19129,N_16267,N_16775);
and U19130 (N_19130,N_17342,N_15618);
or U19131 (N_19131,N_15119,N_16319);
nor U19132 (N_19132,N_16990,N_17052);
xor U19133 (N_19133,N_16134,N_16979);
xor U19134 (N_19134,N_15758,N_16572);
and U19135 (N_19135,N_15757,N_15126);
and U19136 (N_19136,N_15590,N_15983);
xnor U19137 (N_19137,N_15996,N_15433);
and U19138 (N_19138,N_15883,N_16934);
xor U19139 (N_19139,N_16296,N_17324);
xor U19140 (N_19140,N_15800,N_15703);
or U19141 (N_19141,N_17060,N_17013);
and U19142 (N_19142,N_15496,N_16778);
or U19143 (N_19143,N_17267,N_17144);
xor U19144 (N_19144,N_17077,N_16797);
nor U19145 (N_19145,N_17209,N_17123);
nor U19146 (N_19146,N_16896,N_16619);
nand U19147 (N_19147,N_16484,N_15814);
nand U19148 (N_19148,N_15100,N_15858);
xor U19149 (N_19149,N_16869,N_16379);
xor U19150 (N_19150,N_16347,N_16287);
xor U19151 (N_19151,N_15544,N_15766);
nor U19152 (N_19152,N_16284,N_15683);
nand U19153 (N_19153,N_15492,N_16149);
xnor U19154 (N_19154,N_15336,N_15404);
xnor U19155 (N_19155,N_15008,N_16333);
nand U19156 (N_19156,N_15434,N_16581);
or U19157 (N_19157,N_15851,N_15328);
or U19158 (N_19158,N_15931,N_16858);
nor U19159 (N_19159,N_15978,N_16187);
nor U19160 (N_19160,N_15167,N_15383);
xnor U19161 (N_19161,N_17122,N_17339);
or U19162 (N_19162,N_17130,N_15512);
nor U19163 (N_19163,N_17236,N_16962);
nor U19164 (N_19164,N_15202,N_16468);
nor U19165 (N_19165,N_16563,N_16748);
or U19166 (N_19166,N_15662,N_17235);
xnor U19167 (N_19167,N_16042,N_15597);
xor U19168 (N_19168,N_15457,N_15744);
and U19169 (N_19169,N_15626,N_17335);
or U19170 (N_19170,N_15295,N_15397);
and U19171 (N_19171,N_16972,N_16388);
xor U19172 (N_19172,N_15791,N_16743);
xor U19173 (N_19173,N_15022,N_16781);
nand U19174 (N_19174,N_15791,N_17030);
nand U19175 (N_19175,N_15942,N_16698);
nand U19176 (N_19176,N_16354,N_15481);
nor U19177 (N_19177,N_16911,N_16208);
and U19178 (N_19178,N_16366,N_15509);
or U19179 (N_19179,N_16184,N_16136);
nand U19180 (N_19180,N_15485,N_17288);
xor U19181 (N_19181,N_16832,N_16969);
nand U19182 (N_19182,N_16270,N_16057);
and U19183 (N_19183,N_16725,N_16564);
xnor U19184 (N_19184,N_16515,N_15995);
and U19185 (N_19185,N_15365,N_15132);
xor U19186 (N_19186,N_15980,N_15541);
or U19187 (N_19187,N_15416,N_16804);
nand U19188 (N_19188,N_16426,N_15572);
nor U19189 (N_19189,N_16810,N_16982);
xnor U19190 (N_19190,N_15442,N_16031);
nand U19191 (N_19191,N_16949,N_15933);
and U19192 (N_19192,N_16327,N_16633);
xnor U19193 (N_19193,N_17452,N_17464);
xor U19194 (N_19194,N_15822,N_16422);
xor U19195 (N_19195,N_17422,N_16145);
or U19196 (N_19196,N_15645,N_16319);
nor U19197 (N_19197,N_15058,N_16947);
nand U19198 (N_19198,N_15338,N_15470);
xnor U19199 (N_19199,N_16617,N_17115);
nor U19200 (N_19200,N_15416,N_15920);
and U19201 (N_19201,N_15808,N_15379);
xnor U19202 (N_19202,N_16260,N_16003);
or U19203 (N_19203,N_15110,N_17089);
or U19204 (N_19204,N_15001,N_15553);
xnor U19205 (N_19205,N_15838,N_16438);
xor U19206 (N_19206,N_17292,N_16479);
nor U19207 (N_19207,N_16350,N_15993);
and U19208 (N_19208,N_17046,N_15943);
or U19209 (N_19209,N_17123,N_16957);
nor U19210 (N_19210,N_15398,N_15288);
xnor U19211 (N_19211,N_15405,N_16107);
or U19212 (N_19212,N_15669,N_16735);
xnor U19213 (N_19213,N_17211,N_16633);
nor U19214 (N_19214,N_17412,N_16434);
and U19215 (N_19215,N_15705,N_15631);
nor U19216 (N_19216,N_16490,N_15812);
or U19217 (N_19217,N_15848,N_17260);
nor U19218 (N_19218,N_17073,N_15459);
nand U19219 (N_19219,N_16491,N_15803);
and U19220 (N_19220,N_15308,N_16140);
nor U19221 (N_19221,N_15279,N_16255);
nand U19222 (N_19222,N_15333,N_16553);
or U19223 (N_19223,N_16682,N_15526);
nand U19224 (N_19224,N_17236,N_15786);
and U19225 (N_19225,N_17317,N_15664);
and U19226 (N_19226,N_16350,N_16657);
xnor U19227 (N_19227,N_16968,N_15841);
nor U19228 (N_19228,N_17206,N_15151);
or U19229 (N_19229,N_17132,N_15489);
nor U19230 (N_19230,N_15366,N_15147);
and U19231 (N_19231,N_15916,N_16895);
or U19232 (N_19232,N_16936,N_16649);
nand U19233 (N_19233,N_16172,N_16678);
and U19234 (N_19234,N_16937,N_17494);
xor U19235 (N_19235,N_17489,N_15730);
nor U19236 (N_19236,N_15654,N_16371);
nand U19237 (N_19237,N_16291,N_15649);
nor U19238 (N_19238,N_15363,N_17490);
nand U19239 (N_19239,N_16835,N_17226);
or U19240 (N_19240,N_15646,N_15740);
or U19241 (N_19241,N_15909,N_16591);
nor U19242 (N_19242,N_15735,N_15323);
xor U19243 (N_19243,N_15200,N_16905);
and U19244 (N_19244,N_15406,N_15507);
nor U19245 (N_19245,N_15801,N_16949);
or U19246 (N_19246,N_16348,N_16746);
and U19247 (N_19247,N_16717,N_17307);
xnor U19248 (N_19248,N_16186,N_15893);
or U19249 (N_19249,N_16924,N_17086);
xnor U19250 (N_19250,N_17031,N_15191);
or U19251 (N_19251,N_16448,N_15057);
nand U19252 (N_19252,N_16788,N_16378);
or U19253 (N_19253,N_15509,N_15674);
nor U19254 (N_19254,N_15704,N_16456);
nand U19255 (N_19255,N_16155,N_15345);
nand U19256 (N_19256,N_17033,N_15693);
nor U19257 (N_19257,N_16314,N_16711);
nor U19258 (N_19258,N_17405,N_17146);
xor U19259 (N_19259,N_16776,N_15091);
nand U19260 (N_19260,N_16267,N_16389);
xor U19261 (N_19261,N_15165,N_17184);
and U19262 (N_19262,N_16876,N_17207);
xor U19263 (N_19263,N_15395,N_16902);
or U19264 (N_19264,N_17452,N_15708);
or U19265 (N_19265,N_16124,N_15464);
nor U19266 (N_19266,N_16281,N_16231);
nand U19267 (N_19267,N_15852,N_16546);
nor U19268 (N_19268,N_17430,N_15619);
xor U19269 (N_19269,N_15920,N_15987);
nand U19270 (N_19270,N_16199,N_16962);
and U19271 (N_19271,N_16066,N_15603);
or U19272 (N_19272,N_15249,N_16224);
and U19273 (N_19273,N_17376,N_16361);
nor U19274 (N_19274,N_15795,N_16392);
nand U19275 (N_19275,N_16922,N_16144);
and U19276 (N_19276,N_15940,N_16139);
or U19277 (N_19277,N_16498,N_15894);
and U19278 (N_19278,N_17250,N_16726);
xor U19279 (N_19279,N_17031,N_16499);
nor U19280 (N_19280,N_15946,N_15833);
xor U19281 (N_19281,N_15155,N_15925);
or U19282 (N_19282,N_15892,N_15994);
xor U19283 (N_19283,N_15447,N_15637);
or U19284 (N_19284,N_15025,N_15240);
nand U19285 (N_19285,N_16260,N_16972);
or U19286 (N_19286,N_16209,N_15277);
or U19287 (N_19287,N_15127,N_16602);
or U19288 (N_19288,N_16188,N_16194);
nor U19289 (N_19289,N_15800,N_15077);
or U19290 (N_19290,N_17494,N_16753);
nor U19291 (N_19291,N_15097,N_17049);
or U19292 (N_19292,N_16790,N_16480);
xnor U19293 (N_19293,N_16511,N_15418);
nor U19294 (N_19294,N_17041,N_15638);
and U19295 (N_19295,N_15625,N_16016);
and U19296 (N_19296,N_16287,N_16786);
and U19297 (N_19297,N_15575,N_16372);
xnor U19298 (N_19298,N_16605,N_16623);
nor U19299 (N_19299,N_15573,N_16878);
nand U19300 (N_19300,N_16879,N_15072);
nand U19301 (N_19301,N_16531,N_15109);
xnor U19302 (N_19302,N_17291,N_16826);
xnor U19303 (N_19303,N_16992,N_15705);
nand U19304 (N_19304,N_17068,N_15803);
and U19305 (N_19305,N_17047,N_17046);
and U19306 (N_19306,N_16796,N_17286);
nand U19307 (N_19307,N_15248,N_16725);
nor U19308 (N_19308,N_15389,N_15658);
nor U19309 (N_19309,N_15449,N_15962);
xnor U19310 (N_19310,N_15155,N_16848);
xor U19311 (N_19311,N_17229,N_17423);
and U19312 (N_19312,N_15614,N_16588);
xnor U19313 (N_19313,N_15787,N_17166);
xnor U19314 (N_19314,N_15888,N_15028);
or U19315 (N_19315,N_15982,N_16955);
and U19316 (N_19316,N_15944,N_16144);
nand U19317 (N_19317,N_15899,N_16394);
nand U19318 (N_19318,N_15019,N_16297);
or U19319 (N_19319,N_16808,N_15802);
nand U19320 (N_19320,N_16607,N_15502);
and U19321 (N_19321,N_15962,N_15916);
and U19322 (N_19322,N_15069,N_15638);
nor U19323 (N_19323,N_17006,N_17412);
nor U19324 (N_19324,N_16467,N_16749);
nor U19325 (N_19325,N_15764,N_15861);
and U19326 (N_19326,N_15084,N_17057);
and U19327 (N_19327,N_16942,N_15517);
and U19328 (N_19328,N_15787,N_15340);
xnor U19329 (N_19329,N_16747,N_17304);
nor U19330 (N_19330,N_17175,N_16288);
xnor U19331 (N_19331,N_16752,N_16387);
nand U19332 (N_19332,N_15342,N_17395);
and U19333 (N_19333,N_15139,N_17180);
or U19334 (N_19334,N_16750,N_17301);
nand U19335 (N_19335,N_16013,N_16127);
or U19336 (N_19336,N_17341,N_16519);
and U19337 (N_19337,N_16546,N_16538);
nand U19338 (N_19338,N_17084,N_15937);
nand U19339 (N_19339,N_16620,N_15520);
nand U19340 (N_19340,N_15020,N_15276);
xor U19341 (N_19341,N_16362,N_15714);
xnor U19342 (N_19342,N_15047,N_15267);
or U19343 (N_19343,N_15031,N_17336);
nor U19344 (N_19344,N_15136,N_16553);
nor U19345 (N_19345,N_15007,N_15705);
nand U19346 (N_19346,N_15519,N_17274);
nor U19347 (N_19347,N_17317,N_15659);
nor U19348 (N_19348,N_15996,N_15021);
nand U19349 (N_19349,N_16313,N_16916);
nor U19350 (N_19350,N_17054,N_15234);
or U19351 (N_19351,N_15639,N_16671);
and U19352 (N_19352,N_17270,N_15217);
or U19353 (N_19353,N_15560,N_16393);
or U19354 (N_19354,N_16820,N_15082);
nand U19355 (N_19355,N_16823,N_16731);
nor U19356 (N_19356,N_15075,N_16470);
nand U19357 (N_19357,N_16207,N_15828);
or U19358 (N_19358,N_17197,N_16985);
or U19359 (N_19359,N_16591,N_16616);
or U19360 (N_19360,N_17406,N_15396);
or U19361 (N_19361,N_15249,N_15131);
or U19362 (N_19362,N_15358,N_16052);
and U19363 (N_19363,N_16294,N_15080);
nor U19364 (N_19364,N_16449,N_17468);
nand U19365 (N_19365,N_16497,N_15606);
xnor U19366 (N_19366,N_16057,N_15256);
and U19367 (N_19367,N_15943,N_16382);
and U19368 (N_19368,N_16212,N_16749);
xor U19369 (N_19369,N_16543,N_15413);
and U19370 (N_19370,N_15248,N_17178);
and U19371 (N_19371,N_16689,N_15912);
xnor U19372 (N_19372,N_17248,N_17353);
or U19373 (N_19373,N_16418,N_16229);
xnor U19374 (N_19374,N_15047,N_16443);
xnor U19375 (N_19375,N_17168,N_15000);
xnor U19376 (N_19376,N_15658,N_15416);
nor U19377 (N_19377,N_15121,N_15858);
nor U19378 (N_19378,N_15615,N_17070);
and U19379 (N_19379,N_16495,N_16368);
nand U19380 (N_19380,N_15873,N_16242);
nor U19381 (N_19381,N_15196,N_16620);
nor U19382 (N_19382,N_16601,N_17439);
nor U19383 (N_19383,N_16953,N_16701);
nand U19384 (N_19384,N_15027,N_15530);
xnor U19385 (N_19385,N_17097,N_17013);
nor U19386 (N_19386,N_17211,N_15472);
xor U19387 (N_19387,N_15932,N_17439);
nor U19388 (N_19388,N_17259,N_17108);
nor U19389 (N_19389,N_16340,N_15047);
nand U19390 (N_19390,N_15544,N_16268);
or U19391 (N_19391,N_16817,N_16825);
and U19392 (N_19392,N_16632,N_16421);
or U19393 (N_19393,N_16397,N_16410);
or U19394 (N_19394,N_16355,N_16831);
or U19395 (N_19395,N_16108,N_16757);
or U19396 (N_19396,N_17010,N_17438);
nor U19397 (N_19397,N_15426,N_16511);
xor U19398 (N_19398,N_16296,N_15706);
or U19399 (N_19399,N_16524,N_16850);
and U19400 (N_19400,N_17214,N_16562);
xnor U19401 (N_19401,N_16463,N_16958);
nor U19402 (N_19402,N_17373,N_15880);
nor U19403 (N_19403,N_15636,N_16273);
xnor U19404 (N_19404,N_15276,N_16618);
and U19405 (N_19405,N_16147,N_15678);
nor U19406 (N_19406,N_15999,N_16969);
nor U19407 (N_19407,N_16296,N_15400);
nand U19408 (N_19408,N_16679,N_17279);
or U19409 (N_19409,N_15918,N_15247);
nor U19410 (N_19410,N_17098,N_17099);
or U19411 (N_19411,N_15419,N_16122);
and U19412 (N_19412,N_15659,N_17249);
xnor U19413 (N_19413,N_15842,N_16682);
xor U19414 (N_19414,N_15608,N_16821);
and U19415 (N_19415,N_17185,N_17251);
nor U19416 (N_19416,N_15698,N_16061);
nand U19417 (N_19417,N_15120,N_15819);
nand U19418 (N_19418,N_16711,N_15000);
xor U19419 (N_19419,N_15773,N_15154);
and U19420 (N_19420,N_15132,N_16923);
xor U19421 (N_19421,N_17295,N_17305);
nand U19422 (N_19422,N_16653,N_16792);
nand U19423 (N_19423,N_16082,N_16204);
and U19424 (N_19424,N_16368,N_17159);
and U19425 (N_19425,N_15387,N_17269);
nand U19426 (N_19426,N_17237,N_16533);
xnor U19427 (N_19427,N_15701,N_15740);
xor U19428 (N_19428,N_17332,N_16340);
nand U19429 (N_19429,N_16240,N_15751);
nor U19430 (N_19430,N_15366,N_15198);
and U19431 (N_19431,N_16405,N_16174);
nor U19432 (N_19432,N_16192,N_15084);
xor U19433 (N_19433,N_17042,N_15017);
and U19434 (N_19434,N_16232,N_16072);
and U19435 (N_19435,N_15744,N_16850);
nand U19436 (N_19436,N_15853,N_15911);
nor U19437 (N_19437,N_15603,N_17443);
xnor U19438 (N_19438,N_15645,N_15974);
nand U19439 (N_19439,N_16213,N_15493);
nor U19440 (N_19440,N_15780,N_17083);
and U19441 (N_19441,N_17166,N_15294);
or U19442 (N_19442,N_17300,N_17175);
nor U19443 (N_19443,N_15258,N_16773);
nor U19444 (N_19444,N_15696,N_15846);
nand U19445 (N_19445,N_16999,N_16544);
and U19446 (N_19446,N_16278,N_17411);
xnor U19447 (N_19447,N_16533,N_15840);
nor U19448 (N_19448,N_15253,N_15885);
xor U19449 (N_19449,N_16139,N_16831);
nor U19450 (N_19450,N_17277,N_17076);
nor U19451 (N_19451,N_15258,N_16542);
and U19452 (N_19452,N_15436,N_15298);
or U19453 (N_19453,N_17349,N_16182);
or U19454 (N_19454,N_17100,N_15160);
and U19455 (N_19455,N_16873,N_16784);
nor U19456 (N_19456,N_17166,N_15744);
and U19457 (N_19457,N_16403,N_16983);
and U19458 (N_19458,N_15754,N_15932);
nor U19459 (N_19459,N_16049,N_16163);
nand U19460 (N_19460,N_17348,N_16470);
and U19461 (N_19461,N_15804,N_16261);
or U19462 (N_19462,N_16627,N_15989);
nand U19463 (N_19463,N_15061,N_16612);
nand U19464 (N_19464,N_17162,N_17148);
nand U19465 (N_19465,N_16330,N_15061);
nor U19466 (N_19466,N_15626,N_16562);
and U19467 (N_19467,N_15843,N_16114);
xor U19468 (N_19468,N_16573,N_16482);
nor U19469 (N_19469,N_17494,N_15939);
nor U19470 (N_19470,N_17169,N_17207);
and U19471 (N_19471,N_17326,N_15217);
nand U19472 (N_19472,N_15702,N_16521);
nor U19473 (N_19473,N_17045,N_15360);
and U19474 (N_19474,N_15032,N_16054);
or U19475 (N_19475,N_15484,N_16795);
and U19476 (N_19476,N_15298,N_16561);
nor U19477 (N_19477,N_16279,N_15580);
nor U19478 (N_19478,N_16101,N_15998);
nor U19479 (N_19479,N_17193,N_16906);
and U19480 (N_19480,N_16042,N_17375);
nor U19481 (N_19481,N_17310,N_15962);
xnor U19482 (N_19482,N_17303,N_15970);
nand U19483 (N_19483,N_16188,N_15935);
or U19484 (N_19484,N_15877,N_16246);
xor U19485 (N_19485,N_16813,N_16859);
and U19486 (N_19486,N_16956,N_15385);
nand U19487 (N_19487,N_17016,N_17194);
xnor U19488 (N_19488,N_15020,N_16697);
nand U19489 (N_19489,N_16318,N_15212);
or U19490 (N_19490,N_15097,N_16874);
and U19491 (N_19491,N_15352,N_16852);
or U19492 (N_19492,N_17106,N_17336);
nor U19493 (N_19493,N_15746,N_16387);
and U19494 (N_19494,N_15948,N_15190);
nor U19495 (N_19495,N_17297,N_15450);
xnor U19496 (N_19496,N_16594,N_15846);
and U19497 (N_19497,N_17013,N_15461);
xnor U19498 (N_19498,N_16496,N_16781);
nand U19499 (N_19499,N_15839,N_17335);
xnor U19500 (N_19500,N_15496,N_16196);
xor U19501 (N_19501,N_15612,N_17190);
or U19502 (N_19502,N_15045,N_16971);
nor U19503 (N_19503,N_16555,N_17159);
nand U19504 (N_19504,N_15622,N_15620);
nand U19505 (N_19505,N_16738,N_16868);
nor U19506 (N_19506,N_17165,N_15598);
nand U19507 (N_19507,N_15305,N_16952);
nor U19508 (N_19508,N_15297,N_16393);
xor U19509 (N_19509,N_16389,N_15440);
and U19510 (N_19510,N_16998,N_15683);
xnor U19511 (N_19511,N_15417,N_16754);
xor U19512 (N_19512,N_17353,N_15091);
and U19513 (N_19513,N_15619,N_16742);
and U19514 (N_19514,N_15364,N_15098);
and U19515 (N_19515,N_17140,N_15965);
nand U19516 (N_19516,N_15855,N_15895);
nor U19517 (N_19517,N_15248,N_15629);
nor U19518 (N_19518,N_17479,N_15478);
nand U19519 (N_19519,N_15857,N_15235);
nand U19520 (N_19520,N_15947,N_17218);
or U19521 (N_19521,N_15936,N_15918);
xnor U19522 (N_19522,N_16439,N_15548);
nor U19523 (N_19523,N_17214,N_15469);
xnor U19524 (N_19524,N_15707,N_17234);
xnor U19525 (N_19525,N_16422,N_17434);
and U19526 (N_19526,N_16027,N_17051);
xor U19527 (N_19527,N_15133,N_17224);
nor U19528 (N_19528,N_15841,N_16614);
nand U19529 (N_19529,N_16150,N_15170);
nand U19530 (N_19530,N_15865,N_16907);
xor U19531 (N_19531,N_15969,N_17374);
nand U19532 (N_19532,N_15322,N_15267);
xor U19533 (N_19533,N_16066,N_16709);
or U19534 (N_19534,N_15778,N_17475);
or U19535 (N_19535,N_17313,N_16456);
xor U19536 (N_19536,N_15947,N_15637);
and U19537 (N_19537,N_16511,N_15518);
or U19538 (N_19538,N_15951,N_16401);
nand U19539 (N_19539,N_17254,N_16545);
and U19540 (N_19540,N_15165,N_15480);
nor U19541 (N_19541,N_17192,N_15268);
nor U19542 (N_19542,N_16338,N_15770);
and U19543 (N_19543,N_16460,N_16314);
xor U19544 (N_19544,N_15695,N_16706);
nor U19545 (N_19545,N_16643,N_15285);
or U19546 (N_19546,N_15496,N_16490);
and U19547 (N_19547,N_15061,N_17117);
or U19548 (N_19548,N_16481,N_17246);
or U19549 (N_19549,N_16228,N_16811);
nor U19550 (N_19550,N_17147,N_16995);
and U19551 (N_19551,N_17467,N_15820);
nand U19552 (N_19552,N_15663,N_17428);
xor U19553 (N_19553,N_15442,N_16244);
and U19554 (N_19554,N_17258,N_15598);
and U19555 (N_19555,N_15813,N_17330);
and U19556 (N_19556,N_15831,N_16759);
or U19557 (N_19557,N_16145,N_17294);
nand U19558 (N_19558,N_17150,N_16268);
nand U19559 (N_19559,N_17064,N_15826);
nor U19560 (N_19560,N_15841,N_15324);
xor U19561 (N_19561,N_15670,N_15264);
xnor U19562 (N_19562,N_15561,N_16568);
or U19563 (N_19563,N_16831,N_15815);
xor U19564 (N_19564,N_15212,N_15537);
nor U19565 (N_19565,N_16206,N_16911);
nor U19566 (N_19566,N_15408,N_16689);
nor U19567 (N_19567,N_16800,N_15303);
or U19568 (N_19568,N_17168,N_16911);
xor U19569 (N_19569,N_17303,N_15933);
and U19570 (N_19570,N_16798,N_15782);
nand U19571 (N_19571,N_16466,N_15339);
and U19572 (N_19572,N_16368,N_16638);
nand U19573 (N_19573,N_17483,N_15919);
xnor U19574 (N_19574,N_15174,N_15437);
nor U19575 (N_19575,N_15574,N_15378);
nand U19576 (N_19576,N_16630,N_15983);
or U19577 (N_19577,N_15557,N_17316);
nor U19578 (N_19578,N_16777,N_15320);
nor U19579 (N_19579,N_15539,N_16720);
nor U19580 (N_19580,N_15130,N_16341);
and U19581 (N_19581,N_17023,N_15960);
or U19582 (N_19582,N_17332,N_16129);
and U19583 (N_19583,N_15888,N_16627);
nor U19584 (N_19584,N_17422,N_17498);
and U19585 (N_19585,N_16093,N_16803);
nor U19586 (N_19586,N_16774,N_15035);
xnor U19587 (N_19587,N_15683,N_15505);
xnor U19588 (N_19588,N_15567,N_16524);
or U19589 (N_19589,N_16019,N_15531);
xnor U19590 (N_19590,N_17167,N_15974);
nor U19591 (N_19591,N_15280,N_17025);
nand U19592 (N_19592,N_16661,N_16287);
or U19593 (N_19593,N_17350,N_16740);
or U19594 (N_19594,N_15034,N_17389);
and U19595 (N_19595,N_15930,N_16013);
nand U19596 (N_19596,N_16629,N_15301);
nand U19597 (N_19597,N_15756,N_16241);
or U19598 (N_19598,N_15291,N_15204);
nand U19599 (N_19599,N_17131,N_16858);
or U19600 (N_19600,N_16708,N_16408);
nor U19601 (N_19601,N_15591,N_16782);
xnor U19602 (N_19602,N_15409,N_16259);
nand U19603 (N_19603,N_15867,N_16219);
or U19604 (N_19604,N_17331,N_15538);
or U19605 (N_19605,N_16256,N_15371);
nand U19606 (N_19606,N_17393,N_15638);
xor U19607 (N_19607,N_15351,N_16714);
nor U19608 (N_19608,N_15027,N_16478);
and U19609 (N_19609,N_16840,N_15396);
nor U19610 (N_19610,N_15116,N_16064);
nand U19611 (N_19611,N_15880,N_15779);
and U19612 (N_19612,N_16250,N_15131);
nor U19613 (N_19613,N_16648,N_15872);
nor U19614 (N_19614,N_16382,N_16312);
nand U19615 (N_19615,N_15242,N_15391);
and U19616 (N_19616,N_16093,N_16665);
and U19617 (N_19617,N_15816,N_16639);
nor U19618 (N_19618,N_15525,N_15187);
nand U19619 (N_19619,N_16265,N_16254);
nand U19620 (N_19620,N_15243,N_16733);
nand U19621 (N_19621,N_16174,N_16352);
and U19622 (N_19622,N_16026,N_15477);
xnor U19623 (N_19623,N_16176,N_15113);
and U19624 (N_19624,N_15911,N_15336);
xnor U19625 (N_19625,N_16528,N_16918);
xnor U19626 (N_19626,N_15204,N_15974);
or U19627 (N_19627,N_15707,N_15294);
nor U19628 (N_19628,N_15507,N_16836);
and U19629 (N_19629,N_15415,N_15203);
and U19630 (N_19630,N_15348,N_15616);
and U19631 (N_19631,N_15619,N_17391);
nand U19632 (N_19632,N_16830,N_15853);
or U19633 (N_19633,N_16411,N_15591);
nor U19634 (N_19634,N_17149,N_16456);
nor U19635 (N_19635,N_17225,N_16277);
nor U19636 (N_19636,N_16844,N_17309);
nor U19637 (N_19637,N_16052,N_15652);
or U19638 (N_19638,N_15063,N_15274);
xnor U19639 (N_19639,N_16969,N_17380);
or U19640 (N_19640,N_15044,N_16821);
and U19641 (N_19641,N_16790,N_16924);
xnor U19642 (N_19642,N_15026,N_15794);
nor U19643 (N_19643,N_17274,N_16978);
xnor U19644 (N_19644,N_15896,N_15466);
or U19645 (N_19645,N_17384,N_15892);
xnor U19646 (N_19646,N_16028,N_16886);
nor U19647 (N_19647,N_16304,N_16644);
xnor U19648 (N_19648,N_16243,N_16606);
nor U19649 (N_19649,N_15700,N_15366);
and U19650 (N_19650,N_16305,N_16813);
xnor U19651 (N_19651,N_17234,N_15154);
nor U19652 (N_19652,N_16216,N_15021);
xor U19653 (N_19653,N_16453,N_16673);
nand U19654 (N_19654,N_15829,N_16426);
nand U19655 (N_19655,N_17008,N_15055);
nor U19656 (N_19656,N_15392,N_15423);
and U19657 (N_19657,N_17079,N_15406);
nor U19658 (N_19658,N_16563,N_16208);
or U19659 (N_19659,N_16746,N_15680);
xor U19660 (N_19660,N_16417,N_16552);
xnor U19661 (N_19661,N_15798,N_16663);
or U19662 (N_19662,N_15576,N_16120);
xor U19663 (N_19663,N_15213,N_17289);
nand U19664 (N_19664,N_17104,N_16808);
nand U19665 (N_19665,N_15809,N_15324);
nor U19666 (N_19666,N_16950,N_15121);
nand U19667 (N_19667,N_16955,N_16192);
xnor U19668 (N_19668,N_15438,N_15824);
nand U19669 (N_19669,N_15800,N_16375);
nand U19670 (N_19670,N_15868,N_17316);
nor U19671 (N_19671,N_15833,N_17177);
xor U19672 (N_19672,N_17424,N_15882);
xnor U19673 (N_19673,N_17300,N_16183);
and U19674 (N_19674,N_16278,N_16407);
nor U19675 (N_19675,N_15934,N_17314);
or U19676 (N_19676,N_15969,N_17171);
or U19677 (N_19677,N_17448,N_16925);
xnor U19678 (N_19678,N_17211,N_16455);
xor U19679 (N_19679,N_15654,N_16426);
nor U19680 (N_19680,N_17355,N_16281);
xnor U19681 (N_19681,N_16290,N_16060);
nor U19682 (N_19682,N_15165,N_17339);
nor U19683 (N_19683,N_16586,N_15081);
and U19684 (N_19684,N_16586,N_16662);
or U19685 (N_19685,N_15270,N_15048);
nor U19686 (N_19686,N_15354,N_17248);
and U19687 (N_19687,N_15583,N_15163);
and U19688 (N_19688,N_15106,N_16860);
nand U19689 (N_19689,N_17447,N_15015);
xor U19690 (N_19690,N_15326,N_16950);
nor U19691 (N_19691,N_16985,N_15110);
nor U19692 (N_19692,N_17378,N_15905);
and U19693 (N_19693,N_16534,N_17194);
nor U19694 (N_19694,N_16302,N_15210);
and U19695 (N_19695,N_16680,N_15633);
and U19696 (N_19696,N_16875,N_15557);
nor U19697 (N_19697,N_16208,N_15994);
and U19698 (N_19698,N_16447,N_16528);
and U19699 (N_19699,N_15341,N_16557);
and U19700 (N_19700,N_16639,N_17428);
nor U19701 (N_19701,N_15838,N_16733);
xnor U19702 (N_19702,N_16748,N_15021);
xor U19703 (N_19703,N_17212,N_17204);
or U19704 (N_19704,N_16394,N_16178);
and U19705 (N_19705,N_16164,N_15297);
or U19706 (N_19706,N_17157,N_16914);
xnor U19707 (N_19707,N_17247,N_15008);
or U19708 (N_19708,N_15019,N_16592);
and U19709 (N_19709,N_16822,N_17315);
or U19710 (N_19710,N_15815,N_15573);
or U19711 (N_19711,N_17416,N_16099);
xor U19712 (N_19712,N_15980,N_16801);
and U19713 (N_19713,N_15740,N_16627);
nand U19714 (N_19714,N_16463,N_15901);
nand U19715 (N_19715,N_15331,N_17104);
nor U19716 (N_19716,N_16435,N_15722);
nand U19717 (N_19717,N_16832,N_17162);
xor U19718 (N_19718,N_16566,N_15618);
xnor U19719 (N_19719,N_16012,N_16112);
or U19720 (N_19720,N_17090,N_17148);
xnor U19721 (N_19721,N_17195,N_15112);
or U19722 (N_19722,N_15095,N_15499);
or U19723 (N_19723,N_15279,N_15408);
nand U19724 (N_19724,N_17486,N_17188);
nor U19725 (N_19725,N_15667,N_16284);
nor U19726 (N_19726,N_17195,N_16799);
or U19727 (N_19727,N_15188,N_15586);
nand U19728 (N_19728,N_15508,N_16543);
nand U19729 (N_19729,N_16064,N_15684);
xnor U19730 (N_19730,N_15094,N_17340);
nor U19731 (N_19731,N_16772,N_17271);
nand U19732 (N_19732,N_16538,N_16877);
nor U19733 (N_19733,N_17065,N_16534);
nor U19734 (N_19734,N_17410,N_15484);
nor U19735 (N_19735,N_17338,N_15722);
and U19736 (N_19736,N_15758,N_16896);
nand U19737 (N_19737,N_17007,N_15861);
and U19738 (N_19738,N_15573,N_16339);
or U19739 (N_19739,N_16637,N_16431);
nand U19740 (N_19740,N_15028,N_15006);
and U19741 (N_19741,N_16471,N_16704);
nand U19742 (N_19742,N_16043,N_15709);
xor U19743 (N_19743,N_16194,N_15969);
xor U19744 (N_19744,N_17257,N_16233);
xor U19745 (N_19745,N_17454,N_16586);
xnor U19746 (N_19746,N_15385,N_16905);
and U19747 (N_19747,N_16363,N_17143);
xor U19748 (N_19748,N_16206,N_17014);
and U19749 (N_19749,N_15201,N_15735);
or U19750 (N_19750,N_15363,N_16378);
nor U19751 (N_19751,N_17150,N_16865);
and U19752 (N_19752,N_15695,N_16404);
nand U19753 (N_19753,N_17270,N_16150);
nor U19754 (N_19754,N_15270,N_16125);
nand U19755 (N_19755,N_16516,N_16905);
and U19756 (N_19756,N_15722,N_17170);
nand U19757 (N_19757,N_17465,N_16811);
xor U19758 (N_19758,N_17400,N_15930);
nand U19759 (N_19759,N_15954,N_16328);
nand U19760 (N_19760,N_15120,N_15999);
nor U19761 (N_19761,N_15391,N_17394);
nand U19762 (N_19762,N_16694,N_15378);
xnor U19763 (N_19763,N_16546,N_17231);
or U19764 (N_19764,N_16823,N_15163);
nand U19765 (N_19765,N_17435,N_16115);
nor U19766 (N_19766,N_15369,N_16936);
xnor U19767 (N_19767,N_15827,N_16062);
nor U19768 (N_19768,N_16212,N_15413);
and U19769 (N_19769,N_16305,N_15731);
nand U19770 (N_19770,N_16848,N_17106);
and U19771 (N_19771,N_15414,N_16168);
nand U19772 (N_19772,N_17365,N_16413);
xnor U19773 (N_19773,N_15820,N_15255);
xor U19774 (N_19774,N_16942,N_15263);
or U19775 (N_19775,N_17460,N_16063);
nor U19776 (N_19776,N_15492,N_17080);
nand U19777 (N_19777,N_15620,N_17474);
xor U19778 (N_19778,N_15814,N_15916);
xor U19779 (N_19779,N_16954,N_15121);
nor U19780 (N_19780,N_15425,N_15575);
nor U19781 (N_19781,N_15089,N_15813);
and U19782 (N_19782,N_16015,N_17247);
or U19783 (N_19783,N_17079,N_16683);
or U19784 (N_19784,N_16828,N_16466);
xor U19785 (N_19785,N_16485,N_17224);
and U19786 (N_19786,N_15340,N_15580);
or U19787 (N_19787,N_17278,N_17172);
and U19788 (N_19788,N_15207,N_15149);
and U19789 (N_19789,N_15105,N_17470);
or U19790 (N_19790,N_15214,N_15652);
or U19791 (N_19791,N_15492,N_15247);
xnor U19792 (N_19792,N_16528,N_17405);
nand U19793 (N_19793,N_16051,N_17376);
or U19794 (N_19794,N_15942,N_15304);
and U19795 (N_19795,N_15226,N_16570);
or U19796 (N_19796,N_16807,N_15709);
xnor U19797 (N_19797,N_17114,N_16221);
or U19798 (N_19798,N_15123,N_16784);
and U19799 (N_19799,N_17285,N_16917);
nand U19800 (N_19800,N_15336,N_16275);
xor U19801 (N_19801,N_15186,N_17412);
xnor U19802 (N_19802,N_16807,N_15293);
nor U19803 (N_19803,N_15234,N_16269);
xor U19804 (N_19804,N_17438,N_16377);
nor U19805 (N_19805,N_17151,N_17004);
nand U19806 (N_19806,N_16466,N_15923);
nor U19807 (N_19807,N_16832,N_16422);
nand U19808 (N_19808,N_16655,N_16523);
nor U19809 (N_19809,N_15991,N_15966);
and U19810 (N_19810,N_16631,N_17418);
and U19811 (N_19811,N_15468,N_15040);
nor U19812 (N_19812,N_16715,N_15958);
xnor U19813 (N_19813,N_16482,N_17357);
xor U19814 (N_19814,N_16630,N_15308);
or U19815 (N_19815,N_16425,N_17003);
nand U19816 (N_19816,N_15346,N_15016);
nor U19817 (N_19817,N_15737,N_16800);
or U19818 (N_19818,N_16301,N_16498);
xnor U19819 (N_19819,N_16216,N_15914);
nor U19820 (N_19820,N_17317,N_15301);
xnor U19821 (N_19821,N_15422,N_17445);
xnor U19822 (N_19822,N_15841,N_16076);
nand U19823 (N_19823,N_16476,N_15734);
or U19824 (N_19824,N_17477,N_15753);
nor U19825 (N_19825,N_17351,N_17149);
or U19826 (N_19826,N_17253,N_17282);
nor U19827 (N_19827,N_15537,N_15580);
nor U19828 (N_19828,N_16511,N_15470);
or U19829 (N_19829,N_16515,N_15734);
and U19830 (N_19830,N_16145,N_15570);
nand U19831 (N_19831,N_17211,N_15060);
and U19832 (N_19832,N_16194,N_16949);
or U19833 (N_19833,N_17388,N_16557);
or U19834 (N_19834,N_16732,N_17123);
xor U19835 (N_19835,N_16508,N_15878);
xnor U19836 (N_19836,N_17220,N_15446);
xor U19837 (N_19837,N_16914,N_16783);
or U19838 (N_19838,N_17424,N_15040);
and U19839 (N_19839,N_15654,N_17303);
nor U19840 (N_19840,N_17220,N_17306);
nand U19841 (N_19841,N_15838,N_15622);
or U19842 (N_19842,N_15579,N_15598);
and U19843 (N_19843,N_17114,N_17091);
nand U19844 (N_19844,N_17122,N_16826);
nand U19845 (N_19845,N_16591,N_16777);
xnor U19846 (N_19846,N_17268,N_16071);
or U19847 (N_19847,N_17356,N_16356);
nand U19848 (N_19848,N_17062,N_16013);
and U19849 (N_19849,N_17151,N_16717);
and U19850 (N_19850,N_15388,N_16981);
and U19851 (N_19851,N_16834,N_16746);
and U19852 (N_19852,N_15072,N_16842);
and U19853 (N_19853,N_15157,N_16430);
xnor U19854 (N_19854,N_15956,N_16924);
xnor U19855 (N_19855,N_17015,N_17278);
nor U19856 (N_19856,N_17146,N_17088);
nor U19857 (N_19857,N_15501,N_15303);
nand U19858 (N_19858,N_17421,N_16860);
xor U19859 (N_19859,N_16795,N_16101);
nor U19860 (N_19860,N_17092,N_15446);
xnor U19861 (N_19861,N_16112,N_15727);
or U19862 (N_19862,N_17212,N_15491);
nand U19863 (N_19863,N_15680,N_17040);
nand U19864 (N_19864,N_16279,N_16669);
or U19865 (N_19865,N_17192,N_17278);
nor U19866 (N_19866,N_17059,N_15865);
nand U19867 (N_19867,N_15854,N_17107);
nand U19868 (N_19868,N_15280,N_15373);
xnor U19869 (N_19869,N_15396,N_16319);
xor U19870 (N_19870,N_15701,N_16187);
nor U19871 (N_19871,N_15178,N_16104);
nor U19872 (N_19872,N_15848,N_17433);
or U19873 (N_19873,N_16319,N_15809);
nor U19874 (N_19874,N_15198,N_17398);
and U19875 (N_19875,N_16438,N_15484);
or U19876 (N_19876,N_17395,N_17438);
nand U19877 (N_19877,N_16145,N_16157);
xnor U19878 (N_19878,N_16564,N_15786);
and U19879 (N_19879,N_15357,N_17364);
or U19880 (N_19880,N_17442,N_17451);
nand U19881 (N_19881,N_15597,N_16390);
xor U19882 (N_19882,N_16409,N_16233);
or U19883 (N_19883,N_17242,N_16182);
and U19884 (N_19884,N_17210,N_15606);
or U19885 (N_19885,N_17489,N_17292);
or U19886 (N_19886,N_16744,N_15328);
nor U19887 (N_19887,N_15336,N_16566);
xnor U19888 (N_19888,N_16383,N_16696);
nand U19889 (N_19889,N_16635,N_15216);
nor U19890 (N_19890,N_16436,N_17310);
nor U19891 (N_19891,N_16192,N_17047);
xnor U19892 (N_19892,N_16978,N_16456);
and U19893 (N_19893,N_17046,N_16852);
nand U19894 (N_19894,N_15831,N_17444);
nand U19895 (N_19895,N_15439,N_15479);
or U19896 (N_19896,N_16074,N_17123);
and U19897 (N_19897,N_15493,N_15397);
xor U19898 (N_19898,N_16651,N_17315);
xnor U19899 (N_19899,N_17179,N_16909);
nor U19900 (N_19900,N_15742,N_15744);
or U19901 (N_19901,N_16453,N_17155);
and U19902 (N_19902,N_16801,N_16642);
xnor U19903 (N_19903,N_15590,N_16989);
xnor U19904 (N_19904,N_16777,N_16087);
nand U19905 (N_19905,N_15076,N_15269);
or U19906 (N_19906,N_17256,N_15197);
nor U19907 (N_19907,N_16396,N_16369);
xor U19908 (N_19908,N_15454,N_16257);
nand U19909 (N_19909,N_15897,N_17267);
and U19910 (N_19910,N_16603,N_16856);
or U19911 (N_19911,N_15923,N_16877);
xor U19912 (N_19912,N_15371,N_16422);
nand U19913 (N_19913,N_15271,N_16104);
xor U19914 (N_19914,N_15450,N_15254);
nand U19915 (N_19915,N_16133,N_16999);
xor U19916 (N_19916,N_16048,N_15497);
nand U19917 (N_19917,N_16378,N_15806);
nor U19918 (N_19918,N_17240,N_15509);
nor U19919 (N_19919,N_16512,N_15104);
or U19920 (N_19920,N_15701,N_16586);
nand U19921 (N_19921,N_15194,N_16121);
nor U19922 (N_19922,N_15347,N_15640);
nor U19923 (N_19923,N_15734,N_16044);
nor U19924 (N_19924,N_17499,N_17109);
nand U19925 (N_19925,N_15376,N_16074);
and U19926 (N_19926,N_17361,N_17120);
and U19927 (N_19927,N_16823,N_16996);
nand U19928 (N_19928,N_15246,N_16879);
nor U19929 (N_19929,N_15317,N_17041);
nand U19930 (N_19930,N_15567,N_15357);
and U19931 (N_19931,N_17155,N_17445);
xor U19932 (N_19932,N_16406,N_16793);
and U19933 (N_19933,N_16706,N_16357);
and U19934 (N_19934,N_15869,N_15578);
nor U19935 (N_19935,N_16271,N_15084);
xnor U19936 (N_19936,N_17398,N_16611);
nand U19937 (N_19937,N_17163,N_17273);
nor U19938 (N_19938,N_17390,N_15458);
nor U19939 (N_19939,N_17185,N_15318);
nand U19940 (N_19940,N_17268,N_16273);
xor U19941 (N_19941,N_16409,N_15965);
nand U19942 (N_19942,N_17405,N_16462);
nor U19943 (N_19943,N_17087,N_15007);
or U19944 (N_19944,N_15460,N_16784);
nand U19945 (N_19945,N_16584,N_15092);
nor U19946 (N_19946,N_16621,N_16435);
or U19947 (N_19947,N_16014,N_15907);
nand U19948 (N_19948,N_15021,N_16102);
nand U19949 (N_19949,N_17461,N_15188);
or U19950 (N_19950,N_15139,N_16182);
and U19951 (N_19951,N_15344,N_16678);
and U19952 (N_19952,N_17345,N_16892);
nor U19953 (N_19953,N_15597,N_15207);
and U19954 (N_19954,N_15371,N_17320);
and U19955 (N_19955,N_17089,N_15353);
nor U19956 (N_19956,N_16657,N_16333);
and U19957 (N_19957,N_15646,N_16843);
and U19958 (N_19958,N_15063,N_17378);
xnor U19959 (N_19959,N_15884,N_17345);
xor U19960 (N_19960,N_15790,N_15365);
xnor U19961 (N_19961,N_15111,N_15631);
nor U19962 (N_19962,N_17336,N_15653);
xnor U19963 (N_19963,N_15700,N_16585);
xnor U19964 (N_19964,N_17231,N_15030);
and U19965 (N_19965,N_15500,N_15614);
xor U19966 (N_19966,N_17187,N_15892);
or U19967 (N_19967,N_16284,N_15024);
or U19968 (N_19968,N_16780,N_15041);
and U19969 (N_19969,N_16644,N_16611);
xnor U19970 (N_19970,N_15020,N_16338);
or U19971 (N_19971,N_16998,N_16371);
or U19972 (N_19972,N_17032,N_16351);
xnor U19973 (N_19973,N_15192,N_17334);
or U19974 (N_19974,N_16291,N_16797);
xor U19975 (N_19975,N_15874,N_15116);
or U19976 (N_19976,N_15451,N_17018);
nor U19977 (N_19977,N_15260,N_17220);
or U19978 (N_19978,N_15636,N_15744);
xnor U19979 (N_19979,N_15266,N_15056);
nand U19980 (N_19980,N_15612,N_16985);
nor U19981 (N_19981,N_15506,N_16056);
and U19982 (N_19982,N_15729,N_16593);
xnor U19983 (N_19983,N_15003,N_15697);
nor U19984 (N_19984,N_16474,N_15798);
nand U19985 (N_19985,N_16952,N_15890);
and U19986 (N_19986,N_16574,N_15516);
or U19987 (N_19987,N_15680,N_16610);
or U19988 (N_19988,N_15435,N_16746);
and U19989 (N_19989,N_16913,N_16340);
and U19990 (N_19990,N_16686,N_17342);
xnor U19991 (N_19991,N_16493,N_16805);
or U19992 (N_19992,N_15144,N_15553);
or U19993 (N_19993,N_17031,N_15463);
xor U19994 (N_19994,N_16213,N_16393);
nor U19995 (N_19995,N_15015,N_16786);
and U19996 (N_19996,N_15555,N_16974);
and U19997 (N_19997,N_15737,N_17319);
nand U19998 (N_19998,N_16840,N_17207);
or U19999 (N_19999,N_16833,N_16887);
nand U20000 (N_20000,N_19931,N_18315);
or U20001 (N_20001,N_18945,N_18383);
or U20002 (N_20002,N_19123,N_18434);
xnor U20003 (N_20003,N_18177,N_19371);
or U20004 (N_20004,N_19088,N_19994);
nand U20005 (N_20005,N_18998,N_18281);
nand U20006 (N_20006,N_19814,N_19630);
or U20007 (N_20007,N_18296,N_19922);
or U20008 (N_20008,N_17632,N_19685);
nor U20009 (N_20009,N_18543,N_19803);
nand U20010 (N_20010,N_19660,N_19810);
or U20011 (N_20011,N_19645,N_19061);
and U20012 (N_20012,N_18994,N_19380);
and U20013 (N_20013,N_17701,N_18508);
nor U20014 (N_20014,N_19305,N_18507);
and U20015 (N_20015,N_18178,N_19087);
or U20016 (N_20016,N_19782,N_18195);
nand U20017 (N_20017,N_17862,N_18148);
nand U20018 (N_20018,N_18848,N_18878);
nand U20019 (N_20019,N_18786,N_17526);
and U20020 (N_20020,N_19520,N_18966);
xnor U20021 (N_20021,N_19290,N_19640);
xnor U20022 (N_20022,N_17569,N_18175);
or U20023 (N_20023,N_18387,N_17510);
or U20024 (N_20024,N_19908,N_17521);
nand U20025 (N_20025,N_17853,N_19979);
nor U20026 (N_20026,N_19151,N_18759);
xnor U20027 (N_20027,N_19581,N_19323);
xor U20028 (N_20028,N_18411,N_18872);
or U20029 (N_20029,N_18502,N_17574);
or U20030 (N_20030,N_17855,N_17969);
xnor U20031 (N_20031,N_19796,N_19511);
nor U20032 (N_20032,N_18644,N_18634);
nor U20033 (N_20033,N_19066,N_19069);
nand U20034 (N_20034,N_19666,N_18052);
nand U20035 (N_20035,N_19418,N_17509);
nor U20036 (N_20036,N_18865,N_19538);
nor U20037 (N_20037,N_18400,N_19473);
or U20038 (N_20038,N_17629,N_17646);
nand U20039 (N_20039,N_17590,N_18039);
xnor U20040 (N_20040,N_19754,N_17929);
nand U20041 (N_20041,N_19844,N_18883);
nand U20042 (N_20042,N_18196,N_18627);
nand U20043 (N_20043,N_18580,N_19582);
and U20044 (N_20044,N_18896,N_19318);
xnor U20045 (N_20045,N_18763,N_17888);
nor U20046 (N_20046,N_19986,N_19189);
xor U20047 (N_20047,N_18111,N_17966);
and U20048 (N_20048,N_17762,N_17717);
nand U20049 (N_20049,N_18163,N_17640);
and U20050 (N_20050,N_19121,N_18203);
and U20051 (N_20051,N_18625,N_18379);
nand U20052 (N_20052,N_17925,N_18618);
or U20053 (N_20053,N_18446,N_19554);
and U20054 (N_20054,N_18536,N_19054);
and U20055 (N_20055,N_18362,N_19800);
and U20056 (N_20056,N_17690,N_17752);
and U20057 (N_20057,N_17778,N_19542);
nand U20058 (N_20058,N_19879,N_19539);
xnor U20059 (N_20059,N_18079,N_18814);
and U20060 (N_20060,N_19045,N_18220);
nand U20061 (N_20061,N_17621,N_18898);
nand U20062 (N_20062,N_19638,N_18541);
nor U20063 (N_20063,N_19635,N_18230);
nor U20064 (N_20064,N_18675,N_18836);
xor U20065 (N_20065,N_19238,N_17910);
nor U20066 (N_20066,N_19606,N_19627);
nand U20067 (N_20067,N_18073,N_18742);
xor U20068 (N_20068,N_19185,N_18588);
nand U20069 (N_20069,N_19466,N_19383);
nor U20070 (N_20070,N_19722,N_18846);
nor U20071 (N_20071,N_17678,N_19624);
xor U20072 (N_20072,N_18932,N_18859);
nor U20073 (N_20073,N_19326,N_18605);
and U20074 (N_20074,N_18151,N_19234);
xor U20075 (N_20075,N_19029,N_17677);
xor U20076 (N_20076,N_17917,N_19372);
nor U20077 (N_20077,N_18194,N_18869);
and U20078 (N_20078,N_18173,N_19221);
nand U20079 (N_20079,N_19386,N_19619);
nand U20080 (N_20080,N_17829,N_18632);
xor U20081 (N_20081,N_17673,N_19019);
or U20082 (N_20082,N_17767,N_18258);
nand U20083 (N_20083,N_18150,N_19133);
nor U20084 (N_20084,N_17689,N_18562);
nand U20085 (N_20085,N_19052,N_18062);
or U20086 (N_20086,N_19737,N_17962);
and U20087 (N_20087,N_18843,N_18753);
and U20088 (N_20088,N_19250,N_18290);
nand U20089 (N_20089,N_17663,N_18187);
xnor U20090 (N_20090,N_17957,N_19615);
nor U20091 (N_20091,N_19552,N_18950);
nor U20092 (N_20092,N_19304,N_19701);
or U20093 (N_20093,N_19053,N_18352);
or U20094 (N_20094,N_19939,N_19598);
nor U20095 (N_20095,N_17786,N_19572);
nor U20096 (N_20096,N_19090,N_18262);
xor U20097 (N_20097,N_17770,N_18638);
and U20098 (N_20098,N_18834,N_18495);
and U20099 (N_20099,N_17926,N_19159);
nand U20100 (N_20100,N_19881,N_19595);
and U20101 (N_20101,N_18793,N_17593);
xnor U20102 (N_20102,N_19210,N_17906);
xnor U20103 (N_20103,N_19340,N_19845);
xnor U20104 (N_20104,N_19093,N_17980);
xor U20105 (N_20105,N_18467,N_19555);
nor U20106 (N_20106,N_18167,N_18086);
xor U20107 (N_20107,N_18068,N_17742);
or U20108 (N_20108,N_18589,N_18648);
xnor U20109 (N_20109,N_19370,N_17759);
and U20110 (N_20110,N_17603,N_18278);
xnor U20111 (N_20111,N_17530,N_18232);
xnor U20112 (N_20112,N_17923,N_19567);
nor U20113 (N_20113,N_19108,N_19794);
nor U20114 (N_20114,N_19760,N_19763);
nand U20115 (N_20115,N_19601,N_19523);
nand U20116 (N_20116,N_18797,N_18496);
and U20117 (N_20117,N_18683,N_17716);
xor U20118 (N_20118,N_17692,N_17628);
and U20119 (N_20119,N_18445,N_17810);
xnor U20120 (N_20120,N_17713,N_19809);
xor U20121 (N_20121,N_18942,N_19728);
or U20122 (N_20122,N_18581,N_19243);
nor U20123 (N_20123,N_17755,N_18420);
nor U20124 (N_20124,N_19182,N_18478);
or U20125 (N_20125,N_19378,N_18803);
xor U20126 (N_20126,N_18688,N_19697);
nand U20127 (N_20127,N_18840,N_18979);
nand U20128 (N_20128,N_19387,N_18593);
xnor U20129 (N_20129,N_19752,N_18585);
or U20130 (N_20130,N_18987,N_18715);
xnor U20131 (N_20131,N_18565,N_18812);
and U20132 (N_20132,N_19483,N_19876);
xnor U20133 (N_20133,N_17816,N_17706);
xnor U20134 (N_20134,N_18965,N_18686);
or U20135 (N_20135,N_19843,N_19482);
or U20136 (N_20136,N_17991,N_18545);
xor U20137 (N_20137,N_19808,N_19698);
nand U20138 (N_20138,N_18563,N_17736);
and U20139 (N_20139,N_17892,N_18300);
xor U20140 (N_20140,N_19507,N_17782);
or U20141 (N_20141,N_17757,N_19253);
xor U20142 (N_20142,N_18482,N_19330);
and U20143 (N_20143,N_17928,N_19262);
nor U20144 (N_20144,N_18768,N_18805);
nand U20145 (N_20145,N_18515,N_17914);
nor U20146 (N_20146,N_18264,N_18731);
nor U20147 (N_20147,N_18170,N_18384);
nor U20148 (N_20148,N_19166,N_18967);
and U20149 (N_20149,N_19526,N_19670);
and U20150 (N_20150,N_18432,N_18423);
xor U20151 (N_20151,N_17684,N_19625);
nor U20152 (N_20152,N_19109,N_19780);
nor U20153 (N_20153,N_19824,N_18917);
nor U20154 (N_20154,N_19144,N_17572);
xor U20155 (N_20155,N_18261,N_18568);
nand U20156 (N_20156,N_19079,N_18877);
xor U20157 (N_20157,N_17840,N_18540);
nand U20158 (N_20158,N_17769,N_17904);
xor U20159 (N_20159,N_17776,N_18210);
or U20160 (N_20160,N_19329,N_19214);
xnor U20161 (N_20161,N_19333,N_18548);
nor U20162 (N_20162,N_18146,N_19263);
or U20163 (N_20163,N_17505,N_19082);
and U20164 (N_20164,N_18200,N_17664);
nor U20165 (N_20165,N_19802,N_18693);
xnor U20166 (N_20166,N_19911,N_19923);
or U20167 (N_20167,N_18692,N_19279);
or U20168 (N_20168,N_19155,N_19909);
and U20169 (N_20169,N_19900,N_19904);
nand U20170 (N_20170,N_19682,N_17899);
nor U20171 (N_20171,N_19514,N_18864);
or U20172 (N_20172,N_18143,N_19195);
nand U20173 (N_20173,N_19621,N_19367);
nor U20174 (N_20174,N_18449,N_19832);
or U20175 (N_20175,N_18106,N_19616);
and U20176 (N_20176,N_19286,N_18820);
nor U20177 (N_20177,N_17723,N_18019);
or U20178 (N_20178,N_19608,N_17651);
nor U20179 (N_20179,N_17813,N_18041);
or U20180 (N_20180,N_17679,N_18240);
and U20181 (N_20181,N_18154,N_19834);
nand U20182 (N_20182,N_18123,N_19590);
nor U20183 (N_20183,N_18351,N_19348);
or U20184 (N_20184,N_18606,N_18839);
or U20185 (N_20185,N_19235,N_18389);
or U20186 (N_20186,N_17804,N_18852);
or U20187 (N_20187,N_19042,N_18008);
nand U20188 (N_20188,N_18375,N_18301);
or U20189 (N_20189,N_19969,N_18844);
nand U20190 (N_20190,N_18986,N_17841);
and U20191 (N_20191,N_18991,N_17595);
or U20192 (N_20192,N_17922,N_19264);
and U20193 (N_20193,N_19704,N_19711);
nand U20194 (N_20194,N_18224,N_18689);
nor U20195 (N_20195,N_17943,N_19256);
nand U20196 (N_20196,N_19030,N_18798);
nand U20197 (N_20197,N_18271,N_18357);
nor U20198 (N_20198,N_18408,N_17710);
and U20199 (N_20199,N_19416,N_17780);
and U20200 (N_20200,N_18747,N_18845);
and U20201 (N_20201,N_18458,N_17789);
nand U20202 (N_20202,N_19292,N_18102);
nor U20203 (N_20203,N_18671,N_19351);
nor U20204 (N_20204,N_17682,N_19425);
xnor U20205 (N_20205,N_19715,N_19246);
and U20206 (N_20206,N_19532,N_19398);
nor U20207 (N_20207,N_18457,N_18633);
nand U20208 (N_20208,N_17583,N_19048);
nand U20209 (N_20209,N_17758,N_19435);
or U20210 (N_20210,N_18160,N_17790);
or U20211 (N_20211,N_17798,N_19956);
or U20212 (N_20212,N_18342,N_18560);
nand U20213 (N_20213,N_19783,N_17787);
or U20214 (N_20214,N_18356,N_19314);
or U20215 (N_20215,N_19334,N_18863);
nand U20216 (N_20216,N_19219,N_19712);
nand U20217 (N_20217,N_18038,N_17581);
nor U20218 (N_20218,N_18573,N_17675);
nand U20219 (N_20219,N_18021,N_18456);
and U20220 (N_20220,N_17982,N_19460);
or U20221 (N_20221,N_18738,N_17792);
nand U20222 (N_20222,N_18968,N_18460);
and U20223 (N_20223,N_18779,N_17570);
and U20224 (N_20224,N_19709,N_17747);
nor U20225 (N_20225,N_18931,N_19434);
or U20226 (N_20226,N_18244,N_19603);
or U20227 (N_20227,N_19633,N_17618);
nor U20228 (N_20228,N_19374,N_18306);
and U20229 (N_20229,N_19324,N_18144);
or U20230 (N_20230,N_19623,N_19620);
and U20231 (N_20231,N_19441,N_18961);
and U20232 (N_20232,N_19352,N_19164);
nor U20233 (N_20233,N_18533,N_19410);
or U20234 (N_20234,N_19487,N_18586);
nand U20235 (N_20235,N_18801,N_18601);
nor U20236 (N_20236,N_18815,N_18736);
nand U20237 (N_20237,N_18854,N_17584);
and U20238 (N_20238,N_19767,N_18489);
nor U20239 (N_20239,N_19945,N_19848);
and U20240 (N_20240,N_18103,N_17774);
or U20241 (N_20241,N_19871,N_18661);
or U20242 (N_20242,N_18596,N_17815);
and U20243 (N_20243,N_19423,N_18191);
nand U20244 (N_20244,N_17513,N_17911);
nand U20245 (N_20245,N_17616,N_18369);
and U20246 (N_20246,N_17860,N_19774);
or U20247 (N_20247,N_17874,N_18600);
nand U20248 (N_20248,N_19570,N_18424);
xnor U20249 (N_20249,N_18436,N_17764);
nand U20250 (N_20250,N_17585,N_18226);
nand U20251 (N_20251,N_18184,N_18771);
and U20252 (N_20252,N_17726,N_19886);
and U20253 (N_20253,N_18270,N_19591);
nand U20254 (N_20254,N_19963,N_19322);
xnor U20255 (N_20255,N_17958,N_19805);
xor U20256 (N_20256,N_17611,N_19628);
and U20257 (N_20257,N_18181,N_19707);
nor U20258 (N_20258,N_17732,N_18235);
or U20259 (N_20259,N_19202,N_17838);
or U20260 (N_20260,N_18055,N_19756);
and U20261 (N_20261,N_19449,N_19953);
nor U20262 (N_20262,N_17858,N_19962);
xnor U20263 (N_20263,N_17896,N_19091);
xnor U20264 (N_20264,N_18437,N_19336);
nor U20265 (N_20265,N_17971,N_18622);
nor U20266 (N_20266,N_18652,N_19533);
xnor U20267 (N_20267,N_18269,N_17658);
and U20268 (N_20268,N_19585,N_18959);
and U20269 (N_20269,N_19446,N_19359);
xor U20270 (N_20270,N_19674,N_19335);
nand U20271 (N_20271,N_17734,N_19864);
or U20272 (N_20272,N_17970,N_17979);
or U20273 (N_20273,N_18398,N_18957);
nor U20274 (N_20274,N_18288,N_19557);
nor U20275 (N_20275,N_18631,N_19519);
nor U20276 (N_20276,N_18327,N_19749);
nor U20277 (N_20277,N_19165,N_18695);
nor U20278 (N_20278,N_18755,N_19872);
and U20279 (N_20279,N_19394,N_19018);
nand U20280 (N_20280,N_19566,N_18741);
and U20281 (N_20281,N_19642,N_18569);
xnor U20282 (N_20282,N_18292,N_18049);
or U20283 (N_20283,N_19181,N_17671);
nand U20284 (N_20284,N_18228,N_17844);
xnor U20285 (N_20285,N_17848,N_18913);
or U20286 (N_20286,N_19480,N_19580);
nand U20287 (N_20287,N_18721,N_19127);
nor U20288 (N_20288,N_18701,N_19869);
or U20289 (N_20289,N_17919,N_18131);
and U20290 (N_20290,N_18691,N_18268);
and U20291 (N_20291,N_18906,N_18874);
nand U20292 (N_20292,N_17882,N_19431);
and U20293 (N_20293,N_19356,N_19804);
nor U20294 (N_20294,N_17791,N_19186);
nor U20295 (N_20295,N_17733,N_18685);
nor U20296 (N_20296,N_19654,N_18500);
or U20297 (N_20297,N_18992,N_18591);
or U20298 (N_20298,N_17502,N_18713);
xor U20299 (N_20299,N_18129,N_19569);
nand U20300 (N_20300,N_19500,N_19791);
or U20301 (N_20301,N_19610,N_18700);
nor U20302 (N_20302,N_18649,N_19150);
and U20303 (N_20303,N_19980,N_18428);
nand U20304 (N_20304,N_19039,N_17533);
nor U20305 (N_20305,N_17903,N_18023);
nand U20306 (N_20306,N_17676,N_19820);
or U20307 (N_20307,N_19565,N_19187);
nor U20308 (N_20308,N_18450,N_18005);
nor U20309 (N_20309,N_18544,N_19114);
xor U20310 (N_20310,N_19462,N_18476);
or U20311 (N_20311,N_18503,N_19295);
nand U20312 (N_20312,N_19056,N_18418);
nand U20313 (N_20313,N_17609,N_18182);
and U20314 (N_20314,N_18359,N_19901);
and U20315 (N_20315,N_17699,N_17540);
nor U20316 (N_20316,N_19947,N_17607);
and U20317 (N_20317,N_18043,N_18046);
nand U20318 (N_20318,N_18510,N_18413);
nand U20319 (N_20319,N_18838,N_17639);
nand U20320 (N_20320,N_19225,N_17525);
xnor U20321 (N_20321,N_17784,N_18733);
or U20322 (N_20322,N_18130,N_17516);
or U20323 (N_20323,N_18037,N_19490);
and U20324 (N_20324,N_19167,N_18025);
xnor U20325 (N_20325,N_18263,N_19240);
and U20326 (N_20326,N_18169,N_18522);
or U20327 (N_20327,N_17743,N_18980);
xor U20328 (N_20328,N_19694,N_17897);
nand U20329 (N_20329,N_18385,N_19111);
nand U20330 (N_20330,N_18241,N_19083);
nor U20331 (N_20331,N_19512,N_19583);
nand U20332 (N_20332,N_19267,N_19197);
and U20333 (N_20333,N_18925,N_18058);
nor U20334 (N_20334,N_17977,N_18788);
nand U20335 (N_20335,N_19695,N_19223);
nor U20336 (N_20336,N_18745,N_17956);
or U20337 (N_20337,N_17907,N_19850);
or U20338 (N_20338,N_18860,N_19437);
or U20339 (N_20339,N_19903,N_19812);
nand U20340 (N_20340,N_18928,N_18222);
xor U20341 (N_20341,N_18164,N_19815);
xnor U20342 (N_20342,N_18882,N_18772);
or U20343 (N_20343,N_19837,N_17865);
or U20344 (N_20344,N_19556,N_19938);
nand U20345 (N_20345,N_19145,N_17863);
or U20346 (N_20346,N_19935,N_17833);
or U20347 (N_20347,N_17936,N_18572);
xnor U20348 (N_20348,N_18653,N_18523);
and U20349 (N_20349,N_19564,N_18498);
nor U20350 (N_20350,N_19541,N_18211);
nor U20351 (N_20351,N_18372,N_18789);
or U20352 (N_20352,N_18497,N_19893);
nor U20353 (N_20353,N_19152,N_19020);
nand U20354 (N_20354,N_17763,N_17557);
xnor U20355 (N_20355,N_19173,N_19641);
xor U20356 (N_20356,N_19128,N_18934);
or U20357 (N_20357,N_18590,N_19578);
or U20358 (N_20358,N_19971,N_18016);
or U20359 (N_20359,N_18166,N_18775);
nand U20360 (N_20360,N_18579,N_18604);
or U20361 (N_20361,N_18333,N_19308);
nand U20362 (N_20362,N_18748,N_18406);
nand U20363 (N_20363,N_19313,N_19721);
or U20364 (N_20364,N_19933,N_18595);
or U20365 (N_20365,N_19468,N_18371);
nor U20366 (N_20366,N_19459,N_18930);
nor U20367 (N_20367,N_19735,N_17795);
xnor U20368 (N_20368,N_18673,N_17587);
and U20369 (N_20369,N_19798,N_19561);
xnor U20370 (N_20370,N_18116,N_19686);
xnor U20371 (N_20371,N_19992,N_17870);
or U20372 (N_20372,N_18702,N_18804);
and U20373 (N_20373,N_18433,N_17598);
or U20374 (N_20374,N_18421,N_17927);
nand U20375 (N_20375,N_18556,N_18935);
and U20376 (N_20376,N_18105,N_18088);
nand U20377 (N_20377,N_19261,N_18219);
nor U20378 (N_20378,N_17683,N_17672);
nor U20379 (N_20379,N_18238,N_18547);
and U20380 (N_20380,N_19426,N_18993);
nand U20381 (N_20381,N_18245,N_17731);
xnor U20382 (N_20382,N_19631,N_19439);
nand U20383 (N_20383,N_19675,N_19353);
nor U20384 (N_20384,N_18282,N_19696);
nor U20385 (N_20385,N_17568,N_18125);
or U20386 (N_20386,N_17845,N_18350);
or U20387 (N_20387,N_17626,N_19113);
nor U20388 (N_20388,N_18720,N_18750);
nor U20389 (N_20389,N_17947,N_18443);
nor U20390 (N_20390,N_17712,N_19594);
or U20391 (N_20391,N_18363,N_18637);
or U20392 (N_20392,N_17992,N_19649);
or U20393 (N_20393,N_19216,N_17781);
and U20394 (N_20394,N_19702,N_19276);
or U20395 (N_20395,N_17963,N_18977);
and U20396 (N_20396,N_18776,N_19772);
and U20397 (N_20397,N_18287,N_18322);
nand U20398 (N_20398,N_18650,N_19427);
and U20399 (N_20399,N_18310,N_19447);
and U20400 (N_20400,N_19075,N_18842);
xnor U20401 (N_20401,N_19852,N_18465);
or U20402 (N_20402,N_18297,N_19201);
nand U20403 (N_20403,N_19043,N_18463);
nor U20404 (N_20404,N_18654,N_19742);
and U20405 (N_20405,N_18903,N_17631);
nand U20406 (N_20406,N_17974,N_18990);
nor U20407 (N_20407,N_19117,N_18910);
nand U20408 (N_20408,N_17768,N_19160);
or U20409 (N_20409,N_19531,N_19245);
nand U20410 (N_20410,N_19260,N_18795);
nand U20411 (N_20411,N_19445,N_18126);
and U20412 (N_20412,N_18345,N_18147);
nand U20413 (N_20413,N_19716,N_18811);
nor U20414 (N_20414,N_18045,N_17512);
xor U20415 (N_20415,N_19786,N_17552);
xnor U20416 (N_20416,N_17535,N_18555);
xor U20417 (N_20417,N_18137,N_18893);
and U20418 (N_20418,N_19759,N_18902);
or U20419 (N_20419,N_19285,N_19825);
xnor U20420 (N_20420,N_18762,N_19576);
and U20421 (N_20421,N_18321,N_18636);
nand U20422 (N_20422,N_19009,N_18933);
or U20423 (N_20423,N_19148,N_17951);
nand U20424 (N_20424,N_18484,N_19915);
nor U20425 (N_20425,N_19781,N_18353);
nand U20426 (N_20426,N_18997,N_19008);
xor U20427 (N_20427,N_18879,N_18900);
and U20428 (N_20428,N_18635,N_19954);
xnor U20429 (N_20429,N_17744,N_19016);
and U20430 (N_20430,N_17573,N_18093);
or U20431 (N_20431,N_19745,N_18373);
nor U20432 (N_20432,N_17740,N_17688);
and U20433 (N_20433,N_17884,N_17634);
xor U20434 (N_20434,N_17913,N_17534);
nand U20435 (N_20435,N_19443,N_19074);
nor U20436 (N_20436,N_17722,N_18461);
or U20437 (N_20437,N_18911,N_18355);
nand U20438 (N_20438,N_17704,N_18758);
nand U20439 (N_20439,N_19458,N_19743);
nand U20440 (N_20440,N_18361,N_19972);
and U20441 (N_20441,N_19919,N_19489);
xnor U20442 (N_20442,N_19878,N_19977);
nand U20443 (N_20443,N_17602,N_17670);
and U20444 (N_20444,N_17702,N_19254);
nor U20445 (N_20445,N_18391,N_17827);
nand U20446 (N_20446,N_18983,N_18723);
nor U20447 (N_20447,N_18623,N_17832);
nand U20448 (N_20448,N_17567,N_19936);
nand U20449 (N_20449,N_17807,N_18888);
or U20450 (N_20450,N_19924,N_18466);
nor U20451 (N_20451,N_19942,N_19492);
xor U20452 (N_20452,N_18076,N_17693);
nor U20453 (N_20453,N_19966,N_18018);
nor U20454 (N_20454,N_19033,N_18386);
nand U20455 (N_20455,N_19714,N_17964);
or U20456 (N_20456,N_19907,N_19663);
or U20457 (N_20457,N_18441,N_19921);
xor U20458 (N_20458,N_17965,N_19027);
xnor U20459 (N_20459,N_18003,N_18868);
and U20460 (N_20460,N_19239,N_19671);
xor U20461 (N_20461,N_18276,N_19653);
xnor U20462 (N_20462,N_18936,N_17949);
and U20463 (N_20463,N_19790,N_18559);
xnor U20464 (N_20464,N_18974,N_19588);
xor U20465 (N_20465,N_18584,N_19384);
nand U20466 (N_20466,N_17837,N_18087);
nor U20467 (N_20467,N_18853,N_17826);
and U20468 (N_20468,N_19047,N_18380);
and U20469 (N_20469,N_17617,N_18085);
nand U20470 (N_20470,N_17578,N_19661);
nand U20471 (N_20471,N_18481,N_18317);
nand U20472 (N_20472,N_18213,N_19092);
nor U20473 (N_20473,N_19917,N_18072);
or U20474 (N_20474,N_17566,N_17820);
xor U20475 (N_20475,N_19101,N_19301);
and U20476 (N_20476,N_19273,N_17739);
or U20477 (N_20477,N_17830,N_17746);
or U20478 (N_20478,N_19573,N_17539);
and U20479 (N_20479,N_19188,N_19983);
or U20480 (N_20480,N_17729,N_19762);
or U20481 (N_20481,N_19229,N_18651);
nand U20482 (N_20482,N_19455,N_17808);
nor U20483 (N_20483,N_18857,N_19130);
or U20484 (N_20484,N_18074,N_18740);
and U20485 (N_20485,N_19522,N_19502);
xor U20486 (N_20486,N_19788,N_17959);
nor U20487 (N_20487,N_19086,N_19255);
or U20488 (N_20488,N_17511,N_19668);
or U20489 (N_20489,N_18963,N_18153);
nor U20490 (N_20490,N_19821,N_19949);
and U20491 (N_20491,N_19094,N_19041);
xor U20492 (N_20492,N_18311,N_19894);
nand U20493 (N_20493,N_18065,N_18015);
and U20494 (N_20494,N_18599,N_19344);
or U20495 (N_20495,N_18819,N_18982);
or U20496 (N_20496,N_19097,N_19958);
nor U20497 (N_20497,N_17898,N_19571);
nand U20498 (N_20498,N_18698,N_18609);
nand U20499 (N_20499,N_18909,N_19456);
and U20500 (N_20500,N_18973,N_18304);
nand U20501 (N_20501,N_18658,N_17522);
nor U20502 (N_20502,N_18452,N_19310);
xnor U20503 (N_20503,N_18611,N_19428);
nand U20504 (N_20504,N_19354,N_17989);
nand U20505 (N_20505,N_19995,N_19289);
nand U20506 (N_20506,N_17633,N_17915);
and U20507 (N_20507,N_19863,N_19667);
nand U20508 (N_20508,N_18969,N_17749);
xnor U20509 (N_20509,N_17803,N_18782);
and U20510 (N_20510,N_19129,N_18094);
nand U20511 (N_20511,N_18010,N_18266);
or U20512 (N_20512,N_18340,N_18940);
xor U20513 (N_20513,N_19747,N_19122);
xnor U20514 (N_20514,N_17765,N_18112);
and U20515 (N_20515,N_18127,N_19477);
nor U20516 (N_20516,N_18817,N_19385);
nand U20517 (N_20517,N_19085,N_17500);
nor U20518 (N_20518,N_19366,N_18639);
or U20519 (N_20519,N_18620,N_18571);
and U20520 (N_20520,N_19143,N_19673);
nor U20521 (N_20521,N_18455,N_19614);
or U20522 (N_20522,N_17783,N_18628);
nor U20523 (N_20523,N_18118,N_18621);
and U20524 (N_20524,N_18430,N_17937);
nand U20525 (N_20525,N_19194,N_18551);
nand U20526 (N_20526,N_19103,N_17879);
and U20527 (N_20527,N_19251,N_19787);
nor U20528 (N_20528,N_17933,N_19448);
or U20529 (N_20529,N_17987,N_19228);
nor U20530 (N_20530,N_18295,N_18529);
nand U20531 (N_20531,N_19361,N_18115);
nor U20532 (N_20532,N_17591,N_18608);
nand U20533 (N_20533,N_18528,N_18764);
and U20534 (N_20534,N_19328,N_19540);
and U20535 (N_20535,N_17604,N_18862);
xnor U20536 (N_20536,N_19126,N_18946);
nor U20537 (N_20537,N_19764,N_19975);
nand U20538 (N_20538,N_18107,N_19730);
and U20539 (N_20539,N_18880,N_17842);
nor U20540 (N_20540,N_19134,N_18247);
xor U20541 (N_20541,N_19988,N_17894);
nor U20542 (N_20542,N_17501,N_18028);
or U20543 (N_20543,N_17681,N_19636);
nor U20544 (N_20544,N_17993,N_19132);
and U20545 (N_20545,N_17821,N_19600);
or U20546 (N_20546,N_19875,N_19461);
nand U20547 (N_20547,N_17846,N_18676);
or U20548 (N_20548,N_19637,N_19951);
xnor U20549 (N_20549,N_18236,N_18908);
xor U20550 (N_20550,N_18679,N_18855);
nor U20551 (N_20551,N_19925,N_18985);
nand U20552 (N_20552,N_17669,N_18922);
and U20553 (N_20553,N_18616,N_17532);
nand U20554 (N_20554,N_18303,N_18091);
and U20555 (N_20555,N_19952,N_18419);
and U20556 (N_20556,N_18557,N_18615);
or U20557 (N_20557,N_19746,N_19713);
and U20558 (N_20558,N_17944,N_19705);
nor U20559 (N_20559,N_19247,N_17835);
or U20560 (N_20560,N_18850,N_19968);
xor U20561 (N_20561,N_19605,N_19158);
and U20562 (N_20562,N_18491,N_19681);
nor U20563 (N_20563,N_19859,N_18607);
or U20564 (N_20564,N_18447,N_19177);
xnor U20565 (N_20565,N_19537,N_18141);
xor U20566 (N_20566,N_18947,N_17883);
and U20567 (N_20567,N_18337,N_19388);
and U20568 (N_20568,N_17547,N_18577);
nor U20569 (N_20569,N_18610,N_17748);
nand U20570 (N_20570,N_18442,N_19171);
xor U20571 (N_20571,N_19841,N_19017);
nand U20572 (N_20572,N_17779,N_18470);
and U20573 (N_20573,N_18078,N_18225);
xor U20574 (N_20574,N_18197,N_19536);
and U20575 (N_20575,N_19548,N_19277);
xnor U20576 (N_20576,N_19208,N_18064);
xnor U20577 (N_20577,N_17504,N_17869);
nand U20578 (N_20578,N_19300,N_18221);
and U20579 (N_20579,N_19773,N_18212);
or U20580 (N_20580,N_19232,N_18684);
nor U20581 (N_20581,N_19525,N_19319);
xor U20582 (N_20582,N_19718,N_19411);
and U20583 (N_20583,N_18365,N_18624);
or U20584 (N_20584,N_18472,N_17635);
nor U20585 (N_20585,N_19741,N_18155);
and U20586 (N_20586,N_18108,N_18822);
or U20587 (N_20587,N_19156,N_18494);
and U20588 (N_20588,N_17520,N_17794);
nand U20589 (N_20589,N_18867,N_19861);
and U20590 (N_20590,N_19626,N_19226);
xor U20591 (N_20591,N_19391,N_19770);
and U20592 (N_20592,N_18279,N_17895);
nand U20593 (N_20593,N_18554,N_19910);
xor U20594 (N_20594,N_19612,N_18719);
xnor U20595 (N_20595,N_17659,N_19846);
nand U20596 (N_20596,N_19178,N_17796);
or U20597 (N_20597,N_18206,N_18703);
nor U20598 (N_20598,N_17606,N_17686);
nor U20599 (N_20599,N_19175,N_19978);
xor U20600 (N_20600,N_17875,N_17559);
nand U20601 (N_20601,N_19248,N_18128);
xor U20602 (N_20602,N_19475,N_19998);
nand U20603 (N_20603,N_18179,N_17950);
xor U20604 (N_20604,N_18792,N_18527);
or U20605 (N_20605,N_17961,N_18320);
or U20606 (N_20606,N_17756,N_19397);
xor U20607 (N_20607,N_19724,N_18416);
and U20608 (N_20608,N_19689,N_19720);
nor U20609 (N_20609,N_17541,N_19288);
and U20610 (N_20610,N_18717,N_17600);
or U20611 (N_20611,N_19717,N_19390);
and U20612 (N_20612,N_17812,N_19098);
and U20613 (N_20613,N_17721,N_19149);
and U20614 (N_20614,N_17548,N_18981);
or U20615 (N_20615,N_18767,N_19882);
nor U20616 (N_20616,N_17657,N_19296);
xnor U20617 (N_20617,N_19826,N_18090);
nor U20618 (N_20618,N_17945,N_18399);
or U20619 (N_20619,N_19058,N_18783);
nor U20620 (N_20620,N_19454,N_19015);
or U20621 (N_20621,N_17814,N_19577);
xor U20622 (N_20622,N_18907,N_18735);
nor U20623 (N_20623,N_18574,N_19025);
nor U20624 (N_20624,N_17551,N_18561);
and U20625 (N_20625,N_19493,N_18414);
nand U20626 (N_20626,N_18827,N_18535);
and U20627 (N_20627,N_19740,N_17705);
nor U20628 (N_20628,N_17825,N_18316);
nor U20629 (N_20629,N_18035,N_17893);
nor U20630 (N_20630,N_18956,N_19479);
nor U20631 (N_20631,N_18674,N_19183);
or U20632 (N_20632,N_17999,N_19139);
nor U20633 (N_20633,N_18291,N_19609);
nand U20634 (N_20634,N_19659,N_17878);
and U20635 (N_20635,N_19700,N_19154);
or U20636 (N_20636,N_19190,N_19115);
or U20637 (N_20637,N_17564,N_18204);
xor U20638 (N_20638,N_18168,N_19014);
nor U20639 (N_20639,N_17901,N_18439);
nor U20640 (N_20640,N_19022,N_18952);
xnor U20641 (N_20641,N_17967,N_19639);
or U20642 (N_20642,N_19407,N_19867);
xnor U20643 (N_20643,N_19967,N_19586);
and U20644 (N_20644,N_19508,N_19282);
or U20645 (N_20645,N_19753,N_17891);
nand U20646 (N_20646,N_18280,N_18100);
nand U20647 (N_20647,N_19562,N_19829);
nand U20648 (N_20648,N_18697,N_19799);
xor U20649 (N_20649,N_17924,N_18328);
nor U20650 (N_20650,N_18395,N_17655);
nor U20651 (N_20651,N_19847,N_19708);
nor U20652 (N_20652,N_19849,N_19049);
or U20653 (N_20653,N_18978,N_19116);
nand U20654 (N_20654,N_17885,N_19157);
and U20655 (N_20655,N_19424,N_19272);
and U20656 (N_20656,N_18109,N_18749);
nand U20657 (N_20657,N_18215,N_18809);
xor U20658 (N_20658,N_18462,N_18646);
nand U20659 (N_20659,N_17868,N_18512);
and U20660 (N_20660,N_18031,N_18440);
nor U20661 (N_20661,N_19811,N_19692);
xor U20662 (N_20662,N_19222,N_19895);
and U20663 (N_20663,N_18308,N_19119);
nor U20664 (N_20664,N_18294,N_18670);
nor U20665 (N_20665,N_19930,N_19420);
and U20666 (N_20666,N_18504,N_19929);
xnor U20667 (N_20667,N_18254,N_19161);
nand U20668 (N_20668,N_19467,N_19193);
nor U20669 (N_20669,N_17942,N_19912);
or U20670 (N_20670,N_17694,N_18193);
or U20671 (N_20671,N_18256,N_18958);
or U20672 (N_20672,N_17691,N_17737);
nor U20673 (N_20673,N_18207,N_19104);
xnor U20674 (N_20674,N_19976,N_19777);
or U20675 (N_20675,N_18487,N_18598);
nand U20676 (N_20676,N_18286,N_19023);
nor U20677 (N_20677,N_17849,N_18013);
xor U20678 (N_20678,N_19751,N_18505);
or U20679 (N_20679,N_19916,N_19934);
or U20680 (N_20680,N_18253,N_17674);
xnor U20681 (N_20681,N_18403,N_19611);
nand U20682 (N_20682,N_19044,N_18343);
or U20683 (N_20683,N_18681,N_18951);
or U20684 (N_20684,N_17998,N_19024);
nand U20685 (N_20685,N_18760,N_18937);
or U20686 (N_20686,N_18302,N_19607);
or U20687 (N_20687,N_19937,N_18145);
nor U20688 (N_20688,N_18666,N_19430);
and U20689 (N_20689,N_19281,N_18884);
nand U20690 (N_20690,N_18050,N_19220);
and U20691 (N_20691,N_19497,N_18022);
xnor U20692 (N_20692,N_18870,N_18694);
or U20693 (N_20693,N_18597,N_18732);
nand U20694 (N_20694,N_19987,N_19031);
and U20695 (N_20695,N_18012,N_17800);
nand U20696 (N_20696,N_18643,N_19037);
and U20697 (N_20697,N_18218,N_18570);
nand U20698 (N_20698,N_18890,N_17529);
nor U20699 (N_20699,N_18095,N_18806);
or U20700 (N_20700,N_18431,N_17809);
nor U20701 (N_20701,N_19959,N_18664);
xor U20702 (N_20702,N_18077,N_19679);
nand U20703 (N_20703,N_19725,N_19034);
nor U20704 (N_20704,N_19191,N_17909);
or U20705 (N_20705,N_17641,N_18542);
or U20706 (N_20706,N_19550,N_19332);
and U20707 (N_20707,N_17985,N_19233);
and U20708 (N_20708,N_18825,N_18823);
nand U20709 (N_20709,N_17995,N_18017);
nand U20710 (N_20710,N_18323,N_18629);
nor U20711 (N_20711,N_18492,N_18260);
and U20712 (N_20712,N_19270,N_19833);
and U20713 (N_20713,N_19355,N_18641);
or U20714 (N_20714,N_18368,N_19868);
or U20715 (N_20715,N_19828,N_18927);
or U20716 (N_20716,N_18051,N_19236);
or U20717 (N_20717,N_19203,N_18708);
xnor U20718 (N_20718,N_18142,N_18335);
or U20719 (N_20719,N_19906,N_19312);
nand U20720 (N_20720,N_17720,N_18818);
xor U20721 (N_20721,N_18892,N_18097);
or U20722 (N_20722,N_17549,N_19485);
nor U20723 (N_20723,N_17905,N_17773);
nand U20724 (N_20724,N_18135,N_18299);
and U20725 (N_20725,N_18873,N_18897);
xnor U20726 (N_20726,N_17508,N_19529);
xor U20727 (N_20727,N_17981,N_18513);
or U20728 (N_20728,N_19515,N_18665);
or U20729 (N_20729,N_17627,N_18174);
xor U20730 (N_20730,N_18687,N_17847);
and U20731 (N_20731,N_19453,N_17819);
nor U20732 (N_20732,N_17719,N_18227);
xnor U20733 (N_20733,N_18468,N_17653);
xor U20734 (N_20734,N_18216,N_18953);
and U20735 (N_20735,N_19873,N_18480);
or U20736 (N_20736,N_18808,N_19436);
and U20737 (N_20737,N_19648,N_19527);
nor U20738 (N_20738,N_19003,N_18511);
nand U20739 (N_20739,N_19450,N_19006);
nor U20740 (N_20740,N_18099,N_18518);
and U20741 (N_20741,N_19839,N_17697);
or U20742 (N_20742,N_19231,N_18332);
and U20743 (N_20743,N_19891,N_19209);
nand U20744 (N_20744,N_18382,N_18061);
xnor U20745 (N_20745,N_19948,N_18190);
or U20746 (N_20746,N_19269,N_19885);
or U20747 (N_20747,N_19778,N_19429);
xor U20748 (N_20748,N_19213,N_18769);
xor U20749 (N_20749,N_19179,N_19985);
nor U20750 (N_20750,N_18678,N_19010);
nor U20751 (N_20751,N_18119,N_19395);
and U20752 (N_20752,N_18217,N_19080);
nand U20753 (N_20753,N_19646,N_17811);
xor U20754 (N_20754,N_18032,N_18360);
and U20755 (N_20755,N_19866,N_17831);
or U20756 (N_20756,N_18183,N_19153);
nor U20757 (N_20757,N_19984,N_18886);
nor U20758 (N_20758,N_19543,N_17545);
and U20759 (N_20759,N_19488,N_19168);
or U20760 (N_20760,N_18668,N_18004);
or U20761 (N_20761,N_18861,N_19055);
and U20762 (N_20762,N_19941,N_19744);
or U20763 (N_20763,N_19112,N_19451);
nand U20764 (N_20764,N_18471,N_19297);
nand U20765 (N_20765,N_17994,N_18576);
nand U20766 (N_20766,N_18026,N_19283);
and U20767 (N_20767,N_18964,N_18120);
or U20768 (N_20768,N_19278,N_19084);
or U20769 (N_20769,N_19373,N_17614);
nand U20770 (N_20770,N_19258,N_18298);
xnor U20771 (N_20771,N_19307,N_17562);
or U20772 (N_20772,N_18312,N_18881);
nand U20773 (N_20773,N_17975,N_18521);
or U20774 (N_20774,N_19664,N_19180);
nand U20775 (N_20775,N_19699,N_17948);
or U20776 (N_20776,N_18514,N_19199);
nor U20777 (N_20777,N_17724,N_19547);
nor U20778 (N_20778,N_18948,N_17973);
nor U20779 (N_20779,N_19530,N_18233);
xor U20780 (N_20780,N_19831,N_18824);
xor U20781 (N_20781,N_17788,N_18485);
and U20782 (N_20782,N_19558,N_19842);
nand U20783 (N_20783,N_18612,N_17843);
xor U20784 (N_20784,N_17797,N_19506);
and U20785 (N_20785,N_19198,N_19457);
or U20786 (N_20786,N_19051,N_19499);
or U20787 (N_20787,N_17698,N_18202);
or U20788 (N_20788,N_18849,N_17715);
or U20789 (N_20789,N_17550,N_18390);
and U20790 (N_20790,N_17983,N_18284);
nor U20791 (N_20791,N_17649,N_18517);
nor U20792 (N_20792,N_18799,N_18784);
nor U20793 (N_20793,N_19287,N_18889);
xor U20794 (N_20794,N_19516,N_19321);
nor U20795 (N_20795,N_17696,N_17613);
xnor U20796 (N_20796,N_18475,N_19733);
nor U20797 (N_20797,N_19651,N_19946);
nand U20798 (N_20798,N_17900,N_18996);
nand U20799 (N_20799,N_19755,N_19703);
and U20800 (N_20800,N_18746,N_17793);
xor U20801 (N_20801,N_19415,N_18370);
and U20802 (N_20802,N_18830,N_19658);
xnor U20803 (N_20803,N_17619,N_18426);
or U20804 (N_20804,N_19369,N_17514);
xnor U20805 (N_20805,N_17622,N_18378);
and U20806 (N_20806,N_19669,N_19613);
or U20807 (N_20807,N_17527,N_19604);
and U20808 (N_20808,N_19124,N_18157);
nor U20809 (N_20809,N_17608,N_19990);
xnor U20810 (N_20810,N_18724,N_18138);
nand U20811 (N_20811,N_19013,N_19107);
nor U20812 (N_20812,N_18122,N_18660);
nand U20813 (N_20813,N_17887,N_18231);
or U20814 (N_20814,N_18114,N_18690);
xor U20815 (N_20815,N_17889,N_18770);
nand U20816 (N_20816,N_18918,N_19960);
nand U20817 (N_20817,N_17859,N_17687);
or U20818 (N_20818,N_18739,N_17599);
xnor U20819 (N_20819,N_19205,N_19495);
and U20820 (N_20820,N_17856,N_17861);
or U20821 (N_20821,N_19727,N_17517);
and U20822 (N_20822,N_19503,N_18642);
xnor U20823 (N_20823,N_19870,N_18583);
xor U20824 (N_20824,N_18006,N_19955);
nand U20825 (N_20825,N_18250,N_17594);
nor U20826 (N_20826,N_19377,N_19599);
or U20827 (N_20827,N_19147,N_19040);
nand U20828 (N_20828,N_18538,N_18374);
and U20829 (N_20829,N_18895,N_19005);
nor U20830 (N_20830,N_19120,N_19402);
nand U20831 (N_20831,N_19884,N_19241);
nand U20832 (N_20832,N_18459,N_19989);
and U20833 (N_20833,N_19072,N_17908);
and U20834 (N_20834,N_18752,N_18575);
nand U20835 (N_20835,N_19196,N_17750);
nor U20836 (N_20836,N_19224,N_19363);
nor U20837 (N_20837,N_17854,N_19521);
xor U20838 (N_20838,N_19862,N_19096);
nand U20839 (N_20839,N_17524,N_18444);
nand U20840 (N_20840,N_18392,N_18133);
or U20841 (N_20841,N_19364,N_19644);
and U20842 (N_20842,N_18438,N_19257);
xor U20843 (N_20843,N_18630,N_19184);
nor U20844 (N_20844,N_19943,N_18307);
nor U20845 (N_20845,N_19517,N_17886);
xor U20846 (N_20846,N_18659,N_19890);
or U20847 (N_20847,N_19375,N_19032);
xnor U20848 (N_20848,N_19125,N_17536);
nor U20849 (N_20849,N_17760,N_18057);
or U20850 (N_20850,N_19618,N_18984);
nand U20851 (N_20851,N_17668,N_17718);
xnor U20852 (N_20852,N_18923,N_18121);
xnor U20853 (N_20853,N_19393,N_19918);
or U20854 (N_20854,N_18020,N_18796);
and U20855 (N_20855,N_17902,N_19028);
or U20856 (N_20856,N_18790,N_19174);
or U20857 (N_20857,N_18912,N_19719);
and U20858 (N_20858,N_18680,N_18682);
nand U20859 (N_20859,N_19957,N_18347);
and U20860 (N_20860,N_17654,N_17930);
or U20861 (N_20861,N_19887,N_19012);
or U20862 (N_20862,N_18751,N_18875);
nor U20863 (N_20863,N_19100,N_18800);
nand U20864 (N_20864,N_19729,N_18246);
nor U20865 (N_20865,N_18885,N_19553);
nand U20866 (N_20866,N_17986,N_18506);
nand U20867 (N_20867,N_18060,N_17960);
and U20868 (N_20868,N_18728,N_19838);
or U20869 (N_20869,N_18110,N_19899);
nor U20870 (N_20870,N_19389,N_19970);
and U20871 (N_20871,N_19105,N_19940);
xor U20872 (N_20872,N_18552,N_18876);
nand U20873 (N_20873,N_19068,N_18696);
nor U20874 (N_20874,N_18159,N_19237);
nor U20875 (N_20875,N_19974,N_19470);
and U20876 (N_20876,N_19765,N_18780);
nand U20877 (N_20877,N_17990,N_18754);
xnor U20878 (N_20878,N_17596,N_18376);
nand U20879 (N_20879,N_18283,N_18034);
nand U20880 (N_20880,N_19486,N_17968);
or U20881 (N_20881,N_18938,N_19827);
and U20882 (N_20882,N_17685,N_17638);
or U20883 (N_20883,N_17751,N_17921);
nand U20884 (N_20884,N_19902,N_18716);
or U20885 (N_20885,N_19169,N_18988);
or U20886 (N_20886,N_19559,N_19102);
nand U20887 (N_20887,N_18787,N_19316);
and U20888 (N_20888,N_18761,N_18939);
or U20889 (N_20889,N_18080,N_19892);
nor U20890 (N_20890,N_18603,N_18047);
and U20891 (N_20891,N_19339,N_19405);
xnor U20892 (N_20892,N_17938,N_19513);
and U20893 (N_20893,N_19162,N_19579);
or U20894 (N_20894,N_19444,N_19392);
nor U20895 (N_20895,N_19575,N_18901);
and U20896 (N_20896,N_19089,N_17555);
nand U20897 (N_20897,N_19002,N_18539);
or U20898 (N_20898,N_17589,N_19379);
xnor U20899 (N_20899,N_19325,N_18277);
xnor U20900 (N_20900,N_17661,N_18657);
or U20901 (N_20901,N_18036,N_19063);
nand U20902 (N_20902,N_19357,N_17725);
or U20903 (N_20903,N_19771,N_19920);
nand U20904 (N_20904,N_19401,N_19227);
xnor U20905 (N_20905,N_18905,N_19769);
nand U20906 (N_20906,N_19342,N_18092);
nor U20907 (N_20907,N_17528,N_17542);
xnor U20908 (N_20908,N_17941,N_18970);
nand U20909 (N_20909,N_19535,N_18007);
xnor U20910 (N_20910,N_18165,N_18011);
nor U20911 (N_20911,N_19212,N_19748);
nand U20912 (N_20912,N_17612,N_18349);
nor U20913 (N_20913,N_19851,N_19076);
or U20914 (N_20914,N_19472,N_18810);
nand U20915 (N_20915,N_19629,N_19973);
xnor U20916 (N_20916,N_19498,N_17588);
or U20917 (N_20917,N_19860,N_18158);
xnor U20918 (N_20918,N_19442,N_18530);
nand U20919 (N_20919,N_17754,N_19801);
and U20920 (N_20920,N_18712,N_17880);
nand U20921 (N_20921,N_17873,N_18564);
or U20922 (N_20922,N_18833,N_17877);
nand U20923 (N_20923,N_17695,N_19471);
and U20924 (N_20924,N_17553,N_19665);
xnor U20925 (N_20925,N_19856,N_19244);
nand U20926 (N_20926,N_17714,N_18259);
xor U20927 (N_20927,N_17561,N_17625);
nand U20928 (N_20928,N_19806,N_17519);
and U20929 (N_20929,N_18837,N_17775);
nor U20930 (N_20930,N_18915,N_17828);
or U20931 (N_20931,N_18274,N_19889);
xnor U20932 (N_20932,N_17546,N_17708);
or U20933 (N_20933,N_19408,N_19400);
and U20934 (N_20934,N_19944,N_18330);
nand U20935 (N_20935,N_18255,N_17648);
or U20936 (N_20936,N_17556,N_18645);
and U20937 (N_20937,N_19484,N_18943);
nand U20938 (N_20938,N_19035,N_17582);
xor U20939 (N_20939,N_18396,N_18479);
or U20940 (N_20940,N_19710,N_18364);
and U20941 (N_20941,N_18707,N_19163);
nand U20942 (N_20942,N_19927,N_17745);
and U20943 (N_20943,N_18669,N_19589);
nor U20944 (N_20944,N_18319,N_19683);
xor U20945 (N_20945,N_19192,N_18501);
and U20946 (N_20946,N_19897,N_19242);
xor U20947 (N_20947,N_18033,N_18409);
or U20948 (N_20948,N_19215,N_19643);
nand U20949 (N_20949,N_18667,N_18976);
or U20950 (N_20950,N_19280,N_19691);
or U20951 (N_20951,N_19106,N_18188);
or U20952 (N_20952,N_18412,N_17558);
nand U20953 (N_20953,N_17650,N_17652);
and U20954 (N_20954,N_19059,N_17660);
or U20955 (N_20955,N_18891,N_19403);
nand U20956 (N_20956,N_18243,N_19678);
or U20957 (N_20957,N_17805,N_18407);
nor U20958 (N_20958,N_18339,N_19317);
nand U20959 (N_20959,N_18954,N_19291);
xor U20960 (N_20960,N_18354,N_18027);
or U20961 (N_20961,N_18066,N_17575);
and U20962 (N_20962,N_18710,N_17935);
or U20963 (N_20963,N_17946,N_18186);
nand U20964 (N_20964,N_19338,N_18067);
nor U20965 (N_20965,N_18473,N_18367);
nand U20966 (N_20966,N_18662,N_19347);
or U20967 (N_20967,N_18096,N_18709);
nor U20968 (N_20968,N_18293,N_18229);
and U20969 (N_20969,N_18794,N_19587);
or U20970 (N_20970,N_17707,N_19738);
xor U20971 (N_20971,N_17630,N_18546);
or U20972 (N_20972,N_17952,N_19647);
or U20973 (N_20973,N_19650,N_18826);
or U20974 (N_20974,N_17836,N_18044);
or U20975 (N_20975,N_18866,N_17642);
and U20976 (N_20976,N_19732,N_17560);
or U20977 (N_20977,N_19739,N_18171);
nor U20978 (N_20978,N_19265,N_18714);
xnor U20979 (N_20979,N_19818,N_18532);
and U20980 (N_20980,N_18524,N_19465);
nand U20981 (N_20981,N_19789,N_18318);
nand U20982 (N_20982,N_19077,N_17643);
and U20983 (N_20983,N_18030,N_17610);
xor U20984 (N_20984,N_18483,N_17996);
xor U20985 (N_20985,N_19417,N_19078);
xor U20986 (N_20986,N_19346,N_19877);
nor U20987 (N_20987,N_19146,N_19501);
and U20988 (N_20988,N_18989,N_17976);
xor U20989 (N_20989,N_18516,N_18663);
xnor U20990 (N_20990,N_19813,N_18149);
nor U20991 (N_20991,N_18781,N_18081);
nor U20992 (N_20992,N_17988,N_17871);
nand U20993 (N_20993,N_19865,N_19036);
xnor U20994 (N_20994,N_19135,N_18248);
and U20995 (N_20995,N_17636,N_17940);
nor U20996 (N_20996,N_19293,N_18192);
nor U20997 (N_20997,N_19422,N_18189);
nor U20998 (N_20998,N_18729,N_17656);
nor U20999 (N_20999,N_18075,N_19494);
nor U21000 (N_21000,N_17806,N_19551);
xor U21001 (N_21001,N_17918,N_19965);
and U21002 (N_21002,N_18725,N_18509);
and U21003 (N_21003,N_18334,N_18656);
xor U21004 (N_21004,N_18602,N_18887);
xor U21005 (N_21005,N_19524,N_18089);
and U21006 (N_21006,N_19004,N_18626);
nand U21007 (N_21007,N_19464,N_17761);
and U21008 (N_21008,N_19768,N_18205);
nor U21009 (N_21009,N_19294,N_19118);
nor U21010 (N_21010,N_18251,N_17738);
xnor U21011 (N_21011,N_18366,N_18474);
nor U21012 (N_21012,N_19303,N_19622);
or U21013 (N_21013,N_18499,N_18393);
nand U21014 (N_21014,N_19996,N_19534);
nor U21015 (N_21015,N_18132,N_18325);
xnor U21016 (N_21016,N_17644,N_19693);
and U21017 (N_21017,N_19688,N_19438);
nor U21018 (N_21018,N_18346,N_18265);
or U21019 (N_21019,N_18314,N_19252);
xor U21020 (N_21020,N_19099,N_17680);
nand U21021 (N_21021,N_19672,N_19433);
xnor U21022 (N_21022,N_19343,N_19840);
xnor U21023 (N_21023,N_17576,N_17507);
or U21024 (N_21024,N_18777,N_18451);
xnor U21025 (N_21025,N_17984,N_19662);
xnor U21026 (N_21026,N_19544,N_18199);
nand U21027 (N_21027,N_18152,N_18415);
nor U21028 (N_21028,N_19574,N_18002);
and U21029 (N_21029,N_19518,N_18201);
nand U21030 (N_21030,N_17506,N_17972);
nor U21031 (N_21031,N_18009,N_17730);
nand U21032 (N_21032,N_19070,N_17912);
nand U21033 (N_21033,N_17538,N_19734);
nor U21034 (N_21034,N_18531,N_18971);
xor U21035 (N_21035,N_18324,N_19853);
nand U21036 (N_21036,N_18704,N_19057);
nor U21037 (N_21037,N_18730,N_18402);
xnor U21038 (N_21038,N_17666,N_19784);
nor U21039 (N_21039,N_19421,N_18972);
and U21040 (N_21040,N_17777,N_18048);
xnor U21041 (N_21041,N_18774,N_19817);
or U21042 (N_21042,N_17939,N_19073);
or U21043 (N_21043,N_19298,N_19905);
nor U21044 (N_21044,N_19137,N_19997);
and U21045 (N_21045,N_17822,N_19413);
xor U21046 (N_21046,N_18773,N_19545);
xnor U21047 (N_21047,N_18435,N_19350);
and U21048 (N_21048,N_19046,N_18904);
nor U21049 (N_21049,N_19206,N_19060);
nand U21050 (N_21050,N_19874,N_19706);
xnor U21051 (N_21051,N_18156,N_19419);
xor U21052 (N_21052,N_19140,N_17515);
xnor U21053 (N_21053,N_18305,N_19341);
or U21054 (N_21054,N_19593,N_18313);
and U21055 (N_21055,N_18257,N_18785);
and U21056 (N_21056,N_17571,N_17801);
xor U21057 (N_21057,N_17579,N_19680);
and U21058 (N_21058,N_18422,N_18778);
and U21059 (N_21059,N_19549,N_17867);
nand U21060 (N_21060,N_19657,N_19414);
xor U21061 (N_21061,N_18237,N_19200);
nand U21062 (N_21062,N_19358,N_18029);
xor U21063 (N_21063,N_17665,N_19584);
xnor U21064 (N_21064,N_18486,N_19914);
and U21065 (N_21065,N_17876,N_18124);
or U21066 (N_21066,N_18161,N_19249);
xor U21067 (N_21067,N_19136,N_19993);
and U21068 (N_21068,N_18063,N_19396);
nand U21069 (N_21069,N_17785,N_19382);
xnor U21070 (N_21070,N_18331,N_19095);
or U21071 (N_21071,N_18098,N_18162);
xor U21072 (N_21072,N_18929,N_19412);
nand U21073 (N_21073,N_18960,N_19913);
nor U21074 (N_21074,N_18001,N_19474);
nor U21075 (N_21075,N_19652,N_18113);
or U21076 (N_21076,N_18816,N_18566);
nand U21077 (N_21077,N_18706,N_19807);
nand U21078 (N_21078,N_18381,N_19528);
xor U21079 (N_21079,N_18172,N_18828);
xnor U21080 (N_21080,N_19816,N_18404);
or U21081 (N_21081,N_18388,N_17544);
nor U21082 (N_21082,N_18851,N_19656);
or U21083 (N_21083,N_18520,N_18757);
nor U21084 (N_21084,N_18289,N_19775);
nor U21085 (N_21085,N_19271,N_19563);
nor U21086 (N_21086,N_18249,N_18329);
nand U21087 (N_21087,N_18180,N_19597);
and U21088 (N_21088,N_18899,N_19928);
nor U21089 (N_21089,N_18744,N_19510);
and U21090 (N_21090,N_18348,N_18519);
nor U21091 (N_21091,N_18526,N_17537);
nand U21092 (N_21092,N_18054,N_18677);
xnor U21093 (N_21093,N_18252,N_18453);
nand U21094 (N_21094,N_19478,N_18275);
nor U21095 (N_21095,N_17577,N_17866);
or U21096 (N_21096,N_19602,N_19982);
nor U21097 (N_21097,N_19337,N_19723);
nor U21098 (N_21098,N_17597,N_19731);
nand U21099 (N_21099,N_17700,N_19176);
and U21100 (N_21100,N_19560,N_18083);
nor U21101 (N_21101,N_17518,N_19779);
nor U21102 (N_21102,N_19898,N_18394);
and U21103 (N_21103,N_18722,N_18553);
and U21104 (N_21104,N_18949,N_19141);
xnor U21105 (N_21105,N_19880,N_19399);
and U21106 (N_21106,N_19926,N_17916);
xnor U21107 (N_21107,N_18070,N_18813);
and U21108 (N_21108,N_18000,N_19038);
xor U21109 (N_21109,N_19857,N_18209);
or U21110 (N_21110,N_19065,N_19795);
nand U21111 (N_21111,N_17735,N_18856);
xor U21112 (N_21112,N_17741,N_19211);
nand U21113 (N_21113,N_17890,N_19409);
nor U21114 (N_21114,N_19266,N_18807);
xor U21115 (N_21115,N_18208,N_18139);
nand U21116 (N_21116,N_19259,N_19299);
xor U21117 (N_21117,N_19504,N_17851);
nand U21118 (N_21118,N_17703,N_19822);
and U21119 (N_21119,N_18014,N_18962);
and U21120 (N_21120,N_19345,N_18841);
nor U21121 (N_21121,N_17624,N_19888);
or U21122 (N_21122,N_18919,N_17772);
or U21123 (N_21123,N_18040,N_17563);
xnor U21124 (N_21124,N_17834,N_18832);
and U21125 (N_21125,N_18727,N_18448);
or U21126 (N_21126,N_17711,N_18802);
xor U21127 (N_21127,N_19632,N_18272);
xnor U21128 (N_21128,N_18614,N_19797);
nor U21129 (N_21129,N_19138,N_18914);
nand U21130 (N_21130,N_17728,N_19830);
and U21131 (N_21131,N_18578,N_19071);
nor U21132 (N_21132,N_19170,N_18821);
nor U21133 (N_21133,N_18791,N_19062);
xor U21134 (N_21134,N_17824,N_17799);
and U21135 (N_21135,N_18059,N_19432);
and U21136 (N_21136,N_18924,N_17727);
and U21137 (N_21137,N_18464,N_18401);
xnor U21138 (N_21138,N_19592,N_17954);
xor U21139 (N_21139,N_19327,N_18582);
nand U21140 (N_21140,N_18425,N_18734);
and U21141 (N_21141,N_19284,N_19785);
xor U21142 (N_21142,N_17818,N_19268);
and U21143 (N_21143,N_17620,N_18405);
or U21144 (N_21144,N_19676,N_18525);
or U21145 (N_21145,N_17623,N_18619);
and U21146 (N_21146,N_18069,N_19896);
and U21147 (N_21147,N_19476,N_18326);
xor U21148 (N_21148,N_18338,N_18104);
nor U21149 (N_21149,N_18920,N_19858);
nor U21150 (N_21150,N_17802,N_19204);
nor U21151 (N_21151,N_18417,N_19726);
xnor U21152 (N_21152,N_19331,N_19981);
xor U21153 (N_21153,N_18117,N_18534);
nor U21154 (N_21154,N_18377,N_19218);
nand U21155 (N_21155,N_19440,N_17586);
xnor U21156 (N_21156,N_18831,N_19999);
xnor U21157 (N_21157,N_19491,N_18829);
nor U21158 (N_21158,N_18756,N_18336);
or U21159 (N_21159,N_18921,N_18429);
and U21160 (N_21160,N_18134,N_18871);
xnor U21161 (N_21161,N_19463,N_18587);
nand U21162 (N_21162,N_18493,N_18847);
xnor U21163 (N_21163,N_18223,N_19684);
xor U21164 (N_21164,N_19021,N_17920);
xor U21165 (N_21165,N_18975,N_18858);
nor U21166 (N_21166,N_18705,N_17857);
nor U21167 (N_21167,N_19568,N_19217);
and U21168 (N_21168,N_19823,N_17953);
nand U21169 (N_21169,N_18743,N_17647);
nand U21170 (N_21170,N_17645,N_19275);
nor U21171 (N_21171,N_17931,N_17771);
or U21172 (N_21172,N_19067,N_19776);
and U21173 (N_21173,N_19404,N_18234);
nor U21174 (N_21174,N_19050,N_18214);
or U21175 (N_21175,N_19505,N_18344);
and U21176 (N_21176,N_17543,N_19360);
and U21177 (N_21177,N_18427,N_17531);
or U21178 (N_21178,N_17592,N_19011);
nand U21179 (N_21179,N_19309,N_18358);
or U21180 (N_21180,N_19064,N_19362);
or U21181 (N_21181,N_19131,N_19750);
nor U21182 (N_21182,N_18267,N_18397);
xnor U21183 (N_21183,N_18285,N_19991);
nor U21184 (N_21184,N_18944,N_19677);
and U21185 (N_21185,N_19793,N_18140);
nor U21186 (N_21186,N_18198,N_17580);
nand U21187 (N_21187,N_18488,N_18726);
xnor U21188 (N_21188,N_18550,N_18084);
xor U21189 (N_21189,N_19306,N_18558);
or U21190 (N_21190,N_18718,N_18136);
xor U21191 (N_21191,N_17523,N_17615);
nand U21192 (N_21192,N_18053,N_19509);
nor U21193 (N_21193,N_19026,N_19376);
or U21194 (N_21194,N_17978,N_18242);
nor U21195 (N_21195,N_19381,N_19835);
nor U21196 (N_21196,N_19546,N_17881);
or U21197 (N_21197,N_19687,N_19000);
or U21198 (N_21198,N_18655,N_18071);
nand U21199 (N_21199,N_18469,N_19481);
xnor U21200 (N_21200,N_17605,N_18699);
nor U21201 (N_21201,N_17997,N_19302);
nand U21202 (N_21202,N_19617,N_17662);
or U21203 (N_21203,N_18995,N_19655);
or U21204 (N_21204,N_17817,N_19736);
nand U21205 (N_21205,N_18341,N_18410);
xor U21206 (N_21206,N_19142,N_19854);
and U21207 (N_21207,N_18617,N_19883);
nor U21208 (N_21208,N_17839,N_17709);
xnor U21209 (N_21209,N_18916,N_17823);
nor U21210 (N_21210,N_18835,N_19819);
or U21211 (N_21211,N_19311,N_18613);
nor U21212 (N_21212,N_18640,N_17637);
or U21213 (N_21213,N_19496,N_19007);
or U21214 (N_21214,N_19855,N_18549);
nand U21215 (N_21215,N_19315,N_18490);
xnor U21216 (N_21216,N_19766,N_18711);
and U21217 (N_21217,N_18082,N_19172);
and U21218 (N_21218,N_18185,N_18672);
or U21219 (N_21219,N_17766,N_18941);
nor U21220 (N_21220,N_19349,N_19634);
nand U21221 (N_21221,N_19081,N_19365);
and U21222 (N_21222,N_18567,N_18309);
nand U21223 (N_21223,N_18101,N_17667);
nand U21224 (N_21224,N_17934,N_17850);
xnor U21225 (N_21225,N_19274,N_19950);
nor U21226 (N_21226,N_18024,N_18537);
xor U21227 (N_21227,N_19932,N_18955);
nand U21228 (N_21228,N_19964,N_19836);
or U21229 (N_21229,N_18647,N_18592);
nor U21230 (N_21230,N_18765,N_19690);
nand U21231 (N_21231,N_19368,N_18239);
and U21232 (N_21232,N_19761,N_17503);
xnor U21233 (N_21233,N_19792,N_19469);
nor U21234 (N_21234,N_19110,N_17872);
or U21235 (N_21235,N_18273,N_18454);
nand U21236 (N_21236,N_18999,N_19758);
nand U21237 (N_21237,N_19001,N_18926);
and U21238 (N_21238,N_17753,N_17852);
or U21239 (N_21239,N_17955,N_19596);
and U21240 (N_21240,N_17932,N_18056);
xor U21241 (N_21241,N_17554,N_18176);
nor U21242 (N_21242,N_18737,N_18766);
nor U21243 (N_21243,N_18594,N_19207);
and U21244 (N_21244,N_17864,N_19961);
nand U21245 (N_21245,N_19320,N_18042);
and U21246 (N_21246,N_17565,N_19452);
or U21247 (N_21247,N_19406,N_17601);
or U21248 (N_21248,N_18894,N_19230);
or U21249 (N_21249,N_18477,N_19757);
or U21250 (N_21250,N_17733,N_17920);
nor U21251 (N_21251,N_18301,N_19943);
and U21252 (N_21252,N_18061,N_17689);
nor U21253 (N_21253,N_18729,N_18411);
nor U21254 (N_21254,N_17529,N_19318);
or U21255 (N_21255,N_17683,N_19241);
nand U21256 (N_21256,N_19288,N_18953);
or U21257 (N_21257,N_18757,N_17742);
nor U21258 (N_21258,N_17974,N_17785);
nand U21259 (N_21259,N_17651,N_17762);
nand U21260 (N_21260,N_18034,N_18385);
and U21261 (N_21261,N_18269,N_18664);
nand U21262 (N_21262,N_19255,N_17676);
nand U21263 (N_21263,N_18110,N_17895);
nor U21264 (N_21264,N_19930,N_19985);
and U21265 (N_21265,N_17684,N_19272);
xor U21266 (N_21266,N_18222,N_19526);
or U21267 (N_21267,N_17505,N_18811);
xnor U21268 (N_21268,N_18504,N_19552);
nand U21269 (N_21269,N_19945,N_19807);
and U21270 (N_21270,N_17714,N_18600);
and U21271 (N_21271,N_18932,N_17742);
xor U21272 (N_21272,N_19938,N_19162);
nor U21273 (N_21273,N_18348,N_19314);
xnor U21274 (N_21274,N_18226,N_19274);
and U21275 (N_21275,N_18470,N_19245);
nand U21276 (N_21276,N_18594,N_18970);
and U21277 (N_21277,N_17955,N_18171);
xnor U21278 (N_21278,N_19139,N_18286);
and U21279 (N_21279,N_18129,N_19735);
nor U21280 (N_21280,N_18835,N_19274);
nand U21281 (N_21281,N_18252,N_18287);
or U21282 (N_21282,N_18682,N_18288);
nand U21283 (N_21283,N_18090,N_19038);
and U21284 (N_21284,N_19380,N_18182);
and U21285 (N_21285,N_18813,N_17814);
xor U21286 (N_21286,N_18991,N_17937);
or U21287 (N_21287,N_18599,N_19824);
or U21288 (N_21288,N_17611,N_19200);
xor U21289 (N_21289,N_18456,N_17550);
nand U21290 (N_21290,N_18349,N_19634);
nand U21291 (N_21291,N_17694,N_18276);
and U21292 (N_21292,N_18449,N_19426);
or U21293 (N_21293,N_19867,N_19327);
or U21294 (N_21294,N_18958,N_17621);
nor U21295 (N_21295,N_17608,N_17931);
or U21296 (N_21296,N_18334,N_19381);
nand U21297 (N_21297,N_17561,N_18736);
xnor U21298 (N_21298,N_18560,N_18286);
xnor U21299 (N_21299,N_18344,N_18351);
xnor U21300 (N_21300,N_17745,N_18341);
nor U21301 (N_21301,N_17827,N_18383);
and U21302 (N_21302,N_17898,N_19315);
nand U21303 (N_21303,N_19259,N_18029);
or U21304 (N_21304,N_18752,N_17967);
nor U21305 (N_21305,N_19326,N_19902);
or U21306 (N_21306,N_18642,N_19096);
and U21307 (N_21307,N_19365,N_18864);
xor U21308 (N_21308,N_18419,N_19400);
nor U21309 (N_21309,N_18974,N_18952);
or U21310 (N_21310,N_19829,N_19871);
nand U21311 (N_21311,N_18417,N_18657);
nand U21312 (N_21312,N_18815,N_19569);
or U21313 (N_21313,N_19661,N_19663);
nand U21314 (N_21314,N_19543,N_19156);
or U21315 (N_21315,N_17541,N_19986);
nor U21316 (N_21316,N_19445,N_19433);
xnor U21317 (N_21317,N_19897,N_18545);
xor U21318 (N_21318,N_18859,N_18015);
xnor U21319 (N_21319,N_19765,N_18987);
nand U21320 (N_21320,N_18522,N_18606);
nor U21321 (N_21321,N_18796,N_18639);
and U21322 (N_21322,N_18863,N_18676);
nor U21323 (N_21323,N_18250,N_18237);
nor U21324 (N_21324,N_17662,N_19163);
xnor U21325 (N_21325,N_17556,N_19330);
and U21326 (N_21326,N_18556,N_19131);
xor U21327 (N_21327,N_18610,N_17763);
xnor U21328 (N_21328,N_18755,N_19795);
or U21329 (N_21329,N_19297,N_19269);
xor U21330 (N_21330,N_18867,N_19660);
nor U21331 (N_21331,N_17924,N_18773);
or U21332 (N_21332,N_19674,N_19317);
xor U21333 (N_21333,N_18997,N_18581);
or U21334 (N_21334,N_19888,N_17729);
or U21335 (N_21335,N_19005,N_19361);
xnor U21336 (N_21336,N_19707,N_17995);
and U21337 (N_21337,N_19641,N_19447);
and U21338 (N_21338,N_19775,N_18086);
nor U21339 (N_21339,N_19748,N_17624);
and U21340 (N_21340,N_18224,N_18190);
nand U21341 (N_21341,N_18739,N_19816);
xor U21342 (N_21342,N_17699,N_18524);
nand U21343 (N_21343,N_19757,N_19027);
nor U21344 (N_21344,N_19983,N_19299);
nor U21345 (N_21345,N_19281,N_18388);
nand U21346 (N_21346,N_18062,N_17536);
nor U21347 (N_21347,N_18895,N_19081);
nor U21348 (N_21348,N_18581,N_17639);
or U21349 (N_21349,N_18383,N_19285);
xnor U21350 (N_21350,N_17932,N_19257);
and U21351 (N_21351,N_18733,N_18959);
nand U21352 (N_21352,N_19095,N_19790);
or U21353 (N_21353,N_19307,N_19292);
xnor U21354 (N_21354,N_17808,N_18959);
nand U21355 (N_21355,N_18456,N_18045);
or U21356 (N_21356,N_17608,N_17778);
or U21357 (N_21357,N_19551,N_17819);
nand U21358 (N_21358,N_19518,N_18799);
or U21359 (N_21359,N_17722,N_18769);
xnor U21360 (N_21360,N_18701,N_19455);
xnor U21361 (N_21361,N_19417,N_18445);
or U21362 (N_21362,N_18066,N_19021);
and U21363 (N_21363,N_18754,N_17797);
or U21364 (N_21364,N_18897,N_19674);
nand U21365 (N_21365,N_17679,N_19028);
nor U21366 (N_21366,N_18776,N_18074);
nor U21367 (N_21367,N_19516,N_17758);
nor U21368 (N_21368,N_18439,N_19891);
or U21369 (N_21369,N_19121,N_18441);
or U21370 (N_21370,N_19411,N_18572);
and U21371 (N_21371,N_17998,N_18974);
nand U21372 (N_21372,N_19554,N_17617);
xor U21373 (N_21373,N_18082,N_18526);
and U21374 (N_21374,N_18898,N_18418);
or U21375 (N_21375,N_18162,N_17705);
xor U21376 (N_21376,N_19151,N_19575);
nand U21377 (N_21377,N_17580,N_19844);
nor U21378 (N_21378,N_19302,N_18753);
nor U21379 (N_21379,N_17655,N_18418);
xnor U21380 (N_21380,N_18103,N_19330);
or U21381 (N_21381,N_19258,N_19472);
nor U21382 (N_21382,N_19512,N_19380);
or U21383 (N_21383,N_18182,N_18942);
nor U21384 (N_21384,N_18914,N_17912);
nor U21385 (N_21385,N_19275,N_19663);
and U21386 (N_21386,N_19090,N_19159);
xnor U21387 (N_21387,N_18859,N_19487);
nor U21388 (N_21388,N_17802,N_19516);
xor U21389 (N_21389,N_18275,N_18477);
xnor U21390 (N_21390,N_19517,N_18156);
nor U21391 (N_21391,N_19072,N_17702);
nor U21392 (N_21392,N_18600,N_19439);
nor U21393 (N_21393,N_18161,N_19821);
xor U21394 (N_21394,N_18045,N_19519);
xor U21395 (N_21395,N_18982,N_18995);
nand U21396 (N_21396,N_17977,N_18958);
and U21397 (N_21397,N_18995,N_18908);
xor U21398 (N_21398,N_19410,N_19190);
nor U21399 (N_21399,N_18216,N_19269);
and U21400 (N_21400,N_19764,N_19575);
nand U21401 (N_21401,N_19825,N_17700);
nor U21402 (N_21402,N_18425,N_17715);
or U21403 (N_21403,N_18318,N_19277);
and U21404 (N_21404,N_18112,N_18624);
and U21405 (N_21405,N_17775,N_17882);
nand U21406 (N_21406,N_18303,N_18012);
xnor U21407 (N_21407,N_18706,N_17522);
nand U21408 (N_21408,N_18299,N_18624);
xnor U21409 (N_21409,N_18817,N_19796);
nand U21410 (N_21410,N_18704,N_18496);
nand U21411 (N_21411,N_18286,N_18646);
xnor U21412 (N_21412,N_19583,N_19208);
nor U21413 (N_21413,N_17939,N_17940);
xnor U21414 (N_21414,N_17520,N_19994);
and U21415 (N_21415,N_19666,N_18351);
xnor U21416 (N_21416,N_17899,N_18374);
nor U21417 (N_21417,N_19593,N_18763);
and U21418 (N_21418,N_19840,N_18726);
xor U21419 (N_21419,N_19817,N_19773);
xnor U21420 (N_21420,N_18566,N_19955);
xor U21421 (N_21421,N_17819,N_18399);
nand U21422 (N_21422,N_19439,N_18099);
nand U21423 (N_21423,N_18529,N_18310);
or U21424 (N_21424,N_19951,N_18655);
nor U21425 (N_21425,N_17631,N_18476);
xor U21426 (N_21426,N_19823,N_19363);
nand U21427 (N_21427,N_18881,N_17772);
or U21428 (N_21428,N_18846,N_17790);
nand U21429 (N_21429,N_19613,N_18021);
nor U21430 (N_21430,N_19430,N_18271);
nor U21431 (N_21431,N_19545,N_19834);
or U21432 (N_21432,N_19418,N_18926);
or U21433 (N_21433,N_18562,N_19547);
nor U21434 (N_21434,N_18156,N_18590);
nand U21435 (N_21435,N_18456,N_17796);
nor U21436 (N_21436,N_18893,N_17542);
xor U21437 (N_21437,N_19883,N_18685);
xnor U21438 (N_21438,N_19162,N_19583);
and U21439 (N_21439,N_18242,N_17863);
nor U21440 (N_21440,N_19669,N_18854);
nor U21441 (N_21441,N_19840,N_19803);
xnor U21442 (N_21442,N_18251,N_18498);
and U21443 (N_21443,N_18706,N_19299);
xnor U21444 (N_21444,N_19772,N_18686);
nor U21445 (N_21445,N_18201,N_19661);
xor U21446 (N_21446,N_18824,N_19393);
and U21447 (N_21447,N_18007,N_19748);
xor U21448 (N_21448,N_19252,N_19873);
and U21449 (N_21449,N_18279,N_19629);
xnor U21450 (N_21450,N_18452,N_18675);
nor U21451 (N_21451,N_18755,N_18524);
xnor U21452 (N_21452,N_18821,N_19128);
or U21453 (N_21453,N_18638,N_19625);
or U21454 (N_21454,N_19623,N_17526);
nor U21455 (N_21455,N_19737,N_19142);
nand U21456 (N_21456,N_17830,N_17770);
or U21457 (N_21457,N_18095,N_17964);
xnor U21458 (N_21458,N_18775,N_18238);
and U21459 (N_21459,N_17768,N_18497);
nand U21460 (N_21460,N_17694,N_17635);
and U21461 (N_21461,N_18759,N_18340);
nor U21462 (N_21462,N_19623,N_17922);
xnor U21463 (N_21463,N_18786,N_19649);
or U21464 (N_21464,N_18961,N_18259);
nor U21465 (N_21465,N_18794,N_17658);
nand U21466 (N_21466,N_17831,N_18817);
nand U21467 (N_21467,N_18448,N_19678);
xor U21468 (N_21468,N_18944,N_18409);
and U21469 (N_21469,N_19736,N_19385);
and U21470 (N_21470,N_17822,N_17762);
or U21471 (N_21471,N_19937,N_19551);
nand U21472 (N_21472,N_17989,N_18185);
and U21473 (N_21473,N_17618,N_19508);
nand U21474 (N_21474,N_18830,N_17896);
nor U21475 (N_21475,N_18822,N_18444);
or U21476 (N_21476,N_18478,N_18893);
nand U21477 (N_21477,N_19714,N_18303);
nand U21478 (N_21478,N_19264,N_18741);
and U21479 (N_21479,N_19400,N_18424);
and U21480 (N_21480,N_18933,N_18527);
or U21481 (N_21481,N_17829,N_19247);
or U21482 (N_21482,N_18752,N_17993);
and U21483 (N_21483,N_19628,N_18163);
or U21484 (N_21484,N_18179,N_17977);
or U21485 (N_21485,N_17509,N_19492);
nand U21486 (N_21486,N_17749,N_17728);
xnor U21487 (N_21487,N_19215,N_18067);
or U21488 (N_21488,N_17590,N_19451);
nor U21489 (N_21489,N_17507,N_17952);
or U21490 (N_21490,N_17593,N_19650);
xnor U21491 (N_21491,N_18585,N_17926);
nand U21492 (N_21492,N_18504,N_19911);
xor U21493 (N_21493,N_17659,N_18120);
or U21494 (N_21494,N_18451,N_18490);
nand U21495 (N_21495,N_19912,N_19586);
nor U21496 (N_21496,N_19184,N_19538);
nand U21497 (N_21497,N_19011,N_19540);
xor U21498 (N_21498,N_17862,N_17758);
xnor U21499 (N_21499,N_17724,N_19288);
nand U21500 (N_21500,N_19350,N_18330);
nand U21501 (N_21501,N_19517,N_18609);
and U21502 (N_21502,N_19207,N_19839);
and U21503 (N_21503,N_17629,N_18483);
xnor U21504 (N_21504,N_18471,N_18860);
xnor U21505 (N_21505,N_19406,N_19024);
xnor U21506 (N_21506,N_17552,N_18328);
and U21507 (N_21507,N_19294,N_17718);
nor U21508 (N_21508,N_19239,N_18472);
nand U21509 (N_21509,N_18448,N_19199);
nor U21510 (N_21510,N_19083,N_19240);
nand U21511 (N_21511,N_18893,N_19854);
xor U21512 (N_21512,N_18845,N_17775);
nand U21513 (N_21513,N_19283,N_18534);
and U21514 (N_21514,N_19585,N_18898);
xor U21515 (N_21515,N_19407,N_18705);
nand U21516 (N_21516,N_18111,N_19872);
and U21517 (N_21517,N_17703,N_19218);
and U21518 (N_21518,N_19716,N_19864);
nand U21519 (N_21519,N_19207,N_17652);
nor U21520 (N_21520,N_18263,N_18893);
or U21521 (N_21521,N_18338,N_18904);
nand U21522 (N_21522,N_19071,N_18655);
nor U21523 (N_21523,N_19666,N_18545);
nor U21524 (N_21524,N_18553,N_18675);
nand U21525 (N_21525,N_19876,N_17927);
or U21526 (N_21526,N_18160,N_18589);
and U21527 (N_21527,N_19760,N_18333);
nor U21528 (N_21528,N_18002,N_19692);
nand U21529 (N_21529,N_17759,N_19613);
or U21530 (N_21530,N_17551,N_18656);
or U21531 (N_21531,N_18130,N_19285);
nor U21532 (N_21532,N_19694,N_19905);
nand U21533 (N_21533,N_18733,N_19900);
or U21534 (N_21534,N_19146,N_18419);
or U21535 (N_21535,N_19666,N_19860);
xor U21536 (N_21536,N_19257,N_19869);
or U21537 (N_21537,N_19393,N_18287);
xnor U21538 (N_21538,N_19817,N_19729);
xor U21539 (N_21539,N_19644,N_19378);
nand U21540 (N_21540,N_19756,N_18647);
and U21541 (N_21541,N_18273,N_17580);
nand U21542 (N_21542,N_18452,N_18698);
xor U21543 (N_21543,N_18705,N_18089);
and U21544 (N_21544,N_18627,N_17651);
or U21545 (N_21545,N_19524,N_19476);
nor U21546 (N_21546,N_17882,N_19869);
nor U21547 (N_21547,N_17922,N_19194);
or U21548 (N_21548,N_18418,N_18294);
nand U21549 (N_21549,N_18834,N_19317);
nor U21550 (N_21550,N_19583,N_18366);
or U21551 (N_21551,N_18483,N_19282);
nor U21552 (N_21552,N_18600,N_17592);
nand U21553 (N_21553,N_17775,N_18448);
nand U21554 (N_21554,N_19527,N_18846);
xnor U21555 (N_21555,N_18954,N_19370);
or U21556 (N_21556,N_19198,N_19256);
nand U21557 (N_21557,N_18021,N_19363);
nand U21558 (N_21558,N_19966,N_17689);
and U21559 (N_21559,N_19928,N_17655);
nor U21560 (N_21560,N_17692,N_19508);
nor U21561 (N_21561,N_19440,N_19117);
and U21562 (N_21562,N_18349,N_19968);
and U21563 (N_21563,N_19032,N_18050);
or U21564 (N_21564,N_19229,N_19756);
xor U21565 (N_21565,N_19301,N_18825);
nand U21566 (N_21566,N_19587,N_17763);
nand U21567 (N_21567,N_17593,N_17911);
xnor U21568 (N_21568,N_18961,N_18617);
or U21569 (N_21569,N_19299,N_18170);
nor U21570 (N_21570,N_19293,N_18540);
and U21571 (N_21571,N_19206,N_19409);
nand U21572 (N_21572,N_19375,N_18959);
nand U21573 (N_21573,N_19867,N_17982);
xor U21574 (N_21574,N_18189,N_18410);
nor U21575 (N_21575,N_18744,N_19219);
nor U21576 (N_21576,N_18052,N_18184);
or U21577 (N_21577,N_19894,N_19102);
nand U21578 (N_21578,N_18975,N_18630);
nor U21579 (N_21579,N_18268,N_18673);
or U21580 (N_21580,N_18142,N_18126);
nor U21581 (N_21581,N_18033,N_19487);
or U21582 (N_21582,N_18890,N_18527);
or U21583 (N_21583,N_17607,N_18452);
xnor U21584 (N_21584,N_17907,N_18605);
nor U21585 (N_21585,N_17687,N_19274);
nand U21586 (N_21586,N_18106,N_18956);
nand U21587 (N_21587,N_18308,N_19742);
nor U21588 (N_21588,N_19823,N_19153);
nand U21589 (N_21589,N_17700,N_18131);
nand U21590 (N_21590,N_17675,N_18956);
nor U21591 (N_21591,N_18560,N_18371);
and U21592 (N_21592,N_19789,N_19234);
and U21593 (N_21593,N_18036,N_17518);
xnor U21594 (N_21594,N_18227,N_19021);
nand U21595 (N_21595,N_19693,N_19157);
nor U21596 (N_21596,N_17674,N_19020);
or U21597 (N_21597,N_19787,N_17899);
or U21598 (N_21598,N_17957,N_19512);
nor U21599 (N_21599,N_17564,N_19859);
xnor U21600 (N_21600,N_18126,N_19743);
nand U21601 (N_21601,N_19310,N_18954);
xnor U21602 (N_21602,N_18871,N_19393);
nand U21603 (N_21603,N_19563,N_19440);
nor U21604 (N_21604,N_17652,N_19303);
nor U21605 (N_21605,N_18373,N_18876);
xnor U21606 (N_21606,N_18143,N_19362);
xnor U21607 (N_21607,N_19010,N_18163);
xor U21608 (N_21608,N_18067,N_17989);
nand U21609 (N_21609,N_18997,N_18024);
nand U21610 (N_21610,N_17896,N_18730);
nor U21611 (N_21611,N_18822,N_18687);
or U21612 (N_21612,N_18643,N_19555);
or U21613 (N_21613,N_19368,N_19825);
or U21614 (N_21614,N_18228,N_18334);
xnor U21615 (N_21615,N_18130,N_19867);
or U21616 (N_21616,N_19300,N_19435);
nand U21617 (N_21617,N_19945,N_18605);
nor U21618 (N_21618,N_18366,N_18190);
or U21619 (N_21619,N_17572,N_19069);
or U21620 (N_21620,N_17596,N_18585);
xor U21621 (N_21621,N_17668,N_18823);
or U21622 (N_21622,N_18920,N_19036);
and U21623 (N_21623,N_19387,N_19225);
nor U21624 (N_21624,N_18340,N_18981);
and U21625 (N_21625,N_18312,N_17742);
and U21626 (N_21626,N_17627,N_18242);
xnor U21627 (N_21627,N_19942,N_19704);
xor U21628 (N_21628,N_19812,N_19987);
xor U21629 (N_21629,N_18076,N_19058);
nor U21630 (N_21630,N_19609,N_19702);
and U21631 (N_21631,N_19239,N_18695);
and U21632 (N_21632,N_19848,N_18869);
and U21633 (N_21633,N_17591,N_19912);
xor U21634 (N_21634,N_19475,N_18636);
or U21635 (N_21635,N_19162,N_19164);
nor U21636 (N_21636,N_17889,N_17714);
nand U21637 (N_21637,N_19977,N_18375);
and U21638 (N_21638,N_18748,N_18379);
nor U21639 (N_21639,N_18196,N_17590);
nor U21640 (N_21640,N_19897,N_17700);
and U21641 (N_21641,N_18682,N_17517);
and U21642 (N_21642,N_19692,N_19393);
xnor U21643 (N_21643,N_17947,N_18635);
and U21644 (N_21644,N_18493,N_18916);
and U21645 (N_21645,N_19675,N_18251);
nand U21646 (N_21646,N_19277,N_19416);
xor U21647 (N_21647,N_19817,N_19158);
or U21648 (N_21648,N_18402,N_19048);
or U21649 (N_21649,N_19308,N_19459);
xnor U21650 (N_21650,N_18432,N_17909);
xnor U21651 (N_21651,N_19982,N_18104);
xor U21652 (N_21652,N_18910,N_17629);
nor U21653 (N_21653,N_18528,N_17564);
nand U21654 (N_21654,N_18979,N_19088);
nand U21655 (N_21655,N_18646,N_19423);
and U21656 (N_21656,N_18945,N_19407);
xnor U21657 (N_21657,N_19167,N_19302);
or U21658 (N_21658,N_19257,N_19475);
nor U21659 (N_21659,N_19382,N_19213);
nand U21660 (N_21660,N_19547,N_18710);
or U21661 (N_21661,N_19004,N_18250);
and U21662 (N_21662,N_17644,N_18653);
or U21663 (N_21663,N_17578,N_18200);
nand U21664 (N_21664,N_18114,N_18309);
or U21665 (N_21665,N_19084,N_19371);
xnor U21666 (N_21666,N_19808,N_17676);
and U21667 (N_21667,N_19391,N_19323);
xnor U21668 (N_21668,N_19273,N_17997);
nor U21669 (N_21669,N_19667,N_18536);
nor U21670 (N_21670,N_18692,N_17877);
and U21671 (N_21671,N_19029,N_19598);
nand U21672 (N_21672,N_19200,N_18145);
or U21673 (N_21673,N_17747,N_17766);
nor U21674 (N_21674,N_18780,N_19202);
or U21675 (N_21675,N_19416,N_18599);
nand U21676 (N_21676,N_19734,N_19292);
nor U21677 (N_21677,N_18881,N_17927);
xnor U21678 (N_21678,N_19109,N_19479);
nand U21679 (N_21679,N_17663,N_18898);
nor U21680 (N_21680,N_18806,N_19827);
nor U21681 (N_21681,N_18544,N_17682);
or U21682 (N_21682,N_17938,N_18140);
or U21683 (N_21683,N_19830,N_19203);
xor U21684 (N_21684,N_18319,N_17869);
and U21685 (N_21685,N_18409,N_18912);
xnor U21686 (N_21686,N_17816,N_17644);
nor U21687 (N_21687,N_17854,N_17679);
nor U21688 (N_21688,N_17856,N_19647);
and U21689 (N_21689,N_17884,N_18255);
xnor U21690 (N_21690,N_18810,N_19211);
xnor U21691 (N_21691,N_17769,N_17856);
nand U21692 (N_21692,N_18066,N_18104);
nand U21693 (N_21693,N_19680,N_19816);
and U21694 (N_21694,N_18108,N_18589);
and U21695 (N_21695,N_18199,N_19903);
or U21696 (N_21696,N_18936,N_19645);
nor U21697 (N_21697,N_18345,N_19804);
and U21698 (N_21698,N_18081,N_19248);
nand U21699 (N_21699,N_18618,N_19530);
nor U21700 (N_21700,N_19035,N_19795);
nand U21701 (N_21701,N_19114,N_18158);
nor U21702 (N_21702,N_18429,N_17570);
or U21703 (N_21703,N_19235,N_18446);
and U21704 (N_21704,N_19112,N_19238);
xnor U21705 (N_21705,N_18574,N_18291);
nand U21706 (N_21706,N_19896,N_18092);
nor U21707 (N_21707,N_18437,N_19434);
nand U21708 (N_21708,N_19232,N_19956);
or U21709 (N_21709,N_19563,N_18251);
nand U21710 (N_21710,N_18892,N_19374);
and U21711 (N_21711,N_19065,N_18543);
and U21712 (N_21712,N_19413,N_18622);
xor U21713 (N_21713,N_19635,N_17737);
xor U21714 (N_21714,N_18088,N_19899);
nor U21715 (N_21715,N_18150,N_19861);
nand U21716 (N_21716,N_18945,N_19581);
or U21717 (N_21717,N_17952,N_17763);
xor U21718 (N_21718,N_19717,N_19285);
nor U21719 (N_21719,N_18474,N_17521);
or U21720 (N_21720,N_18393,N_19371);
nand U21721 (N_21721,N_17639,N_19400);
nand U21722 (N_21722,N_17960,N_18452);
nand U21723 (N_21723,N_19978,N_19785);
or U21724 (N_21724,N_18016,N_17582);
and U21725 (N_21725,N_17720,N_18171);
and U21726 (N_21726,N_18960,N_18846);
and U21727 (N_21727,N_17846,N_18004);
nand U21728 (N_21728,N_19647,N_19431);
xnor U21729 (N_21729,N_19816,N_17521);
or U21730 (N_21730,N_18781,N_19541);
nand U21731 (N_21731,N_18400,N_18496);
nand U21732 (N_21732,N_18559,N_18259);
nand U21733 (N_21733,N_19825,N_17803);
nor U21734 (N_21734,N_19981,N_18507);
xor U21735 (N_21735,N_19373,N_18968);
or U21736 (N_21736,N_19112,N_18084);
or U21737 (N_21737,N_18694,N_18101);
or U21738 (N_21738,N_18435,N_18741);
nand U21739 (N_21739,N_19776,N_17902);
nor U21740 (N_21740,N_17588,N_18602);
xor U21741 (N_21741,N_19789,N_17893);
nand U21742 (N_21742,N_18917,N_18102);
xor U21743 (N_21743,N_19500,N_18376);
and U21744 (N_21744,N_19879,N_17847);
nand U21745 (N_21745,N_18714,N_17594);
and U21746 (N_21746,N_17863,N_18091);
and U21747 (N_21747,N_19799,N_17773);
nand U21748 (N_21748,N_19603,N_19179);
and U21749 (N_21749,N_17920,N_18397);
and U21750 (N_21750,N_18827,N_19521);
or U21751 (N_21751,N_18054,N_18695);
or U21752 (N_21752,N_18802,N_18292);
xnor U21753 (N_21753,N_17540,N_18407);
nor U21754 (N_21754,N_18359,N_18033);
and U21755 (N_21755,N_18443,N_17565);
nor U21756 (N_21756,N_19141,N_19718);
and U21757 (N_21757,N_17859,N_19866);
nor U21758 (N_21758,N_18734,N_19243);
and U21759 (N_21759,N_17526,N_19839);
and U21760 (N_21760,N_17796,N_19024);
and U21761 (N_21761,N_18035,N_18871);
or U21762 (N_21762,N_19037,N_17744);
and U21763 (N_21763,N_19043,N_19596);
nand U21764 (N_21764,N_18847,N_18350);
xor U21765 (N_21765,N_18458,N_18565);
and U21766 (N_21766,N_18691,N_19134);
or U21767 (N_21767,N_19962,N_18395);
xnor U21768 (N_21768,N_19436,N_19915);
nand U21769 (N_21769,N_19250,N_18168);
xnor U21770 (N_21770,N_19587,N_19846);
nand U21771 (N_21771,N_18536,N_18002);
or U21772 (N_21772,N_18113,N_18001);
xor U21773 (N_21773,N_17907,N_19324);
xnor U21774 (N_21774,N_19489,N_18183);
nand U21775 (N_21775,N_19479,N_18167);
or U21776 (N_21776,N_19957,N_19164);
or U21777 (N_21777,N_19499,N_19702);
or U21778 (N_21778,N_18388,N_19472);
nor U21779 (N_21779,N_19274,N_19967);
nand U21780 (N_21780,N_19803,N_17608);
xor U21781 (N_21781,N_19170,N_19581);
or U21782 (N_21782,N_18228,N_17934);
nand U21783 (N_21783,N_17657,N_18537);
and U21784 (N_21784,N_17779,N_18961);
nand U21785 (N_21785,N_17861,N_19612);
and U21786 (N_21786,N_19400,N_18514);
or U21787 (N_21787,N_19687,N_17528);
nand U21788 (N_21788,N_18819,N_19111);
xor U21789 (N_21789,N_19520,N_17616);
xor U21790 (N_21790,N_18995,N_19922);
nand U21791 (N_21791,N_17781,N_19851);
or U21792 (N_21792,N_19105,N_17671);
nor U21793 (N_21793,N_19133,N_18621);
or U21794 (N_21794,N_18617,N_18219);
or U21795 (N_21795,N_18841,N_18299);
nor U21796 (N_21796,N_19712,N_18978);
xnor U21797 (N_21797,N_19076,N_19701);
and U21798 (N_21798,N_17766,N_18776);
or U21799 (N_21799,N_19749,N_18688);
or U21800 (N_21800,N_19253,N_17707);
nand U21801 (N_21801,N_19850,N_18821);
nand U21802 (N_21802,N_19128,N_17655);
and U21803 (N_21803,N_17815,N_19335);
nand U21804 (N_21804,N_18994,N_18266);
xor U21805 (N_21805,N_18843,N_19144);
and U21806 (N_21806,N_19580,N_18710);
and U21807 (N_21807,N_18647,N_19738);
nor U21808 (N_21808,N_17581,N_19786);
and U21809 (N_21809,N_19461,N_17766);
xor U21810 (N_21810,N_19893,N_19354);
or U21811 (N_21811,N_18178,N_17746);
or U21812 (N_21812,N_18666,N_19139);
xnor U21813 (N_21813,N_18157,N_17668);
nand U21814 (N_21814,N_18995,N_17830);
nor U21815 (N_21815,N_17506,N_18977);
or U21816 (N_21816,N_18981,N_18887);
nand U21817 (N_21817,N_19570,N_17833);
and U21818 (N_21818,N_19220,N_18190);
xnor U21819 (N_21819,N_19833,N_19775);
or U21820 (N_21820,N_17572,N_18827);
xnor U21821 (N_21821,N_17872,N_17873);
and U21822 (N_21822,N_19813,N_19908);
and U21823 (N_21823,N_19620,N_17680);
nand U21824 (N_21824,N_17531,N_19224);
xor U21825 (N_21825,N_17998,N_18437);
and U21826 (N_21826,N_17886,N_17723);
nand U21827 (N_21827,N_18029,N_17627);
and U21828 (N_21828,N_19556,N_18413);
xor U21829 (N_21829,N_19250,N_18753);
nand U21830 (N_21830,N_18153,N_17949);
nand U21831 (N_21831,N_18843,N_18932);
or U21832 (N_21832,N_18410,N_17841);
xor U21833 (N_21833,N_19706,N_17881);
nor U21834 (N_21834,N_18593,N_19170);
and U21835 (N_21835,N_19247,N_18709);
xor U21836 (N_21836,N_18502,N_17667);
xor U21837 (N_21837,N_18770,N_17916);
and U21838 (N_21838,N_18215,N_19954);
xnor U21839 (N_21839,N_17601,N_18708);
nor U21840 (N_21840,N_18829,N_18404);
nor U21841 (N_21841,N_17554,N_18061);
nor U21842 (N_21842,N_17648,N_19790);
or U21843 (N_21843,N_19670,N_19507);
and U21844 (N_21844,N_18414,N_19610);
xnor U21845 (N_21845,N_19359,N_18353);
or U21846 (N_21846,N_17770,N_19803);
or U21847 (N_21847,N_17592,N_19659);
nand U21848 (N_21848,N_19597,N_19416);
xor U21849 (N_21849,N_18534,N_18258);
nor U21850 (N_21850,N_18941,N_18581);
nor U21851 (N_21851,N_18099,N_17790);
and U21852 (N_21852,N_19834,N_19404);
or U21853 (N_21853,N_19061,N_19454);
or U21854 (N_21854,N_18734,N_18621);
or U21855 (N_21855,N_18578,N_17856);
nand U21856 (N_21856,N_18023,N_19855);
and U21857 (N_21857,N_17953,N_19389);
nand U21858 (N_21858,N_18734,N_19919);
nand U21859 (N_21859,N_17503,N_18824);
or U21860 (N_21860,N_18292,N_18523);
and U21861 (N_21861,N_18698,N_18866);
or U21862 (N_21862,N_19419,N_18871);
xnor U21863 (N_21863,N_18983,N_18002);
xnor U21864 (N_21864,N_18384,N_19234);
nor U21865 (N_21865,N_18503,N_17835);
and U21866 (N_21866,N_19577,N_17546);
nand U21867 (N_21867,N_18967,N_17802);
nand U21868 (N_21868,N_18860,N_18382);
or U21869 (N_21869,N_18605,N_17852);
xor U21870 (N_21870,N_19198,N_19201);
nand U21871 (N_21871,N_17600,N_18591);
nor U21872 (N_21872,N_19184,N_18282);
and U21873 (N_21873,N_19073,N_19477);
xor U21874 (N_21874,N_19564,N_18114);
xnor U21875 (N_21875,N_17617,N_19814);
nand U21876 (N_21876,N_18373,N_18015);
nand U21877 (N_21877,N_19462,N_17605);
nor U21878 (N_21878,N_17786,N_17794);
xnor U21879 (N_21879,N_18849,N_19172);
nor U21880 (N_21880,N_18326,N_19733);
and U21881 (N_21881,N_18920,N_18956);
nor U21882 (N_21882,N_18635,N_19117);
nand U21883 (N_21883,N_19286,N_18909);
or U21884 (N_21884,N_19367,N_17861);
or U21885 (N_21885,N_19827,N_19412);
nand U21886 (N_21886,N_17826,N_17687);
xnor U21887 (N_21887,N_18666,N_17905);
or U21888 (N_21888,N_19554,N_18445);
or U21889 (N_21889,N_18141,N_17618);
and U21890 (N_21890,N_19136,N_17859);
or U21891 (N_21891,N_18764,N_17793);
or U21892 (N_21892,N_19480,N_17908);
nor U21893 (N_21893,N_18627,N_18526);
nand U21894 (N_21894,N_17993,N_18178);
and U21895 (N_21895,N_18830,N_19223);
nand U21896 (N_21896,N_18593,N_19335);
and U21897 (N_21897,N_18270,N_18273);
xor U21898 (N_21898,N_18165,N_18308);
xor U21899 (N_21899,N_19680,N_18406);
nand U21900 (N_21900,N_18817,N_18008);
nand U21901 (N_21901,N_17634,N_17652);
or U21902 (N_21902,N_19521,N_18783);
nand U21903 (N_21903,N_18148,N_18650);
nor U21904 (N_21904,N_18487,N_18989);
and U21905 (N_21905,N_18476,N_19346);
or U21906 (N_21906,N_18312,N_18167);
xor U21907 (N_21907,N_19521,N_19420);
and U21908 (N_21908,N_19189,N_19175);
and U21909 (N_21909,N_17629,N_18784);
nand U21910 (N_21910,N_19007,N_18928);
and U21911 (N_21911,N_18101,N_18742);
or U21912 (N_21912,N_18834,N_19664);
nor U21913 (N_21913,N_18969,N_17621);
xor U21914 (N_21914,N_19441,N_17690);
xor U21915 (N_21915,N_19386,N_19032);
or U21916 (N_21916,N_18282,N_17732);
nor U21917 (N_21917,N_19866,N_19062);
nand U21918 (N_21918,N_18417,N_17598);
nand U21919 (N_21919,N_19073,N_19232);
nand U21920 (N_21920,N_18811,N_17872);
nand U21921 (N_21921,N_18574,N_17500);
nand U21922 (N_21922,N_17825,N_17513);
nor U21923 (N_21923,N_18546,N_19101);
and U21924 (N_21924,N_18646,N_19730);
nor U21925 (N_21925,N_18356,N_19649);
nor U21926 (N_21926,N_17512,N_19950);
xnor U21927 (N_21927,N_17746,N_18719);
and U21928 (N_21928,N_18665,N_19435);
xnor U21929 (N_21929,N_18419,N_17889);
nor U21930 (N_21930,N_19367,N_18143);
nand U21931 (N_21931,N_18343,N_19056);
and U21932 (N_21932,N_18332,N_19259);
nand U21933 (N_21933,N_19215,N_18854);
xor U21934 (N_21934,N_19212,N_19389);
nand U21935 (N_21935,N_18698,N_18271);
nor U21936 (N_21936,N_18880,N_18580);
nand U21937 (N_21937,N_19021,N_17749);
nand U21938 (N_21938,N_19466,N_17748);
nor U21939 (N_21939,N_19569,N_17677);
or U21940 (N_21940,N_19028,N_17546);
and U21941 (N_21941,N_18372,N_18672);
nor U21942 (N_21942,N_18838,N_18002);
and U21943 (N_21943,N_19421,N_17972);
or U21944 (N_21944,N_18516,N_18166);
nor U21945 (N_21945,N_18327,N_19514);
nand U21946 (N_21946,N_18855,N_19023);
nand U21947 (N_21947,N_17867,N_19027);
nand U21948 (N_21948,N_19084,N_18534);
xnor U21949 (N_21949,N_18066,N_19845);
nor U21950 (N_21950,N_19074,N_18757);
xnor U21951 (N_21951,N_19053,N_18137);
and U21952 (N_21952,N_19091,N_17949);
xnor U21953 (N_21953,N_18726,N_18197);
nor U21954 (N_21954,N_17666,N_17941);
xor U21955 (N_21955,N_17553,N_18062);
nor U21956 (N_21956,N_18564,N_17962);
nor U21957 (N_21957,N_18548,N_18882);
nor U21958 (N_21958,N_17721,N_18203);
xnor U21959 (N_21959,N_18589,N_19755);
xor U21960 (N_21960,N_19973,N_17789);
nor U21961 (N_21961,N_19621,N_19489);
or U21962 (N_21962,N_17995,N_19017);
xor U21963 (N_21963,N_18427,N_19391);
xnor U21964 (N_21964,N_18129,N_18355);
nand U21965 (N_21965,N_18143,N_18865);
nand U21966 (N_21966,N_17578,N_19373);
nor U21967 (N_21967,N_19864,N_18376);
nand U21968 (N_21968,N_18938,N_19313);
nor U21969 (N_21969,N_19050,N_18961);
xor U21970 (N_21970,N_17743,N_18061);
and U21971 (N_21971,N_18024,N_19954);
xor U21972 (N_21972,N_19164,N_19613);
nor U21973 (N_21973,N_19440,N_18103);
or U21974 (N_21974,N_18192,N_18260);
nand U21975 (N_21975,N_19707,N_19406);
or U21976 (N_21976,N_19691,N_18902);
or U21977 (N_21977,N_19496,N_18296);
nor U21978 (N_21978,N_18051,N_17639);
nand U21979 (N_21979,N_17798,N_17817);
nor U21980 (N_21980,N_18711,N_18440);
xor U21981 (N_21981,N_19800,N_19160);
nand U21982 (N_21982,N_19140,N_18756);
nand U21983 (N_21983,N_19229,N_18692);
and U21984 (N_21984,N_19233,N_19275);
nor U21985 (N_21985,N_19954,N_19604);
and U21986 (N_21986,N_19471,N_18164);
nor U21987 (N_21987,N_18647,N_19482);
nor U21988 (N_21988,N_18965,N_18541);
nand U21989 (N_21989,N_19883,N_19604);
xnor U21990 (N_21990,N_18618,N_19388);
or U21991 (N_21991,N_17711,N_19688);
nor U21992 (N_21992,N_19923,N_17820);
nor U21993 (N_21993,N_17858,N_18850);
or U21994 (N_21994,N_17748,N_18571);
or U21995 (N_21995,N_19547,N_19243);
and U21996 (N_21996,N_17965,N_17747);
xnor U21997 (N_21997,N_18610,N_17966);
nor U21998 (N_21998,N_19005,N_17566);
nand U21999 (N_21999,N_19892,N_18916);
xor U22000 (N_22000,N_17571,N_19522);
and U22001 (N_22001,N_17877,N_17978);
or U22002 (N_22002,N_18488,N_18711);
nand U22003 (N_22003,N_17509,N_19049);
nor U22004 (N_22004,N_19008,N_19958);
nor U22005 (N_22005,N_19907,N_17923);
nor U22006 (N_22006,N_17984,N_19836);
or U22007 (N_22007,N_18093,N_17969);
nor U22008 (N_22008,N_19994,N_18694);
xnor U22009 (N_22009,N_19097,N_18207);
xnor U22010 (N_22010,N_19422,N_18529);
and U22011 (N_22011,N_18517,N_18783);
xor U22012 (N_22012,N_19916,N_18427);
xnor U22013 (N_22013,N_19827,N_19899);
or U22014 (N_22014,N_18566,N_17688);
or U22015 (N_22015,N_18050,N_19857);
nand U22016 (N_22016,N_19161,N_18768);
nand U22017 (N_22017,N_19843,N_18724);
xnor U22018 (N_22018,N_19531,N_18591);
xor U22019 (N_22019,N_18822,N_19970);
and U22020 (N_22020,N_18391,N_18316);
nor U22021 (N_22021,N_19624,N_19046);
and U22022 (N_22022,N_19465,N_17575);
nand U22023 (N_22023,N_19427,N_19309);
or U22024 (N_22024,N_19453,N_18823);
xnor U22025 (N_22025,N_17530,N_19499);
xnor U22026 (N_22026,N_19080,N_17834);
xnor U22027 (N_22027,N_18865,N_17775);
nor U22028 (N_22028,N_19390,N_19476);
xnor U22029 (N_22029,N_19014,N_19286);
xor U22030 (N_22030,N_18878,N_18401);
and U22031 (N_22031,N_17512,N_17508);
and U22032 (N_22032,N_19908,N_19416);
nand U22033 (N_22033,N_18879,N_17549);
nand U22034 (N_22034,N_18791,N_18718);
nand U22035 (N_22035,N_19950,N_19241);
or U22036 (N_22036,N_19219,N_18956);
and U22037 (N_22037,N_17757,N_19584);
xor U22038 (N_22038,N_18567,N_19638);
xor U22039 (N_22039,N_17629,N_18168);
nand U22040 (N_22040,N_17793,N_19635);
and U22041 (N_22041,N_18838,N_17578);
nor U22042 (N_22042,N_17579,N_19325);
nor U22043 (N_22043,N_19192,N_18770);
or U22044 (N_22044,N_18205,N_18441);
nand U22045 (N_22045,N_18550,N_17889);
nand U22046 (N_22046,N_18985,N_18668);
xnor U22047 (N_22047,N_18111,N_19593);
and U22048 (N_22048,N_19654,N_19168);
nand U22049 (N_22049,N_19119,N_17556);
or U22050 (N_22050,N_19301,N_19819);
nand U22051 (N_22051,N_19938,N_17631);
xor U22052 (N_22052,N_18826,N_17843);
nand U22053 (N_22053,N_18002,N_19071);
nand U22054 (N_22054,N_19491,N_17603);
xor U22055 (N_22055,N_17885,N_17829);
xnor U22056 (N_22056,N_18908,N_19445);
nor U22057 (N_22057,N_19628,N_18254);
or U22058 (N_22058,N_19579,N_18225);
xor U22059 (N_22059,N_19672,N_17639);
nor U22060 (N_22060,N_17607,N_17790);
and U22061 (N_22061,N_17809,N_19576);
nand U22062 (N_22062,N_19034,N_19011);
xor U22063 (N_22063,N_19226,N_19687);
nor U22064 (N_22064,N_19450,N_18551);
nor U22065 (N_22065,N_19653,N_17997);
xnor U22066 (N_22066,N_19473,N_18151);
or U22067 (N_22067,N_19627,N_17681);
nor U22068 (N_22068,N_18787,N_19941);
nand U22069 (N_22069,N_18974,N_17515);
xor U22070 (N_22070,N_18438,N_19564);
and U22071 (N_22071,N_17669,N_19153);
nor U22072 (N_22072,N_17701,N_18675);
xor U22073 (N_22073,N_18270,N_19474);
xnor U22074 (N_22074,N_17625,N_17672);
and U22075 (N_22075,N_19713,N_17632);
nand U22076 (N_22076,N_19839,N_18458);
and U22077 (N_22077,N_18384,N_18663);
nand U22078 (N_22078,N_19787,N_19577);
or U22079 (N_22079,N_19544,N_18945);
nor U22080 (N_22080,N_18588,N_17788);
and U22081 (N_22081,N_19893,N_18291);
or U22082 (N_22082,N_18861,N_18152);
xnor U22083 (N_22083,N_17899,N_18064);
nor U22084 (N_22084,N_18693,N_17681);
or U22085 (N_22085,N_19982,N_18944);
nand U22086 (N_22086,N_18766,N_18410);
nand U22087 (N_22087,N_18323,N_18781);
xor U22088 (N_22088,N_17984,N_18454);
nand U22089 (N_22089,N_17786,N_18568);
xor U22090 (N_22090,N_19142,N_19097);
xnor U22091 (N_22091,N_17868,N_18253);
and U22092 (N_22092,N_19323,N_19507);
xor U22093 (N_22093,N_18255,N_17907);
xnor U22094 (N_22094,N_18102,N_18415);
or U22095 (N_22095,N_17583,N_17670);
nand U22096 (N_22096,N_18070,N_18502);
nand U22097 (N_22097,N_18011,N_17890);
or U22098 (N_22098,N_18780,N_18518);
nand U22099 (N_22099,N_17954,N_18800);
or U22100 (N_22100,N_18691,N_17951);
or U22101 (N_22101,N_17546,N_18178);
nor U22102 (N_22102,N_18759,N_18314);
nor U22103 (N_22103,N_19834,N_19009);
and U22104 (N_22104,N_18118,N_17778);
nor U22105 (N_22105,N_18457,N_18875);
or U22106 (N_22106,N_19051,N_17571);
nand U22107 (N_22107,N_19489,N_17532);
nand U22108 (N_22108,N_18295,N_18422);
nand U22109 (N_22109,N_19188,N_19178);
or U22110 (N_22110,N_18042,N_18266);
nor U22111 (N_22111,N_18188,N_19174);
nand U22112 (N_22112,N_18275,N_19105);
nor U22113 (N_22113,N_17798,N_17847);
nand U22114 (N_22114,N_18801,N_17775);
and U22115 (N_22115,N_19111,N_18615);
and U22116 (N_22116,N_17761,N_19035);
nor U22117 (N_22117,N_19558,N_19976);
or U22118 (N_22118,N_19068,N_18618);
xor U22119 (N_22119,N_18936,N_18254);
nor U22120 (N_22120,N_18347,N_18315);
and U22121 (N_22121,N_18726,N_18386);
xnor U22122 (N_22122,N_19164,N_19842);
nand U22123 (N_22123,N_18356,N_18508);
xor U22124 (N_22124,N_18610,N_18456);
nand U22125 (N_22125,N_17593,N_19916);
and U22126 (N_22126,N_19016,N_17520);
nand U22127 (N_22127,N_17522,N_19373);
and U22128 (N_22128,N_18413,N_18273);
nand U22129 (N_22129,N_18719,N_18783);
and U22130 (N_22130,N_18471,N_19945);
and U22131 (N_22131,N_18314,N_19179);
xnor U22132 (N_22132,N_18453,N_18635);
nor U22133 (N_22133,N_17656,N_18714);
and U22134 (N_22134,N_19377,N_19083);
nor U22135 (N_22135,N_18782,N_17943);
nor U22136 (N_22136,N_18231,N_18370);
or U22137 (N_22137,N_18318,N_18309);
or U22138 (N_22138,N_18155,N_19232);
nor U22139 (N_22139,N_19123,N_18630);
nand U22140 (N_22140,N_19618,N_18485);
or U22141 (N_22141,N_18142,N_19210);
and U22142 (N_22142,N_17826,N_18905);
or U22143 (N_22143,N_17835,N_18720);
xnor U22144 (N_22144,N_18245,N_19112);
and U22145 (N_22145,N_19748,N_18181);
and U22146 (N_22146,N_19880,N_19755);
nor U22147 (N_22147,N_18206,N_18293);
nand U22148 (N_22148,N_19807,N_18325);
nor U22149 (N_22149,N_17972,N_18874);
nor U22150 (N_22150,N_18033,N_19722);
or U22151 (N_22151,N_18348,N_18801);
nor U22152 (N_22152,N_19513,N_18958);
nand U22153 (N_22153,N_19352,N_19423);
nand U22154 (N_22154,N_19171,N_18601);
xnor U22155 (N_22155,N_19000,N_17670);
nor U22156 (N_22156,N_18113,N_19750);
nor U22157 (N_22157,N_18775,N_18007);
nor U22158 (N_22158,N_19055,N_18123);
and U22159 (N_22159,N_18979,N_19383);
and U22160 (N_22160,N_19478,N_17524);
nand U22161 (N_22161,N_17513,N_17986);
nand U22162 (N_22162,N_19020,N_19817);
or U22163 (N_22163,N_17566,N_17678);
and U22164 (N_22164,N_17577,N_18655);
xor U22165 (N_22165,N_18766,N_17797);
nor U22166 (N_22166,N_17844,N_19677);
or U22167 (N_22167,N_18413,N_18628);
xnor U22168 (N_22168,N_19822,N_18005);
or U22169 (N_22169,N_18002,N_19591);
nand U22170 (N_22170,N_18409,N_19571);
or U22171 (N_22171,N_18873,N_17548);
nor U22172 (N_22172,N_19232,N_18225);
or U22173 (N_22173,N_18911,N_19220);
nand U22174 (N_22174,N_17968,N_18126);
xnor U22175 (N_22175,N_18611,N_17989);
or U22176 (N_22176,N_19420,N_17776);
and U22177 (N_22177,N_18712,N_18942);
and U22178 (N_22178,N_18039,N_18880);
and U22179 (N_22179,N_18481,N_19856);
and U22180 (N_22180,N_19192,N_19055);
nand U22181 (N_22181,N_18157,N_17827);
xor U22182 (N_22182,N_18869,N_17995);
and U22183 (N_22183,N_17764,N_18402);
xor U22184 (N_22184,N_18534,N_18019);
and U22185 (N_22185,N_19853,N_17662);
or U22186 (N_22186,N_19287,N_19852);
xor U22187 (N_22187,N_18106,N_19286);
nand U22188 (N_22188,N_17607,N_18323);
nand U22189 (N_22189,N_19328,N_19473);
nor U22190 (N_22190,N_19505,N_19720);
or U22191 (N_22191,N_17683,N_18024);
and U22192 (N_22192,N_19916,N_19641);
or U22193 (N_22193,N_18945,N_17925);
nor U22194 (N_22194,N_19423,N_18036);
or U22195 (N_22195,N_19409,N_19895);
and U22196 (N_22196,N_18186,N_18452);
xnor U22197 (N_22197,N_18119,N_18046);
nor U22198 (N_22198,N_18685,N_18243);
nand U22199 (N_22199,N_17953,N_18793);
or U22200 (N_22200,N_17848,N_19654);
and U22201 (N_22201,N_18438,N_19889);
and U22202 (N_22202,N_19960,N_19710);
nor U22203 (N_22203,N_18578,N_18386);
xor U22204 (N_22204,N_18709,N_19533);
xor U22205 (N_22205,N_18692,N_19444);
nand U22206 (N_22206,N_18437,N_18562);
or U22207 (N_22207,N_18428,N_18595);
xnor U22208 (N_22208,N_19845,N_18946);
or U22209 (N_22209,N_19931,N_19830);
or U22210 (N_22210,N_18639,N_18302);
or U22211 (N_22211,N_19516,N_18955);
xnor U22212 (N_22212,N_19601,N_17651);
nor U22213 (N_22213,N_18756,N_18631);
nand U22214 (N_22214,N_18383,N_17518);
and U22215 (N_22215,N_19647,N_19862);
nand U22216 (N_22216,N_18432,N_19743);
xor U22217 (N_22217,N_19994,N_19443);
xnor U22218 (N_22218,N_19785,N_17945);
and U22219 (N_22219,N_18504,N_18431);
nand U22220 (N_22220,N_18990,N_18907);
nand U22221 (N_22221,N_18238,N_17835);
or U22222 (N_22222,N_18643,N_18075);
xnor U22223 (N_22223,N_18574,N_17796);
xnor U22224 (N_22224,N_19039,N_19675);
and U22225 (N_22225,N_18679,N_19949);
nor U22226 (N_22226,N_19278,N_18492);
and U22227 (N_22227,N_19963,N_19504);
nor U22228 (N_22228,N_18389,N_18972);
and U22229 (N_22229,N_18403,N_18809);
or U22230 (N_22230,N_17776,N_19935);
xnor U22231 (N_22231,N_19137,N_18099);
nand U22232 (N_22232,N_17918,N_17674);
or U22233 (N_22233,N_19758,N_18162);
nand U22234 (N_22234,N_19929,N_19811);
nand U22235 (N_22235,N_17787,N_19305);
or U22236 (N_22236,N_18360,N_19631);
or U22237 (N_22237,N_18715,N_19172);
nor U22238 (N_22238,N_17978,N_17836);
xor U22239 (N_22239,N_18380,N_19665);
xor U22240 (N_22240,N_18584,N_19808);
and U22241 (N_22241,N_19638,N_17949);
nand U22242 (N_22242,N_18305,N_18015);
and U22243 (N_22243,N_18880,N_18892);
nor U22244 (N_22244,N_19608,N_18790);
and U22245 (N_22245,N_18465,N_18271);
nor U22246 (N_22246,N_19916,N_19844);
or U22247 (N_22247,N_17708,N_18768);
nor U22248 (N_22248,N_18418,N_18990);
nand U22249 (N_22249,N_19871,N_18397);
nor U22250 (N_22250,N_18647,N_19680);
nand U22251 (N_22251,N_18736,N_17602);
or U22252 (N_22252,N_19160,N_19275);
xor U22253 (N_22253,N_17626,N_18408);
and U22254 (N_22254,N_19893,N_19327);
and U22255 (N_22255,N_19281,N_18131);
xor U22256 (N_22256,N_17976,N_19886);
nor U22257 (N_22257,N_19944,N_17818);
or U22258 (N_22258,N_18886,N_19761);
nor U22259 (N_22259,N_18241,N_18302);
or U22260 (N_22260,N_19465,N_19326);
or U22261 (N_22261,N_18737,N_19255);
or U22262 (N_22262,N_19273,N_18084);
or U22263 (N_22263,N_18891,N_17861);
xnor U22264 (N_22264,N_17603,N_19237);
or U22265 (N_22265,N_18329,N_19198);
nand U22266 (N_22266,N_18880,N_18890);
nor U22267 (N_22267,N_17748,N_19246);
and U22268 (N_22268,N_19197,N_18228);
nor U22269 (N_22269,N_19885,N_18614);
nand U22270 (N_22270,N_19502,N_18697);
nand U22271 (N_22271,N_17629,N_17603);
nand U22272 (N_22272,N_18794,N_19271);
xnor U22273 (N_22273,N_19284,N_18331);
xor U22274 (N_22274,N_19764,N_19945);
and U22275 (N_22275,N_19628,N_19116);
xnor U22276 (N_22276,N_19469,N_17772);
or U22277 (N_22277,N_19318,N_19617);
nand U22278 (N_22278,N_17632,N_18269);
nand U22279 (N_22279,N_19259,N_19934);
nor U22280 (N_22280,N_18392,N_18041);
xnor U22281 (N_22281,N_18812,N_18366);
or U22282 (N_22282,N_18430,N_18120);
nand U22283 (N_22283,N_18043,N_19316);
and U22284 (N_22284,N_18802,N_18820);
nand U22285 (N_22285,N_19825,N_19753);
and U22286 (N_22286,N_19774,N_18026);
nor U22287 (N_22287,N_19071,N_18933);
or U22288 (N_22288,N_18403,N_19495);
nor U22289 (N_22289,N_17951,N_18025);
or U22290 (N_22290,N_18561,N_19690);
nand U22291 (N_22291,N_19229,N_18278);
or U22292 (N_22292,N_18096,N_18421);
or U22293 (N_22293,N_19366,N_17663);
and U22294 (N_22294,N_19978,N_18082);
xor U22295 (N_22295,N_19911,N_19924);
xor U22296 (N_22296,N_19888,N_19605);
nand U22297 (N_22297,N_18706,N_19173);
or U22298 (N_22298,N_19834,N_19395);
nor U22299 (N_22299,N_19105,N_17971);
nand U22300 (N_22300,N_18029,N_19448);
or U22301 (N_22301,N_17701,N_19398);
or U22302 (N_22302,N_19008,N_18541);
or U22303 (N_22303,N_19570,N_18845);
xnor U22304 (N_22304,N_18483,N_18423);
and U22305 (N_22305,N_19173,N_18864);
or U22306 (N_22306,N_17819,N_18367);
or U22307 (N_22307,N_19762,N_19592);
nand U22308 (N_22308,N_18751,N_19799);
nand U22309 (N_22309,N_19439,N_19515);
nand U22310 (N_22310,N_18798,N_19126);
xnor U22311 (N_22311,N_18550,N_18777);
and U22312 (N_22312,N_19113,N_18655);
nand U22313 (N_22313,N_18419,N_18580);
xnor U22314 (N_22314,N_19225,N_18429);
or U22315 (N_22315,N_18861,N_18736);
and U22316 (N_22316,N_18395,N_19742);
nand U22317 (N_22317,N_18292,N_18393);
and U22318 (N_22318,N_18393,N_19539);
nand U22319 (N_22319,N_18785,N_19005);
xnor U22320 (N_22320,N_18130,N_19060);
and U22321 (N_22321,N_18120,N_19842);
xor U22322 (N_22322,N_18497,N_19052);
nand U22323 (N_22323,N_19179,N_18195);
nand U22324 (N_22324,N_19103,N_19622);
nor U22325 (N_22325,N_17875,N_17893);
nand U22326 (N_22326,N_19246,N_17601);
nor U22327 (N_22327,N_17797,N_17525);
nand U22328 (N_22328,N_19409,N_18576);
or U22329 (N_22329,N_19918,N_19321);
or U22330 (N_22330,N_18420,N_19983);
and U22331 (N_22331,N_19370,N_17960);
or U22332 (N_22332,N_17636,N_17620);
nand U22333 (N_22333,N_19851,N_18053);
nor U22334 (N_22334,N_19218,N_19887);
xnor U22335 (N_22335,N_17854,N_18342);
and U22336 (N_22336,N_18423,N_17518);
xnor U22337 (N_22337,N_18020,N_19174);
nor U22338 (N_22338,N_19366,N_19469);
nor U22339 (N_22339,N_18769,N_18644);
nand U22340 (N_22340,N_18399,N_18117);
or U22341 (N_22341,N_17612,N_17738);
and U22342 (N_22342,N_17817,N_19537);
xor U22343 (N_22343,N_18320,N_18713);
or U22344 (N_22344,N_17522,N_19878);
nand U22345 (N_22345,N_17996,N_17890);
and U22346 (N_22346,N_18791,N_19119);
or U22347 (N_22347,N_19763,N_17837);
nand U22348 (N_22348,N_18853,N_17702);
and U22349 (N_22349,N_19961,N_19354);
and U22350 (N_22350,N_18373,N_17747);
and U22351 (N_22351,N_18295,N_18116);
nor U22352 (N_22352,N_19483,N_19319);
nor U22353 (N_22353,N_17637,N_19881);
and U22354 (N_22354,N_19776,N_18054);
xnor U22355 (N_22355,N_19010,N_18024);
nor U22356 (N_22356,N_17510,N_19824);
nor U22357 (N_22357,N_17643,N_18876);
nor U22358 (N_22358,N_19844,N_19329);
nor U22359 (N_22359,N_18505,N_18884);
and U22360 (N_22360,N_19787,N_17623);
nand U22361 (N_22361,N_17746,N_19478);
nor U22362 (N_22362,N_19535,N_18826);
nand U22363 (N_22363,N_19327,N_17966);
and U22364 (N_22364,N_18429,N_18223);
nand U22365 (N_22365,N_19682,N_18570);
xnor U22366 (N_22366,N_18272,N_18450);
and U22367 (N_22367,N_19421,N_17755);
nand U22368 (N_22368,N_18184,N_18230);
or U22369 (N_22369,N_17576,N_17514);
xor U22370 (N_22370,N_18942,N_19644);
or U22371 (N_22371,N_17845,N_18885);
and U22372 (N_22372,N_19472,N_18815);
xor U22373 (N_22373,N_17664,N_19535);
nor U22374 (N_22374,N_19616,N_17970);
or U22375 (N_22375,N_18814,N_19853);
and U22376 (N_22376,N_19752,N_19675);
nand U22377 (N_22377,N_17701,N_18693);
nor U22378 (N_22378,N_19504,N_18459);
or U22379 (N_22379,N_17733,N_19042);
nand U22380 (N_22380,N_17683,N_18684);
and U22381 (N_22381,N_19946,N_18266);
nand U22382 (N_22382,N_19787,N_18304);
or U22383 (N_22383,N_19239,N_17536);
and U22384 (N_22384,N_19353,N_18187);
xor U22385 (N_22385,N_18547,N_19134);
or U22386 (N_22386,N_18191,N_19127);
xnor U22387 (N_22387,N_19393,N_18288);
nor U22388 (N_22388,N_17617,N_18363);
nand U22389 (N_22389,N_18396,N_19616);
nand U22390 (N_22390,N_18245,N_18687);
nor U22391 (N_22391,N_18383,N_19539);
or U22392 (N_22392,N_17618,N_19864);
nor U22393 (N_22393,N_18761,N_18088);
and U22394 (N_22394,N_18703,N_17675);
and U22395 (N_22395,N_19817,N_18581);
or U22396 (N_22396,N_18793,N_17606);
and U22397 (N_22397,N_19314,N_19548);
nand U22398 (N_22398,N_19985,N_19099);
xor U22399 (N_22399,N_18142,N_18934);
nor U22400 (N_22400,N_19366,N_18947);
and U22401 (N_22401,N_19774,N_18506);
xnor U22402 (N_22402,N_18565,N_18068);
nor U22403 (N_22403,N_19703,N_19052);
nand U22404 (N_22404,N_18467,N_17610);
or U22405 (N_22405,N_19497,N_17848);
xnor U22406 (N_22406,N_17799,N_17761);
xor U22407 (N_22407,N_19473,N_19738);
and U22408 (N_22408,N_17789,N_19636);
nor U22409 (N_22409,N_18391,N_19359);
or U22410 (N_22410,N_19969,N_19807);
nor U22411 (N_22411,N_17679,N_18631);
nand U22412 (N_22412,N_19862,N_18076);
nand U22413 (N_22413,N_18580,N_19153);
nor U22414 (N_22414,N_19168,N_18603);
nor U22415 (N_22415,N_17738,N_18688);
and U22416 (N_22416,N_17575,N_19972);
and U22417 (N_22417,N_19142,N_18672);
nor U22418 (N_22418,N_19473,N_17941);
nor U22419 (N_22419,N_19337,N_18695);
or U22420 (N_22420,N_17981,N_17684);
or U22421 (N_22421,N_19399,N_19802);
or U22422 (N_22422,N_18582,N_19908);
or U22423 (N_22423,N_18319,N_18519);
xor U22424 (N_22424,N_19124,N_19085);
and U22425 (N_22425,N_18156,N_17748);
nand U22426 (N_22426,N_18623,N_17633);
xnor U22427 (N_22427,N_18583,N_19746);
xor U22428 (N_22428,N_18803,N_18988);
xor U22429 (N_22429,N_19619,N_18721);
and U22430 (N_22430,N_18613,N_18927);
nand U22431 (N_22431,N_18804,N_19929);
and U22432 (N_22432,N_19932,N_18544);
nor U22433 (N_22433,N_18276,N_19142);
nand U22434 (N_22434,N_17978,N_18769);
xor U22435 (N_22435,N_17623,N_19272);
or U22436 (N_22436,N_17617,N_18669);
xnor U22437 (N_22437,N_19423,N_18791);
or U22438 (N_22438,N_19164,N_19716);
and U22439 (N_22439,N_18112,N_19396);
nand U22440 (N_22440,N_19224,N_18782);
or U22441 (N_22441,N_17985,N_18817);
and U22442 (N_22442,N_19230,N_17650);
nand U22443 (N_22443,N_17846,N_18738);
xnor U22444 (N_22444,N_17667,N_19193);
or U22445 (N_22445,N_19071,N_18428);
or U22446 (N_22446,N_17862,N_18997);
xor U22447 (N_22447,N_18290,N_17786);
xnor U22448 (N_22448,N_17697,N_19997);
xor U22449 (N_22449,N_17754,N_19705);
nor U22450 (N_22450,N_17871,N_18387);
xnor U22451 (N_22451,N_17812,N_18141);
xor U22452 (N_22452,N_19918,N_19567);
nor U22453 (N_22453,N_19206,N_18875);
xor U22454 (N_22454,N_19300,N_19383);
xor U22455 (N_22455,N_17562,N_17501);
or U22456 (N_22456,N_18504,N_19071);
nor U22457 (N_22457,N_18495,N_18151);
and U22458 (N_22458,N_17542,N_19168);
and U22459 (N_22459,N_18770,N_19522);
or U22460 (N_22460,N_19750,N_18052);
nand U22461 (N_22461,N_19604,N_17986);
nand U22462 (N_22462,N_18341,N_18887);
or U22463 (N_22463,N_18539,N_18712);
nor U22464 (N_22464,N_18326,N_17750);
xor U22465 (N_22465,N_19355,N_17941);
nand U22466 (N_22466,N_18439,N_18684);
nor U22467 (N_22467,N_17966,N_19615);
xor U22468 (N_22468,N_17673,N_18385);
xor U22469 (N_22469,N_17657,N_17946);
nor U22470 (N_22470,N_17924,N_18007);
and U22471 (N_22471,N_19969,N_19592);
or U22472 (N_22472,N_19137,N_19870);
and U22473 (N_22473,N_19797,N_18811);
xnor U22474 (N_22474,N_17625,N_18865);
xnor U22475 (N_22475,N_18758,N_18006);
or U22476 (N_22476,N_17884,N_19524);
nand U22477 (N_22477,N_19232,N_17570);
and U22478 (N_22478,N_17776,N_18024);
nor U22479 (N_22479,N_19241,N_19619);
xor U22480 (N_22480,N_18442,N_19484);
xor U22481 (N_22481,N_18987,N_19485);
and U22482 (N_22482,N_19498,N_19557);
xor U22483 (N_22483,N_19546,N_17748);
and U22484 (N_22484,N_17588,N_17914);
or U22485 (N_22485,N_19151,N_17986);
xnor U22486 (N_22486,N_17558,N_18213);
xnor U22487 (N_22487,N_18734,N_17768);
xnor U22488 (N_22488,N_18457,N_18622);
xor U22489 (N_22489,N_19464,N_18343);
nor U22490 (N_22490,N_18370,N_17797);
or U22491 (N_22491,N_18660,N_18938);
nand U22492 (N_22492,N_18719,N_18955);
and U22493 (N_22493,N_18430,N_19021);
and U22494 (N_22494,N_18427,N_18659);
nand U22495 (N_22495,N_18408,N_18825);
xnor U22496 (N_22496,N_18921,N_17937);
or U22497 (N_22497,N_17878,N_18585);
or U22498 (N_22498,N_19621,N_19934);
and U22499 (N_22499,N_19188,N_17897);
nand U22500 (N_22500,N_20376,N_20512);
nor U22501 (N_22501,N_21880,N_21910);
and U22502 (N_22502,N_22345,N_21932);
nor U22503 (N_22503,N_22299,N_21726);
xor U22504 (N_22504,N_20067,N_20349);
nor U22505 (N_22505,N_21897,N_20088);
xor U22506 (N_22506,N_21667,N_20078);
xor U22507 (N_22507,N_21048,N_21207);
nand U22508 (N_22508,N_20283,N_21798);
nand U22509 (N_22509,N_20487,N_21883);
xnor U22510 (N_22510,N_22424,N_21109);
nand U22511 (N_22511,N_20548,N_22004);
xor U22512 (N_22512,N_21082,N_22455);
xor U22513 (N_22513,N_21478,N_21532);
nor U22514 (N_22514,N_20143,N_20360);
and U22515 (N_22515,N_20290,N_22491);
or U22516 (N_22516,N_21878,N_20506);
xor U22517 (N_22517,N_20800,N_21855);
nor U22518 (N_22518,N_20797,N_20665);
nor U22519 (N_22519,N_21830,N_21133);
xnor U22520 (N_22520,N_21906,N_20079);
xnor U22521 (N_22521,N_21837,N_22362);
xor U22522 (N_22522,N_20835,N_21891);
or U22523 (N_22523,N_22217,N_21571);
xnor U22524 (N_22524,N_21709,N_20302);
nor U22525 (N_22525,N_21378,N_20101);
nor U22526 (N_22526,N_21523,N_21688);
xor U22527 (N_22527,N_22085,N_20920);
or U22528 (N_22528,N_21131,N_21947);
and U22529 (N_22529,N_22141,N_20123);
or U22530 (N_22530,N_21490,N_20683);
nand U22531 (N_22531,N_21093,N_20644);
xor U22532 (N_22532,N_20323,N_20267);
nor U22533 (N_22533,N_20266,N_21811);
nand U22534 (N_22534,N_21911,N_20457);
nor U22535 (N_22535,N_22021,N_20784);
or U22536 (N_22536,N_20397,N_21029);
and U22537 (N_22537,N_21994,N_22340);
nand U22538 (N_22538,N_20869,N_22445);
xor U22539 (N_22539,N_22151,N_21261);
and U22540 (N_22540,N_22118,N_22297);
nand U22541 (N_22541,N_21405,N_21442);
xnor U22542 (N_22542,N_21300,N_20870);
xor U22543 (N_22543,N_20031,N_22155);
or U22544 (N_22544,N_22153,N_22440);
nor U22545 (N_22545,N_21139,N_20113);
nand U22546 (N_22546,N_21354,N_20362);
or U22547 (N_22547,N_20825,N_20263);
nor U22548 (N_22548,N_21853,N_22460);
and U22549 (N_22549,N_21651,N_21495);
xnor U22550 (N_22550,N_21736,N_22111);
or U22551 (N_22551,N_20764,N_20697);
and U22552 (N_22552,N_21665,N_21597);
nor U22553 (N_22553,N_21999,N_20020);
xnor U22554 (N_22554,N_20517,N_21874);
or U22555 (N_22555,N_20104,N_21611);
or U22556 (N_22556,N_21307,N_20610);
xnor U22557 (N_22557,N_21987,N_20798);
xor U22558 (N_22558,N_20236,N_21330);
and U22559 (N_22559,N_20214,N_20367);
and U22560 (N_22560,N_21744,N_21190);
nand U22561 (N_22561,N_20727,N_20515);
nand U22562 (N_22562,N_20966,N_21452);
xnor U22563 (N_22563,N_21011,N_20530);
or U22564 (N_22564,N_20448,N_20698);
nor U22565 (N_22565,N_21526,N_21149);
xnor U22566 (N_22566,N_21695,N_20091);
nor U22567 (N_22567,N_20897,N_20488);
or U22568 (N_22568,N_20040,N_20299);
or U22569 (N_22569,N_21635,N_21181);
nand U22570 (N_22570,N_22385,N_20977);
or U22571 (N_22571,N_22072,N_20285);
nand U22572 (N_22572,N_22047,N_21625);
and U22573 (N_22573,N_21770,N_22376);
and U22574 (N_22574,N_22074,N_20099);
or U22575 (N_22575,N_22177,N_20243);
xor U22576 (N_22576,N_22339,N_20630);
xor U22577 (N_22577,N_20057,N_20799);
xor U22578 (N_22578,N_21958,N_20674);
nor U22579 (N_22579,N_20297,N_20444);
xnor U22580 (N_22580,N_22466,N_21989);
xnor U22581 (N_22581,N_20898,N_20199);
and U22582 (N_22582,N_21338,N_20000);
nor U22583 (N_22583,N_21374,N_21385);
and U22584 (N_22584,N_22233,N_20623);
nand U22585 (N_22585,N_22036,N_21185);
and U22586 (N_22586,N_20089,N_22066);
nand U22587 (N_22587,N_22380,N_20370);
nor U22588 (N_22588,N_21273,N_20423);
and U22589 (N_22589,N_22169,N_22022);
xor U22590 (N_22590,N_20066,N_21521);
nor U22591 (N_22591,N_21633,N_20968);
or U22592 (N_22592,N_21828,N_20436);
or U22593 (N_22593,N_20042,N_21714);
nor U22594 (N_22594,N_21324,N_22312);
or U22595 (N_22595,N_21802,N_20307);
nor U22596 (N_22596,N_20076,N_21541);
or U22597 (N_22597,N_21851,N_21650);
or U22598 (N_22598,N_20303,N_20719);
or U22599 (N_22599,N_22418,N_21603);
xor U22600 (N_22600,N_20287,N_22069);
nand U22601 (N_22601,N_20751,N_20492);
and U22602 (N_22602,N_22325,N_20760);
xor U22603 (N_22603,N_21716,N_21416);
xor U22604 (N_22604,N_22116,N_21843);
or U22605 (N_22605,N_21609,N_21247);
nand U22606 (N_22606,N_21009,N_21661);
nand U22607 (N_22607,N_22480,N_20095);
or U22608 (N_22608,N_20818,N_21809);
xnor U22609 (N_22609,N_20176,N_20442);
xnor U22610 (N_22610,N_20552,N_21923);
nor U22611 (N_22611,N_21114,N_21846);
or U22612 (N_22612,N_21964,N_21441);
nand U22613 (N_22613,N_20363,N_22368);
xnor U22614 (N_22614,N_21510,N_20980);
nand U22615 (N_22615,N_22114,N_22175);
or U22616 (N_22616,N_20958,N_21970);
xnor U22617 (N_22617,N_21220,N_21288);
nor U22618 (N_22618,N_21108,N_20007);
nand U22619 (N_22619,N_20331,N_20725);
nand U22620 (N_22620,N_20785,N_21046);
nand U22621 (N_22621,N_21540,N_21382);
or U22622 (N_22622,N_20938,N_21389);
nand U22623 (N_22623,N_21615,N_21227);
nor U22624 (N_22624,N_20445,N_20813);
nand U22625 (N_22625,N_22145,N_20246);
or U22626 (N_22626,N_22163,N_20666);
xor U22627 (N_22627,N_22484,N_22432);
or U22628 (N_22628,N_21852,N_20282);
nand U22629 (N_22629,N_21555,N_20879);
and U22630 (N_22630,N_22499,N_20860);
nand U22631 (N_22631,N_21259,N_20296);
and U22632 (N_22632,N_21723,N_20748);
xnor U22633 (N_22633,N_22434,N_21610);
xor U22634 (N_22634,N_22497,N_20269);
or U22635 (N_22635,N_21920,N_20865);
nand U22636 (N_22636,N_21805,N_20636);
xnor U22637 (N_22637,N_21125,N_22468);
xor U22638 (N_22638,N_20194,N_20841);
and U22639 (N_22639,N_20659,N_21687);
nand U22640 (N_22640,N_20171,N_22411);
or U22641 (N_22641,N_21907,N_21411);
nand U22642 (N_22642,N_20858,N_22307);
or U22643 (N_22643,N_21499,N_20153);
and U22644 (N_22644,N_21905,N_20301);
nor U22645 (N_22645,N_20461,N_22053);
xor U22646 (N_22646,N_22203,N_22355);
xnor U22647 (N_22647,N_22478,N_22238);
nand U22648 (N_22648,N_20514,N_21569);
nand U22649 (N_22649,N_21993,N_22056);
nor U22650 (N_22650,N_20503,N_22446);
xor U22651 (N_22651,N_22241,N_20223);
xnor U22652 (N_22652,N_20033,N_21545);
xnor U22653 (N_22653,N_20446,N_20563);
xor U22654 (N_22654,N_22240,N_21547);
nand U22655 (N_22655,N_21713,N_20589);
or U22656 (N_22656,N_21772,N_21895);
nor U22657 (N_22657,N_21771,N_22356);
or U22658 (N_22658,N_20775,N_20872);
xor U22659 (N_22659,N_21194,N_21360);
and U22660 (N_22660,N_20649,N_20677);
xor U22661 (N_22661,N_21289,N_20422);
nand U22662 (N_22662,N_22332,N_22413);
nand U22663 (N_22663,N_21347,N_20051);
and U22664 (N_22664,N_22398,N_21572);
or U22665 (N_22665,N_20703,N_21570);
and U22666 (N_22666,N_21038,N_20888);
or U22667 (N_22667,N_22142,N_21141);
and U22668 (N_22668,N_21636,N_22373);
xor U22669 (N_22669,N_21019,N_21000);
or U22670 (N_22670,N_21514,N_20239);
xnor U22671 (N_22671,N_20616,N_21388);
nor U22672 (N_22672,N_20689,N_22094);
nor U22673 (N_22673,N_21161,N_22442);
xor U22674 (N_22674,N_22462,N_21804);
xor U22675 (N_22675,N_22101,N_22437);
nor U22676 (N_22676,N_21395,N_20276);
or U22677 (N_22677,N_20161,N_20274);
or U22678 (N_22678,N_21335,N_20867);
and U22679 (N_22679,N_20452,N_21466);
nand U22680 (N_22680,N_22205,N_21094);
and U22681 (N_22681,N_20187,N_20516);
nor U22682 (N_22682,N_22453,N_22439);
or U22683 (N_22683,N_21949,N_21806);
and U22684 (N_22684,N_20651,N_20288);
or U22685 (N_22685,N_20310,N_22079);
xnor U22686 (N_22686,N_21642,N_20178);
and U22687 (N_22687,N_21053,N_21278);
xnor U22688 (N_22688,N_20691,N_21256);
nor U22689 (N_22689,N_20568,N_21175);
and U22690 (N_22690,N_21329,N_22333);
or U22691 (N_22691,N_20570,N_20746);
and U22692 (N_22692,N_20038,N_22092);
nor U22693 (N_22693,N_20017,N_20672);
and U22694 (N_22694,N_21575,N_20468);
or U22695 (N_22695,N_20964,N_20407);
or U22696 (N_22696,N_20391,N_20336);
and U22697 (N_22697,N_20365,N_20179);
and U22698 (N_22698,N_20553,N_22102);
nand U22699 (N_22699,N_22134,N_21888);
and U22700 (N_22700,N_22482,N_22430);
nor U22701 (N_22701,N_20894,N_22009);
or U22702 (N_22702,N_20174,N_20930);
or U22703 (N_22703,N_21464,N_21430);
xnor U22704 (N_22704,N_22336,N_21777);
xnor U22705 (N_22705,N_20714,N_20379);
nor U22706 (N_22706,N_21332,N_21410);
xor U22707 (N_22707,N_21435,N_21015);
or U22708 (N_22708,N_20502,N_20700);
xnor U22709 (N_22709,N_22078,N_22387);
and U22710 (N_22710,N_21944,N_21312);
and U22711 (N_22711,N_21063,N_21304);
xor U22712 (N_22712,N_21043,N_21414);
nor U22713 (N_22713,N_21601,N_22378);
nand U22714 (N_22714,N_20692,N_21104);
or U22715 (N_22715,N_20022,N_20357);
nand U22716 (N_22716,N_22086,N_22032);
nand U22717 (N_22717,N_21833,N_21810);
nand U22718 (N_22718,N_21254,N_22223);
xor U22719 (N_22719,N_22495,N_20994);
xor U22720 (N_22720,N_21244,N_21145);
xor U22721 (N_22721,N_21251,N_20169);
nand U22722 (N_22722,N_20158,N_20893);
nand U22723 (N_22723,N_22041,N_21560);
nor U22724 (N_22724,N_21404,N_20188);
or U22725 (N_22725,N_22262,N_20284);
nand U22726 (N_22726,N_20388,N_22181);
nor U22727 (N_22727,N_20682,N_20587);
xnor U22728 (N_22728,N_22375,N_20193);
and U22729 (N_22729,N_21458,N_22052);
nor U22730 (N_22730,N_21098,N_20062);
and U22731 (N_22731,N_22451,N_20092);
or U22732 (N_22732,N_20647,N_21815);
nor U22733 (N_22733,N_20624,N_20633);
nor U22734 (N_22734,N_22138,N_20549);
xnor U22735 (N_22735,N_22013,N_22279);
or U22736 (N_22736,N_21336,N_22003);
nand U22737 (N_22737,N_20929,N_21129);
xnor U22738 (N_22738,N_21327,N_20011);
or U22739 (N_22739,N_22199,N_22459);
nand U22740 (N_22740,N_21755,N_20910);
nand U22741 (N_22741,N_22443,N_20424);
nand U22742 (N_22742,N_21350,N_20988);
nand U22743 (N_22743,N_20612,N_21275);
and U22744 (N_22744,N_22379,N_21432);
nor U22745 (N_22745,N_21144,N_21459);
nor U22746 (N_22746,N_20747,N_22167);
nor U22747 (N_22747,N_21102,N_20475);
nor U22748 (N_22748,N_21599,N_21072);
nor U22749 (N_22749,N_20375,N_21240);
xor U22750 (N_22750,N_21107,N_22259);
xnor U22751 (N_22751,N_21218,N_22146);
nand U22752 (N_22752,N_22033,N_22230);
nor U22753 (N_22753,N_22208,N_22382);
or U22754 (N_22754,N_20386,N_20704);
nor U22755 (N_22755,N_20394,N_21689);
or U22756 (N_22756,N_21269,N_22469);
nand U22757 (N_22757,N_21487,N_20029);
xor U22758 (N_22758,N_22492,N_21525);
or U22759 (N_22759,N_20971,N_21213);
xnor U22760 (N_22760,N_21444,N_20013);
and U22761 (N_22761,N_21731,N_21208);
or U22762 (N_22762,N_21574,N_21033);
nand U22763 (N_22763,N_20716,N_22269);
xnor U22764 (N_22764,N_22174,N_22300);
nand U22765 (N_22765,N_20655,N_21583);
or U22766 (N_22766,N_20440,N_21553);
and U22767 (N_22767,N_21861,N_21516);
or U22768 (N_22768,N_21059,N_21073);
or U22769 (N_22769,N_21018,N_20795);
nor U22770 (N_22770,N_21120,N_21658);
or U22771 (N_22771,N_20069,N_20690);
nor U22772 (N_22772,N_22293,N_21252);
xnor U22773 (N_22773,N_20262,N_21858);
xor U22774 (N_22774,N_20505,N_20392);
and U22775 (N_22775,N_21303,N_20545);
or U22776 (N_22776,N_21155,N_22272);
nor U22777 (N_22777,N_22343,N_20044);
nand U22778 (N_22778,N_20884,N_21638);
xnor U22779 (N_22779,N_22211,N_21042);
or U22780 (N_22780,N_21103,N_21715);
xnor U22781 (N_22781,N_20945,N_20270);
or U22782 (N_22782,N_20769,N_20839);
nand U22783 (N_22783,N_20831,N_21050);
nor U22784 (N_22784,N_20710,N_22028);
or U22785 (N_22785,N_21076,N_20410);
and U22786 (N_22786,N_21649,N_22067);
and U22787 (N_22787,N_20264,N_20431);
nor U22788 (N_22788,N_20573,N_20707);
nor U22789 (N_22789,N_20686,N_22048);
nand U22790 (N_22790,N_20399,N_22317);
xor U22791 (N_22791,N_22065,N_20170);
nand U22792 (N_22792,N_21720,N_20983);
or U22793 (N_22793,N_20763,N_20138);
xnor U22794 (N_22794,N_21505,N_20100);
nand U22795 (N_22795,N_21097,N_21561);
nor U22796 (N_22796,N_20576,N_20511);
nand U22797 (N_22797,N_21562,N_21566);
nand U22798 (N_22798,N_21438,N_21694);
xor U22799 (N_22799,N_22038,N_20354);
and U22800 (N_22800,N_22235,N_21451);
xor U22801 (N_22801,N_22049,N_20905);
and U22802 (N_22802,N_20960,N_21573);
nand U22803 (N_22803,N_21316,N_21100);
nand U22804 (N_22804,N_20862,N_21533);
or U22805 (N_22805,N_22128,N_21877);
nor U22806 (N_22806,N_22422,N_22131);
and U22807 (N_22807,N_22148,N_20721);
nor U22808 (N_22808,N_21169,N_20742);
nor U22809 (N_22809,N_20081,N_20404);
and U22810 (N_22810,N_22346,N_21243);
or U22811 (N_22811,N_20998,N_22018);
nand U22812 (N_22812,N_21531,N_22105);
nor U22813 (N_22813,N_20183,N_22404);
nor U22814 (N_22814,N_22000,N_21346);
and U22815 (N_22815,N_22447,N_21283);
xnor U22816 (N_22816,N_20372,N_21886);
xnor U22817 (N_22817,N_20737,N_20319);
and U22818 (N_22818,N_20213,N_20579);
nand U22819 (N_22819,N_21189,N_20050);
nand U22820 (N_22820,N_21969,N_22386);
nor U22821 (N_22821,N_21831,N_22185);
xnor U22822 (N_22822,N_20030,N_21365);
xnor U22823 (N_22823,N_21276,N_20796);
or U22824 (N_22824,N_20513,N_20032);
or U22825 (N_22825,N_20874,N_22410);
nand U22826 (N_22826,N_21670,N_22420);
nor U22827 (N_22827,N_21004,N_21622);
xor U22828 (N_22828,N_21342,N_21422);
or U22829 (N_22829,N_22154,N_20871);
nand U22830 (N_22830,N_21749,N_21210);
xnor U22831 (N_22831,N_20412,N_20248);
nor U22832 (N_22832,N_20973,N_21138);
nor U22833 (N_22833,N_21361,N_21126);
and U22834 (N_22834,N_20259,N_21750);
or U22835 (N_22835,N_20509,N_20359);
and U22836 (N_22836,N_21260,N_20421);
nand U22837 (N_22837,N_22318,N_21871);
nor U22838 (N_22838,N_21954,N_20129);
nand U22839 (N_22839,N_20478,N_21899);
nor U22840 (N_22840,N_20827,N_20896);
nand U22841 (N_22841,N_21272,N_21051);
xor U22842 (N_22842,N_22302,N_22286);
or U22843 (N_22843,N_21513,N_22393);
or U22844 (N_22844,N_21475,N_21201);
nand U22845 (N_22845,N_20318,N_20026);
xnor U22846 (N_22846,N_21473,N_20177);
nand U22847 (N_22847,N_20396,N_21439);
nand U22848 (N_22848,N_22489,N_22054);
nor U22849 (N_22849,N_20922,N_21578);
nand U22850 (N_22850,N_21854,N_20271);
nand U22851 (N_22851,N_21445,N_21463);
xor U22852 (N_22852,N_22465,N_21509);
nor U22853 (N_22853,N_21468,N_22096);
or U22854 (N_22854,N_20631,N_20112);
nor U22855 (N_22855,N_22010,N_20901);
or U22856 (N_22856,N_20851,N_21682);
and U22857 (N_22857,N_21448,N_21988);
nand U22858 (N_22858,N_20565,N_20476);
and U22859 (N_22859,N_21081,N_20383);
nor U22860 (N_22860,N_22361,N_20317);
nor U22861 (N_22861,N_21331,N_22209);
nand U22862 (N_22862,N_20167,N_21974);
nor U22863 (N_22863,N_22347,N_21202);
xnor U22864 (N_22864,N_20992,N_21299);
and U22865 (N_22865,N_21710,N_21310);
or U22866 (N_22866,N_20149,N_21902);
nor U22867 (N_22867,N_21068,N_22412);
or U22868 (N_22868,N_21328,N_21934);
nor U22869 (N_22869,N_20217,N_20915);
or U22870 (N_22870,N_21701,N_20669);
and U22871 (N_22871,N_20205,N_20060);
nor U22872 (N_22872,N_20997,N_20961);
or U22873 (N_22873,N_22168,N_21693);
xor U22874 (N_22874,N_20275,N_22456);
nor U22875 (N_22875,N_22110,N_21423);
or U22876 (N_22876,N_21768,N_21061);
xor U22877 (N_22877,N_20991,N_21669);
nand U22878 (N_22878,N_21677,N_22156);
and U22879 (N_22879,N_20738,N_21297);
nor U22880 (N_22880,N_21676,N_21472);
or U22881 (N_22881,N_21270,N_20472);
and U22882 (N_22882,N_20969,N_21730);
nand U22883 (N_22883,N_21616,N_20572);
nand U22884 (N_22884,N_20504,N_20406);
nor U22885 (N_22885,N_20249,N_20417);
or U22886 (N_22886,N_22149,N_21363);
nand U22887 (N_22887,N_22257,N_20965);
xor U22888 (N_22888,N_21140,N_20838);
nor U22889 (N_22889,N_20401,N_21674);
and U22890 (N_22890,N_20215,N_20393);
nor U22891 (N_22891,N_21937,N_20590);
xnor U22892 (N_22892,N_20168,N_20643);
xnor U22893 (N_22893,N_21844,N_20462);
and U22894 (N_22894,N_20895,N_20277);
xor U22895 (N_22895,N_21591,N_20024);
nor U22896 (N_22896,N_22483,N_21074);
and U22897 (N_22897,N_22188,N_20739);
or U22898 (N_22898,N_22403,N_21485);
or U22899 (N_22899,N_22161,N_20508);
or U22900 (N_22900,N_21391,N_21807);
or U22901 (N_22901,N_20306,N_20510);
or U22902 (N_22902,N_21418,N_20434);
or U22903 (N_22903,N_21985,N_20708);
or U22904 (N_22904,N_21228,N_20524);
nand U22905 (N_22905,N_21953,N_22425);
xnor U22906 (N_22906,N_20904,N_21795);
nor U22907 (N_22907,N_20157,N_20857);
or U22908 (N_22908,N_20315,N_22275);
or U22909 (N_22909,N_21034,N_20449);
nand U22910 (N_22910,N_20280,N_20935);
or U22911 (N_22911,N_21956,N_22159);
or U22912 (N_22912,N_20684,N_20008);
or U22913 (N_22913,N_20597,N_20909);
and U22914 (N_22914,N_22005,N_22215);
or U22915 (N_22915,N_21172,N_22113);
and U22916 (N_22916,N_22352,N_20889);
nand U22917 (N_22917,N_21963,N_22370);
and U22918 (N_22918,N_20483,N_22081);
xnor U22919 (N_22919,N_20558,N_21150);
nor U22920 (N_22920,N_21241,N_22281);
xnor U22921 (N_22921,N_22354,N_21428);
and U22922 (N_22922,N_20660,N_20629);
and U22923 (N_22923,N_22255,N_20611);
nand U22924 (N_22924,N_20046,N_22416);
nor U22925 (N_22925,N_22397,N_22409);
and U22926 (N_22926,N_20976,N_22187);
or U22927 (N_22927,N_21176,N_21800);
or U22928 (N_22928,N_22458,N_22419);
xnor U22929 (N_22929,N_21538,N_20054);
and U22930 (N_22930,N_20699,N_21862);
or U22931 (N_22931,N_21044,N_21832);
nor U22932 (N_22932,N_21402,N_21453);
xor U22933 (N_22933,N_20566,N_22031);
nor U22934 (N_22934,N_20162,N_20731);
nor U22935 (N_22935,N_20844,N_21216);
nand U22936 (N_22936,N_22042,N_21398);
and U22937 (N_22937,N_21023,N_20772);
or U22938 (N_22938,N_22027,N_20543);
and U22939 (N_22939,N_21685,N_22098);
and U22940 (N_22940,N_21734,N_22248);
nand U22941 (N_22941,N_21727,N_21757);
xor U22942 (N_22942,N_21640,N_21829);
or U22943 (N_22943,N_22225,N_21535);
or U22944 (N_22944,N_20286,N_21142);
xnor U22945 (N_22945,N_22408,N_21412);
nor U22946 (N_22946,N_20148,N_20564);
nor U22947 (N_22947,N_20529,N_22219);
nand U22948 (N_22948,N_20822,N_20115);
or U22949 (N_22949,N_22170,N_21582);
nor U22950 (N_22950,N_21700,N_20428);
nor U22951 (N_22951,N_21612,N_21083);
or U22952 (N_22952,N_21699,N_21116);
nand U22953 (N_22953,N_20160,N_21349);
nor U22954 (N_22954,N_20923,N_20141);
or U22955 (N_22955,N_20789,N_22457);
nand U22956 (N_22956,N_20812,N_21062);
nor U22957 (N_22957,N_21186,N_20773);
xor U22958 (N_22958,N_21778,N_21580);
nand U22959 (N_22959,N_20150,N_21747);
xor U22960 (N_22960,N_20864,N_21501);
nor U22961 (N_22961,N_21719,N_21457);
xor U22962 (N_22962,N_22319,N_21596);
nand U22963 (N_22963,N_20202,N_20124);
nor U22964 (N_22964,N_21340,N_21819);
nand U22965 (N_22965,N_21409,N_22202);
or U22966 (N_22966,N_20451,N_22133);
or U22967 (N_22967,N_20729,N_22401);
nand U22968 (N_22968,N_21668,N_20438);
nor U22969 (N_22969,N_20103,N_20722);
xnor U22970 (N_22970,N_20546,N_20637);
and U22971 (N_22971,N_21318,N_20569);
and U22972 (N_22972,N_21197,N_21864);
or U22973 (N_22973,N_21047,N_20414);
or U22974 (N_22974,N_21787,N_20845);
nand U22975 (N_22975,N_21357,N_21976);
xor U22976 (N_22976,N_22320,N_20768);
nor U22977 (N_22977,N_22076,N_20327);
xnor U22978 (N_22978,N_20544,N_21069);
or U22979 (N_22979,N_20912,N_20028);
xnor U22980 (N_22980,N_21752,N_20485);
and U22981 (N_22981,N_20837,N_20120);
nor U22982 (N_22982,N_20783,N_21762);
and U22983 (N_22983,N_21781,N_20418);
and U22984 (N_22984,N_22206,N_20518);
and U22985 (N_22985,N_20863,N_21941);
xnor U22986 (N_22986,N_21306,N_20940);
nand U22987 (N_22987,N_21222,N_22016);
xnor U22988 (N_22988,N_21766,N_20875);
nand U22989 (N_22989,N_21427,N_22080);
xor U22990 (N_22990,N_20490,N_20928);
or U22991 (N_22991,N_22073,N_21166);
nand U22992 (N_22992,N_21027,N_21882);
and U22993 (N_22993,N_20776,N_21503);
and U22994 (N_22994,N_20650,N_20238);
and U22995 (N_22995,N_21587,N_21746);
or U22996 (N_22996,N_21519,N_21654);
nor U22997 (N_22997,N_21095,N_21170);
nand U22998 (N_22998,N_22197,N_20450);
or U22999 (N_22999,N_20254,N_22474);
xnor U23000 (N_23000,N_21697,N_20094);
nand U23001 (N_23001,N_21784,N_21199);
nand U23002 (N_23002,N_21950,N_21500);
or U23003 (N_23003,N_20606,N_21977);
nand U23004 (N_23004,N_20480,N_20353);
xnor U23005 (N_23005,N_20715,N_22189);
and U23006 (N_23006,N_22119,N_22367);
or U23007 (N_23007,N_22198,N_22093);
and U23008 (N_23008,N_20951,N_21052);
or U23009 (N_23009,N_20163,N_21122);
nand U23010 (N_23010,N_20724,N_22251);
or U23011 (N_23011,N_20580,N_21659);
or U23012 (N_23012,N_20134,N_20500);
or U23013 (N_23013,N_21743,N_20229);
and U23014 (N_23014,N_22481,N_21075);
nand U23015 (N_23015,N_20679,N_22288);
or U23016 (N_23016,N_21392,N_20197);
and U23017 (N_23017,N_22112,N_21966);
or U23018 (N_23018,N_20279,N_22353);
xor U23019 (N_23019,N_20899,N_21112);
xnor U23020 (N_23020,N_20903,N_20185);
xor U23021 (N_23021,N_20970,N_21291);
nor U23022 (N_23022,N_20937,N_21737);
and U23023 (N_23023,N_21265,N_20528);
xor U23024 (N_23024,N_22444,N_22123);
nand U23025 (N_23025,N_20782,N_22358);
nor U23026 (N_23026,N_20240,N_21823);
and U23027 (N_23027,N_21631,N_22173);
xor U23028 (N_23028,N_21707,N_20626);
or U23029 (N_23029,N_20374,N_20642);
and U23030 (N_23030,N_20657,N_20435);
nor U23031 (N_23031,N_21086,N_22280);
and U23032 (N_23032,N_21264,N_21588);
xnor U23033 (N_23033,N_22087,N_20539);
nor U23034 (N_23034,N_22147,N_21021);
nor U23035 (N_23035,N_22195,N_20256);
nand U23036 (N_23036,N_21991,N_20493);
or U23037 (N_23037,N_20974,N_21756);
or U23038 (N_23038,N_21147,N_21420);
or U23039 (N_23039,N_20987,N_20826);
nor U23040 (N_23040,N_21825,N_21753);
or U23041 (N_23041,N_20664,N_20473);
xor U23042 (N_23042,N_20661,N_22239);
or U23043 (N_23043,N_21364,N_20314);
or U23044 (N_23044,N_21971,N_21286);
nor U23045 (N_23045,N_20615,N_20726);
and U23046 (N_23046,N_22470,N_20368);
nand U23047 (N_23047,N_22231,N_22476);
nor U23048 (N_23048,N_20709,N_20364);
nand U23049 (N_23049,N_20944,N_21704);
xnor U23050 (N_23050,N_22229,N_21173);
nand U23051 (N_23051,N_21511,N_20653);
and U23052 (N_23052,N_21443,N_22126);
or U23053 (N_23053,N_21366,N_20021);
nand U23054 (N_23054,N_21177,N_21188);
nor U23055 (N_23055,N_21396,N_20599);
and U23056 (N_23056,N_20577,N_21552);
and U23057 (N_23057,N_20823,N_21184);
nand U23058 (N_23058,N_20191,N_20433);
nand U23059 (N_23059,N_21775,N_20770);
or U23060 (N_23060,N_21014,N_22285);
and U23061 (N_23061,N_20016,N_20403);
nand U23062 (N_23062,N_21776,N_20766);
xnor U23063 (N_23063,N_20460,N_20931);
or U23064 (N_23064,N_21118,N_20550);
and U23065 (N_23065,N_20087,N_22323);
nand U23066 (N_23066,N_21493,N_22363);
nand U23067 (N_23067,N_21191,N_20430);
and U23068 (N_23068,N_22043,N_21078);
nor U23069 (N_23069,N_21797,N_21728);
xor U23070 (N_23070,N_21317,N_20588);
xnor U23071 (N_23071,N_21980,N_20950);
xor U23072 (N_23072,N_21137,N_21030);
and U23073 (N_23073,N_21494,N_22190);
nand U23074 (N_23074,N_20982,N_21986);
xnor U23075 (N_23075,N_21071,N_21065);
xnor U23076 (N_23076,N_21678,N_21817);
or U23077 (N_23077,N_22267,N_21314);
nor U23078 (N_23078,N_20332,N_20990);
nand U23079 (N_23079,N_21037,N_21554);
xor U23080 (N_23080,N_21106,N_22282);
xor U23081 (N_23081,N_20334,N_20618);
nand U23082 (N_23082,N_20497,N_20300);
nor U23083 (N_23083,N_20192,N_21579);
xor U23084 (N_23084,N_21930,N_21632);
nor U23085 (N_23085,N_21779,N_20762);
nor U23086 (N_23086,N_21653,N_22383);
nor U23087 (N_23087,N_21568,N_21066);
or U23088 (N_23088,N_21231,N_20211);
xnor U23089 (N_23089,N_20146,N_20233);
or U23090 (N_23090,N_20859,N_20322);
or U23091 (N_23091,N_21245,N_22256);
nor U23092 (N_23092,N_20972,N_21267);
xor U23093 (N_23093,N_21146,N_20911);
xnor U23094 (N_23094,N_22019,N_20219);
nor U23095 (N_23095,N_22026,N_20757);
or U23096 (N_23096,N_21308,N_21528);
nor U23097 (N_23097,N_21972,N_21232);
nand U23098 (N_23098,N_20405,N_21824);
or U23099 (N_23099,N_22107,N_20891);
nor U23100 (N_23100,N_20562,N_21159);
nand U23101 (N_23101,N_21151,N_22338);
and U23102 (N_23102,N_22150,N_20328);
nand U23103 (N_23103,N_21648,N_21036);
or U23104 (N_23104,N_20880,N_20519);
or U23105 (N_23105,N_22284,N_22454);
xnor U23106 (N_23106,N_21959,N_21325);
or U23107 (N_23107,N_21206,N_22322);
xnor U23108 (N_23108,N_22436,N_22226);
nor U23109 (N_23109,N_21226,N_20114);
and U23110 (N_23110,N_21606,N_21896);
nor U23111 (N_23111,N_21292,N_20463);
and U23112 (N_23112,N_22166,N_22461);
nand U23113 (N_23113,N_20887,N_20761);
nor U23114 (N_23114,N_21132,N_22271);
xnor U23115 (N_23115,N_20220,N_20701);
and U23116 (N_23116,N_22292,N_20750);
nor U23117 (N_23117,N_22467,N_21408);
nor U23118 (N_23118,N_22157,N_22283);
or U23119 (N_23119,N_22260,N_20196);
nor U23120 (N_23120,N_22310,N_21915);
nand U23121 (N_23121,N_21522,N_21725);
nor U23122 (N_23122,N_20173,N_21960);
nor U23123 (N_23123,N_21373,N_20201);
nand U23124 (N_23124,N_20936,N_20836);
or U23125 (N_23125,N_21470,N_21914);
nor U23126 (N_23126,N_21751,N_20145);
nand U23127 (N_23127,N_22244,N_21761);
and U23128 (N_23128,N_22136,N_20272);
or U23129 (N_23129,N_21281,N_21482);
and U23130 (N_23130,N_22077,N_20584);
nor U23131 (N_23131,N_22108,N_21742);
nor U23132 (N_23132,N_22008,N_21355);
and U23133 (N_23133,N_21376,N_20395);
and U23134 (N_23134,N_20603,N_20458);
and U23135 (N_23135,N_20257,N_22095);
xor U23136 (N_23136,N_22139,N_20978);
nor U23137 (N_23137,N_21353,N_20846);
and U23138 (N_23138,N_22037,N_20890);
nand U23139 (N_23139,N_20154,N_21556);
xnor U23140 (N_23140,N_21995,N_21827);
nor U23141 (N_23141,N_20304,N_20361);
and U23142 (N_23142,N_20996,N_21656);
nand U23143 (N_23143,N_20678,N_20126);
nand U23144 (N_23144,N_22124,N_21796);
or U23145 (N_23145,N_20481,N_21399);
nor U23146 (N_23146,N_20342,N_21491);
and U23147 (N_23147,N_21646,N_20045);
xor U23148 (N_23148,N_21602,N_21339);
xnor U23149 (N_23149,N_21156,N_20556);
and U23150 (N_23150,N_22423,N_20064);
nand U23151 (N_23151,N_21925,N_22394);
or U23152 (N_23152,N_20047,N_21168);
and U23153 (N_23153,N_22261,N_20258);
nor U23154 (N_23154,N_20883,N_20495);
nand U23155 (N_23155,N_21792,N_20420);
nand U23156 (N_23156,N_21359,N_22486);
and U23157 (N_23157,N_22210,N_20609);
and U23158 (N_23158,N_20130,N_21544);
xnor U23159 (N_23159,N_21683,N_21087);
or U23160 (N_23160,N_22127,N_21124);
xnor U23161 (N_23161,N_21386,N_21564);
or U23162 (N_23162,N_20116,N_22182);
xor U23163 (N_23163,N_22324,N_22030);
and U23164 (N_23164,N_20876,N_21157);
and U23165 (N_23165,N_20614,N_21869);
or U23166 (N_23166,N_22106,N_22220);
nor U23167 (N_23167,N_22303,N_20625);
or U23168 (N_23168,N_22274,N_21952);
or U23169 (N_23169,N_21032,N_20470);
or U23170 (N_23170,N_22143,N_21508);
xor U23171 (N_23171,N_21900,N_21961);
xor U23172 (N_23172,N_20413,N_20753);
and U23173 (N_23173,N_20012,N_20809);
xnor U23174 (N_23174,N_21760,N_20226);
and U23175 (N_23175,N_21456,N_21708);
and U23176 (N_23176,N_20132,N_22046);
or U23177 (N_23177,N_21916,N_20740);
nor U23178 (N_23178,N_20097,N_22463);
or U23179 (N_23179,N_20207,N_21436);
xnor U23180 (N_23180,N_20819,N_22306);
and U23181 (N_23181,N_21135,N_20242);
xnor U23182 (N_23182,N_21724,N_21866);
xnor U23183 (N_23183,N_20355,N_20946);
or U23184 (N_23184,N_21238,N_21948);
nor U23185 (N_23185,N_21909,N_22417);
and U23186 (N_23186,N_20377,N_21617);
and U23187 (N_23187,N_21835,N_20914);
or U23188 (N_23188,N_21857,N_20156);
nand U23189 (N_23189,N_20068,N_20052);
nor U23190 (N_23190,N_22331,N_20833);
xnor U23191 (N_23191,N_21613,N_20037);
nor U23192 (N_23192,N_20681,N_21618);
nand U23193 (N_23193,N_21165,N_22015);
or U23194 (N_23194,N_20072,N_21028);
and U23195 (N_23195,N_21041,N_22207);
nor U23196 (N_23196,N_21894,N_21884);
xor U23197 (N_23197,N_21060,N_21913);
nor U23198 (N_23198,N_21225,N_20437);
nand U23199 (N_23199,N_20730,N_20203);
or U23200 (N_23200,N_20919,N_20411);
nor U23201 (N_23201,N_20767,N_21007);
and U23202 (N_23202,N_20814,N_20535);
and U23203 (N_23203,N_21876,N_21279);
nor U23204 (N_23204,N_21480,N_21341);
nor U23205 (N_23205,N_21319,N_20855);
nor U23206 (N_23206,N_20425,N_21219);
or U23207 (N_23207,N_22390,N_21735);
and U23208 (N_23208,N_22301,N_20198);
xor U23209 (N_23209,N_21856,N_21629);
and U23210 (N_23210,N_22396,N_20015);
nand U23211 (N_23211,N_21195,N_21039);
nor U23212 (N_23212,N_21982,N_21549);
and U23213 (N_23213,N_21250,N_21924);
or U23214 (N_23214,N_21598,N_21287);
and U23215 (N_23215,N_20489,N_22213);
nand U23216 (N_23216,N_20989,N_21460);
or U23217 (N_23217,N_20019,N_20245);
and U23218 (N_23218,N_21242,N_20695);
nand U23219 (N_23219,N_22277,N_20253);
or U23220 (N_23220,N_20454,N_21105);
and U23221 (N_23221,N_21025,N_21111);
nor U23222 (N_23222,N_21117,N_21431);
and U23223 (N_23223,N_20531,N_20218);
and U23224 (N_23224,N_22122,N_21313);
nand U23225 (N_23225,N_20804,N_20065);
xor U23226 (N_23226,N_21221,N_20640);
nand U23227 (N_23227,N_20706,N_20184);
xor U23228 (N_23228,N_20080,N_20427);
xnor U23229 (N_23229,N_22428,N_21984);
or U23230 (N_23230,N_21057,N_20073);
nor U23231 (N_23231,N_21738,N_21022);
or U23232 (N_23232,N_20477,N_21630);
or U23233 (N_23233,N_20494,N_21527);
nor U23234 (N_23234,N_20540,N_21397);
or U23235 (N_23235,N_20852,N_22247);
and U23236 (N_23236,N_21469,N_21808);
xor U23237 (N_23237,N_20155,N_21164);
and U23238 (N_23238,N_21239,N_21001);
or U23239 (N_23239,N_22001,N_21012);
or U23240 (N_23240,N_20696,N_21178);
nand U23241 (N_23241,N_20415,N_21506);
nand U23242 (N_23242,N_21530,N_21008);
xnor U23243 (N_23243,N_22350,N_22017);
xnor U23244 (N_23244,N_21193,N_21290);
xnor U23245 (N_23245,N_21031,N_20137);
and U23246 (N_23246,N_20107,N_21371);
nand U23247 (N_23247,N_22222,N_21998);
or U23248 (N_23248,N_22291,N_22140);
or U23249 (N_23249,N_21337,N_22485);
nand U23250 (N_23250,N_21774,N_20268);
xor U23251 (N_23251,N_21951,N_20853);
and U23252 (N_23252,N_20109,N_21446);
xor U23253 (N_23253,N_21983,N_20778);
and U23254 (N_23254,N_20224,N_21927);
nor U23255 (N_23255,N_21706,N_21127);
nand U23256 (N_23256,N_21875,N_22103);
and U23257 (N_23257,N_22071,N_22011);
nand U23258 (N_23258,N_21623,N_21608);
nor U23259 (N_23259,N_21628,N_22084);
nor U23260 (N_23260,N_22389,N_21079);
or U23261 (N_23261,N_21826,N_22221);
nor U23262 (N_23262,N_20082,N_21326);
and U23263 (N_23263,N_20947,N_21148);
nor U23264 (N_23264,N_21358,N_20781);
xnor U23265 (N_23265,N_21055,N_21449);
xnor U23266 (N_23266,N_20547,N_21437);
or U23267 (N_23267,N_21054,N_20351);
or U23268 (N_23268,N_20526,N_21489);
xor U23269 (N_23269,N_21058,N_20986);
nand U23270 (N_23270,N_21285,N_20181);
or U23271 (N_23271,N_21885,N_21235);
and U23272 (N_23272,N_20210,N_22218);
nor U23273 (N_23273,N_21465,N_20190);
and U23274 (N_23274,N_22258,N_20005);
and U23275 (N_23275,N_20252,N_20824);
and U23276 (N_23276,N_20627,N_21394);
nor U23277 (N_23277,N_21722,N_20829);
nand U23278 (N_23278,N_21476,N_21758);
nor U23279 (N_23279,N_21088,N_21383);
and U23280 (N_23280,N_21788,N_21666);
nand U23281 (N_23281,N_21548,N_21978);
or U23282 (N_23282,N_20907,N_22162);
and U23283 (N_23283,N_20952,N_20702);
xnor U23284 (N_23284,N_22204,N_21152);
nor U23285 (N_23285,N_21223,N_21483);
or U23286 (N_23286,N_20409,N_22471);
nand U23287 (N_23287,N_20491,N_21005);
or U23288 (N_23288,N_22496,N_21565);
or U23289 (N_23289,N_20467,N_20443);
nor U23290 (N_23290,N_22304,N_20802);
or U23291 (N_23291,N_22097,N_20538);
nand U23292 (N_23292,N_20265,N_21684);
nor U23293 (N_23293,N_20204,N_21214);
nor U23294 (N_23294,N_20232,N_21745);
nor U23295 (N_23295,N_21455,N_20208);
and U23296 (N_23296,N_21946,N_20847);
nand U23297 (N_23297,N_22090,N_21790);
xnor U23298 (N_23298,N_22035,N_21090);
nor U23299 (N_23299,N_21154,N_21248);
or U23300 (N_23300,N_21153,N_22176);
or U23301 (N_23301,N_20330,N_20369);
xor U23302 (N_23302,N_21035,N_21791);
xor U23303 (N_23303,N_21813,N_21537);
xnor U23304 (N_23304,N_20464,N_20771);
nor U23305 (N_23305,N_21863,N_22082);
nor U23306 (N_23306,N_20456,N_20744);
nor U23307 (N_23307,N_20594,N_21624);
nor U23308 (N_23308,N_21492,N_20906);
or U23309 (N_23309,N_22024,N_20736);
nor U23310 (N_23310,N_20711,N_21679);
or U23311 (N_23311,N_22044,N_21979);
nand U23312 (N_23312,N_20638,N_22120);
or U23313 (N_23313,N_20231,N_20093);
or U23314 (N_23314,N_22371,N_20765);
or U23315 (N_23315,N_22344,N_21965);
and U23316 (N_23316,N_20039,N_21918);
and U23317 (N_23317,N_20096,N_21415);
nand U23318 (N_23318,N_21429,N_20759);
nor U23319 (N_23319,N_20607,N_21217);
and U23320 (N_23320,N_22365,N_21237);
nand U23321 (N_23321,N_21763,N_20658);
and U23322 (N_23322,N_21479,N_21056);
xor U23323 (N_23323,N_22184,N_21294);
nor U23324 (N_23324,N_21794,N_20628);
nand U23325 (N_23325,N_20581,N_20004);
nand U23326 (N_23326,N_21904,N_20601);
or U23327 (N_23327,N_20261,N_20598);
nand U23328 (N_23328,N_20820,N_22063);
or U23329 (N_23329,N_22357,N_20419);
and U23330 (N_23330,N_21113,N_22224);
nand U23331 (N_23331,N_20320,N_20118);
and U23332 (N_23332,N_21996,N_21049);
xor U23333 (N_23333,N_22414,N_21536);
nor U23334 (N_23334,N_20641,N_20142);
nor U23335 (N_23335,N_20324,N_21119);
nor U23336 (N_23336,N_22290,N_21401);
xor U23337 (N_23337,N_20723,N_20358);
xnor U23338 (N_23338,N_21822,N_21639);
nor U23339 (N_23339,N_20604,N_21017);
nor U23340 (N_23340,N_20645,N_21769);
nor U23341 (N_23341,N_22473,N_22061);
or U23342 (N_23342,N_21387,N_20595);
or U23343 (N_23343,N_21253,N_22012);
nand U23344 (N_23344,N_20559,N_21298);
and U23345 (N_23345,N_20745,N_20484);
nor U23346 (N_23346,N_21657,N_22214);
nor U23347 (N_23347,N_21921,N_21284);
nand U23348 (N_23348,N_20525,N_21230);
and U23349 (N_23349,N_21085,N_21024);
nor U23350 (N_23350,N_21892,N_21070);
nand U23351 (N_23351,N_20886,N_21183);
nor U23352 (N_23352,N_21003,N_20041);
xnor U23353 (N_23353,N_21484,N_21064);
or U23354 (N_23354,N_22493,N_20617);
and U23355 (N_23355,N_20533,N_22487);
and U23356 (N_23356,N_21406,N_20340);
nor U23357 (N_23357,N_21377,N_22152);
nand U23358 (N_23358,N_21301,N_22007);
nand U23359 (N_23359,N_20866,N_21801);
nand U23360 (N_23360,N_21868,N_21271);
xor U23361 (N_23361,N_20622,N_21692);
nand U23362 (N_23362,N_21077,N_20378);
and U23363 (N_23363,N_20648,N_20371);
nand U23364 (N_23364,N_21322,N_21433);
or U23365 (N_23365,N_21013,N_20346);
nand U23366 (N_23366,N_20189,N_20878);
xnor U23367 (N_23367,N_20200,N_22391);
nand U23368 (N_23368,N_21662,N_22326);
or U23369 (N_23369,N_20806,N_20278);
and U23370 (N_23370,N_21939,N_21733);
or U23371 (N_23371,N_20063,N_20447);
xnor U23372 (N_23372,N_20542,N_20499);
or U23373 (N_23373,N_22421,N_22178);
or U23374 (N_23374,N_20244,N_20635);
and U23375 (N_23375,N_21711,N_22099);
nand U23376 (N_23376,N_21690,N_21504);
or U23377 (N_23377,N_20981,N_21696);
nor U23378 (N_23378,N_20343,N_21614);
and U23379 (N_23379,N_21589,N_20832);
and U23380 (N_23380,N_21785,N_21205);
xnor U23381 (N_23381,N_21417,N_20326);
nand U23382 (N_23382,N_22464,N_21010);
nor U23383 (N_23383,N_20925,N_21200);
or U23384 (N_23384,N_20321,N_22392);
nand U23385 (N_23385,N_22313,N_20250);
xnor U23386 (N_23386,N_22289,N_20541);
or U23387 (N_23387,N_20995,N_20956);
and U23388 (N_23388,N_22186,N_22064);
xor U23389 (N_23389,N_21563,N_20216);
or U23390 (N_23390,N_21663,N_21981);
xnor U23391 (N_23391,N_21233,N_22266);
xor U23392 (N_23392,N_22045,N_20305);
or U23393 (N_23393,N_20380,N_20125);
xnor U23394 (N_23394,N_20152,N_20941);
xnor U23395 (N_23395,N_21997,N_22298);
or U23396 (N_23396,N_21084,N_20127);
xor U23397 (N_23397,N_21296,N_20975);
or U23398 (N_23398,N_22254,N_21542);
nand U23399 (N_23399,N_21634,N_21262);
and U23400 (N_23400,N_22494,N_20780);
and U23401 (N_23401,N_20734,N_21847);
and U23402 (N_23402,N_20131,N_22243);
xnor U23403 (N_23403,N_21302,N_22121);
and U23404 (N_23404,N_20234,N_21680);
nor U23405 (N_23405,N_20675,N_21619);
nor U23406 (N_23406,N_20151,N_22200);
or U23407 (N_23407,N_21257,N_21246);
xnor U23408 (N_23408,N_22193,N_21375);
or U23409 (N_23409,N_21323,N_20713);
nand U23410 (N_23410,N_22183,N_21179);
nand U23411 (N_23411,N_20416,N_21931);
nor U23412 (N_23412,N_21764,N_22196);
nor U23413 (N_23413,N_20848,N_20632);
nor U23414 (N_23414,N_20237,N_21258);
or U23415 (N_23415,N_20933,N_22431);
or U23416 (N_23416,N_21799,N_21295);
nand U23417 (N_23417,N_21645,N_21450);
nor U23418 (N_23418,N_20465,N_21236);
nor U23419 (N_23419,N_20522,N_21517);
xnor U23420 (N_23420,N_22025,N_22498);
xnor U23421 (N_23421,N_20387,N_22216);
xnor U23422 (N_23422,N_21607,N_21092);
and U23423 (N_23423,N_21873,N_21524);
or U23424 (N_23424,N_21134,N_21973);
or U23425 (N_23425,N_20133,N_20743);
nor U23426 (N_23426,N_21903,N_21515);
or U23427 (N_23427,N_21425,N_20908);
nor U23428 (N_23428,N_20673,N_21783);
or U23429 (N_23429,N_20059,N_21812);
or U23430 (N_23430,N_20861,N_21765);
nand U23431 (N_23431,N_20333,N_21293);
nor U23432 (N_23432,N_20943,N_22232);
or U23433 (N_23433,N_21040,N_22068);
and U23434 (N_23434,N_20613,N_20273);
xor U23435 (N_23435,N_22006,N_21748);
nor U23436 (N_23436,N_20111,N_20159);
nor U23437 (N_23437,N_20140,N_22115);
nor U23438 (N_23438,N_20344,N_20591);
xnor U23439 (N_23439,N_20298,N_20119);
nor U23440 (N_23440,N_22360,N_22278);
xor U23441 (N_23441,N_20345,N_21454);
nand U23442 (N_23442,N_22334,N_21786);
nor U23443 (N_23443,N_20551,N_21620);
xnor U23444 (N_23444,N_20805,N_22330);
nor U23445 (N_23445,N_21249,N_20791);
xor U23446 (N_23446,N_20792,N_20939);
xnor U23447 (N_23447,N_20786,N_20917);
nor U23448 (N_23448,N_20608,N_20984);
xor U23449 (N_23449,N_22250,N_21263);
nor U23450 (N_23450,N_21546,N_21577);
or U23451 (N_23451,N_20955,N_21912);
nor U23452 (N_23452,N_21718,N_20180);
or U23453 (N_23453,N_21928,N_21089);
nor U23454 (N_23454,N_21128,N_22050);
and U23455 (N_23455,N_20356,N_21917);
nand U23456 (N_23456,N_21158,N_20921);
and U23457 (N_23457,N_21424,N_20496);
and U23458 (N_23458,N_22433,N_22449);
and U23459 (N_23459,N_20408,N_20090);
nand U23460 (N_23460,N_20868,N_22117);
xor U23461 (N_23461,N_21234,N_21975);
xnor U23462 (N_23462,N_21627,N_20733);
and U23463 (N_23463,N_21671,N_20680);
or U23464 (N_23464,N_21502,N_20002);
or U23465 (N_23465,N_21721,N_20957);
nor U23466 (N_23466,N_20003,N_21362);
nor U23467 (N_23467,N_20293,N_22268);
nor U23468 (N_23468,N_21229,N_20793);
nand U23469 (N_23469,N_20582,N_21780);
or U23470 (N_23470,N_20398,N_20400);
nor U23471 (N_23471,N_21413,N_22349);
nand U23472 (N_23472,N_21344,N_20106);
or U23473 (N_23473,N_20662,N_21215);
and U23474 (N_23474,N_20441,N_20754);
xnor U23475 (N_23475,N_21955,N_21782);
nor U23476 (N_23476,N_20717,N_21926);
nand U23477 (N_23477,N_20209,N_20329);
xor U23478 (N_23478,N_21712,N_20312);
nand U23479 (N_23479,N_21604,N_20779);
nor U23480 (N_23480,N_21203,N_20752);
xor U23481 (N_23481,N_22137,N_20390);
and U23482 (N_23482,N_20561,N_21321);
and U23483 (N_23483,N_20292,N_20195);
nand U23484 (N_23484,N_22479,N_22135);
or U23485 (N_23485,N_20498,N_21793);
xnor U23486 (N_23486,N_21182,N_21938);
nor U23487 (N_23487,N_22132,N_21026);
nor U23488 (N_23488,N_20241,N_21163);
or U23489 (N_23489,N_22448,N_20840);
xnor U23490 (N_23490,N_21067,N_22328);
or U23491 (N_23491,N_21462,N_21860);
nor U23492 (N_23492,N_22014,N_22384);
nand U23493 (N_23493,N_21002,N_21839);
and U23494 (N_23494,N_20882,N_20164);
nand U23495 (N_23495,N_22308,N_20139);
nor U23496 (N_23496,N_21702,N_20482);
xnor U23497 (N_23497,N_21351,N_21277);
or U23498 (N_23498,N_21655,N_20110);
and U23499 (N_23499,N_20166,N_22020);
nand U23500 (N_23500,N_21315,N_21198);
nor U23501 (N_23501,N_20206,N_20807);
nand U23502 (N_23502,N_20309,N_22429);
nor U23503 (N_23503,N_20575,N_20985);
xnor U23504 (N_23504,N_22129,N_22051);
or U23505 (N_23505,N_20121,N_20816);
nor U23506 (N_23506,N_22245,N_20774);
xnor U23507 (N_23507,N_21908,N_21096);
xor U23508 (N_23508,N_21872,N_20560);
nand U23509 (N_23509,N_21110,N_20122);
or U23510 (N_23510,N_20756,N_22348);
nor U23511 (N_23511,N_22088,N_21268);
xnor U23512 (N_23512,N_20555,N_22377);
nand U23513 (N_23513,N_22160,N_21558);
xor U23514 (N_23514,N_22253,N_20055);
xnor U23515 (N_23515,N_20172,N_21767);
nor U23516 (N_23516,N_20230,N_20366);
nor U23517 (N_23517,N_20918,N_22083);
and U23518 (N_23518,N_21320,N_21348);
nor U23519 (N_23519,N_20843,N_21224);
and U23520 (N_23520,N_20453,N_21739);
nor U23521 (N_23521,N_21204,N_20338);
and U23522 (N_23522,N_20182,N_21673);
and U23523 (N_23523,N_22477,N_22165);
nand U23524 (N_23524,N_20429,N_20705);
or U23525 (N_23525,N_21968,N_20507);
nand U23526 (N_23526,N_21551,N_21836);
and U23527 (N_23527,N_22441,N_22236);
nor U23528 (N_23528,N_21016,N_20520);
nor U23529 (N_23529,N_20954,N_21898);
or U23530 (N_23530,N_21020,N_20693);
and U23531 (N_23531,N_22452,N_20341);
and U23532 (N_23532,N_21595,N_21421);
nand U23533 (N_23533,N_21539,N_20999);
and U23534 (N_23534,N_20567,N_20070);
nand U23535 (N_23535,N_21136,N_21557);
nand U23536 (N_23536,N_21367,N_20654);
nand U23537 (N_23537,N_22321,N_22130);
and U23538 (N_23538,N_21641,N_22438);
or U23539 (N_23539,N_21933,N_22234);
nor U23540 (N_23540,N_21600,N_20186);
xor U23541 (N_23541,N_20749,N_20381);
nand U23542 (N_23542,N_20536,N_20281);
nor U23543 (N_23543,N_21586,N_20586);
nand U23544 (N_23544,N_21840,N_20534);
or U23545 (N_23545,N_20600,N_20758);
nor U23546 (N_23546,N_21890,N_21818);
and U23547 (N_23547,N_21849,N_21935);
nor U23548 (N_23548,N_20527,N_22374);
and U23549 (N_23549,N_22070,N_20621);
or U23550 (N_23550,N_21543,N_20074);
nand U23551 (N_23551,N_20942,N_21496);
nand U23552 (N_23552,N_20085,N_20075);
nand U23553 (N_23553,N_20136,N_21834);
nor U23554 (N_23554,N_20934,N_20471);
xnor U23555 (N_23555,N_20885,N_20634);
and U23556 (N_23556,N_20810,N_20668);
or U23557 (N_23557,N_20788,N_21867);
nand U23558 (N_23558,N_20834,N_21481);
nor U23559 (N_23559,N_21967,N_21879);
nor U23560 (N_23560,N_22246,N_22057);
xor U23561 (N_23561,N_22270,N_22315);
xnor U23562 (N_23562,N_21426,N_20474);
nor U23563 (N_23563,N_21334,N_21419);
xnor U23564 (N_23564,N_21647,N_22450);
or U23565 (N_23565,N_22075,N_20718);
nand U23566 (N_23566,N_22294,N_21859);
nor U23567 (N_23567,N_21845,N_21345);
xor U23568 (N_23568,N_21380,N_22472);
and U23569 (N_23569,N_20339,N_20803);
and U23570 (N_23570,N_20325,N_21660);
and U23571 (N_23571,N_22335,N_21045);
or U23572 (N_23572,N_21006,N_20571);
nand U23573 (N_23573,N_21507,N_20916);
or U23574 (N_23574,N_21370,N_21520);
nand U23575 (N_23575,N_22164,N_22252);
xor U23576 (N_23576,N_21192,N_22475);
and U23577 (N_23577,N_20023,N_21584);
nand U23578 (N_23578,N_22351,N_21196);
nor U23579 (N_23579,N_21121,N_21576);
or U23580 (N_23580,N_21729,N_21940);
and U23581 (N_23581,N_21497,N_20426);
nor U23582 (N_23582,N_20663,N_20523);
nor U23583 (N_23583,N_20036,N_20830);
nand U23584 (N_23584,N_20963,N_22341);
nor U23585 (N_23585,N_20212,N_22059);
nand U23586 (N_23586,N_20043,N_20962);
nand U23587 (N_23587,N_20712,N_20850);
nand U23588 (N_23588,N_21652,N_22402);
nand U23589 (N_23589,N_20777,N_20308);
nor U23590 (N_23590,N_22060,N_21080);
or U23591 (N_23591,N_21773,N_20932);
nand U23592 (N_23592,N_21850,N_21488);
or U23593 (N_23593,N_21474,N_21789);
or U23594 (N_23594,N_20670,N_22327);
nor U23595 (N_23595,N_22100,N_20466);
nand U23596 (N_23596,N_21841,N_21936);
nand U23597 (N_23597,N_22263,N_21848);
and U23598 (N_23598,N_20652,N_20165);
or U23599 (N_23599,N_21741,N_20794);
or U23600 (N_23600,N_22388,N_20384);
nand U23601 (N_23601,N_20993,N_22237);
or U23602 (N_23602,N_20849,N_22287);
xnor U23603 (N_23603,N_22366,N_22295);
nand U23604 (N_23604,N_20105,N_21282);
nand U23605 (N_23605,N_20025,N_22029);
nand U23606 (N_23606,N_21162,N_21816);
and U23607 (N_23607,N_22490,N_20856);
nor U23608 (N_23608,N_20083,N_20347);
and U23609 (N_23609,N_21467,N_20602);
and U23610 (N_23610,N_21672,N_22314);
xnor U23611 (N_23611,N_20455,N_22062);
xnor U23612 (N_23612,N_21821,N_20225);
xnor U23613 (N_23613,N_21962,N_20913);
nand U23614 (N_23614,N_20385,N_21115);
nand U23615 (N_23615,N_21592,N_21889);
xnor U23616 (N_23616,N_21605,N_20222);
and U23617 (N_23617,N_20741,N_20316);
nand U23618 (N_23618,N_20817,N_21590);
nor U23619 (N_23619,N_20688,N_22228);
nand U23620 (N_23620,N_20382,N_20979);
xnor U23621 (N_23621,N_22264,N_20728);
xnor U23622 (N_23622,N_21919,N_21529);
and U23623 (N_23623,N_21167,N_20291);
xor U23624 (N_23624,N_20289,N_21686);
xnor U23625 (N_23625,N_20735,N_21732);
or U23626 (N_23626,N_21393,N_22395);
xor U23627 (N_23627,N_20313,N_20058);
and U23628 (N_23628,N_20335,N_22180);
or U23629 (N_23629,N_21356,N_21814);
and U23630 (N_23630,N_21585,N_21717);
xnor U23631 (N_23631,N_20295,N_20350);
nand U23632 (N_23632,N_20389,N_20578);
and U23633 (N_23633,N_21703,N_20056);
nand U23634 (N_23634,N_20469,N_21486);
nand U23635 (N_23635,N_22179,N_20147);
nand U23636 (N_23636,N_20821,N_20646);
and U23637 (N_23637,N_20009,N_20790);
nor U23638 (N_23638,N_20667,N_22242);
nand U23639 (N_23639,N_21400,N_20900);
nand U23640 (N_23640,N_22194,N_22435);
nand U23641 (N_23641,N_20583,N_20479);
xor U23642 (N_23642,N_22359,N_21820);
nor U23643 (N_23643,N_21929,N_20071);
or U23644 (N_23644,N_21870,N_20251);
and U23645 (N_23645,N_20924,N_21637);
and U23646 (N_23646,N_20128,N_20881);
xor U23647 (N_23647,N_22273,N_22337);
xor U23648 (N_23648,N_20348,N_21698);
or U23649 (N_23649,N_21922,N_22406);
nor U23650 (N_23650,N_22400,N_21274);
xor U23651 (N_23651,N_20337,N_21581);
and U23652 (N_23652,N_21143,N_20815);
nor U23653 (N_23653,N_21343,N_22125);
nand U23654 (N_23654,N_20086,N_20235);
xor U23655 (N_23655,N_22109,N_21160);
and U23656 (N_23656,N_20228,N_20854);
and U23657 (N_23657,N_22034,N_22039);
xnor U23658 (N_23658,N_20084,N_20557);
nor U23659 (N_23659,N_21266,N_21803);
nor U23660 (N_23660,N_21381,N_21559);
nand U23661 (N_23661,N_21447,N_22172);
and U23662 (N_23662,N_20676,N_21333);
nand U23663 (N_23663,N_20755,N_20554);
or U23664 (N_23664,N_21957,N_21461);
xor U23665 (N_23665,N_22158,N_21754);
or U23666 (N_23666,N_22249,N_20048);
xor U23667 (N_23667,N_21945,N_20135);
nor U23668 (N_23668,N_21838,N_22023);
and U23669 (N_23669,N_22311,N_20175);
or U23670 (N_23670,N_20596,N_22488);
and U23671 (N_23671,N_22381,N_20459);
or U23672 (N_23672,N_21644,N_21434);
and U23673 (N_23673,N_20877,N_22276);
nor U23674 (N_23674,N_21390,N_20227);
or U23675 (N_23675,N_21865,N_20311);
nand U23676 (N_23676,N_20102,N_20927);
and U23677 (N_23677,N_20402,N_22058);
nor U23678 (N_23678,N_20010,N_20948);
nor U23679 (N_23679,N_22055,N_21842);
and U23680 (N_23680,N_21887,N_20732);
nand U23681 (N_23681,N_20053,N_21990);
or U23682 (N_23682,N_22144,N_20486);
or U23683 (N_23683,N_21691,N_21384);
xnor U23684 (N_23684,N_21174,N_21171);
nor U23685 (N_23685,N_22372,N_22212);
and U23686 (N_23686,N_20532,N_21309);
nand U23687 (N_23687,N_20352,N_22426);
nand U23688 (N_23688,N_22040,N_20260);
and U23689 (N_23689,N_20811,N_20061);
xor U23690 (N_23690,N_20098,N_21593);
nor U23691 (N_23691,N_20953,N_21091);
xnor U23692 (N_23692,N_20687,N_21881);
nand U23693 (N_23693,N_21477,N_21943);
nor U23694 (N_23694,N_22104,N_22342);
and U23695 (N_23695,N_20117,N_22191);
nand U23696 (N_23696,N_21101,N_21550);
nand U23697 (N_23697,N_21372,N_21352);
xnor U23698 (N_23698,N_21407,N_22399);
xor U23699 (N_23699,N_21471,N_21440);
nor U23700 (N_23700,N_20001,N_21992);
xnor U23701 (N_23701,N_21567,N_20801);
xnor U23702 (N_23702,N_20842,N_21534);
xnor U23703 (N_23703,N_20671,N_20656);
nor U23704 (N_23704,N_21123,N_22201);
or U23705 (N_23705,N_20873,N_21130);
nand U23706 (N_23706,N_22305,N_20949);
nand U23707 (N_23707,N_20585,N_20685);
and U23708 (N_23708,N_22002,N_20967);
and U23709 (N_23709,N_20720,N_21705);
and U23710 (N_23710,N_22091,N_20620);
nor U23711 (N_23711,N_21675,N_21403);
or U23712 (N_23712,N_20787,N_20694);
xor U23713 (N_23713,N_20221,N_22089);
nor U23714 (N_23714,N_20521,N_21368);
and U23715 (N_23715,N_21311,N_21187);
or U23716 (N_23716,N_20537,N_21369);
xor U23717 (N_23717,N_20639,N_21901);
nand U23718 (N_23718,N_21643,N_20108);
nand U23719 (N_23719,N_21498,N_20034);
or U23720 (N_23720,N_20014,N_20501);
nor U23721 (N_23721,N_20605,N_20018);
xor U23722 (N_23722,N_21212,N_20006);
nor U23723 (N_23723,N_21280,N_22296);
nand U23724 (N_23724,N_21211,N_21518);
and U23725 (N_23725,N_20959,N_20828);
nand U23726 (N_23726,N_20035,N_22192);
and U23727 (N_23727,N_20439,N_21099);
or U23728 (N_23728,N_22415,N_22407);
xnor U23729 (N_23729,N_20144,N_20892);
nor U23730 (N_23730,N_20808,N_20027);
or U23731 (N_23731,N_21255,N_21740);
and U23732 (N_23732,N_21209,N_21512);
nor U23733 (N_23733,N_21664,N_22369);
nor U23734 (N_23734,N_22316,N_20593);
or U23735 (N_23735,N_20926,N_20373);
nand U23736 (N_23736,N_20247,N_20592);
xor U23737 (N_23737,N_22427,N_21626);
xor U23738 (N_23738,N_21893,N_21942);
and U23739 (N_23739,N_21759,N_20049);
or U23740 (N_23740,N_22309,N_22364);
or U23741 (N_23741,N_20255,N_20574);
and U23742 (N_23742,N_21180,N_22265);
and U23743 (N_23743,N_21594,N_21305);
nand U23744 (N_23744,N_20902,N_21621);
xor U23745 (N_23745,N_20619,N_20077);
and U23746 (N_23746,N_22329,N_22227);
xor U23747 (N_23747,N_21379,N_20432);
xnor U23748 (N_23748,N_20294,N_21681);
nand U23749 (N_23749,N_22171,N_22405);
nor U23750 (N_23750,N_20436,N_21083);
nor U23751 (N_23751,N_21598,N_21657);
and U23752 (N_23752,N_22144,N_20210);
nand U23753 (N_23753,N_20415,N_21004);
nand U23754 (N_23754,N_21035,N_20046);
xor U23755 (N_23755,N_20640,N_20148);
nor U23756 (N_23756,N_21526,N_21878);
or U23757 (N_23757,N_21804,N_20601);
xor U23758 (N_23758,N_21348,N_21958);
or U23759 (N_23759,N_20419,N_20696);
nand U23760 (N_23760,N_20250,N_22010);
nor U23761 (N_23761,N_20994,N_21349);
nand U23762 (N_23762,N_22182,N_22195);
and U23763 (N_23763,N_22031,N_21787);
or U23764 (N_23764,N_21369,N_21691);
xnor U23765 (N_23765,N_20847,N_20706);
or U23766 (N_23766,N_20737,N_21601);
or U23767 (N_23767,N_22158,N_20593);
xor U23768 (N_23768,N_21054,N_21242);
nor U23769 (N_23769,N_22404,N_22479);
and U23770 (N_23770,N_21467,N_20325);
xnor U23771 (N_23771,N_22387,N_20760);
nand U23772 (N_23772,N_21386,N_22227);
nand U23773 (N_23773,N_21013,N_20928);
xnor U23774 (N_23774,N_20674,N_20132);
xnor U23775 (N_23775,N_20735,N_22174);
and U23776 (N_23776,N_21234,N_22278);
xor U23777 (N_23777,N_21503,N_20963);
or U23778 (N_23778,N_20711,N_21826);
and U23779 (N_23779,N_21224,N_21162);
and U23780 (N_23780,N_20463,N_21792);
and U23781 (N_23781,N_20411,N_21556);
xnor U23782 (N_23782,N_20090,N_22023);
or U23783 (N_23783,N_20334,N_20944);
xnor U23784 (N_23784,N_21102,N_20893);
and U23785 (N_23785,N_22075,N_22482);
or U23786 (N_23786,N_20526,N_20776);
xor U23787 (N_23787,N_20874,N_21560);
and U23788 (N_23788,N_22488,N_21395);
nand U23789 (N_23789,N_21741,N_21745);
and U23790 (N_23790,N_21762,N_21514);
nand U23791 (N_23791,N_21906,N_21432);
or U23792 (N_23792,N_21856,N_22122);
nor U23793 (N_23793,N_21410,N_21700);
nand U23794 (N_23794,N_21046,N_20833);
nor U23795 (N_23795,N_21437,N_21661);
and U23796 (N_23796,N_20518,N_20013);
or U23797 (N_23797,N_21974,N_20268);
or U23798 (N_23798,N_20158,N_20387);
xor U23799 (N_23799,N_20504,N_21928);
or U23800 (N_23800,N_20871,N_22282);
nand U23801 (N_23801,N_21543,N_22399);
nor U23802 (N_23802,N_22240,N_21969);
nor U23803 (N_23803,N_21595,N_22376);
nand U23804 (N_23804,N_21597,N_21868);
xor U23805 (N_23805,N_20359,N_20582);
or U23806 (N_23806,N_22184,N_22102);
xnor U23807 (N_23807,N_22071,N_21253);
or U23808 (N_23808,N_20564,N_20454);
or U23809 (N_23809,N_21496,N_21022);
nor U23810 (N_23810,N_21786,N_20093);
nand U23811 (N_23811,N_20098,N_20973);
nand U23812 (N_23812,N_20816,N_20166);
and U23813 (N_23813,N_20997,N_21194);
nor U23814 (N_23814,N_21025,N_20109);
and U23815 (N_23815,N_21519,N_22260);
nor U23816 (N_23816,N_20148,N_21948);
xnor U23817 (N_23817,N_20859,N_20396);
nand U23818 (N_23818,N_22241,N_21430);
or U23819 (N_23819,N_21106,N_20267);
nand U23820 (N_23820,N_20396,N_20160);
nor U23821 (N_23821,N_21003,N_21901);
xnor U23822 (N_23822,N_21007,N_20044);
nand U23823 (N_23823,N_20272,N_20763);
nand U23824 (N_23824,N_21594,N_21069);
nor U23825 (N_23825,N_21619,N_20457);
or U23826 (N_23826,N_21146,N_20102);
and U23827 (N_23827,N_21227,N_20628);
or U23828 (N_23828,N_20037,N_20554);
and U23829 (N_23829,N_21290,N_21151);
and U23830 (N_23830,N_21561,N_22406);
or U23831 (N_23831,N_20466,N_21503);
or U23832 (N_23832,N_20975,N_20364);
xor U23833 (N_23833,N_21452,N_22030);
xor U23834 (N_23834,N_22303,N_22352);
nor U23835 (N_23835,N_20751,N_20214);
nand U23836 (N_23836,N_22346,N_20759);
and U23837 (N_23837,N_21772,N_22405);
nand U23838 (N_23838,N_20298,N_21862);
or U23839 (N_23839,N_22002,N_21314);
nor U23840 (N_23840,N_20629,N_20899);
xor U23841 (N_23841,N_20887,N_20866);
nand U23842 (N_23842,N_21977,N_22024);
or U23843 (N_23843,N_20123,N_21672);
nand U23844 (N_23844,N_21437,N_22001);
nand U23845 (N_23845,N_22098,N_20750);
nor U23846 (N_23846,N_21408,N_20762);
xor U23847 (N_23847,N_20392,N_22430);
xnor U23848 (N_23848,N_20732,N_21189);
nor U23849 (N_23849,N_21865,N_21857);
nor U23850 (N_23850,N_20955,N_20443);
nand U23851 (N_23851,N_20102,N_20819);
nor U23852 (N_23852,N_20777,N_21262);
or U23853 (N_23853,N_21230,N_21857);
nand U23854 (N_23854,N_20920,N_20578);
or U23855 (N_23855,N_21040,N_21128);
or U23856 (N_23856,N_22205,N_20132);
nand U23857 (N_23857,N_21115,N_20124);
nor U23858 (N_23858,N_20715,N_21584);
xnor U23859 (N_23859,N_21445,N_20021);
nor U23860 (N_23860,N_20492,N_20534);
nand U23861 (N_23861,N_21444,N_21873);
xor U23862 (N_23862,N_22095,N_21990);
xor U23863 (N_23863,N_20767,N_21999);
and U23864 (N_23864,N_21383,N_22312);
or U23865 (N_23865,N_20924,N_21029);
xnor U23866 (N_23866,N_22342,N_21114);
or U23867 (N_23867,N_20513,N_20576);
nand U23868 (N_23868,N_20582,N_20706);
nor U23869 (N_23869,N_20236,N_21711);
xor U23870 (N_23870,N_22238,N_20876);
xnor U23871 (N_23871,N_21259,N_22161);
nor U23872 (N_23872,N_20610,N_20662);
and U23873 (N_23873,N_20100,N_20999);
or U23874 (N_23874,N_20156,N_21914);
xor U23875 (N_23875,N_20263,N_21389);
and U23876 (N_23876,N_21556,N_21395);
nor U23877 (N_23877,N_21689,N_20903);
and U23878 (N_23878,N_21561,N_22185);
nand U23879 (N_23879,N_21602,N_22320);
and U23880 (N_23880,N_21675,N_21773);
xnor U23881 (N_23881,N_21911,N_20082);
and U23882 (N_23882,N_20062,N_22428);
or U23883 (N_23883,N_20345,N_22180);
nand U23884 (N_23884,N_20580,N_20581);
nor U23885 (N_23885,N_20653,N_20329);
xor U23886 (N_23886,N_21890,N_20379);
and U23887 (N_23887,N_20420,N_21644);
nor U23888 (N_23888,N_20787,N_20458);
and U23889 (N_23889,N_21659,N_22335);
xnor U23890 (N_23890,N_22479,N_21116);
and U23891 (N_23891,N_20352,N_22392);
nor U23892 (N_23892,N_20809,N_20808);
nand U23893 (N_23893,N_20420,N_22210);
and U23894 (N_23894,N_21166,N_22191);
and U23895 (N_23895,N_20439,N_20893);
or U23896 (N_23896,N_21439,N_20532);
xor U23897 (N_23897,N_20647,N_20364);
xnor U23898 (N_23898,N_20922,N_21191);
and U23899 (N_23899,N_20180,N_20761);
xnor U23900 (N_23900,N_21809,N_20357);
and U23901 (N_23901,N_21781,N_21303);
and U23902 (N_23902,N_20768,N_20945);
nor U23903 (N_23903,N_20437,N_21606);
nor U23904 (N_23904,N_20003,N_20065);
or U23905 (N_23905,N_21591,N_20901);
nand U23906 (N_23906,N_20703,N_20081);
nor U23907 (N_23907,N_20044,N_20505);
or U23908 (N_23908,N_20868,N_21022);
and U23909 (N_23909,N_22443,N_20618);
and U23910 (N_23910,N_20074,N_21127);
or U23911 (N_23911,N_21075,N_20283);
nand U23912 (N_23912,N_20651,N_22365);
nand U23913 (N_23913,N_20137,N_20545);
nor U23914 (N_23914,N_22473,N_20623);
nand U23915 (N_23915,N_20863,N_22382);
xor U23916 (N_23916,N_21848,N_22318);
xor U23917 (N_23917,N_20778,N_21258);
xor U23918 (N_23918,N_22033,N_21982);
xor U23919 (N_23919,N_21794,N_21880);
nand U23920 (N_23920,N_21426,N_21567);
xnor U23921 (N_23921,N_21425,N_20775);
xor U23922 (N_23922,N_21682,N_20522);
xor U23923 (N_23923,N_21488,N_20616);
or U23924 (N_23924,N_20167,N_21646);
nor U23925 (N_23925,N_20978,N_21793);
and U23926 (N_23926,N_22018,N_20630);
and U23927 (N_23927,N_20320,N_21540);
nand U23928 (N_23928,N_22436,N_20714);
and U23929 (N_23929,N_22067,N_20495);
xnor U23930 (N_23930,N_20423,N_20404);
nor U23931 (N_23931,N_20949,N_21507);
xor U23932 (N_23932,N_20048,N_21818);
or U23933 (N_23933,N_22415,N_22432);
and U23934 (N_23934,N_20650,N_20835);
nand U23935 (N_23935,N_21636,N_20545);
and U23936 (N_23936,N_20745,N_20346);
and U23937 (N_23937,N_21132,N_21356);
nor U23938 (N_23938,N_20725,N_21717);
nor U23939 (N_23939,N_20179,N_21065);
nand U23940 (N_23940,N_21370,N_21274);
nand U23941 (N_23941,N_20598,N_21494);
xor U23942 (N_23942,N_21200,N_20184);
and U23943 (N_23943,N_20550,N_20754);
nand U23944 (N_23944,N_20128,N_21967);
and U23945 (N_23945,N_22300,N_21744);
xor U23946 (N_23946,N_21267,N_21062);
or U23947 (N_23947,N_20024,N_21251);
nand U23948 (N_23948,N_21755,N_21604);
and U23949 (N_23949,N_21510,N_21818);
nand U23950 (N_23950,N_21336,N_20453);
xnor U23951 (N_23951,N_20181,N_20276);
nor U23952 (N_23952,N_20247,N_20052);
and U23953 (N_23953,N_22452,N_22231);
nor U23954 (N_23954,N_21860,N_20448);
nand U23955 (N_23955,N_21631,N_22067);
or U23956 (N_23956,N_21291,N_22399);
and U23957 (N_23957,N_21431,N_20875);
nand U23958 (N_23958,N_22276,N_20444);
nand U23959 (N_23959,N_21760,N_22079);
nor U23960 (N_23960,N_20333,N_21689);
nand U23961 (N_23961,N_22258,N_20626);
xnor U23962 (N_23962,N_20724,N_22185);
or U23963 (N_23963,N_21270,N_20469);
xor U23964 (N_23964,N_22094,N_21820);
xor U23965 (N_23965,N_21576,N_22126);
nor U23966 (N_23966,N_22100,N_20204);
and U23967 (N_23967,N_20014,N_21417);
nor U23968 (N_23968,N_21979,N_21294);
or U23969 (N_23969,N_20106,N_20986);
xor U23970 (N_23970,N_20985,N_20257);
nor U23971 (N_23971,N_20900,N_20444);
xor U23972 (N_23972,N_21237,N_20981);
and U23973 (N_23973,N_21201,N_21681);
nor U23974 (N_23974,N_21011,N_20252);
or U23975 (N_23975,N_20011,N_21376);
nor U23976 (N_23976,N_21720,N_20369);
xnor U23977 (N_23977,N_20448,N_20694);
xnor U23978 (N_23978,N_22078,N_20001);
xnor U23979 (N_23979,N_21202,N_20459);
and U23980 (N_23980,N_20288,N_20190);
or U23981 (N_23981,N_22065,N_20454);
xnor U23982 (N_23982,N_20397,N_21933);
xor U23983 (N_23983,N_20914,N_22490);
nand U23984 (N_23984,N_22061,N_21873);
nand U23985 (N_23985,N_22170,N_22050);
xnor U23986 (N_23986,N_22017,N_21616);
and U23987 (N_23987,N_21220,N_21983);
nor U23988 (N_23988,N_20675,N_20506);
and U23989 (N_23989,N_21483,N_21506);
nand U23990 (N_23990,N_22104,N_22463);
or U23991 (N_23991,N_21332,N_20244);
and U23992 (N_23992,N_21986,N_21804);
nand U23993 (N_23993,N_22377,N_21864);
nor U23994 (N_23994,N_20795,N_20056);
or U23995 (N_23995,N_20888,N_21564);
and U23996 (N_23996,N_20120,N_20572);
or U23997 (N_23997,N_21025,N_21492);
xor U23998 (N_23998,N_21798,N_22058);
nand U23999 (N_23999,N_20941,N_20428);
xnor U24000 (N_24000,N_21731,N_20203);
and U24001 (N_24001,N_20387,N_20153);
nor U24002 (N_24002,N_21053,N_21677);
nor U24003 (N_24003,N_21777,N_21349);
xnor U24004 (N_24004,N_20186,N_20307);
xnor U24005 (N_24005,N_22338,N_20560);
nand U24006 (N_24006,N_21240,N_22452);
xnor U24007 (N_24007,N_21752,N_22441);
and U24008 (N_24008,N_21285,N_22430);
and U24009 (N_24009,N_21252,N_21640);
and U24010 (N_24010,N_21158,N_20259);
nand U24011 (N_24011,N_21868,N_22055);
nand U24012 (N_24012,N_21437,N_20931);
and U24013 (N_24013,N_20127,N_22275);
nand U24014 (N_24014,N_20289,N_21808);
xor U24015 (N_24015,N_21308,N_22177);
xor U24016 (N_24016,N_22426,N_22496);
nor U24017 (N_24017,N_21593,N_22035);
or U24018 (N_24018,N_21625,N_20406);
nor U24019 (N_24019,N_21661,N_22017);
nand U24020 (N_24020,N_22391,N_21123);
and U24021 (N_24021,N_20389,N_21353);
nor U24022 (N_24022,N_20941,N_20917);
and U24023 (N_24023,N_21559,N_20797);
nor U24024 (N_24024,N_22278,N_21849);
and U24025 (N_24025,N_20556,N_22131);
nand U24026 (N_24026,N_20743,N_22189);
and U24027 (N_24027,N_20167,N_21139);
and U24028 (N_24028,N_20057,N_20335);
nor U24029 (N_24029,N_21944,N_21702);
or U24030 (N_24030,N_21803,N_21196);
or U24031 (N_24031,N_21313,N_22249);
nor U24032 (N_24032,N_21131,N_21780);
xor U24033 (N_24033,N_20546,N_21007);
xor U24034 (N_24034,N_21798,N_21138);
and U24035 (N_24035,N_20404,N_21327);
nor U24036 (N_24036,N_21194,N_20447);
nand U24037 (N_24037,N_20167,N_21103);
xor U24038 (N_24038,N_20587,N_21437);
or U24039 (N_24039,N_21834,N_20636);
or U24040 (N_24040,N_22364,N_21710);
and U24041 (N_24041,N_21944,N_20917);
nand U24042 (N_24042,N_21409,N_21331);
or U24043 (N_24043,N_21075,N_20995);
xor U24044 (N_24044,N_21893,N_21253);
nand U24045 (N_24045,N_21705,N_22286);
and U24046 (N_24046,N_20249,N_20926);
xnor U24047 (N_24047,N_21401,N_21430);
xor U24048 (N_24048,N_20905,N_20045);
and U24049 (N_24049,N_21297,N_20736);
or U24050 (N_24050,N_21887,N_21513);
nor U24051 (N_24051,N_22199,N_20211);
nand U24052 (N_24052,N_20294,N_20668);
nor U24053 (N_24053,N_20267,N_20927);
xnor U24054 (N_24054,N_22466,N_21531);
nor U24055 (N_24055,N_21106,N_21309);
and U24056 (N_24056,N_22369,N_22079);
or U24057 (N_24057,N_21749,N_22440);
nor U24058 (N_24058,N_20333,N_22275);
xor U24059 (N_24059,N_22029,N_22359);
xnor U24060 (N_24060,N_22465,N_21093);
xor U24061 (N_24061,N_20285,N_21037);
or U24062 (N_24062,N_20881,N_20002);
and U24063 (N_24063,N_20570,N_21183);
nand U24064 (N_24064,N_21100,N_20014);
xor U24065 (N_24065,N_21823,N_22436);
nand U24066 (N_24066,N_22390,N_20832);
nand U24067 (N_24067,N_20871,N_20682);
or U24068 (N_24068,N_20692,N_22479);
or U24069 (N_24069,N_20917,N_22003);
and U24070 (N_24070,N_22087,N_22407);
or U24071 (N_24071,N_20347,N_20837);
nand U24072 (N_24072,N_20094,N_21117);
or U24073 (N_24073,N_21158,N_21319);
nand U24074 (N_24074,N_20815,N_21606);
and U24075 (N_24075,N_22318,N_22276);
xor U24076 (N_24076,N_22378,N_20684);
and U24077 (N_24077,N_20546,N_22002);
and U24078 (N_24078,N_20454,N_21125);
or U24079 (N_24079,N_21701,N_21715);
nor U24080 (N_24080,N_20408,N_20226);
and U24081 (N_24081,N_20874,N_21383);
nor U24082 (N_24082,N_20778,N_20355);
xor U24083 (N_24083,N_21129,N_22444);
xor U24084 (N_24084,N_21127,N_22041);
and U24085 (N_24085,N_20642,N_20467);
or U24086 (N_24086,N_21954,N_22464);
nor U24087 (N_24087,N_20555,N_21662);
xor U24088 (N_24088,N_20603,N_22139);
nor U24089 (N_24089,N_20616,N_22281);
and U24090 (N_24090,N_21866,N_22472);
xor U24091 (N_24091,N_20799,N_21935);
and U24092 (N_24092,N_20207,N_20054);
nand U24093 (N_24093,N_20365,N_21302);
nand U24094 (N_24094,N_20419,N_20912);
or U24095 (N_24095,N_21890,N_20473);
or U24096 (N_24096,N_20586,N_20049);
nand U24097 (N_24097,N_21629,N_20722);
nor U24098 (N_24098,N_21674,N_20474);
nand U24099 (N_24099,N_20622,N_20634);
nand U24100 (N_24100,N_21974,N_21370);
xnor U24101 (N_24101,N_20982,N_20432);
or U24102 (N_24102,N_21842,N_21976);
nor U24103 (N_24103,N_22403,N_21582);
nor U24104 (N_24104,N_21882,N_20682);
and U24105 (N_24105,N_22335,N_21507);
nand U24106 (N_24106,N_21418,N_22392);
and U24107 (N_24107,N_22460,N_21501);
and U24108 (N_24108,N_20265,N_20320);
and U24109 (N_24109,N_22241,N_22182);
nor U24110 (N_24110,N_20374,N_21101);
xnor U24111 (N_24111,N_21747,N_22137);
nor U24112 (N_24112,N_20015,N_21089);
or U24113 (N_24113,N_20664,N_22334);
or U24114 (N_24114,N_21267,N_21194);
nor U24115 (N_24115,N_21958,N_20116);
or U24116 (N_24116,N_21562,N_22345);
and U24117 (N_24117,N_21006,N_20520);
or U24118 (N_24118,N_20111,N_21963);
xnor U24119 (N_24119,N_20933,N_22065);
xnor U24120 (N_24120,N_20747,N_21334);
and U24121 (N_24121,N_21097,N_22078);
nor U24122 (N_24122,N_22398,N_21972);
nor U24123 (N_24123,N_22331,N_22313);
nor U24124 (N_24124,N_21112,N_20809);
nor U24125 (N_24125,N_20842,N_20560);
xor U24126 (N_24126,N_21864,N_20506);
and U24127 (N_24127,N_20284,N_21523);
nor U24128 (N_24128,N_21113,N_20604);
and U24129 (N_24129,N_22484,N_21160);
nor U24130 (N_24130,N_22441,N_20434);
and U24131 (N_24131,N_20947,N_21292);
nand U24132 (N_24132,N_21668,N_21899);
nor U24133 (N_24133,N_21467,N_21807);
or U24134 (N_24134,N_22274,N_21709);
nor U24135 (N_24135,N_20069,N_20033);
or U24136 (N_24136,N_21571,N_21644);
nand U24137 (N_24137,N_20423,N_22083);
xor U24138 (N_24138,N_21324,N_20903);
and U24139 (N_24139,N_20624,N_22069);
nor U24140 (N_24140,N_21835,N_20837);
xnor U24141 (N_24141,N_22241,N_20537);
and U24142 (N_24142,N_20093,N_20303);
and U24143 (N_24143,N_20186,N_21154);
nand U24144 (N_24144,N_22380,N_20848);
nor U24145 (N_24145,N_20244,N_20670);
xor U24146 (N_24146,N_20246,N_21686);
nand U24147 (N_24147,N_21452,N_20132);
or U24148 (N_24148,N_22469,N_21493);
nor U24149 (N_24149,N_21111,N_21004);
nor U24150 (N_24150,N_20796,N_21051);
or U24151 (N_24151,N_22209,N_22481);
and U24152 (N_24152,N_21110,N_21153);
nor U24153 (N_24153,N_20076,N_20057);
or U24154 (N_24154,N_21691,N_21143);
nor U24155 (N_24155,N_22285,N_20581);
and U24156 (N_24156,N_21076,N_20683);
nand U24157 (N_24157,N_22275,N_21073);
nand U24158 (N_24158,N_21624,N_20927);
nor U24159 (N_24159,N_20370,N_20366);
nor U24160 (N_24160,N_22241,N_20803);
and U24161 (N_24161,N_20296,N_20683);
xnor U24162 (N_24162,N_21562,N_20677);
nand U24163 (N_24163,N_20788,N_21455);
or U24164 (N_24164,N_21427,N_20858);
nand U24165 (N_24165,N_20443,N_22325);
or U24166 (N_24166,N_21354,N_21065);
xnor U24167 (N_24167,N_21606,N_20935);
nor U24168 (N_24168,N_20776,N_21667);
or U24169 (N_24169,N_21423,N_20192);
nor U24170 (N_24170,N_20059,N_20265);
nand U24171 (N_24171,N_21070,N_20465);
nor U24172 (N_24172,N_20343,N_21890);
nand U24173 (N_24173,N_21062,N_22437);
and U24174 (N_24174,N_22340,N_20659);
or U24175 (N_24175,N_20009,N_22124);
and U24176 (N_24176,N_22104,N_22368);
nand U24177 (N_24177,N_22284,N_20526);
and U24178 (N_24178,N_20291,N_20345);
nand U24179 (N_24179,N_21734,N_22461);
and U24180 (N_24180,N_20333,N_20085);
nor U24181 (N_24181,N_22376,N_20419);
xnor U24182 (N_24182,N_22219,N_21058);
nor U24183 (N_24183,N_21585,N_22084);
xnor U24184 (N_24184,N_21755,N_20240);
nand U24185 (N_24185,N_22120,N_21522);
nor U24186 (N_24186,N_20744,N_20871);
or U24187 (N_24187,N_20029,N_20296);
nand U24188 (N_24188,N_21278,N_22413);
or U24189 (N_24189,N_21271,N_21765);
nand U24190 (N_24190,N_21015,N_20229);
and U24191 (N_24191,N_21330,N_20254);
and U24192 (N_24192,N_20551,N_20870);
or U24193 (N_24193,N_20496,N_21093);
xnor U24194 (N_24194,N_21676,N_21749);
nand U24195 (N_24195,N_21093,N_21675);
xor U24196 (N_24196,N_22309,N_20587);
and U24197 (N_24197,N_21193,N_21727);
and U24198 (N_24198,N_21380,N_22454);
xor U24199 (N_24199,N_22010,N_22455);
nor U24200 (N_24200,N_21221,N_20266);
and U24201 (N_24201,N_20448,N_21059);
nand U24202 (N_24202,N_20019,N_21841);
or U24203 (N_24203,N_21745,N_21815);
xnor U24204 (N_24204,N_20694,N_21860);
or U24205 (N_24205,N_21469,N_21758);
nand U24206 (N_24206,N_22106,N_20447);
nor U24207 (N_24207,N_20396,N_21786);
nor U24208 (N_24208,N_21207,N_22156);
nand U24209 (N_24209,N_20991,N_20016);
nor U24210 (N_24210,N_22431,N_21272);
nand U24211 (N_24211,N_20189,N_20080);
xor U24212 (N_24212,N_21430,N_20450);
or U24213 (N_24213,N_22302,N_22231);
xnor U24214 (N_24214,N_21615,N_20200);
nand U24215 (N_24215,N_21588,N_21051);
or U24216 (N_24216,N_21127,N_21659);
or U24217 (N_24217,N_22406,N_20590);
nand U24218 (N_24218,N_20465,N_22041);
and U24219 (N_24219,N_20603,N_20113);
nand U24220 (N_24220,N_21206,N_20922);
and U24221 (N_24221,N_20737,N_22459);
nand U24222 (N_24222,N_21781,N_22354);
and U24223 (N_24223,N_20780,N_20020);
and U24224 (N_24224,N_21287,N_20644);
xnor U24225 (N_24225,N_21315,N_20964);
nand U24226 (N_24226,N_20718,N_21018);
or U24227 (N_24227,N_21135,N_22374);
nand U24228 (N_24228,N_20294,N_20330);
nand U24229 (N_24229,N_20713,N_22347);
or U24230 (N_24230,N_22368,N_20355);
and U24231 (N_24231,N_20726,N_22072);
xnor U24232 (N_24232,N_22309,N_20521);
or U24233 (N_24233,N_22231,N_20581);
xnor U24234 (N_24234,N_22289,N_20029);
xnor U24235 (N_24235,N_20374,N_22313);
or U24236 (N_24236,N_22497,N_20283);
and U24237 (N_24237,N_20439,N_21955);
and U24238 (N_24238,N_20970,N_21424);
and U24239 (N_24239,N_22138,N_20655);
nand U24240 (N_24240,N_22099,N_21544);
and U24241 (N_24241,N_21086,N_20263);
xnor U24242 (N_24242,N_21355,N_22265);
or U24243 (N_24243,N_21975,N_21430);
nor U24244 (N_24244,N_22175,N_22249);
or U24245 (N_24245,N_21894,N_21855);
xor U24246 (N_24246,N_21926,N_22423);
and U24247 (N_24247,N_21935,N_22159);
nand U24248 (N_24248,N_21057,N_20990);
and U24249 (N_24249,N_20945,N_21480);
nor U24250 (N_24250,N_21909,N_22090);
nand U24251 (N_24251,N_21565,N_21772);
or U24252 (N_24252,N_21831,N_21170);
nor U24253 (N_24253,N_20075,N_20101);
nand U24254 (N_24254,N_21718,N_22485);
nand U24255 (N_24255,N_22335,N_20471);
or U24256 (N_24256,N_22426,N_21190);
xor U24257 (N_24257,N_22092,N_22211);
xor U24258 (N_24258,N_20777,N_20804);
nor U24259 (N_24259,N_20811,N_22397);
nand U24260 (N_24260,N_21918,N_21161);
or U24261 (N_24261,N_22210,N_21488);
and U24262 (N_24262,N_20901,N_21432);
xnor U24263 (N_24263,N_20165,N_22043);
and U24264 (N_24264,N_21313,N_22361);
and U24265 (N_24265,N_21775,N_21854);
or U24266 (N_24266,N_21428,N_20227);
nand U24267 (N_24267,N_22077,N_20882);
nor U24268 (N_24268,N_21111,N_22355);
nor U24269 (N_24269,N_21150,N_20170);
xnor U24270 (N_24270,N_21001,N_22108);
and U24271 (N_24271,N_20292,N_22270);
xor U24272 (N_24272,N_20913,N_20244);
nand U24273 (N_24273,N_21896,N_20132);
and U24274 (N_24274,N_21557,N_22077);
and U24275 (N_24275,N_22107,N_22131);
or U24276 (N_24276,N_20487,N_22370);
nand U24277 (N_24277,N_22174,N_21454);
nor U24278 (N_24278,N_21823,N_22421);
nor U24279 (N_24279,N_21959,N_22230);
or U24280 (N_24280,N_22085,N_22239);
or U24281 (N_24281,N_21268,N_20779);
and U24282 (N_24282,N_20749,N_22033);
nand U24283 (N_24283,N_21281,N_21105);
or U24284 (N_24284,N_21146,N_21609);
and U24285 (N_24285,N_20503,N_21656);
and U24286 (N_24286,N_21026,N_20440);
xnor U24287 (N_24287,N_21543,N_22479);
nand U24288 (N_24288,N_22286,N_20386);
or U24289 (N_24289,N_20410,N_22077);
xor U24290 (N_24290,N_22032,N_21916);
nand U24291 (N_24291,N_21253,N_21421);
xor U24292 (N_24292,N_22267,N_21242);
and U24293 (N_24293,N_21800,N_21609);
and U24294 (N_24294,N_20529,N_20922);
and U24295 (N_24295,N_20814,N_20445);
nor U24296 (N_24296,N_22167,N_22352);
nand U24297 (N_24297,N_22114,N_20939);
xor U24298 (N_24298,N_21766,N_22173);
nor U24299 (N_24299,N_21307,N_20827);
nand U24300 (N_24300,N_20175,N_21751);
and U24301 (N_24301,N_20808,N_22489);
xor U24302 (N_24302,N_22166,N_20470);
nor U24303 (N_24303,N_21376,N_20353);
xor U24304 (N_24304,N_22055,N_20249);
nand U24305 (N_24305,N_21684,N_21876);
nor U24306 (N_24306,N_21047,N_20720);
xor U24307 (N_24307,N_21876,N_21780);
or U24308 (N_24308,N_20928,N_22122);
nand U24309 (N_24309,N_22200,N_20126);
and U24310 (N_24310,N_20856,N_21250);
nor U24311 (N_24311,N_20668,N_22002);
nand U24312 (N_24312,N_22335,N_22374);
xor U24313 (N_24313,N_21157,N_21292);
nor U24314 (N_24314,N_20175,N_21199);
and U24315 (N_24315,N_21341,N_20528);
and U24316 (N_24316,N_21936,N_22272);
nand U24317 (N_24317,N_20464,N_20248);
nand U24318 (N_24318,N_20689,N_21161);
or U24319 (N_24319,N_20059,N_21219);
and U24320 (N_24320,N_20636,N_22003);
xnor U24321 (N_24321,N_21736,N_21641);
nor U24322 (N_24322,N_21880,N_20283);
and U24323 (N_24323,N_20941,N_21748);
nand U24324 (N_24324,N_21004,N_22495);
or U24325 (N_24325,N_20586,N_20198);
nor U24326 (N_24326,N_20266,N_21671);
or U24327 (N_24327,N_22498,N_22265);
and U24328 (N_24328,N_20560,N_20092);
or U24329 (N_24329,N_20171,N_22230);
nand U24330 (N_24330,N_20055,N_20668);
nor U24331 (N_24331,N_21762,N_21265);
nor U24332 (N_24332,N_20090,N_20653);
and U24333 (N_24333,N_20346,N_20746);
xor U24334 (N_24334,N_21929,N_20408);
xor U24335 (N_24335,N_20046,N_20508);
and U24336 (N_24336,N_22312,N_21665);
xnor U24337 (N_24337,N_22375,N_21697);
and U24338 (N_24338,N_20972,N_21570);
xnor U24339 (N_24339,N_20139,N_21525);
xnor U24340 (N_24340,N_20228,N_20694);
xnor U24341 (N_24341,N_21441,N_21060);
or U24342 (N_24342,N_20534,N_20338);
xnor U24343 (N_24343,N_20213,N_21486);
xnor U24344 (N_24344,N_20363,N_20356);
nor U24345 (N_24345,N_21745,N_21812);
or U24346 (N_24346,N_21994,N_20051);
and U24347 (N_24347,N_22448,N_21011);
and U24348 (N_24348,N_20941,N_20558);
or U24349 (N_24349,N_20479,N_20380);
and U24350 (N_24350,N_20505,N_20723);
or U24351 (N_24351,N_21324,N_21528);
or U24352 (N_24352,N_21989,N_21142);
and U24353 (N_24353,N_20850,N_20600);
and U24354 (N_24354,N_20721,N_21259);
xor U24355 (N_24355,N_21724,N_20116);
nor U24356 (N_24356,N_20092,N_21940);
nor U24357 (N_24357,N_21369,N_20913);
xnor U24358 (N_24358,N_22104,N_22493);
xor U24359 (N_24359,N_20090,N_21957);
nand U24360 (N_24360,N_21626,N_22401);
or U24361 (N_24361,N_20651,N_21173);
nand U24362 (N_24362,N_21881,N_21537);
xnor U24363 (N_24363,N_22250,N_22111);
nand U24364 (N_24364,N_22419,N_20783);
xor U24365 (N_24365,N_20306,N_21856);
or U24366 (N_24366,N_20673,N_21181);
nand U24367 (N_24367,N_20798,N_22089);
xor U24368 (N_24368,N_22250,N_21529);
or U24369 (N_24369,N_22155,N_21596);
xor U24370 (N_24370,N_21028,N_21227);
or U24371 (N_24371,N_20669,N_22041);
nand U24372 (N_24372,N_22238,N_20711);
nor U24373 (N_24373,N_21437,N_20262);
nand U24374 (N_24374,N_21323,N_22475);
and U24375 (N_24375,N_20290,N_20422);
and U24376 (N_24376,N_22188,N_22424);
xnor U24377 (N_24377,N_21066,N_22145);
or U24378 (N_24378,N_21064,N_20973);
nor U24379 (N_24379,N_20476,N_20683);
xnor U24380 (N_24380,N_21001,N_21498);
and U24381 (N_24381,N_22114,N_21421);
xnor U24382 (N_24382,N_21002,N_20791);
and U24383 (N_24383,N_21348,N_20934);
nor U24384 (N_24384,N_20016,N_20350);
nand U24385 (N_24385,N_21639,N_20840);
nor U24386 (N_24386,N_21655,N_20871);
nor U24387 (N_24387,N_20571,N_20484);
or U24388 (N_24388,N_21568,N_21001);
and U24389 (N_24389,N_21621,N_22356);
nand U24390 (N_24390,N_20629,N_20566);
and U24391 (N_24391,N_20232,N_20766);
xnor U24392 (N_24392,N_22461,N_20785);
and U24393 (N_24393,N_20272,N_20237);
or U24394 (N_24394,N_20663,N_22252);
nor U24395 (N_24395,N_21985,N_20651);
nand U24396 (N_24396,N_21356,N_20771);
and U24397 (N_24397,N_21701,N_20874);
xnor U24398 (N_24398,N_22423,N_21614);
nor U24399 (N_24399,N_22398,N_20406);
xor U24400 (N_24400,N_20613,N_21144);
nand U24401 (N_24401,N_20369,N_20060);
and U24402 (N_24402,N_21691,N_20695);
or U24403 (N_24403,N_22006,N_20919);
nand U24404 (N_24404,N_21179,N_21318);
xor U24405 (N_24405,N_22139,N_22318);
nor U24406 (N_24406,N_20820,N_20575);
nor U24407 (N_24407,N_22101,N_21416);
nor U24408 (N_24408,N_20577,N_21745);
nor U24409 (N_24409,N_22489,N_20903);
xor U24410 (N_24410,N_21884,N_21185);
xor U24411 (N_24411,N_21355,N_21962);
or U24412 (N_24412,N_21389,N_21013);
xor U24413 (N_24413,N_20226,N_21995);
nor U24414 (N_24414,N_20804,N_21369);
nor U24415 (N_24415,N_21279,N_20433);
or U24416 (N_24416,N_20921,N_22113);
nand U24417 (N_24417,N_21904,N_22344);
nand U24418 (N_24418,N_21729,N_21397);
nand U24419 (N_24419,N_20933,N_20848);
xnor U24420 (N_24420,N_22340,N_20772);
nor U24421 (N_24421,N_21543,N_20618);
and U24422 (N_24422,N_21304,N_20977);
nor U24423 (N_24423,N_21806,N_20994);
xor U24424 (N_24424,N_21724,N_22096);
nand U24425 (N_24425,N_21567,N_22229);
nor U24426 (N_24426,N_22098,N_20316);
xor U24427 (N_24427,N_20311,N_20410);
nor U24428 (N_24428,N_20518,N_20411);
nor U24429 (N_24429,N_21979,N_20302);
nor U24430 (N_24430,N_20280,N_20736);
and U24431 (N_24431,N_20607,N_20838);
or U24432 (N_24432,N_20767,N_20895);
or U24433 (N_24433,N_20241,N_20553);
or U24434 (N_24434,N_21829,N_21557);
nor U24435 (N_24435,N_20663,N_21938);
or U24436 (N_24436,N_20742,N_21572);
xor U24437 (N_24437,N_20714,N_21011);
or U24438 (N_24438,N_21439,N_20034);
nor U24439 (N_24439,N_21416,N_20342);
xor U24440 (N_24440,N_20497,N_21419);
nor U24441 (N_24441,N_21166,N_21404);
and U24442 (N_24442,N_22202,N_21215);
and U24443 (N_24443,N_21934,N_22473);
xnor U24444 (N_24444,N_21194,N_21233);
or U24445 (N_24445,N_20625,N_21586);
nor U24446 (N_24446,N_20808,N_22399);
and U24447 (N_24447,N_22254,N_20767);
or U24448 (N_24448,N_22413,N_20089);
xnor U24449 (N_24449,N_20979,N_20640);
and U24450 (N_24450,N_21530,N_20027);
nor U24451 (N_24451,N_21575,N_22470);
xor U24452 (N_24452,N_21999,N_20119);
xnor U24453 (N_24453,N_21725,N_21055);
or U24454 (N_24454,N_22259,N_20236);
or U24455 (N_24455,N_20891,N_22037);
or U24456 (N_24456,N_21511,N_20634);
xnor U24457 (N_24457,N_20943,N_21304);
nand U24458 (N_24458,N_20415,N_21179);
or U24459 (N_24459,N_22256,N_20695);
nand U24460 (N_24460,N_21956,N_21995);
nor U24461 (N_24461,N_21049,N_20062);
and U24462 (N_24462,N_22364,N_20325);
and U24463 (N_24463,N_21039,N_21495);
or U24464 (N_24464,N_22440,N_20836);
or U24465 (N_24465,N_22235,N_21555);
and U24466 (N_24466,N_21400,N_20765);
nand U24467 (N_24467,N_21835,N_20505);
or U24468 (N_24468,N_22008,N_21313);
and U24469 (N_24469,N_20082,N_21583);
xor U24470 (N_24470,N_21450,N_20043);
nor U24471 (N_24471,N_22127,N_22359);
nor U24472 (N_24472,N_22391,N_21510);
xnor U24473 (N_24473,N_21066,N_21635);
or U24474 (N_24474,N_21469,N_21700);
nand U24475 (N_24475,N_20625,N_20558);
and U24476 (N_24476,N_20700,N_21173);
nand U24477 (N_24477,N_21492,N_20745);
nor U24478 (N_24478,N_20586,N_22405);
and U24479 (N_24479,N_21924,N_20023);
or U24480 (N_24480,N_22484,N_20444);
or U24481 (N_24481,N_22127,N_21555);
xnor U24482 (N_24482,N_21943,N_21199);
xnor U24483 (N_24483,N_20320,N_20524);
nand U24484 (N_24484,N_22176,N_22084);
nand U24485 (N_24485,N_20212,N_21844);
nor U24486 (N_24486,N_20192,N_21037);
xor U24487 (N_24487,N_20090,N_22254);
and U24488 (N_24488,N_20244,N_21779);
nor U24489 (N_24489,N_21885,N_21010);
nand U24490 (N_24490,N_22164,N_22202);
nor U24491 (N_24491,N_21262,N_22115);
xnor U24492 (N_24492,N_21197,N_22102);
nor U24493 (N_24493,N_20554,N_21138);
nand U24494 (N_24494,N_21062,N_22378);
or U24495 (N_24495,N_21239,N_21225);
nand U24496 (N_24496,N_21465,N_20972);
or U24497 (N_24497,N_21365,N_21338);
nand U24498 (N_24498,N_21820,N_22305);
nor U24499 (N_24499,N_20271,N_20268);
and U24500 (N_24500,N_21055,N_20771);
and U24501 (N_24501,N_20765,N_20797);
nor U24502 (N_24502,N_21348,N_22260);
and U24503 (N_24503,N_21660,N_22490);
xnor U24504 (N_24504,N_22264,N_21517);
nand U24505 (N_24505,N_21979,N_20776);
or U24506 (N_24506,N_21338,N_21584);
nor U24507 (N_24507,N_21340,N_20862);
xnor U24508 (N_24508,N_20591,N_22109);
and U24509 (N_24509,N_20544,N_21088);
nor U24510 (N_24510,N_21059,N_21632);
xor U24511 (N_24511,N_21217,N_22273);
nor U24512 (N_24512,N_20746,N_22395);
or U24513 (N_24513,N_21341,N_21584);
nor U24514 (N_24514,N_20693,N_21766);
or U24515 (N_24515,N_21919,N_21348);
or U24516 (N_24516,N_20769,N_20066);
xnor U24517 (N_24517,N_20407,N_21848);
xor U24518 (N_24518,N_22093,N_21862);
or U24519 (N_24519,N_20295,N_20944);
or U24520 (N_24520,N_22436,N_20462);
xnor U24521 (N_24521,N_20354,N_21997);
nand U24522 (N_24522,N_20406,N_20493);
xnor U24523 (N_24523,N_20262,N_20167);
and U24524 (N_24524,N_21558,N_20369);
nor U24525 (N_24525,N_22254,N_21697);
nand U24526 (N_24526,N_21944,N_22046);
or U24527 (N_24527,N_21805,N_21469);
nor U24528 (N_24528,N_22124,N_20539);
or U24529 (N_24529,N_21463,N_21315);
nand U24530 (N_24530,N_20260,N_21263);
nand U24531 (N_24531,N_20605,N_22274);
or U24532 (N_24532,N_20387,N_20558);
and U24533 (N_24533,N_22482,N_21199);
nor U24534 (N_24534,N_20744,N_22330);
and U24535 (N_24535,N_21142,N_22326);
xnor U24536 (N_24536,N_21587,N_21150);
and U24537 (N_24537,N_20587,N_21024);
and U24538 (N_24538,N_20055,N_20446);
or U24539 (N_24539,N_22237,N_20099);
nor U24540 (N_24540,N_22308,N_22428);
nor U24541 (N_24541,N_22472,N_20168);
and U24542 (N_24542,N_20454,N_21186);
or U24543 (N_24543,N_21903,N_20185);
nand U24544 (N_24544,N_21028,N_20734);
and U24545 (N_24545,N_21443,N_21222);
nand U24546 (N_24546,N_21193,N_21251);
nand U24547 (N_24547,N_21906,N_20050);
xor U24548 (N_24548,N_21952,N_20946);
and U24549 (N_24549,N_21776,N_20312);
or U24550 (N_24550,N_20334,N_20088);
nor U24551 (N_24551,N_20707,N_21715);
nand U24552 (N_24552,N_21148,N_21506);
and U24553 (N_24553,N_20699,N_21445);
xor U24554 (N_24554,N_20653,N_20637);
nor U24555 (N_24555,N_20214,N_21651);
nand U24556 (N_24556,N_22015,N_20699);
and U24557 (N_24557,N_20652,N_20582);
nand U24558 (N_24558,N_21510,N_20102);
and U24559 (N_24559,N_20405,N_21147);
xor U24560 (N_24560,N_21691,N_22466);
nand U24561 (N_24561,N_21645,N_22165);
or U24562 (N_24562,N_20243,N_20597);
nand U24563 (N_24563,N_22027,N_22168);
xor U24564 (N_24564,N_21927,N_20631);
xnor U24565 (N_24565,N_21001,N_22080);
xor U24566 (N_24566,N_21652,N_20973);
nand U24567 (N_24567,N_21252,N_21083);
nand U24568 (N_24568,N_22277,N_20068);
nand U24569 (N_24569,N_22359,N_21513);
nand U24570 (N_24570,N_20566,N_20795);
and U24571 (N_24571,N_20829,N_20979);
xnor U24572 (N_24572,N_21270,N_21000);
and U24573 (N_24573,N_22003,N_20263);
nor U24574 (N_24574,N_20385,N_20725);
and U24575 (N_24575,N_20407,N_22139);
or U24576 (N_24576,N_20358,N_21358);
and U24577 (N_24577,N_21416,N_20687);
or U24578 (N_24578,N_20179,N_22451);
or U24579 (N_24579,N_22334,N_20722);
or U24580 (N_24580,N_21322,N_21163);
nand U24581 (N_24581,N_20798,N_20706);
or U24582 (N_24582,N_21352,N_20024);
nand U24583 (N_24583,N_20165,N_20089);
and U24584 (N_24584,N_20228,N_22187);
nand U24585 (N_24585,N_20071,N_21596);
or U24586 (N_24586,N_22382,N_20992);
nor U24587 (N_24587,N_20218,N_21646);
xor U24588 (N_24588,N_20590,N_21459);
nand U24589 (N_24589,N_20305,N_21162);
nand U24590 (N_24590,N_20133,N_21319);
and U24591 (N_24591,N_21822,N_20200);
nand U24592 (N_24592,N_20201,N_20448);
or U24593 (N_24593,N_21343,N_21210);
xor U24594 (N_24594,N_20025,N_22226);
or U24595 (N_24595,N_21017,N_20664);
nand U24596 (N_24596,N_21704,N_20390);
nor U24597 (N_24597,N_22022,N_20248);
nand U24598 (N_24598,N_20978,N_20272);
or U24599 (N_24599,N_20241,N_20699);
xnor U24600 (N_24600,N_21756,N_21226);
nand U24601 (N_24601,N_21351,N_22025);
nand U24602 (N_24602,N_20069,N_20708);
nand U24603 (N_24603,N_21983,N_22434);
xnor U24604 (N_24604,N_20526,N_21275);
nor U24605 (N_24605,N_21834,N_21743);
xnor U24606 (N_24606,N_21020,N_20695);
and U24607 (N_24607,N_21369,N_20610);
xnor U24608 (N_24608,N_20493,N_20028);
nor U24609 (N_24609,N_20140,N_21722);
and U24610 (N_24610,N_21853,N_22485);
and U24611 (N_24611,N_21281,N_21565);
or U24612 (N_24612,N_21266,N_21492);
xor U24613 (N_24613,N_20439,N_21378);
or U24614 (N_24614,N_22365,N_21297);
or U24615 (N_24615,N_22319,N_20390);
or U24616 (N_24616,N_21405,N_21942);
xor U24617 (N_24617,N_20747,N_21589);
or U24618 (N_24618,N_22172,N_20932);
nand U24619 (N_24619,N_20908,N_20548);
xor U24620 (N_24620,N_22077,N_21174);
nor U24621 (N_24621,N_22087,N_22031);
or U24622 (N_24622,N_22366,N_22250);
and U24623 (N_24623,N_21641,N_20050);
and U24624 (N_24624,N_20480,N_20884);
xor U24625 (N_24625,N_22436,N_21008);
and U24626 (N_24626,N_20660,N_20747);
xnor U24627 (N_24627,N_20023,N_20577);
xnor U24628 (N_24628,N_21095,N_20916);
xor U24629 (N_24629,N_20833,N_20496);
nand U24630 (N_24630,N_20381,N_21334);
and U24631 (N_24631,N_21705,N_21293);
xnor U24632 (N_24632,N_20986,N_22030);
xor U24633 (N_24633,N_20794,N_20274);
and U24634 (N_24634,N_20663,N_22321);
xnor U24635 (N_24635,N_21847,N_21386);
or U24636 (N_24636,N_22415,N_20062);
nor U24637 (N_24637,N_22257,N_21039);
or U24638 (N_24638,N_20963,N_21990);
and U24639 (N_24639,N_21246,N_21455);
nand U24640 (N_24640,N_22204,N_21758);
nor U24641 (N_24641,N_20905,N_20900);
nor U24642 (N_24642,N_21692,N_21167);
nand U24643 (N_24643,N_21545,N_21757);
nor U24644 (N_24644,N_20976,N_20166);
and U24645 (N_24645,N_20052,N_21019);
nor U24646 (N_24646,N_22065,N_21752);
nand U24647 (N_24647,N_22387,N_20856);
or U24648 (N_24648,N_20875,N_22170);
nand U24649 (N_24649,N_21962,N_22350);
nor U24650 (N_24650,N_21058,N_21140);
nor U24651 (N_24651,N_20280,N_20163);
or U24652 (N_24652,N_20426,N_20868);
nand U24653 (N_24653,N_22266,N_22102);
nand U24654 (N_24654,N_21023,N_20909);
nor U24655 (N_24655,N_21304,N_20439);
xor U24656 (N_24656,N_20984,N_20095);
and U24657 (N_24657,N_21136,N_20213);
nand U24658 (N_24658,N_21327,N_21167);
nand U24659 (N_24659,N_20721,N_20880);
and U24660 (N_24660,N_22363,N_20268);
nand U24661 (N_24661,N_21920,N_21678);
nor U24662 (N_24662,N_21512,N_20403);
nand U24663 (N_24663,N_21639,N_20588);
nand U24664 (N_24664,N_21076,N_20746);
nor U24665 (N_24665,N_21390,N_20170);
or U24666 (N_24666,N_20687,N_21381);
and U24667 (N_24667,N_21204,N_21533);
nand U24668 (N_24668,N_20665,N_20519);
xnor U24669 (N_24669,N_21875,N_20054);
and U24670 (N_24670,N_20406,N_20625);
nand U24671 (N_24671,N_21170,N_20865);
xor U24672 (N_24672,N_20497,N_20444);
or U24673 (N_24673,N_21957,N_20975);
and U24674 (N_24674,N_20763,N_22375);
xnor U24675 (N_24675,N_21808,N_21648);
and U24676 (N_24676,N_21366,N_20092);
nor U24677 (N_24677,N_21955,N_20302);
or U24678 (N_24678,N_22482,N_20652);
or U24679 (N_24679,N_21938,N_20178);
nand U24680 (N_24680,N_21359,N_20958);
or U24681 (N_24681,N_22005,N_20515);
nor U24682 (N_24682,N_22091,N_20944);
nand U24683 (N_24683,N_20551,N_22364);
nor U24684 (N_24684,N_21538,N_21374);
and U24685 (N_24685,N_20746,N_22221);
nor U24686 (N_24686,N_21610,N_22061);
nand U24687 (N_24687,N_21355,N_21356);
or U24688 (N_24688,N_20517,N_22264);
xor U24689 (N_24689,N_20347,N_22403);
nor U24690 (N_24690,N_20375,N_21937);
nand U24691 (N_24691,N_21240,N_21376);
or U24692 (N_24692,N_20309,N_21910);
or U24693 (N_24693,N_21135,N_21381);
xor U24694 (N_24694,N_21082,N_21967);
nor U24695 (N_24695,N_20216,N_21437);
nand U24696 (N_24696,N_21872,N_22256);
nand U24697 (N_24697,N_20375,N_20255);
and U24698 (N_24698,N_21902,N_20242);
or U24699 (N_24699,N_21161,N_21358);
and U24700 (N_24700,N_21602,N_20105);
xnor U24701 (N_24701,N_21448,N_21338);
nand U24702 (N_24702,N_21605,N_20702);
and U24703 (N_24703,N_21972,N_20378);
and U24704 (N_24704,N_21272,N_21785);
or U24705 (N_24705,N_20802,N_21064);
and U24706 (N_24706,N_20974,N_21270);
xor U24707 (N_24707,N_22367,N_22371);
xnor U24708 (N_24708,N_21945,N_22050);
nand U24709 (N_24709,N_20457,N_22157);
nor U24710 (N_24710,N_20205,N_22154);
nor U24711 (N_24711,N_20059,N_21074);
or U24712 (N_24712,N_20543,N_20251);
and U24713 (N_24713,N_20731,N_22145);
nor U24714 (N_24714,N_22030,N_21892);
nand U24715 (N_24715,N_22276,N_21566);
xnor U24716 (N_24716,N_20242,N_21148);
xnor U24717 (N_24717,N_20914,N_20819);
nor U24718 (N_24718,N_21244,N_21924);
or U24719 (N_24719,N_21814,N_20028);
nor U24720 (N_24720,N_20579,N_21868);
nand U24721 (N_24721,N_22205,N_21592);
and U24722 (N_24722,N_21937,N_21212);
xor U24723 (N_24723,N_20951,N_21267);
nor U24724 (N_24724,N_22233,N_20431);
and U24725 (N_24725,N_20847,N_20720);
xnor U24726 (N_24726,N_22172,N_22450);
xnor U24727 (N_24727,N_21840,N_20142);
and U24728 (N_24728,N_22367,N_21371);
xnor U24729 (N_24729,N_21007,N_21985);
xor U24730 (N_24730,N_22203,N_22023);
nand U24731 (N_24731,N_21234,N_21499);
or U24732 (N_24732,N_20653,N_20386);
or U24733 (N_24733,N_20358,N_20498);
xnor U24734 (N_24734,N_21172,N_20171);
and U24735 (N_24735,N_22099,N_22279);
xor U24736 (N_24736,N_20644,N_20155);
nand U24737 (N_24737,N_20349,N_21354);
and U24738 (N_24738,N_22471,N_22359);
nor U24739 (N_24739,N_22273,N_20252);
nor U24740 (N_24740,N_20684,N_21802);
nand U24741 (N_24741,N_20961,N_21718);
and U24742 (N_24742,N_22345,N_20971);
nor U24743 (N_24743,N_21784,N_20476);
and U24744 (N_24744,N_21269,N_20884);
nor U24745 (N_24745,N_22435,N_20190);
nor U24746 (N_24746,N_22233,N_20473);
or U24747 (N_24747,N_20974,N_20080);
xnor U24748 (N_24748,N_21582,N_20732);
xnor U24749 (N_24749,N_21950,N_20976);
xor U24750 (N_24750,N_21541,N_22423);
or U24751 (N_24751,N_20405,N_20942);
xor U24752 (N_24752,N_21370,N_22208);
nor U24753 (N_24753,N_21501,N_21877);
and U24754 (N_24754,N_20006,N_20636);
nand U24755 (N_24755,N_21953,N_21693);
and U24756 (N_24756,N_21834,N_20505);
nand U24757 (N_24757,N_22274,N_21909);
nand U24758 (N_24758,N_22317,N_20899);
xor U24759 (N_24759,N_21349,N_21855);
or U24760 (N_24760,N_21582,N_22215);
nand U24761 (N_24761,N_20485,N_20566);
and U24762 (N_24762,N_20308,N_22462);
or U24763 (N_24763,N_20815,N_20555);
and U24764 (N_24764,N_20298,N_21752);
nor U24765 (N_24765,N_20942,N_22342);
nand U24766 (N_24766,N_21409,N_20121);
nand U24767 (N_24767,N_20896,N_21888);
and U24768 (N_24768,N_20885,N_21972);
xor U24769 (N_24769,N_21159,N_21586);
and U24770 (N_24770,N_20225,N_22377);
nand U24771 (N_24771,N_22360,N_20557);
xor U24772 (N_24772,N_21929,N_21587);
xnor U24773 (N_24773,N_20910,N_22450);
and U24774 (N_24774,N_20156,N_22398);
and U24775 (N_24775,N_22454,N_22067);
and U24776 (N_24776,N_20927,N_21265);
xnor U24777 (N_24777,N_20038,N_21707);
or U24778 (N_24778,N_20439,N_20685);
xor U24779 (N_24779,N_20980,N_21520);
xnor U24780 (N_24780,N_20027,N_20585);
nor U24781 (N_24781,N_22258,N_20904);
nand U24782 (N_24782,N_20157,N_21020);
and U24783 (N_24783,N_21090,N_20260);
or U24784 (N_24784,N_21627,N_20113);
nand U24785 (N_24785,N_22436,N_20282);
nand U24786 (N_24786,N_20449,N_21239);
nand U24787 (N_24787,N_20243,N_20817);
nor U24788 (N_24788,N_21403,N_22468);
and U24789 (N_24789,N_20973,N_22144);
or U24790 (N_24790,N_20574,N_20125);
and U24791 (N_24791,N_20989,N_22037);
or U24792 (N_24792,N_21083,N_21549);
xnor U24793 (N_24793,N_20080,N_21278);
and U24794 (N_24794,N_21395,N_20646);
nand U24795 (N_24795,N_21837,N_21460);
nand U24796 (N_24796,N_20411,N_20714);
nand U24797 (N_24797,N_22072,N_21230);
xor U24798 (N_24798,N_21589,N_21453);
xnor U24799 (N_24799,N_20344,N_20780);
xor U24800 (N_24800,N_22432,N_20602);
nand U24801 (N_24801,N_20019,N_20673);
and U24802 (N_24802,N_20563,N_20994);
nand U24803 (N_24803,N_21649,N_21710);
nand U24804 (N_24804,N_22028,N_20508);
nand U24805 (N_24805,N_20304,N_20070);
or U24806 (N_24806,N_20704,N_22383);
nand U24807 (N_24807,N_22446,N_20353);
xor U24808 (N_24808,N_20143,N_21799);
or U24809 (N_24809,N_21399,N_21815);
xnor U24810 (N_24810,N_20420,N_20201);
or U24811 (N_24811,N_20107,N_20194);
nor U24812 (N_24812,N_20618,N_21515);
nor U24813 (N_24813,N_20968,N_20628);
xor U24814 (N_24814,N_21980,N_22420);
nor U24815 (N_24815,N_22490,N_20391);
nor U24816 (N_24816,N_21662,N_20223);
and U24817 (N_24817,N_20929,N_20841);
nor U24818 (N_24818,N_20433,N_20859);
nand U24819 (N_24819,N_20509,N_20171);
xnor U24820 (N_24820,N_21718,N_21506);
and U24821 (N_24821,N_20792,N_20165);
nand U24822 (N_24822,N_21513,N_21651);
xnor U24823 (N_24823,N_20267,N_21455);
and U24824 (N_24824,N_22392,N_22247);
and U24825 (N_24825,N_21915,N_20450);
or U24826 (N_24826,N_22295,N_22494);
xor U24827 (N_24827,N_22212,N_21887);
xor U24828 (N_24828,N_20782,N_22427);
xor U24829 (N_24829,N_22386,N_20138);
nand U24830 (N_24830,N_22475,N_20407);
xnor U24831 (N_24831,N_21266,N_21454);
and U24832 (N_24832,N_21234,N_21344);
nand U24833 (N_24833,N_22375,N_20569);
or U24834 (N_24834,N_20055,N_21507);
and U24835 (N_24835,N_20584,N_22312);
or U24836 (N_24836,N_21276,N_21778);
nand U24837 (N_24837,N_20478,N_20527);
xor U24838 (N_24838,N_22170,N_20092);
and U24839 (N_24839,N_20202,N_20846);
nand U24840 (N_24840,N_21845,N_22160);
or U24841 (N_24841,N_20518,N_22026);
nand U24842 (N_24842,N_22459,N_20601);
xor U24843 (N_24843,N_21156,N_20180);
xor U24844 (N_24844,N_20647,N_20286);
or U24845 (N_24845,N_20742,N_20866);
nor U24846 (N_24846,N_21071,N_21874);
nor U24847 (N_24847,N_22101,N_21885);
xor U24848 (N_24848,N_22234,N_20032);
or U24849 (N_24849,N_20316,N_20074);
nor U24850 (N_24850,N_20947,N_22271);
nand U24851 (N_24851,N_20749,N_20230);
or U24852 (N_24852,N_21532,N_21097);
xnor U24853 (N_24853,N_20024,N_20817);
xnor U24854 (N_24854,N_20678,N_22186);
nand U24855 (N_24855,N_20816,N_21535);
nand U24856 (N_24856,N_20686,N_20946);
or U24857 (N_24857,N_22016,N_20473);
nand U24858 (N_24858,N_21276,N_21509);
xor U24859 (N_24859,N_20059,N_22248);
nor U24860 (N_24860,N_20149,N_21795);
and U24861 (N_24861,N_21356,N_20797);
and U24862 (N_24862,N_22026,N_20545);
and U24863 (N_24863,N_20811,N_21054);
xnor U24864 (N_24864,N_20849,N_22075);
and U24865 (N_24865,N_21386,N_20641);
nor U24866 (N_24866,N_20911,N_21552);
nand U24867 (N_24867,N_20256,N_20051);
nand U24868 (N_24868,N_22262,N_21642);
nand U24869 (N_24869,N_20208,N_20761);
and U24870 (N_24870,N_22470,N_22499);
and U24871 (N_24871,N_22458,N_22074);
nor U24872 (N_24872,N_20497,N_21593);
nand U24873 (N_24873,N_20958,N_22334);
xor U24874 (N_24874,N_20338,N_21174);
xor U24875 (N_24875,N_20299,N_20380);
and U24876 (N_24876,N_21588,N_20798);
and U24877 (N_24877,N_22019,N_21082);
or U24878 (N_24878,N_21588,N_20438);
nor U24879 (N_24879,N_20281,N_22270);
and U24880 (N_24880,N_21091,N_22047);
and U24881 (N_24881,N_21764,N_20909);
xnor U24882 (N_24882,N_20614,N_21977);
nand U24883 (N_24883,N_21767,N_20998);
nand U24884 (N_24884,N_22405,N_22359);
or U24885 (N_24885,N_21068,N_22430);
and U24886 (N_24886,N_21793,N_21377);
nor U24887 (N_24887,N_22132,N_21874);
nor U24888 (N_24888,N_20290,N_21116);
and U24889 (N_24889,N_22080,N_22125);
or U24890 (N_24890,N_20473,N_21292);
nand U24891 (N_24891,N_21326,N_20630);
and U24892 (N_24892,N_20730,N_21020);
nand U24893 (N_24893,N_21364,N_20958);
or U24894 (N_24894,N_22019,N_20924);
xnor U24895 (N_24895,N_21700,N_22418);
or U24896 (N_24896,N_20416,N_22374);
or U24897 (N_24897,N_21792,N_21584);
or U24898 (N_24898,N_21461,N_20589);
nand U24899 (N_24899,N_20882,N_22163);
and U24900 (N_24900,N_20877,N_22258);
nand U24901 (N_24901,N_22398,N_21726);
xor U24902 (N_24902,N_20550,N_20878);
and U24903 (N_24903,N_20024,N_20517);
and U24904 (N_24904,N_21715,N_20744);
nand U24905 (N_24905,N_22125,N_20963);
xor U24906 (N_24906,N_21406,N_20618);
xnor U24907 (N_24907,N_22113,N_22245);
nand U24908 (N_24908,N_21372,N_20038);
nor U24909 (N_24909,N_22237,N_20069);
and U24910 (N_24910,N_21256,N_21936);
or U24911 (N_24911,N_21816,N_22496);
and U24912 (N_24912,N_20870,N_20313);
nor U24913 (N_24913,N_20608,N_21999);
nor U24914 (N_24914,N_22432,N_21491);
nor U24915 (N_24915,N_20543,N_22061);
and U24916 (N_24916,N_20879,N_21998);
nor U24917 (N_24917,N_21054,N_21035);
or U24918 (N_24918,N_21933,N_20734);
nand U24919 (N_24919,N_21995,N_20296);
and U24920 (N_24920,N_20319,N_21038);
xnor U24921 (N_24921,N_20271,N_22228);
nor U24922 (N_24922,N_21528,N_21772);
nand U24923 (N_24923,N_21491,N_20242);
and U24924 (N_24924,N_22329,N_20182);
nor U24925 (N_24925,N_20003,N_20120);
and U24926 (N_24926,N_21634,N_20759);
nor U24927 (N_24927,N_20669,N_20089);
xor U24928 (N_24928,N_20518,N_22444);
xor U24929 (N_24929,N_20024,N_20065);
and U24930 (N_24930,N_22306,N_22015);
and U24931 (N_24931,N_22385,N_20975);
or U24932 (N_24932,N_21707,N_21088);
or U24933 (N_24933,N_22095,N_22145);
nor U24934 (N_24934,N_20912,N_21237);
xnor U24935 (N_24935,N_21122,N_21567);
nand U24936 (N_24936,N_20668,N_21912);
nor U24937 (N_24937,N_22141,N_21387);
or U24938 (N_24938,N_21398,N_22273);
xnor U24939 (N_24939,N_22261,N_20857);
xnor U24940 (N_24940,N_20125,N_20473);
nand U24941 (N_24941,N_20911,N_22094);
xnor U24942 (N_24942,N_20839,N_20094);
or U24943 (N_24943,N_21321,N_21228);
and U24944 (N_24944,N_21610,N_21926);
and U24945 (N_24945,N_22402,N_20121);
xor U24946 (N_24946,N_20970,N_21275);
and U24947 (N_24947,N_22342,N_20656);
nor U24948 (N_24948,N_20172,N_21925);
nor U24949 (N_24949,N_21541,N_21099);
or U24950 (N_24950,N_21598,N_21452);
or U24951 (N_24951,N_20674,N_22337);
or U24952 (N_24952,N_21624,N_20448);
nor U24953 (N_24953,N_21559,N_20586);
nand U24954 (N_24954,N_20943,N_20327);
or U24955 (N_24955,N_21390,N_21052);
and U24956 (N_24956,N_21983,N_20311);
nor U24957 (N_24957,N_20359,N_20668);
xnor U24958 (N_24958,N_21691,N_22458);
and U24959 (N_24959,N_22319,N_21747);
nand U24960 (N_24960,N_21594,N_20669);
xor U24961 (N_24961,N_20793,N_21358);
or U24962 (N_24962,N_21195,N_21690);
and U24963 (N_24963,N_21258,N_20683);
xor U24964 (N_24964,N_20902,N_22150);
xnor U24965 (N_24965,N_21796,N_22052);
nor U24966 (N_24966,N_20890,N_22244);
xnor U24967 (N_24967,N_21368,N_22460);
nor U24968 (N_24968,N_20477,N_20359);
or U24969 (N_24969,N_22006,N_21239);
nand U24970 (N_24970,N_21509,N_20994);
and U24971 (N_24971,N_21735,N_22250);
and U24972 (N_24972,N_20317,N_21107);
nand U24973 (N_24973,N_22280,N_20580);
xor U24974 (N_24974,N_22313,N_21558);
nand U24975 (N_24975,N_21536,N_20715);
nor U24976 (N_24976,N_22098,N_20547);
xor U24977 (N_24977,N_20970,N_22204);
nand U24978 (N_24978,N_21579,N_20872);
xor U24979 (N_24979,N_21882,N_21192);
nand U24980 (N_24980,N_21357,N_22195);
and U24981 (N_24981,N_20179,N_21546);
xor U24982 (N_24982,N_22428,N_20048);
nor U24983 (N_24983,N_22019,N_21310);
xnor U24984 (N_24984,N_21630,N_21746);
nand U24985 (N_24985,N_21177,N_20122);
nand U24986 (N_24986,N_21010,N_20111);
or U24987 (N_24987,N_20549,N_21551);
nor U24988 (N_24988,N_21204,N_21046);
xnor U24989 (N_24989,N_21983,N_21081);
or U24990 (N_24990,N_20700,N_22379);
and U24991 (N_24991,N_20033,N_20428);
or U24992 (N_24992,N_20445,N_22078);
or U24993 (N_24993,N_20365,N_20879);
or U24994 (N_24994,N_20875,N_20642);
xor U24995 (N_24995,N_22185,N_21739);
nand U24996 (N_24996,N_20167,N_20672);
nand U24997 (N_24997,N_20079,N_21653);
nand U24998 (N_24998,N_21329,N_22246);
nand U24999 (N_24999,N_21599,N_21615);
or UO_0 (O_0,N_24143,N_23303);
and UO_1 (O_1,N_23964,N_24519);
and UO_2 (O_2,N_23106,N_24673);
nand UO_3 (O_3,N_24189,N_22665);
or UO_4 (O_4,N_22681,N_23068);
nand UO_5 (O_5,N_24719,N_24176);
xnor UO_6 (O_6,N_23879,N_24395);
nor UO_7 (O_7,N_24550,N_23852);
and UO_8 (O_8,N_22946,N_23823);
and UO_9 (O_9,N_24931,N_22589);
nor UO_10 (O_10,N_22969,N_23772);
or UO_11 (O_11,N_22661,N_23388);
or UO_12 (O_12,N_24067,N_24145);
and UO_13 (O_13,N_24841,N_22749);
or UO_14 (O_14,N_22535,N_22725);
nor UO_15 (O_15,N_23005,N_23024);
xnor UO_16 (O_16,N_24574,N_23988);
and UO_17 (O_17,N_23966,N_23075);
nand UO_18 (O_18,N_23523,N_23034);
and UO_19 (O_19,N_24182,N_24029);
and UO_20 (O_20,N_24650,N_22837);
nor UO_21 (O_21,N_22640,N_24955);
nor UO_22 (O_22,N_22682,N_23037);
xor UO_23 (O_23,N_22819,N_22518);
and UO_24 (O_24,N_23796,N_24591);
xor UO_25 (O_25,N_24798,N_22773);
nand UO_26 (O_26,N_24575,N_22543);
nor UO_27 (O_27,N_22525,N_24496);
or UO_28 (O_28,N_23397,N_23612);
and UO_29 (O_29,N_22656,N_22724);
nor UO_30 (O_30,N_23732,N_24262);
nand UO_31 (O_31,N_24526,N_23582);
or UO_32 (O_32,N_24943,N_23228);
xor UO_33 (O_33,N_24066,N_22975);
nand UO_34 (O_34,N_24459,N_23477);
nand UO_35 (O_35,N_24102,N_24859);
and UO_36 (O_36,N_24226,N_24241);
nor UO_37 (O_37,N_24708,N_24071);
xnor UO_38 (O_38,N_24092,N_22613);
nor UO_39 (O_39,N_23422,N_24499);
nand UO_40 (O_40,N_23892,N_24439);
nand UO_41 (O_41,N_23583,N_23284);
xnor UO_42 (O_42,N_22949,N_24249);
or UO_43 (O_43,N_24737,N_24918);
and UO_44 (O_44,N_23437,N_22532);
or UO_45 (O_45,N_23475,N_23585);
xor UO_46 (O_46,N_24528,N_22838);
nand UO_47 (O_47,N_22978,N_23781);
and UO_48 (O_48,N_24529,N_23900);
or UO_49 (O_49,N_23280,N_24299);
nand UO_50 (O_50,N_23077,N_22654);
xor UO_51 (O_51,N_23872,N_23141);
or UO_52 (O_52,N_23450,N_24018);
nor UO_53 (O_53,N_23384,N_24015);
nor UO_54 (O_54,N_24876,N_24979);
and UO_55 (O_55,N_24214,N_23276);
or UO_56 (O_56,N_24588,N_24073);
or UO_57 (O_57,N_24573,N_23937);
xor UO_58 (O_58,N_22973,N_23036);
or UO_59 (O_59,N_24829,N_23263);
and UO_60 (O_60,N_24340,N_23807);
or UO_61 (O_61,N_24361,N_24794);
or UO_62 (O_62,N_22897,N_24111);
and UO_63 (O_63,N_22998,N_22933);
and UO_64 (O_64,N_24987,N_22855);
xnor UO_65 (O_65,N_24056,N_23294);
nand UO_66 (O_66,N_24784,N_24722);
nor UO_67 (O_67,N_23833,N_24374);
xnor UO_68 (O_68,N_24305,N_22805);
nand UO_69 (O_69,N_22792,N_22777);
and UO_70 (O_70,N_23500,N_23884);
or UO_71 (O_71,N_24233,N_22726);
nor UO_72 (O_72,N_24925,N_24264);
nand UO_73 (O_73,N_23288,N_24203);
nor UO_74 (O_74,N_23677,N_23190);
nand UO_75 (O_75,N_22573,N_24831);
nor UO_76 (O_76,N_22506,N_22999);
nand UO_77 (O_77,N_24744,N_24595);
nor UO_78 (O_78,N_23264,N_22655);
nand UO_79 (O_79,N_23650,N_24124);
or UO_80 (O_80,N_22699,N_24272);
or UO_81 (O_81,N_22785,N_23110);
nor UO_82 (O_82,N_23274,N_23579);
and UO_83 (O_83,N_23121,N_24070);
nor UO_84 (O_84,N_24576,N_24122);
xnor UO_85 (O_85,N_23390,N_24509);
nand UO_86 (O_86,N_24845,N_24676);
nor UO_87 (O_87,N_22616,N_23347);
nand UO_88 (O_88,N_24540,N_23491);
nor UO_89 (O_89,N_24287,N_23688);
nand UO_90 (O_90,N_23752,N_24052);
and UO_91 (O_91,N_24202,N_24043);
or UO_92 (O_92,N_23358,N_22541);
or UO_93 (O_93,N_24022,N_24332);
or UO_94 (O_94,N_24711,N_24545);
and UO_95 (O_95,N_23853,N_24805);
nand UO_96 (O_96,N_22937,N_24270);
xnor UO_97 (O_97,N_22686,N_24833);
and UO_98 (O_98,N_22923,N_23158);
or UO_99 (O_99,N_22818,N_23766);
nand UO_100 (O_100,N_23980,N_23600);
or UO_101 (O_101,N_24953,N_23260);
nand UO_102 (O_102,N_23604,N_24587);
nor UO_103 (O_103,N_23154,N_24606);
nor UO_104 (O_104,N_23527,N_24410);
xor UO_105 (O_105,N_22717,N_23040);
nand UO_106 (O_106,N_23241,N_22789);
nand UO_107 (O_107,N_22846,N_23267);
xnor UO_108 (O_108,N_22559,N_23044);
xor UO_109 (O_109,N_24154,N_23730);
nand UO_110 (O_110,N_24238,N_23888);
nand UO_111 (O_111,N_22971,N_24080);
xnor UO_112 (O_112,N_24635,N_24517);
nand UO_113 (O_113,N_23392,N_23117);
or UO_114 (O_114,N_24341,N_23953);
or UO_115 (O_115,N_24563,N_24271);
nor UO_116 (O_116,N_24342,N_23939);
nand UO_117 (O_117,N_24157,N_23842);
xnor UO_118 (O_118,N_23972,N_23671);
and UO_119 (O_119,N_23769,N_24791);
and UO_120 (O_120,N_24471,N_23530);
xor UO_121 (O_121,N_24914,N_23919);
or UO_122 (O_122,N_24725,N_24462);
or UO_123 (O_123,N_23237,N_22956);
nor UO_124 (O_124,N_22642,N_23365);
nand UO_125 (O_125,N_23969,N_22731);
or UO_126 (O_126,N_24454,N_22555);
or UO_127 (O_127,N_22505,N_24907);
xor UO_128 (O_128,N_23038,N_22683);
xor UO_129 (O_129,N_23349,N_23925);
nand UO_130 (O_130,N_24922,N_23759);
nand UO_131 (O_131,N_24594,N_24856);
and UO_132 (O_132,N_23004,N_23101);
nor UO_133 (O_133,N_23584,N_23314);
and UO_134 (O_134,N_24551,N_22893);
or UO_135 (O_135,N_23447,N_23663);
and UO_136 (O_136,N_23587,N_23809);
nor UO_137 (O_137,N_22840,N_23719);
nand UO_138 (O_138,N_24893,N_22844);
nor UO_139 (O_139,N_24755,N_22934);
xor UO_140 (O_140,N_23277,N_23748);
or UO_141 (O_141,N_23750,N_23291);
xor UO_142 (O_142,N_24243,N_23637);
nand UO_143 (O_143,N_23640,N_24050);
and UO_144 (O_144,N_24826,N_24417);
xnor UO_145 (O_145,N_24348,N_23982);
nor UO_146 (O_146,N_24218,N_23103);
xor UO_147 (O_147,N_23393,N_24012);
nand UO_148 (O_148,N_23409,N_23448);
xnor UO_149 (O_149,N_24713,N_24780);
xor UO_150 (O_150,N_24198,N_24220);
xnor UO_151 (O_151,N_22542,N_24866);
and UO_152 (O_152,N_24633,N_22500);
and UO_153 (O_153,N_22631,N_22585);
or UO_154 (O_154,N_24490,N_23548);
xor UO_155 (O_155,N_23742,N_22925);
nor UO_156 (O_156,N_22502,N_23028);
nor UO_157 (O_157,N_23296,N_22877);
nand UO_158 (O_158,N_24438,N_22641);
nand UO_159 (O_159,N_24685,N_23931);
and UO_160 (O_160,N_23346,N_24852);
nor UO_161 (O_161,N_24399,N_24631);
nand UO_162 (O_162,N_24892,N_23091);
and UO_163 (O_163,N_24019,N_23062);
xnor UO_164 (O_164,N_22887,N_24774);
xor UO_165 (O_165,N_24853,N_23078);
xor UO_166 (O_166,N_23856,N_24387);
xnor UO_167 (O_167,N_24771,N_23696);
xnor UO_168 (O_168,N_24473,N_22827);
or UO_169 (O_169,N_22888,N_22797);
xnor UO_170 (O_170,N_22571,N_22754);
nor UO_171 (O_171,N_24620,N_23309);
and UO_172 (O_172,N_22760,N_23261);
nand UO_173 (O_173,N_22938,N_22637);
nand UO_174 (O_174,N_22741,N_23381);
and UO_175 (O_175,N_24166,N_23130);
and UO_176 (O_176,N_22578,N_24937);
nand UO_177 (O_177,N_23985,N_24195);
nand UO_178 (O_178,N_24846,N_24107);
nor UO_179 (O_179,N_24824,N_24707);
or UO_180 (O_180,N_23461,N_24174);
nand UO_181 (O_181,N_23735,N_24658);
xor UO_182 (O_182,N_24184,N_23271);
or UO_183 (O_183,N_24649,N_23569);
and UO_184 (O_184,N_22733,N_24729);
or UO_185 (O_185,N_24084,N_23188);
nand UO_186 (O_186,N_24413,N_24141);
or UO_187 (O_187,N_23245,N_24643);
nand UO_188 (O_188,N_23147,N_24186);
and UO_189 (O_189,N_24915,N_23764);
nand UO_190 (O_190,N_24873,N_24038);
xor UO_191 (O_191,N_24760,N_23387);
nor UO_192 (O_192,N_24242,N_23191);
nand UO_193 (O_193,N_24133,N_24730);
or UO_194 (O_194,N_23981,N_23518);
nor UO_195 (O_195,N_22746,N_22562);
xnor UO_196 (O_196,N_24695,N_23832);
or UO_197 (O_197,N_24571,N_24169);
or UO_198 (O_198,N_24059,N_22990);
nor UO_199 (O_199,N_23557,N_24261);
xor UO_200 (O_200,N_22873,N_23380);
xor UO_201 (O_201,N_24608,N_23176);
and UO_202 (O_202,N_23208,N_22790);
nand UO_203 (O_203,N_23070,N_24208);
nand UO_204 (O_204,N_22638,N_22703);
or UO_205 (O_205,N_22581,N_23090);
xor UO_206 (O_206,N_23834,N_23921);
and UO_207 (O_207,N_24512,N_23869);
nand UO_208 (O_208,N_22700,N_23107);
or UO_209 (O_209,N_24349,N_23410);
nor UO_210 (O_210,N_24162,N_22904);
nor UO_211 (O_211,N_22663,N_24449);
and UO_212 (O_212,N_24160,N_24093);
nor UO_213 (O_213,N_22895,N_22940);
nor UO_214 (O_214,N_23354,N_22714);
or UO_215 (O_215,N_23161,N_23416);
or UO_216 (O_216,N_22776,N_22859);
or UO_217 (O_217,N_23670,N_24781);
xnor UO_218 (O_218,N_23702,N_23368);
nand UO_219 (O_219,N_24662,N_22566);
nand UO_220 (O_220,N_24148,N_22950);
nand UO_221 (O_221,N_24675,N_24338);
xor UO_222 (O_222,N_23767,N_24848);
and UO_223 (O_223,N_22503,N_23425);
and UO_224 (O_224,N_23882,N_23076);
nor UO_225 (O_225,N_24373,N_23496);
or UO_226 (O_226,N_22926,N_24355);
xnor UO_227 (O_227,N_23114,N_24127);
nand UO_228 (O_228,N_24855,N_24165);
xor UO_229 (O_229,N_23444,N_22786);
and UO_230 (O_230,N_23345,N_23229);
or UO_231 (O_231,N_24328,N_23200);
nand UO_232 (O_232,N_23064,N_24803);
xnor UO_233 (O_233,N_24615,N_22899);
xnor UO_234 (O_234,N_23166,N_24319);
nor UO_235 (O_235,N_24753,N_22890);
and UO_236 (O_236,N_24516,N_24508);
or UO_237 (O_237,N_22929,N_23621);
xnor UO_238 (O_238,N_24583,N_23306);
or UO_239 (O_239,N_22698,N_24054);
xnor UO_240 (O_240,N_24391,N_24201);
nand UO_241 (O_241,N_24240,N_23338);
xor UO_242 (O_242,N_23348,N_24069);
or UO_243 (O_243,N_23510,N_22708);
nand UO_244 (O_244,N_24554,N_24627);
nor UO_245 (O_245,N_24721,N_24644);
nand UO_246 (O_246,N_22924,N_23227);
nand UO_247 (O_247,N_22602,N_22551);
nor UO_248 (O_248,N_22539,N_23638);
nor UO_249 (O_249,N_22830,N_24874);
or UO_250 (O_250,N_22951,N_23083);
xor UO_251 (O_251,N_23223,N_23300);
xor UO_252 (O_252,N_24311,N_23812);
xor UO_253 (O_253,N_24756,N_24634);
or UO_254 (O_254,N_23802,N_23613);
nand UO_255 (O_255,N_24382,N_24538);
and UO_256 (O_256,N_24652,N_23403);
nor UO_257 (O_257,N_24983,N_22565);
nor UO_258 (O_258,N_22643,N_23019);
nand UO_259 (O_259,N_23813,N_24369);
nor UO_260 (O_260,N_24933,N_24468);
xor UO_261 (O_261,N_23443,N_24096);
or UO_262 (O_262,N_24881,N_22531);
and UO_263 (O_263,N_23849,N_24535);
xnor UO_264 (O_264,N_23170,N_23421);
xor UO_265 (O_265,N_22530,N_23597);
or UO_266 (O_266,N_23698,N_23377);
or UO_267 (O_267,N_23924,N_23171);
or UO_268 (O_268,N_23249,N_24995);
xnor UO_269 (O_269,N_24191,N_24228);
nand UO_270 (O_270,N_24916,N_23343);
and UO_271 (O_271,N_24014,N_23041);
or UO_272 (O_272,N_23353,N_23687);
or UO_273 (O_273,N_23538,N_23187);
xor UO_274 (O_274,N_22875,N_24539);
and UO_275 (O_275,N_24706,N_23434);
and UO_276 (O_276,N_24068,N_23887);
nor UO_277 (O_277,N_23289,N_24592);
nor UO_278 (O_278,N_24209,N_24739);
nor UO_279 (O_279,N_23479,N_24281);
nor UO_280 (O_280,N_23873,N_23533);
and UO_281 (O_281,N_22764,N_23133);
xnor UO_282 (O_282,N_24702,N_24932);
nand UO_283 (O_283,N_23578,N_24295);
nand UO_284 (O_284,N_24078,N_23991);
and UO_285 (O_285,N_23466,N_23279);
xor UO_286 (O_286,N_23727,N_23693);
xnor UO_287 (O_287,N_24236,N_24447);
or UO_288 (O_288,N_24075,N_24385);
nand UO_289 (O_289,N_23554,N_22534);
nand UO_290 (O_290,N_23027,N_23428);
nor UO_291 (O_291,N_24904,N_22845);
nor UO_292 (O_292,N_23224,N_23895);
nand UO_293 (O_293,N_23559,N_24333);
nor UO_294 (O_294,N_24021,N_23630);
or UO_295 (O_295,N_23737,N_23148);
nand UO_296 (O_296,N_23283,N_22809);
and UO_297 (O_297,N_22958,N_24365);
xnor UO_298 (O_298,N_24742,N_22516);
and UO_299 (O_299,N_23993,N_24344);
and UO_300 (O_300,N_23020,N_24911);
nand UO_301 (O_301,N_24619,N_24809);
xor UO_302 (O_302,N_23625,N_22861);
or UO_303 (O_303,N_24398,N_22979);
nor UO_304 (O_304,N_24183,N_23015);
and UO_305 (O_305,N_22996,N_24677);
xnor UO_306 (O_306,N_23493,N_22507);
or UO_307 (O_307,N_24764,N_24950);
nand UO_308 (O_308,N_23927,N_24890);
nand UO_309 (O_309,N_22902,N_23747);
and UO_310 (O_310,N_23516,N_22753);
nor UO_311 (O_311,N_24642,N_23675);
xor UO_312 (O_312,N_22848,N_23344);
nand UO_313 (O_313,N_23456,N_22833);
xnor UO_314 (O_314,N_23499,N_22652);
and UO_315 (O_315,N_24007,N_22671);
and UO_316 (O_316,N_23374,N_24762);
xnor UO_317 (O_317,N_23486,N_22928);
xor UO_318 (O_318,N_23645,N_23143);
nor UO_319 (O_319,N_22992,N_22782);
nor UO_320 (O_320,N_23478,N_24980);
xnor UO_321 (O_321,N_24358,N_23618);
and UO_322 (O_322,N_23940,N_22916);
or UO_323 (O_323,N_24777,N_23626);
xor UO_324 (O_324,N_23646,N_24106);
nor UO_325 (O_325,N_22868,N_24322);
nor UO_326 (O_326,N_24320,N_24057);
or UO_327 (O_327,N_23945,N_24787);
nor UO_328 (O_328,N_23893,N_24278);
or UO_329 (O_329,N_23647,N_24337);
nand UO_330 (O_330,N_24546,N_24735);
nor UO_331 (O_331,N_22592,N_23438);
nor UO_332 (O_332,N_23045,N_22560);
xor UO_333 (O_333,N_22694,N_22743);
nand UO_334 (O_334,N_22501,N_24416);
nor UO_335 (O_335,N_23672,N_23053);
nor UO_336 (O_336,N_24232,N_23868);
and UO_337 (O_337,N_23960,N_24408);
or UO_338 (O_338,N_22907,N_23692);
nor UO_339 (O_339,N_24611,N_22801);
and UO_340 (O_340,N_24610,N_23104);
nand UO_341 (O_341,N_23631,N_22906);
nand UO_342 (O_342,N_23903,N_24171);
nor UO_343 (O_343,N_24577,N_23731);
or UO_344 (O_344,N_24108,N_24894);
and UO_345 (O_345,N_24375,N_23485);
and UO_346 (O_346,N_23494,N_23278);
nand UO_347 (O_347,N_24135,N_23861);
nor UO_348 (O_348,N_23476,N_22612);
or UO_349 (O_349,N_22954,N_24974);
nor UO_350 (O_350,N_23971,N_23897);
and UO_351 (O_351,N_23460,N_23048);
xnor UO_352 (O_352,N_23060,N_22599);
nand UO_353 (O_353,N_24090,N_24193);
nand UO_354 (O_354,N_22752,N_24260);
nor UO_355 (O_355,N_22715,N_23285);
nand UO_356 (O_356,N_23679,N_23446);
xor UO_357 (O_357,N_23620,N_24625);
xor UO_358 (O_358,N_24982,N_23016);
xnor UO_359 (O_359,N_23705,N_22751);
xor UO_360 (O_360,N_24210,N_23576);
nor UO_361 (O_361,N_24808,N_23412);
nor UO_362 (O_362,N_24568,N_23168);
xor UO_363 (O_363,N_24119,N_23525);
and UO_364 (O_364,N_24750,N_24248);
nor UO_365 (O_365,N_24971,N_23907);
and UO_366 (O_366,N_22762,N_22705);
xor UO_367 (O_367,N_24871,N_23838);
or UO_368 (O_368,N_23093,N_22811);
and UO_369 (O_369,N_22993,N_24103);
or UO_370 (O_370,N_22968,N_24996);
nand UO_371 (O_371,N_22882,N_23911);
or UO_372 (O_372,N_23127,N_22966);
xnor UO_373 (O_373,N_23482,N_24800);
xor UO_374 (O_374,N_23001,N_23366);
xnor UO_375 (O_375,N_24268,N_23965);
xnor UO_376 (O_376,N_24682,N_23811);
nand UO_377 (O_377,N_23762,N_24788);
nor UO_378 (O_378,N_23032,N_23754);
or UO_379 (O_379,N_24415,N_24088);
xnor UO_380 (O_380,N_23949,N_23956);
and UO_381 (O_381,N_24547,N_24020);
nor UO_382 (O_382,N_24616,N_23257);
or UO_383 (O_383,N_22997,N_22898);
nor UO_384 (O_384,N_22630,N_23259);
nor UO_385 (O_385,N_24993,N_24830);
or UO_386 (O_386,N_24356,N_23420);
or UO_387 (O_387,N_23023,N_23791);
xor UO_388 (O_388,N_23411,N_23634);
and UO_389 (O_389,N_22563,N_22546);
nand UO_390 (O_390,N_24301,N_23866);
nand UO_391 (O_391,N_23788,N_24807);
nand UO_392 (O_392,N_23871,N_23863);
or UO_393 (O_393,N_22552,N_23877);
and UO_394 (O_394,N_24469,N_22672);
xor UO_395 (O_395,N_22965,N_23627);
or UO_396 (O_396,N_23094,N_22635);
nor UO_397 (O_397,N_23607,N_24079);
nor UO_398 (O_398,N_24053,N_24992);
nand UO_399 (O_399,N_22981,N_24006);
nand UO_400 (O_400,N_23550,N_23322);
nor UO_401 (O_401,N_24474,N_24674);
nor UO_402 (O_402,N_23361,N_23653);
xor UO_403 (O_403,N_22988,N_22945);
nor UO_404 (O_404,N_23622,N_23826);
nand UO_405 (O_405,N_24476,N_24857);
nand UO_406 (O_406,N_23617,N_22570);
nand UO_407 (O_407,N_23898,N_24827);
xor UO_408 (O_408,N_24282,N_24666);
nor UO_409 (O_409,N_22884,N_24041);
xnor UO_410 (O_410,N_24500,N_23112);
nand UO_411 (O_411,N_24956,N_24255);
nand UO_412 (O_412,N_22930,N_23978);
xnor UO_413 (O_413,N_23857,N_22567);
nor UO_414 (O_414,N_24003,N_24976);
and UO_415 (O_415,N_24370,N_24645);
xor UO_416 (O_416,N_23102,N_24968);
nor UO_417 (O_417,N_24741,N_24734);
xor UO_418 (O_418,N_22696,N_24430);
or UO_419 (O_419,N_24265,N_24294);
and UO_420 (O_420,N_24244,N_22540);
or UO_421 (O_421,N_22727,N_22866);
nand UO_422 (O_422,N_23035,N_23398);
or UO_423 (O_423,N_24909,N_22621);
nor UO_424 (O_424,N_24085,N_22995);
and UO_425 (O_425,N_22678,N_24900);
nor UO_426 (O_426,N_24903,N_23383);
or UO_427 (O_427,N_23707,N_24076);
or UO_428 (O_428,N_23321,N_23920);
nand UO_429 (O_429,N_24795,N_23574);
xor UO_430 (O_430,N_22863,N_22759);
and UO_431 (O_431,N_22739,N_23994);
nor UO_432 (O_432,N_24661,N_22852);
nor UO_433 (O_433,N_22679,N_24432);
xnor UO_434 (O_434,N_24558,N_23058);
or UO_435 (O_435,N_22829,N_24495);
xnor UO_436 (O_436,N_24728,N_23069);
or UO_437 (O_437,N_23814,N_23656);
or UO_438 (O_438,N_22835,N_24033);
or UO_439 (O_439,N_23445,N_23801);
nand UO_440 (O_440,N_22834,N_23149);
or UO_441 (O_441,N_24697,N_24194);
xnor UO_442 (O_442,N_22927,N_23218);
or UO_443 (O_443,N_22912,N_23736);
or UO_444 (O_444,N_23673,N_22823);
and UO_445 (O_445,N_23441,N_24283);
and UO_446 (O_446,N_22794,N_24276);
xnor UO_447 (O_447,N_23449,N_24738);
nand UO_448 (O_448,N_24680,N_23596);
nand UO_449 (O_449,N_23235,N_22883);
or UO_450 (O_450,N_22594,N_24110);
xnor UO_451 (O_451,N_22947,N_24843);
nand UO_452 (O_452,N_22849,N_22847);
or UO_453 (O_453,N_23676,N_22879);
or UO_454 (O_454,N_24197,N_24440);
xnor UO_455 (O_455,N_24797,N_23598);
xnor UO_456 (O_456,N_22985,N_22688);
nand UO_457 (O_457,N_24040,N_24289);
and UO_458 (O_458,N_23498,N_22524);
xnor UO_459 (O_459,N_23363,N_22885);
xor UO_460 (O_460,N_24990,N_22817);
nand UO_461 (O_461,N_24152,N_22986);
xnor UO_462 (O_462,N_23402,N_24530);
nor UO_463 (O_463,N_23082,N_24754);
xor UO_464 (O_464,N_24331,N_23396);
xnor UO_465 (O_465,N_22821,N_22521);
nand UO_466 (O_466,N_24969,N_23529);
nand UO_467 (O_467,N_23139,N_24223);
nand UO_468 (O_468,N_23657,N_24670);
nand UO_469 (O_469,N_23184,N_23744);
and UO_470 (O_470,N_23194,N_24025);
or UO_471 (O_471,N_23591,N_22720);
nor UO_472 (O_472,N_23599,N_24882);
and UO_473 (O_473,N_23890,N_23706);
or UO_474 (O_474,N_24061,N_24823);
nand UO_475 (O_475,N_24884,N_23508);
xnor UO_476 (O_476,N_23544,N_24745);
nor UO_477 (O_477,N_23097,N_24889);
or UO_478 (O_478,N_23787,N_24930);
nand UO_479 (O_479,N_24441,N_23662);
or UO_480 (O_480,N_24589,N_23841);
nand UO_481 (O_481,N_22788,N_24134);
and UO_482 (O_482,N_23021,N_23963);
nor UO_483 (O_483,N_22948,N_23385);
nor UO_484 (O_484,N_23105,N_22583);
xnor UO_485 (O_485,N_24854,N_23153);
nand UO_486 (O_486,N_23932,N_23360);
nor UO_487 (O_487,N_22803,N_23836);
or UO_488 (O_488,N_24604,N_24603);
nand UO_489 (O_489,N_23014,N_23367);
nand UO_490 (O_490,N_22557,N_24752);
nand UO_491 (O_491,N_24696,N_22769);
xor UO_492 (O_492,N_24304,N_23968);
and UO_493 (O_493,N_24074,N_22972);
nor UO_494 (O_494,N_23172,N_22693);
xnor UO_495 (O_495,N_24277,N_23116);
nor UO_496 (O_496,N_22796,N_22771);
xnor UO_497 (O_497,N_24775,N_22677);
or UO_498 (O_498,N_23197,N_24504);
nand UO_499 (O_499,N_23896,N_24151);
and UO_500 (O_500,N_24518,N_23619);
xnor UO_501 (O_501,N_23717,N_24548);
xnor UO_502 (O_502,N_24351,N_23844);
xor UO_503 (O_503,N_23975,N_23225);
nor UO_504 (O_504,N_23547,N_24091);
xor UO_505 (O_505,N_23751,N_22577);
nor UO_506 (O_506,N_24751,N_24569);
or UO_507 (O_507,N_24027,N_23209);
nand UO_508 (O_508,N_24222,N_24487);
nand UO_509 (O_509,N_23710,N_23457);
and UO_510 (O_510,N_24310,N_24199);
nand UO_511 (O_511,N_23669,N_22590);
nor UO_512 (O_512,N_23183,N_23572);
xor UO_513 (O_513,N_22646,N_23770);
xor UO_514 (O_514,N_23250,N_23055);
nand UO_515 (O_515,N_24896,N_24446);
or UO_516 (O_516,N_23111,N_24380);
nand UO_517 (O_517,N_24164,N_24617);
and UO_518 (O_518,N_23240,N_23386);
nand UO_519 (O_519,N_24403,N_24307);
or UO_520 (O_520,N_24104,N_22862);
nor UO_521 (O_521,N_23575,N_24396);
xor UO_522 (O_522,N_22894,N_23961);
nor UO_523 (O_523,N_24180,N_24175);
xor UO_524 (O_524,N_22553,N_24460);
xnor UO_525 (O_525,N_23370,N_23126);
or UO_526 (O_526,N_22704,N_23934);
nor UO_527 (O_527,N_23986,N_22721);
and UO_528 (O_528,N_24689,N_24280);
nor UO_529 (O_529,N_24804,N_23815);
nor UO_530 (O_530,N_24624,N_24654);
or UO_531 (O_531,N_22527,N_24115);
xor UO_532 (O_532,N_24527,N_23088);
xnor UO_533 (O_533,N_23269,N_23308);
and UO_534 (O_534,N_22549,N_23375);
xnor UO_535 (O_535,N_23124,N_23660);
xor UO_536 (O_536,N_22728,N_24405);
xor UO_537 (O_537,N_23685,N_24790);
nor UO_538 (O_538,N_23885,N_22660);
or UO_539 (O_539,N_23511,N_22610);
nor UO_540 (O_540,N_24443,N_24023);
or UO_541 (O_541,N_24452,N_23605);
or UO_542 (O_542,N_24580,N_24811);
nand UO_543 (O_543,N_24688,N_24028);
nor UO_544 (O_544,N_23287,N_24818);
or UO_545 (O_545,N_24414,N_22941);
or UO_546 (O_546,N_24851,N_24407);
nand UO_547 (O_547,N_23341,N_24561);
nand UO_548 (O_548,N_24312,N_22629);
and UO_549 (O_549,N_24748,N_23092);
nor UO_550 (O_550,N_24986,N_23536);
nor UO_551 (O_551,N_22510,N_23442);
nand UO_552 (O_552,N_22509,N_23327);
xnor UO_553 (O_553,N_23481,N_23186);
or UO_554 (O_554,N_24783,N_23816);
nand UO_555 (O_555,N_24258,N_23955);
or UO_556 (O_556,N_23236,N_23189);
xor UO_557 (O_557,N_24936,N_23192);
nor UO_558 (O_558,N_22676,N_24559);
and UO_559 (O_559,N_24521,N_24653);
and UO_560 (O_560,N_23755,N_23545);
xnor UO_561 (O_561,N_22730,N_23213);
nand UO_562 (O_562,N_24300,N_24792);
xor UO_563 (O_563,N_24371,N_22983);
and UO_564 (O_564,N_23255,N_23253);
nand UO_565 (O_565,N_23950,N_23320);
xor UO_566 (O_566,N_22798,N_23681);
nand UO_567 (O_567,N_22900,N_23889);
and UO_568 (O_568,N_23201,N_23821);
and UO_569 (O_569,N_23081,N_23025);
and UO_570 (O_570,N_24799,N_23242);
or UO_571 (O_571,N_23824,N_23256);
nand UO_572 (O_572,N_22784,N_23318);
or UO_573 (O_573,N_24227,N_23565);
xor UO_574 (O_574,N_23983,N_24315);
or UO_575 (O_575,N_23029,N_24567);
nor UO_576 (O_576,N_23305,N_24534);
nand UO_577 (O_577,N_23506,N_24947);
xnor UO_578 (O_578,N_24039,N_23495);
nand UO_579 (O_579,N_22619,N_23938);
and UO_580 (O_580,N_23151,N_22634);
or UO_581 (O_581,N_23215,N_22709);
nand UO_582 (O_582,N_24327,N_24161);
nor UO_583 (O_583,N_22582,N_23178);
and UO_584 (O_584,N_24318,N_22627);
nand UO_585 (O_585,N_24118,N_24699);
xnor UO_586 (O_586,N_24231,N_23908);
nor UO_587 (O_587,N_24743,N_22575);
or UO_588 (O_588,N_23757,N_24378);
nor UO_589 (O_589,N_24705,N_23246);
xnor UO_590 (O_590,N_23408,N_23913);
nand UO_591 (O_591,N_22922,N_23883);
nor UO_592 (O_592,N_24221,N_23394);
nand UO_593 (O_593,N_23142,N_24772);
or UO_594 (O_594,N_22872,N_24770);
nand UO_595 (O_595,N_23723,N_24806);
nand UO_596 (O_596,N_23795,N_24457);
xnor UO_597 (O_597,N_24814,N_22808);
xor UO_598 (O_598,N_24044,N_22812);
xor UO_599 (O_599,N_22891,N_23593);
and UO_600 (O_600,N_24844,N_24481);
and UO_601 (O_601,N_23570,N_24065);
or UO_602 (O_602,N_23455,N_23997);
xor UO_603 (O_603,N_22822,N_22804);
nor UO_604 (O_604,N_24585,N_23614);
and UO_605 (O_605,N_22675,N_22963);
nor UO_606 (O_606,N_24724,N_22851);
nand UO_607 (O_607,N_23204,N_22920);
and UO_608 (O_608,N_23756,N_23268);
or UO_609 (O_609,N_22931,N_24207);
nor UO_610 (O_610,N_23085,N_24431);
nor UO_611 (O_611,N_24060,N_22860);
nor UO_612 (O_612,N_22617,N_23419);
nor UO_613 (O_613,N_23221,N_23079);
or UO_614 (O_614,N_22668,N_24786);
nor UO_615 (O_615,N_24087,N_23109);
xnor UO_616 (O_616,N_23517,N_24684);
or UO_617 (O_617,N_24556,N_22967);
nor UO_618 (O_618,N_24448,N_23159);
xor UO_619 (O_619,N_23490,N_24350);
or UO_620 (O_620,N_24215,N_24732);
xnor UO_621 (O_621,N_23451,N_23629);
and UO_622 (O_622,N_22917,N_22639);
nor UO_623 (O_623,N_22701,N_23382);
nand UO_624 (O_624,N_22806,N_23173);
nand UO_625 (O_625,N_24949,N_22734);
or UO_626 (O_626,N_24144,N_24196);
nand UO_627 (O_627,N_24694,N_24200);
xor UO_628 (O_628,N_23876,N_24599);
or UO_629 (O_629,N_23552,N_22952);
xnor UO_630 (O_630,N_22514,N_24759);
and UO_631 (O_631,N_24557,N_23659);
xnor UO_632 (O_632,N_24842,N_22586);
nor UO_633 (O_633,N_23022,N_22713);
nand UO_634 (O_634,N_23123,N_24723);
nor UO_635 (O_635,N_22901,N_23065);
and UO_636 (O_636,N_24626,N_24681);
and UO_637 (O_637,N_23886,N_23047);
nor UO_638 (O_638,N_22504,N_24832);
xnor UO_639 (O_639,N_23691,N_23155);
nor UO_640 (O_640,N_22903,N_22667);
nand UO_641 (O_641,N_23878,N_23134);
or UO_642 (O_642,N_24239,N_24622);
nand UO_643 (O_643,N_22778,N_24878);
xnor UO_644 (O_644,N_24095,N_23864);
xor UO_645 (O_645,N_23328,N_23128);
and UO_646 (O_646,N_24442,N_22609);
and UO_647 (O_647,N_24746,N_23252);
xor UO_648 (O_648,N_22526,N_22779);
xor UO_649 (O_649,N_23573,N_22970);
nor UO_650 (O_650,N_24389,N_22712);
xor UO_651 (O_651,N_23608,N_24273);
nor UO_652 (O_652,N_22666,N_23137);
or UO_653 (O_653,N_24834,N_24325);
and UO_654 (O_654,N_23914,N_23711);
nor UO_655 (O_655,N_22780,N_23658);
xnor UO_656 (O_656,N_24989,N_24466);
xnor UO_657 (O_657,N_24426,N_24155);
or UO_658 (O_658,N_23697,N_24031);
nor UO_659 (O_659,N_23648,N_23413);
nand UO_660 (O_660,N_23198,N_23534);
xnor UO_661 (O_661,N_23610,N_23943);
nor UO_662 (O_662,N_22685,N_22670);
nor UO_663 (O_663,N_24206,N_22657);
or UO_664 (O_664,N_23568,N_23129);
and UO_665 (O_665,N_23912,N_24923);
xnor UO_666 (O_666,N_24479,N_22523);
xor UO_667 (O_667,N_24701,N_23404);
nor UO_668 (O_668,N_24009,N_22889);
nand UO_669 (O_669,N_24648,N_24926);
nor UO_670 (O_670,N_24747,N_23715);
nor UO_671 (O_671,N_23541,N_23761);
xnor UO_672 (O_672,N_23440,N_22611);
and UO_673 (O_673,N_23655,N_23738);
xnor UO_674 (O_674,N_24498,N_24377);
or UO_675 (O_675,N_24364,N_23782);
and UO_676 (O_676,N_23431,N_24941);
nor UO_677 (O_677,N_22604,N_24376);
and UO_678 (O_678,N_23008,N_22799);
and UO_679 (O_679,N_23266,N_24112);
nor UO_680 (O_680,N_24284,N_24946);
or UO_681 (O_681,N_23210,N_23870);
xor UO_682 (O_682,N_23334,N_24423);
and UO_683 (O_683,N_23247,N_23917);
or UO_684 (O_684,N_23526,N_24114);
nand UO_685 (O_685,N_23244,N_24727);
or UO_686 (O_686,N_23776,N_22826);
or UO_687 (O_687,N_24101,N_24422);
and UO_688 (O_688,N_24510,N_24895);
nor UO_689 (O_689,N_23577,N_23828);
xor UO_690 (O_690,N_22558,N_24146);
nor UO_691 (O_691,N_24934,N_23714);
nor UO_692 (O_692,N_24817,N_23930);
and UO_693 (O_693,N_22732,N_22710);
or UO_694 (O_694,N_22982,N_24717);
or UO_695 (O_695,N_23906,N_24883);
and UO_696 (O_696,N_23043,N_23910);
nor UO_697 (O_697,N_23865,N_24138);
or UO_698 (O_698,N_24862,N_23400);
xor UO_699 (O_699,N_24597,N_24555);
nand UO_700 (O_700,N_22783,N_23317);
xnor UO_701 (O_701,N_22750,N_22596);
or UO_702 (O_702,N_24531,N_23426);
or UO_703 (O_703,N_22774,N_22684);
xor UO_704 (O_704,N_24924,N_22974);
and UO_705 (O_705,N_23003,N_23310);
nor UO_706 (O_706,N_24293,N_22991);
or UO_707 (O_707,N_23316,N_23039);
or UO_708 (O_708,N_23628,N_24444);
nor UO_709 (O_709,N_24864,N_23054);
nor UO_710 (O_710,N_23902,N_22942);
xnor UO_711 (O_711,N_23286,N_24776);
nand UO_712 (O_712,N_24607,N_23635);
xnor UO_713 (O_713,N_23463,N_23904);
nor UO_714 (O_714,N_23721,N_24590);
nand UO_715 (O_715,N_24973,N_23131);
or UO_716 (O_716,N_23459,N_24977);
nand UO_717 (O_717,N_23323,N_24153);
xor UO_718 (O_718,N_22548,N_22651);
xor UO_719 (O_719,N_22689,N_23592);
nand UO_720 (O_720,N_22706,N_24421);
or UO_721 (O_721,N_22691,N_23984);
nor UO_722 (O_722,N_24605,N_22569);
xor UO_723 (O_723,N_23649,N_23336);
nand UO_724 (O_724,N_22781,N_24970);
or UO_725 (O_725,N_24150,N_23531);
xnor UO_726 (O_726,N_24159,N_23785);
xor UO_727 (O_727,N_23728,N_22614);
nand UO_728 (O_728,N_23720,N_23990);
xor UO_729 (O_729,N_24334,N_24951);
xor UO_730 (O_730,N_24921,N_23453);
nor UO_731 (O_731,N_24975,N_24507);
xnor UO_732 (O_732,N_23678,N_24726);
or UO_733 (O_733,N_22768,N_22791);
xnor UO_734 (O_734,N_24126,N_24254);
and UO_735 (O_735,N_22836,N_22987);
xnor UO_736 (O_736,N_23084,N_22718);
and UO_737 (O_737,N_23973,N_22513);
nor UO_738 (O_738,N_22869,N_23674);
xor UO_739 (O_739,N_23709,N_23976);
and UO_740 (O_740,N_24130,N_23819);
nor UO_741 (O_741,N_23216,N_24346);
xnor UO_742 (O_742,N_24641,N_23169);
nand UO_743 (O_743,N_24314,N_23829);
xor UO_744 (O_744,N_23469,N_23489);
nand UO_745 (O_745,N_24802,N_24177);
xor UO_746 (O_746,N_24400,N_24793);
nand UO_747 (O_747,N_24156,N_22748);
nand UO_748 (O_748,N_22915,N_23080);
and UO_749 (O_749,N_22989,N_22758);
xnor UO_750 (O_750,N_23503,N_24586);
xor UO_751 (O_751,N_23423,N_23272);
or UO_752 (O_752,N_23207,N_24213);
and UO_753 (O_753,N_23642,N_22645);
and UO_754 (O_754,N_23540,N_24089);
or UO_755 (O_755,N_23974,N_23616);
xor UO_756 (O_756,N_23415,N_22892);
and UO_757 (O_757,N_24275,N_24323);
and UO_758 (O_758,N_23473,N_24757);
and UO_759 (O_759,N_23641,N_22737);
nor UO_760 (O_760,N_24458,N_23433);
and UO_761 (O_761,N_23067,N_24663);
nor UO_762 (O_762,N_23716,N_24445);
xor UO_763 (O_763,N_24420,N_24286);
nor UO_764 (O_764,N_24105,N_22858);
nand UO_765 (O_765,N_23429,N_23018);
or UO_766 (O_766,N_23100,N_24288);
nor UO_767 (O_767,N_24940,N_22765);
and UO_768 (O_768,N_23611,N_24187);
nor UO_769 (O_769,N_23232,N_24929);
and UO_770 (O_770,N_23603,N_24565);
and UO_771 (O_771,N_23957,N_24292);
nor UO_772 (O_772,N_24815,N_23389);
or UO_773 (O_773,N_23946,N_23615);
nor UO_774 (O_774,N_24712,N_24397);
or UO_775 (O_775,N_23765,N_23667);
xnor UO_776 (O_776,N_23099,N_23050);
or UO_777 (O_777,N_23556,N_24920);
nand UO_778 (O_778,N_24478,N_24836);
nor UO_779 (O_779,N_22649,N_24579);
and UO_780 (O_780,N_22878,N_23145);
nor UO_781 (O_781,N_22735,N_24560);
nand UO_782 (O_782,N_23195,N_23528);
nor UO_783 (O_783,N_24427,N_23254);
nand UO_784 (O_784,N_23301,N_23474);
xor UO_785 (O_785,N_23202,N_23808);
nor UO_786 (O_786,N_23509,N_24816);
nor UO_787 (O_787,N_23006,N_23108);
or UO_788 (O_788,N_24082,N_23239);
xor UO_789 (O_789,N_23880,N_23017);
and UO_790 (O_790,N_23790,N_24656);
nor UO_791 (O_791,N_24488,N_24668);
nand UO_792 (O_792,N_22795,N_23418);
nand UO_793 (O_793,N_23464,N_24928);
xnor UO_794 (O_794,N_23571,N_23595);
and UO_795 (O_795,N_22512,N_22632);
or UO_796 (O_796,N_24109,N_23794);
nand UO_797 (O_797,N_24406,N_23909);
or UO_798 (O_798,N_24779,N_24637);
or UO_799 (O_799,N_24778,N_24672);
or UO_800 (O_800,N_23734,N_23800);
or UO_801 (O_801,N_22905,N_23230);
or UO_802 (O_802,N_23797,N_24543);
nand UO_803 (O_803,N_24113,N_23703);
nand UO_804 (O_804,N_24886,N_24917);
xor UO_805 (O_805,N_23951,N_24368);
nor UO_806 (O_806,N_24326,N_22716);
or UO_807 (O_807,N_23512,N_23839);
or UO_808 (O_808,N_23535,N_23848);
nor UO_809 (O_809,N_24533,N_24083);
nand UO_810 (O_810,N_24216,N_24763);
nand UO_811 (O_811,N_23248,N_23804);
xnor UO_812 (O_812,N_24525,N_24948);
or UO_813 (O_813,N_23546,N_23846);
or UO_814 (O_814,N_23664,N_24959);
and UO_815 (O_815,N_23602,N_22723);
and UO_816 (O_816,N_23837,N_23779);
and UO_817 (O_817,N_22828,N_24503);
nand UO_818 (O_818,N_24055,N_23471);
nand UO_819 (O_819,N_23468,N_23522);
or UO_820 (O_820,N_22864,N_24913);
nor UO_821 (O_821,N_23689,N_24505);
nor UO_822 (O_822,N_23214,N_24906);
and UO_823 (O_823,N_23746,N_24957);
and UO_824 (O_824,N_23330,N_23740);
nand UO_825 (O_825,N_23146,N_23532);
and UO_826 (O_826,N_24016,N_23786);
nand UO_827 (O_827,N_24163,N_24192);
or UO_828 (O_828,N_24502,N_23825);
nand UO_829 (O_829,N_24497,N_23970);
nand UO_830 (O_830,N_24939,N_24049);
nand UO_831 (O_831,N_24718,N_23935);
nand UO_832 (O_832,N_23063,N_23820);
or UO_833 (O_833,N_23514,N_24347);
nand UO_834 (O_834,N_24984,N_23160);
nand UO_835 (O_835,N_22561,N_22568);
nand UO_836 (O_836,N_23926,N_23948);
xnor UO_837 (O_837,N_24434,N_24037);
and UO_838 (O_838,N_24245,N_23722);
nor UO_839 (O_839,N_24392,N_24693);
xor UO_840 (O_840,N_23051,N_24524);
nor UO_841 (O_841,N_24285,N_24715);
and UO_842 (O_842,N_24769,N_22747);
nand UO_843 (O_843,N_24901,N_23098);
nor UO_844 (O_844,N_24048,N_23012);
nor UO_845 (O_845,N_23684,N_24897);
nand UO_846 (O_846,N_23302,N_23071);
nand UO_847 (O_847,N_24360,N_24885);
nor UO_848 (O_848,N_22857,N_24291);
xor UO_849 (O_849,N_23066,N_23843);
nor UO_850 (O_850,N_24698,N_24219);
or UO_851 (O_851,N_23515,N_24298);
nand UO_852 (O_852,N_24450,N_24173);
or UO_853 (O_853,N_24544,N_23962);
and UO_854 (O_854,N_23331,N_22865);
nor UO_855 (O_855,N_24514,N_24279);
nor UO_856 (O_856,N_24600,N_24047);
nor UO_857 (O_857,N_23567,N_22842);
or UO_858 (O_858,N_24679,N_24046);
nand UO_859 (O_859,N_24801,N_22976);
and UO_860 (O_860,N_22697,N_24665);
and UO_861 (O_861,N_24353,N_22673);
xnor UO_862 (O_862,N_24224,N_23929);
xnor UO_863 (O_863,N_24785,N_24632);
nor UO_864 (O_864,N_23157,N_23805);
and UO_865 (O_865,N_24664,N_23998);
and UO_866 (O_866,N_24419,N_23524);
xor UO_867 (O_867,N_23427,N_23010);
or UO_868 (O_868,N_24190,N_24463);
or UO_869 (O_869,N_24062,N_24552);
and UO_870 (O_870,N_22825,N_22692);
nor UO_871 (O_871,N_24297,N_22824);
and UO_872 (O_872,N_23505,N_22953);
or UO_873 (O_873,N_23977,N_23594);
xnor UO_874 (O_874,N_23061,N_22711);
and UO_875 (O_875,N_24703,N_23609);
xnor UO_876 (O_876,N_23399,N_24167);
nand UO_877 (O_877,N_23581,N_22815);
xnor UO_878 (O_878,N_24352,N_23414);
xnor UO_879 (O_879,N_23665,N_22729);
and UO_880 (O_880,N_23733,N_23792);
or UO_881 (O_881,N_23297,N_24687);
xor UO_882 (O_882,N_24178,N_24418);
nand UO_883 (O_883,N_23156,N_24296);
and UO_884 (O_884,N_22959,N_22775);
and UO_885 (O_885,N_24181,N_23967);
nand UO_886 (O_886,N_23211,N_24962);
or UO_887 (O_887,N_23119,N_23258);
nor UO_888 (O_888,N_23007,N_24902);
or UO_889 (O_889,N_23203,N_24253);
nor UO_890 (O_890,N_23150,N_24491);
nand UO_891 (O_891,N_24324,N_22910);
xnor UO_892 (O_892,N_24343,N_24849);
or UO_893 (O_893,N_24099,N_24880);
nor UO_894 (O_894,N_23580,N_23369);
xor UO_895 (O_895,N_23700,N_24250);
or UO_896 (O_896,N_22544,N_23115);
nand UO_897 (O_897,N_23319,N_24372);
nand UO_898 (O_898,N_24553,N_24136);
xor UO_899 (O_899,N_23226,N_23056);
nand UO_900 (O_900,N_22772,N_24891);
nand UO_901 (O_901,N_23089,N_24011);
nor UO_902 (O_902,N_24366,N_24229);
nor UO_903 (O_903,N_24961,N_23923);
xnor UO_904 (O_904,N_23136,N_24782);
and UO_905 (O_905,N_23352,N_24710);
nor UO_906 (O_906,N_24132,N_24621);
or UO_907 (O_907,N_23299,N_24967);
nor UO_908 (O_908,N_24690,N_23704);
or UO_909 (O_909,N_23270,N_24669);
nor UO_910 (O_910,N_22547,N_24390);
nand UO_911 (O_911,N_23881,N_24667);
nor UO_912 (O_912,N_24456,N_22909);
or UO_913 (O_913,N_22647,N_24437);
nand UO_914 (O_914,N_23295,N_24647);
xor UO_915 (O_915,N_23763,N_24247);
or UO_916 (O_916,N_22919,N_22807);
xnor UO_917 (O_917,N_22608,N_23031);
xnor UO_918 (O_918,N_24123,N_24686);
nand UO_919 (O_919,N_24086,N_24609);
xnor UO_920 (O_920,N_22580,N_23586);
xnor UO_921 (O_921,N_23162,N_23560);
xnor UO_922 (O_922,N_23954,N_24453);
xnor UO_923 (O_923,N_23959,N_23875);
xor UO_924 (O_924,N_23894,N_23979);
nand UO_925 (O_925,N_22814,N_24905);
and UO_926 (O_926,N_24257,N_24875);
and UO_927 (O_927,N_23561,N_23831);
nor UO_928 (O_928,N_24125,N_23231);
or UO_929 (O_929,N_24246,N_24766);
or UO_930 (O_930,N_24919,N_24329);
nor UO_931 (O_931,N_23862,N_23830);
xor UO_932 (O_932,N_23690,N_22921);
xnor UO_933 (O_933,N_23424,N_23454);
xnor UO_934 (O_934,N_23095,N_23589);
or UO_935 (O_935,N_24010,N_24837);
nand UO_936 (O_936,N_24094,N_24596);
and UO_937 (O_937,N_24302,N_22935);
nor UO_938 (O_938,N_22850,N_24290);
or UO_939 (O_939,N_24861,N_23666);
nor UO_940 (O_940,N_23177,N_23458);
nand UO_941 (O_941,N_23652,N_24630);
nor UO_942 (O_942,N_24828,N_23724);
or UO_943 (O_943,N_24640,N_23140);
xnor UO_944 (O_944,N_24034,N_23026);
nand UO_945 (O_945,N_23417,N_23680);
nor UO_946 (O_946,N_24230,N_24870);
and UO_947 (O_947,N_23465,N_23307);
nor UO_948 (O_948,N_22736,N_23840);
xor UO_949 (O_949,N_24958,N_24035);
or UO_950 (O_950,N_24172,N_22745);
xnor UO_951 (O_951,N_24639,N_23521);
nor UO_952 (O_952,N_22650,N_23163);
nand UO_953 (O_953,N_23125,N_24467);
or UO_954 (O_954,N_24472,N_22695);
and UO_955 (O_955,N_24234,N_24835);
or UO_956 (O_956,N_22911,N_22601);
xnor UO_957 (O_957,N_24120,N_22633);
and UO_958 (O_958,N_23439,N_23799);
and UO_959 (O_959,N_23947,N_23989);
and UO_960 (O_960,N_24072,N_23661);
nor UO_961 (O_961,N_24486,N_22687);
or UO_962 (O_962,N_23739,N_23233);
xnor UO_963 (O_963,N_24981,N_22980);
or UO_964 (O_964,N_24179,N_24205);
or UO_965 (O_965,N_24629,N_23113);
nand UO_966 (O_966,N_24819,N_24128);
xor UO_967 (O_967,N_24736,N_22984);
or UO_968 (O_968,N_24536,N_23144);
xnor UO_969 (O_969,N_24511,N_24005);
nand UO_970 (O_970,N_23185,N_23002);
xnor UO_971 (O_971,N_24097,N_24691);
and UO_972 (O_972,N_23372,N_23633);
nand UO_973 (O_973,N_24256,N_24978);
xor UO_974 (O_974,N_24572,N_24898);
nand UO_975 (O_975,N_23753,N_24424);
and UO_976 (O_976,N_24030,N_22763);
or UO_977 (O_977,N_23132,N_24212);
and UO_978 (O_978,N_23783,N_22528);
or UO_979 (O_979,N_23196,N_23563);
nand UO_980 (O_980,N_22936,N_22766);
nand UO_981 (O_981,N_24623,N_24601);
nand UO_982 (O_982,N_23773,N_23542);
nor UO_983 (O_983,N_22603,N_22943);
or UO_984 (O_984,N_22588,N_24731);
nor UO_985 (O_985,N_24520,N_23916);
or UO_986 (O_986,N_24860,N_22644);
nor UO_987 (O_987,N_24613,N_24002);
or UO_988 (O_988,N_23212,N_24383);
and UO_989 (O_989,N_23324,N_23281);
xor UO_990 (O_990,N_23712,N_23467);
and UO_991 (O_991,N_23784,N_24998);
or UO_992 (O_992,N_23234,N_23699);
xor UO_993 (O_993,N_24935,N_24850);
nand UO_994 (O_994,N_23850,N_24966);
nor UO_995 (O_995,N_22977,N_22690);
xor UO_996 (O_996,N_22854,N_24363);
or UO_997 (O_997,N_23928,N_24646);
and UO_998 (O_998,N_23588,N_22913);
xor UO_999 (O_999,N_24749,N_22598);
xor UO_1000 (O_1000,N_24899,N_24308);
xnor UO_1001 (O_1001,N_24593,N_24740);
nor UO_1002 (O_1002,N_24584,N_22939);
nand UO_1003 (O_1003,N_24908,N_22564);
xnor UO_1004 (O_1004,N_23359,N_23072);
nand UO_1005 (O_1005,N_24582,N_24211);
and UO_1006 (O_1006,N_23918,N_24428);
nor UO_1007 (O_1007,N_24513,N_23768);
or UO_1008 (O_1008,N_24204,N_23395);
and UO_1009 (O_1009,N_24628,N_24578);
xor UO_1010 (O_1010,N_24451,N_24537);
xor UO_1011 (O_1011,N_22843,N_24655);
or UO_1012 (O_1012,N_24714,N_23555);
and UO_1013 (O_1013,N_24541,N_24796);
nand UO_1014 (O_1014,N_24464,N_22522);
nor UO_1015 (O_1015,N_24566,N_23729);
nand UO_1016 (O_1016,N_23789,N_23430);
xnor UO_1017 (O_1017,N_23513,N_22742);
nand UO_1018 (O_1018,N_24564,N_23339);
or UO_1019 (O_1019,N_24765,N_24362);
or UO_1020 (O_1020,N_24483,N_24058);
and UO_1021 (O_1021,N_22755,N_22674);
nand UO_1022 (O_1022,N_23483,N_23606);
or UO_1023 (O_1023,N_22886,N_23052);
and UO_1024 (O_1024,N_23165,N_24839);
xor UO_1025 (O_1025,N_22722,N_24379);
or UO_1026 (O_1026,N_23472,N_24077);
xor UO_1027 (O_1027,N_24042,N_23683);
nor UO_1028 (O_1028,N_24820,N_24716);
nor UO_1029 (O_1029,N_24985,N_22628);
nor UO_1030 (O_1030,N_23644,N_23030);
nand UO_1031 (O_1031,N_23537,N_23312);
or UO_1032 (O_1032,N_24317,N_24912);
or UO_1033 (O_1033,N_24789,N_23519);
xor UO_1034 (O_1034,N_24598,N_22597);
nor UO_1035 (O_1035,N_22964,N_23193);
nor UO_1036 (O_1036,N_24678,N_22605);
and UO_1037 (O_1037,N_22961,N_24602);
nor UO_1038 (O_1038,N_24704,N_22955);
and UO_1039 (O_1039,N_23298,N_24997);
xnor UO_1040 (O_1040,N_24773,N_23562);
and UO_1041 (O_1041,N_24767,N_24384);
or UO_1042 (O_1042,N_23933,N_23854);
and UO_1043 (O_1043,N_24045,N_22800);
or UO_1044 (O_1044,N_23749,N_22719);
or UO_1045 (O_1045,N_22767,N_22606);
and UO_1046 (O_1046,N_23436,N_22556);
nand UO_1047 (O_1047,N_24863,N_23484);
xor UO_1048 (O_1048,N_24170,N_22626);
nor UO_1049 (O_1049,N_24024,N_24081);
xor UO_1050 (O_1050,N_23682,N_24321);
xor UO_1051 (O_1051,N_23624,N_23325);
or UO_1052 (O_1052,N_24470,N_23401);
or UO_1053 (O_1053,N_23164,N_24357);
and UO_1054 (O_1054,N_23987,N_22896);
xnor UO_1055 (O_1055,N_23220,N_24810);
or UO_1056 (O_1056,N_23775,N_22738);
or UO_1057 (O_1057,N_24359,N_23356);
xnor UO_1058 (O_1058,N_23899,N_24303);
xor UO_1059 (O_1059,N_24158,N_22624);
nand UO_1060 (O_1060,N_22881,N_23452);
and UO_1061 (O_1061,N_24872,N_23745);
and UO_1062 (O_1062,N_23009,N_23941);
xor UO_1063 (O_1063,N_24455,N_22962);
nand UO_1064 (O_1064,N_24339,N_23992);
or UO_1065 (O_1065,N_23803,N_24393);
xnor UO_1066 (O_1066,N_22550,N_24367);
and UO_1067 (O_1067,N_22744,N_23936);
xnor UO_1068 (O_1068,N_24000,N_24869);
xnor UO_1069 (O_1069,N_24252,N_23539);
nor UO_1070 (O_1070,N_23643,N_24139);
nor UO_1071 (O_1071,N_22653,N_23504);
nor UO_1072 (O_1072,N_24618,N_23958);
or UO_1073 (O_1073,N_22515,N_22918);
or UO_1074 (O_1074,N_24306,N_24266);
nand UO_1075 (O_1075,N_22874,N_23798);
and UO_1076 (O_1076,N_24168,N_22793);
or UO_1077 (O_1077,N_23855,N_23371);
nor UO_1078 (O_1078,N_23152,N_23780);
nor UO_1079 (O_1079,N_24494,N_23340);
nor UO_1080 (O_1080,N_23337,N_22595);
xor UO_1081 (O_1081,N_22511,N_24465);
xor UO_1082 (O_1082,N_24523,N_23138);
xnor UO_1083 (O_1083,N_22579,N_22839);
xnor UO_1084 (O_1084,N_24142,N_22664);
and UO_1085 (O_1085,N_22841,N_23000);
nand UO_1086 (O_1086,N_22593,N_23333);
and UO_1087 (O_1087,N_24952,N_23501);
xor UO_1088 (O_1088,N_23013,N_23217);
nand UO_1089 (O_1089,N_23405,N_23206);
nand UO_1090 (O_1090,N_22620,N_23551);
nor UO_1091 (O_1091,N_23432,N_23180);
nand UO_1092 (O_1092,N_23793,N_23373);
and UO_1093 (O_1093,N_22554,N_22944);
and UO_1094 (O_1094,N_23342,N_24263);
nor UO_1095 (O_1095,N_23329,N_24542);
nor UO_1096 (O_1096,N_23376,N_24963);
nor UO_1097 (O_1097,N_24858,N_24485);
nand UO_1098 (O_1098,N_23326,N_23480);
or UO_1099 (O_1099,N_24954,N_23668);
and UO_1100 (O_1100,N_24825,N_22871);
xnor UO_1101 (O_1101,N_24354,N_24477);
nor UO_1102 (O_1102,N_24433,N_22810);
xor UO_1103 (O_1103,N_22876,N_24812);
or UO_1104 (O_1104,N_22659,N_24700);
xor UO_1105 (O_1105,N_24098,N_24235);
nor UO_1106 (O_1106,N_24480,N_24879);
or UO_1107 (O_1107,N_22856,N_23686);
and UO_1108 (O_1108,N_24013,N_24032);
and UO_1109 (O_1109,N_23282,N_24004);
or UO_1110 (O_1110,N_24401,N_22707);
and UO_1111 (O_1111,N_24394,N_23601);
nand UO_1112 (O_1112,N_24994,N_24821);
nor UO_1113 (O_1113,N_23120,N_23847);
nand UO_1114 (O_1114,N_23874,N_24888);
nand UO_1115 (O_1115,N_24709,N_22529);
nand UO_1116 (O_1116,N_22960,N_23901);
or UO_1117 (O_1117,N_24651,N_22832);
xor UO_1118 (O_1118,N_23057,N_24867);
xnor UO_1119 (O_1119,N_22574,N_24822);
or UO_1120 (O_1120,N_23827,N_23351);
xnor UO_1121 (O_1121,N_24313,N_23182);
xnor UO_1122 (O_1122,N_23219,N_24562);
or UO_1123 (O_1123,N_23743,N_24614);
nand UO_1124 (O_1124,N_24964,N_24522);
and UO_1125 (O_1125,N_23391,N_24269);
nor UO_1126 (O_1126,N_24657,N_22813);
nand UO_1127 (O_1127,N_22787,N_24549);
nor UO_1128 (O_1128,N_23818,N_23777);
nand UO_1129 (O_1129,N_24945,N_24570);
nand UO_1130 (O_1130,N_24991,N_22537);
or UO_1131 (O_1131,N_24017,N_24515);
and UO_1132 (O_1132,N_24910,N_23492);
or UO_1133 (O_1133,N_22702,N_23407);
nor UO_1134 (O_1134,N_24887,N_24404);
nand UO_1135 (O_1135,N_23205,N_22831);
nor UO_1136 (O_1136,N_23502,N_24137);
nor UO_1137 (O_1137,N_23073,N_23199);
and UO_1138 (O_1138,N_24117,N_23851);
and UO_1139 (O_1139,N_23290,N_23915);
nand UO_1140 (O_1140,N_22584,N_24267);
and UO_1141 (O_1141,N_24001,N_23406);
xor UO_1142 (O_1142,N_22994,N_24345);
nor UO_1143 (O_1143,N_22618,N_24237);
nor UO_1144 (O_1144,N_23867,N_24506);
or UO_1145 (O_1145,N_22740,N_23251);
or UO_1146 (O_1146,N_23222,N_23175);
nor UO_1147 (O_1147,N_24868,N_22545);
or UO_1148 (O_1148,N_24036,N_24484);
nand UO_1149 (O_1149,N_22662,N_23096);
nor UO_1150 (O_1150,N_23507,N_23778);
and UO_1151 (O_1151,N_22867,N_24492);
nand UO_1152 (O_1152,N_24386,N_22533);
and UO_1153 (O_1153,N_24140,N_23355);
nor UO_1154 (O_1154,N_24336,N_24259);
nand UO_1155 (O_1155,N_24461,N_24149);
nor UO_1156 (O_1156,N_23332,N_23315);
or UO_1157 (O_1157,N_24381,N_23694);
nand UO_1158 (O_1158,N_23654,N_22957);
xor UO_1159 (O_1159,N_24733,N_22761);
or UO_1160 (O_1160,N_24482,N_23364);
nand UO_1161 (O_1161,N_23181,N_23952);
nand UO_1162 (O_1162,N_22636,N_22591);
nor UO_1163 (O_1163,N_24865,N_24840);
and UO_1164 (O_1164,N_23167,N_24972);
xor UO_1165 (O_1165,N_24938,N_22607);
and UO_1166 (O_1166,N_22587,N_22756);
and UO_1167 (O_1167,N_23033,N_23543);
xor UO_1168 (O_1168,N_23549,N_22757);
xor UO_1169 (O_1169,N_23860,N_23996);
xnor UO_1170 (O_1170,N_24435,N_23995);
xor UO_1171 (O_1171,N_24309,N_24388);
or UO_1172 (O_1172,N_22880,N_24412);
nand UO_1173 (O_1173,N_23042,N_24638);
xnor UO_1174 (O_1174,N_22816,N_23243);
or UO_1175 (O_1175,N_23462,N_23566);
and UO_1176 (O_1176,N_22908,N_23758);
and UO_1177 (O_1177,N_24188,N_24671);
nor UO_1178 (O_1178,N_22914,N_23760);
and UO_1179 (O_1179,N_23179,N_23701);
and UO_1180 (O_1180,N_23350,N_24942);
and UO_1181 (O_1181,N_23311,N_23806);
xnor UO_1182 (O_1182,N_23087,N_22625);
or UO_1183 (O_1183,N_23497,N_24051);
xnor UO_1184 (O_1184,N_24692,N_24100);
nand UO_1185 (O_1185,N_23135,N_24581);
nor UO_1186 (O_1186,N_23845,N_23822);
xnor UO_1187 (O_1187,N_23590,N_23487);
nand UO_1188 (O_1188,N_24274,N_23817);
nand UO_1189 (O_1189,N_23273,N_24965);
nand UO_1190 (O_1190,N_23922,N_24402);
and UO_1191 (O_1191,N_24429,N_22870);
nor UO_1192 (O_1192,N_22648,N_23835);
and UO_1193 (O_1193,N_24999,N_23558);
and UO_1194 (O_1194,N_24225,N_23357);
nor UO_1195 (O_1195,N_22572,N_24636);
or UO_1196 (O_1196,N_24129,N_24436);
nand UO_1197 (O_1197,N_23632,N_24813);
nor UO_1198 (O_1198,N_24501,N_22520);
nor UO_1199 (O_1199,N_24217,N_23858);
and UO_1200 (O_1200,N_23774,N_22538);
or UO_1201 (O_1201,N_24944,N_23049);
and UO_1202 (O_1202,N_23011,N_24838);
and UO_1203 (O_1203,N_22600,N_23725);
and UO_1204 (O_1204,N_24121,N_24927);
and UO_1205 (O_1205,N_24877,N_23942);
and UO_1206 (O_1206,N_24147,N_24720);
and UO_1207 (O_1207,N_24532,N_24847);
xnor UO_1208 (O_1208,N_23891,N_23623);
xor UO_1209 (O_1209,N_23713,N_24988);
xor UO_1210 (O_1210,N_24761,N_23695);
nand UO_1211 (O_1211,N_23636,N_23520);
nor UO_1212 (O_1212,N_22517,N_23639);
nor UO_1213 (O_1213,N_23859,N_24026);
nor UO_1214 (O_1214,N_22658,N_23118);
xor UO_1215 (O_1215,N_23362,N_23810);
xnor UO_1216 (O_1216,N_23488,N_23379);
xor UO_1217 (O_1217,N_24335,N_23174);
and UO_1218 (O_1218,N_23553,N_23265);
nand UO_1219 (O_1219,N_23378,N_23086);
nor UO_1220 (O_1220,N_22853,N_23122);
nand UO_1221 (O_1221,N_24185,N_23470);
or UO_1222 (O_1222,N_24659,N_23651);
and UO_1223 (O_1223,N_22576,N_24768);
nor UO_1224 (O_1224,N_23335,N_24489);
and UO_1225 (O_1225,N_22680,N_23238);
and UO_1226 (O_1226,N_22519,N_22615);
xnor UO_1227 (O_1227,N_24493,N_23741);
nand UO_1228 (O_1228,N_24683,N_24425);
nand UO_1229 (O_1229,N_24064,N_22622);
nor UO_1230 (O_1230,N_23074,N_24758);
xor UO_1231 (O_1231,N_23435,N_23059);
and UO_1232 (O_1232,N_23771,N_23293);
or UO_1233 (O_1233,N_24660,N_22820);
nor UO_1234 (O_1234,N_23262,N_24612);
nand UO_1235 (O_1235,N_23564,N_24008);
xor UO_1236 (O_1236,N_22669,N_23708);
xnor UO_1237 (O_1237,N_24475,N_24316);
xnor UO_1238 (O_1238,N_23313,N_24409);
or UO_1239 (O_1239,N_24063,N_23999);
xnor UO_1240 (O_1240,N_24251,N_22802);
nand UO_1241 (O_1241,N_22508,N_23292);
nor UO_1242 (O_1242,N_23726,N_24116);
and UO_1243 (O_1243,N_23944,N_23304);
or UO_1244 (O_1244,N_22536,N_24131);
nor UO_1245 (O_1245,N_24330,N_23275);
xor UO_1246 (O_1246,N_22932,N_23046);
or UO_1247 (O_1247,N_23718,N_23905);
xnor UO_1248 (O_1248,N_22770,N_24411);
and UO_1249 (O_1249,N_24960,N_22623);
nand UO_1250 (O_1250,N_23273,N_23985);
or UO_1251 (O_1251,N_22585,N_23309);
or UO_1252 (O_1252,N_22677,N_23492);
nand UO_1253 (O_1253,N_22511,N_23539);
or UO_1254 (O_1254,N_23079,N_23413);
nor UO_1255 (O_1255,N_24180,N_23660);
xnor UO_1256 (O_1256,N_23860,N_23950);
or UO_1257 (O_1257,N_24872,N_22675);
xor UO_1258 (O_1258,N_23072,N_23104);
nor UO_1259 (O_1259,N_22817,N_23995);
or UO_1260 (O_1260,N_24350,N_24130);
or UO_1261 (O_1261,N_22886,N_22828);
xor UO_1262 (O_1262,N_24008,N_24786);
nor UO_1263 (O_1263,N_22759,N_23088);
nor UO_1264 (O_1264,N_23968,N_23477);
xnor UO_1265 (O_1265,N_24673,N_24640);
and UO_1266 (O_1266,N_23920,N_24509);
nor UO_1267 (O_1267,N_24013,N_24646);
or UO_1268 (O_1268,N_24654,N_24233);
or UO_1269 (O_1269,N_23983,N_24945);
xor UO_1270 (O_1270,N_24837,N_22775);
nor UO_1271 (O_1271,N_23198,N_22606);
nor UO_1272 (O_1272,N_23082,N_23754);
and UO_1273 (O_1273,N_22864,N_23529);
and UO_1274 (O_1274,N_23790,N_24134);
xnor UO_1275 (O_1275,N_22732,N_23228);
xnor UO_1276 (O_1276,N_24041,N_24381);
xnor UO_1277 (O_1277,N_24098,N_24015);
nand UO_1278 (O_1278,N_24817,N_24340);
nor UO_1279 (O_1279,N_24528,N_24839);
or UO_1280 (O_1280,N_24984,N_22777);
nand UO_1281 (O_1281,N_23280,N_23176);
nand UO_1282 (O_1282,N_22873,N_24257);
nor UO_1283 (O_1283,N_23880,N_23738);
and UO_1284 (O_1284,N_24905,N_24944);
nor UO_1285 (O_1285,N_22521,N_23567);
and UO_1286 (O_1286,N_24418,N_23483);
or UO_1287 (O_1287,N_22584,N_23603);
and UO_1288 (O_1288,N_23979,N_23521);
and UO_1289 (O_1289,N_23786,N_23311);
xor UO_1290 (O_1290,N_22874,N_24299);
nand UO_1291 (O_1291,N_24250,N_23611);
or UO_1292 (O_1292,N_24027,N_23225);
xor UO_1293 (O_1293,N_24579,N_23613);
and UO_1294 (O_1294,N_22548,N_24793);
or UO_1295 (O_1295,N_24035,N_23683);
nor UO_1296 (O_1296,N_24386,N_23398);
or UO_1297 (O_1297,N_22510,N_24988);
and UO_1298 (O_1298,N_24117,N_23118);
nand UO_1299 (O_1299,N_24137,N_23386);
nor UO_1300 (O_1300,N_24013,N_24931);
or UO_1301 (O_1301,N_23623,N_24025);
or UO_1302 (O_1302,N_23771,N_22526);
nor UO_1303 (O_1303,N_24781,N_23103);
and UO_1304 (O_1304,N_22736,N_24244);
nor UO_1305 (O_1305,N_24258,N_24399);
and UO_1306 (O_1306,N_24640,N_23117);
xor UO_1307 (O_1307,N_23430,N_23176);
nor UO_1308 (O_1308,N_24275,N_23071);
nor UO_1309 (O_1309,N_22735,N_24910);
nor UO_1310 (O_1310,N_23760,N_24193);
or UO_1311 (O_1311,N_23621,N_23687);
xor UO_1312 (O_1312,N_24335,N_22572);
nand UO_1313 (O_1313,N_24427,N_24441);
nor UO_1314 (O_1314,N_24822,N_22924);
nand UO_1315 (O_1315,N_24262,N_24337);
and UO_1316 (O_1316,N_23126,N_22621);
and UO_1317 (O_1317,N_24336,N_22593);
nand UO_1318 (O_1318,N_22660,N_23157);
and UO_1319 (O_1319,N_24031,N_23493);
xnor UO_1320 (O_1320,N_22873,N_24193);
or UO_1321 (O_1321,N_24505,N_23105);
nor UO_1322 (O_1322,N_23147,N_22972);
nor UO_1323 (O_1323,N_24748,N_24081);
xnor UO_1324 (O_1324,N_24044,N_23596);
nand UO_1325 (O_1325,N_24445,N_23830);
and UO_1326 (O_1326,N_24127,N_22571);
xnor UO_1327 (O_1327,N_23722,N_23185);
xor UO_1328 (O_1328,N_24263,N_24726);
and UO_1329 (O_1329,N_24901,N_24953);
nor UO_1330 (O_1330,N_22571,N_23109);
nor UO_1331 (O_1331,N_24730,N_24626);
and UO_1332 (O_1332,N_23712,N_22757);
nand UO_1333 (O_1333,N_24985,N_23911);
and UO_1334 (O_1334,N_24313,N_24505);
nor UO_1335 (O_1335,N_24356,N_23271);
nor UO_1336 (O_1336,N_24017,N_23302);
xnor UO_1337 (O_1337,N_23909,N_23222);
or UO_1338 (O_1338,N_22632,N_24377);
nor UO_1339 (O_1339,N_24461,N_24138);
nor UO_1340 (O_1340,N_23957,N_23984);
xnor UO_1341 (O_1341,N_22514,N_24607);
nor UO_1342 (O_1342,N_24683,N_24625);
and UO_1343 (O_1343,N_23140,N_23735);
nand UO_1344 (O_1344,N_22538,N_23627);
xor UO_1345 (O_1345,N_22798,N_24890);
and UO_1346 (O_1346,N_23703,N_24949);
or UO_1347 (O_1347,N_23082,N_23002);
nand UO_1348 (O_1348,N_22518,N_22683);
nor UO_1349 (O_1349,N_24014,N_24552);
and UO_1350 (O_1350,N_23896,N_24854);
nand UO_1351 (O_1351,N_22795,N_24713);
nor UO_1352 (O_1352,N_23854,N_23518);
xor UO_1353 (O_1353,N_24989,N_22627);
and UO_1354 (O_1354,N_22569,N_23482);
nand UO_1355 (O_1355,N_23942,N_22540);
xnor UO_1356 (O_1356,N_23944,N_24259);
nor UO_1357 (O_1357,N_23417,N_23500);
nor UO_1358 (O_1358,N_23311,N_24483);
nor UO_1359 (O_1359,N_23872,N_23876);
nand UO_1360 (O_1360,N_24042,N_22582);
and UO_1361 (O_1361,N_23336,N_24979);
nor UO_1362 (O_1362,N_24159,N_23071);
and UO_1363 (O_1363,N_24595,N_24225);
xnor UO_1364 (O_1364,N_22569,N_23903);
or UO_1365 (O_1365,N_22574,N_23867);
or UO_1366 (O_1366,N_23812,N_24031);
and UO_1367 (O_1367,N_22843,N_23165);
nand UO_1368 (O_1368,N_22967,N_24180);
and UO_1369 (O_1369,N_22905,N_24566);
xnor UO_1370 (O_1370,N_24293,N_23893);
nand UO_1371 (O_1371,N_22914,N_23763);
or UO_1372 (O_1372,N_24824,N_22553);
nor UO_1373 (O_1373,N_22740,N_24462);
nor UO_1374 (O_1374,N_23003,N_22768);
nand UO_1375 (O_1375,N_22552,N_22572);
and UO_1376 (O_1376,N_23408,N_23139);
and UO_1377 (O_1377,N_24636,N_24570);
nand UO_1378 (O_1378,N_24369,N_24810);
nor UO_1379 (O_1379,N_24037,N_24972);
nor UO_1380 (O_1380,N_23823,N_24480);
and UO_1381 (O_1381,N_24280,N_22848);
and UO_1382 (O_1382,N_22988,N_24231);
and UO_1383 (O_1383,N_23717,N_24088);
or UO_1384 (O_1384,N_23078,N_23576);
nor UO_1385 (O_1385,N_24774,N_24080);
xor UO_1386 (O_1386,N_23345,N_23600);
xnor UO_1387 (O_1387,N_24635,N_22954);
nor UO_1388 (O_1388,N_23874,N_22517);
nor UO_1389 (O_1389,N_23175,N_24650);
nand UO_1390 (O_1390,N_23500,N_23445);
xnor UO_1391 (O_1391,N_23714,N_22657);
or UO_1392 (O_1392,N_24199,N_24888);
nor UO_1393 (O_1393,N_24892,N_23246);
xor UO_1394 (O_1394,N_24751,N_24065);
xnor UO_1395 (O_1395,N_22514,N_22693);
nand UO_1396 (O_1396,N_23239,N_22874);
xnor UO_1397 (O_1397,N_24314,N_23763);
nand UO_1398 (O_1398,N_22716,N_24153);
and UO_1399 (O_1399,N_24266,N_22896);
nand UO_1400 (O_1400,N_24515,N_24898);
or UO_1401 (O_1401,N_22971,N_24796);
or UO_1402 (O_1402,N_23761,N_24978);
nor UO_1403 (O_1403,N_23310,N_24052);
xor UO_1404 (O_1404,N_23949,N_23254);
xor UO_1405 (O_1405,N_23377,N_24781);
and UO_1406 (O_1406,N_23505,N_24183);
xor UO_1407 (O_1407,N_24531,N_23678);
xnor UO_1408 (O_1408,N_23748,N_22697);
and UO_1409 (O_1409,N_24295,N_23493);
xor UO_1410 (O_1410,N_23452,N_24479);
nand UO_1411 (O_1411,N_22583,N_22919);
nor UO_1412 (O_1412,N_24370,N_22569);
and UO_1413 (O_1413,N_22597,N_22964);
nand UO_1414 (O_1414,N_24188,N_23601);
nor UO_1415 (O_1415,N_22717,N_24418);
nor UO_1416 (O_1416,N_24393,N_22827);
xnor UO_1417 (O_1417,N_24520,N_23753);
nor UO_1418 (O_1418,N_22657,N_23419);
and UO_1419 (O_1419,N_23681,N_22884);
and UO_1420 (O_1420,N_24606,N_22506);
xor UO_1421 (O_1421,N_24983,N_24741);
xor UO_1422 (O_1422,N_24934,N_24664);
and UO_1423 (O_1423,N_23726,N_23498);
xor UO_1424 (O_1424,N_22586,N_23283);
nand UO_1425 (O_1425,N_24736,N_22592);
xnor UO_1426 (O_1426,N_23065,N_23858);
xor UO_1427 (O_1427,N_22694,N_24410);
and UO_1428 (O_1428,N_24175,N_24830);
or UO_1429 (O_1429,N_22903,N_23925);
or UO_1430 (O_1430,N_23953,N_24495);
xnor UO_1431 (O_1431,N_23360,N_23295);
or UO_1432 (O_1432,N_22737,N_23551);
nand UO_1433 (O_1433,N_23404,N_24770);
xor UO_1434 (O_1434,N_23993,N_24302);
xor UO_1435 (O_1435,N_24444,N_23838);
xnor UO_1436 (O_1436,N_24344,N_24816);
nor UO_1437 (O_1437,N_22927,N_23880);
or UO_1438 (O_1438,N_24204,N_23639);
nand UO_1439 (O_1439,N_24357,N_23733);
nor UO_1440 (O_1440,N_24410,N_24133);
and UO_1441 (O_1441,N_23298,N_23128);
nor UO_1442 (O_1442,N_24602,N_23489);
nor UO_1443 (O_1443,N_24544,N_24976);
nor UO_1444 (O_1444,N_22501,N_24996);
nand UO_1445 (O_1445,N_24091,N_22624);
nor UO_1446 (O_1446,N_22615,N_23666);
nand UO_1447 (O_1447,N_23817,N_23876);
and UO_1448 (O_1448,N_23460,N_23376);
and UO_1449 (O_1449,N_22631,N_23593);
and UO_1450 (O_1450,N_23233,N_24652);
xor UO_1451 (O_1451,N_23543,N_23499);
xnor UO_1452 (O_1452,N_23520,N_22925);
xnor UO_1453 (O_1453,N_24551,N_24844);
nand UO_1454 (O_1454,N_23387,N_24367);
nand UO_1455 (O_1455,N_24068,N_22822);
or UO_1456 (O_1456,N_24964,N_23070);
and UO_1457 (O_1457,N_23392,N_24077);
nand UO_1458 (O_1458,N_24140,N_24975);
or UO_1459 (O_1459,N_24983,N_22588);
and UO_1460 (O_1460,N_23606,N_23610);
or UO_1461 (O_1461,N_22551,N_24620);
or UO_1462 (O_1462,N_23551,N_24737);
and UO_1463 (O_1463,N_23075,N_23817);
nor UO_1464 (O_1464,N_23920,N_24702);
xor UO_1465 (O_1465,N_24637,N_22914);
and UO_1466 (O_1466,N_23760,N_22968);
and UO_1467 (O_1467,N_23160,N_22739);
or UO_1468 (O_1468,N_23889,N_24837);
or UO_1469 (O_1469,N_24144,N_24840);
or UO_1470 (O_1470,N_23257,N_23071);
nor UO_1471 (O_1471,N_23454,N_23268);
xnor UO_1472 (O_1472,N_22688,N_24786);
and UO_1473 (O_1473,N_22667,N_22740);
nand UO_1474 (O_1474,N_23048,N_23922);
or UO_1475 (O_1475,N_23081,N_24277);
nor UO_1476 (O_1476,N_24435,N_23376);
xor UO_1477 (O_1477,N_24844,N_24276);
and UO_1478 (O_1478,N_24146,N_23828);
nor UO_1479 (O_1479,N_24438,N_24144);
and UO_1480 (O_1480,N_24007,N_23137);
xor UO_1481 (O_1481,N_23511,N_23523);
or UO_1482 (O_1482,N_23943,N_23296);
nand UO_1483 (O_1483,N_23413,N_24461);
nand UO_1484 (O_1484,N_23431,N_23233);
nand UO_1485 (O_1485,N_22789,N_24773);
and UO_1486 (O_1486,N_24824,N_24363);
nor UO_1487 (O_1487,N_23827,N_24827);
nand UO_1488 (O_1488,N_24394,N_23674);
nand UO_1489 (O_1489,N_24767,N_23031);
nand UO_1490 (O_1490,N_24581,N_23078);
and UO_1491 (O_1491,N_22612,N_23033);
nand UO_1492 (O_1492,N_23346,N_22517);
or UO_1493 (O_1493,N_23521,N_23231);
nor UO_1494 (O_1494,N_24957,N_22965);
nand UO_1495 (O_1495,N_23552,N_23474);
nor UO_1496 (O_1496,N_22640,N_22680);
nand UO_1497 (O_1497,N_22964,N_23216);
xor UO_1498 (O_1498,N_24935,N_23304);
nand UO_1499 (O_1499,N_24232,N_24154);
nand UO_1500 (O_1500,N_24331,N_24372);
or UO_1501 (O_1501,N_23729,N_24555);
nand UO_1502 (O_1502,N_22794,N_22616);
xnor UO_1503 (O_1503,N_23276,N_24527);
xnor UO_1504 (O_1504,N_24387,N_23489);
or UO_1505 (O_1505,N_23988,N_24558);
and UO_1506 (O_1506,N_23302,N_23493);
or UO_1507 (O_1507,N_23524,N_23539);
nand UO_1508 (O_1508,N_23322,N_24130);
nand UO_1509 (O_1509,N_23795,N_22604);
xnor UO_1510 (O_1510,N_23151,N_23652);
nand UO_1511 (O_1511,N_23115,N_23129);
xor UO_1512 (O_1512,N_23749,N_24705);
nand UO_1513 (O_1513,N_22748,N_23600);
nor UO_1514 (O_1514,N_24563,N_24248);
xor UO_1515 (O_1515,N_22986,N_23605);
or UO_1516 (O_1516,N_24120,N_24579);
and UO_1517 (O_1517,N_23170,N_24098);
xnor UO_1518 (O_1518,N_24409,N_24819);
nor UO_1519 (O_1519,N_24551,N_24889);
xor UO_1520 (O_1520,N_22992,N_24451);
nor UO_1521 (O_1521,N_22786,N_23324);
nand UO_1522 (O_1522,N_24337,N_24394);
or UO_1523 (O_1523,N_24887,N_23284);
nand UO_1524 (O_1524,N_22695,N_23271);
nand UO_1525 (O_1525,N_24824,N_23110);
or UO_1526 (O_1526,N_23612,N_22971);
nand UO_1527 (O_1527,N_22716,N_24752);
or UO_1528 (O_1528,N_23269,N_23643);
xor UO_1529 (O_1529,N_23480,N_24900);
xnor UO_1530 (O_1530,N_23555,N_24389);
and UO_1531 (O_1531,N_24344,N_23192);
xor UO_1532 (O_1532,N_22805,N_24842);
and UO_1533 (O_1533,N_24533,N_22845);
and UO_1534 (O_1534,N_23897,N_24250);
nor UO_1535 (O_1535,N_22657,N_23741);
or UO_1536 (O_1536,N_23542,N_24998);
nor UO_1537 (O_1537,N_24474,N_24120);
nand UO_1538 (O_1538,N_23031,N_24802);
or UO_1539 (O_1539,N_23187,N_23580);
and UO_1540 (O_1540,N_24007,N_23094);
nor UO_1541 (O_1541,N_23660,N_22994);
xnor UO_1542 (O_1542,N_22636,N_24934);
or UO_1543 (O_1543,N_24198,N_23454);
or UO_1544 (O_1544,N_23613,N_23507);
xor UO_1545 (O_1545,N_24410,N_23488);
or UO_1546 (O_1546,N_22919,N_24510);
nor UO_1547 (O_1547,N_23022,N_23985);
nand UO_1548 (O_1548,N_24290,N_23762);
xnor UO_1549 (O_1549,N_22831,N_24325);
nor UO_1550 (O_1550,N_22794,N_24865);
nand UO_1551 (O_1551,N_22698,N_23530);
or UO_1552 (O_1552,N_22792,N_24463);
nand UO_1553 (O_1553,N_23408,N_22997);
nor UO_1554 (O_1554,N_24807,N_24170);
or UO_1555 (O_1555,N_24088,N_23151);
or UO_1556 (O_1556,N_24699,N_23071);
nand UO_1557 (O_1557,N_24581,N_23117);
and UO_1558 (O_1558,N_22809,N_23631);
and UO_1559 (O_1559,N_22524,N_24908);
nand UO_1560 (O_1560,N_23654,N_23819);
xor UO_1561 (O_1561,N_24781,N_23734);
or UO_1562 (O_1562,N_24951,N_24734);
xnor UO_1563 (O_1563,N_22840,N_23306);
nor UO_1564 (O_1564,N_22887,N_24118);
nand UO_1565 (O_1565,N_22639,N_23203);
or UO_1566 (O_1566,N_22796,N_23043);
or UO_1567 (O_1567,N_23326,N_23770);
or UO_1568 (O_1568,N_23606,N_24050);
or UO_1569 (O_1569,N_22528,N_23516);
and UO_1570 (O_1570,N_24054,N_23514);
nor UO_1571 (O_1571,N_23882,N_24586);
nor UO_1572 (O_1572,N_23404,N_24891);
or UO_1573 (O_1573,N_22941,N_24974);
nand UO_1574 (O_1574,N_23798,N_23327);
nor UO_1575 (O_1575,N_22550,N_23904);
and UO_1576 (O_1576,N_24835,N_24860);
nor UO_1577 (O_1577,N_24684,N_24079);
and UO_1578 (O_1578,N_24470,N_24399);
or UO_1579 (O_1579,N_22506,N_24192);
xnor UO_1580 (O_1580,N_23511,N_24161);
nor UO_1581 (O_1581,N_24457,N_24355);
nand UO_1582 (O_1582,N_23917,N_24782);
and UO_1583 (O_1583,N_23547,N_23740);
xnor UO_1584 (O_1584,N_23570,N_22859);
xor UO_1585 (O_1585,N_23432,N_24321);
nor UO_1586 (O_1586,N_24062,N_22963);
and UO_1587 (O_1587,N_24042,N_22513);
xnor UO_1588 (O_1588,N_24229,N_24183);
and UO_1589 (O_1589,N_22989,N_22933);
nand UO_1590 (O_1590,N_23853,N_24851);
xnor UO_1591 (O_1591,N_23105,N_24945);
nand UO_1592 (O_1592,N_24370,N_22896);
xnor UO_1593 (O_1593,N_23629,N_22804);
nand UO_1594 (O_1594,N_24876,N_24975);
nand UO_1595 (O_1595,N_22927,N_24195);
and UO_1596 (O_1596,N_22766,N_24014);
nor UO_1597 (O_1597,N_24822,N_24562);
nor UO_1598 (O_1598,N_23428,N_23132);
xor UO_1599 (O_1599,N_23808,N_24700);
nor UO_1600 (O_1600,N_24496,N_24128);
or UO_1601 (O_1601,N_23275,N_24137);
xor UO_1602 (O_1602,N_24642,N_24853);
xor UO_1603 (O_1603,N_24184,N_22973);
or UO_1604 (O_1604,N_24054,N_22601);
and UO_1605 (O_1605,N_23227,N_23943);
xor UO_1606 (O_1606,N_23035,N_23213);
nand UO_1607 (O_1607,N_23736,N_24897);
and UO_1608 (O_1608,N_24894,N_24146);
or UO_1609 (O_1609,N_24933,N_22626);
nor UO_1610 (O_1610,N_23166,N_23014);
or UO_1611 (O_1611,N_23969,N_23485);
and UO_1612 (O_1612,N_24525,N_23091);
nand UO_1613 (O_1613,N_23288,N_23107);
nand UO_1614 (O_1614,N_22608,N_24896);
nand UO_1615 (O_1615,N_24659,N_22870);
nor UO_1616 (O_1616,N_24935,N_23265);
and UO_1617 (O_1617,N_24467,N_23273);
or UO_1618 (O_1618,N_23292,N_23119);
nand UO_1619 (O_1619,N_24545,N_22967);
xnor UO_1620 (O_1620,N_24766,N_24120);
and UO_1621 (O_1621,N_22901,N_24255);
or UO_1622 (O_1622,N_23268,N_24762);
xor UO_1623 (O_1623,N_24751,N_23817);
nor UO_1624 (O_1624,N_24922,N_23856);
nand UO_1625 (O_1625,N_22955,N_24220);
nor UO_1626 (O_1626,N_22686,N_22628);
nand UO_1627 (O_1627,N_24980,N_22887);
xor UO_1628 (O_1628,N_24725,N_23251);
nand UO_1629 (O_1629,N_24603,N_24542);
and UO_1630 (O_1630,N_24512,N_24926);
nor UO_1631 (O_1631,N_22538,N_24476);
or UO_1632 (O_1632,N_24164,N_22832);
nor UO_1633 (O_1633,N_24473,N_24898);
nor UO_1634 (O_1634,N_23443,N_23133);
or UO_1635 (O_1635,N_24765,N_24592);
xnor UO_1636 (O_1636,N_22723,N_23514);
and UO_1637 (O_1637,N_22592,N_23080);
nand UO_1638 (O_1638,N_24924,N_24675);
nand UO_1639 (O_1639,N_24059,N_24408);
nand UO_1640 (O_1640,N_23594,N_23432);
nand UO_1641 (O_1641,N_24962,N_23750);
nor UO_1642 (O_1642,N_23458,N_23283);
xnor UO_1643 (O_1643,N_22763,N_23235);
nand UO_1644 (O_1644,N_23503,N_23241);
and UO_1645 (O_1645,N_24196,N_23830);
nor UO_1646 (O_1646,N_23958,N_23687);
nor UO_1647 (O_1647,N_24610,N_22693);
nand UO_1648 (O_1648,N_22548,N_24516);
nor UO_1649 (O_1649,N_23869,N_22762);
or UO_1650 (O_1650,N_23924,N_23622);
nor UO_1651 (O_1651,N_23043,N_23580);
and UO_1652 (O_1652,N_23579,N_24769);
or UO_1653 (O_1653,N_24102,N_24113);
nor UO_1654 (O_1654,N_23965,N_23665);
xor UO_1655 (O_1655,N_22505,N_23518);
and UO_1656 (O_1656,N_24708,N_22926);
xnor UO_1657 (O_1657,N_22529,N_23523);
xor UO_1658 (O_1658,N_23492,N_23025);
nor UO_1659 (O_1659,N_24721,N_24559);
and UO_1660 (O_1660,N_23355,N_23353);
xor UO_1661 (O_1661,N_24592,N_24285);
xor UO_1662 (O_1662,N_24560,N_23218);
and UO_1663 (O_1663,N_22535,N_23936);
nor UO_1664 (O_1664,N_24825,N_22802);
xor UO_1665 (O_1665,N_23120,N_23044);
or UO_1666 (O_1666,N_23624,N_23024);
nor UO_1667 (O_1667,N_23891,N_23340);
nand UO_1668 (O_1668,N_23985,N_23905);
or UO_1669 (O_1669,N_24741,N_24237);
and UO_1670 (O_1670,N_24934,N_24287);
nand UO_1671 (O_1671,N_22688,N_23038);
nand UO_1672 (O_1672,N_23135,N_23261);
or UO_1673 (O_1673,N_22937,N_24871);
nor UO_1674 (O_1674,N_24620,N_22911);
xor UO_1675 (O_1675,N_22586,N_24546);
xnor UO_1676 (O_1676,N_23637,N_23693);
and UO_1677 (O_1677,N_23736,N_24586);
and UO_1678 (O_1678,N_23583,N_22831);
nand UO_1679 (O_1679,N_23238,N_24078);
and UO_1680 (O_1680,N_22973,N_23857);
and UO_1681 (O_1681,N_23753,N_23183);
xnor UO_1682 (O_1682,N_23344,N_22813);
and UO_1683 (O_1683,N_23730,N_23554);
and UO_1684 (O_1684,N_24465,N_22795);
and UO_1685 (O_1685,N_22789,N_22608);
xor UO_1686 (O_1686,N_24680,N_23702);
nand UO_1687 (O_1687,N_23109,N_24155);
xor UO_1688 (O_1688,N_24605,N_22623);
and UO_1689 (O_1689,N_23935,N_23262);
and UO_1690 (O_1690,N_24338,N_23034);
nand UO_1691 (O_1691,N_23140,N_22737);
and UO_1692 (O_1692,N_24164,N_22754);
nand UO_1693 (O_1693,N_23593,N_23991);
nand UO_1694 (O_1694,N_23810,N_22727);
nand UO_1695 (O_1695,N_23705,N_24168);
xor UO_1696 (O_1696,N_23171,N_23741);
nand UO_1697 (O_1697,N_22934,N_23665);
nand UO_1698 (O_1698,N_22869,N_23378);
nor UO_1699 (O_1699,N_23425,N_22547);
nand UO_1700 (O_1700,N_24195,N_23451);
nand UO_1701 (O_1701,N_24696,N_23400);
or UO_1702 (O_1702,N_23327,N_24914);
nor UO_1703 (O_1703,N_24860,N_23909);
nand UO_1704 (O_1704,N_24409,N_24904);
xnor UO_1705 (O_1705,N_23769,N_22960);
and UO_1706 (O_1706,N_24395,N_24901);
xnor UO_1707 (O_1707,N_22899,N_23618);
and UO_1708 (O_1708,N_24147,N_23678);
and UO_1709 (O_1709,N_23638,N_24576);
nand UO_1710 (O_1710,N_24430,N_23631);
nand UO_1711 (O_1711,N_22631,N_22721);
and UO_1712 (O_1712,N_24022,N_24502);
nand UO_1713 (O_1713,N_22752,N_24478);
or UO_1714 (O_1714,N_22882,N_24991);
xnor UO_1715 (O_1715,N_23217,N_22672);
nor UO_1716 (O_1716,N_24209,N_22587);
nor UO_1717 (O_1717,N_23697,N_23962);
xor UO_1718 (O_1718,N_23764,N_24742);
nor UO_1719 (O_1719,N_23403,N_24798);
xnor UO_1720 (O_1720,N_23522,N_23688);
nand UO_1721 (O_1721,N_24953,N_23247);
nand UO_1722 (O_1722,N_24349,N_22742);
nand UO_1723 (O_1723,N_22820,N_24093);
and UO_1724 (O_1724,N_22652,N_24409);
nor UO_1725 (O_1725,N_22904,N_23508);
nand UO_1726 (O_1726,N_24118,N_23178);
nand UO_1727 (O_1727,N_23758,N_22543);
xnor UO_1728 (O_1728,N_22608,N_23700);
or UO_1729 (O_1729,N_23633,N_23705);
or UO_1730 (O_1730,N_23656,N_24513);
and UO_1731 (O_1731,N_24974,N_24591);
nor UO_1732 (O_1732,N_24787,N_22686);
and UO_1733 (O_1733,N_23348,N_23848);
nand UO_1734 (O_1734,N_24319,N_24823);
nand UO_1735 (O_1735,N_23885,N_24618);
and UO_1736 (O_1736,N_23422,N_22829);
or UO_1737 (O_1737,N_22752,N_23664);
xnor UO_1738 (O_1738,N_24002,N_22527);
xor UO_1739 (O_1739,N_22960,N_24689);
nand UO_1740 (O_1740,N_23587,N_23958);
nand UO_1741 (O_1741,N_24914,N_23995);
nor UO_1742 (O_1742,N_22964,N_22615);
and UO_1743 (O_1743,N_22668,N_22905);
nor UO_1744 (O_1744,N_23851,N_22937);
nor UO_1745 (O_1745,N_22966,N_22823);
nor UO_1746 (O_1746,N_22891,N_24855);
nor UO_1747 (O_1747,N_22942,N_24273);
nor UO_1748 (O_1748,N_23165,N_23967);
nor UO_1749 (O_1749,N_23816,N_22778);
xor UO_1750 (O_1750,N_24700,N_23845);
nor UO_1751 (O_1751,N_22783,N_24894);
or UO_1752 (O_1752,N_23002,N_23168);
and UO_1753 (O_1753,N_23892,N_22703);
xnor UO_1754 (O_1754,N_23030,N_24345);
and UO_1755 (O_1755,N_23970,N_22789);
nor UO_1756 (O_1756,N_24327,N_23608);
and UO_1757 (O_1757,N_23397,N_23526);
or UO_1758 (O_1758,N_23025,N_24173);
and UO_1759 (O_1759,N_23397,N_23351);
or UO_1760 (O_1760,N_23094,N_22868);
nor UO_1761 (O_1761,N_22527,N_23625);
or UO_1762 (O_1762,N_24581,N_23420);
or UO_1763 (O_1763,N_24199,N_22850);
nand UO_1764 (O_1764,N_24979,N_22698);
and UO_1765 (O_1765,N_24168,N_23793);
nand UO_1766 (O_1766,N_24694,N_24966);
and UO_1767 (O_1767,N_24932,N_24501);
nor UO_1768 (O_1768,N_23006,N_24979);
xor UO_1769 (O_1769,N_24480,N_22828);
nor UO_1770 (O_1770,N_24021,N_23220);
or UO_1771 (O_1771,N_23848,N_23322);
nor UO_1772 (O_1772,N_24545,N_23354);
nand UO_1773 (O_1773,N_22524,N_24379);
or UO_1774 (O_1774,N_22526,N_22550);
or UO_1775 (O_1775,N_23170,N_24703);
nor UO_1776 (O_1776,N_24616,N_23460);
nor UO_1777 (O_1777,N_24933,N_23540);
xor UO_1778 (O_1778,N_23663,N_24352);
or UO_1779 (O_1779,N_23477,N_22742);
and UO_1780 (O_1780,N_23361,N_23695);
nand UO_1781 (O_1781,N_24518,N_22667);
and UO_1782 (O_1782,N_24305,N_22933);
and UO_1783 (O_1783,N_23151,N_24991);
xor UO_1784 (O_1784,N_24229,N_24544);
nor UO_1785 (O_1785,N_23621,N_23674);
or UO_1786 (O_1786,N_22864,N_24323);
or UO_1787 (O_1787,N_23124,N_24399);
or UO_1788 (O_1788,N_24286,N_23179);
nand UO_1789 (O_1789,N_23051,N_24921);
nor UO_1790 (O_1790,N_22985,N_24705);
nand UO_1791 (O_1791,N_23477,N_23919);
nand UO_1792 (O_1792,N_23594,N_23210);
or UO_1793 (O_1793,N_24705,N_24339);
nor UO_1794 (O_1794,N_24956,N_24990);
xor UO_1795 (O_1795,N_24560,N_23143);
nor UO_1796 (O_1796,N_23059,N_24098);
xor UO_1797 (O_1797,N_24247,N_23872);
nor UO_1798 (O_1798,N_24969,N_24787);
and UO_1799 (O_1799,N_24862,N_22750);
nand UO_1800 (O_1800,N_24402,N_22844);
xnor UO_1801 (O_1801,N_24004,N_23626);
nand UO_1802 (O_1802,N_23899,N_23452);
and UO_1803 (O_1803,N_24150,N_24888);
and UO_1804 (O_1804,N_23593,N_24415);
nor UO_1805 (O_1805,N_22800,N_24768);
or UO_1806 (O_1806,N_23185,N_23890);
xnor UO_1807 (O_1807,N_24724,N_23226);
nor UO_1808 (O_1808,N_24652,N_23089);
nand UO_1809 (O_1809,N_22903,N_23476);
xnor UO_1810 (O_1810,N_24429,N_22699);
and UO_1811 (O_1811,N_23686,N_23234);
nand UO_1812 (O_1812,N_23797,N_23149);
xor UO_1813 (O_1813,N_24924,N_23156);
xor UO_1814 (O_1814,N_23785,N_22691);
and UO_1815 (O_1815,N_23342,N_24974);
and UO_1816 (O_1816,N_23333,N_22554);
or UO_1817 (O_1817,N_23215,N_23488);
or UO_1818 (O_1818,N_22743,N_23278);
nor UO_1819 (O_1819,N_23934,N_24400);
xor UO_1820 (O_1820,N_24194,N_24580);
xnor UO_1821 (O_1821,N_24774,N_22799);
xor UO_1822 (O_1822,N_24966,N_23413);
and UO_1823 (O_1823,N_22593,N_23018);
nor UO_1824 (O_1824,N_22823,N_24784);
nor UO_1825 (O_1825,N_24217,N_24107);
and UO_1826 (O_1826,N_22847,N_23861);
xnor UO_1827 (O_1827,N_24575,N_22808);
xor UO_1828 (O_1828,N_24458,N_23501);
nand UO_1829 (O_1829,N_24263,N_24078);
nor UO_1830 (O_1830,N_23495,N_24842);
nor UO_1831 (O_1831,N_24378,N_23436);
or UO_1832 (O_1832,N_23079,N_23850);
or UO_1833 (O_1833,N_24151,N_24044);
and UO_1834 (O_1834,N_23491,N_23816);
and UO_1835 (O_1835,N_23322,N_24177);
nor UO_1836 (O_1836,N_24734,N_23372);
xnor UO_1837 (O_1837,N_24892,N_23533);
or UO_1838 (O_1838,N_22659,N_24261);
and UO_1839 (O_1839,N_22890,N_24922);
nand UO_1840 (O_1840,N_24135,N_23241);
nor UO_1841 (O_1841,N_24400,N_23990);
and UO_1842 (O_1842,N_24404,N_24965);
xnor UO_1843 (O_1843,N_22928,N_23288);
nand UO_1844 (O_1844,N_23065,N_24094);
or UO_1845 (O_1845,N_24213,N_24138);
nor UO_1846 (O_1846,N_24813,N_24028);
or UO_1847 (O_1847,N_23874,N_22580);
and UO_1848 (O_1848,N_23485,N_24743);
nand UO_1849 (O_1849,N_22592,N_24949);
or UO_1850 (O_1850,N_24948,N_22512);
nand UO_1851 (O_1851,N_24575,N_24260);
xor UO_1852 (O_1852,N_22619,N_23121);
nand UO_1853 (O_1853,N_22911,N_22807);
nor UO_1854 (O_1854,N_23704,N_23684);
nand UO_1855 (O_1855,N_24002,N_23097);
or UO_1856 (O_1856,N_24697,N_23492);
or UO_1857 (O_1857,N_22646,N_22501);
or UO_1858 (O_1858,N_23730,N_23505);
nor UO_1859 (O_1859,N_24092,N_23899);
or UO_1860 (O_1860,N_24830,N_23407);
and UO_1861 (O_1861,N_24174,N_24604);
nand UO_1862 (O_1862,N_23876,N_24983);
nand UO_1863 (O_1863,N_23985,N_23665);
nor UO_1864 (O_1864,N_24759,N_23072);
or UO_1865 (O_1865,N_22773,N_23152);
or UO_1866 (O_1866,N_24841,N_23989);
nand UO_1867 (O_1867,N_24591,N_22572);
nand UO_1868 (O_1868,N_23857,N_23778);
nor UO_1869 (O_1869,N_24115,N_23476);
and UO_1870 (O_1870,N_22910,N_23149);
nor UO_1871 (O_1871,N_22870,N_24854);
nand UO_1872 (O_1872,N_24237,N_24427);
xor UO_1873 (O_1873,N_23134,N_24684);
and UO_1874 (O_1874,N_24960,N_24839);
or UO_1875 (O_1875,N_23507,N_24883);
nand UO_1876 (O_1876,N_24253,N_23905);
nor UO_1877 (O_1877,N_23200,N_22749);
or UO_1878 (O_1878,N_24773,N_23938);
nand UO_1879 (O_1879,N_23285,N_23744);
nand UO_1880 (O_1880,N_24726,N_22790);
nor UO_1881 (O_1881,N_23008,N_24729);
nand UO_1882 (O_1882,N_22618,N_24539);
or UO_1883 (O_1883,N_22706,N_24470);
or UO_1884 (O_1884,N_23573,N_23538);
and UO_1885 (O_1885,N_24285,N_23530);
and UO_1886 (O_1886,N_24491,N_23240);
and UO_1887 (O_1887,N_24784,N_23150);
nor UO_1888 (O_1888,N_24264,N_22918);
nand UO_1889 (O_1889,N_22877,N_24643);
or UO_1890 (O_1890,N_22666,N_23894);
nor UO_1891 (O_1891,N_24893,N_22744);
xor UO_1892 (O_1892,N_22857,N_23367);
and UO_1893 (O_1893,N_23242,N_23850);
nor UO_1894 (O_1894,N_23052,N_23819);
xnor UO_1895 (O_1895,N_24831,N_23605);
and UO_1896 (O_1896,N_24599,N_24058);
or UO_1897 (O_1897,N_24961,N_24919);
xor UO_1898 (O_1898,N_23777,N_23586);
xnor UO_1899 (O_1899,N_24870,N_23050);
and UO_1900 (O_1900,N_24571,N_24303);
nand UO_1901 (O_1901,N_23333,N_24581);
xor UO_1902 (O_1902,N_23296,N_23956);
or UO_1903 (O_1903,N_22951,N_24192);
nand UO_1904 (O_1904,N_23843,N_23531);
nand UO_1905 (O_1905,N_23927,N_23018);
nand UO_1906 (O_1906,N_22564,N_23906);
and UO_1907 (O_1907,N_22645,N_24951);
nand UO_1908 (O_1908,N_23900,N_24547);
xnor UO_1909 (O_1909,N_22703,N_23561);
or UO_1910 (O_1910,N_23644,N_22657);
or UO_1911 (O_1911,N_24158,N_24329);
and UO_1912 (O_1912,N_23491,N_23382);
or UO_1913 (O_1913,N_22961,N_24352);
or UO_1914 (O_1914,N_22683,N_22772);
xnor UO_1915 (O_1915,N_23546,N_23642);
or UO_1916 (O_1916,N_23814,N_24187);
nor UO_1917 (O_1917,N_23239,N_23006);
nand UO_1918 (O_1918,N_22739,N_23428);
nor UO_1919 (O_1919,N_22849,N_24091);
nor UO_1920 (O_1920,N_24577,N_24429);
nand UO_1921 (O_1921,N_23936,N_24680);
or UO_1922 (O_1922,N_24393,N_22688);
and UO_1923 (O_1923,N_24048,N_23024);
or UO_1924 (O_1924,N_23794,N_24701);
nand UO_1925 (O_1925,N_24427,N_22562);
nand UO_1926 (O_1926,N_23116,N_24394);
nor UO_1927 (O_1927,N_24032,N_23059);
or UO_1928 (O_1928,N_22649,N_23143);
and UO_1929 (O_1929,N_23091,N_23632);
or UO_1930 (O_1930,N_23521,N_23417);
or UO_1931 (O_1931,N_22616,N_22748);
xor UO_1932 (O_1932,N_23704,N_24820);
xnor UO_1933 (O_1933,N_24381,N_23257);
and UO_1934 (O_1934,N_24581,N_24878);
xnor UO_1935 (O_1935,N_24136,N_23559);
or UO_1936 (O_1936,N_23371,N_22887);
xnor UO_1937 (O_1937,N_24682,N_23774);
nor UO_1938 (O_1938,N_24936,N_23996);
nand UO_1939 (O_1939,N_24174,N_23545);
and UO_1940 (O_1940,N_24600,N_23439);
nor UO_1941 (O_1941,N_24894,N_23491);
nor UO_1942 (O_1942,N_23691,N_24078);
and UO_1943 (O_1943,N_24035,N_24405);
xor UO_1944 (O_1944,N_23000,N_24839);
and UO_1945 (O_1945,N_24725,N_24275);
nor UO_1946 (O_1946,N_22566,N_22536);
and UO_1947 (O_1947,N_23195,N_24067);
nand UO_1948 (O_1948,N_23545,N_22996);
nor UO_1949 (O_1949,N_23016,N_22727);
nand UO_1950 (O_1950,N_24551,N_23631);
xor UO_1951 (O_1951,N_23089,N_23845);
nor UO_1952 (O_1952,N_24754,N_23024);
nor UO_1953 (O_1953,N_22676,N_23509);
nand UO_1954 (O_1954,N_23889,N_23176);
or UO_1955 (O_1955,N_22552,N_23508);
or UO_1956 (O_1956,N_23318,N_24553);
and UO_1957 (O_1957,N_23282,N_22748);
nor UO_1958 (O_1958,N_22656,N_24853);
nand UO_1959 (O_1959,N_23266,N_23212);
xor UO_1960 (O_1960,N_22653,N_24246);
and UO_1961 (O_1961,N_24947,N_23498);
and UO_1962 (O_1962,N_24218,N_24071);
nand UO_1963 (O_1963,N_22916,N_23770);
or UO_1964 (O_1964,N_22670,N_23137);
and UO_1965 (O_1965,N_24013,N_23328);
nor UO_1966 (O_1966,N_22725,N_23092);
or UO_1967 (O_1967,N_24606,N_22865);
and UO_1968 (O_1968,N_24830,N_23365);
nor UO_1969 (O_1969,N_23152,N_23630);
xnor UO_1970 (O_1970,N_23596,N_23458);
and UO_1971 (O_1971,N_24072,N_23036);
nor UO_1972 (O_1972,N_24672,N_24911);
xnor UO_1973 (O_1973,N_23695,N_24175);
or UO_1974 (O_1974,N_24838,N_24827);
and UO_1975 (O_1975,N_23543,N_23934);
xor UO_1976 (O_1976,N_24467,N_23562);
nand UO_1977 (O_1977,N_24720,N_24574);
nand UO_1978 (O_1978,N_23126,N_24413);
xor UO_1979 (O_1979,N_24517,N_23521);
nor UO_1980 (O_1980,N_23025,N_23945);
and UO_1981 (O_1981,N_24486,N_23352);
and UO_1982 (O_1982,N_23622,N_24825);
nand UO_1983 (O_1983,N_24408,N_24079);
nor UO_1984 (O_1984,N_23879,N_23705);
and UO_1985 (O_1985,N_24446,N_22807);
or UO_1986 (O_1986,N_23321,N_23448);
nor UO_1987 (O_1987,N_24609,N_24916);
or UO_1988 (O_1988,N_22751,N_24591);
and UO_1989 (O_1989,N_23849,N_24644);
nand UO_1990 (O_1990,N_23511,N_24649);
and UO_1991 (O_1991,N_24514,N_24869);
and UO_1992 (O_1992,N_22514,N_24647);
xnor UO_1993 (O_1993,N_24703,N_24067);
nand UO_1994 (O_1994,N_22599,N_24189);
nor UO_1995 (O_1995,N_24615,N_23917);
and UO_1996 (O_1996,N_24123,N_24415);
nand UO_1997 (O_1997,N_22772,N_22760);
xor UO_1998 (O_1998,N_24308,N_22656);
nor UO_1999 (O_1999,N_22961,N_22869);
nor UO_2000 (O_2000,N_24425,N_22543);
xnor UO_2001 (O_2001,N_22542,N_23892);
and UO_2002 (O_2002,N_24229,N_22774);
nand UO_2003 (O_2003,N_24332,N_23826);
xnor UO_2004 (O_2004,N_23761,N_23267);
xor UO_2005 (O_2005,N_22992,N_23547);
nor UO_2006 (O_2006,N_24657,N_23128);
nor UO_2007 (O_2007,N_22701,N_24248);
nand UO_2008 (O_2008,N_23360,N_22863);
nand UO_2009 (O_2009,N_23853,N_22571);
or UO_2010 (O_2010,N_24067,N_23077);
nor UO_2011 (O_2011,N_23107,N_23003);
nor UO_2012 (O_2012,N_23434,N_23036);
nand UO_2013 (O_2013,N_22644,N_22859);
nor UO_2014 (O_2014,N_23827,N_23899);
nand UO_2015 (O_2015,N_23829,N_24279);
or UO_2016 (O_2016,N_23755,N_23326);
or UO_2017 (O_2017,N_24665,N_24953);
and UO_2018 (O_2018,N_24055,N_23976);
xnor UO_2019 (O_2019,N_24077,N_23985);
and UO_2020 (O_2020,N_23050,N_24512);
or UO_2021 (O_2021,N_22973,N_23438);
xor UO_2022 (O_2022,N_23013,N_24907);
nand UO_2023 (O_2023,N_24879,N_24578);
nand UO_2024 (O_2024,N_24478,N_24115);
xor UO_2025 (O_2025,N_23081,N_23626);
nand UO_2026 (O_2026,N_23201,N_23778);
nand UO_2027 (O_2027,N_22913,N_24314);
and UO_2028 (O_2028,N_24491,N_23926);
nand UO_2029 (O_2029,N_24433,N_23211);
nor UO_2030 (O_2030,N_23985,N_22661);
xnor UO_2031 (O_2031,N_22753,N_24600);
nor UO_2032 (O_2032,N_22799,N_23347);
and UO_2033 (O_2033,N_23809,N_24314);
nand UO_2034 (O_2034,N_22742,N_22843);
nand UO_2035 (O_2035,N_23658,N_22662);
nand UO_2036 (O_2036,N_24851,N_24866);
nand UO_2037 (O_2037,N_24005,N_23150);
and UO_2038 (O_2038,N_24140,N_22622);
xor UO_2039 (O_2039,N_23373,N_23784);
or UO_2040 (O_2040,N_24017,N_22930);
nand UO_2041 (O_2041,N_23172,N_22664);
nor UO_2042 (O_2042,N_23902,N_24542);
nor UO_2043 (O_2043,N_23169,N_22624);
nand UO_2044 (O_2044,N_24016,N_22912);
and UO_2045 (O_2045,N_24683,N_24346);
nand UO_2046 (O_2046,N_24478,N_24729);
nand UO_2047 (O_2047,N_24183,N_24447);
xnor UO_2048 (O_2048,N_24511,N_22846);
or UO_2049 (O_2049,N_23894,N_23562);
and UO_2050 (O_2050,N_23712,N_22879);
xnor UO_2051 (O_2051,N_23596,N_23359);
and UO_2052 (O_2052,N_23522,N_23940);
and UO_2053 (O_2053,N_23473,N_23098);
or UO_2054 (O_2054,N_22535,N_23457);
nand UO_2055 (O_2055,N_22823,N_23685);
or UO_2056 (O_2056,N_23636,N_24678);
nand UO_2057 (O_2057,N_22871,N_24264);
xor UO_2058 (O_2058,N_22530,N_24705);
and UO_2059 (O_2059,N_24407,N_23986);
nor UO_2060 (O_2060,N_23278,N_24094);
or UO_2061 (O_2061,N_23906,N_23188);
nor UO_2062 (O_2062,N_23199,N_23676);
xor UO_2063 (O_2063,N_24086,N_22588);
nor UO_2064 (O_2064,N_24278,N_24683);
and UO_2065 (O_2065,N_22670,N_23989);
and UO_2066 (O_2066,N_24767,N_23993);
or UO_2067 (O_2067,N_22716,N_24232);
xor UO_2068 (O_2068,N_24315,N_22945);
or UO_2069 (O_2069,N_23943,N_24041);
xor UO_2070 (O_2070,N_24464,N_23032);
xnor UO_2071 (O_2071,N_24617,N_23862);
xnor UO_2072 (O_2072,N_22504,N_24056);
xnor UO_2073 (O_2073,N_24357,N_23200);
nor UO_2074 (O_2074,N_23320,N_24699);
nor UO_2075 (O_2075,N_24394,N_23379);
and UO_2076 (O_2076,N_23316,N_22858);
or UO_2077 (O_2077,N_24270,N_24579);
xnor UO_2078 (O_2078,N_23527,N_23436);
or UO_2079 (O_2079,N_24598,N_24334);
nor UO_2080 (O_2080,N_24170,N_24095);
and UO_2081 (O_2081,N_23754,N_24047);
or UO_2082 (O_2082,N_23323,N_24154);
xnor UO_2083 (O_2083,N_23835,N_22943);
and UO_2084 (O_2084,N_23100,N_24425);
and UO_2085 (O_2085,N_24071,N_23917);
nor UO_2086 (O_2086,N_24151,N_24695);
nor UO_2087 (O_2087,N_22624,N_23670);
and UO_2088 (O_2088,N_23767,N_24842);
nor UO_2089 (O_2089,N_24474,N_24942);
and UO_2090 (O_2090,N_24891,N_24079);
nand UO_2091 (O_2091,N_22711,N_23527);
xor UO_2092 (O_2092,N_23625,N_23762);
nor UO_2093 (O_2093,N_22552,N_23764);
or UO_2094 (O_2094,N_24739,N_24927);
nand UO_2095 (O_2095,N_23038,N_23806);
xor UO_2096 (O_2096,N_22695,N_22668);
and UO_2097 (O_2097,N_23526,N_24103);
nor UO_2098 (O_2098,N_23508,N_24324);
nand UO_2099 (O_2099,N_23273,N_22833);
xor UO_2100 (O_2100,N_22539,N_24628);
or UO_2101 (O_2101,N_24260,N_23335);
xor UO_2102 (O_2102,N_23925,N_22918);
and UO_2103 (O_2103,N_24192,N_22929);
and UO_2104 (O_2104,N_23275,N_24892);
nand UO_2105 (O_2105,N_24808,N_23931);
and UO_2106 (O_2106,N_24791,N_22707);
or UO_2107 (O_2107,N_23622,N_23683);
and UO_2108 (O_2108,N_24342,N_22872);
nand UO_2109 (O_2109,N_23205,N_23793);
or UO_2110 (O_2110,N_22958,N_22683);
xnor UO_2111 (O_2111,N_23486,N_24538);
xor UO_2112 (O_2112,N_22740,N_24834);
nand UO_2113 (O_2113,N_23449,N_23100);
nor UO_2114 (O_2114,N_22957,N_24191);
and UO_2115 (O_2115,N_23804,N_23467);
or UO_2116 (O_2116,N_24932,N_24760);
nor UO_2117 (O_2117,N_24657,N_23271);
nor UO_2118 (O_2118,N_23573,N_23006);
or UO_2119 (O_2119,N_22588,N_23195);
xor UO_2120 (O_2120,N_23001,N_24849);
nand UO_2121 (O_2121,N_24892,N_22761);
nor UO_2122 (O_2122,N_23393,N_24995);
xor UO_2123 (O_2123,N_23978,N_22900);
xnor UO_2124 (O_2124,N_23759,N_23675);
or UO_2125 (O_2125,N_24756,N_22794);
nor UO_2126 (O_2126,N_24498,N_22799);
xnor UO_2127 (O_2127,N_23673,N_24252);
nand UO_2128 (O_2128,N_22806,N_24665);
and UO_2129 (O_2129,N_23161,N_24423);
nor UO_2130 (O_2130,N_22767,N_22931);
or UO_2131 (O_2131,N_24735,N_22631);
nand UO_2132 (O_2132,N_24882,N_24366);
xnor UO_2133 (O_2133,N_23931,N_22997);
or UO_2134 (O_2134,N_22562,N_23155);
nor UO_2135 (O_2135,N_24975,N_24733);
nor UO_2136 (O_2136,N_24371,N_24955);
or UO_2137 (O_2137,N_22871,N_22978);
and UO_2138 (O_2138,N_24611,N_24001);
xnor UO_2139 (O_2139,N_22544,N_22992);
and UO_2140 (O_2140,N_23053,N_24815);
nand UO_2141 (O_2141,N_22817,N_24449);
xor UO_2142 (O_2142,N_22735,N_24460);
nand UO_2143 (O_2143,N_23182,N_23542);
nand UO_2144 (O_2144,N_24422,N_22893);
nand UO_2145 (O_2145,N_24815,N_23291);
xor UO_2146 (O_2146,N_24032,N_22541);
nand UO_2147 (O_2147,N_24530,N_24406);
xnor UO_2148 (O_2148,N_24312,N_24443);
nand UO_2149 (O_2149,N_22787,N_22925);
or UO_2150 (O_2150,N_23655,N_23626);
or UO_2151 (O_2151,N_22717,N_22680);
and UO_2152 (O_2152,N_23658,N_24049);
and UO_2153 (O_2153,N_23656,N_24284);
nand UO_2154 (O_2154,N_24309,N_24450);
nor UO_2155 (O_2155,N_23210,N_24088);
nor UO_2156 (O_2156,N_24111,N_23880);
or UO_2157 (O_2157,N_24910,N_22889);
and UO_2158 (O_2158,N_22534,N_23219);
nand UO_2159 (O_2159,N_23031,N_23830);
and UO_2160 (O_2160,N_24379,N_23591);
and UO_2161 (O_2161,N_24927,N_24527);
or UO_2162 (O_2162,N_22583,N_24877);
xnor UO_2163 (O_2163,N_22729,N_24806);
or UO_2164 (O_2164,N_23439,N_22771);
and UO_2165 (O_2165,N_23282,N_22678);
or UO_2166 (O_2166,N_23416,N_23914);
or UO_2167 (O_2167,N_24562,N_22763);
xnor UO_2168 (O_2168,N_23167,N_24528);
nor UO_2169 (O_2169,N_24298,N_23064);
nor UO_2170 (O_2170,N_23582,N_22992);
nor UO_2171 (O_2171,N_22850,N_24308);
nand UO_2172 (O_2172,N_24495,N_22517);
xor UO_2173 (O_2173,N_22830,N_24430);
or UO_2174 (O_2174,N_24729,N_23400);
and UO_2175 (O_2175,N_23372,N_23275);
xnor UO_2176 (O_2176,N_23656,N_24696);
xor UO_2177 (O_2177,N_24820,N_24949);
xnor UO_2178 (O_2178,N_23311,N_24005);
and UO_2179 (O_2179,N_23225,N_23374);
nor UO_2180 (O_2180,N_23685,N_23313);
xor UO_2181 (O_2181,N_24227,N_24296);
or UO_2182 (O_2182,N_24078,N_23689);
nand UO_2183 (O_2183,N_23590,N_23344);
or UO_2184 (O_2184,N_24946,N_24153);
and UO_2185 (O_2185,N_23554,N_24294);
and UO_2186 (O_2186,N_24265,N_22690);
and UO_2187 (O_2187,N_23815,N_24587);
xnor UO_2188 (O_2188,N_22644,N_24745);
xor UO_2189 (O_2189,N_23477,N_24945);
nor UO_2190 (O_2190,N_24683,N_23013);
nor UO_2191 (O_2191,N_23215,N_23007);
xnor UO_2192 (O_2192,N_24292,N_23664);
nor UO_2193 (O_2193,N_23372,N_23395);
nand UO_2194 (O_2194,N_24058,N_22906);
or UO_2195 (O_2195,N_23351,N_23773);
or UO_2196 (O_2196,N_23982,N_24169);
nor UO_2197 (O_2197,N_23047,N_23319);
or UO_2198 (O_2198,N_24430,N_23083);
or UO_2199 (O_2199,N_23365,N_24049);
nand UO_2200 (O_2200,N_23674,N_24843);
xor UO_2201 (O_2201,N_22601,N_23925);
or UO_2202 (O_2202,N_24236,N_24779);
nor UO_2203 (O_2203,N_23355,N_24454);
or UO_2204 (O_2204,N_24411,N_24507);
nand UO_2205 (O_2205,N_22957,N_24427);
nand UO_2206 (O_2206,N_24183,N_22887);
or UO_2207 (O_2207,N_23955,N_22816);
xnor UO_2208 (O_2208,N_23099,N_23709);
nor UO_2209 (O_2209,N_24615,N_22894);
nor UO_2210 (O_2210,N_22776,N_23388);
nand UO_2211 (O_2211,N_23001,N_24024);
and UO_2212 (O_2212,N_24728,N_23635);
or UO_2213 (O_2213,N_23396,N_24099);
nand UO_2214 (O_2214,N_23841,N_23770);
and UO_2215 (O_2215,N_23458,N_24104);
and UO_2216 (O_2216,N_24983,N_23357);
xnor UO_2217 (O_2217,N_24176,N_23911);
nor UO_2218 (O_2218,N_24291,N_24762);
or UO_2219 (O_2219,N_23011,N_23818);
and UO_2220 (O_2220,N_24604,N_22690);
and UO_2221 (O_2221,N_24432,N_23028);
or UO_2222 (O_2222,N_23496,N_24160);
nand UO_2223 (O_2223,N_24078,N_24123);
nor UO_2224 (O_2224,N_23203,N_24885);
nor UO_2225 (O_2225,N_24539,N_22943);
and UO_2226 (O_2226,N_23928,N_23351);
or UO_2227 (O_2227,N_24834,N_22660);
or UO_2228 (O_2228,N_23046,N_22977);
nand UO_2229 (O_2229,N_22513,N_24523);
xor UO_2230 (O_2230,N_24445,N_23460);
or UO_2231 (O_2231,N_23027,N_24279);
nor UO_2232 (O_2232,N_22604,N_22548);
nor UO_2233 (O_2233,N_24253,N_22808);
nor UO_2234 (O_2234,N_24078,N_24431);
and UO_2235 (O_2235,N_22915,N_23573);
xnor UO_2236 (O_2236,N_22871,N_24937);
nand UO_2237 (O_2237,N_24405,N_23513);
nand UO_2238 (O_2238,N_24295,N_23293);
and UO_2239 (O_2239,N_24508,N_23103);
nand UO_2240 (O_2240,N_23601,N_22566);
and UO_2241 (O_2241,N_24251,N_24731);
nand UO_2242 (O_2242,N_23904,N_24785);
and UO_2243 (O_2243,N_23996,N_24997);
nand UO_2244 (O_2244,N_23470,N_24127);
or UO_2245 (O_2245,N_24675,N_24239);
nor UO_2246 (O_2246,N_22517,N_24515);
nor UO_2247 (O_2247,N_24379,N_22962);
nor UO_2248 (O_2248,N_22775,N_23657);
xor UO_2249 (O_2249,N_23927,N_22929);
or UO_2250 (O_2250,N_23232,N_24439);
xnor UO_2251 (O_2251,N_23517,N_24406);
and UO_2252 (O_2252,N_24535,N_24881);
xnor UO_2253 (O_2253,N_24749,N_22724);
xnor UO_2254 (O_2254,N_24291,N_24674);
nand UO_2255 (O_2255,N_23985,N_23724);
or UO_2256 (O_2256,N_24258,N_22576);
and UO_2257 (O_2257,N_24929,N_23678);
and UO_2258 (O_2258,N_23311,N_23393);
nand UO_2259 (O_2259,N_22519,N_24936);
nand UO_2260 (O_2260,N_24973,N_24607);
nand UO_2261 (O_2261,N_23991,N_24865);
xnor UO_2262 (O_2262,N_22601,N_23444);
nor UO_2263 (O_2263,N_24698,N_22976);
and UO_2264 (O_2264,N_23793,N_22866);
or UO_2265 (O_2265,N_24424,N_22514);
xor UO_2266 (O_2266,N_24167,N_23205);
nor UO_2267 (O_2267,N_24884,N_24442);
xor UO_2268 (O_2268,N_23858,N_23179);
and UO_2269 (O_2269,N_24627,N_23739);
or UO_2270 (O_2270,N_22813,N_24641);
nor UO_2271 (O_2271,N_24110,N_23440);
and UO_2272 (O_2272,N_22738,N_23617);
xnor UO_2273 (O_2273,N_22654,N_22764);
and UO_2274 (O_2274,N_24697,N_23357);
and UO_2275 (O_2275,N_23292,N_23662);
and UO_2276 (O_2276,N_24048,N_23617);
xnor UO_2277 (O_2277,N_24322,N_23724);
nor UO_2278 (O_2278,N_23644,N_24903);
nor UO_2279 (O_2279,N_24087,N_23260);
and UO_2280 (O_2280,N_23938,N_24045);
nor UO_2281 (O_2281,N_23137,N_23047);
nand UO_2282 (O_2282,N_22664,N_24718);
nand UO_2283 (O_2283,N_23522,N_23492);
or UO_2284 (O_2284,N_23214,N_22913);
nand UO_2285 (O_2285,N_23612,N_22603);
nand UO_2286 (O_2286,N_22575,N_22902);
or UO_2287 (O_2287,N_23060,N_23592);
nor UO_2288 (O_2288,N_24554,N_24874);
nand UO_2289 (O_2289,N_24135,N_24303);
and UO_2290 (O_2290,N_23054,N_24513);
nand UO_2291 (O_2291,N_23999,N_23779);
nor UO_2292 (O_2292,N_24368,N_23314);
nand UO_2293 (O_2293,N_24514,N_24120);
nand UO_2294 (O_2294,N_24799,N_23720);
and UO_2295 (O_2295,N_24510,N_23591);
nor UO_2296 (O_2296,N_24849,N_23152);
nand UO_2297 (O_2297,N_23148,N_24259);
nor UO_2298 (O_2298,N_23443,N_22768);
nand UO_2299 (O_2299,N_24456,N_24551);
or UO_2300 (O_2300,N_23860,N_22799);
or UO_2301 (O_2301,N_23596,N_23031);
nor UO_2302 (O_2302,N_22662,N_24063);
or UO_2303 (O_2303,N_24738,N_22615);
nor UO_2304 (O_2304,N_24303,N_24924);
xnor UO_2305 (O_2305,N_23557,N_22996);
or UO_2306 (O_2306,N_23531,N_24983);
nand UO_2307 (O_2307,N_23413,N_22626);
xnor UO_2308 (O_2308,N_22832,N_24183);
or UO_2309 (O_2309,N_23571,N_23537);
xor UO_2310 (O_2310,N_22804,N_23855);
and UO_2311 (O_2311,N_24578,N_23870);
nand UO_2312 (O_2312,N_24648,N_24164);
or UO_2313 (O_2313,N_24691,N_24266);
nor UO_2314 (O_2314,N_23580,N_23533);
nor UO_2315 (O_2315,N_24280,N_22971);
and UO_2316 (O_2316,N_24374,N_23141);
xor UO_2317 (O_2317,N_24420,N_24648);
xor UO_2318 (O_2318,N_23761,N_23794);
and UO_2319 (O_2319,N_24256,N_24456);
nor UO_2320 (O_2320,N_23211,N_23166);
xnor UO_2321 (O_2321,N_22511,N_23270);
nor UO_2322 (O_2322,N_24225,N_23509);
xor UO_2323 (O_2323,N_23164,N_24313);
nor UO_2324 (O_2324,N_24655,N_22554);
and UO_2325 (O_2325,N_23014,N_22725);
and UO_2326 (O_2326,N_22502,N_24868);
or UO_2327 (O_2327,N_24392,N_23906);
or UO_2328 (O_2328,N_23648,N_23003);
xor UO_2329 (O_2329,N_24575,N_22938);
and UO_2330 (O_2330,N_23982,N_24936);
nor UO_2331 (O_2331,N_24073,N_24017);
and UO_2332 (O_2332,N_23642,N_23871);
or UO_2333 (O_2333,N_24832,N_23118);
or UO_2334 (O_2334,N_23710,N_23984);
nand UO_2335 (O_2335,N_24935,N_24142);
nand UO_2336 (O_2336,N_24431,N_23366);
nand UO_2337 (O_2337,N_23289,N_24526);
xor UO_2338 (O_2338,N_23942,N_23971);
nor UO_2339 (O_2339,N_23743,N_24924);
and UO_2340 (O_2340,N_23617,N_22708);
xnor UO_2341 (O_2341,N_23799,N_24638);
xor UO_2342 (O_2342,N_23336,N_23623);
nor UO_2343 (O_2343,N_23448,N_24413);
and UO_2344 (O_2344,N_23970,N_22547);
and UO_2345 (O_2345,N_22852,N_22905);
nor UO_2346 (O_2346,N_22726,N_23715);
nor UO_2347 (O_2347,N_23734,N_24161);
xnor UO_2348 (O_2348,N_22948,N_24482);
and UO_2349 (O_2349,N_23263,N_23503);
nor UO_2350 (O_2350,N_24600,N_22709);
nor UO_2351 (O_2351,N_22539,N_24791);
or UO_2352 (O_2352,N_24195,N_23422);
or UO_2353 (O_2353,N_24341,N_24661);
xnor UO_2354 (O_2354,N_24509,N_23886);
xnor UO_2355 (O_2355,N_24864,N_24808);
xor UO_2356 (O_2356,N_23478,N_23367);
nand UO_2357 (O_2357,N_24755,N_24485);
xor UO_2358 (O_2358,N_24590,N_22517);
xor UO_2359 (O_2359,N_22743,N_23236);
and UO_2360 (O_2360,N_24254,N_24948);
and UO_2361 (O_2361,N_22712,N_24780);
nor UO_2362 (O_2362,N_24600,N_24123);
nand UO_2363 (O_2363,N_22810,N_24877);
nor UO_2364 (O_2364,N_24829,N_24168);
or UO_2365 (O_2365,N_23138,N_23664);
nor UO_2366 (O_2366,N_24301,N_23348);
or UO_2367 (O_2367,N_24851,N_23455);
nand UO_2368 (O_2368,N_23416,N_24030);
nor UO_2369 (O_2369,N_23538,N_24875);
or UO_2370 (O_2370,N_24393,N_24170);
nor UO_2371 (O_2371,N_23423,N_24566);
nand UO_2372 (O_2372,N_24728,N_22505);
nand UO_2373 (O_2373,N_23987,N_23839);
nor UO_2374 (O_2374,N_24897,N_24008);
and UO_2375 (O_2375,N_24044,N_23368);
nor UO_2376 (O_2376,N_23867,N_24826);
nand UO_2377 (O_2377,N_23506,N_24076);
nor UO_2378 (O_2378,N_23045,N_24108);
nand UO_2379 (O_2379,N_24163,N_23480);
xnor UO_2380 (O_2380,N_22582,N_22563);
or UO_2381 (O_2381,N_24410,N_23393);
and UO_2382 (O_2382,N_24053,N_24524);
or UO_2383 (O_2383,N_22915,N_24214);
or UO_2384 (O_2384,N_24772,N_22634);
xnor UO_2385 (O_2385,N_23021,N_23747);
nand UO_2386 (O_2386,N_23854,N_23231);
nor UO_2387 (O_2387,N_24531,N_24972);
xor UO_2388 (O_2388,N_22766,N_22668);
xor UO_2389 (O_2389,N_24507,N_24401);
nor UO_2390 (O_2390,N_24066,N_23604);
or UO_2391 (O_2391,N_23658,N_23465);
or UO_2392 (O_2392,N_24780,N_23867);
nor UO_2393 (O_2393,N_22989,N_24448);
xor UO_2394 (O_2394,N_22802,N_24750);
nand UO_2395 (O_2395,N_24579,N_23700);
or UO_2396 (O_2396,N_24697,N_23820);
xnor UO_2397 (O_2397,N_24289,N_24882);
or UO_2398 (O_2398,N_23644,N_24797);
nand UO_2399 (O_2399,N_23862,N_24370);
xnor UO_2400 (O_2400,N_22625,N_24373);
or UO_2401 (O_2401,N_24140,N_22718);
or UO_2402 (O_2402,N_24836,N_24229);
xor UO_2403 (O_2403,N_24560,N_24667);
nor UO_2404 (O_2404,N_23467,N_24601);
xor UO_2405 (O_2405,N_23949,N_23853);
or UO_2406 (O_2406,N_24068,N_23982);
or UO_2407 (O_2407,N_24971,N_24396);
or UO_2408 (O_2408,N_24561,N_24235);
xnor UO_2409 (O_2409,N_23779,N_23335);
or UO_2410 (O_2410,N_23186,N_24772);
and UO_2411 (O_2411,N_23010,N_24195);
xor UO_2412 (O_2412,N_23194,N_24806);
and UO_2413 (O_2413,N_22556,N_24139);
xnor UO_2414 (O_2414,N_24408,N_24108);
nor UO_2415 (O_2415,N_24332,N_22849);
xnor UO_2416 (O_2416,N_22566,N_23506);
xnor UO_2417 (O_2417,N_22522,N_24339);
or UO_2418 (O_2418,N_24347,N_24711);
xnor UO_2419 (O_2419,N_22682,N_24153);
or UO_2420 (O_2420,N_23567,N_24403);
xor UO_2421 (O_2421,N_24965,N_22992);
xor UO_2422 (O_2422,N_23366,N_24749);
nand UO_2423 (O_2423,N_22838,N_23748);
xor UO_2424 (O_2424,N_22684,N_24617);
or UO_2425 (O_2425,N_24154,N_23095);
and UO_2426 (O_2426,N_22790,N_24934);
xnor UO_2427 (O_2427,N_23398,N_23820);
and UO_2428 (O_2428,N_22536,N_22600);
or UO_2429 (O_2429,N_23873,N_23908);
xnor UO_2430 (O_2430,N_24303,N_24997);
or UO_2431 (O_2431,N_23469,N_23775);
nand UO_2432 (O_2432,N_24005,N_23926);
or UO_2433 (O_2433,N_24691,N_23028);
nor UO_2434 (O_2434,N_23479,N_22888);
xor UO_2435 (O_2435,N_22811,N_23621);
or UO_2436 (O_2436,N_23460,N_22717);
nand UO_2437 (O_2437,N_24534,N_23830);
xor UO_2438 (O_2438,N_24726,N_22578);
xor UO_2439 (O_2439,N_24438,N_22666);
xor UO_2440 (O_2440,N_22726,N_23782);
or UO_2441 (O_2441,N_22707,N_23177);
nand UO_2442 (O_2442,N_24674,N_23700);
and UO_2443 (O_2443,N_23813,N_24387);
nor UO_2444 (O_2444,N_24817,N_22939);
and UO_2445 (O_2445,N_22735,N_22974);
xnor UO_2446 (O_2446,N_23921,N_22818);
nand UO_2447 (O_2447,N_24392,N_24075);
nor UO_2448 (O_2448,N_23697,N_22930);
and UO_2449 (O_2449,N_23460,N_22832);
xnor UO_2450 (O_2450,N_23740,N_24013);
and UO_2451 (O_2451,N_23577,N_24986);
and UO_2452 (O_2452,N_23262,N_24731);
nor UO_2453 (O_2453,N_24167,N_23788);
and UO_2454 (O_2454,N_24175,N_24844);
nand UO_2455 (O_2455,N_23982,N_24506);
nand UO_2456 (O_2456,N_23176,N_24350);
and UO_2457 (O_2457,N_23870,N_24486);
nor UO_2458 (O_2458,N_24658,N_24766);
nand UO_2459 (O_2459,N_23609,N_24423);
and UO_2460 (O_2460,N_23847,N_22969);
nand UO_2461 (O_2461,N_23090,N_23212);
xnor UO_2462 (O_2462,N_24146,N_24716);
xnor UO_2463 (O_2463,N_23598,N_24830);
nor UO_2464 (O_2464,N_23440,N_23225);
and UO_2465 (O_2465,N_22652,N_24606);
nand UO_2466 (O_2466,N_23447,N_24917);
nand UO_2467 (O_2467,N_23025,N_24180);
or UO_2468 (O_2468,N_23736,N_23462);
xnor UO_2469 (O_2469,N_24582,N_24278);
and UO_2470 (O_2470,N_23611,N_24219);
or UO_2471 (O_2471,N_24439,N_24017);
xor UO_2472 (O_2472,N_23389,N_22820);
xnor UO_2473 (O_2473,N_23489,N_23422);
xor UO_2474 (O_2474,N_24259,N_23575);
nor UO_2475 (O_2475,N_24707,N_22974);
nand UO_2476 (O_2476,N_24002,N_24720);
nor UO_2477 (O_2477,N_24861,N_24459);
nor UO_2478 (O_2478,N_24911,N_22830);
nor UO_2479 (O_2479,N_24706,N_24880);
nand UO_2480 (O_2480,N_24789,N_24618);
and UO_2481 (O_2481,N_24493,N_23956);
or UO_2482 (O_2482,N_23711,N_24558);
or UO_2483 (O_2483,N_22854,N_24716);
nor UO_2484 (O_2484,N_22963,N_24933);
or UO_2485 (O_2485,N_22531,N_24920);
nand UO_2486 (O_2486,N_23865,N_23007);
nand UO_2487 (O_2487,N_22713,N_22832);
xor UO_2488 (O_2488,N_22525,N_24462);
or UO_2489 (O_2489,N_23686,N_24431);
nand UO_2490 (O_2490,N_23082,N_24938);
and UO_2491 (O_2491,N_23399,N_24472);
nand UO_2492 (O_2492,N_24450,N_24382);
xor UO_2493 (O_2493,N_24539,N_23330);
xor UO_2494 (O_2494,N_23373,N_23344);
nor UO_2495 (O_2495,N_22528,N_23173);
and UO_2496 (O_2496,N_24745,N_22721);
or UO_2497 (O_2497,N_23107,N_24437);
nand UO_2498 (O_2498,N_23642,N_23580);
nand UO_2499 (O_2499,N_22727,N_23144);
nor UO_2500 (O_2500,N_23359,N_24811);
and UO_2501 (O_2501,N_24478,N_23421);
nand UO_2502 (O_2502,N_23483,N_24757);
nand UO_2503 (O_2503,N_23888,N_23712);
xnor UO_2504 (O_2504,N_23612,N_23263);
nand UO_2505 (O_2505,N_24579,N_24169);
nand UO_2506 (O_2506,N_24020,N_23799);
and UO_2507 (O_2507,N_24631,N_23052);
nor UO_2508 (O_2508,N_24371,N_22789);
nor UO_2509 (O_2509,N_23322,N_23907);
or UO_2510 (O_2510,N_24900,N_23201);
or UO_2511 (O_2511,N_24224,N_23454);
xor UO_2512 (O_2512,N_23177,N_22566);
nand UO_2513 (O_2513,N_24665,N_23716);
xnor UO_2514 (O_2514,N_23759,N_23637);
nand UO_2515 (O_2515,N_23445,N_23184);
and UO_2516 (O_2516,N_24499,N_24862);
and UO_2517 (O_2517,N_23950,N_22793);
and UO_2518 (O_2518,N_23722,N_22913);
and UO_2519 (O_2519,N_24522,N_24333);
nand UO_2520 (O_2520,N_23941,N_23591);
nor UO_2521 (O_2521,N_23940,N_24400);
nor UO_2522 (O_2522,N_23977,N_23691);
nor UO_2523 (O_2523,N_24529,N_24053);
and UO_2524 (O_2524,N_23893,N_23789);
nor UO_2525 (O_2525,N_24532,N_22932);
nand UO_2526 (O_2526,N_23258,N_23567);
nand UO_2527 (O_2527,N_24461,N_22800);
nor UO_2528 (O_2528,N_24272,N_24537);
nand UO_2529 (O_2529,N_23346,N_24368);
nand UO_2530 (O_2530,N_23040,N_22834);
nand UO_2531 (O_2531,N_24872,N_22766);
or UO_2532 (O_2532,N_24027,N_23809);
or UO_2533 (O_2533,N_22749,N_23868);
and UO_2534 (O_2534,N_23449,N_24719);
xor UO_2535 (O_2535,N_23176,N_23369);
or UO_2536 (O_2536,N_22737,N_24814);
nor UO_2537 (O_2537,N_24388,N_23302);
xor UO_2538 (O_2538,N_24104,N_24554);
and UO_2539 (O_2539,N_23556,N_22547);
nor UO_2540 (O_2540,N_24791,N_24549);
and UO_2541 (O_2541,N_23088,N_24471);
nand UO_2542 (O_2542,N_24300,N_23619);
or UO_2543 (O_2543,N_23427,N_23537);
and UO_2544 (O_2544,N_22511,N_23264);
and UO_2545 (O_2545,N_24967,N_24113);
nor UO_2546 (O_2546,N_22977,N_24185);
and UO_2547 (O_2547,N_23168,N_23817);
xnor UO_2548 (O_2548,N_23453,N_24325);
or UO_2549 (O_2549,N_23208,N_23978);
xor UO_2550 (O_2550,N_22602,N_23340);
nand UO_2551 (O_2551,N_23627,N_23749);
and UO_2552 (O_2552,N_22750,N_22859);
nand UO_2553 (O_2553,N_24110,N_22802);
and UO_2554 (O_2554,N_24023,N_23030);
or UO_2555 (O_2555,N_22737,N_23238);
or UO_2556 (O_2556,N_23423,N_24026);
nor UO_2557 (O_2557,N_24937,N_22708);
xor UO_2558 (O_2558,N_24306,N_23396);
nand UO_2559 (O_2559,N_24139,N_24508);
or UO_2560 (O_2560,N_24947,N_23183);
xnor UO_2561 (O_2561,N_23347,N_24380);
xor UO_2562 (O_2562,N_23061,N_23715);
and UO_2563 (O_2563,N_24442,N_23968);
nand UO_2564 (O_2564,N_22597,N_24562);
nand UO_2565 (O_2565,N_22959,N_23334);
or UO_2566 (O_2566,N_22532,N_24736);
xnor UO_2567 (O_2567,N_22657,N_23464);
and UO_2568 (O_2568,N_24319,N_22811);
nor UO_2569 (O_2569,N_23000,N_22931);
or UO_2570 (O_2570,N_24244,N_23837);
xnor UO_2571 (O_2571,N_23764,N_22891);
or UO_2572 (O_2572,N_23532,N_24284);
nor UO_2573 (O_2573,N_23352,N_23895);
or UO_2574 (O_2574,N_23054,N_24422);
xnor UO_2575 (O_2575,N_24446,N_22788);
nand UO_2576 (O_2576,N_24736,N_22700);
xnor UO_2577 (O_2577,N_23084,N_24248);
or UO_2578 (O_2578,N_24527,N_22537);
nor UO_2579 (O_2579,N_24454,N_24087);
xnor UO_2580 (O_2580,N_24401,N_24106);
nor UO_2581 (O_2581,N_22941,N_24529);
nand UO_2582 (O_2582,N_23711,N_22580);
nand UO_2583 (O_2583,N_24050,N_22986);
nand UO_2584 (O_2584,N_24674,N_22686);
xor UO_2585 (O_2585,N_23793,N_23700);
or UO_2586 (O_2586,N_24372,N_24397);
xor UO_2587 (O_2587,N_24572,N_23646);
nor UO_2588 (O_2588,N_23266,N_24685);
nor UO_2589 (O_2589,N_23720,N_24384);
or UO_2590 (O_2590,N_24058,N_24250);
or UO_2591 (O_2591,N_24881,N_23003);
and UO_2592 (O_2592,N_23539,N_23055);
nand UO_2593 (O_2593,N_23449,N_24041);
nor UO_2594 (O_2594,N_23292,N_24162);
xor UO_2595 (O_2595,N_23488,N_23602);
or UO_2596 (O_2596,N_22991,N_22946);
and UO_2597 (O_2597,N_24097,N_24620);
xor UO_2598 (O_2598,N_24964,N_24034);
or UO_2599 (O_2599,N_22850,N_23402);
nor UO_2600 (O_2600,N_24099,N_22557);
or UO_2601 (O_2601,N_23654,N_22604);
xor UO_2602 (O_2602,N_22604,N_24530);
nor UO_2603 (O_2603,N_24343,N_23438);
and UO_2604 (O_2604,N_24010,N_24262);
and UO_2605 (O_2605,N_24773,N_24202);
xor UO_2606 (O_2606,N_23151,N_24800);
nand UO_2607 (O_2607,N_24331,N_22735);
nand UO_2608 (O_2608,N_24809,N_22919);
and UO_2609 (O_2609,N_22643,N_24323);
or UO_2610 (O_2610,N_23468,N_23210);
or UO_2611 (O_2611,N_24870,N_22584);
and UO_2612 (O_2612,N_24601,N_23526);
nand UO_2613 (O_2613,N_22873,N_24366);
xor UO_2614 (O_2614,N_24869,N_23342);
and UO_2615 (O_2615,N_23040,N_24418);
xnor UO_2616 (O_2616,N_23299,N_23675);
xor UO_2617 (O_2617,N_22757,N_22504);
or UO_2618 (O_2618,N_24284,N_24170);
nor UO_2619 (O_2619,N_23367,N_22507);
nor UO_2620 (O_2620,N_24038,N_23777);
and UO_2621 (O_2621,N_23526,N_24327);
xor UO_2622 (O_2622,N_24769,N_23022);
and UO_2623 (O_2623,N_23592,N_24564);
nor UO_2624 (O_2624,N_24499,N_23395);
and UO_2625 (O_2625,N_24240,N_22808);
and UO_2626 (O_2626,N_22887,N_24748);
and UO_2627 (O_2627,N_24935,N_24508);
xor UO_2628 (O_2628,N_24101,N_24376);
or UO_2629 (O_2629,N_24530,N_23099);
and UO_2630 (O_2630,N_22860,N_24993);
and UO_2631 (O_2631,N_24309,N_23331);
and UO_2632 (O_2632,N_24638,N_23323);
xnor UO_2633 (O_2633,N_24808,N_24222);
and UO_2634 (O_2634,N_22873,N_24962);
nor UO_2635 (O_2635,N_24594,N_24704);
xor UO_2636 (O_2636,N_24593,N_24672);
nand UO_2637 (O_2637,N_22952,N_23527);
and UO_2638 (O_2638,N_24536,N_24202);
nor UO_2639 (O_2639,N_23448,N_23389);
xnor UO_2640 (O_2640,N_24326,N_23252);
xor UO_2641 (O_2641,N_24096,N_24022);
and UO_2642 (O_2642,N_24042,N_24863);
nor UO_2643 (O_2643,N_22710,N_23199);
and UO_2644 (O_2644,N_22561,N_24155);
and UO_2645 (O_2645,N_22976,N_23507);
nand UO_2646 (O_2646,N_24803,N_24110);
nand UO_2647 (O_2647,N_22813,N_22864);
xnor UO_2648 (O_2648,N_22774,N_24496);
nor UO_2649 (O_2649,N_24730,N_22691);
xnor UO_2650 (O_2650,N_24400,N_23528);
xor UO_2651 (O_2651,N_22992,N_22963);
nand UO_2652 (O_2652,N_24512,N_23859);
and UO_2653 (O_2653,N_23324,N_22840);
xnor UO_2654 (O_2654,N_24764,N_24020);
and UO_2655 (O_2655,N_23748,N_23487);
and UO_2656 (O_2656,N_22902,N_22698);
xor UO_2657 (O_2657,N_24123,N_22783);
nand UO_2658 (O_2658,N_24240,N_23757);
xnor UO_2659 (O_2659,N_24306,N_24901);
or UO_2660 (O_2660,N_24365,N_23364);
xor UO_2661 (O_2661,N_22998,N_23347);
nand UO_2662 (O_2662,N_22829,N_22596);
xnor UO_2663 (O_2663,N_23887,N_24574);
or UO_2664 (O_2664,N_24834,N_24336);
and UO_2665 (O_2665,N_22694,N_23857);
or UO_2666 (O_2666,N_24853,N_24134);
and UO_2667 (O_2667,N_23856,N_24231);
and UO_2668 (O_2668,N_23159,N_23232);
or UO_2669 (O_2669,N_23107,N_22985);
or UO_2670 (O_2670,N_24315,N_24745);
nor UO_2671 (O_2671,N_22529,N_24552);
or UO_2672 (O_2672,N_24363,N_23690);
nor UO_2673 (O_2673,N_23118,N_23630);
nor UO_2674 (O_2674,N_22924,N_24851);
and UO_2675 (O_2675,N_24412,N_24641);
nor UO_2676 (O_2676,N_22761,N_23083);
or UO_2677 (O_2677,N_23100,N_23565);
and UO_2678 (O_2678,N_23639,N_23052);
xor UO_2679 (O_2679,N_23919,N_24722);
xor UO_2680 (O_2680,N_23877,N_24969);
xnor UO_2681 (O_2681,N_24776,N_22625);
and UO_2682 (O_2682,N_23785,N_22704);
or UO_2683 (O_2683,N_23828,N_24489);
nand UO_2684 (O_2684,N_23477,N_24339);
or UO_2685 (O_2685,N_23553,N_24300);
xor UO_2686 (O_2686,N_23764,N_22737);
or UO_2687 (O_2687,N_22836,N_22656);
nand UO_2688 (O_2688,N_24617,N_24043);
and UO_2689 (O_2689,N_24926,N_24950);
or UO_2690 (O_2690,N_24644,N_23737);
and UO_2691 (O_2691,N_23192,N_23982);
nand UO_2692 (O_2692,N_22796,N_22762);
nor UO_2693 (O_2693,N_24850,N_24842);
nand UO_2694 (O_2694,N_24917,N_23348);
xor UO_2695 (O_2695,N_24734,N_24242);
and UO_2696 (O_2696,N_24442,N_23188);
nand UO_2697 (O_2697,N_22671,N_24065);
nor UO_2698 (O_2698,N_24749,N_22602);
nand UO_2699 (O_2699,N_23617,N_23989);
nor UO_2700 (O_2700,N_22953,N_22613);
or UO_2701 (O_2701,N_23020,N_24216);
and UO_2702 (O_2702,N_23796,N_24034);
or UO_2703 (O_2703,N_24741,N_24967);
nor UO_2704 (O_2704,N_24947,N_23476);
nand UO_2705 (O_2705,N_24026,N_24229);
xor UO_2706 (O_2706,N_23791,N_24573);
nand UO_2707 (O_2707,N_24097,N_23048);
nand UO_2708 (O_2708,N_24172,N_24762);
and UO_2709 (O_2709,N_23710,N_22923);
xnor UO_2710 (O_2710,N_23039,N_23034);
nor UO_2711 (O_2711,N_23159,N_22640);
nand UO_2712 (O_2712,N_24840,N_23409);
nand UO_2713 (O_2713,N_23461,N_24127);
and UO_2714 (O_2714,N_22546,N_24186);
or UO_2715 (O_2715,N_22953,N_23877);
nand UO_2716 (O_2716,N_24373,N_23416);
xor UO_2717 (O_2717,N_23676,N_24100);
xor UO_2718 (O_2718,N_23472,N_24932);
and UO_2719 (O_2719,N_24721,N_24686);
nand UO_2720 (O_2720,N_23983,N_24026);
or UO_2721 (O_2721,N_23758,N_23622);
nor UO_2722 (O_2722,N_24655,N_23319);
or UO_2723 (O_2723,N_22627,N_24886);
nand UO_2724 (O_2724,N_23510,N_22591);
or UO_2725 (O_2725,N_22554,N_22507);
and UO_2726 (O_2726,N_24604,N_23877);
nor UO_2727 (O_2727,N_23200,N_24314);
and UO_2728 (O_2728,N_24232,N_22727);
xnor UO_2729 (O_2729,N_22548,N_22970);
and UO_2730 (O_2730,N_23690,N_23365);
nand UO_2731 (O_2731,N_24145,N_24065);
nand UO_2732 (O_2732,N_23097,N_24709);
xor UO_2733 (O_2733,N_23134,N_22508);
xnor UO_2734 (O_2734,N_23251,N_23600);
nor UO_2735 (O_2735,N_24314,N_23573);
nand UO_2736 (O_2736,N_23802,N_23010);
nand UO_2737 (O_2737,N_22664,N_24977);
nand UO_2738 (O_2738,N_24311,N_23774);
xor UO_2739 (O_2739,N_24372,N_24087);
nand UO_2740 (O_2740,N_23467,N_23861);
or UO_2741 (O_2741,N_22996,N_24889);
and UO_2742 (O_2742,N_23241,N_23402);
xnor UO_2743 (O_2743,N_23674,N_23752);
xnor UO_2744 (O_2744,N_22933,N_22524);
nor UO_2745 (O_2745,N_24832,N_24391);
nor UO_2746 (O_2746,N_22713,N_22620);
and UO_2747 (O_2747,N_22552,N_22978);
or UO_2748 (O_2748,N_24345,N_24902);
and UO_2749 (O_2749,N_22549,N_23222);
and UO_2750 (O_2750,N_23474,N_24446);
or UO_2751 (O_2751,N_22610,N_23144);
xor UO_2752 (O_2752,N_23357,N_23286);
or UO_2753 (O_2753,N_24208,N_22975);
or UO_2754 (O_2754,N_22525,N_23444);
nor UO_2755 (O_2755,N_24634,N_22628);
or UO_2756 (O_2756,N_23609,N_23335);
nand UO_2757 (O_2757,N_24192,N_22680);
nand UO_2758 (O_2758,N_22835,N_23373);
xnor UO_2759 (O_2759,N_24319,N_23478);
or UO_2760 (O_2760,N_23543,N_24700);
nor UO_2761 (O_2761,N_22742,N_23508);
nand UO_2762 (O_2762,N_23552,N_23302);
or UO_2763 (O_2763,N_23977,N_22744);
nor UO_2764 (O_2764,N_23295,N_24793);
nand UO_2765 (O_2765,N_23668,N_23703);
and UO_2766 (O_2766,N_24970,N_24350);
nand UO_2767 (O_2767,N_23926,N_24544);
and UO_2768 (O_2768,N_23198,N_22908);
nor UO_2769 (O_2769,N_24697,N_23167);
nor UO_2770 (O_2770,N_24381,N_24074);
or UO_2771 (O_2771,N_24048,N_24928);
and UO_2772 (O_2772,N_24357,N_24903);
or UO_2773 (O_2773,N_23601,N_24950);
xnor UO_2774 (O_2774,N_24387,N_24558);
nand UO_2775 (O_2775,N_24610,N_23059);
or UO_2776 (O_2776,N_22665,N_22750);
xnor UO_2777 (O_2777,N_24884,N_22887);
xnor UO_2778 (O_2778,N_22934,N_24300);
nor UO_2779 (O_2779,N_23227,N_22709);
xnor UO_2780 (O_2780,N_24582,N_22746);
nand UO_2781 (O_2781,N_22656,N_23076);
nand UO_2782 (O_2782,N_23685,N_23865);
xor UO_2783 (O_2783,N_24603,N_23334);
or UO_2784 (O_2784,N_24034,N_23673);
nand UO_2785 (O_2785,N_23060,N_23605);
and UO_2786 (O_2786,N_23809,N_24231);
nor UO_2787 (O_2787,N_23272,N_23841);
or UO_2788 (O_2788,N_24093,N_23179);
or UO_2789 (O_2789,N_22673,N_24461);
nor UO_2790 (O_2790,N_24321,N_23812);
or UO_2791 (O_2791,N_24408,N_23184);
and UO_2792 (O_2792,N_22596,N_24666);
nand UO_2793 (O_2793,N_24510,N_23595);
nor UO_2794 (O_2794,N_24174,N_24921);
nand UO_2795 (O_2795,N_24050,N_23630);
xor UO_2796 (O_2796,N_24267,N_24300);
nor UO_2797 (O_2797,N_24889,N_23348);
and UO_2798 (O_2798,N_24057,N_22992);
nor UO_2799 (O_2799,N_24904,N_24233);
xor UO_2800 (O_2800,N_24833,N_23475);
or UO_2801 (O_2801,N_24096,N_22886);
xnor UO_2802 (O_2802,N_24800,N_23138);
xnor UO_2803 (O_2803,N_24331,N_23290);
nand UO_2804 (O_2804,N_23784,N_24759);
or UO_2805 (O_2805,N_23513,N_22932);
nand UO_2806 (O_2806,N_23461,N_24689);
xor UO_2807 (O_2807,N_22653,N_23348);
or UO_2808 (O_2808,N_23873,N_24180);
xor UO_2809 (O_2809,N_24340,N_23166);
nor UO_2810 (O_2810,N_22616,N_24939);
and UO_2811 (O_2811,N_23076,N_24012);
xnor UO_2812 (O_2812,N_23634,N_24282);
or UO_2813 (O_2813,N_23769,N_24874);
or UO_2814 (O_2814,N_23397,N_24107);
nor UO_2815 (O_2815,N_24028,N_24773);
and UO_2816 (O_2816,N_24886,N_22843);
xnor UO_2817 (O_2817,N_24089,N_23678);
and UO_2818 (O_2818,N_22529,N_24445);
xor UO_2819 (O_2819,N_23632,N_23345);
xnor UO_2820 (O_2820,N_23161,N_22679);
nor UO_2821 (O_2821,N_22645,N_24058);
and UO_2822 (O_2822,N_24781,N_24223);
or UO_2823 (O_2823,N_22889,N_23662);
or UO_2824 (O_2824,N_24731,N_23299);
or UO_2825 (O_2825,N_24941,N_24406);
nor UO_2826 (O_2826,N_23804,N_22813);
nor UO_2827 (O_2827,N_24512,N_24300);
nand UO_2828 (O_2828,N_24599,N_24069);
nor UO_2829 (O_2829,N_24077,N_24205);
nand UO_2830 (O_2830,N_23478,N_22619);
nor UO_2831 (O_2831,N_23261,N_24544);
nor UO_2832 (O_2832,N_23918,N_23691);
nand UO_2833 (O_2833,N_23758,N_24083);
nand UO_2834 (O_2834,N_23740,N_24188);
or UO_2835 (O_2835,N_24574,N_23503);
xor UO_2836 (O_2836,N_23567,N_23787);
xor UO_2837 (O_2837,N_23624,N_24603);
nor UO_2838 (O_2838,N_23049,N_24308);
or UO_2839 (O_2839,N_23620,N_23059);
nand UO_2840 (O_2840,N_23235,N_23183);
nor UO_2841 (O_2841,N_24777,N_22610);
xnor UO_2842 (O_2842,N_23196,N_24317);
and UO_2843 (O_2843,N_24350,N_23233);
nor UO_2844 (O_2844,N_24268,N_22884);
nand UO_2845 (O_2845,N_23080,N_23696);
or UO_2846 (O_2846,N_24160,N_23536);
and UO_2847 (O_2847,N_24496,N_22950);
or UO_2848 (O_2848,N_23641,N_23976);
xor UO_2849 (O_2849,N_22681,N_24490);
nand UO_2850 (O_2850,N_23549,N_23590);
and UO_2851 (O_2851,N_24314,N_24759);
or UO_2852 (O_2852,N_22828,N_23389);
and UO_2853 (O_2853,N_24888,N_22589);
nand UO_2854 (O_2854,N_24512,N_23105);
nand UO_2855 (O_2855,N_23427,N_23851);
xnor UO_2856 (O_2856,N_24201,N_24743);
xor UO_2857 (O_2857,N_22661,N_23570);
and UO_2858 (O_2858,N_23936,N_23162);
xnor UO_2859 (O_2859,N_22552,N_23922);
xor UO_2860 (O_2860,N_23029,N_23207);
xnor UO_2861 (O_2861,N_23226,N_22532);
nor UO_2862 (O_2862,N_24235,N_23144);
or UO_2863 (O_2863,N_23992,N_24299);
nand UO_2864 (O_2864,N_24663,N_23859);
and UO_2865 (O_2865,N_22836,N_24412);
or UO_2866 (O_2866,N_23034,N_23387);
nor UO_2867 (O_2867,N_23014,N_22903);
xnor UO_2868 (O_2868,N_24702,N_24183);
and UO_2869 (O_2869,N_23849,N_22596);
nand UO_2870 (O_2870,N_24879,N_23992);
nand UO_2871 (O_2871,N_23155,N_23838);
or UO_2872 (O_2872,N_23961,N_23827);
xor UO_2873 (O_2873,N_24261,N_23975);
nand UO_2874 (O_2874,N_23172,N_23592);
nor UO_2875 (O_2875,N_22538,N_22771);
and UO_2876 (O_2876,N_24675,N_24396);
or UO_2877 (O_2877,N_24027,N_22768);
and UO_2878 (O_2878,N_23804,N_24222);
xor UO_2879 (O_2879,N_23710,N_23727);
and UO_2880 (O_2880,N_23090,N_22834);
or UO_2881 (O_2881,N_23943,N_23051);
nor UO_2882 (O_2882,N_24020,N_23008);
xor UO_2883 (O_2883,N_23859,N_24562);
or UO_2884 (O_2884,N_23035,N_23584);
and UO_2885 (O_2885,N_23494,N_23175);
or UO_2886 (O_2886,N_23820,N_24535);
or UO_2887 (O_2887,N_22995,N_22639);
nor UO_2888 (O_2888,N_23900,N_24189);
nand UO_2889 (O_2889,N_24502,N_23517);
and UO_2890 (O_2890,N_22696,N_22919);
and UO_2891 (O_2891,N_24635,N_24445);
nand UO_2892 (O_2892,N_23173,N_23501);
nor UO_2893 (O_2893,N_24868,N_22984);
and UO_2894 (O_2894,N_23588,N_23348);
nand UO_2895 (O_2895,N_23577,N_24617);
xnor UO_2896 (O_2896,N_23987,N_24472);
nand UO_2897 (O_2897,N_23433,N_24978);
and UO_2898 (O_2898,N_24368,N_23893);
xor UO_2899 (O_2899,N_23930,N_24358);
and UO_2900 (O_2900,N_23324,N_23838);
and UO_2901 (O_2901,N_23840,N_24642);
nand UO_2902 (O_2902,N_23357,N_23508);
xnor UO_2903 (O_2903,N_22516,N_23554);
and UO_2904 (O_2904,N_23022,N_22915);
xnor UO_2905 (O_2905,N_23147,N_24771);
and UO_2906 (O_2906,N_22670,N_23461);
nand UO_2907 (O_2907,N_23495,N_23292);
nand UO_2908 (O_2908,N_22936,N_23823);
nor UO_2909 (O_2909,N_23985,N_23365);
nor UO_2910 (O_2910,N_24449,N_24512);
nor UO_2911 (O_2911,N_23374,N_24045);
and UO_2912 (O_2912,N_22984,N_24550);
xnor UO_2913 (O_2913,N_24405,N_24096);
nor UO_2914 (O_2914,N_22867,N_23755);
nor UO_2915 (O_2915,N_23169,N_24453);
and UO_2916 (O_2916,N_22709,N_24675);
nand UO_2917 (O_2917,N_23202,N_23900);
nand UO_2918 (O_2918,N_24720,N_22520);
nor UO_2919 (O_2919,N_22786,N_23572);
nor UO_2920 (O_2920,N_22716,N_24305);
or UO_2921 (O_2921,N_24928,N_24512);
nor UO_2922 (O_2922,N_22524,N_24005);
nand UO_2923 (O_2923,N_22624,N_24063);
nor UO_2924 (O_2924,N_22917,N_22800);
nand UO_2925 (O_2925,N_24099,N_22686);
nor UO_2926 (O_2926,N_24376,N_23685);
nor UO_2927 (O_2927,N_23074,N_24615);
or UO_2928 (O_2928,N_24417,N_23640);
or UO_2929 (O_2929,N_22512,N_24804);
nor UO_2930 (O_2930,N_24263,N_24928);
xnor UO_2931 (O_2931,N_24473,N_23344);
or UO_2932 (O_2932,N_23006,N_24712);
xnor UO_2933 (O_2933,N_22573,N_24353);
nand UO_2934 (O_2934,N_22721,N_22913);
nand UO_2935 (O_2935,N_24190,N_23172);
nor UO_2936 (O_2936,N_22511,N_22981);
or UO_2937 (O_2937,N_24541,N_24007);
nand UO_2938 (O_2938,N_23334,N_23328);
and UO_2939 (O_2939,N_22861,N_23281);
xor UO_2940 (O_2940,N_23088,N_22580);
xnor UO_2941 (O_2941,N_23658,N_24773);
or UO_2942 (O_2942,N_24484,N_23299);
or UO_2943 (O_2943,N_23607,N_24792);
xor UO_2944 (O_2944,N_22899,N_23184);
xor UO_2945 (O_2945,N_24098,N_22602);
xor UO_2946 (O_2946,N_24030,N_24450);
nor UO_2947 (O_2947,N_23230,N_24695);
nand UO_2948 (O_2948,N_22985,N_22880);
nor UO_2949 (O_2949,N_22738,N_24720);
nor UO_2950 (O_2950,N_24442,N_24893);
nor UO_2951 (O_2951,N_23120,N_22734);
xor UO_2952 (O_2952,N_23326,N_23687);
xnor UO_2953 (O_2953,N_24486,N_23647);
nand UO_2954 (O_2954,N_24100,N_23348);
nand UO_2955 (O_2955,N_23524,N_24632);
nand UO_2956 (O_2956,N_22852,N_23321);
and UO_2957 (O_2957,N_23429,N_24863);
nor UO_2958 (O_2958,N_23630,N_23814);
or UO_2959 (O_2959,N_22584,N_22755);
xor UO_2960 (O_2960,N_22635,N_23586);
nor UO_2961 (O_2961,N_23458,N_23153);
xor UO_2962 (O_2962,N_24920,N_24983);
or UO_2963 (O_2963,N_24571,N_24284);
xnor UO_2964 (O_2964,N_24771,N_24749);
nor UO_2965 (O_2965,N_24236,N_24551);
xor UO_2966 (O_2966,N_23511,N_23420);
nand UO_2967 (O_2967,N_24359,N_24538);
or UO_2968 (O_2968,N_24923,N_23364);
nand UO_2969 (O_2969,N_23566,N_23954);
xor UO_2970 (O_2970,N_23091,N_24496);
nand UO_2971 (O_2971,N_24575,N_23869);
xor UO_2972 (O_2972,N_24596,N_24585);
and UO_2973 (O_2973,N_23026,N_24787);
xor UO_2974 (O_2974,N_24936,N_23119);
nor UO_2975 (O_2975,N_22819,N_23542);
nand UO_2976 (O_2976,N_24146,N_24478);
xnor UO_2977 (O_2977,N_24516,N_24175);
and UO_2978 (O_2978,N_22644,N_23853);
nor UO_2979 (O_2979,N_24938,N_23528);
or UO_2980 (O_2980,N_22716,N_23328);
nand UO_2981 (O_2981,N_23017,N_24926);
or UO_2982 (O_2982,N_23521,N_23210);
nand UO_2983 (O_2983,N_24625,N_23444);
or UO_2984 (O_2984,N_22846,N_23647);
and UO_2985 (O_2985,N_23090,N_24447);
nand UO_2986 (O_2986,N_24448,N_23892);
xor UO_2987 (O_2987,N_23123,N_24867);
xnor UO_2988 (O_2988,N_23489,N_24968);
nand UO_2989 (O_2989,N_23062,N_22748);
xnor UO_2990 (O_2990,N_24546,N_23095);
or UO_2991 (O_2991,N_24118,N_24162);
nor UO_2992 (O_2992,N_23233,N_24838);
or UO_2993 (O_2993,N_23817,N_23884);
nand UO_2994 (O_2994,N_22738,N_24460);
or UO_2995 (O_2995,N_23697,N_23967);
and UO_2996 (O_2996,N_24566,N_24909);
and UO_2997 (O_2997,N_23170,N_22823);
nand UO_2998 (O_2998,N_23226,N_23199);
and UO_2999 (O_2999,N_23833,N_22691);
endmodule