module basic_1000_10000_1500_5_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_216,In_504);
or U1 (N_1,In_72,In_715);
nor U2 (N_2,In_171,In_344);
nor U3 (N_3,In_60,In_672);
nor U4 (N_4,In_142,In_986);
or U5 (N_5,In_104,In_463);
or U6 (N_6,In_961,In_567);
and U7 (N_7,In_134,In_212);
nand U8 (N_8,In_230,In_856);
or U9 (N_9,In_647,In_424);
nor U10 (N_10,In_107,In_288);
nor U11 (N_11,In_55,In_488);
or U12 (N_12,In_250,In_997);
and U13 (N_13,In_612,In_678);
and U14 (N_14,In_81,In_983);
and U15 (N_15,In_246,In_176);
nand U16 (N_16,In_234,In_347);
nor U17 (N_17,In_450,In_293);
and U18 (N_18,In_361,In_712);
nand U19 (N_19,In_823,In_659);
and U20 (N_20,In_272,In_987);
nor U21 (N_21,In_181,In_422);
nor U22 (N_22,In_337,In_137);
nor U23 (N_23,In_566,In_39);
and U24 (N_24,In_694,In_487);
xnor U25 (N_25,In_590,In_41);
xor U26 (N_26,In_928,In_313);
nor U27 (N_27,In_904,In_453);
nor U28 (N_28,In_906,In_756);
nor U29 (N_29,In_128,In_430);
xor U30 (N_30,In_839,In_535);
and U31 (N_31,In_692,In_820);
nand U32 (N_32,In_609,In_315);
nor U33 (N_33,In_243,In_218);
and U34 (N_34,In_975,In_27);
or U35 (N_35,In_653,In_934);
nor U36 (N_36,In_335,In_263);
or U37 (N_37,In_338,In_911);
and U38 (N_38,In_570,In_664);
nand U39 (N_39,In_371,In_561);
nand U40 (N_40,In_539,In_891);
and U41 (N_41,In_318,In_482);
xor U42 (N_42,In_403,In_22);
or U43 (N_43,In_349,In_679);
nand U44 (N_44,In_989,In_931);
or U45 (N_45,In_866,In_873);
or U46 (N_46,In_362,In_600);
and U47 (N_47,In_784,In_491);
or U48 (N_48,In_620,In_919);
and U49 (N_49,In_256,In_173);
nand U50 (N_50,In_690,In_435);
and U51 (N_51,In_348,In_414);
nor U52 (N_52,In_733,In_200);
nand U53 (N_53,In_990,In_373);
nor U54 (N_54,In_448,In_201);
or U55 (N_55,In_656,In_381);
nor U56 (N_56,In_155,In_452);
or U57 (N_57,In_193,In_202);
nor U58 (N_58,In_747,In_816);
nor U59 (N_59,In_550,In_970);
nor U60 (N_60,In_75,In_386);
nand U61 (N_61,In_459,In_251);
or U62 (N_62,In_164,In_541);
and U63 (N_63,In_133,In_864);
and U64 (N_64,In_749,In_761);
or U65 (N_65,In_291,In_506);
nand U66 (N_66,In_812,In_196);
and U67 (N_67,In_56,In_358);
nand U68 (N_68,In_262,In_392);
and U69 (N_69,In_775,In_227);
and U70 (N_70,In_443,In_462);
and U71 (N_71,In_937,In_648);
or U72 (N_72,In_545,In_966);
nand U73 (N_73,In_458,In_411);
nand U74 (N_74,In_180,In_169);
and U75 (N_75,In_682,In_351);
or U76 (N_76,In_2,In_851);
nor U77 (N_77,In_350,In_404);
nand U78 (N_78,In_905,In_719);
nor U79 (N_79,In_456,In_611);
nor U80 (N_80,In_252,In_902);
nand U81 (N_81,In_255,In_86);
nand U82 (N_82,In_45,In_304);
or U83 (N_83,In_689,In_190);
or U84 (N_84,In_325,In_810);
xnor U85 (N_85,In_857,In_298);
nand U86 (N_86,In_330,In_862);
nor U87 (N_87,In_714,In_881);
nand U88 (N_88,In_575,In_863);
nor U89 (N_89,In_882,In_825);
or U90 (N_90,In_215,In_633);
nand U91 (N_91,In_644,In_25);
and U92 (N_92,In_356,In_375);
nand U93 (N_93,In_743,In_923);
or U94 (N_94,In_419,In_476);
and U95 (N_95,In_853,In_593);
and U96 (N_96,In_223,In_716);
nand U97 (N_97,In_945,In_523);
and U98 (N_98,In_793,In_898);
or U99 (N_99,In_768,In_62);
or U100 (N_100,In_57,In_241);
nand U101 (N_101,In_493,In_13);
nand U102 (N_102,In_108,In_584);
nor U103 (N_103,In_106,In_595);
or U104 (N_104,In_401,In_811);
or U105 (N_105,In_936,In_306);
or U106 (N_106,In_82,In_179);
or U107 (N_107,In_977,In_726);
and U108 (N_108,In_292,In_307);
xnor U109 (N_109,In_354,In_433);
nand U110 (N_110,In_929,In_310);
and U111 (N_111,In_260,In_80);
nor U112 (N_112,In_870,In_867);
nor U113 (N_113,In_237,In_290);
nor U114 (N_114,In_925,In_814);
or U115 (N_115,In_554,In_996);
and U116 (N_116,In_529,In_16);
or U117 (N_117,In_489,In_877);
or U118 (N_118,In_739,In_296);
nor U119 (N_119,In_666,In_817);
nand U120 (N_120,In_168,In_156);
nand U121 (N_121,In_832,In_229);
nor U122 (N_122,In_829,In_469);
or U123 (N_123,In_117,In_380);
or U124 (N_124,In_819,In_159);
and U125 (N_125,In_577,In_467);
nor U126 (N_126,In_398,In_445);
nor U127 (N_127,In_594,In_933);
xor U128 (N_128,In_167,In_324);
xor U129 (N_129,In_789,In_652);
or U130 (N_130,In_622,In_267);
nand U131 (N_131,In_157,In_172);
or U132 (N_132,In_175,In_264);
and U133 (N_133,In_681,In_160);
nor U134 (N_134,In_855,In_591);
nor U135 (N_135,In_572,In_831);
and U136 (N_136,In_395,In_47);
nor U137 (N_137,In_843,In_6);
xor U138 (N_138,In_568,In_367);
or U139 (N_139,In_532,In_943);
and U140 (N_140,In_94,In_626);
nand U141 (N_141,In_518,In_231);
nand U142 (N_142,In_368,In_76);
or U143 (N_143,In_903,In_766);
nand U144 (N_144,In_14,In_40);
or U145 (N_145,In_492,In_511);
nand U146 (N_146,In_470,In_507);
and U147 (N_147,In_608,In_70);
and U148 (N_148,In_186,In_444);
and U149 (N_149,In_259,In_490);
nand U150 (N_150,In_198,In_702);
and U151 (N_151,In_299,In_346);
or U152 (N_152,In_979,In_822);
and U153 (N_153,In_885,In_317);
nand U154 (N_154,In_236,In_334);
and U155 (N_155,In_951,In_763);
and U156 (N_156,In_625,In_432);
and U157 (N_157,In_782,In_725);
nand U158 (N_158,In_161,In_24);
nand U159 (N_159,In_43,In_895);
and U160 (N_160,In_824,In_418);
nand U161 (N_161,In_676,In_805);
or U162 (N_162,In_145,In_558);
nand U163 (N_163,In_606,In_195);
or U164 (N_164,In_191,In_760);
nand U165 (N_165,In_68,In_232);
xnor U166 (N_166,In_302,In_438);
or U167 (N_167,In_410,In_520);
nor U168 (N_168,In_828,In_607);
nand U169 (N_169,In_124,In_872);
or U170 (N_170,In_571,In_93);
nand U171 (N_171,In_602,In_637);
xnor U172 (N_172,In_826,In_883);
nor U173 (N_173,In_240,In_205);
and U174 (N_174,In_278,In_846);
nand U175 (N_175,In_974,In_589);
or U176 (N_176,In_804,In_50);
and U177 (N_177,In_484,In_616);
nand U178 (N_178,In_412,In_673);
and U179 (N_179,In_203,In_147);
or U180 (N_180,In_918,In_224);
nand U181 (N_181,In_665,In_512);
nand U182 (N_182,In_222,In_848);
or U183 (N_183,In_818,In_509);
nand U184 (N_184,In_51,In_603);
nor U185 (N_185,In_295,In_728);
and U186 (N_186,In_700,In_294);
and U187 (N_187,In_954,In_79);
nand U188 (N_188,In_377,In_695);
nor U189 (N_189,In_683,In_274);
nor U190 (N_190,In_868,In_900);
and U191 (N_191,In_64,In_384);
nor U192 (N_192,In_516,In_757);
or U193 (N_193,In_613,In_12);
nand U194 (N_194,In_980,In_396);
xnor U195 (N_195,In_960,In_809);
or U196 (N_196,In_420,In_140);
and U197 (N_197,In_429,In_573);
and U198 (N_198,In_208,In_661);
and U199 (N_199,In_991,In_604);
and U200 (N_200,In_786,In_130);
or U201 (N_201,In_751,In_752);
and U202 (N_202,In_618,In_799);
or U203 (N_203,In_184,In_235);
nor U204 (N_204,In_519,In_807);
or U205 (N_205,In_115,In_649);
nand U206 (N_206,In_408,In_699);
nand U207 (N_207,In_813,In_99);
xor U208 (N_208,In_220,In_907);
or U209 (N_209,In_769,In_788);
xor U210 (N_210,In_889,In_771);
or U211 (N_211,In_632,In_671);
and U212 (N_212,In_780,In_153);
nor U213 (N_213,In_527,In_54);
or U214 (N_214,In_3,In_29);
nor U215 (N_215,In_783,In_720);
xor U216 (N_216,In_580,In_559);
nor U217 (N_217,In_913,In_485);
nor U218 (N_218,In_38,In_998);
nor U219 (N_219,In_283,In_400);
nand U220 (N_220,In_582,In_326);
or U221 (N_221,In_800,In_439);
nor U222 (N_222,In_583,In_724);
nor U223 (N_223,In_875,In_393);
xor U224 (N_224,In_275,In_765);
xor U225 (N_225,In_4,In_736);
nor U226 (N_226,In_266,In_333);
or U227 (N_227,In_538,In_314);
or U228 (N_228,In_691,In_74);
nor U229 (N_229,In_887,In_586);
and U230 (N_230,In_976,In_854);
nor U231 (N_231,In_697,In_947);
xor U232 (N_232,In_792,In_31);
xor U233 (N_233,In_286,In_20);
nor U234 (N_234,In_741,In_935);
nand U235 (N_235,In_847,In_217);
nand U236 (N_236,In_34,In_63);
and U237 (N_237,In_98,In_655);
nor U238 (N_238,In_542,In_734);
or U239 (N_239,In_442,In_667);
and U240 (N_240,In_131,In_543);
nand U241 (N_241,In_233,In_119);
nor U242 (N_242,In_930,In_61);
xnor U243 (N_243,In_537,In_546);
xnor U244 (N_244,In_711,In_364);
nand U245 (N_245,In_84,In_921);
nand U246 (N_246,In_879,In_845);
or U247 (N_247,In_674,In_696);
nor U248 (N_248,In_801,In_103);
nand U249 (N_249,In_745,In_908);
nor U250 (N_250,In_343,In_440);
nand U251 (N_251,In_552,In_964);
nor U252 (N_252,In_920,In_750);
nand U253 (N_253,In_588,In_758);
and U254 (N_254,In_383,In_97);
and U255 (N_255,In_513,In_526);
nand U256 (N_256,In_312,In_709);
nand U257 (N_257,In_496,In_623);
nor U258 (N_258,In_844,In_922);
nand U259 (N_259,In_457,In_194);
or U260 (N_260,In_698,In_610);
nor U261 (N_261,In_717,In_636);
and U262 (N_262,In_985,In_858);
xor U263 (N_263,In_394,In_564);
or U264 (N_264,In_949,In_406);
and U265 (N_265,In_576,In_654);
or U266 (N_266,In_44,In_495);
or U267 (N_267,In_796,In_451);
nand U268 (N_268,In_833,In_287);
xnor U269 (N_269,In_87,In_503);
nand U270 (N_270,In_185,In_525);
and U271 (N_271,In_423,In_65);
or U272 (N_272,In_500,In_806);
and U273 (N_273,In_138,In_556);
and U274 (N_274,In_37,In_308);
nor U275 (N_275,In_912,In_226);
nor U276 (N_276,In_309,In_981);
nand U277 (N_277,In_994,In_468);
or U278 (N_278,In_982,In_365);
and U279 (N_279,In_409,In_953);
nor U280 (N_280,In_100,In_701);
nor U281 (N_281,In_66,In_340);
and U282 (N_282,In_407,In_869);
and U283 (N_283,In_165,In_643);
nand U284 (N_284,In_281,In_28);
and U285 (N_285,In_239,In_940);
or U286 (N_286,In_927,In_723);
or U287 (N_287,In_650,In_0);
xor U288 (N_288,In_269,In_821);
nand U289 (N_289,In_148,In_102);
xnor U290 (N_290,In_533,In_544);
and U291 (N_291,In_101,In_662);
nor U292 (N_292,In_472,In_790);
nor U293 (N_293,In_515,In_827);
nand U294 (N_294,In_69,In_36);
and U295 (N_295,In_548,In_53);
and U296 (N_296,In_727,In_950);
nor U297 (N_297,In_305,In_841);
nor U298 (N_298,In_89,In_737);
xnor U299 (N_299,In_668,In_563);
xor U300 (N_300,In_268,In_26);
or U301 (N_301,In_316,In_703);
nand U302 (N_302,In_860,In_635);
nor U303 (N_303,In_273,In_17);
xor U304 (N_304,In_686,In_547);
or U305 (N_305,In_878,In_261);
or U306 (N_306,In_791,In_58);
and U307 (N_307,In_454,In_23);
or U308 (N_308,In_886,In_178);
and U309 (N_309,In_342,In_917);
nand U310 (N_310,In_551,In_963);
nor U311 (N_311,In_969,In_15);
xnor U312 (N_312,In_328,In_242);
nand U313 (N_313,In_182,In_188);
nand U314 (N_314,In_522,In_596);
or U315 (N_315,In_416,In_540);
nand U316 (N_316,In_721,In_893);
xor U317 (N_317,In_798,In_968);
nor U318 (N_318,In_640,In_83);
nor U319 (N_319,In_280,In_957);
and U320 (N_320,In_118,In_289);
nand U321 (N_321,In_587,In_494);
and U322 (N_322,In_865,In_376);
or U323 (N_323,In_499,In_932);
and U324 (N_324,In_238,In_78);
nor U325 (N_325,In_151,In_105);
and U326 (N_326,In_221,In_311);
nand U327 (N_327,In_748,In_258);
nand U328 (N_328,In_122,In_219);
nand U329 (N_329,In_508,In_713);
or U330 (N_330,In_486,In_327);
or U331 (N_331,In_651,In_42);
nor U332 (N_332,In_213,In_871);
nand U333 (N_333,In_803,In_9);
and U334 (N_334,In_329,In_189);
xor U335 (N_335,In_303,In_323);
xnor U336 (N_336,In_471,In_955);
nand U337 (N_337,In_874,In_387);
xnor U338 (N_338,In_385,In_759);
nor U339 (N_339,In_849,In_685);
nor U340 (N_340,In_764,In_627);
or U341 (N_341,In_111,In_658);
and U342 (N_342,In_706,In_5);
and U343 (N_343,In_211,In_815);
xor U344 (N_344,In_92,In_352);
and U345 (N_345,In_112,In_840);
nor U346 (N_346,In_524,In_753);
nand U347 (N_347,In_777,In_332);
or U348 (N_348,In_355,In_152);
or U349 (N_349,In_248,In_425);
nor U350 (N_350,In_560,In_531);
nand U351 (N_351,In_732,In_279);
and U352 (N_352,In_120,In_146);
and U353 (N_353,In_958,In_730);
nor U354 (N_354,In_770,In_154);
nand U355 (N_355,In_46,In_253);
nor U356 (N_356,In_884,In_892);
nand U357 (N_357,In_621,In_132);
or U358 (N_358,In_619,In_708);
nand U359 (N_359,In_477,In_129);
nor U360 (N_360,In_773,In_740);
nand U361 (N_361,In_464,In_399);
nand U362 (N_362,In_630,In_245);
nor U363 (N_363,In_30,In_710);
and U364 (N_364,In_746,In_437);
or U365 (N_365,In_319,In_984);
and U366 (N_366,In_441,In_669);
nand U367 (N_367,In_776,In_924);
nor U368 (N_368,In_534,In_956);
or U369 (N_369,In_48,In_510);
or U370 (N_370,In_521,In_722);
nand U371 (N_371,In_225,In_687);
or U372 (N_372,In_378,In_52);
or U373 (N_373,In_341,In_677);
nand U374 (N_374,In_562,In_139);
xor U375 (N_375,In_372,In_121);
or U376 (N_376,In_718,In_113);
and U377 (N_377,In_729,In_939);
nor U378 (N_378,In_85,In_73);
and U379 (N_379,In_434,In_428);
nor U380 (N_380,In_896,In_207);
or U381 (N_381,In_938,In_498);
nand U382 (N_382,In_11,In_474);
or U383 (N_383,In_599,In_914);
nand U384 (N_384,In_565,In_941);
nor U385 (N_385,In_501,In_282);
nor U386 (N_386,In_461,In_466);
nor U387 (N_387,In_794,In_894);
or U388 (N_388,In_549,In_553);
nor U389 (N_389,In_370,In_842);
and U390 (N_390,In_8,In_754);
nor U391 (N_391,In_71,In_123);
or U392 (N_392,In_973,In_369);
nor U393 (N_393,In_95,In_21);
and U394 (N_394,In_688,In_774);
and U395 (N_395,In_483,In_639);
nand U396 (N_396,In_645,In_336);
nand U397 (N_397,In_779,In_177);
nand U398 (N_398,In_767,In_447);
nand U399 (N_399,In_88,In_465);
xor U400 (N_400,In_942,In_276);
xnor U401 (N_401,In_397,In_642);
or U402 (N_402,In_693,In_897);
nand U403 (N_403,In_802,In_388);
and U404 (N_404,In_127,In_379);
nor U405 (N_405,In_90,In_244);
or U406 (N_406,In_993,In_926);
nand U407 (N_407,In_852,In_528);
and U408 (N_408,In_557,In_366);
and U409 (N_409,In_624,In_836);
xnor U410 (N_410,In_143,In_657);
or U411 (N_411,In_967,In_163);
or U412 (N_412,In_7,In_663);
or U413 (N_413,In_944,In_210);
nor U414 (N_414,In_808,In_995);
nor U415 (N_415,In_284,In_988);
nor U416 (N_416,In_876,In_345);
or U417 (N_417,In_285,In_838);
nand U418 (N_418,In_992,In_436);
xnor U419 (N_419,In_320,In_402);
nor U420 (N_420,In_675,In_257);
nor U421 (N_421,In_135,In_174);
nand U422 (N_422,In_578,In_670);
xor U423 (N_423,In_959,In_778);
or U424 (N_424,In_166,In_859);
nor U425 (N_425,In_965,In_597);
or U426 (N_426,In_204,In_136);
nand U427 (N_427,In_405,In_359);
or U428 (N_428,In_144,In_480);
or U429 (N_429,In_880,In_254);
or U430 (N_430,In_49,In_742);
nor U431 (N_431,In_427,In_772);
xor U432 (N_432,In_149,In_382);
nor U433 (N_433,In_481,In_514);
and U434 (N_434,In_426,In_249);
nand U435 (N_435,In_629,In_910);
and U436 (N_436,In_363,In_192);
or U437 (N_437,In_555,In_91);
or U438 (N_438,In_787,In_158);
or U439 (N_439,In_971,In_150);
or U440 (N_440,In_605,In_187);
or U441 (N_441,In_888,In_449);
xor U442 (N_442,In_18,In_321);
or U443 (N_443,In_530,In_141);
or U444 (N_444,In_415,In_646);
nand U445 (N_445,In_199,In_77);
nand U446 (N_446,In_948,In_762);
and U447 (N_447,In_301,In_277);
and U448 (N_448,In_478,In_109);
or U449 (N_449,In_899,In_585);
and U450 (N_450,In_634,In_265);
or U451 (N_451,In_614,In_850);
nand U452 (N_452,In_628,In_660);
nor U453 (N_453,In_781,In_617);
or U454 (N_454,In_455,In_389);
nor U455 (N_455,In_446,In_116);
nand U456 (N_456,In_579,In_574);
nand U457 (N_457,In_126,In_125);
or U458 (N_458,In_497,In_705);
or U459 (N_459,In_901,In_228);
nor U460 (N_460,In_598,In_505);
nor U461 (N_461,In_183,In_374);
nand U462 (N_462,In_19,In_707);
nand U463 (N_463,In_952,In_360);
and U464 (N_464,In_797,In_431);
nand U465 (N_465,In_391,In_322);
nor U466 (N_466,In_502,In_536);
or U467 (N_467,In_738,In_962);
or U468 (N_468,In_297,In_735);
xor U469 (N_469,In_353,In_680);
nor U470 (N_470,In_909,In_413);
nor U471 (N_471,In_641,In_247);
nand U472 (N_472,In_460,In_10);
and U473 (N_473,In_785,In_339);
or U474 (N_474,In_592,In_390);
and U475 (N_475,In_300,In_331);
nand U476 (N_476,In_206,In_33);
nor U477 (N_477,In_834,In_110);
and U478 (N_478,In_162,In_35);
and U479 (N_479,In_114,In_473);
or U480 (N_480,In_357,In_615);
nor U481 (N_481,In_830,In_209);
nand U482 (N_482,In_601,In_421);
nor U483 (N_483,In_631,In_744);
nor U484 (N_484,In_214,In_517);
or U485 (N_485,In_67,In_837);
or U486 (N_486,In_96,In_271);
or U487 (N_487,In_569,In_197);
nor U488 (N_488,In_270,In_1);
or U489 (N_489,In_684,In_972);
or U490 (N_490,In_861,In_581);
nor U491 (N_491,In_479,In_835);
nor U492 (N_492,In_638,In_755);
or U493 (N_493,In_417,In_475);
and U494 (N_494,In_704,In_916);
nor U495 (N_495,In_978,In_795);
or U496 (N_496,In_915,In_59);
and U497 (N_497,In_731,In_170);
and U498 (N_498,In_890,In_32);
or U499 (N_499,In_946,In_999);
or U500 (N_500,In_138,In_85);
and U501 (N_501,In_243,In_943);
and U502 (N_502,In_742,In_430);
or U503 (N_503,In_47,In_625);
nand U504 (N_504,In_315,In_88);
nor U505 (N_505,In_150,In_935);
or U506 (N_506,In_177,In_240);
nor U507 (N_507,In_893,In_217);
or U508 (N_508,In_341,In_680);
nand U509 (N_509,In_169,In_552);
or U510 (N_510,In_568,In_874);
xor U511 (N_511,In_191,In_310);
or U512 (N_512,In_43,In_527);
nand U513 (N_513,In_278,In_467);
or U514 (N_514,In_401,In_106);
or U515 (N_515,In_445,In_309);
and U516 (N_516,In_9,In_191);
nor U517 (N_517,In_400,In_731);
nand U518 (N_518,In_974,In_519);
and U519 (N_519,In_422,In_826);
and U520 (N_520,In_296,In_501);
or U521 (N_521,In_214,In_964);
or U522 (N_522,In_914,In_43);
nand U523 (N_523,In_578,In_459);
or U524 (N_524,In_923,In_489);
nor U525 (N_525,In_3,In_756);
xor U526 (N_526,In_30,In_307);
nand U527 (N_527,In_180,In_3);
or U528 (N_528,In_860,In_916);
or U529 (N_529,In_605,In_214);
or U530 (N_530,In_412,In_494);
or U531 (N_531,In_238,In_411);
or U532 (N_532,In_426,In_694);
and U533 (N_533,In_986,In_894);
and U534 (N_534,In_289,In_246);
and U535 (N_535,In_335,In_956);
nor U536 (N_536,In_709,In_657);
xnor U537 (N_537,In_235,In_341);
or U538 (N_538,In_78,In_231);
or U539 (N_539,In_957,In_888);
or U540 (N_540,In_190,In_955);
nor U541 (N_541,In_182,In_220);
or U542 (N_542,In_806,In_176);
or U543 (N_543,In_286,In_781);
nand U544 (N_544,In_883,In_364);
or U545 (N_545,In_27,In_537);
and U546 (N_546,In_865,In_972);
nor U547 (N_547,In_107,In_513);
nand U548 (N_548,In_99,In_142);
nand U549 (N_549,In_734,In_781);
nor U550 (N_550,In_352,In_541);
and U551 (N_551,In_717,In_332);
or U552 (N_552,In_740,In_952);
or U553 (N_553,In_598,In_449);
xnor U554 (N_554,In_3,In_817);
xor U555 (N_555,In_498,In_673);
or U556 (N_556,In_174,In_295);
nor U557 (N_557,In_720,In_828);
nand U558 (N_558,In_725,In_919);
xor U559 (N_559,In_902,In_508);
or U560 (N_560,In_948,In_922);
nor U561 (N_561,In_644,In_326);
nand U562 (N_562,In_408,In_576);
nor U563 (N_563,In_444,In_293);
xnor U564 (N_564,In_748,In_839);
or U565 (N_565,In_543,In_975);
or U566 (N_566,In_295,In_419);
xnor U567 (N_567,In_541,In_513);
or U568 (N_568,In_478,In_154);
nor U569 (N_569,In_934,In_834);
or U570 (N_570,In_66,In_16);
nor U571 (N_571,In_436,In_967);
or U572 (N_572,In_642,In_843);
nand U573 (N_573,In_74,In_246);
and U574 (N_574,In_73,In_577);
and U575 (N_575,In_789,In_267);
xor U576 (N_576,In_894,In_506);
or U577 (N_577,In_431,In_642);
nor U578 (N_578,In_927,In_21);
nor U579 (N_579,In_190,In_686);
and U580 (N_580,In_322,In_919);
or U581 (N_581,In_831,In_786);
or U582 (N_582,In_137,In_876);
nor U583 (N_583,In_857,In_149);
nor U584 (N_584,In_924,In_933);
nand U585 (N_585,In_718,In_733);
nand U586 (N_586,In_116,In_414);
nor U587 (N_587,In_876,In_524);
nand U588 (N_588,In_573,In_400);
or U589 (N_589,In_155,In_856);
and U590 (N_590,In_319,In_510);
or U591 (N_591,In_334,In_980);
or U592 (N_592,In_817,In_663);
and U593 (N_593,In_679,In_573);
or U594 (N_594,In_140,In_421);
and U595 (N_595,In_631,In_972);
nor U596 (N_596,In_333,In_817);
nand U597 (N_597,In_959,In_22);
nand U598 (N_598,In_870,In_583);
xnor U599 (N_599,In_87,In_873);
nand U600 (N_600,In_501,In_408);
and U601 (N_601,In_395,In_926);
nand U602 (N_602,In_309,In_641);
and U603 (N_603,In_49,In_331);
nand U604 (N_604,In_647,In_284);
xnor U605 (N_605,In_157,In_439);
nand U606 (N_606,In_852,In_954);
or U607 (N_607,In_308,In_85);
or U608 (N_608,In_667,In_697);
nor U609 (N_609,In_937,In_636);
or U610 (N_610,In_396,In_710);
nor U611 (N_611,In_637,In_558);
nand U612 (N_612,In_585,In_40);
or U613 (N_613,In_751,In_152);
nor U614 (N_614,In_342,In_395);
nor U615 (N_615,In_783,In_499);
nor U616 (N_616,In_808,In_835);
or U617 (N_617,In_907,In_784);
nor U618 (N_618,In_610,In_822);
nor U619 (N_619,In_558,In_616);
or U620 (N_620,In_887,In_668);
or U621 (N_621,In_279,In_544);
and U622 (N_622,In_662,In_307);
or U623 (N_623,In_61,In_88);
or U624 (N_624,In_772,In_801);
nor U625 (N_625,In_451,In_250);
or U626 (N_626,In_207,In_246);
or U627 (N_627,In_212,In_788);
and U628 (N_628,In_994,In_83);
and U629 (N_629,In_835,In_169);
nand U630 (N_630,In_59,In_80);
nor U631 (N_631,In_754,In_381);
and U632 (N_632,In_760,In_223);
nor U633 (N_633,In_728,In_843);
and U634 (N_634,In_54,In_871);
nand U635 (N_635,In_6,In_417);
and U636 (N_636,In_387,In_982);
and U637 (N_637,In_182,In_680);
nand U638 (N_638,In_823,In_676);
or U639 (N_639,In_434,In_852);
nand U640 (N_640,In_276,In_580);
and U641 (N_641,In_626,In_476);
nand U642 (N_642,In_569,In_386);
and U643 (N_643,In_537,In_343);
nand U644 (N_644,In_753,In_599);
nand U645 (N_645,In_580,In_756);
xnor U646 (N_646,In_573,In_735);
xnor U647 (N_647,In_925,In_71);
nor U648 (N_648,In_988,In_614);
xnor U649 (N_649,In_710,In_257);
or U650 (N_650,In_925,In_144);
and U651 (N_651,In_734,In_391);
xnor U652 (N_652,In_486,In_194);
nor U653 (N_653,In_552,In_793);
xnor U654 (N_654,In_534,In_319);
nand U655 (N_655,In_736,In_615);
or U656 (N_656,In_554,In_983);
or U657 (N_657,In_792,In_532);
xor U658 (N_658,In_244,In_137);
nor U659 (N_659,In_987,In_420);
or U660 (N_660,In_375,In_621);
nand U661 (N_661,In_760,In_639);
or U662 (N_662,In_699,In_875);
or U663 (N_663,In_540,In_939);
xor U664 (N_664,In_302,In_416);
or U665 (N_665,In_914,In_782);
xor U666 (N_666,In_578,In_699);
nor U667 (N_667,In_464,In_140);
or U668 (N_668,In_966,In_299);
xnor U669 (N_669,In_700,In_27);
nor U670 (N_670,In_55,In_429);
nor U671 (N_671,In_776,In_74);
nor U672 (N_672,In_619,In_881);
nor U673 (N_673,In_473,In_720);
xnor U674 (N_674,In_212,In_666);
and U675 (N_675,In_814,In_811);
nand U676 (N_676,In_699,In_500);
xor U677 (N_677,In_715,In_634);
or U678 (N_678,In_646,In_951);
or U679 (N_679,In_291,In_13);
nand U680 (N_680,In_83,In_669);
or U681 (N_681,In_163,In_835);
nand U682 (N_682,In_237,In_461);
nor U683 (N_683,In_304,In_479);
or U684 (N_684,In_856,In_562);
or U685 (N_685,In_862,In_746);
nand U686 (N_686,In_141,In_83);
nor U687 (N_687,In_577,In_834);
nor U688 (N_688,In_53,In_457);
nor U689 (N_689,In_410,In_229);
and U690 (N_690,In_160,In_780);
nand U691 (N_691,In_442,In_84);
nand U692 (N_692,In_716,In_553);
nand U693 (N_693,In_756,In_864);
or U694 (N_694,In_768,In_589);
or U695 (N_695,In_777,In_742);
and U696 (N_696,In_367,In_718);
nor U697 (N_697,In_456,In_739);
and U698 (N_698,In_308,In_816);
nand U699 (N_699,In_828,In_745);
nand U700 (N_700,In_274,In_733);
nor U701 (N_701,In_857,In_513);
nand U702 (N_702,In_764,In_631);
nand U703 (N_703,In_588,In_455);
nand U704 (N_704,In_913,In_840);
nand U705 (N_705,In_55,In_746);
or U706 (N_706,In_805,In_706);
nand U707 (N_707,In_69,In_177);
nand U708 (N_708,In_544,In_488);
nor U709 (N_709,In_139,In_763);
nor U710 (N_710,In_346,In_248);
or U711 (N_711,In_819,In_534);
nor U712 (N_712,In_404,In_203);
or U713 (N_713,In_587,In_84);
and U714 (N_714,In_104,In_474);
or U715 (N_715,In_819,In_631);
or U716 (N_716,In_214,In_469);
and U717 (N_717,In_125,In_418);
nand U718 (N_718,In_620,In_520);
nand U719 (N_719,In_178,In_907);
or U720 (N_720,In_584,In_517);
or U721 (N_721,In_684,In_815);
nor U722 (N_722,In_848,In_962);
and U723 (N_723,In_784,In_857);
or U724 (N_724,In_299,In_26);
and U725 (N_725,In_330,In_469);
nor U726 (N_726,In_350,In_742);
nand U727 (N_727,In_854,In_741);
and U728 (N_728,In_353,In_876);
nor U729 (N_729,In_394,In_740);
nor U730 (N_730,In_425,In_156);
and U731 (N_731,In_77,In_529);
xnor U732 (N_732,In_667,In_999);
or U733 (N_733,In_780,In_918);
or U734 (N_734,In_21,In_972);
nor U735 (N_735,In_830,In_51);
and U736 (N_736,In_377,In_474);
nor U737 (N_737,In_548,In_238);
and U738 (N_738,In_57,In_334);
or U739 (N_739,In_375,In_358);
or U740 (N_740,In_96,In_274);
xnor U741 (N_741,In_115,In_459);
xnor U742 (N_742,In_983,In_892);
xnor U743 (N_743,In_932,In_777);
or U744 (N_744,In_543,In_682);
nand U745 (N_745,In_878,In_212);
nand U746 (N_746,In_162,In_765);
nor U747 (N_747,In_285,In_561);
and U748 (N_748,In_979,In_133);
or U749 (N_749,In_405,In_384);
nor U750 (N_750,In_516,In_788);
nor U751 (N_751,In_604,In_287);
nand U752 (N_752,In_507,In_857);
and U753 (N_753,In_637,In_208);
nor U754 (N_754,In_529,In_571);
or U755 (N_755,In_678,In_695);
nand U756 (N_756,In_978,In_832);
nor U757 (N_757,In_65,In_777);
and U758 (N_758,In_822,In_282);
xor U759 (N_759,In_767,In_789);
nor U760 (N_760,In_639,In_146);
and U761 (N_761,In_632,In_23);
nor U762 (N_762,In_407,In_738);
nor U763 (N_763,In_989,In_241);
and U764 (N_764,In_498,In_58);
or U765 (N_765,In_18,In_53);
nor U766 (N_766,In_61,In_210);
xor U767 (N_767,In_227,In_340);
nor U768 (N_768,In_16,In_961);
nand U769 (N_769,In_251,In_448);
nor U770 (N_770,In_582,In_157);
and U771 (N_771,In_374,In_667);
and U772 (N_772,In_68,In_376);
nand U773 (N_773,In_304,In_822);
and U774 (N_774,In_88,In_666);
and U775 (N_775,In_835,In_753);
or U776 (N_776,In_936,In_380);
and U777 (N_777,In_982,In_306);
nand U778 (N_778,In_393,In_484);
or U779 (N_779,In_239,In_365);
nand U780 (N_780,In_75,In_615);
or U781 (N_781,In_588,In_93);
xnor U782 (N_782,In_88,In_929);
and U783 (N_783,In_580,In_187);
or U784 (N_784,In_638,In_336);
nand U785 (N_785,In_341,In_944);
nor U786 (N_786,In_692,In_637);
and U787 (N_787,In_837,In_780);
xnor U788 (N_788,In_352,In_256);
and U789 (N_789,In_144,In_79);
or U790 (N_790,In_113,In_956);
or U791 (N_791,In_29,In_713);
nor U792 (N_792,In_767,In_820);
or U793 (N_793,In_777,In_256);
xor U794 (N_794,In_452,In_131);
and U795 (N_795,In_804,In_957);
and U796 (N_796,In_899,In_446);
xor U797 (N_797,In_188,In_484);
or U798 (N_798,In_927,In_500);
xor U799 (N_799,In_904,In_723);
or U800 (N_800,In_524,In_934);
xnor U801 (N_801,In_942,In_241);
xor U802 (N_802,In_174,In_254);
xnor U803 (N_803,In_491,In_388);
xnor U804 (N_804,In_359,In_738);
and U805 (N_805,In_935,In_257);
or U806 (N_806,In_831,In_318);
and U807 (N_807,In_690,In_684);
nand U808 (N_808,In_693,In_47);
or U809 (N_809,In_61,In_871);
and U810 (N_810,In_33,In_15);
or U811 (N_811,In_852,In_407);
nor U812 (N_812,In_519,In_125);
xnor U813 (N_813,In_984,In_159);
and U814 (N_814,In_223,In_866);
and U815 (N_815,In_629,In_624);
nor U816 (N_816,In_374,In_782);
or U817 (N_817,In_131,In_164);
nor U818 (N_818,In_677,In_183);
or U819 (N_819,In_330,In_962);
xnor U820 (N_820,In_677,In_798);
nor U821 (N_821,In_419,In_281);
or U822 (N_822,In_146,In_983);
and U823 (N_823,In_453,In_94);
nand U824 (N_824,In_463,In_664);
nand U825 (N_825,In_753,In_994);
xnor U826 (N_826,In_182,In_439);
or U827 (N_827,In_419,In_713);
or U828 (N_828,In_273,In_959);
nor U829 (N_829,In_326,In_744);
or U830 (N_830,In_227,In_183);
nand U831 (N_831,In_264,In_93);
or U832 (N_832,In_40,In_801);
nand U833 (N_833,In_953,In_593);
nor U834 (N_834,In_25,In_921);
nor U835 (N_835,In_64,In_100);
nor U836 (N_836,In_870,In_657);
or U837 (N_837,In_639,In_524);
and U838 (N_838,In_125,In_249);
xor U839 (N_839,In_417,In_496);
and U840 (N_840,In_293,In_566);
xnor U841 (N_841,In_262,In_890);
nor U842 (N_842,In_710,In_293);
or U843 (N_843,In_380,In_922);
nand U844 (N_844,In_94,In_687);
or U845 (N_845,In_189,In_878);
nor U846 (N_846,In_474,In_613);
xnor U847 (N_847,In_378,In_322);
and U848 (N_848,In_317,In_987);
and U849 (N_849,In_188,In_525);
and U850 (N_850,In_64,In_402);
or U851 (N_851,In_451,In_286);
and U852 (N_852,In_369,In_87);
and U853 (N_853,In_162,In_540);
and U854 (N_854,In_872,In_878);
nand U855 (N_855,In_129,In_968);
nor U856 (N_856,In_87,In_885);
or U857 (N_857,In_240,In_738);
nor U858 (N_858,In_629,In_772);
or U859 (N_859,In_24,In_15);
and U860 (N_860,In_746,In_111);
xor U861 (N_861,In_570,In_39);
nand U862 (N_862,In_924,In_436);
xnor U863 (N_863,In_788,In_223);
nor U864 (N_864,In_957,In_314);
nor U865 (N_865,In_657,In_633);
nor U866 (N_866,In_213,In_455);
nor U867 (N_867,In_538,In_523);
nor U868 (N_868,In_859,In_18);
nand U869 (N_869,In_985,In_300);
and U870 (N_870,In_581,In_566);
nand U871 (N_871,In_302,In_665);
and U872 (N_872,In_890,In_27);
nor U873 (N_873,In_693,In_35);
nand U874 (N_874,In_69,In_647);
xnor U875 (N_875,In_723,In_45);
nand U876 (N_876,In_318,In_818);
or U877 (N_877,In_385,In_290);
nand U878 (N_878,In_294,In_980);
or U879 (N_879,In_970,In_986);
nor U880 (N_880,In_988,In_864);
nand U881 (N_881,In_152,In_547);
and U882 (N_882,In_322,In_194);
xnor U883 (N_883,In_79,In_867);
or U884 (N_884,In_661,In_780);
nor U885 (N_885,In_865,In_963);
and U886 (N_886,In_847,In_457);
and U887 (N_887,In_186,In_112);
nand U888 (N_888,In_4,In_149);
xor U889 (N_889,In_23,In_481);
or U890 (N_890,In_209,In_441);
nor U891 (N_891,In_950,In_236);
nand U892 (N_892,In_246,In_657);
nor U893 (N_893,In_83,In_982);
nor U894 (N_894,In_384,In_83);
or U895 (N_895,In_246,In_156);
and U896 (N_896,In_760,In_20);
or U897 (N_897,In_436,In_219);
or U898 (N_898,In_526,In_254);
xnor U899 (N_899,In_776,In_17);
nor U900 (N_900,In_386,In_697);
nand U901 (N_901,In_907,In_158);
nand U902 (N_902,In_953,In_783);
xnor U903 (N_903,In_738,In_752);
nor U904 (N_904,In_357,In_933);
nor U905 (N_905,In_953,In_978);
and U906 (N_906,In_568,In_801);
nor U907 (N_907,In_421,In_89);
and U908 (N_908,In_28,In_978);
nor U909 (N_909,In_390,In_508);
and U910 (N_910,In_957,In_435);
nor U911 (N_911,In_959,In_650);
xor U912 (N_912,In_614,In_69);
nand U913 (N_913,In_658,In_875);
xor U914 (N_914,In_675,In_774);
or U915 (N_915,In_753,In_149);
or U916 (N_916,In_509,In_524);
nand U917 (N_917,In_747,In_369);
or U918 (N_918,In_386,In_538);
nand U919 (N_919,In_513,In_670);
and U920 (N_920,In_206,In_929);
or U921 (N_921,In_904,In_202);
nand U922 (N_922,In_756,In_985);
xnor U923 (N_923,In_96,In_866);
nand U924 (N_924,In_717,In_683);
xnor U925 (N_925,In_977,In_817);
nand U926 (N_926,In_717,In_749);
and U927 (N_927,In_521,In_162);
xnor U928 (N_928,In_290,In_392);
or U929 (N_929,In_479,In_363);
nor U930 (N_930,In_972,In_628);
nand U931 (N_931,In_747,In_859);
or U932 (N_932,In_277,In_823);
or U933 (N_933,In_715,In_223);
nand U934 (N_934,In_590,In_303);
or U935 (N_935,In_17,In_267);
or U936 (N_936,In_617,In_508);
and U937 (N_937,In_447,In_156);
nor U938 (N_938,In_932,In_124);
and U939 (N_939,In_768,In_700);
xor U940 (N_940,In_605,In_794);
xnor U941 (N_941,In_259,In_943);
nand U942 (N_942,In_862,In_370);
and U943 (N_943,In_448,In_467);
nand U944 (N_944,In_932,In_155);
nand U945 (N_945,In_722,In_461);
or U946 (N_946,In_600,In_517);
or U947 (N_947,In_88,In_835);
nand U948 (N_948,In_952,In_347);
and U949 (N_949,In_700,In_436);
or U950 (N_950,In_704,In_720);
nand U951 (N_951,In_959,In_924);
or U952 (N_952,In_181,In_970);
nand U953 (N_953,In_452,In_12);
and U954 (N_954,In_200,In_875);
nand U955 (N_955,In_373,In_27);
nor U956 (N_956,In_585,In_788);
and U957 (N_957,In_62,In_72);
xor U958 (N_958,In_346,In_307);
and U959 (N_959,In_930,In_980);
or U960 (N_960,In_950,In_119);
and U961 (N_961,In_59,In_877);
nor U962 (N_962,In_445,In_648);
nor U963 (N_963,In_282,In_840);
nand U964 (N_964,In_371,In_313);
xnor U965 (N_965,In_377,In_241);
and U966 (N_966,In_440,In_122);
or U967 (N_967,In_37,In_927);
and U968 (N_968,In_477,In_795);
nor U969 (N_969,In_849,In_818);
or U970 (N_970,In_743,In_875);
nor U971 (N_971,In_695,In_637);
or U972 (N_972,In_976,In_279);
nor U973 (N_973,In_462,In_570);
xnor U974 (N_974,In_728,In_648);
nor U975 (N_975,In_420,In_688);
and U976 (N_976,In_966,In_186);
nand U977 (N_977,In_55,In_392);
and U978 (N_978,In_422,In_781);
or U979 (N_979,In_751,In_629);
nand U980 (N_980,In_828,In_723);
or U981 (N_981,In_209,In_158);
nor U982 (N_982,In_90,In_68);
or U983 (N_983,In_798,In_616);
and U984 (N_984,In_643,In_882);
and U985 (N_985,In_84,In_402);
nand U986 (N_986,In_888,In_255);
nand U987 (N_987,In_794,In_645);
and U988 (N_988,In_645,In_449);
or U989 (N_989,In_63,In_284);
and U990 (N_990,In_854,In_690);
and U991 (N_991,In_985,In_612);
or U992 (N_992,In_419,In_584);
and U993 (N_993,In_353,In_617);
or U994 (N_994,In_190,In_614);
and U995 (N_995,In_607,In_67);
or U996 (N_996,In_672,In_72);
xor U997 (N_997,In_313,In_882);
and U998 (N_998,In_727,In_80);
and U999 (N_999,In_454,In_62);
nor U1000 (N_1000,In_556,In_472);
or U1001 (N_1001,In_520,In_357);
nor U1002 (N_1002,In_202,In_853);
nor U1003 (N_1003,In_783,In_518);
and U1004 (N_1004,In_976,In_905);
nor U1005 (N_1005,In_633,In_167);
nor U1006 (N_1006,In_413,In_515);
and U1007 (N_1007,In_18,In_252);
or U1008 (N_1008,In_889,In_971);
nor U1009 (N_1009,In_651,In_848);
nand U1010 (N_1010,In_53,In_433);
nor U1011 (N_1011,In_137,In_832);
xnor U1012 (N_1012,In_92,In_720);
or U1013 (N_1013,In_758,In_55);
nand U1014 (N_1014,In_429,In_60);
nor U1015 (N_1015,In_205,In_42);
nor U1016 (N_1016,In_925,In_885);
nand U1017 (N_1017,In_703,In_189);
and U1018 (N_1018,In_140,In_231);
nand U1019 (N_1019,In_748,In_699);
xor U1020 (N_1020,In_999,In_45);
nand U1021 (N_1021,In_432,In_352);
nor U1022 (N_1022,In_179,In_529);
and U1023 (N_1023,In_916,In_598);
nand U1024 (N_1024,In_282,In_21);
and U1025 (N_1025,In_818,In_254);
and U1026 (N_1026,In_105,In_245);
xor U1027 (N_1027,In_512,In_235);
nand U1028 (N_1028,In_852,In_854);
nor U1029 (N_1029,In_114,In_699);
or U1030 (N_1030,In_370,In_843);
nand U1031 (N_1031,In_259,In_454);
or U1032 (N_1032,In_462,In_893);
or U1033 (N_1033,In_157,In_175);
or U1034 (N_1034,In_317,In_636);
nand U1035 (N_1035,In_747,In_635);
nand U1036 (N_1036,In_531,In_288);
nor U1037 (N_1037,In_150,In_402);
or U1038 (N_1038,In_839,In_902);
and U1039 (N_1039,In_266,In_551);
or U1040 (N_1040,In_667,In_291);
nand U1041 (N_1041,In_887,In_124);
nor U1042 (N_1042,In_575,In_54);
nor U1043 (N_1043,In_685,In_878);
and U1044 (N_1044,In_775,In_442);
or U1045 (N_1045,In_77,In_984);
or U1046 (N_1046,In_192,In_938);
or U1047 (N_1047,In_413,In_414);
xnor U1048 (N_1048,In_942,In_340);
and U1049 (N_1049,In_489,In_573);
nand U1050 (N_1050,In_970,In_717);
nor U1051 (N_1051,In_392,In_502);
or U1052 (N_1052,In_269,In_214);
nor U1053 (N_1053,In_338,In_333);
or U1054 (N_1054,In_473,In_36);
nand U1055 (N_1055,In_323,In_532);
nor U1056 (N_1056,In_370,In_435);
or U1057 (N_1057,In_459,In_827);
nand U1058 (N_1058,In_192,In_622);
nor U1059 (N_1059,In_145,In_641);
and U1060 (N_1060,In_748,In_654);
or U1061 (N_1061,In_636,In_220);
and U1062 (N_1062,In_310,In_762);
and U1063 (N_1063,In_352,In_531);
nand U1064 (N_1064,In_104,In_392);
nor U1065 (N_1065,In_815,In_338);
or U1066 (N_1066,In_359,In_537);
or U1067 (N_1067,In_379,In_243);
or U1068 (N_1068,In_540,In_970);
and U1069 (N_1069,In_185,In_883);
xnor U1070 (N_1070,In_29,In_236);
nand U1071 (N_1071,In_273,In_522);
and U1072 (N_1072,In_451,In_862);
and U1073 (N_1073,In_805,In_527);
nor U1074 (N_1074,In_715,In_496);
or U1075 (N_1075,In_962,In_667);
nor U1076 (N_1076,In_157,In_732);
or U1077 (N_1077,In_445,In_839);
or U1078 (N_1078,In_942,In_837);
nand U1079 (N_1079,In_463,In_1);
nor U1080 (N_1080,In_971,In_730);
or U1081 (N_1081,In_400,In_64);
nor U1082 (N_1082,In_924,In_131);
xnor U1083 (N_1083,In_394,In_986);
or U1084 (N_1084,In_42,In_812);
nand U1085 (N_1085,In_793,In_523);
and U1086 (N_1086,In_186,In_28);
nand U1087 (N_1087,In_329,In_160);
nand U1088 (N_1088,In_79,In_256);
nor U1089 (N_1089,In_255,In_259);
nand U1090 (N_1090,In_823,In_854);
and U1091 (N_1091,In_480,In_479);
nand U1092 (N_1092,In_538,In_280);
and U1093 (N_1093,In_656,In_458);
nor U1094 (N_1094,In_974,In_527);
xor U1095 (N_1095,In_401,In_971);
nor U1096 (N_1096,In_758,In_882);
and U1097 (N_1097,In_512,In_965);
xnor U1098 (N_1098,In_228,In_628);
xnor U1099 (N_1099,In_978,In_882);
xnor U1100 (N_1100,In_276,In_72);
nor U1101 (N_1101,In_848,In_170);
and U1102 (N_1102,In_944,In_247);
nor U1103 (N_1103,In_503,In_450);
or U1104 (N_1104,In_984,In_577);
nor U1105 (N_1105,In_954,In_128);
nand U1106 (N_1106,In_237,In_338);
nand U1107 (N_1107,In_327,In_707);
nor U1108 (N_1108,In_60,In_899);
and U1109 (N_1109,In_583,In_885);
or U1110 (N_1110,In_919,In_256);
and U1111 (N_1111,In_80,In_101);
nand U1112 (N_1112,In_195,In_897);
and U1113 (N_1113,In_550,In_231);
nor U1114 (N_1114,In_27,In_112);
or U1115 (N_1115,In_264,In_183);
nor U1116 (N_1116,In_232,In_886);
and U1117 (N_1117,In_534,In_405);
nand U1118 (N_1118,In_804,In_453);
and U1119 (N_1119,In_105,In_657);
nor U1120 (N_1120,In_151,In_797);
and U1121 (N_1121,In_894,In_752);
and U1122 (N_1122,In_435,In_697);
nand U1123 (N_1123,In_941,In_144);
xnor U1124 (N_1124,In_41,In_913);
and U1125 (N_1125,In_257,In_989);
nor U1126 (N_1126,In_379,In_525);
and U1127 (N_1127,In_627,In_503);
xor U1128 (N_1128,In_552,In_80);
nand U1129 (N_1129,In_107,In_280);
nand U1130 (N_1130,In_326,In_432);
or U1131 (N_1131,In_342,In_875);
or U1132 (N_1132,In_938,In_698);
or U1133 (N_1133,In_745,In_687);
nor U1134 (N_1134,In_431,In_336);
or U1135 (N_1135,In_484,In_150);
and U1136 (N_1136,In_740,In_537);
or U1137 (N_1137,In_112,In_923);
nand U1138 (N_1138,In_163,In_674);
xor U1139 (N_1139,In_67,In_987);
nand U1140 (N_1140,In_40,In_858);
or U1141 (N_1141,In_902,In_9);
nor U1142 (N_1142,In_3,In_190);
and U1143 (N_1143,In_787,In_92);
nand U1144 (N_1144,In_209,In_117);
nor U1145 (N_1145,In_156,In_668);
or U1146 (N_1146,In_217,In_67);
or U1147 (N_1147,In_417,In_444);
and U1148 (N_1148,In_979,In_703);
and U1149 (N_1149,In_645,In_930);
nor U1150 (N_1150,In_198,In_980);
and U1151 (N_1151,In_402,In_764);
or U1152 (N_1152,In_454,In_590);
and U1153 (N_1153,In_398,In_9);
nor U1154 (N_1154,In_375,In_172);
and U1155 (N_1155,In_217,In_477);
and U1156 (N_1156,In_836,In_488);
nor U1157 (N_1157,In_498,In_176);
nand U1158 (N_1158,In_910,In_732);
nor U1159 (N_1159,In_632,In_294);
or U1160 (N_1160,In_279,In_798);
nor U1161 (N_1161,In_940,In_139);
nor U1162 (N_1162,In_923,In_700);
and U1163 (N_1163,In_998,In_177);
and U1164 (N_1164,In_501,In_306);
nand U1165 (N_1165,In_672,In_480);
xor U1166 (N_1166,In_207,In_707);
nand U1167 (N_1167,In_820,In_206);
or U1168 (N_1168,In_970,In_264);
or U1169 (N_1169,In_821,In_445);
nor U1170 (N_1170,In_868,In_892);
or U1171 (N_1171,In_21,In_904);
and U1172 (N_1172,In_363,In_610);
and U1173 (N_1173,In_820,In_468);
or U1174 (N_1174,In_203,In_617);
and U1175 (N_1175,In_98,In_977);
and U1176 (N_1176,In_567,In_587);
nand U1177 (N_1177,In_947,In_198);
and U1178 (N_1178,In_64,In_263);
and U1179 (N_1179,In_359,In_0);
nor U1180 (N_1180,In_453,In_539);
nor U1181 (N_1181,In_310,In_651);
nand U1182 (N_1182,In_793,In_162);
nand U1183 (N_1183,In_95,In_534);
and U1184 (N_1184,In_462,In_507);
nand U1185 (N_1185,In_461,In_649);
and U1186 (N_1186,In_388,In_621);
nand U1187 (N_1187,In_30,In_448);
and U1188 (N_1188,In_956,In_506);
nor U1189 (N_1189,In_698,In_97);
nand U1190 (N_1190,In_859,In_842);
or U1191 (N_1191,In_84,In_90);
xnor U1192 (N_1192,In_266,In_415);
and U1193 (N_1193,In_620,In_167);
nor U1194 (N_1194,In_392,In_222);
nor U1195 (N_1195,In_128,In_765);
or U1196 (N_1196,In_352,In_433);
nor U1197 (N_1197,In_939,In_304);
or U1198 (N_1198,In_950,In_437);
or U1199 (N_1199,In_645,In_139);
xor U1200 (N_1200,In_452,In_787);
xor U1201 (N_1201,In_997,In_678);
or U1202 (N_1202,In_764,In_61);
nor U1203 (N_1203,In_588,In_202);
nand U1204 (N_1204,In_336,In_750);
and U1205 (N_1205,In_30,In_957);
nand U1206 (N_1206,In_357,In_952);
nor U1207 (N_1207,In_478,In_796);
or U1208 (N_1208,In_70,In_679);
nand U1209 (N_1209,In_334,In_896);
and U1210 (N_1210,In_226,In_84);
nand U1211 (N_1211,In_466,In_766);
and U1212 (N_1212,In_140,In_163);
xnor U1213 (N_1213,In_487,In_971);
xor U1214 (N_1214,In_17,In_966);
nand U1215 (N_1215,In_610,In_966);
nand U1216 (N_1216,In_582,In_772);
nor U1217 (N_1217,In_920,In_35);
or U1218 (N_1218,In_243,In_154);
nor U1219 (N_1219,In_655,In_676);
nor U1220 (N_1220,In_863,In_318);
or U1221 (N_1221,In_937,In_657);
nor U1222 (N_1222,In_246,In_31);
nor U1223 (N_1223,In_89,In_450);
nand U1224 (N_1224,In_166,In_444);
nand U1225 (N_1225,In_370,In_891);
nor U1226 (N_1226,In_91,In_651);
or U1227 (N_1227,In_491,In_316);
nand U1228 (N_1228,In_340,In_717);
nand U1229 (N_1229,In_649,In_551);
nor U1230 (N_1230,In_772,In_893);
nor U1231 (N_1231,In_142,In_414);
nand U1232 (N_1232,In_10,In_68);
and U1233 (N_1233,In_716,In_213);
xnor U1234 (N_1234,In_211,In_114);
nor U1235 (N_1235,In_208,In_589);
nor U1236 (N_1236,In_77,In_141);
and U1237 (N_1237,In_917,In_52);
or U1238 (N_1238,In_410,In_203);
nor U1239 (N_1239,In_58,In_42);
or U1240 (N_1240,In_355,In_938);
nand U1241 (N_1241,In_323,In_598);
nor U1242 (N_1242,In_363,In_856);
nor U1243 (N_1243,In_747,In_599);
and U1244 (N_1244,In_363,In_120);
xor U1245 (N_1245,In_716,In_66);
and U1246 (N_1246,In_462,In_943);
xor U1247 (N_1247,In_166,In_841);
nand U1248 (N_1248,In_248,In_748);
nand U1249 (N_1249,In_752,In_706);
nor U1250 (N_1250,In_190,In_908);
or U1251 (N_1251,In_527,In_477);
or U1252 (N_1252,In_213,In_114);
xor U1253 (N_1253,In_684,In_910);
or U1254 (N_1254,In_94,In_128);
and U1255 (N_1255,In_604,In_739);
and U1256 (N_1256,In_25,In_930);
nand U1257 (N_1257,In_114,In_160);
and U1258 (N_1258,In_66,In_278);
nand U1259 (N_1259,In_706,In_311);
or U1260 (N_1260,In_880,In_133);
and U1261 (N_1261,In_666,In_567);
xnor U1262 (N_1262,In_51,In_856);
or U1263 (N_1263,In_73,In_557);
or U1264 (N_1264,In_658,In_800);
and U1265 (N_1265,In_930,In_830);
nor U1266 (N_1266,In_227,In_762);
or U1267 (N_1267,In_648,In_96);
or U1268 (N_1268,In_955,In_591);
and U1269 (N_1269,In_486,In_638);
and U1270 (N_1270,In_633,In_119);
nand U1271 (N_1271,In_98,In_605);
and U1272 (N_1272,In_772,In_226);
nor U1273 (N_1273,In_261,In_39);
nand U1274 (N_1274,In_904,In_716);
or U1275 (N_1275,In_207,In_356);
or U1276 (N_1276,In_352,In_744);
xnor U1277 (N_1277,In_321,In_519);
or U1278 (N_1278,In_181,In_457);
nand U1279 (N_1279,In_269,In_490);
nor U1280 (N_1280,In_877,In_774);
or U1281 (N_1281,In_897,In_721);
nor U1282 (N_1282,In_562,In_338);
nand U1283 (N_1283,In_984,In_8);
and U1284 (N_1284,In_948,In_194);
nor U1285 (N_1285,In_526,In_805);
nand U1286 (N_1286,In_420,In_504);
xnor U1287 (N_1287,In_973,In_920);
nor U1288 (N_1288,In_270,In_770);
nor U1289 (N_1289,In_901,In_884);
or U1290 (N_1290,In_109,In_977);
and U1291 (N_1291,In_30,In_920);
nand U1292 (N_1292,In_536,In_733);
and U1293 (N_1293,In_299,In_97);
and U1294 (N_1294,In_797,In_696);
or U1295 (N_1295,In_653,In_830);
nand U1296 (N_1296,In_26,In_116);
and U1297 (N_1297,In_935,In_870);
and U1298 (N_1298,In_445,In_207);
nor U1299 (N_1299,In_937,In_255);
nand U1300 (N_1300,In_398,In_351);
nor U1301 (N_1301,In_823,In_615);
nand U1302 (N_1302,In_924,In_245);
and U1303 (N_1303,In_755,In_470);
nand U1304 (N_1304,In_677,In_502);
or U1305 (N_1305,In_693,In_98);
nor U1306 (N_1306,In_571,In_712);
or U1307 (N_1307,In_492,In_819);
and U1308 (N_1308,In_306,In_653);
nand U1309 (N_1309,In_348,In_598);
or U1310 (N_1310,In_748,In_358);
xnor U1311 (N_1311,In_46,In_702);
or U1312 (N_1312,In_658,In_884);
xor U1313 (N_1313,In_239,In_927);
or U1314 (N_1314,In_77,In_530);
nor U1315 (N_1315,In_939,In_81);
nor U1316 (N_1316,In_202,In_610);
and U1317 (N_1317,In_958,In_165);
or U1318 (N_1318,In_990,In_834);
nor U1319 (N_1319,In_268,In_952);
nor U1320 (N_1320,In_621,In_545);
or U1321 (N_1321,In_776,In_964);
and U1322 (N_1322,In_355,In_599);
nand U1323 (N_1323,In_417,In_321);
or U1324 (N_1324,In_68,In_250);
xnor U1325 (N_1325,In_153,In_632);
nor U1326 (N_1326,In_244,In_511);
xor U1327 (N_1327,In_240,In_700);
or U1328 (N_1328,In_920,In_316);
and U1329 (N_1329,In_714,In_942);
nand U1330 (N_1330,In_574,In_102);
xor U1331 (N_1331,In_956,In_544);
or U1332 (N_1332,In_231,In_443);
xor U1333 (N_1333,In_759,In_160);
and U1334 (N_1334,In_574,In_70);
or U1335 (N_1335,In_986,In_260);
nand U1336 (N_1336,In_338,In_611);
nand U1337 (N_1337,In_141,In_507);
nor U1338 (N_1338,In_427,In_804);
or U1339 (N_1339,In_422,In_380);
or U1340 (N_1340,In_146,In_67);
nor U1341 (N_1341,In_775,In_964);
xnor U1342 (N_1342,In_131,In_940);
and U1343 (N_1343,In_287,In_151);
nor U1344 (N_1344,In_411,In_355);
nand U1345 (N_1345,In_152,In_476);
nor U1346 (N_1346,In_17,In_520);
or U1347 (N_1347,In_109,In_740);
nor U1348 (N_1348,In_226,In_255);
and U1349 (N_1349,In_750,In_865);
or U1350 (N_1350,In_797,In_269);
and U1351 (N_1351,In_639,In_717);
nor U1352 (N_1352,In_660,In_821);
and U1353 (N_1353,In_76,In_511);
nor U1354 (N_1354,In_666,In_923);
or U1355 (N_1355,In_707,In_740);
and U1356 (N_1356,In_7,In_569);
and U1357 (N_1357,In_157,In_920);
or U1358 (N_1358,In_437,In_229);
xor U1359 (N_1359,In_478,In_936);
and U1360 (N_1360,In_5,In_100);
xnor U1361 (N_1361,In_654,In_632);
nand U1362 (N_1362,In_963,In_354);
and U1363 (N_1363,In_974,In_606);
or U1364 (N_1364,In_506,In_358);
or U1365 (N_1365,In_379,In_224);
nand U1366 (N_1366,In_348,In_168);
nand U1367 (N_1367,In_162,In_40);
or U1368 (N_1368,In_785,In_833);
nor U1369 (N_1369,In_878,In_253);
nand U1370 (N_1370,In_468,In_989);
nand U1371 (N_1371,In_152,In_607);
nor U1372 (N_1372,In_800,In_423);
and U1373 (N_1373,In_401,In_309);
nand U1374 (N_1374,In_128,In_147);
nand U1375 (N_1375,In_78,In_717);
or U1376 (N_1376,In_655,In_184);
nand U1377 (N_1377,In_193,In_572);
nor U1378 (N_1378,In_229,In_372);
nor U1379 (N_1379,In_917,In_102);
and U1380 (N_1380,In_152,In_698);
or U1381 (N_1381,In_907,In_353);
and U1382 (N_1382,In_654,In_47);
or U1383 (N_1383,In_93,In_545);
nor U1384 (N_1384,In_19,In_779);
nor U1385 (N_1385,In_880,In_178);
nand U1386 (N_1386,In_123,In_190);
or U1387 (N_1387,In_886,In_978);
nor U1388 (N_1388,In_334,In_985);
nand U1389 (N_1389,In_513,In_538);
and U1390 (N_1390,In_223,In_55);
nor U1391 (N_1391,In_741,In_929);
and U1392 (N_1392,In_68,In_86);
or U1393 (N_1393,In_791,In_117);
xnor U1394 (N_1394,In_484,In_682);
and U1395 (N_1395,In_332,In_997);
and U1396 (N_1396,In_792,In_603);
nand U1397 (N_1397,In_174,In_511);
and U1398 (N_1398,In_654,In_329);
and U1399 (N_1399,In_355,In_132);
nand U1400 (N_1400,In_851,In_218);
nor U1401 (N_1401,In_535,In_508);
or U1402 (N_1402,In_802,In_56);
nand U1403 (N_1403,In_784,In_909);
nor U1404 (N_1404,In_973,In_180);
nor U1405 (N_1405,In_828,In_345);
nor U1406 (N_1406,In_265,In_916);
nor U1407 (N_1407,In_859,In_449);
and U1408 (N_1408,In_43,In_759);
nand U1409 (N_1409,In_928,In_877);
or U1410 (N_1410,In_308,In_619);
xnor U1411 (N_1411,In_413,In_581);
and U1412 (N_1412,In_589,In_486);
nor U1413 (N_1413,In_408,In_599);
nor U1414 (N_1414,In_946,In_468);
nor U1415 (N_1415,In_556,In_295);
nor U1416 (N_1416,In_756,In_916);
and U1417 (N_1417,In_73,In_123);
nor U1418 (N_1418,In_863,In_739);
nor U1419 (N_1419,In_889,In_748);
and U1420 (N_1420,In_722,In_377);
nand U1421 (N_1421,In_209,In_898);
nor U1422 (N_1422,In_875,In_583);
nand U1423 (N_1423,In_172,In_799);
and U1424 (N_1424,In_127,In_77);
nand U1425 (N_1425,In_219,In_666);
or U1426 (N_1426,In_314,In_812);
or U1427 (N_1427,In_116,In_972);
nand U1428 (N_1428,In_547,In_120);
nor U1429 (N_1429,In_185,In_940);
or U1430 (N_1430,In_289,In_505);
and U1431 (N_1431,In_435,In_287);
and U1432 (N_1432,In_38,In_593);
nand U1433 (N_1433,In_347,In_75);
or U1434 (N_1434,In_217,In_992);
nand U1435 (N_1435,In_436,In_826);
nand U1436 (N_1436,In_14,In_279);
xnor U1437 (N_1437,In_104,In_935);
nor U1438 (N_1438,In_775,In_425);
nand U1439 (N_1439,In_165,In_457);
and U1440 (N_1440,In_882,In_397);
nor U1441 (N_1441,In_943,In_104);
nand U1442 (N_1442,In_959,In_330);
nor U1443 (N_1443,In_677,In_580);
nor U1444 (N_1444,In_189,In_578);
xnor U1445 (N_1445,In_28,In_373);
nor U1446 (N_1446,In_67,In_852);
nand U1447 (N_1447,In_969,In_921);
nor U1448 (N_1448,In_130,In_542);
or U1449 (N_1449,In_162,In_756);
or U1450 (N_1450,In_511,In_461);
nor U1451 (N_1451,In_630,In_763);
xnor U1452 (N_1452,In_379,In_943);
or U1453 (N_1453,In_959,In_93);
nand U1454 (N_1454,In_498,In_640);
or U1455 (N_1455,In_742,In_685);
nand U1456 (N_1456,In_760,In_418);
or U1457 (N_1457,In_264,In_900);
and U1458 (N_1458,In_771,In_298);
nor U1459 (N_1459,In_114,In_248);
nor U1460 (N_1460,In_832,In_516);
and U1461 (N_1461,In_52,In_969);
or U1462 (N_1462,In_567,In_103);
or U1463 (N_1463,In_488,In_601);
or U1464 (N_1464,In_368,In_93);
nor U1465 (N_1465,In_246,In_972);
nor U1466 (N_1466,In_301,In_161);
nor U1467 (N_1467,In_982,In_263);
nor U1468 (N_1468,In_158,In_817);
nor U1469 (N_1469,In_906,In_521);
and U1470 (N_1470,In_924,In_311);
nand U1471 (N_1471,In_731,In_422);
nand U1472 (N_1472,In_259,In_633);
or U1473 (N_1473,In_78,In_611);
nand U1474 (N_1474,In_537,In_548);
xnor U1475 (N_1475,In_836,In_323);
and U1476 (N_1476,In_164,In_220);
nand U1477 (N_1477,In_232,In_423);
nand U1478 (N_1478,In_836,In_893);
and U1479 (N_1479,In_936,In_337);
nand U1480 (N_1480,In_792,In_324);
nor U1481 (N_1481,In_719,In_519);
nor U1482 (N_1482,In_505,In_75);
or U1483 (N_1483,In_163,In_616);
nor U1484 (N_1484,In_645,In_326);
nor U1485 (N_1485,In_794,In_118);
and U1486 (N_1486,In_563,In_199);
nor U1487 (N_1487,In_292,In_291);
nand U1488 (N_1488,In_537,In_211);
nor U1489 (N_1489,In_100,In_56);
nand U1490 (N_1490,In_447,In_610);
nor U1491 (N_1491,In_581,In_584);
and U1492 (N_1492,In_821,In_950);
nand U1493 (N_1493,In_889,In_800);
or U1494 (N_1494,In_260,In_582);
nor U1495 (N_1495,In_947,In_673);
or U1496 (N_1496,In_0,In_134);
and U1497 (N_1497,In_540,In_518);
xnor U1498 (N_1498,In_821,In_357);
nand U1499 (N_1499,In_111,In_613);
or U1500 (N_1500,In_26,In_106);
and U1501 (N_1501,In_377,In_684);
or U1502 (N_1502,In_739,In_809);
and U1503 (N_1503,In_130,In_882);
and U1504 (N_1504,In_697,In_145);
or U1505 (N_1505,In_85,In_743);
xnor U1506 (N_1506,In_952,In_391);
nor U1507 (N_1507,In_242,In_287);
nor U1508 (N_1508,In_209,In_961);
and U1509 (N_1509,In_444,In_219);
and U1510 (N_1510,In_637,In_88);
and U1511 (N_1511,In_178,In_381);
nor U1512 (N_1512,In_378,In_777);
nand U1513 (N_1513,In_235,In_73);
nand U1514 (N_1514,In_862,In_887);
nor U1515 (N_1515,In_334,In_537);
nor U1516 (N_1516,In_616,In_968);
nand U1517 (N_1517,In_212,In_913);
nor U1518 (N_1518,In_766,In_752);
nand U1519 (N_1519,In_616,In_648);
or U1520 (N_1520,In_831,In_258);
nor U1521 (N_1521,In_686,In_779);
or U1522 (N_1522,In_412,In_187);
nor U1523 (N_1523,In_326,In_191);
nand U1524 (N_1524,In_668,In_765);
nand U1525 (N_1525,In_773,In_519);
nand U1526 (N_1526,In_420,In_37);
or U1527 (N_1527,In_310,In_736);
xor U1528 (N_1528,In_353,In_980);
nor U1529 (N_1529,In_415,In_308);
and U1530 (N_1530,In_946,In_664);
nor U1531 (N_1531,In_781,In_991);
and U1532 (N_1532,In_116,In_259);
nor U1533 (N_1533,In_449,In_563);
nand U1534 (N_1534,In_753,In_126);
and U1535 (N_1535,In_472,In_709);
or U1536 (N_1536,In_882,In_104);
and U1537 (N_1537,In_634,In_788);
or U1538 (N_1538,In_171,In_178);
and U1539 (N_1539,In_818,In_843);
nand U1540 (N_1540,In_758,In_330);
nand U1541 (N_1541,In_68,In_500);
and U1542 (N_1542,In_940,In_481);
nor U1543 (N_1543,In_885,In_157);
nand U1544 (N_1544,In_205,In_604);
nand U1545 (N_1545,In_147,In_212);
and U1546 (N_1546,In_695,In_164);
nor U1547 (N_1547,In_893,In_941);
nor U1548 (N_1548,In_796,In_429);
or U1549 (N_1549,In_121,In_480);
and U1550 (N_1550,In_521,In_834);
xor U1551 (N_1551,In_84,In_758);
or U1552 (N_1552,In_752,In_6);
nand U1553 (N_1553,In_259,In_666);
nand U1554 (N_1554,In_386,In_19);
nand U1555 (N_1555,In_144,In_793);
and U1556 (N_1556,In_605,In_992);
and U1557 (N_1557,In_641,In_412);
nor U1558 (N_1558,In_544,In_125);
xor U1559 (N_1559,In_997,In_297);
and U1560 (N_1560,In_476,In_35);
xor U1561 (N_1561,In_87,In_387);
nand U1562 (N_1562,In_283,In_27);
nand U1563 (N_1563,In_887,In_163);
or U1564 (N_1564,In_53,In_236);
and U1565 (N_1565,In_642,In_425);
and U1566 (N_1566,In_509,In_471);
nor U1567 (N_1567,In_854,In_508);
nand U1568 (N_1568,In_485,In_866);
and U1569 (N_1569,In_234,In_701);
nand U1570 (N_1570,In_76,In_720);
or U1571 (N_1571,In_598,In_136);
xor U1572 (N_1572,In_450,In_132);
and U1573 (N_1573,In_357,In_778);
nor U1574 (N_1574,In_220,In_177);
or U1575 (N_1575,In_428,In_530);
nor U1576 (N_1576,In_343,In_361);
or U1577 (N_1577,In_488,In_440);
or U1578 (N_1578,In_513,In_357);
xor U1579 (N_1579,In_211,In_545);
nor U1580 (N_1580,In_696,In_693);
nor U1581 (N_1581,In_556,In_65);
nand U1582 (N_1582,In_94,In_104);
and U1583 (N_1583,In_919,In_686);
nand U1584 (N_1584,In_322,In_723);
nor U1585 (N_1585,In_815,In_362);
nor U1586 (N_1586,In_323,In_153);
nor U1587 (N_1587,In_476,In_28);
or U1588 (N_1588,In_612,In_962);
nand U1589 (N_1589,In_397,In_578);
xor U1590 (N_1590,In_126,In_773);
or U1591 (N_1591,In_339,In_999);
and U1592 (N_1592,In_984,In_931);
nand U1593 (N_1593,In_820,In_618);
xnor U1594 (N_1594,In_487,In_920);
or U1595 (N_1595,In_764,In_21);
and U1596 (N_1596,In_272,In_526);
xnor U1597 (N_1597,In_496,In_317);
or U1598 (N_1598,In_303,In_227);
nand U1599 (N_1599,In_379,In_614);
nor U1600 (N_1600,In_238,In_413);
xor U1601 (N_1601,In_129,In_77);
and U1602 (N_1602,In_82,In_458);
nand U1603 (N_1603,In_904,In_821);
nor U1604 (N_1604,In_689,In_64);
or U1605 (N_1605,In_52,In_691);
xor U1606 (N_1606,In_604,In_46);
nand U1607 (N_1607,In_476,In_136);
xor U1608 (N_1608,In_904,In_915);
nor U1609 (N_1609,In_292,In_220);
or U1610 (N_1610,In_264,In_245);
or U1611 (N_1611,In_575,In_970);
xor U1612 (N_1612,In_887,In_414);
or U1613 (N_1613,In_154,In_584);
nor U1614 (N_1614,In_254,In_676);
nand U1615 (N_1615,In_359,In_354);
and U1616 (N_1616,In_383,In_517);
nor U1617 (N_1617,In_803,In_192);
xor U1618 (N_1618,In_960,In_354);
and U1619 (N_1619,In_699,In_353);
nor U1620 (N_1620,In_869,In_553);
or U1621 (N_1621,In_314,In_99);
or U1622 (N_1622,In_460,In_617);
or U1623 (N_1623,In_196,In_396);
xor U1624 (N_1624,In_57,In_790);
nand U1625 (N_1625,In_255,In_658);
or U1626 (N_1626,In_759,In_500);
xor U1627 (N_1627,In_990,In_217);
nand U1628 (N_1628,In_923,In_67);
or U1629 (N_1629,In_73,In_839);
or U1630 (N_1630,In_326,In_9);
or U1631 (N_1631,In_642,In_727);
nor U1632 (N_1632,In_972,In_354);
or U1633 (N_1633,In_860,In_799);
nand U1634 (N_1634,In_245,In_546);
xor U1635 (N_1635,In_79,In_339);
and U1636 (N_1636,In_820,In_743);
or U1637 (N_1637,In_831,In_429);
xnor U1638 (N_1638,In_8,In_541);
nor U1639 (N_1639,In_519,In_750);
and U1640 (N_1640,In_816,In_13);
xnor U1641 (N_1641,In_565,In_380);
or U1642 (N_1642,In_411,In_906);
or U1643 (N_1643,In_494,In_971);
nand U1644 (N_1644,In_1,In_139);
xor U1645 (N_1645,In_717,In_319);
xor U1646 (N_1646,In_704,In_11);
xnor U1647 (N_1647,In_683,In_147);
or U1648 (N_1648,In_47,In_345);
nand U1649 (N_1649,In_220,In_534);
nor U1650 (N_1650,In_865,In_749);
and U1651 (N_1651,In_722,In_869);
and U1652 (N_1652,In_946,In_952);
or U1653 (N_1653,In_290,In_908);
nand U1654 (N_1654,In_398,In_45);
and U1655 (N_1655,In_451,In_210);
xnor U1656 (N_1656,In_825,In_891);
and U1657 (N_1657,In_888,In_818);
xor U1658 (N_1658,In_780,In_909);
nand U1659 (N_1659,In_853,In_875);
or U1660 (N_1660,In_737,In_994);
or U1661 (N_1661,In_251,In_528);
nand U1662 (N_1662,In_899,In_736);
nand U1663 (N_1663,In_544,In_660);
nor U1664 (N_1664,In_567,In_250);
xnor U1665 (N_1665,In_781,In_870);
nor U1666 (N_1666,In_230,In_96);
nor U1667 (N_1667,In_330,In_799);
or U1668 (N_1668,In_21,In_961);
or U1669 (N_1669,In_137,In_390);
nor U1670 (N_1670,In_450,In_695);
nand U1671 (N_1671,In_170,In_62);
or U1672 (N_1672,In_336,In_176);
and U1673 (N_1673,In_7,In_792);
xnor U1674 (N_1674,In_523,In_111);
nand U1675 (N_1675,In_918,In_877);
nand U1676 (N_1676,In_851,In_874);
and U1677 (N_1677,In_784,In_440);
nor U1678 (N_1678,In_322,In_939);
nor U1679 (N_1679,In_124,In_871);
nand U1680 (N_1680,In_61,In_678);
and U1681 (N_1681,In_38,In_516);
nor U1682 (N_1682,In_483,In_640);
nand U1683 (N_1683,In_278,In_529);
or U1684 (N_1684,In_333,In_119);
nor U1685 (N_1685,In_756,In_912);
and U1686 (N_1686,In_549,In_336);
xnor U1687 (N_1687,In_949,In_932);
nand U1688 (N_1688,In_821,In_348);
nand U1689 (N_1689,In_354,In_803);
or U1690 (N_1690,In_363,In_287);
or U1691 (N_1691,In_696,In_491);
and U1692 (N_1692,In_371,In_503);
and U1693 (N_1693,In_667,In_792);
or U1694 (N_1694,In_362,In_978);
and U1695 (N_1695,In_189,In_517);
or U1696 (N_1696,In_818,In_690);
and U1697 (N_1697,In_973,In_640);
nand U1698 (N_1698,In_17,In_911);
nor U1699 (N_1699,In_582,In_198);
nand U1700 (N_1700,In_249,In_750);
nor U1701 (N_1701,In_424,In_243);
xor U1702 (N_1702,In_230,In_165);
and U1703 (N_1703,In_301,In_652);
nor U1704 (N_1704,In_418,In_183);
xnor U1705 (N_1705,In_447,In_931);
nor U1706 (N_1706,In_916,In_575);
nand U1707 (N_1707,In_455,In_587);
or U1708 (N_1708,In_229,In_590);
and U1709 (N_1709,In_463,In_85);
xnor U1710 (N_1710,In_372,In_326);
or U1711 (N_1711,In_438,In_926);
nor U1712 (N_1712,In_944,In_914);
and U1713 (N_1713,In_656,In_885);
and U1714 (N_1714,In_25,In_840);
and U1715 (N_1715,In_10,In_616);
nor U1716 (N_1716,In_384,In_797);
nor U1717 (N_1717,In_866,In_56);
and U1718 (N_1718,In_783,In_756);
nand U1719 (N_1719,In_115,In_367);
nor U1720 (N_1720,In_442,In_470);
or U1721 (N_1721,In_647,In_628);
xor U1722 (N_1722,In_48,In_977);
and U1723 (N_1723,In_69,In_266);
and U1724 (N_1724,In_422,In_260);
nand U1725 (N_1725,In_489,In_369);
nor U1726 (N_1726,In_63,In_942);
or U1727 (N_1727,In_328,In_429);
or U1728 (N_1728,In_568,In_772);
nor U1729 (N_1729,In_202,In_901);
or U1730 (N_1730,In_240,In_7);
nand U1731 (N_1731,In_104,In_932);
nand U1732 (N_1732,In_184,In_779);
or U1733 (N_1733,In_330,In_305);
or U1734 (N_1734,In_947,In_616);
nand U1735 (N_1735,In_867,In_368);
nor U1736 (N_1736,In_269,In_637);
or U1737 (N_1737,In_927,In_292);
and U1738 (N_1738,In_313,In_12);
and U1739 (N_1739,In_515,In_84);
xor U1740 (N_1740,In_80,In_384);
nor U1741 (N_1741,In_682,In_725);
nand U1742 (N_1742,In_738,In_420);
nor U1743 (N_1743,In_551,In_928);
and U1744 (N_1744,In_167,In_130);
and U1745 (N_1745,In_980,In_269);
or U1746 (N_1746,In_244,In_862);
nand U1747 (N_1747,In_168,In_823);
nand U1748 (N_1748,In_428,In_874);
or U1749 (N_1749,In_59,In_866);
nor U1750 (N_1750,In_861,In_75);
nand U1751 (N_1751,In_902,In_852);
or U1752 (N_1752,In_622,In_583);
nand U1753 (N_1753,In_219,In_460);
or U1754 (N_1754,In_522,In_528);
and U1755 (N_1755,In_165,In_549);
nor U1756 (N_1756,In_343,In_794);
nor U1757 (N_1757,In_847,In_964);
or U1758 (N_1758,In_501,In_119);
nand U1759 (N_1759,In_86,In_95);
and U1760 (N_1760,In_122,In_324);
nor U1761 (N_1761,In_268,In_14);
nor U1762 (N_1762,In_349,In_215);
or U1763 (N_1763,In_454,In_668);
nand U1764 (N_1764,In_119,In_205);
and U1765 (N_1765,In_169,In_516);
nand U1766 (N_1766,In_513,In_676);
nand U1767 (N_1767,In_703,In_957);
nor U1768 (N_1768,In_292,In_751);
or U1769 (N_1769,In_454,In_786);
or U1770 (N_1770,In_493,In_898);
and U1771 (N_1771,In_572,In_312);
and U1772 (N_1772,In_154,In_924);
nand U1773 (N_1773,In_104,In_723);
nand U1774 (N_1774,In_210,In_913);
nand U1775 (N_1775,In_62,In_157);
xnor U1776 (N_1776,In_212,In_736);
nand U1777 (N_1777,In_341,In_823);
and U1778 (N_1778,In_474,In_46);
nor U1779 (N_1779,In_399,In_878);
or U1780 (N_1780,In_923,In_93);
nor U1781 (N_1781,In_709,In_332);
or U1782 (N_1782,In_382,In_818);
nor U1783 (N_1783,In_791,In_761);
nor U1784 (N_1784,In_992,In_351);
xnor U1785 (N_1785,In_626,In_853);
and U1786 (N_1786,In_385,In_43);
nor U1787 (N_1787,In_21,In_541);
xor U1788 (N_1788,In_885,In_128);
and U1789 (N_1789,In_715,In_474);
and U1790 (N_1790,In_489,In_466);
xnor U1791 (N_1791,In_21,In_243);
or U1792 (N_1792,In_366,In_786);
or U1793 (N_1793,In_911,In_954);
nor U1794 (N_1794,In_449,In_825);
nor U1795 (N_1795,In_106,In_947);
and U1796 (N_1796,In_686,In_606);
and U1797 (N_1797,In_310,In_549);
nand U1798 (N_1798,In_412,In_661);
xor U1799 (N_1799,In_630,In_86);
nor U1800 (N_1800,In_560,In_595);
or U1801 (N_1801,In_933,In_739);
nor U1802 (N_1802,In_652,In_833);
or U1803 (N_1803,In_832,In_336);
nor U1804 (N_1804,In_274,In_836);
nand U1805 (N_1805,In_621,In_433);
or U1806 (N_1806,In_200,In_181);
or U1807 (N_1807,In_625,In_24);
nand U1808 (N_1808,In_215,In_253);
or U1809 (N_1809,In_361,In_201);
nand U1810 (N_1810,In_754,In_942);
or U1811 (N_1811,In_370,In_289);
nand U1812 (N_1812,In_787,In_170);
nand U1813 (N_1813,In_765,In_594);
and U1814 (N_1814,In_566,In_77);
or U1815 (N_1815,In_233,In_393);
or U1816 (N_1816,In_755,In_539);
or U1817 (N_1817,In_989,In_880);
and U1818 (N_1818,In_259,In_828);
or U1819 (N_1819,In_551,In_908);
and U1820 (N_1820,In_471,In_711);
xnor U1821 (N_1821,In_706,In_382);
nand U1822 (N_1822,In_298,In_559);
or U1823 (N_1823,In_172,In_184);
and U1824 (N_1824,In_670,In_941);
nor U1825 (N_1825,In_836,In_756);
nor U1826 (N_1826,In_51,In_762);
or U1827 (N_1827,In_326,In_167);
or U1828 (N_1828,In_807,In_670);
nand U1829 (N_1829,In_442,In_144);
nand U1830 (N_1830,In_654,In_946);
nor U1831 (N_1831,In_854,In_928);
and U1832 (N_1832,In_581,In_632);
nand U1833 (N_1833,In_447,In_372);
nor U1834 (N_1834,In_84,In_391);
or U1835 (N_1835,In_599,In_919);
and U1836 (N_1836,In_285,In_491);
nand U1837 (N_1837,In_116,In_187);
nor U1838 (N_1838,In_518,In_414);
xor U1839 (N_1839,In_545,In_771);
and U1840 (N_1840,In_137,In_829);
and U1841 (N_1841,In_727,In_232);
xor U1842 (N_1842,In_363,In_405);
or U1843 (N_1843,In_622,In_203);
nand U1844 (N_1844,In_609,In_882);
nor U1845 (N_1845,In_998,In_740);
and U1846 (N_1846,In_842,In_483);
and U1847 (N_1847,In_465,In_132);
and U1848 (N_1848,In_537,In_685);
or U1849 (N_1849,In_959,In_152);
or U1850 (N_1850,In_849,In_804);
or U1851 (N_1851,In_886,In_3);
and U1852 (N_1852,In_624,In_199);
and U1853 (N_1853,In_179,In_429);
xnor U1854 (N_1854,In_233,In_764);
nand U1855 (N_1855,In_57,In_8);
xor U1856 (N_1856,In_943,In_301);
nor U1857 (N_1857,In_128,In_196);
nor U1858 (N_1858,In_263,In_714);
nor U1859 (N_1859,In_78,In_247);
and U1860 (N_1860,In_557,In_817);
and U1861 (N_1861,In_502,In_733);
and U1862 (N_1862,In_776,In_419);
or U1863 (N_1863,In_687,In_556);
nand U1864 (N_1864,In_863,In_346);
or U1865 (N_1865,In_708,In_740);
nor U1866 (N_1866,In_308,In_431);
or U1867 (N_1867,In_857,In_280);
nand U1868 (N_1868,In_511,In_414);
or U1869 (N_1869,In_892,In_606);
or U1870 (N_1870,In_430,In_677);
xor U1871 (N_1871,In_577,In_969);
or U1872 (N_1872,In_933,In_588);
nor U1873 (N_1873,In_874,In_38);
and U1874 (N_1874,In_330,In_20);
xor U1875 (N_1875,In_179,In_860);
nor U1876 (N_1876,In_456,In_836);
nand U1877 (N_1877,In_466,In_200);
xor U1878 (N_1878,In_135,In_555);
or U1879 (N_1879,In_58,In_298);
nor U1880 (N_1880,In_826,In_936);
nand U1881 (N_1881,In_319,In_421);
nand U1882 (N_1882,In_606,In_120);
nor U1883 (N_1883,In_156,In_871);
nor U1884 (N_1884,In_645,In_971);
and U1885 (N_1885,In_432,In_134);
nor U1886 (N_1886,In_74,In_704);
or U1887 (N_1887,In_925,In_563);
nand U1888 (N_1888,In_169,In_480);
nor U1889 (N_1889,In_121,In_263);
and U1890 (N_1890,In_154,In_27);
nand U1891 (N_1891,In_115,In_54);
nor U1892 (N_1892,In_311,In_901);
xnor U1893 (N_1893,In_60,In_179);
and U1894 (N_1894,In_113,In_269);
nor U1895 (N_1895,In_834,In_873);
or U1896 (N_1896,In_262,In_662);
nor U1897 (N_1897,In_143,In_622);
or U1898 (N_1898,In_158,In_553);
and U1899 (N_1899,In_767,In_781);
nand U1900 (N_1900,In_972,In_122);
xor U1901 (N_1901,In_314,In_3);
nor U1902 (N_1902,In_541,In_150);
nand U1903 (N_1903,In_467,In_816);
or U1904 (N_1904,In_153,In_158);
or U1905 (N_1905,In_697,In_174);
nor U1906 (N_1906,In_875,In_912);
nor U1907 (N_1907,In_518,In_467);
or U1908 (N_1908,In_647,In_149);
nor U1909 (N_1909,In_736,In_953);
nor U1910 (N_1910,In_68,In_24);
nor U1911 (N_1911,In_984,In_827);
or U1912 (N_1912,In_965,In_507);
nor U1913 (N_1913,In_333,In_598);
nand U1914 (N_1914,In_84,In_677);
nand U1915 (N_1915,In_767,In_852);
xnor U1916 (N_1916,In_287,In_408);
or U1917 (N_1917,In_489,In_656);
xor U1918 (N_1918,In_276,In_95);
and U1919 (N_1919,In_295,In_21);
and U1920 (N_1920,In_356,In_738);
nand U1921 (N_1921,In_273,In_745);
nand U1922 (N_1922,In_509,In_993);
nor U1923 (N_1923,In_104,In_992);
or U1924 (N_1924,In_832,In_818);
nor U1925 (N_1925,In_693,In_44);
nand U1926 (N_1926,In_789,In_487);
nor U1927 (N_1927,In_274,In_52);
and U1928 (N_1928,In_898,In_241);
nor U1929 (N_1929,In_296,In_273);
nor U1930 (N_1930,In_691,In_89);
nor U1931 (N_1931,In_309,In_638);
nor U1932 (N_1932,In_275,In_456);
or U1933 (N_1933,In_866,In_562);
nand U1934 (N_1934,In_259,In_328);
or U1935 (N_1935,In_898,In_104);
and U1936 (N_1936,In_44,In_389);
and U1937 (N_1937,In_537,In_182);
nor U1938 (N_1938,In_355,In_268);
or U1939 (N_1939,In_671,In_620);
xor U1940 (N_1940,In_953,In_50);
and U1941 (N_1941,In_411,In_944);
nor U1942 (N_1942,In_94,In_459);
xnor U1943 (N_1943,In_145,In_775);
or U1944 (N_1944,In_581,In_784);
nor U1945 (N_1945,In_344,In_758);
nand U1946 (N_1946,In_786,In_254);
nand U1947 (N_1947,In_278,In_874);
or U1948 (N_1948,In_768,In_897);
nor U1949 (N_1949,In_741,In_983);
and U1950 (N_1950,In_351,In_822);
and U1951 (N_1951,In_400,In_143);
or U1952 (N_1952,In_878,In_887);
nor U1953 (N_1953,In_214,In_575);
nor U1954 (N_1954,In_72,In_449);
or U1955 (N_1955,In_228,In_182);
nor U1956 (N_1956,In_395,In_56);
and U1957 (N_1957,In_218,In_60);
nand U1958 (N_1958,In_860,In_117);
or U1959 (N_1959,In_231,In_761);
nor U1960 (N_1960,In_274,In_688);
nor U1961 (N_1961,In_654,In_678);
nor U1962 (N_1962,In_722,In_354);
and U1963 (N_1963,In_325,In_272);
xor U1964 (N_1964,In_23,In_568);
nor U1965 (N_1965,In_557,In_720);
or U1966 (N_1966,In_645,In_909);
nor U1967 (N_1967,In_462,In_140);
and U1968 (N_1968,In_304,In_635);
and U1969 (N_1969,In_801,In_430);
or U1970 (N_1970,In_647,In_579);
nor U1971 (N_1971,In_953,In_490);
nand U1972 (N_1972,In_545,In_790);
nand U1973 (N_1973,In_677,In_840);
and U1974 (N_1974,In_715,In_67);
and U1975 (N_1975,In_516,In_331);
nand U1976 (N_1976,In_198,In_695);
or U1977 (N_1977,In_634,In_866);
nor U1978 (N_1978,In_751,In_278);
nor U1979 (N_1979,In_466,In_780);
and U1980 (N_1980,In_460,In_662);
nor U1981 (N_1981,In_117,In_629);
or U1982 (N_1982,In_116,In_561);
and U1983 (N_1983,In_810,In_714);
nand U1984 (N_1984,In_752,In_205);
nand U1985 (N_1985,In_970,In_56);
or U1986 (N_1986,In_274,In_331);
nor U1987 (N_1987,In_438,In_258);
nor U1988 (N_1988,In_365,In_501);
and U1989 (N_1989,In_297,In_386);
or U1990 (N_1990,In_126,In_958);
and U1991 (N_1991,In_688,In_861);
and U1992 (N_1992,In_103,In_392);
nand U1993 (N_1993,In_443,In_96);
nand U1994 (N_1994,In_491,In_349);
or U1995 (N_1995,In_928,In_130);
xnor U1996 (N_1996,In_629,In_582);
and U1997 (N_1997,In_267,In_475);
nand U1998 (N_1998,In_116,In_179);
nand U1999 (N_1999,In_712,In_936);
and U2000 (N_2000,N_782,N_202);
nand U2001 (N_2001,N_1312,N_559);
and U2002 (N_2002,N_1498,N_707);
nor U2003 (N_2003,N_1641,N_1910);
nand U2004 (N_2004,N_258,N_712);
nor U2005 (N_2005,N_1194,N_1866);
nand U2006 (N_2006,N_1882,N_848);
nor U2007 (N_2007,N_506,N_588);
nor U2008 (N_2008,N_1255,N_408);
xor U2009 (N_2009,N_355,N_1804);
nand U2010 (N_2010,N_1577,N_553);
xor U2011 (N_2011,N_1684,N_179);
and U2012 (N_2012,N_665,N_141);
and U2013 (N_2013,N_226,N_1770);
or U2014 (N_2014,N_1940,N_1747);
xnor U2015 (N_2015,N_514,N_805);
or U2016 (N_2016,N_1693,N_490);
xnor U2017 (N_2017,N_422,N_1774);
nand U2018 (N_2018,N_872,N_1254);
nand U2019 (N_2019,N_1829,N_1298);
nor U2020 (N_2020,N_458,N_1619);
nand U2021 (N_2021,N_115,N_1314);
nand U2022 (N_2022,N_390,N_1405);
xor U2023 (N_2023,N_1607,N_522);
and U2024 (N_2024,N_239,N_1943);
nor U2025 (N_2025,N_1341,N_1425);
nand U2026 (N_2026,N_1566,N_806);
xnor U2027 (N_2027,N_1777,N_146);
nand U2028 (N_2028,N_352,N_1749);
nor U2029 (N_2029,N_619,N_338);
and U2030 (N_2030,N_1233,N_1685);
nand U2031 (N_2031,N_1987,N_1570);
nor U2032 (N_2032,N_1784,N_1841);
and U2033 (N_2033,N_1675,N_1129);
and U2034 (N_2034,N_1480,N_1152);
nand U2035 (N_2035,N_1980,N_1883);
or U2036 (N_2036,N_995,N_1632);
or U2037 (N_2037,N_613,N_108);
or U2038 (N_2038,N_384,N_1592);
nand U2039 (N_2039,N_1855,N_1831);
or U2040 (N_2040,N_201,N_574);
or U2041 (N_2041,N_66,N_1115);
nand U2042 (N_2042,N_519,N_1308);
nor U2043 (N_2043,N_394,N_1064);
nand U2044 (N_2044,N_1297,N_1960);
and U2045 (N_2045,N_1726,N_130);
nand U2046 (N_2046,N_38,N_16);
and U2047 (N_2047,N_1966,N_247);
xnor U2048 (N_2048,N_18,N_708);
or U2049 (N_2049,N_710,N_1005);
and U2050 (N_2050,N_1635,N_253);
nand U2051 (N_2051,N_77,N_109);
and U2052 (N_2052,N_630,N_1328);
nor U2053 (N_2053,N_614,N_891);
nor U2054 (N_2054,N_794,N_1089);
nand U2055 (N_2055,N_1846,N_402);
xor U2056 (N_2056,N_1216,N_699);
nand U2057 (N_2057,N_1847,N_1088);
nand U2058 (N_2058,N_1549,N_1168);
or U2059 (N_2059,N_902,N_1440);
or U2060 (N_2060,N_1256,N_494);
nor U2061 (N_2061,N_549,N_579);
and U2062 (N_2062,N_807,N_1914);
nor U2063 (N_2063,N_564,N_1184);
xnor U2064 (N_2064,N_1271,N_748);
nor U2065 (N_2065,N_628,N_1240);
and U2066 (N_2066,N_1106,N_1460);
and U2067 (N_2067,N_1172,N_1895);
or U2068 (N_2068,N_1019,N_1273);
or U2069 (N_2069,N_962,N_1718);
or U2070 (N_2070,N_627,N_1043);
or U2071 (N_2071,N_298,N_1588);
nand U2072 (N_2072,N_971,N_438);
nand U2073 (N_2073,N_1180,N_1560);
and U2074 (N_2074,N_40,N_334);
nor U2075 (N_2075,N_1664,N_974);
nand U2076 (N_2076,N_1579,N_1530);
nand U2077 (N_2077,N_263,N_1683);
and U2078 (N_2078,N_1125,N_1374);
or U2079 (N_2079,N_1080,N_1844);
nand U2080 (N_2080,N_1617,N_456);
nor U2081 (N_2081,N_119,N_575);
nor U2082 (N_2082,N_1919,N_606);
and U2083 (N_2083,N_1660,N_544);
nor U2084 (N_2084,N_155,N_1113);
nor U2085 (N_2085,N_137,N_1536);
nand U2086 (N_2086,N_1176,N_445);
and U2087 (N_2087,N_498,N_188);
nand U2088 (N_2088,N_593,N_1791);
xnor U2089 (N_2089,N_1996,N_1157);
xor U2090 (N_2090,N_819,N_436);
or U2091 (N_2091,N_735,N_1786);
nor U2092 (N_2092,N_1992,N_124);
and U2093 (N_2093,N_252,N_1020);
nor U2094 (N_2094,N_845,N_1410);
or U2095 (N_2095,N_1833,N_901);
and U2096 (N_2096,N_1821,N_1346);
xor U2097 (N_2097,N_80,N_1959);
and U2098 (N_2098,N_752,N_878);
nand U2099 (N_2099,N_1404,N_1528);
or U2100 (N_2100,N_364,N_26);
and U2101 (N_2101,N_1171,N_361);
nor U2102 (N_2102,N_620,N_1776);
or U2103 (N_2103,N_599,N_1396);
nand U2104 (N_2104,N_1487,N_1699);
nand U2105 (N_2105,N_883,N_660);
and U2106 (N_2106,N_111,N_1923);
xnor U2107 (N_2107,N_407,N_1659);
nand U2108 (N_2108,N_1542,N_272);
nor U2109 (N_2109,N_1287,N_860);
nand U2110 (N_2110,N_885,N_44);
or U2111 (N_2111,N_687,N_1525);
and U2112 (N_2112,N_1739,N_153);
nand U2113 (N_2113,N_193,N_739);
and U2114 (N_2114,N_597,N_766);
xor U2115 (N_2115,N_488,N_656);
or U2116 (N_2116,N_576,N_114);
and U2117 (N_2117,N_74,N_6);
or U2118 (N_2118,N_777,N_1488);
and U2119 (N_2119,N_1433,N_404);
or U2120 (N_2120,N_615,N_1672);
nor U2121 (N_2121,N_1290,N_870);
xor U2122 (N_2122,N_1642,N_1413);
xor U2123 (N_2123,N_1518,N_42);
nor U2124 (N_2124,N_432,N_1834);
nor U2125 (N_2125,N_1403,N_1419);
and U2126 (N_2126,N_1486,N_288);
nand U2127 (N_2127,N_1337,N_526);
or U2128 (N_2128,N_686,N_1070);
nor U2129 (N_2129,N_154,N_1463);
nor U2130 (N_2130,N_1942,N_461);
and U2131 (N_2131,N_1873,N_1384);
and U2132 (N_2132,N_975,N_688);
and U2133 (N_2133,N_1623,N_1954);
and U2134 (N_2134,N_1760,N_251);
nor U2135 (N_2135,N_1059,N_388);
nor U2136 (N_2136,N_530,N_24);
nor U2137 (N_2137,N_822,N_340);
nor U2138 (N_2138,N_983,N_747);
and U2139 (N_2139,N_411,N_1727);
xnor U2140 (N_2140,N_1681,N_1012);
and U2141 (N_2141,N_89,N_1357);
or U2142 (N_2142,N_1908,N_1021);
and U2143 (N_2143,N_668,N_48);
nor U2144 (N_2144,N_1250,N_25);
and U2145 (N_2145,N_909,N_493);
and U2146 (N_2146,N_1514,N_396);
xor U2147 (N_2147,N_1674,N_1949);
and U2148 (N_2148,N_186,N_1852);
nor U2149 (N_2149,N_1995,N_1808);
or U2150 (N_2150,N_992,N_383);
or U2151 (N_2151,N_967,N_1792);
and U2152 (N_2152,N_1838,N_1779);
nand U2153 (N_2153,N_472,N_309);
xnor U2154 (N_2154,N_545,N_1751);
or U2155 (N_2155,N_1851,N_296);
nor U2156 (N_2156,N_1906,N_152);
xor U2157 (N_2157,N_851,N_287);
nand U2158 (N_2158,N_1961,N_1169);
xnor U2159 (N_2159,N_1745,N_1267);
and U2160 (N_2160,N_212,N_1884);
xnor U2161 (N_2161,N_934,N_774);
nor U2162 (N_2162,N_1225,N_0);
or U2163 (N_2163,N_1587,N_1615);
nand U2164 (N_2164,N_643,N_359);
or U2165 (N_2165,N_43,N_324);
nand U2166 (N_2166,N_1340,N_304);
xnor U2167 (N_2167,N_561,N_1277);
nand U2168 (N_2168,N_631,N_199);
or U2169 (N_2169,N_601,N_277);
or U2170 (N_2170,N_103,N_1775);
and U2171 (N_2171,N_1618,N_1666);
nor U2172 (N_2172,N_1014,N_1097);
or U2173 (N_2173,N_462,N_637);
nand U2174 (N_2174,N_594,N_636);
nor U2175 (N_2175,N_1416,N_1969);
nor U2176 (N_2176,N_1188,N_1448);
or U2177 (N_2177,N_1878,N_329);
and U2178 (N_2178,N_1058,N_1686);
nor U2179 (N_2179,N_621,N_1437);
nor U2180 (N_2180,N_1761,N_398);
nor U2181 (N_2181,N_999,N_1670);
or U2182 (N_2182,N_837,N_426);
xnor U2183 (N_2183,N_641,N_107);
or U2184 (N_2184,N_1561,N_1178);
nor U2185 (N_2185,N_79,N_1937);
or U2186 (N_2186,N_1108,N_280);
and U2187 (N_2187,N_311,N_93);
and U2188 (N_2188,N_497,N_802);
nand U2189 (N_2189,N_122,N_227);
nand U2190 (N_2190,N_240,N_1471);
and U2191 (N_2191,N_69,N_920);
nand U2192 (N_2192,N_421,N_1067);
and U2193 (N_2193,N_368,N_742);
nor U2194 (N_2194,N_166,N_788);
or U2195 (N_2195,N_1797,N_1511);
or U2196 (N_2196,N_804,N_1033);
and U2197 (N_2197,N_1719,N_640);
or U2198 (N_2198,N_333,N_959);
and U2199 (N_2199,N_1015,N_832);
nor U2200 (N_2200,N_21,N_1093);
nand U2201 (N_2201,N_197,N_428);
and U2202 (N_2202,N_1904,N_816);
or U2203 (N_2203,N_413,N_546);
nor U2204 (N_2204,N_1028,N_419);
or U2205 (N_2205,N_1372,N_1636);
nand U2206 (N_2206,N_161,N_741);
nand U2207 (N_2207,N_1717,N_1105);
nand U2208 (N_2208,N_163,N_1643);
nor U2209 (N_2209,N_290,N_1722);
or U2210 (N_2210,N_1075,N_1546);
or U2211 (N_2211,N_1701,N_976);
nor U2212 (N_2212,N_1343,N_417);
xor U2213 (N_2213,N_765,N_1427);
nor U2214 (N_2214,N_572,N_1212);
nor U2215 (N_2215,N_276,N_457);
and U2216 (N_2216,N_1687,N_1163);
and U2217 (N_2217,N_1072,N_230);
or U2218 (N_2218,N_1902,N_243);
nor U2219 (N_2219,N_265,N_125);
and U2220 (N_2220,N_612,N_1832);
and U2221 (N_2221,N_841,N_134);
nand U2222 (N_2222,N_1513,N_1263);
xor U2223 (N_2223,N_833,N_459);
and U2224 (N_2224,N_1462,N_618);
nor U2225 (N_2225,N_165,N_144);
nand U2226 (N_2226,N_1046,N_779);
and U2227 (N_2227,N_715,N_1605);
nand U2228 (N_2228,N_1262,N_1359);
nor U2229 (N_2229,N_377,N_1226);
nand U2230 (N_2230,N_1069,N_634);
nor U2231 (N_2231,N_1063,N_1383);
nand U2232 (N_2232,N_349,N_1754);
xor U2233 (N_2233,N_1925,N_1794);
or U2234 (N_2234,N_360,N_956);
and U2235 (N_2235,N_916,N_1252);
or U2236 (N_2236,N_1202,N_1266);
xor U2237 (N_2237,N_843,N_724);
nand U2238 (N_2238,N_1648,N_964);
and U2239 (N_2239,N_1096,N_1723);
or U2240 (N_2240,N_84,N_915);
or U2241 (N_2241,N_221,N_370);
nor U2242 (N_2242,N_1270,N_27);
or U2243 (N_2243,N_1426,N_483);
and U2244 (N_2244,N_1522,N_1634);
xor U2245 (N_2245,N_1442,N_1752);
and U2246 (N_2246,N_61,N_527);
nand U2247 (N_2247,N_538,N_881);
or U2248 (N_2248,N_449,N_1496);
nor U2249 (N_2249,N_1977,N_1978);
xnor U2250 (N_2250,N_1692,N_1568);
and U2251 (N_2251,N_1633,N_1799);
nand U2252 (N_2252,N_171,N_1493);
xnor U2253 (N_2253,N_550,N_681);
nand U2254 (N_2254,N_356,N_242);
nand U2255 (N_2255,N_993,N_362);
nand U2256 (N_2256,N_1247,N_196);
and U2257 (N_2257,N_1690,N_1933);
and U2258 (N_2258,N_1502,N_1339);
nand U2259 (N_2259,N_1235,N_1510);
nor U2260 (N_2260,N_1531,N_695);
or U2261 (N_2261,N_1104,N_672);
nand U2262 (N_2262,N_745,N_824);
and U2263 (N_2263,N_1470,N_312);
or U2264 (N_2264,N_1915,N_1616);
or U2265 (N_2265,N_1305,N_1393);
nand U2266 (N_2266,N_539,N_502);
or U2267 (N_2267,N_1612,N_577);
and U2268 (N_2268,N_1210,N_1620);
and U2269 (N_2269,N_1946,N_75);
and U2270 (N_2270,N_1482,N_444);
xnor U2271 (N_2271,N_205,N_50);
xnor U2272 (N_2272,N_1785,N_580);
xor U2273 (N_2273,N_1334,N_1092);
and U2274 (N_2274,N_467,N_773);
and U2275 (N_2275,N_351,N_293);
nor U2276 (N_2276,N_68,N_923);
nor U2277 (N_2277,N_1736,N_1845);
nor U2278 (N_2278,N_1519,N_1807);
or U2279 (N_2279,N_1564,N_143);
and U2280 (N_2280,N_1229,N_71);
or U2281 (N_2281,N_1815,N_718);
nand U2282 (N_2282,N_571,N_924);
or U2283 (N_2283,N_1999,N_305);
nor U2284 (N_2284,N_725,N_127);
xor U2285 (N_2285,N_799,N_1888);
or U2286 (N_2286,N_1947,N_1386);
nor U2287 (N_2287,N_596,N_292);
and U2288 (N_2288,N_129,N_1816);
or U2289 (N_2289,N_1865,N_590);
or U2290 (N_2290,N_584,N_301);
and U2291 (N_2291,N_323,N_274);
nor U2292 (N_2292,N_917,N_1243);
nor U2293 (N_2293,N_1557,N_229);
and U2294 (N_2294,N_512,N_1166);
or U2295 (N_2295,N_524,N_1483);
and U2296 (N_2296,N_1134,N_198);
or U2297 (N_2297,N_877,N_1051);
or U2298 (N_2298,N_11,N_605);
nand U2299 (N_2299,N_116,N_1899);
xnor U2300 (N_2300,N_1205,N_768);
nor U2301 (N_2301,N_1732,N_1452);
nor U2302 (N_2302,N_1191,N_880);
xor U2303 (N_2303,N_138,N_1830);
nand U2304 (N_2304,N_158,N_679);
or U2305 (N_2305,N_1881,N_948);
nor U2306 (N_2306,N_1302,N_1221);
and U2307 (N_2307,N_1868,N_507);
xnor U2308 (N_2308,N_961,N_1753);
nand U2309 (N_2309,N_142,N_73);
nand U2310 (N_2310,N_1661,N_874);
nor U2311 (N_2311,N_300,N_1897);
and U2312 (N_2312,N_393,N_1321);
nand U2313 (N_2313,N_800,N_719);
xor U2314 (N_2314,N_267,N_1351);
and U2315 (N_2315,N_446,N_1590);
and U2316 (N_2316,N_1121,N_790);
nand U2317 (N_2317,N_439,N_217);
nor U2318 (N_2318,N_128,N_1354);
and U2319 (N_2319,N_1668,N_1325);
xnor U2320 (N_2320,N_1200,N_1280);
or U2321 (N_2321,N_1209,N_1820);
xnor U2322 (N_2322,N_1715,N_1926);
and U2323 (N_2323,N_906,N_1466);
and U2324 (N_2324,N_1074,N_1869);
nand U2325 (N_2325,N_34,N_565);
or U2326 (N_2326,N_1391,N_416);
and U2327 (N_2327,N_126,N_783);
or U2328 (N_2328,N_1856,N_1697);
nor U2329 (N_2329,N_556,N_1936);
nor U2330 (N_2330,N_1465,N_381);
nand U2331 (N_2331,N_873,N_1958);
nor U2332 (N_2332,N_37,N_131);
nand U2333 (N_2333,N_1927,N_1602);
nor U2334 (N_2334,N_1653,N_776);
nor U2335 (N_2335,N_336,N_1700);
nor U2336 (N_2336,N_893,N_1430);
nand U2337 (N_2337,N_908,N_1197);
xor U2338 (N_2338,N_913,N_1757);
or U2339 (N_2339,N_391,N_1490);
nand U2340 (N_2340,N_187,N_1447);
nand U2341 (N_2341,N_847,N_1309);
or U2342 (N_2342,N_448,N_140);
xnor U2343 (N_2343,N_1503,N_1147);
xor U2344 (N_2344,N_216,N_1728);
and U2345 (N_2345,N_1812,N_757);
nor U2346 (N_2346,N_1957,N_844);
xnor U2347 (N_2347,N_1972,N_926);
and U2348 (N_2348,N_1161,N_460);
nor U2349 (N_2349,N_90,N_1068);
nand U2350 (N_2350,N_865,N_476);
and U2351 (N_2351,N_1573,N_1232);
nand U2352 (N_2352,N_1026,N_1931);
nor U2353 (N_2353,N_1165,N_1101);
nand U2354 (N_2354,N_1842,N_1030);
nor U2355 (N_2355,N_1547,N_1464);
nand U2356 (N_2356,N_261,N_1025);
xor U2357 (N_2357,N_1190,N_256);
nor U2358 (N_2358,N_425,N_245);
nor U2359 (N_2359,N_736,N_1491);
nor U2360 (N_2360,N_1932,N_1342);
and U2361 (N_2361,N_307,N_500);
or U2362 (N_2362,N_1017,N_1246);
nor U2363 (N_2363,N_1789,N_224);
nand U2364 (N_2364,N_1045,N_147);
nor U2365 (N_2365,N_470,N_1008);
xnor U2366 (N_2366,N_1278,N_1712);
xor U2367 (N_2367,N_1392,N_1819);
xnor U2368 (N_2368,N_1311,N_1604);
and U2369 (N_2369,N_156,N_234);
nand U2370 (N_2370,N_495,N_1504);
and U2371 (N_2371,N_289,N_884);
and U2372 (N_2372,N_1095,N_657);
or U2373 (N_2373,N_722,N_1721);
nand U2374 (N_2374,N_271,N_587);
nand U2375 (N_2375,N_1850,N_1976);
or U2376 (N_2376,N_1253,N_1611);
and U2377 (N_2377,N_347,N_753);
and U2378 (N_2378,N_1900,N_132);
nor U2379 (N_2379,N_1408,N_914);
nand U2380 (N_2380,N_1939,N_864);
nor U2381 (N_2381,N_1421,N_1242);
and U2382 (N_2382,N_750,N_1762);
nand U2383 (N_2383,N_331,N_1175);
xor U2384 (N_2384,N_45,N_1508);
and U2385 (N_2385,N_1296,N_1551);
and U2386 (N_2386,N_905,N_731);
nand U2387 (N_2387,N_22,N_1187);
xnor U2388 (N_2388,N_392,N_809);
and U2389 (N_2389,N_1474,N_1373);
and U2390 (N_2390,N_1454,N_573);
and U2391 (N_2391,N_395,N_775);
and U2392 (N_2392,N_1580,N_386);
nor U2393 (N_2393,N_1185,N_1562);
or U2394 (N_2394,N_886,N_644);
and U2395 (N_2395,N_475,N_1887);
and U2396 (N_2396,N_1679,N_478);
nor U2397 (N_2397,N_1120,N_246);
nor U2398 (N_2398,N_1432,N_1206);
and U2399 (N_2399,N_897,N_452);
xnor U2400 (N_2400,N_378,N_249);
nand U2401 (N_2401,N_178,N_551);
xnor U2402 (N_2402,N_958,N_1627);
xnor U2403 (N_2403,N_1239,N_1159);
nor U2404 (N_2404,N_738,N_1769);
or U2405 (N_2405,N_1153,N_1137);
nand U2406 (N_2406,N_1824,N_1554);
nor U2407 (N_2407,N_1521,N_808);
nor U2408 (N_2408,N_353,N_1128);
and U2409 (N_2409,N_443,N_996);
or U2410 (N_2410,N_986,N_898);
and U2411 (N_2411,N_1965,N_1222);
xor U2412 (N_2412,N_582,N_1505);
and U2413 (N_2413,N_1130,N_1730);
nand U2414 (N_2414,N_1705,N_397);
and U2415 (N_2415,N_690,N_1533);
nand U2416 (N_2416,N_1920,N_1414);
nor U2417 (N_2417,N_1889,N_308);
and U2418 (N_2418,N_876,N_1609);
nor U2419 (N_2419,N_56,N_1827);
or U2420 (N_2420,N_208,N_52);
nor U2421 (N_2421,N_570,N_685);
nand U2422 (N_2422,N_1800,N_568);
nor U2423 (N_2423,N_433,N_47);
or U2424 (N_2424,N_1553,N_1282);
or U2425 (N_2425,N_1938,N_1795);
nor U2426 (N_2426,N_1307,N_1327);
nor U2427 (N_2427,N_318,N_1858);
nor U2428 (N_2428,N_521,N_1467);
and U2429 (N_2429,N_1081,N_339);
nand U2430 (N_2430,N_814,N_367);
and U2431 (N_2431,N_162,N_1928);
nand U2432 (N_2432,N_925,N_30);
nand U2433 (N_2433,N_499,N_994);
nand U2434 (N_2434,N_1640,N_379);
or U2435 (N_2435,N_321,N_49);
or U2436 (N_2436,N_1787,N_858);
nor U2437 (N_2437,N_1485,N_1086);
nand U2438 (N_2438,N_283,N_257);
or U2439 (N_2439,N_1288,N_469);
and U2440 (N_2440,N_1407,N_1365);
nand U2441 (N_2441,N_602,N_1993);
or U2442 (N_2442,N_1967,N_1767);
nand U2443 (N_2443,N_737,N_1929);
and U2444 (N_2444,N_784,N_1556);
nor U2445 (N_2445,N_41,N_1338);
nor U2446 (N_2446,N_326,N_1515);
or U2447 (N_2447,N_1136,N_3);
or U2448 (N_2448,N_659,N_1772);
nand U2449 (N_2449,N_180,N_429);
or U2450 (N_2450,N_705,N_648);
or U2451 (N_2451,N_1335,N_358);
or U2452 (N_2452,N_1763,N_1898);
and U2453 (N_2453,N_1355,N_693);
or U2454 (N_2454,N_871,N_1224);
or U2455 (N_2455,N_1315,N_441);
nand U2456 (N_2456,N_1424,N_64);
xnor U2457 (N_2457,N_314,N_899);
and U2458 (N_2458,N_1652,N_167);
and U2459 (N_2459,N_791,N_1099);
and U2460 (N_2460,N_1901,N_303);
nand U2461 (N_2461,N_1657,N_555);
nand U2462 (N_2462,N_1650,N_1249);
or U2463 (N_2463,N_929,N_623);
or U2464 (N_2464,N_1118,N_523);
or U2465 (N_2465,N_1991,N_1286);
nor U2466 (N_2466,N_567,N_485);
nor U2467 (N_2467,N_836,N_215);
nor U2468 (N_2468,N_1874,N_1143);
and U2469 (N_2469,N_1945,N_5);
nand U2470 (N_2470,N_1597,N_1645);
nand U2471 (N_2471,N_1179,N_1524);
nor U2472 (N_2472,N_1294,N_664);
and U2473 (N_2473,N_991,N_1150);
nand U2474 (N_2474,N_1085,N_1608);
nor U2475 (N_2475,N_1078,N_23);
xor U2476 (N_2476,N_746,N_1741);
nand U2477 (N_2477,N_172,N_1671);
and U2478 (N_2478,N_1420,N_486);
nor U2479 (N_2479,N_270,N_59);
nor U2480 (N_2480,N_795,N_1731);
and U2481 (N_2481,N_888,N_92);
nand U2482 (N_2482,N_529,N_984);
or U2483 (N_2483,N_709,N_1916);
and U2484 (N_2484,N_464,N_262);
nand U2485 (N_2485,N_412,N_857);
nor U2486 (N_2486,N_740,N_62);
nor U2487 (N_2487,N_1541,N_447);
and U2488 (N_2488,N_1848,N_813);
or U2489 (N_2489,N_988,N_1771);
and U2490 (N_2490,N_1479,N_1859);
or U2491 (N_2491,N_531,N_855);
xor U2492 (N_2492,N_829,N_279);
nand U2493 (N_2493,N_667,N_734);
nor U2494 (N_2494,N_581,N_1796);
nand U2495 (N_2495,N_14,N_1177);
nor U2496 (N_2496,N_214,N_1151);
nand U2497 (N_2497,N_540,N_82);
nand U2498 (N_2498,N_951,N_453);
nand U2499 (N_2499,N_51,N_319);
nor U2500 (N_2500,N_985,N_626);
nor U2501 (N_2501,N_427,N_496);
or U2502 (N_2502,N_701,N_1698);
and U2503 (N_2503,N_1116,N_1501);
nand U2504 (N_2504,N_604,N_1011);
and U2505 (N_2505,N_1052,N_1406);
or U2506 (N_2506,N_1411,N_87);
nand U2507 (N_2507,N_517,N_1495);
xor U2508 (N_2508,N_919,N_730);
nor U2509 (N_2509,N_1737,N_320);
nor U2510 (N_2510,N_941,N_1537);
or U2511 (N_2511,N_1649,N_889);
nor U2512 (N_2512,N_633,N_1622);
or U2513 (N_2513,N_474,N_1861);
or U2514 (N_2514,N_297,N_1057);
nand U2515 (N_2515,N_1245,N_204);
or U2516 (N_2516,N_1548,N_431);
nor U2517 (N_2517,N_181,N_1704);
nand U2518 (N_2518,N_1512,N_1663);
and U2519 (N_2519,N_1990,N_518);
and U2520 (N_2520,N_1186,N_603);
xor U2521 (N_2521,N_1441,N_1429);
nor U2522 (N_2522,N_110,N_1055);
and U2523 (N_2523,N_1003,N_55);
and U2524 (N_2524,N_284,N_1532);
and U2525 (N_2525,N_838,N_1720);
or U2526 (N_2526,N_481,N_585);
or U2527 (N_2527,N_1457,N_1292);
nand U2528 (N_2528,N_159,N_1768);
nand U2529 (N_2529,N_1835,N_1639);
nor U2530 (N_2530,N_169,N_1313);
nand U2531 (N_2531,N_65,N_1973);
or U2532 (N_2532,N_1825,N_706);
nand U2533 (N_2533,N_1638,N_1048);
nor U2534 (N_2534,N_1228,N_1366);
nor U2535 (N_2535,N_1922,N_1475);
and U2536 (N_2536,N_1376,N_442);
nand U2537 (N_2537,N_595,N_375);
nor U2538 (N_2538,N_420,N_1007);
nand U2539 (N_2539,N_927,N_1912);
and U2540 (N_2540,N_1738,N_81);
or U2541 (N_2541,N_1469,N_952);
and U2542 (N_2542,N_1535,N_468);
and U2543 (N_2543,N_1765,N_1318);
nand U2544 (N_2544,N_772,N_135);
nor U2545 (N_2545,N_1436,N_1023);
and U2546 (N_2546,N_970,N_894);
or U2547 (N_2547,N_1195,N_818);
nor U2548 (N_2548,N_9,N_1822);
nor U2549 (N_2549,N_756,N_535);
or U2550 (N_2550,N_1654,N_1581);
nand U2551 (N_2551,N_1237,N_1886);
nand U2552 (N_2552,N_1455,N_542);
nand U2553 (N_2553,N_189,N_1039);
nand U2554 (N_2554,N_1155,N_939);
nand U2555 (N_2555,N_717,N_1084);
or U2556 (N_2556,N_671,N_879);
nand U2557 (N_2557,N_801,N_281);
nor U2558 (N_2558,N_1836,N_473);
nor U2559 (N_2559,N_1378,N_1127);
or U2560 (N_2560,N_825,N_414);
nand U2561 (N_2561,N_781,N_133);
nand U2562 (N_2562,N_1924,N_998);
nor U2563 (N_2563,N_1135,N_978);
nand U2564 (N_2564,N_1952,N_291);
nand U2565 (N_2565,N_831,N_1154);
nor U2566 (N_2566,N_911,N_1809);
or U2567 (N_2567,N_385,N_763);
nand U2568 (N_2568,N_1098,N_1324);
nor U2569 (N_2569,N_760,N_1823);
nor U2570 (N_2570,N_350,N_2);
and U2571 (N_2571,N_1673,N_210);
or U2572 (N_2572,N_1711,N_1905);
nor U2573 (N_2573,N_513,N_1415);
nor U2574 (N_2574,N_60,N_173);
xnor U2575 (N_2575,N_558,N_946);
nand U2576 (N_2576,N_409,N_697);
nand U2577 (N_2577,N_299,N_1259);
nand U2578 (N_2578,N_1329,N_98);
and U2579 (N_2579,N_1203,N_780);
and U2580 (N_2580,N_211,N_1103);
or U2581 (N_2581,N_1667,N_1276);
xnor U2582 (N_2582,N_1658,N_528);
and U2583 (N_2583,N_102,N_237);
or U2584 (N_2584,N_617,N_1241);
and U2585 (N_2585,N_583,N_1369);
or U2586 (N_2586,N_1102,N_1813);
nand U2587 (N_2587,N_1230,N_1941);
or U2588 (N_2588,N_830,N_525);
or U2589 (N_2589,N_184,N_1603);
or U2590 (N_2590,N_1132,N_1506);
nor U2591 (N_2591,N_139,N_1544);
nand U2592 (N_2592,N_1035,N_1911);
xor U2593 (N_2593,N_337,N_1087);
and U2594 (N_2594,N_1569,N_862);
xor U2595 (N_2595,N_223,N_248);
and U2596 (N_2596,N_136,N_1631);
nand U2597 (N_2597,N_653,N_895);
or U2598 (N_2598,N_1268,N_1451);
and U2599 (N_2599,N_405,N_1211);
nor U2600 (N_2600,N_1892,N_151);
or U2601 (N_2601,N_53,N_1002);
nand U2602 (N_2602,N_1540,N_1559);
nor U2603 (N_2603,N_651,N_1837);
and U2604 (N_2604,N_933,N_1598);
xor U2605 (N_2605,N_1526,N_1709);
xnor U2606 (N_2606,N_406,N_646);
nand U2607 (N_2607,N_1803,N_1412);
xor U2608 (N_2608,N_1100,N_1422);
or U2609 (N_2609,N_616,N_1867);
and U2610 (N_2610,N_1390,N_815);
xnor U2611 (N_2611,N_907,N_900);
or U2612 (N_2612,N_645,N_1759);
nand U2613 (N_2613,N_95,N_859);
nand U2614 (N_2614,N_1840,N_1893);
or U2615 (N_2615,N_826,N_1997);
and U2616 (N_2616,N_1193,N_213);
nor U2617 (N_2617,N_1382,N_1090);
nand U2618 (N_2618,N_185,N_105);
and U2619 (N_2619,N_1336,N_120);
nor U2620 (N_2620,N_1385,N_209);
and U2621 (N_2621,N_1449,N_1782);
nor U2622 (N_2622,N_1181,N_113);
or U2623 (N_2623,N_654,N_255);
nand U2624 (N_2624,N_1065,N_315);
nor U2625 (N_2625,N_692,N_1713);
and U2626 (N_2626,N_578,N_1400);
and U2627 (N_2627,N_1788,N_1979);
nand U2628 (N_2628,N_1299,N_839);
or U2629 (N_2629,N_785,N_1356);
xor U2630 (N_2630,N_1094,N_1742);
or U2631 (N_2631,N_503,N_332);
nand U2632 (N_2632,N_942,N_980);
and U2633 (N_2633,N_1624,N_440);
and U2634 (N_2634,N_346,N_1810);
or U2635 (N_2635,N_1647,N_997);
xnor U2636 (N_2636,N_767,N_1585);
and U2637 (N_2637,N_786,N_1481);
and U2638 (N_2638,N_1428,N_1921);
or U2639 (N_2639,N_1944,N_1423);
or U2640 (N_2640,N_1748,N_1853);
nand U2641 (N_2641,N_1706,N_850);
nand U2642 (N_2642,N_1164,N_1213);
or U2643 (N_2643,N_793,N_1814);
nand U2644 (N_2644,N_1839,N_1935);
xor U2645 (N_2645,N_828,N_1646);
and U2646 (N_2646,N_762,N_275);
and U2647 (N_2647,N_399,N_674);
and U2648 (N_2648,N_57,N_680);
and U2649 (N_2649,N_1934,N_1204);
and U2650 (N_2650,N_344,N_1798);
nand U2651 (N_2651,N_1907,N_1691);
or U2652 (N_2652,N_1275,N_1499);
nand U2653 (N_2653,N_78,N_1142);
and U2654 (N_2654,N_1144,N_1117);
or U2655 (N_2655,N_1708,N_1801);
xnor U2656 (N_2656,N_1994,N_1478);
and U2657 (N_2657,N_1534,N_749);
or U2658 (N_2658,N_1182,N_1284);
and U2659 (N_2659,N_728,N_591);
and U2660 (N_2660,N_938,N_1285);
or U2661 (N_2661,N_480,N_684);
nand U2662 (N_2662,N_536,N_607);
xor U2663 (N_2663,N_1009,N_376);
and U2664 (N_2664,N_1326,N_1628);
nor U2665 (N_2665,N_533,N_953);
nor U2666 (N_2666,N_273,N_164);
nor U2667 (N_2667,N_1260,N_1207);
nor U2668 (N_2668,N_1218,N_658);
and U2669 (N_2669,N_1214,N_1332);
nand U2670 (N_2670,N_678,N_1353);
or U2671 (N_2671,N_666,N_1744);
nor U2672 (N_2672,N_823,N_1484);
and U2673 (N_2673,N_1773,N_922);
and U2674 (N_2674,N_1790,N_1849);
or U2675 (N_2675,N_1930,N_1955);
or U2676 (N_2676,N_1037,N_673);
nor U2677 (N_2677,N_435,N_236);
or U2678 (N_2678,N_1109,N_1053);
or U2679 (N_2679,N_380,N_316);
nor U2680 (N_2680,N_649,N_1140);
nor U2681 (N_2681,N_1662,N_1555);
nand U2682 (N_2682,N_973,N_1368);
nor U2683 (N_2683,N_1688,N_13);
or U2684 (N_2684,N_190,N_1606);
or U2685 (N_2685,N_195,N_121);
and U2686 (N_2686,N_940,N_1971);
or U2687 (N_2687,N_1138,N_714);
xnor U2688 (N_2688,N_17,N_1707);
and U2689 (N_2689,N_94,N_1310);
nor U2690 (N_2690,N_635,N_29);
nand U2691 (N_2691,N_504,N_1545);
xnor U2692 (N_2692,N_1217,N_1877);
nand U2693 (N_2693,N_1950,N_206);
and U2694 (N_2694,N_764,N_341);
and U2695 (N_2695,N_455,N_1388);
and U2696 (N_2696,N_1621,N_15);
or U2697 (N_2697,N_629,N_510);
and U2698 (N_2698,N_990,N_325);
nand U2699 (N_2699,N_912,N_803);
xor U2700 (N_2700,N_1476,N_1347);
nor U2701 (N_2701,N_1122,N_935);
and U2702 (N_2702,N_1111,N_191);
and U2703 (N_2703,N_1871,N_403);
nor U2704 (N_2704,N_1231,N_733);
nor U2705 (N_2705,N_703,N_1196);
nor U2706 (N_2706,N_20,N_1459);
or U2707 (N_2707,N_1446,N_744);
nor U2708 (N_2708,N_1360,N_560);
and U2709 (N_2709,N_1817,N_759);
nor U2710 (N_2710,N_1517,N_1317);
or U2711 (N_2711,N_1872,N_543);
nand U2712 (N_2712,N_268,N_1112);
nand U2713 (N_2713,N_532,N_853);
and U2714 (N_2714,N_1962,N_1507);
or U2715 (N_2715,N_727,N_1119);
xnor U2716 (N_2716,N_1780,N_389);
nand U2717 (N_2717,N_1880,N_511);
xor U2718 (N_2718,N_1402,N_1027);
and U2719 (N_2719,N_1576,N_856);
nand U2720 (N_2720,N_1272,N_566);
xor U2721 (N_2721,N_1703,N_1060);
and U2722 (N_2722,N_250,N_1963);
nor U2723 (N_2723,N_1445,N_751);
nor U2724 (N_2724,N_1201,N_866);
or U2725 (N_2725,N_282,N_1375);
nand U2726 (N_2726,N_1637,N_1083);
xnor U2727 (N_2727,N_1783,N_99);
nand U2728 (N_2728,N_157,N_1367);
nor U2729 (N_2729,N_1714,N_423);
or U2730 (N_2730,N_609,N_1040);
nand U2731 (N_2731,N_944,N_1073);
or U2732 (N_2732,N_1149,N_1300);
and U2733 (N_2733,N_1583,N_101);
nor U2734 (N_2734,N_875,N_516);
and U2735 (N_2735,N_1778,N_28);
or U2736 (N_2736,N_363,N_1781);
nor U2737 (N_2737,N_704,N_1600);
and U2738 (N_2738,N_1001,N_1953);
nand U2739 (N_2739,N_1725,N_798);
nand U2740 (N_2740,N_610,N_1956);
nand U2741 (N_2741,N_960,N_812);
nand U2742 (N_2742,N_1543,N_868);
and U2743 (N_2743,N_1656,N_264);
nor U2744 (N_2744,N_1071,N_854);
nand U2745 (N_2745,N_244,N_910);
or U2746 (N_2746,N_232,N_1198);
and U2747 (N_2747,N_1344,N_145);
or U2748 (N_2748,N_1018,N_608);
nand U2749 (N_2749,N_36,N_937);
and U2750 (N_2750,N_987,N_72);
nor U2751 (N_2751,N_1192,N_400);
xnor U2752 (N_2752,N_1295,N_743);
nor U2753 (N_2753,N_505,N_313);
and U2754 (N_2754,N_1107,N_638);
nand U2755 (N_2755,N_969,N_662);
and U2756 (N_2756,N_1843,N_33);
or U2757 (N_2757,N_1626,N_437);
or U2758 (N_2758,N_1538,N_792);
nor U2759 (N_2759,N_1434,N_1435);
nand U2760 (N_2760,N_771,N_1695);
nand U2761 (N_2761,N_1401,N_1625);
or U2762 (N_2762,N_1077,N_1750);
nor U2763 (N_2763,N_537,N_1167);
nor U2764 (N_2764,N_1669,N_31);
and U2765 (N_2765,N_1473,N_35);
nand U2766 (N_2766,N_1805,N_1133);
nor U2767 (N_2767,N_541,N_302);
or U2768 (N_2768,N_1141,N_1896);
nand U2769 (N_2769,N_177,N_327);
and U2770 (N_2770,N_477,N_515);
nor U2771 (N_2771,N_827,N_1380);
nand U2772 (N_2772,N_1131,N_371);
or U2773 (N_2773,N_1894,N_1755);
xor U2774 (N_2774,N_867,N_1062);
and U2775 (N_2775,N_811,N_834);
nand U2776 (N_2776,N_1461,N_451);
xnor U2777 (N_2777,N_1875,N_175);
and U2778 (N_2778,N_401,N_1395);
xnor U2779 (N_2779,N_655,N_1860);
xor U2780 (N_2780,N_1079,N_1456);
and U2781 (N_2781,N_1584,N_354);
nor U2782 (N_2782,N_484,N_1574);
nor U2783 (N_2783,N_869,N_1306);
nor U2784 (N_2784,N_1970,N_508);
and U2785 (N_2785,N_963,N_1265);
nor U2786 (N_2786,N_849,N_1236);
nand U2787 (N_2787,N_1523,N_1054);
or U2788 (N_2788,N_1162,N_563);
nor U2789 (N_2789,N_1509,N_238);
nor U2790 (N_2790,N_1988,N_32);
xor U2791 (N_2791,N_650,N_1975);
nor U2792 (N_2792,N_965,N_1599);
nor U2793 (N_2793,N_1806,N_702);
nor U2794 (N_2794,N_1811,N_1350);
and U2795 (N_2795,N_387,N_835);
nand U2796 (N_2796,N_950,N_70);
and U2797 (N_2797,N_1431,N_1909);
or U2798 (N_2798,N_228,N_778);
or U2799 (N_2799,N_1319,N_1497);
and U2800 (N_2800,N_1399,N_1746);
nand U2801 (N_2801,N_1985,N_1322);
or U2802 (N_2802,N_1610,N_520);
nor U2803 (N_2803,N_1578,N_1316);
nand U2804 (N_2804,N_1126,N_1041);
and U2805 (N_2805,N_882,N_1264);
nand U2806 (N_2806,N_357,N_797);
nor U2807 (N_2807,N_1248,N_266);
nand U2808 (N_2808,N_1489,N_1857);
nor U2809 (N_2809,N_1362,N_1364);
and U2810 (N_2810,N_1029,N_1379);
or U2811 (N_2811,N_1,N_1323);
nand U2812 (N_2812,N_97,N_982);
or U2813 (N_2813,N_691,N_123);
nand U2814 (N_2814,N_1044,N_1261);
xor U2815 (N_2815,N_1913,N_968);
or U2816 (N_2816,N_1183,N_85);
nand U2817 (N_2817,N_966,N_489);
nor U2818 (N_2818,N_663,N_1145);
nand U2819 (N_2819,N_1494,N_726);
nor U2820 (N_2820,N_479,N_1689);
and U2821 (N_2821,N_1031,N_233);
nand U2822 (N_2822,N_1740,N_254);
xor U2823 (N_2823,N_1998,N_1199);
and U2824 (N_2824,N_149,N_160);
or U2825 (N_2825,N_1472,N_1863);
or U2826 (N_2826,N_661,N_1630);
nand U2827 (N_2827,N_501,N_295);
and U2828 (N_2828,N_1733,N_345);
or U2829 (N_2829,N_1238,N_1758);
nor U2830 (N_2830,N_921,N_1890);
xnor U2831 (N_2831,N_487,N_677);
xnor U2832 (N_2832,N_7,N_207);
and U2833 (N_2833,N_758,N_1891);
and U2834 (N_2834,N_1864,N_203);
or U2835 (N_2835,N_720,N_977);
and U2836 (N_2836,N_1734,N_1885);
and U2837 (N_2837,N_1333,N_1696);
or U2838 (N_2838,N_1320,N_1826);
or U2839 (N_2839,N_1234,N_821);
xnor U2840 (N_2840,N_789,N_1283);
nand U2841 (N_2841,N_1492,N_1593);
xor U2842 (N_2842,N_8,N_1289);
nand U2843 (N_2843,N_1601,N_1274);
and U2844 (N_2844,N_330,N_1409);
nand U2845 (N_2845,N_76,N_1047);
or U2846 (N_2846,N_769,N_1034);
xor U2847 (N_2847,N_1951,N_1591);
nor U2848 (N_2848,N_755,N_112);
xor U2849 (N_2849,N_1443,N_96);
nor U2850 (N_2850,N_716,N_682);
nand U2851 (N_2851,N_1082,N_4);
nor U2852 (N_2852,N_863,N_1571);
nor U2853 (N_2853,N_259,N_1529);
nor U2854 (N_2854,N_1349,N_1394);
and U2855 (N_2855,N_611,N_1756);
nor U2856 (N_2856,N_86,N_88);
nand U2857 (N_2857,N_1398,N_632);
nand U2858 (N_2858,N_1879,N_91);
nor U2859 (N_2859,N_382,N_1258);
and U2860 (N_2860,N_600,N_1964);
nor U2861 (N_2861,N_1572,N_372);
and U2862 (N_2862,N_787,N_183);
nor U2863 (N_2863,N_491,N_1629);
or U2864 (N_2864,N_1038,N_698);
or U2865 (N_2865,N_83,N_1743);
nand U2866 (N_2866,N_1215,N_840);
nor U2867 (N_2867,N_1006,N_949);
nand U2868 (N_2868,N_1139,N_652);
nor U2869 (N_2869,N_1174,N_1361);
nand U2870 (N_2870,N_322,N_846);
nor U2871 (N_2871,N_713,N_260);
nor U2872 (N_2872,N_932,N_328);
and U2873 (N_2873,N_1303,N_46);
nor U2874 (N_2874,N_1917,N_1982);
nand U2875 (N_2875,N_1678,N_1173);
nor U2876 (N_2876,N_1870,N_1281);
xnor U2877 (N_2877,N_1257,N_269);
and U2878 (N_2878,N_366,N_106);
or U2879 (N_2879,N_557,N_711);
or U2880 (N_2880,N_552,N_1061);
or U2881 (N_2881,N_471,N_1651);
nand U2882 (N_2882,N_1219,N_1387);
and U2883 (N_2883,N_904,N_696);
or U2884 (N_2884,N_118,N_592);
nor U2885 (N_2885,N_1986,N_220);
and U2886 (N_2886,N_1024,N_100);
nor U2887 (N_2887,N_547,N_1363);
nand U2888 (N_2888,N_1468,N_1004);
and U2889 (N_2889,N_1439,N_374);
nand U2890 (N_2890,N_1552,N_1677);
and U2891 (N_2891,N_890,N_1269);
nand U2892 (N_2892,N_1348,N_1244);
nor U2893 (N_2893,N_694,N_554);
and U2894 (N_2894,N_981,N_1903);
nand U2895 (N_2895,N_1358,N_979);
and U2896 (N_2896,N_1589,N_1066);
nor U2897 (N_2897,N_1110,N_861);
and U2898 (N_2898,N_1984,N_1735);
nor U2899 (N_2899,N_642,N_1123);
nand U2900 (N_2900,N_930,N_1527);
and U2901 (N_2901,N_1655,N_482);
nand U2902 (N_2902,N_647,N_342);
nand U2903 (N_2903,N_285,N_817);
nand U2904 (N_2904,N_1500,N_1114);
nand U2905 (N_2905,N_418,N_989);
nand U2906 (N_2906,N_410,N_1458);
and U2907 (N_2907,N_1220,N_235);
xnor U2908 (N_2908,N_1989,N_194);
or U2909 (N_2909,N_1304,N_218);
nor U2910 (N_2910,N_1983,N_1000);
and U2911 (N_2911,N_343,N_729);
and U2912 (N_2912,N_1227,N_176);
or U2913 (N_2913,N_1948,N_1170);
nand U2914 (N_2914,N_700,N_1567);
and U2915 (N_2915,N_936,N_1418);
and U2916 (N_2916,N_770,N_1389);
or U2917 (N_2917,N_1397,N_1146);
and U2918 (N_2918,N_222,N_1301);
nand U2919 (N_2919,N_1981,N_624);
and U2920 (N_2920,N_1520,N_1330);
and U2921 (N_2921,N_1345,N_454);
nand U2922 (N_2922,N_1582,N_1575);
nand U2923 (N_2923,N_1293,N_1279);
xnor U2924 (N_2924,N_928,N_1862);
nand U2925 (N_2925,N_918,N_168);
and U2926 (N_2926,N_373,N_598);
xor U2927 (N_2927,N_1918,N_317);
or U2928 (N_2928,N_1594,N_1595);
nand U2929 (N_2929,N_365,N_1022);
and U2930 (N_2930,N_931,N_434);
nand U2931 (N_2931,N_1818,N_669);
nand U2932 (N_2932,N_1724,N_1453);
nand U2933 (N_2933,N_842,N_1056);
nand U2934 (N_2934,N_1444,N_1676);
nand U2935 (N_2935,N_1854,N_947);
and U2936 (N_2936,N_1050,N_430);
or U2937 (N_2937,N_1766,N_586);
nor U2938 (N_2938,N_1291,N_1539);
nand U2939 (N_2939,N_625,N_1352);
nand U2940 (N_2940,N_1764,N_463);
nand U2941 (N_2941,N_1710,N_683);
and U2942 (N_2942,N_1968,N_562);
nand U2943 (N_2943,N_1148,N_1828);
or U2944 (N_2944,N_424,N_796);
and U2945 (N_2945,N_63,N_1694);
and U2946 (N_2946,N_754,N_200);
nand U2947 (N_2947,N_548,N_945);
and U2948 (N_2948,N_1036,N_1563);
or U2949 (N_2949,N_1076,N_1381);
nor U2950 (N_2950,N_1438,N_1558);
and U2951 (N_2951,N_415,N_219);
nor U2952 (N_2952,N_1702,N_192);
nor U2953 (N_2953,N_286,N_1189);
xor U2954 (N_2954,N_104,N_174);
nor U2955 (N_2955,N_148,N_670);
and U2956 (N_2956,N_1032,N_954);
nor U2957 (N_2957,N_896,N_887);
nand U2958 (N_2958,N_1477,N_1665);
nor U2959 (N_2959,N_1613,N_1550);
nor U2960 (N_2960,N_957,N_509);
nor U2961 (N_2961,N_676,N_1802);
or U2962 (N_2962,N_1450,N_1680);
and U2963 (N_2963,N_1876,N_852);
and U2964 (N_2964,N_182,N_569);
or U2965 (N_2965,N_1010,N_1251);
and U2966 (N_2966,N_58,N_335);
nand U2967 (N_2967,N_943,N_1042);
and U2968 (N_2968,N_10,N_67);
nand U2969 (N_2969,N_721,N_1208);
or U2970 (N_2970,N_1223,N_639);
or U2971 (N_2971,N_19,N_892);
or U2972 (N_2972,N_1377,N_1565);
nand U2973 (N_2973,N_170,N_1793);
or U2974 (N_2974,N_1614,N_1331);
nor U2975 (N_2975,N_1158,N_1586);
nand U2976 (N_2976,N_492,N_278);
nor U2977 (N_2977,N_1016,N_450);
nor U2978 (N_2978,N_589,N_1417);
or U2979 (N_2979,N_732,N_294);
nor U2980 (N_2980,N_1371,N_1370);
nand U2981 (N_2981,N_310,N_689);
or U2982 (N_2982,N_1124,N_955);
and U2983 (N_2983,N_225,N_1974);
nor U2984 (N_2984,N_150,N_723);
and U2985 (N_2985,N_1644,N_810);
xor U2986 (N_2986,N_761,N_231);
and U2987 (N_2987,N_1682,N_1716);
or U2988 (N_2988,N_1156,N_348);
and U2989 (N_2989,N_820,N_972);
or U2990 (N_2990,N_1596,N_1091);
xor U2991 (N_2991,N_622,N_12);
nor U2992 (N_2992,N_1516,N_903);
or U2993 (N_2993,N_465,N_1729);
or U2994 (N_2994,N_1013,N_54);
nor U2995 (N_2995,N_241,N_675);
and U2996 (N_2996,N_306,N_466);
or U2997 (N_2997,N_117,N_39);
or U2998 (N_2998,N_534,N_1049);
or U2999 (N_2999,N_369,N_1160);
xnor U3000 (N_3000,N_1683,N_411);
and U3001 (N_3001,N_952,N_1313);
or U3002 (N_3002,N_1991,N_489);
or U3003 (N_3003,N_1737,N_614);
xor U3004 (N_3004,N_1148,N_710);
nor U3005 (N_3005,N_475,N_430);
and U3006 (N_3006,N_1540,N_250);
nand U3007 (N_3007,N_141,N_39);
and U3008 (N_3008,N_596,N_1436);
nand U3009 (N_3009,N_1683,N_921);
nand U3010 (N_3010,N_725,N_196);
or U3011 (N_3011,N_1076,N_561);
or U3012 (N_3012,N_1797,N_1600);
nand U3013 (N_3013,N_147,N_1972);
nor U3014 (N_3014,N_1113,N_188);
nor U3015 (N_3015,N_1035,N_1493);
nand U3016 (N_3016,N_1769,N_326);
nor U3017 (N_3017,N_1383,N_894);
and U3018 (N_3018,N_1193,N_1796);
or U3019 (N_3019,N_184,N_1764);
nor U3020 (N_3020,N_1542,N_1996);
xor U3021 (N_3021,N_1507,N_1238);
nand U3022 (N_3022,N_1237,N_585);
or U3023 (N_3023,N_65,N_1165);
or U3024 (N_3024,N_520,N_1248);
nor U3025 (N_3025,N_1008,N_578);
nand U3026 (N_3026,N_41,N_922);
xnor U3027 (N_3027,N_1697,N_1309);
nand U3028 (N_3028,N_1823,N_304);
and U3029 (N_3029,N_1452,N_1796);
xor U3030 (N_3030,N_1726,N_823);
xor U3031 (N_3031,N_1653,N_1304);
and U3032 (N_3032,N_801,N_62);
xor U3033 (N_3033,N_1998,N_958);
nand U3034 (N_3034,N_1145,N_1960);
or U3035 (N_3035,N_1988,N_397);
nor U3036 (N_3036,N_62,N_1415);
xnor U3037 (N_3037,N_52,N_810);
and U3038 (N_3038,N_1939,N_1559);
nor U3039 (N_3039,N_342,N_571);
xor U3040 (N_3040,N_1704,N_885);
and U3041 (N_3041,N_97,N_453);
xor U3042 (N_3042,N_1035,N_1987);
nand U3043 (N_3043,N_293,N_882);
xor U3044 (N_3044,N_16,N_1533);
and U3045 (N_3045,N_450,N_1073);
nor U3046 (N_3046,N_1658,N_1332);
and U3047 (N_3047,N_1052,N_616);
xor U3048 (N_3048,N_1059,N_810);
nor U3049 (N_3049,N_1382,N_1255);
or U3050 (N_3050,N_1073,N_1731);
or U3051 (N_3051,N_1255,N_1416);
nand U3052 (N_3052,N_1050,N_568);
nor U3053 (N_3053,N_207,N_960);
nor U3054 (N_3054,N_1111,N_1237);
nand U3055 (N_3055,N_568,N_1512);
nand U3056 (N_3056,N_1732,N_492);
and U3057 (N_3057,N_1375,N_1908);
nand U3058 (N_3058,N_1860,N_144);
xnor U3059 (N_3059,N_1534,N_1737);
nand U3060 (N_3060,N_785,N_361);
or U3061 (N_3061,N_381,N_1626);
nand U3062 (N_3062,N_398,N_1270);
nor U3063 (N_3063,N_1277,N_1336);
nand U3064 (N_3064,N_33,N_1021);
xor U3065 (N_3065,N_707,N_1276);
or U3066 (N_3066,N_428,N_167);
and U3067 (N_3067,N_898,N_1854);
and U3068 (N_3068,N_1942,N_424);
and U3069 (N_3069,N_1415,N_1709);
and U3070 (N_3070,N_1994,N_1836);
nand U3071 (N_3071,N_571,N_351);
xnor U3072 (N_3072,N_1669,N_677);
and U3073 (N_3073,N_262,N_241);
or U3074 (N_3074,N_1948,N_870);
or U3075 (N_3075,N_155,N_659);
xnor U3076 (N_3076,N_1004,N_1893);
and U3077 (N_3077,N_1358,N_102);
nor U3078 (N_3078,N_37,N_1890);
and U3079 (N_3079,N_1199,N_1641);
or U3080 (N_3080,N_1312,N_1657);
or U3081 (N_3081,N_451,N_315);
nand U3082 (N_3082,N_391,N_481);
nor U3083 (N_3083,N_1545,N_1539);
or U3084 (N_3084,N_111,N_1370);
xnor U3085 (N_3085,N_645,N_1808);
nand U3086 (N_3086,N_960,N_1659);
and U3087 (N_3087,N_1867,N_1748);
and U3088 (N_3088,N_13,N_1700);
nor U3089 (N_3089,N_405,N_481);
nor U3090 (N_3090,N_990,N_1408);
nor U3091 (N_3091,N_466,N_1528);
or U3092 (N_3092,N_1072,N_816);
nand U3093 (N_3093,N_968,N_142);
and U3094 (N_3094,N_1081,N_953);
xor U3095 (N_3095,N_823,N_151);
nand U3096 (N_3096,N_1551,N_617);
or U3097 (N_3097,N_435,N_384);
nor U3098 (N_3098,N_1692,N_1778);
and U3099 (N_3099,N_1097,N_19);
and U3100 (N_3100,N_1519,N_303);
or U3101 (N_3101,N_400,N_1084);
or U3102 (N_3102,N_399,N_716);
or U3103 (N_3103,N_1784,N_523);
or U3104 (N_3104,N_718,N_1313);
or U3105 (N_3105,N_520,N_293);
or U3106 (N_3106,N_261,N_1961);
nand U3107 (N_3107,N_1812,N_974);
or U3108 (N_3108,N_1800,N_1568);
or U3109 (N_3109,N_377,N_586);
or U3110 (N_3110,N_1173,N_990);
nand U3111 (N_3111,N_1279,N_531);
and U3112 (N_3112,N_1261,N_818);
xnor U3113 (N_3113,N_1946,N_549);
and U3114 (N_3114,N_354,N_1336);
and U3115 (N_3115,N_786,N_1170);
xnor U3116 (N_3116,N_1501,N_564);
or U3117 (N_3117,N_463,N_758);
nor U3118 (N_3118,N_1872,N_29);
or U3119 (N_3119,N_1385,N_1005);
or U3120 (N_3120,N_534,N_524);
nor U3121 (N_3121,N_892,N_1701);
or U3122 (N_3122,N_862,N_826);
nor U3123 (N_3123,N_1858,N_1217);
xnor U3124 (N_3124,N_1808,N_521);
or U3125 (N_3125,N_40,N_362);
nand U3126 (N_3126,N_721,N_795);
nand U3127 (N_3127,N_1764,N_1314);
nor U3128 (N_3128,N_1911,N_666);
or U3129 (N_3129,N_159,N_811);
nor U3130 (N_3130,N_812,N_478);
nand U3131 (N_3131,N_194,N_1668);
and U3132 (N_3132,N_146,N_1885);
nand U3133 (N_3133,N_1384,N_1266);
and U3134 (N_3134,N_1609,N_84);
or U3135 (N_3135,N_890,N_486);
xor U3136 (N_3136,N_730,N_1295);
and U3137 (N_3137,N_357,N_847);
nor U3138 (N_3138,N_639,N_351);
or U3139 (N_3139,N_518,N_1251);
nand U3140 (N_3140,N_1009,N_1251);
nor U3141 (N_3141,N_67,N_351);
and U3142 (N_3142,N_876,N_908);
or U3143 (N_3143,N_1057,N_1525);
nand U3144 (N_3144,N_1440,N_1974);
or U3145 (N_3145,N_459,N_547);
or U3146 (N_3146,N_1495,N_709);
xnor U3147 (N_3147,N_1424,N_1427);
nand U3148 (N_3148,N_1571,N_1807);
nor U3149 (N_3149,N_1864,N_434);
nor U3150 (N_3150,N_894,N_781);
or U3151 (N_3151,N_671,N_796);
nor U3152 (N_3152,N_976,N_1971);
or U3153 (N_3153,N_58,N_1847);
or U3154 (N_3154,N_631,N_1342);
and U3155 (N_3155,N_1773,N_1334);
nand U3156 (N_3156,N_1930,N_1619);
and U3157 (N_3157,N_1328,N_1729);
xnor U3158 (N_3158,N_379,N_1566);
nor U3159 (N_3159,N_1565,N_1257);
nor U3160 (N_3160,N_1890,N_856);
or U3161 (N_3161,N_622,N_709);
or U3162 (N_3162,N_1123,N_691);
and U3163 (N_3163,N_1777,N_1206);
nand U3164 (N_3164,N_1667,N_122);
or U3165 (N_3165,N_954,N_1046);
nor U3166 (N_3166,N_1898,N_1273);
nor U3167 (N_3167,N_145,N_1777);
nor U3168 (N_3168,N_756,N_1612);
nand U3169 (N_3169,N_1307,N_946);
and U3170 (N_3170,N_601,N_1977);
xor U3171 (N_3171,N_1655,N_1422);
and U3172 (N_3172,N_1467,N_305);
nand U3173 (N_3173,N_960,N_351);
nand U3174 (N_3174,N_434,N_414);
nand U3175 (N_3175,N_903,N_92);
or U3176 (N_3176,N_164,N_227);
xor U3177 (N_3177,N_1699,N_1718);
nor U3178 (N_3178,N_1512,N_1115);
nand U3179 (N_3179,N_684,N_40);
nor U3180 (N_3180,N_533,N_276);
nor U3181 (N_3181,N_1102,N_707);
nand U3182 (N_3182,N_595,N_1324);
or U3183 (N_3183,N_400,N_574);
xnor U3184 (N_3184,N_1434,N_1649);
nor U3185 (N_3185,N_806,N_786);
xor U3186 (N_3186,N_119,N_1426);
nor U3187 (N_3187,N_408,N_187);
nor U3188 (N_3188,N_406,N_160);
and U3189 (N_3189,N_566,N_75);
nand U3190 (N_3190,N_636,N_1005);
nor U3191 (N_3191,N_1749,N_294);
and U3192 (N_3192,N_91,N_473);
or U3193 (N_3193,N_1639,N_371);
nand U3194 (N_3194,N_1725,N_1359);
nor U3195 (N_3195,N_57,N_675);
xnor U3196 (N_3196,N_1637,N_1044);
nand U3197 (N_3197,N_961,N_611);
or U3198 (N_3198,N_1976,N_1317);
and U3199 (N_3199,N_884,N_1055);
nand U3200 (N_3200,N_306,N_1223);
nor U3201 (N_3201,N_1010,N_656);
nor U3202 (N_3202,N_1626,N_1866);
or U3203 (N_3203,N_1959,N_1268);
or U3204 (N_3204,N_1307,N_1684);
or U3205 (N_3205,N_1312,N_1160);
nor U3206 (N_3206,N_323,N_1571);
nand U3207 (N_3207,N_1236,N_1453);
nand U3208 (N_3208,N_462,N_787);
or U3209 (N_3209,N_128,N_1157);
xnor U3210 (N_3210,N_1728,N_692);
nand U3211 (N_3211,N_639,N_1099);
or U3212 (N_3212,N_694,N_1681);
nand U3213 (N_3213,N_1242,N_1100);
or U3214 (N_3214,N_118,N_1552);
nor U3215 (N_3215,N_311,N_983);
and U3216 (N_3216,N_1790,N_464);
xnor U3217 (N_3217,N_975,N_1289);
or U3218 (N_3218,N_878,N_1001);
xnor U3219 (N_3219,N_343,N_623);
nand U3220 (N_3220,N_142,N_978);
nor U3221 (N_3221,N_1436,N_1859);
and U3222 (N_3222,N_1862,N_263);
and U3223 (N_3223,N_322,N_686);
or U3224 (N_3224,N_1370,N_39);
nand U3225 (N_3225,N_1347,N_1705);
nor U3226 (N_3226,N_1369,N_1517);
and U3227 (N_3227,N_1842,N_1706);
and U3228 (N_3228,N_1599,N_1208);
and U3229 (N_3229,N_1222,N_1895);
or U3230 (N_3230,N_1619,N_592);
nand U3231 (N_3231,N_622,N_1837);
and U3232 (N_3232,N_682,N_645);
and U3233 (N_3233,N_893,N_1764);
or U3234 (N_3234,N_1217,N_132);
or U3235 (N_3235,N_927,N_1070);
and U3236 (N_3236,N_1848,N_841);
and U3237 (N_3237,N_1786,N_1411);
nor U3238 (N_3238,N_791,N_544);
or U3239 (N_3239,N_1309,N_901);
nand U3240 (N_3240,N_1507,N_1653);
and U3241 (N_3241,N_1881,N_1823);
nor U3242 (N_3242,N_1105,N_637);
xor U3243 (N_3243,N_620,N_1265);
xnor U3244 (N_3244,N_1781,N_1182);
nor U3245 (N_3245,N_204,N_678);
and U3246 (N_3246,N_105,N_1246);
or U3247 (N_3247,N_1195,N_712);
and U3248 (N_3248,N_119,N_836);
and U3249 (N_3249,N_873,N_192);
or U3250 (N_3250,N_1757,N_229);
nor U3251 (N_3251,N_557,N_1525);
nor U3252 (N_3252,N_1890,N_75);
or U3253 (N_3253,N_326,N_839);
xor U3254 (N_3254,N_1881,N_682);
nand U3255 (N_3255,N_640,N_1838);
or U3256 (N_3256,N_191,N_889);
and U3257 (N_3257,N_889,N_1481);
and U3258 (N_3258,N_886,N_1949);
or U3259 (N_3259,N_431,N_825);
and U3260 (N_3260,N_590,N_441);
xnor U3261 (N_3261,N_1985,N_1662);
and U3262 (N_3262,N_1539,N_69);
nor U3263 (N_3263,N_601,N_1912);
nand U3264 (N_3264,N_1574,N_1747);
or U3265 (N_3265,N_561,N_1504);
and U3266 (N_3266,N_1563,N_12);
and U3267 (N_3267,N_240,N_1668);
or U3268 (N_3268,N_1634,N_101);
nand U3269 (N_3269,N_1589,N_749);
or U3270 (N_3270,N_660,N_1757);
nand U3271 (N_3271,N_774,N_1490);
and U3272 (N_3272,N_1453,N_1982);
nor U3273 (N_3273,N_1987,N_181);
nor U3274 (N_3274,N_434,N_1326);
nand U3275 (N_3275,N_1509,N_633);
nor U3276 (N_3276,N_89,N_1132);
and U3277 (N_3277,N_1694,N_166);
and U3278 (N_3278,N_35,N_112);
nand U3279 (N_3279,N_1238,N_692);
and U3280 (N_3280,N_1942,N_200);
nand U3281 (N_3281,N_1422,N_1356);
nand U3282 (N_3282,N_94,N_1931);
or U3283 (N_3283,N_1536,N_503);
or U3284 (N_3284,N_842,N_1514);
and U3285 (N_3285,N_129,N_450);
and U3286 (N_3286,N_1167,N_460);
or U3287 (N_3287,N_339,N_1602);
or U3288 (N_3288,N_1393,N_1638);
and U3289 (N_3289,N_806,N_1362);
or U3290 (N_3290,N_694,N_613);
and U3291 (N_3291,N_1055,N_925);
nand U3292 (N_3292,N_258,N_69);
nor U3293 (N_3293,N_505,N_45);
nor U3294 (N_3294,N_1556,N_372);
or U3295 (N_3295,N_1931,N_199);
nor U3296 (N_3296,N_1707,N_1752);
and U3297 (N_3297,N_1,N_1634);
and U3298 (N_3298,N_344,N_959);
xnor U3299 (N_3299,N_1404,N_903);
nor U3300 (N_3300,N_1103,N_755);
or U3301 (N_3301,N_1761,N_420);
and U3302 (N_3302,N_648,N_1524);
and U3303 (N_3303,N_714,N_940);
nand U3304 (N_3304,N_1998,N_590);
xor U3305 (N_3305,N_1698,N_449);
and U3306 (N_3306,N_1348,N_1136);
nand U3307 (N_3307,N_110,N_669);
nor U3308 (N_3308,N_1518,N_1600);
nand U3309 (N_3309,N_1149,N_1070);
xnor U3310 (N_3310,N_66,N_1002);
and U3311 (N_3311,N_387,N_1941);
or U3312 (N_3312,N_566,N_1570);
nand U3313 (N_3313,N_1105,N_232);
nand U3314 (N_3314,N_301,N_328);
and U3315 (N_3315,N_1675,N_34);
or U3316 (N_3316,N_1261,N_472);
xnor U3317 (N_3317,N_57,N_1749);
nand U3318 (N_3318,N_611,N_1135);
nor U3319 (N_3319,N_813,N_1844);
nand U3320 (N_3320,N_221,N_1659);
nand U3321 (N_3321,N_870,N_672);
and U3322 (N_3322,N_289,N_1412);
and U3323 (N_3323,N_1976,N_1922);
nor U3324 (N_3324,N_832,N_773);
nand U3325 (N_3325,N_75,N_54);
or U3326 (N_3326,N_945,N_367);
and U3327 (N_3327,N_278,N_1900);
nand U3328 (N_3328,N_1748,N_920);
nor U3329 (N_3329,N_1658,N_1770);
xnor U3330 (N_3330,N_751,N_732);
nor U3331 (N_3331,N_756,N_1180);
or U3332 (N_3332,N_1171,N_464);
nand U3333 (N_3333,N_1215,N_1989);
nand U3334 (N_3334,N_1393,N_1588);
nor U3335 (N_3335,N_503,N_1213);
nor U3336 (N_3336,N_362,N_1759);
nand U3337 (N_3337,N_727,N_1522);
nand U3338 (N_3338,N_524,N_894);
nor U3339 (N_3339,N_194,N_1644);
xnor U3340 (N_3340,N_335,N_1231);
nand U3341 (N_3341,N_185,N_812);
nor U3342 (N_3342,N_1281,N_1976);
nor U3343 (N_3343,N_140,N_910);
or U3344 (N_3344,N_1338,N_1328);
and U3345 (N_3345,N_1084,N_1429);
nor U3346 (N_3346,N_1451,N_1690);
xor U3347 (N_3347,N_164,N_126);
and U3348 (N_3348,N_1474,N_1353);
xor U3349 (N_3349,N_1522,N_378);
nor U3350 (N_3350,N_1517,N_1513);
nor U3351 (N_3351,N_1974,N_1585);
and U3352 (N_3352,N_1300,N_1790);
or U3353 (N_3353,N_202,N_1897);
and U3354 (N_3354,N_1947,N_1727);
xor U3355 (N_3355,N_1551,N_860);
or U3356 (N_3356,N_139,N_1633);
or U3357 (N_3357,N_1589,N_760);
or U3358 (N_3358,N_1544,N_1683);
or U3359 (N_3359,N_533,N_682);
and U3360 (N_3360,N_664,N_505);
and U3361 (N_3361,N_970,N_1158);
nor U3362 (N_3362,N_1311,N_1407);
xor U3363 (N_3363,N_1250,N_397);
or U3364 (N_3364,N_1569,N_1186);
or U3365 (N_3365,N_38,N_783);
nand U3366 (N_3366,N_958,N_89);
nor U3367 (N_3367,N_691,N_327);
xnor U3368 (N_3368,N_123,N_1277);
nor U3369 (N_3369,N_1420,N_1909);
or U3370 (N_3370,N_481,N_1468);
nand U3371 (N_3371,N_1797,N_1830);
nor U3372 (N_3372,N_154,N_686);
nor U3373 (N_3373,N_58,N_1151);
nor U3374 (N_3374,N_743,N_1816);
nand U3375 (N_3375,N_1838,N_1543);
or U3376 (N_3376,N_293,N_1933);
nand U3377 (N_3377,N_1445,N_201);
nor U3378 (N_3378,N_1826,N_873);
nor U3379 (N_3379,N_1109,N_84);
or U3380 (N_3380,N_279,N_511);
or U3381 (N_3381,N_1780,N_397);
and U3382 (N_3382,N_1941,N_1134);
xor U3383 (N_3383,N_1536,N_211);
or U3384 (N_3384,N_443,N_1360);
or U3385 (N_3385,N_767,N_1862);
nand U3386 (N_3386,N_153,N_708);
and U3387 (N_3387,N_1769,N_430);
nor U3388 (N_3388,N_1228,N_1829);
nand U3389 (N_3389,N_285,N_1970);
nand U3390 (N_3390,N_578,N_1771);
and U3391 (N_3391,N_244,N_1429);
nor U3392 (N_3392,N_536,N_1525);
or U3393 (N_3393,N_1186,N_846);
or U3394 (N_3394,N_476,N_186);
nand U3395 (N_3395,N_501,N_1266);
or U3396 (N_3396,N_1665,N_677);
or U3397 (N_3397,N_1456,N_1670);
or U3398 (N_3398,N_1853,N_935);
nor U3399 (N_3399,N_901,N_154);
nand U3400 (N_3400,N_317,N_878);
and U3401 (N_3401,N_1819,N_422);
or U3402 (N_3402,N_1131,N_1260);
or U3403 (N_3403,N_1547,N_1918);
xnor U3404 (N_3404,N_561,N_677);
nor U3405 (N_3405,N_1587,N_1470);
nand U3406 (N_3406,N_1733,N_445);
nor U3407 (N_3407,N_505,N_12);
and U3408 (N_3408,N_387,N_476);
and U3409 (N_3409,N_1785,N_15);
or U3410 (N_3410,N_1917,N_1461);
nand U3411 (N_3411,N_1541,N_68);
and U3412 (N_3412,N_199,N_126);
or U3413 (N_3413,N_1228,N_1288);
and U3414 (N_3414,N_1524,N_1700);
or U3415 (N_3415,N_1533,N_216);
or U3416 (N_3416,N_86,N_525);
nor U3417 (N_3417,N_446,N_126);
and U3418 (N_3418,N_1385,N_455);
nand U3419 (N_3419,N_332,N_1347);
nand U3420 (N_3420,N_74,N_1432);
and U3421 (N_3421,N_967,N_1387);
nand U3422 (N_3422,N_1208,N_269);
or U3423 (N_3423,N_1287,N_356);
and U3424 (N_3424,N_1785,N_1382);
nor U3425 (N_3425,N_475,N_903);
or U3426 (N_3426,N_292,N_1286);
and U3427 (N_3427,N_1666,N_1642);
and U3428 (N_3428,N_126,N_1574);
or U3429 (N_3429,N_1090,N_402);
nor U3430 (N_3430,N_434,N_604);
and U3431 (N_3431,N_1731,N_736);
and U3432 (N_3432,N_1308,N_528);
xnor U3433 (N_3433,N_1803,N_0);
and U3434 (N_3434,N_97,N_103);
xnor U3435 (N_3435,N_1011,N_110);
xnor U3436 (N_3436,N_684,N_79);
and U3437 (N_3437,N_1327,N_1507);
or U3438 (N_3438,N_955,N_1167);
nand U3439 (N_3439,N_335,N_439);
nor U3440 (N_3440,N_1552,N_301);
nor U3441 (N_3441,N_1631,N_905);
and U3442 (N_3442,N_1797,N_1448);
nand U3443 (N_3443,N_1381,N_679);
and U3444 (N_3444,N_1009,N_438);
nor U3445 (N_3445,N_457,N_1107);
nand U3446 (N_3446,N_1794,N_1932);
nand U3447 (N_3447,N_922,N_1320);
nor U3448 (N_3448,N_804,N_1743);
nand U3449 (N_3449,N_1740,N_1014);
xor U3450 (N_3450,N_1008,N_349);
and U3451 (N_3451,N_119,N_754);
xor U3452 (N_3452,N_1201,N_1747);
nor U3453 (N_3453,N_1912,N_760);
or U3454 (N_3454,N_674,N_1904);
xnor U3455 (N_3455,N_68,N_526);
or U3456 (N_3456,N_1091,N_1475);
xnor U3457 (N_3457,N_1631,N_1801);
xor U3458 (N_3458,N_650,N_1354);
xnor U3459 (N_3459,N_791,N_1927);
nor U3460 (N_3460,N_1569,N_561);
or U3461 (N_3461,N_179,N_1904);
nand U3462 (N_3462,N_1168,N_150);
xnor U3463 (N_3463,N_1674,N_915);
nor U3464 (N_3464,N_1828,N_1536);
and U3465 (N_3465,N_1760,N_624);
nor U3466 (N_3466,N_857,N_762);
nor U3467 (N_3467,N_446,N_1462);
and U3468 (N_3468,N_202,N_736);
nor U3469 (N_3469,N_352,N_643);
or U3470 (N_3470,N_1989,N_1272);
and U3471 (N_3471,N_891,N_920);
or U3472 (N_3472,N_459,N_1447);
nand U3473 (N_3473,N_393,N_846);
and U3474 (N_3474,N_1327,N_1013);
nand U3475 (N_3475,N_1716,N_691);
or U3476 (N_3476,N_1183,N_241);
or U3477 (N_3477,N_269,N_80);
and U3478 (N_3478,N_1750,N_114);
nor U3479 (N_3479,N_480,N_70);
nand U3480 (N_3480,N_1826,N_265);
nor U3481 (N_3481,N_1733,N_373);
xnor U3482 (N_3482,N_532,N_386);
nand U3483 (N_3483,N_1167,N_122);
nor U3484 (N_3484,N_1295,N_1183);
xnor U3485 (N_3485,N_1760,N_318);
nor U3486 (N_3486,N_323,N_1639);
nand U3487 (N_3487,N_60,N_1828);
nor U3488 (N_3488,N_598,N_458);
nor U3489 (N_3489,N_686,N_1170);
and U3490 (N_3490,N_1912,N_766);
or U3491 (N_3491,N_157,N_1276);
or U3492 (N_3492,N_772,N_752);
or U3493 (N_3493,N_1815,N_1527);
nand U3494 (N_3494,N_1973,N_1187);
or U3495 (N_3495,N_1484,N_78);
and U3496 (N_3496,N_1811,N_801);
nor U3497 (N_3497,N_1138,N_1693);
nand U3498 (N_3498,N_1539,N_1645);
and U3499 (N_3499,N_430,N_434);
and U3500 (N_3500,N_1124,N_1749);
nor U3501 (N_3501,N_49,N_1369);
xnor U3502 (N_3502,N_1686,N_1188);
or U3503 (N_3503,N_864,N_236);
nor U3504 (N_3504,N_430,N_1114);
or U3505 (N_3505,N_1145,N_1885);
nor U3506 (N_3506,N_520,N_310);
and U3507 (N_3507,N_1783,N_186);
and U3508 (N_3508,N_1985,N_1791);
nor U3509 (N_3509,N_817,N_227);
xor U3510 (N_3510,N_374,N_1077);
and U3511 (N_3511,N_1060,N_363);
or U3512 (N_3512,N_1593,N_1404);
or U3513 (N_3513,N_196,N_382);
or U3514 (N_3514,N_996,N_1085);
nand U3515 (N_3515,N_145,N_85);
nor U3516 (N_3516,N_1075,N_556);
and U3517 (N_3517,N_744,N_964);
nor U3518 (N_3518,N_1482,N_1839);
nor U3519 (N_3519,N_1811,N_1359);
nor U3520 (N_3520,N_921,N_1387);
and U3521 (N_3521,N_1202,N_1100);
nand U3522 (N_3522,N_1098,N_492);
nor U3523 (N_3523,N_1360,N_1258);
nand U3524 (N_3524,N_193,N_1226);
and U3525 (N_3525,N_1294,N_228);
nand U3526 (N_3526,N_1723,N_717);
and U3527 (N_3527,N_249,N_1786);
nor U3528 (N_3528,N_1413,N_599);
nand U3529 (N_3529,N_1427,N_1246);
nor U3530 (N_3530,N_180,N_1095);
and U3531 (N_3531,N_1558,N_802);
xnor U3532 (N_3532,N_588,N_1720);
nand U3533 (N_3533,N_1963,N_1259);
nor U3534 (N_3534,N_335,N_499);
or U3535 (N_3535,N_1781,N_1121);
or U3536 (N_3536,N_1808,N_167);
or U3537 (N_3537,N_1247,N_475);
nand U3538 (N_3538,N_1934,N_526);
nand U3539 (N_3539,N_1120,N_475);
nor U3540 (N_3540,N_277,N_406);
or U3541 (N_3541,N_1107,N_1365);
or U3542 (N_3542,N_1830,N_1058);
nor U3543 (N_3543,N_291,N_1663);
nand U3544 (N_3544,N_1673,N_1334);
and U3545 (N_3545,N_565,N_1392);
and U3546 (N_3546,N_1541,N_943);
nand U3547 (N_3547,N_672,N_1482);
nand U3548 (N_3548,N_646,N_1259);
or U3549 (N_3549,N_1876,N_491);
or U3550 (N_3550,N_1587,N_1613);
nor U3551 (N_3551,N_1331,N_1055);
and U3552 (N_3552,N_506,N_240);
and U3553 (N_3553,N_567,N_352);
and U3554 (N_3554,N_471,N_1835);
nor U3555 (N_3555,N_1791,N_1617);
xnor U3556 (N_3556,N_1842,N_1562);
or U3557 (N_3557,N_221,N_1921);
nor U3558 (N_3558,N_1702,N_1055);
nor U3559 (N_3559,N_1204,N_1732);
nor U3560 (N_3560,N_1202,N_594);
or U3561 (N_3561,N_704,N_1737);
and U3562 (N_3562,N_1987,N_1484);
nand U3563 (N_3563,N_1537,N_232);
and U3564 (N_3564,N_967,N_725);
nor U3565 (N_3565,N_1806,N_1059);
or U3566 (N_3566,N_469,N_1717);
or U3567 (N_3567,N_1790,N_1204);
nor U3568 (N_3568,N_1480,N_558);
or U3569 (N_3569,N_765,N_725);
nor U3570 (N_3570,N_1218,N_80);
nand U3571 (N_3571,N_327,N_1387);
nor U3572 (N_3572,N_1360,N_1959);
or U3573 (N_3573,N_636,N_1135);
nand U3574 (N_3574,N_1482,N_1551);
nand U3575 (N_3575,N_524,N_1536);
or U3576 (N_3576,N_42,N_1173);
and U3577 (N_3577,N_548,N_118);
xnor U3578 (N_3578,N_688,N_317);
and U3579 (N_3579,N_1915,N_1836);
nand U3580 (N_3580,N_61,N_521);
nor U3581 (N_3581,N_668,N_1517);
and U3582 (N_3582,N_123,N_1365);
or U3583 (N_3583,N_1898,N_791);
nor U3584 (N_3584,N_1392,N_827);
and U3585 (N_3585,N_1124,N_1242);
and U3586 (N_3586,N_1324,N_542);
nor U3587 (N_3587,N_1415,N_1581);
nand U3588 (N_3588,N_1110,N_1001);
and U3589 (N_3589,N_1092,N_1835);
nor U3590 (N_3590,N_461,N_977);
and U3591 (N_3591,N_1413,N_1599);
nor U3592 (N_3592,N_1825,N_936);
and U3593 (N_3593,N_177,N_1065);
xnor U3594 (N_3594,N_77,N_1302);
or U3595 (N_3595,N_1093,N_793);
nand U3596 (N_3596,N_1077,N_551);
and U3597 (N_3597,N_1207,N_666);
and U3598 (N_3598,N_348,N_909);
nand U3599 (N_3599,N_1895,N_1091);
or U3600 (N_3600,N_553,N_571);
nand U3601 (N_3601,N_977,N_1494);
nand U3602 (N_3602,N_1813,N_1570);
nor U3603 (N_3603,N_1949,N_454);
nor U3604 (N_3604,N_1657,N_919);
nor U3605 (N_3605,N_1755,N_1997);
xnor U3606 (N_3606,N_1162,N_222);
or U3607 (N_3607,N_873,N_94);
and U3608 (N_3608,N_102,N_1357);
or U3609 (N_3609,N_1843,N_989);
nor U3610 (N_3610,N_283,N_619);
nor U3611 (N_3611,N_394,N_450);
and U3612 (N_3612,N_1393,N_1274);
nand U3613 (N_3613,N_1019,N_1858);
nor U3614 (N_3614,N_1114,N_988);
and U3615 (N_3615,N_1893,N_803);
nor U3616 (N_3616,N_965,N_622);
and U3617 (N_3617,N_1028,N_594);
and U3618 (N_3618,N_1417,N_1301);
and U3619 (N_3619,N_1863,N_168);
and U3620 (N_3620,N_1512,N_1066);
nand U3621 (N_3621,N_1567,N_551);
nor U3622 (N_3622,N_1872,N_1529);
nand U3623 (N_3623,N_1991,N_133);
nor U3624 (N_3624,N_523,N_1320);
nor U3625 (N_3625,N_693,N_107);
nor U3626 (N_3626,N_1645,N_310);
nor U3627 (N_3627,N_1042,N_1029);
and U3628 (N_3628,N_1324,N_782);
and U3629 (N_3629,N_1793,N_354);
nand U3630 (N_3630,N_310,N_953);
nand U3631 (N_3631,N_1981,N_201);
xor U3632 (N_3632,N_1640,N_503);
nor U3633 (N_3633,N_1425,N_767);
and U3634 (N_3634,N_343,N_59);
nor U3635 (N_3635,N_305,N_1173);
nor U3636 (N_3636,N_1590,N_1690);
nand U3637 (N_3637,N_5,N_472);
nor U3638 (N_3638,N_1766,N_591);
nand U3639 (N_3639,N_1495,N_756);
xnor U3640 (N_3640,N_762,N_1595);
and U3641 (N_3641,N_942,N_1519);
nand U3642 (N_3642,N_1380,N_1213);
nor U3643 (N_3643,N_1451,N_1816);
xor U3644 (N_3644,N_25,N_1932);
nand U3645 (N_3645,N_1141,N_1114);
and U3646 (N_3646,N_422,N_861);
and U3647 (N_3647,N_628,N_650);
xnor U3648 (N_3648,N_177,N_281);
nor U3649 (N_3649,N_1154,N_1987);
or U3650 (N_3650,N_1290,N_1170);
and U3651 (N_3651,N_1400,N_1779);
nand U3652 (N_3652,N_1946,N_896);
nand U3653 (N_3653,N_713,N_1309);
and U3654 (N_3654,N_1471,N_1699);
nand U3655 (N_3655,N_1212,N_889);
and U3656 (N_3656,N_1928,N_466);
and U3657 (N_3657,N_1019,N_1374);
and U3658 (N_3658,N_1438,N_814);
and U3659 (N_3659,N_479,N_466);
and U3660 (N_3660,N_700,N_678);
or U3661 (N_3661,N_971,N_582);
and U3662 (N_3662,N_1995,N_574);
and U3663 (N_3663,N_1121,N_1549);
and U3664 (N_3664,N_874,N_1309);
and U3665 (N_3665,N_1970,N_1983);
or U3666 (N_3666,N_1886,N_1209);
or U3667 (N_3667,N_1236,N_1217);
nor U3668 (N_3668,N_1977,N_1154);
nor U3669 (N_3669,N_517,N_1581);
nor U3670 (N_3670,N_334,N_1792);
nand U3671 (N_3671,N_1927,N_1760);
nor U3672 (N_3672,N_313,N_1498);
or U3673 (N_3673,N_1607,N_1938);
nor U3674 (N_3674,N_9,N_1350);
or U3675 (N_3675,N_222,N_1316);
nand U3676 (N_3676,N_1696,N_765);
or U3677 (N_3677,N_1367,N_1436);
and U3678 (N_3678,N_1677,N_91);
xor U3679 (N_3679,N_936,N_1300);
nor U3680 (N_3680,N_1859,N_1264);
or U3681 (N_3681,N_802,N_1006);
nor U3682 (N_3682,N_96,N_1806);
or U3683 (N_3683,N_765,N_1127);
and U3684 (N_3684,N_1298,N_712);
nand U3685 (N_3685,N_549,N_344);
or U3686 (N_3686,N_1015,N_974);
xnor U3687 (N_3687,N_976,N_663);
nor U3688 (N_3688,N_1638,N_1467);
or U3689 (N_3689,N_550,N_460);
and U3690 (N_3690,N_416,N_1661);
xnor U3691 (N_3691,N_695,N_1042);
and U3692 (N_3692,N_1411,N_987);
or U3693 (N_3693,N_398,N_1670);
or U3694 (N_3694,N_805,N_413);
nor U3695 (N_3695,N_1416,N_1328);
xor U3696 (N_3696,N_1017,N_1776);
xor U3697 (N_3697,N_1362,N_900);
or U3698 (N_3698,N_1155,N_1276);
and U3699 (N_3699,N_1419,N_1112);
and U3700 (N_3700,N_1972,N_1053);
xor U3701 (N_3701,N_1442,N_1318);
xor U3702 (N_3702,N_954,N_829);
nand U3703 (N_3703,N_963,N_403);
and U3704 (N_3704,N_1778,N_855);
and U3705 (N_3705,N_438,N_769);
or U3706 (N_3706,N_104,N_1580);
or U3707 (N_3707,N_354,N_1493);
nand U3708 (N_3708,N_1364,N_1721);
nand U3709 (N_3709,N_744,N_175);
and U3710 (N_3710,N_984,N_1076);
or U3711 (N_3711,N_1642,N_1778);
and U3712 (N_3712,N_198,N_1297);
xnor U3713 (N_3713,N_1924,N_1338);
or U3714 (N_3714,N_117,N_303);
and U3715 (N_3715,N_413,N_1697);
and U3716 (N_3716,N_1502,N_380);
or U3717 (N_3717,N_48,N_1269);
nor U3718 (N_3718,N_1722,N_33);
nand U3719 (N_3719,N_458,N_150);
xnor U3720 (N_3720,N_593,N_666);
nor U3721 (N_3721,N_1997,N_242);
xnor U3722 (N_3722,N_333,N_1016);
and U3723 (N_3723,N_1249,N_979);
xnor U3724 (N_3724,N_700,N_580);
or U3725 (N_3725,N_273,N_1680);
and U3726 (N_3726,N_1137,N_361);
and U3727 (N_3727,N_1490,N_178);
or U3728 (N_3728,N_1781,N_529);
nor U3729 (N_3729,N_159,N_919);
nand U3730 (N_3730,N_680,N_76);
nand U3731 (N_3731,N_10,N_735);
nand U3732 (N_3732,N_1086,N_964);
xnor U3733 (N_3733,N_1333,N_901);
nand U3734 (N_3734,N_1791,N_1023);
and U3735 (N_3735,N_593,N_910);
nor U3736 (N_3736,N_1289,N_1420);
or U3737 (N_3737,N_1167,N_1044);
or U3738 (N_3738,N_1325,N_1789);
nor U3739 (N_3739,N_627,N_389);
and U3740 (N_3740,N_1117,N_1977);
or U3741 (N_3741,N_871,N_424);
and U3742 (N_3742,N_1656,N_698);
nand U3743 (N_3743,N_1124,N_211);
or U3744 (N_3744,N_331,N_1527);
or U3745 (N_3745,N_1845,N_1306);
nor U3746 (N_3746,N_47,N_791);
or U3747 (N_3747,N_718,N_592);
nor U3748 (N_3748,N_1219,N_329);
nand U3749 (N_3749,N_1661,N_962);
xor U3750 (N_3750,N_70,N_1535);
nor U3751 (N_3751,N_341,N_4);
and U3752 (N_3752,N_1449,N_1329);
and U3753 (N_3753,N_1904,N_28);
xor U3754 (N_3754,N_1022,N_300);
nor U3755 (N_3755,N_297,N_193);
or U3756 (N_3756,N_376,N_1466);
or U3757 (N_3757,N_63,N_449);
or U3758 (N_3758,N_572,N_1524);
nand U3759 (N_3759,N_1042,N_305);
nor U3760 (N_3760,N_564,N_1351);
or U3761 (N_3761,N_1100,N_1796);
xor U3762 (N_3762,N_396,N_839);
nor U3763 (N_3763,N_1266,N_27);
nor U3764 (N_3764,N_1798,N_1450);
or U3765 (N_3765,N_1827,N_234);
and U3766 (N_3766,N_461,N_1297);
and U3767 (N_3767,N_1752,N_1275);
nor U3768 (N_3768,N_107,N_1745);
or U3769 (N_3769,N_506,N_1179);
nand U3770 (N_3770,N_1930,N_759);
nor U3771 (N_3771,N_1724,N_1159);
or U3772 (N_3772,N_1100,N_300);
and U3773 (N_3773,N_639,N_1059);
nand U3774 (N_3774,N_1836,N_1581);
and U3775 (N_3775,N_893,N_1546);
and U3776 (N_3776,N_1954,N_1998);
nor U3777 (N_3777,N_1655,N_1385);
and U3778 (N_3778,N_1361,N_102);
nand U3779 (N_3779,N_1458,N_920);
and U3780 (N_3780,N_844,N_1863);
and U3781 (N_3781,N_225,N_876);
nor U3782 (N_3782,N_719,N_1705);
or U3783 (N_3783,N_512,N_247);
nand U3784 (N_3784,N_1347,N_1890);
nand U3785 (N_3785,N_1293,N_1818);
nor U3786 (N_3786,N_1644,N_1400);
and U3787 (N_3787,N_1018,N_1789);
nor U3788 (N_3788,N_225,N_406);
xnor U3789 (N_3789,N_829,N_1905);
or U3790 (N_3790,N_732,N_320);
nand U3791 (N_3791,N_1107,N_70);
and U3792 (N_3792,N_99,N_1977);
nand U3793 (N_3793,N_1382,N_1771);
xnor U3794 (N_3794,N_1472,N_1253);
or U3795 (N_3795,N_1987,N_666);
or U3796 (N_3796,N_1473,N_1052);
and U3797 (N_3797,N_1202,N_1709);
xnor U3798 (N_3798,N_1247,N_1764);
and U3799 (N_3799,N_1043,N_1962);
and U3800 (N_3800,N_1074,N_503);
nand U3801 (N_3801,N_1965,N_1985);
nand U3802 (N_3802,N_1457,N_33);
and U3803 (N_3803,N_247,N_1082);
and U3804 (N_3804,N_895,N_945);
and U3805 (N_3805,N_490,N_1678);
and U3806 (N_3806,N_1765,N_1608);
and U3807 (N_3807,N_889,N_710);
xnor U3808 (N_3808,N_793,N_815);
or U3809 (N_3809,N_1120,N_651);
and U3810 (N_3810,N_1275,N_875);
nand U3811 (N_3811,N_322,N_1708);
nor U3812 (N_3812,N_837,N_1599);
xor U3813 (N_3813,N_1641,N_605);
nor U3814 (N_3814,N_1882,N_755);
or U3815 (N_3815,N_1273,N_720);
and U3816 (N_3816,N_388,N_997);
nor U3817 (N_3817,N_1601,N_1046);
nor U3818 (N_3818,N_1213,N_1822);
nor U3819 (N_3819,N_1241,N_210);
or U3820 (N_3820,N_622,N_100);
or U3821 (N_3821,N_377,N_693);
xor U3822 (N_3822,N_1840,N_115);
and U3823 (N_3823,N_856,N_401);
or U3824 (N_3824,N_311,N_1868);
nand U3825 (N_3825,N_1841,N_1737);
or U3826 (N_3826,N_260,N_1704);
nand U3827 (N_3827,N_1504,N_1407);
and U3828 (N_3828,N_1728,N_1312);
nand U3829 (N_3829,N_1000,N_289);
nor U3830 (N_3830,N_1238,N_1292);
and U3831 (N_3831,N_503,N_1436);
nor U3832 (N_3832,N_768,N_593);
or U3833 (N_3833,N_400,N_362);
nor U3834 (N_3834,N_1909,N_1407);
or U3835 (N_3835,N_1357,N_1954);
and U3836 (N_3836,N_1483,N_137);
xor U3837 (N_3837,N_1522,N_1061);
nor U3838 (N_3838,N_1392,N_138);
and U3839 (N_3839,N_1231,N_1239);
or U3840 (N_3840,N_1612,N_1102);
nor U3841 (N_3841,N_1876,N_50);
or U3842 (N_3842,N_515,N_1697);
nor U3843 (N_3843,N_637,N_302);
or U3844 (N_3844,N_815,N_1476);
and U3845 (N_3845,N_1493,N_70);
nand U3846 (N_3846,N_1884,N_733);
nor U3847 (N_3847,N_1766,N_893);
and U3848 (N_3848,N_1951,N_113);
nand U3849 (N_3849,N_1890,N_396);
or U3850 (N_3850,N_335,N_639);
or U3851 (N_3851,N_1827,N_1667);
or U3852 (N_3852,N_1198,N_1970);
nand U3853 (N_3853,N_1000,N_897);
and U3854 (N_3854,N_1954,N_1020);
and U3855 (N_3855,N_747,N_331);
or U3856 (N_3856,N_870,N_447);
nor U3857 (N_3857,N_105,N_563);
nor U3858 (N_3858,N_1453,N_1828);
nor U3859 (N_3859,N_1112,N_966);
or U3860 (N_3860,N_96,N_264);
or U3861 (N_3861,N_636,N_1580);
xnor U3862 (N_3862,N_1908,N_327);
nand U3863 (N_3863,N_1459,N_1902);
or U3864 (N_3864,N_576,N_720);
or U3865 (N_3865,N_1309,N_520);
nor U3866 (N_3866,N_1554,N_28);
or U3867 (N_3867,N_1231,N_644);
xor U3868 (N_3868,N_1727,N_1313);
xor U3869 (N_3869,N_638,N_1318);
nand U3870 (N_3870,N_1084,N_1921);
and U3871 (N_3871,N_1063,N_694);
nand U3872 (N_3872,N_335,N_1794);
nor U3873 (N_3873,N_873,N_1624);
nand U3874 (N_3874,N_689,N_240);
xnor U3875 (N_3875,N_53,N_1642);
nand U3876 (N_3876,N_1895,N_1326);
and U3877 (N_3877,N_1655,N_1195);
and U3878 (N_3878,N_1318,N_184);
nand U3879 (N_3879,N_41,N_1638);
xnor U3880 (N_3880,N_280,N_859);
xnor U3881 (N_3881,N_970,N_819);
nand U3882 (N_3882,N_860,N_1241);
nand U3883 (N_3883,N_1982,N_336);
xor U3884 (N_3884,N_718,N_712);
nand U3885 (N_3885,N_1606,N_263);
or U3886 (N_3886,N_786,N_71);
nand U3887 (N_3887,N_1027,N_865);
and U3888 (N_3888,N_279,N_822);
or U3889 (N_3889,N_436,N_1053);
nand U3890 (N_3890,N_1411,N_1380);
or U3891 (N_3891,N_627,N_1453);
xor U3892 (N_3892,N_1448,N_717);
nand U3893 (N_3893,N_862,N_824);
nor U3894 (N_3894,N_1888,N_404);
or U3895 (N_3895,N_1932,N_1817);
nand U3896 (N_3896,N_0,N_1279);
nand U3897 (N_3897,N_1836,N_290);
nor U3898 (N_3898,N_1877,N_1129);
nand U3899 (N_3899,N_362,N_1481);
and U3900 (N_3900,N_1907,N_420);
nand U3901 (N_3901,N_795,N_1352);
nand U3902 (N_3902,N_1303,N_1197);
nand U3903 (N_3903,N_215,N_407);
and U3904 (N_3904,N_272,N_1594);
nor U3905 (N_3905,N_16,N_143);
and U3906 (N_3906,N_398,N_280);
or U3907 (N_3907,N_656,N_1924);
nand U3908 (N_3908,N_1503,N_478);
xor U3909 (N_3909,N_1927,N_94);
nand U3910 (N_3910,N_254,N_1247);
nand U3911 (N_3911,N_897,N_291);
nand U3912 (N_3912,N_169,N_1887);
or U3913 (N_3913,N_495,N_462);
and U3914 (N_3914,N_965,N_972);
or U3915 (N_3915,N_742,N_1445);
nor U3916 (N_3916,N_112,N_1910);
xor U3917 (N_3917,N_104,N_1533);
xnor U3918 (N_3918,N_453,N_1561);
and U3919 (N_3919,N_884,N_878);
or U3920 (N_3920,N_1724,N_1127);
nand U3921 (N_3921,N_435,N_225);
nand U3922 (N_3922,N_1603,N_738);
and U3923 (N_3923,N_837,N_1666);
or U3924 (N_3924,N_1959,N_1072);
nor U3925 (N_3925,N_1584,N_522);
and U3926 (N_3926,N_605,N_80);
and U3927 (N_3927,N_272,N_1728);
xnor U3928 (N_3928,N_526,N_1665);
nand U3929 (N_3929,N_848,N_0);
nor U3930 (N_3930,N_220,N_118);
or U3931 (N_3931,N_308,N_1595);
nor U3932 (N_3932,N_434,N_1294);
and U3933 (N_3933,N_1865,N_1271);
and U3934 (N_3934,N_803,N_120);
nand U3935 (N_3935,N_1211,N_1392);
nand U3936 (N_3936,N_526,N_618);
nand U3937 (N_3937,N_764,N_33);
xor U3938 (N_3938,N_700,N_1170);
nand U3939 (N_3939,N_369,N_990);
or U3940 (N_3940,N_1485,N_439);
or U3941 (N_3941,N_1426,N_837);
and U3942 (N_3942,N_262,N_1988);
nor U3943 (N_3943,N_1643,N_553);
nor U3944 (N_3944,N_1895,N_1581);
and U3945 (N_3945,N_1437,N_1403);
xnor U3946 (N_3946,N_715,N_1583);
and U3947 (N_3947,N_529,N_411);
or U3948 (N_3948,N_501,N_1402);
or U3949 (N_3949,N_1310,N_717);
or U3950 (N_3950,N_222,N_485);
nand U3951 (N_3951,N_372,N_1978);
nor U3952 (N_3952,N_692,N_63);
nor U3953 (N_3953,N_1823,N_1077);
nor U3954 (N_3954,N_593,N_492);
and U3955 (N_3955,N_260,N_1302);
nand U3956 (N_3956,N_1904,N_502);
and U3957 (N_3957,N_1062,N_79);
nand U3958 (N_3958,N_1033,N_635);
and U3959 (N_3959,N_482,N_1491);
or U3960 (N_3960,N_1206,N_1615);
nor U3961 (N_3961,N_1736,N_461);
nand U3962 (N_3962,N_1751,N_1191);
and U3963 (N_3963,N_1963,N_1176);
or U3964 (N_3964,N_598,N_488);
or U3965 (N_3965,N_160,N_720);
or U3966 (N_3966,N_421,N_1461);
nor U3967 (N_3967,N_1118,N_507);
nand U3968 (N_3968,N_631,N_433);
nor U3969 (N_3969,N_1033,N_1696);
nand U3970 (N_3970,N_1303,N_1767);
and U3971 (N_3971,N_317,N_224);
nor U3972 (N_3972,N_1198,N_771);
xnor U3973 (N_3973,N_1703,N_826);
and U3974 (N_3974,N_376,N_1522);
nand U3975 (N_3975,N_1244,N_1097);
nand U3976 (N_3976,N_1569,N_422);
xor U3977 (N_3977,N_1705,N_1879);
xnor U3978 (N_3978,N_315,N_730);
nand U3979 (N_3979,N_110,N_438);
or U3980 (N_3980,N_884,N_1587);
or U3981 (N_3981,N_454,N_1032);
or U3982 (N_3982,N_31,N_962);
and U3983 (N_3983,N_1721,N_707);
and U3984 (N_3984,N_1505,N_1950);
and U3985 (N_3985,N_1749,N_1121);
xor U3986 (N_3986,N_70,N_108);
nor U3987 (N_3987,N_552,N_643);
nor U3988 (N_3988,N_1729,N_1627);
xor U3989 (N_3989,N_1079,N_906);
xnor U3990 (N_3990,N_1555,N_1259);
nor U3991 (N_3991,N_878,N_869);
nor U3992 (N_3992,N_663,N_679);
nor U3993 (N_3993,N_385,N_1643);
xnor U3994 (N_3994,N_1077,N_196);
and U3995 (N_3995,N_747,N_1908);
and U3996 (N_3996,N_213,N_379);
xor U3997 (N_3997,N_71,N_1015);
or U3998 (N_3998,N_198,N_1905);
and U3999 (N_3999,N_1274,N_1108);
nand U4000 (N_4000,N_3894,N_2161);
xnor U4001 (N_4001,N_2034,N_2255);
nand U4002 (N_4002,N_3554,N_2741);
xor U4003 (N_4003,N_2253,N_2261);
and U4004 (N_4004,N_2274,N_3816);
nor U4005 (N_4005,N_3908,N_2493);
or U4006 (N_4006,N_3099,N_2409);
and U4007 (N_4007,N_3448,N_3662);
xor U4008 (N_4008,N_2656,N_3735);
or U4009 (N_4009,N_3836,N_2170);
nand U4010 (N_4010,N_3486,N_3502);
and U4011 (N_4011,N_3244,N_2003);
nor U4012 (N_4012,N_3074,N_2878);
xor U4013 (N_4013,N_2452,N_2421);
and U4014 (N_4014,N_2084,N_2527);
and U4015 (N_4015,N_3699,N_2224);
xnor U4016 (N_4016,N_3854,N_3346);
or U4017 (N_4017,N_3784,N_3593);
nand U4018 (N_4018,N_3056,N_3451);
nor U4019 (N_4019,N_3700,N_3557);
and U4020 (N_4020,N_3417,N_3209);
or U4021 (N_4021,N_2806,N_2987);
nor U4022 (N_4022,N_2174,N_2047);
nand U4023 (N_4023,N_3691,N_3131);
or U4024 (N_4024,N_2761,N_3727);
and U4025 (N_4025,N_2635,N_2734);
nor U4026 (N_4026,N_3479,N_3634);
nand U4027 (N_4027,N_2980,N_3145);
nand U4028 (N_4028,N_2881,N_3198);
or U4029 (N_4029,N_2615,N_3420);
and U4030 (N_4030,N_2554,N_3200);
nand U4031 (N_4031,N_2584,N_2521);
or U4032 (N_4032,N_3339,N_3967);
nand U4033 (N_4033,N_2233,N_3891);
and U4034 (N_4034,N_2422,N_2115);
or U4035 (N_4035,N_2473,N_2925);
nor U4036 (N_4036,N_3710,N_2279);
nor U4037 (N_4037,N_3280,N_2860);
nand U4038 (N_4038,N_3228,N_2789);
and U4039 (N_4039,N_2348,N_3819);
nand U4040 (N_4040,N_3302,N_3000);
or U4041 (N_4041,N_2306,N_3626);
or U4042 (N_4042,N_2549,N_2378);
xor U4043 (N_4043,N_2616,N_3912);
and U4044 (N_4044,N_2623,N_3284);
and U4045 (N_4045,N_3064,N_2105);
nor U4046 (N_4046,N_2686,N_3273);
nand U4047 (N_4047,N_2198,N_2964);
nor U4048 (N_4048,N_2710,N_3948);
or U4049 (N_4049,N_3919,N_2642);
nor U4050 (N_4050,N_2441,N_2829);
or U4051 (N_4051,N_3324,N_2337);
nand U4052 (N_4052,N_3125,N_3372);
nor U4053 (N_4053,N_3184,N_2858);
xor U4054 (N_4054,N_3680,N_2329);
nor U4055 (N_4055,N_2703,N_2309);
or U4056 (N_4056,N_2842,N_2499);
nand U4057 (N_4057,N_2326,N_2978);
and U4058 (N_4058,N_3872,N_2235);
and U4059 (N_4059,N_2366,N_3437);
and U4060 (N_4060,N_2672,N_3380);
or U4061 (N_4061,N_2577,N_2874);
and U4062 (N_4062,N_2677,N_3647);
and U4063 (N_4063,N_3589,N_2974);
or U4064 (N_4064,N_2924,N_2432);
and U4065 (N_4065,N_3797,N_2598);
nor U4066 (N_4066,N_2230,N_2317);
or U4067 (N_4067,N_3938,N_2712);
nor U4068 (N_4068,N_2190,N_3286);
nand U4069 (N_4069,N_3134,N_2620);
nand U4070 (N_4070,N_3195,N_3594);
nand U4071 (N_4071,N_2334,N_3164);
and U4072 (N_4072,N_2485,N_3500);
nand U4073 (N_4073,N_2681,N_2475);
nand U4074 (N_4074,N_2424,N_2026);
and U4075 (N_4075,N_2423,N_3325);
nor U4076 (N_4076,N_2088,N_2377);
xnor U4077 (N_4077,N_2655,N_2061);
xnor U4078 (N_4078,N_2612,N_3965);
and U4079 (N_4079,N_2833,N_3254);
or U4080 (N_4080,N_2639,N_3588);
nand U4081 (N_4081,N_2060,N_2586);
and U4082 (N_4082,N_2533,N_2567);
or U4083 (N_4083,N_3600,N_2123);
nor U4084 (N_4084,N_3845,N_3535);
or U4085 (N_4085,N_2178,N_2213);
and U4086 (N_4086,N_3037,N_3107);
nand U4087 (N_4087,N_2665,N_2205);
nand U4088 (N_4088,N_2937,N_2495);
nand U4089 (N_4089,N_3030,N_2585);
and U4090 (N_4090,N_2217,N_3127);
nor U4091 (N_4091,N_3016,N_2621);
nand U4092 (N_4092,N_3736,N_2905);
nor U4093 (N_4093,N_3641,N_2376);
and U4094 (N_4094,N_3860,N_3987);
and U4095 (N_4095,N_3213,N_2315);
and U4096 (N_4096,N_2735,N_3459);
or U4097 (N_4097,N_2831,N_3211);
and U4098 (N_4098,N_2406,N_2919);
xnor U4099 (N_4099,N_3690,N_2759);
xnor U4100 (N_4100,N_3330,N_3876);
nand U4101 (N_4101,N_3875,N_2625);
nor U4102 (N_4102,N_2752,N_2263);
and U4103 (N_4103,N_2412,N_2374);
nor U4104 (N_4104,N_2595,N_3068);
xor U4105 (N_4105,N_3087,N_2965);
xor U4106 (N_4106,N_2573,N_2512);
nand U4107 (N_4107,N_2393,N_2888);
nor U4108 (N_4108,N_3676,N_3970);
or U4109 (N_4109,N_3091,N_3288);
or U4110 (N_4110,N_2242,N_2568);
nand U4111 (N_4111,N_3017,N_2040);
nand U4112 (N_4112,N_3899,N_3985);
or U4113 (N_4113,N_2469,N_2841);
or U4114 (N_4114,N_2877,N_3962);
xnor U4115 (N_4115,N_3115,N_2617);
nand U4116 (N_4116,N_2767,N_3260);
nor U4117 (N_4117,N_3586,N_3309);
nor U4118 (N_4118,N_2226,N_2962);
and U4119 (N_4119,N_2561,N_2870);
nor U4120 (N_4120,N_2117,N_3685);
xnor U4121 (N_4121,N_2151,N_3754);
or U4122 (N_4122,N_3665,N_2289);
or U4123 (N_4123,N_3999,N_3666);
nor U4124 (N_4124,N_3078,N_2085);
and U4125 (N_4125,N_2222,N_3842);
or U4126 (N_4126,N_2529,N_3981);
or U4127 (N_4127,N_3823,N_3106);
and U4128 (N_4128,N_2094,N_3674);
nand U4129 (N_4129,N_3864,N_3751);
or U4130 (N_4130,N_2514,N_2748);
nand U4131 (N_4131,N_2975,N_2323);
and U4132 (N_4132,N_2551,N_3896);
nand U4133 (N_4133,N_2508,N_3971);
nand U4134 (N_4134,N_2572,N_2254);
or U4135 (N_4135,N_2520,N_3282);
nand U4136 (N_4136,N_2845,N_3397);
or U4137 (N_4137,N_3765,N_3522);
and U4138 (N_4138,N_3436,N_3222);
and U4139 (N_4139,N_2774,N_3455);
xor U4140 (N_4140,N_3974,N_2375);
and U4141 (N_4141,N_2714,N_3454);
xor U4142 (N_4142,N_3098,N_3250);
nand U4143 (N_4143,N_3741,N_3543);
nor U4144 (N_4144,N_2792,N_3932);
and U4145 (N_4145,N_2679,N_2737);
nand U4146 (N_4146,N_2384,N_3314);
and U4147 (N_4147,N_2356,N_3568);
nand U4148 (N_4148,N_3749,N_2398);
nand U4149 (N_4149,N_3539,N_3722);
or U4150 (N_4150,N_2054,N_3572);
nor U4151 (N_4151,N_3713,N_3161);
and U4152 (N_4152,N_2697,N_3524);
or U4153 (N_4153,N_2405,N_2654);
or U4154 (N_4154,N_2588,N_3728);
nand U4155 (N_4155,N_3959,N_3954);
and U4156 (N_4156,N_2451,N_3995);
or U4157 (N_4157,N_3423,N_3060);
and U4158 (N_4158,N_3071,N_2608);
nor U4159 (N_4159,N_3787,N_3780);
nor U4160 (N_4160,N_2918,N_2211);
nand U4161 (N_4161,N_2536,N_2091);
and U4162 (N_4162,N_2401,N_2304);
nand U4163 (N_4163,N_3677,N_2130);
nor U4164 (N_4164,N_2180,N_2004);
nand U4165 (N_4165,N_3988,N_3224);
or U4166 (N_4166,N_3259,N_2808);
or U4167 (N_4167,N_3367,N_2185);
and U4168 (N_4168,N_2866,N_2717);
nand U4169 (N_4169,N_2603,N_3581);
nor U4170 (N_4170,N_2597,N_2660);
or U4171 (N_4171,N_3483,N_2044);
nand U4172 (N_4172,N_2576,N_2896);
nor U4173 (N_4173,N_3705,N_3384);
and U4174 (N_4174,N_3698,N_2943);
nand U4175 (N_4175,N_3857,N_3430);
xnor U4176 (N_4176,N_2383,N_3345);
nand U4177 (N_4177,N_3612,N_3824);
xor U4178 (N_4178,N_2388,N_3267);
and U4179 (N_4179,N_2435,N_2641);
and U4180 (N_4180,N_3412,N_3587);
and U4181 (N_4181,N_2020,N_3838);
xnor U4182 (N_4182,N_3445,N_2191);
nand U4183 (N_4183,N_2522,N_3117);
xor U4184 (N_4184,N_2619,N_3435);
nor U4185 (N_4185,N_3122,N_3553);
or U4186 (N_4186,N_2966,N_3584);
nand U4187 (N_4187,N_3208,N_3050);
nor U4188 (N_4188,N_2815,N_2555);
nand U4189 (N_4189,N_2777,N_3047);
or U4190 (N_4190,N_2601,N_2327);
nor U4191 (N_4191,N_3968,N_3811);
nand U4192 (N_4192,N_2515,N_2682);
or U4193 (N_4193,N_3807,N_3510);
or U4194 (N_4194,N_2359,N_2360);
nor U4195 (N_4195,N_2313,N_2237);
nor U4196 (N_4196,N_3444,N_2241);
or U4197 (N_4197,N_2025,N_3310);
xnor U4198 (N_4198,N_2019,N_3810);
nand U4199 (N_4199,N_2364,N_2751);
nand U4200 (N_4200,N_2922,N_3015);
or U4201 (N_4201,N_3373,N_2702);
and U4202 (N_4202,N_2935,N_3179);
nor U4203 (N_4203,N_3137,N_3307);
nor U4204 (N_4204,N_2893,N_2556);
or U4205 (N_4205,N_3177,N_2442);
nor U4206 (N_4206,N_3979,N_3764);
and U4207 (N_4207,N_2238,N_2208);
and U4208 (N_4208,N_2780,N_2753);
nor U4209 (N_4209,N_3365,N_3389);
nor U4210 (N_4210,N_2016,N_2622);
or U4211 (N_4211,N_3591,N_3269);
nor U4212 (N_4212,N_3348,N_3359);
nor U4213 (N_4213,N_2387,N_2219);
and U4214 (N_4214,N_2855,N_3742);
nand U4215 (N_4215,N_2221,N_2290);
nor U4216 (N_4216,N_3206,N_3619);
and U4217 (N_4217,N_2914,N_3096);
and U4218 (N_4218,N_2370,N_2179);
nand U4219 (N_4219,N_3799,N_2611);
or U4220 (N_4220,N_3172,N_3242);
or U4221 (N_4221,N_3093,N_3322);
and U4222 (N_4222,N_3453,N_2143);
or U4223 (N_4223,N_2769,N_2827);
nor U4224 (N_4224,N_3283,N_3388);
or U4225 (N_4225,N_3418,N_3048);
nor U4226 (N_4226,N_3475,N_2590);
and U4227 (N_4227,N_2535,N_3083);
nand U4228 (N_4228,N_3993,N_2828);
or U4229 (N_4229,N_3303,N_2504);
or U4230 (N_4230,N_3731,N_2429);
and U4231 (N_4231,N_2784,N_3154);
nor U4232 (N_4232,N_3776,N_2911);
nand U4233 (N_4233,N_3419,N_2743);
nand U4234 (N_4234,N_3667,N_2122);
nand U4235 (N_4235,N_2981,N_2357);
nand U4236 (N_4236,N_3792,N_3552);
nand U4237 (N_4237,N_3396,N_3187);
nor U4238 (N_4238,N_3934,N_2381);
nand U4239 (N_4239,N_2813,N_2256);
nor U4240 (N_4240,N_3333,N_3318);
nor U4241 (N_4241,N_2407,N_3602);
and U4242 (N_4242,N_2781,N_2927);
or U4243 (N_4243,N_3212,N_3529);
and U4244 (N_4244,N_3752,N_2444);
xnor U4245 (N_4245,N_2474,N_2145);
xnor U4246 (N_4246,N_2229,N_2252);
and U4247 (N_4247,N_2873,N_2571);
and U4248 (N_4248,N_2605,N_2404);
nand U4249 (N_4249,N_3920,N_2899);
nor U4250 (N_4250,N_3001,N_3852);
nand U4251 (N_4251,N_2022,N_3334);
and U4252 (N_4252,N_3051,N_2156);
or U4253 (N_4253,N_2671,N_2129);
and U4254 (N_4254,N_3331,N_2402);
and U4255 (N_4255,N_2299,N_3121);
nor U4256 (N_4256,N_2725,N_3519);
and U4257 (N_4257,N_2167,N_3230);
and U4258 (N_4258,N_2417,N_2760);
and U4259 (N_4259,N_2394,N_3844);
or U4260 (N_4260,N_2148,N_3335);
xor U4261 (N_4261,N_2644,N_3110);
nor U4262 (N_4262,N_3077,N_3404);
nor U4263 (N_4263,N_2455,N_3936);
or U4264 (N_4264,N_2107,N_3013);
nor U4265 (N_4265,N_2552,N_3781);
nor U4266 (N_4266,N_2318,N_3471);
and U4267 (N_4267,N_3571,N_2258);
nor U4268 (N_4268,N_2321,N_3723);
nand U4269 (N_4269,N_3942,N_2545);
or U4270 (N_4270,N_2168,N_3977);
xnor U4271 (N_4271,N_3002,N_3748);
nand U4272 (N_4272,N_2463,N_2108);
nand U4273 (N_4273,N_2645,N_2562);
and U4274 (N_4274,N_2745,N_3009);
nand U4275 (N_4275,N_3075,N_3018);
or U4276 (N_4276,N_2816,N_2494);
nor U4277 (N_4277,N_3923,N_3336);
nand U4278 (N_4278,N_2472,N_3186);
nor U4279 (N_4279,N_3049,N_2723);
and U4280 (N_4280,N_3140,N_2102);
nand U4281 (N_4281,N_2465,N_2443);
and U4282 (N_4282,N_2915,N_3544);
or U4283 (N_4283,N_2868,N_2668);
or U4284 (N_4284,N_2786,N_2064);
nand U4285 (N_4285,N_2872,N_3065);
nand U4286 (N_4286,N_2270,N_3344);
nor U4287 (N_4287,N_2204,N_3827);
nor U4288 (N_4288,N_3306,N_3785);
or U4289 (N_4289,N_2311,N_3944);
xor U4290 (N_4290,N_3608,N_3234);
nor U4291 (N_4291,N_3243,N_3003);
nor U4292 (N_4292,N_3277,N_3489);
or U4293 (N_4293,N_2320,N_2667);
nand U4294 (N_4294,N_2430,N_2453);
and U4295 (N_4295,N_2691,N_3966);
nand U4296 (N_4296,N_3498,N_3614);
nor U4297 (N_4297,N_2916,N_2719);
nor U4298 (N_4298,N_2236,N_2754);
xnor U4299 (N_4299,N_2464,N_3036);
and U4300 (N_4300,N_3462,N_2477);
nor U4301 (N_4301,N_3627,N_2460);
and U4302 (N_4302,N_3173,N_3364);
nor U4303 (N_4303,N_2343,N_3300);
and U4304 (N_4304,N_3235,N_2142);
and U4305 (N_4305,N_3007,N_2166);
nor U4306 (N_4306,N_3452,N_2822);
nand U4307 (N_4307,N_3887,N_2125);
and U4308 (N_4308,N_2507,N_2673);
nand U4309 (N_4309,N_2373,N_2581);
and U4310 (N_4310,N_2209,N_2250);
or U4311 (N_4311,N_3055,N_2534);
and U4312 (N_4312,N_2724,N_3375);
or U4313 (N_4313,N_3290,N_2192);
nand U4314 (N_4314,N_2438,N_2565);
and U4315 (N_4315,N_3343,N_3381);
nor U4316 (N_4316,N_2969,N_2251);
nand U4317 (N_4317,N_3879,N_3762);
and U4318 (N_4318,N_2103,N_3616);
nand U4319 (N_4319,N_3889,N_3661);
and U4320 (N_4320,N_2196,N_3080);
xnor U4321 (N_4321,N_2248,N_3996);
nand U4322 (N_4322,N_3382,N_3814);
nor U4323 (N_4323,N_3621,N_3658);
and U4324 (N_4324,N_2910,N_3297);
or U4325 (N_4325,N_2324,N_2303);
nand U4326 (N_4326,N_2014,N_2150);
nand U4327 (N_4327,N_3292,N_2807);
nor U4328 (N_4328,N_2067,N_2368);
xnor U4329 (N_4329,N_3426,N_2092);
nor U4330 (N_4330,N_3928,N_2292);
and U4331 (N_4331,N_2403,N_3856);
nor U4332 (N_4332,N_2550,N_2693);
or U4333 (N_4333,N_2481,N_2502);
nor U4334 (N_4334,N_3193,N_3265);
and U4335 (N_4335,N_2716,N_3983);
or U4336 (N_4336,N_3880,N_3246);
or U4337 (N_4337,N_2247,N_2880);
xor U4338 (N_4338,N_3969,N_3538);
nand U4339 (N_4339,N_2037,N_2835);
nand U4340 (N_4340,N_2901,N_3513);
nor U4341 (N_4341,N_2766,N_3841);
nor U4342 (N_4342,N_2995,N_2482);
and U4343 (N_4343,N_3255,N_3405);
or U4344 (N_4344,N_3644,N_3984);
nand U4345 (N_4345,N_3044,N_3369);
and U4346 (N_4346,N_2232,N_2503);
or U4347 (N_4347,N_2649,N_3561);
and U4348 (N_4348,N_3102,N_2342);
nor U4349 (N_4349,N_2532,N_3394);
nand U4350 (N_4350,N_3090,N_3374);
nor U4351 (N_4351,N_2264,N_2923);
nor U4352 (N_4352,N_3668,N_3566);
nand U4353 (N_4353,N_2476,N_3356);
nor U4354 (N_4354,N_3155,N_2498);
or U4355 (N_4355,N_3066,N_2856);
nor U4356 (N_4356,N_2811,N_2566);
nand U4357 (N_4357,N_3555,N_3663);
and U4358 (N_4358,N_3832,N_3181);
or U4359 (N_4359,N_2570,N_2834);
or U4360 (N_4360,N_3848,N_3963);
nor U4361 (N_4361,N_2269,N_2553);
and U4362 (N_4362,N_3415,N_2763);
xor U4363 (N_4363,N_3769,N_2750);
nand U4364 (N_4364,N_2967,N_2670);
nand U4365 (N_4365,N_2903,N_3960);
xor U4366 (N_4366,N_3101,N_3358);
or U4367 (N_4367,N_2659,N_3694);
nand U4368 (N_4368,N_3238,N_2963);
nand U4369 (N_4369,N_2904,N_2713);
or U4370 (N_4370,N_2518,N_2846);
or U4371 (N_4371,N_3601,N_2266);
nand U4372 (N_4372,N_2116,N_2489);
nand U4373 (N_4373,N_2852,N_3756);
nand U4374 (N_4374,N_2731,N_3081);
nand U4375 (N_4375,N_3393,N_3463);
nor U4376 (N_4376,N_3596,N_2193);
or U4377 (N_4377,N_3032,N_3688);
nor U4378 (N_4378,N_2462,N_3360);
nor U4379 (N_4379,N_3192,N_2948);
xor U4380 (N_4380,N_2316,N_2281);
nor U4381 (N_4381,N_3025,N_2330);
and U4382 (N_4382,N_3625,N_3103);
and U4383 (N_4383,N_3472,N_2450);
xor U4384 (N_4384,N_3576,N_2559);
nand U4385 (N_4385,N_3556,N_2996);
nor U4386 (N_4386,N_2257,N_3682);
nor U4387 (N_4387,N_2528,N_3693);
and U4388 (N_4388,N_2413,N_3877);
nand U4389 (N_4389,N_2804,N_2991);
nand U4390 (N_4390,N_2669,N_3189);
or U4391 (N_4391,N_3109,N_3329);
nor U4392 (N_4392,N_2484,N_3862);
nand U4393 (N_4393,N_3327,N_2207);
nand U4394 (N_4394,N_3350,N_2971);
or U4395 (N_4395,N_2121,N_3416);
nand U4396 (N_4396,N_2613,N_2272);
and U4397 (N_4397,N_2500,N_3028);
nand U4398 (N_4398,N_3760,N_3499);
or U4399 (N_4399,N_3817,N_2496);
or U4400 (N_4400,N_3903,N_3818);
or U4401 (N_4401,N_3869,N_3153);
and U4402 (N_4402,N_3672,N_3162);
or U4403 (N_4403,N_3905,N_2945);
and U4404 (N_4404,N_2887,N_3537);
or U4405 (N_4405,N_3163,N_2560);
and U4406 (N_4406,N_3266,N_3460);
or U4407 (N_4407,N_3620,N_2081);
or U4408 (N_4408,N_2159,N_3505);
and U4409 (N_4409,N_3684,N_2200);
and U4410 (N_4410,N_3005,N_2291);
xor U4411 (N_4411,N_2517,N_2640);
and U4412 (N_4412,N_3709,N_2839);
and U4413 (N_4413,N_3871,N_3158);
or U4414 (N_4414,N_3440,N_3205);
nand U4415 (N_4415,N_3149,N_3402);
nor U4416 (N_4416,N_3400,N_3136);
nor U4417 (N_4417,N_3809,N_2140);
nand U4418 (N_4418,N_2956,N_2575);
xor U4419 (N_4419,N_2853,N_3795);
and U4420 (N_4420,N_3227,N_3716);
nand U4421 (N_4421,N_3395,N_3223);
nor U4422 (N_4422,N_3095,N_2867);
nand U4423 (N_4423,N_2810,N_2414);
and U4424 (N_4424,N_3245,N_3918);
nor U4425 (N_4425,N_3403,N_3421);
and U4426 (N_4426,N_2931,N_2280);
xnor U4427 (N_4427,N_2859,N_2696);
nand U4428 (N_4428,N_2847,N_2580);
nor U4429 (N_4429,N_2596,N_2341);
and U4430 (N_4430,N_3837,N_3886);
nor U4431 (N_4431,N_2764,N_2689);
nor U4432 (N_4432,N_3449,N_2920);
or U4433 (N_4433,N_3635,N_3916);
and U4434 (N_4434,N_2591,N_3387);
nand U4435 (N_4435,N_3994,N_3947);
nand U4436 (N_4436,N_3738,N_3564);
nand U4437 (N_4437,N_3116,N_3111);
and U4438 (N_4438,N_2801,N_2283);
nand U4439 (N_4439,N_2483,N_3020);
and U4440 (N_4440,N_2706,N_2814);
nand U4441 (N_4441,N_2926,N_2411);
nor U4442 (N_4442,N_2433,N_3835);
and U4443 (N_4443,N_3517,N_3520);
or U4444 (N_4444,N_2415,N_2799);
and U4445 (N_4445,N_3484,N_3704);
nor U4446 (N_4446,N_3160,N_2038);
nand U4447 (N_4447,N_3829,N_2961);
nor U4448 (N_4448,N_3045,N_2643);
or U4449 (N_4449,N_2154,N_3536);
and U4450 (N_4450,N_3450,N_3933);
and U4451 (N_4451,N_2039,N_3683);
nand U4452 (N_4452,N_3560,N_3915);
and U4453 (N_4453,N_2346,N_2757);
and U4454 (N_4454,N_3431,N_3138);
and U4455 (N_4455,N_2467,N_3910);
and U4456 (N_4456,N_3401,N_2011);
and U4457 (N_4457,N_3800,N_2787);
nor U4458 (N_4458,N_2440,N_3058);
and U4459 (N_4459,N_2095,N_2069);
nor U4460 (N_4460,N_2297,N_3907);
xor U4461 (N_4461,N_2400,N_3441);
or U4462 (N_4462,N_2891,N_3258);
nand U4463 (N_4463,N_2097,N_2066);
nor U4464 (N_4464,N_3174,N_3474);
nand U4465 (N_4465,N_3806,N_3312);
or U4466 (N_4466,N_2803,N_3866);
nand U4467 (N_4467,N_2036,N_3660);
and U4468 (N_4468,N_3305,N_3196);
nor U4469 (N_4469,N_3642,N_3465);
nor U4470 (N_4470,N_2583,N_2322);
nor U4471 (N_4471,N_3038,N_2371);
nor U4472 (N_4472,N_3457,N_2854);
or U4473 (N_4473,N_2307,N_3317);
nor U4474 (N_4474,N_3681,N_2942);
xnor U4475 (N_4475,N_3152,N_2558);
and U4476 (N_4476,N_2052,N_3812);
nor U4477 (N_4477,N_2369,N_3408);
or U4478 (N_4478,N_2820,N_3469);
or U4479 (N_4479,N_2135,N_3008);
nand U4480 (N_4480,N_3826,N_3755);
nand U4481 (N_4481,N_2073,N_3574);
nor U4482 (N_4482,N_2086,N_2126);
nand U4483 (N_4483,N_3446,N_3308);
and U4484 (N_4484,N_3104,N_2933);
and U4485 (N_4485,N_2694,N_2875);
nor U4486 (N_4486,N_2758,N_2998);
xnor U4487 (N_4487,N_3178,N_2162);
nor U4488 (N_4488,N_3914,N_2007);
and U4489 (N_4489,N_2138,N_2990);
nor U4490 (N_4490,N_2218,N_3029);
nand U4491 (N_4491,N_3758,N_3183);
or U4492 (N_4492,N_3893,N_3467);
and U4493 (N_4493,N_3708,N_2090);
nor U4494 (N_4494,N_2246,N_2361);
and U4495 (N_4495,N_3113,N_2898);
xor U4496 (N_4496,N_3833,N_3147);
nand U4497 (N_4497,N_3386,N_3262);
nand U4498 (N_4498,N_3873,N_2249);
and U4499 (N_4499,N_3248,N_2487);
nand U4500 (N_4500,N_2711,N_2325);
nor U4501 (N_4501,N_2685,N_3692);
and U4502 (N_4502,N_2530,N_3654);
xnor U4503 (N_4503,N_3157,N_3617);
xnor U4504 (N_4504,N_3531,N_2053);
or U4505 (N_4505,N_2546,N_3883);
xor U4506 (N_4506,N_3295,N_2187);
or U4507 (N_4507,N_3257,N_2788);
or U4508 (N_4508,N_2663,N_3805);
nor U4509 (N_4509,N_2486,N_3802);
nand U4510 (N_4510,N_2825,N_2812);
nor U4511 (N_4511,N_2111,N_3014);
and U4512 (N_4512,N_3379,N_2946);
nor U4513 (N_4513,N_3707,N_3820);
nor U4514 (N_4514,N_3130,N_3126);
and U4515 (N_4515,N_3629,N_2785);
or U4516 (N_4516,N_2906,N_2220);
nand U4517 (N_4517,N_3411,N_3937);
nand U4518 (N_4518,N_3711,N_3233);
nand U4519 (N_4519,N_2890,N_3034);
nand U4520 (N_4520,N_2349,N_3719);
xor U4521 (N_4521,N_2794,N_2305);
nand U4522 (N_4522,N_2118,N_2652);
nor U4523 (N_4523,N_2626,N_2390);
or U4524 (N_4524,N_2772,N_3926);
and U4525 (N_4525,N_2186,N_2296);
nand U4526 (N_4526,N_2100,N_2077);
and U4527 (N_4527,N_2199,N_2516);
nand U4528 (N_4528,N_3291,N_2594);
xnor U4529 (N_4529,N_3461,N_3207);
and U4530 (N_4530,N_2680,N_2968);
xor U4531 (N_4531,N_3825,N_3882);
nor U4532 (N_4532,N_3263,N_2312);
and U4533 (N_4533,N_2079,N_3767);
or U4534 (N_4534,N_3583,N_2314);
or U4535 (N_4535,N_2295,N_3424);
nand U4536 (N_4536,N_2797,N_3225);
or U4537 (N_4537,N_2756,N_3429);
nor U4538 (N_4538,N_2944,N_3547);
nand U4539 (N_4539,N_3664,N_2049);
or U4540 (N_4540,N_2372,N_2796);
and U4541 (N_4541,N_3390,N_3689);
nor U4542 (N_4542,N_3362,N_2439);
or U4543 (N_4543,N_3226,N_3311);
xor U4544 (N_4544,N_3956,N_3830);
and U4545 (N_4545,N_2240,N_3532);
nor U4546 (N_4546,N_3900,N_2093);
or U4547 (N_4547,N_2634,N_3464);
and U4548 (N_4548,N_2675,N_2068);
or U4549 (N_4549,N_2164,N_3961);
nor U4550 (N_4550,N_3898,N_3821);
nand U4551 (N_4551,N_3112,N_3219);
nand U4552 (N_4552,N_3342,N_2354);
nor U4553 (N_4553,N_3046,N_3801);
nand U4554 (N_4554,N_2865,N_3851);
nor U4555 (N_4555,N_3427,N_2087);
nand U4556 (N_4556,N_3275,N_3782);
xor U4557 (N_4557,N_3846,N_3351);
nor U4558 (N_4558,N_3929,N_2630);
or U4559 (N_4559,N_2447,N_3190);
nand U4560 (N_4560,N_2268,N_2599);
nand U4561 (N_4561,N_2137,N_3957);
nor U4562 (N_4562,N_2153,N_2849);
or U4563 (N_4563,N_3545,N_2287);
nor U4564 (N_4564,N_3582,N_2001);
nand U4565 (N_4565,N_2738,N_3737);
or U4566 (N_4566,N_3953,N_2177);
nor U4567 (N_4567,N_2426,N_2434);
xnor U4568 (N_4568,N_3730,N_2189);
or U4569 (N_4569,N_3328,N_3714);
or U4570 (N_4570,N_2478,N_2173);
or U4571 (N_4571,N_2070,N_2857);
or U4572 (N_4572,N_2993,N_3268);
and U4573 (N_4573,N_2009,N_3012);
nand U4574 (N_4574,N_3470,N_2722);
nand U4575 (N_4575,N_3558,N_2817);
nand U4576 (N_4576,N_3480,N_3338);
and U4577 (N_4577,N_3671,N_3272);
nand U4578 (N_4578,N_2683,N_3563);
nand U4579 (N_4579,N_2033,N_3231);
nor U4580 (N_4580,N_3182,N_3599);
nor U4581 (N_4581,N_2892,N_3442);
and U4582 (N_4582,N_2490,N_2908);
nor U4583 (N_4583,N_2013,N_3170);
xor U4584 (N_4584,N_2885,N_2762);
or U4585 (N_4585,N_2350,N_3019);
nand U4586 (N_4586,N_2479,N_3648);
xnor U4587 (N_4587,N_3636,N_2952);
nand U4588 (N_4588,N_2339,N_2418);
nor U4589 (N_4589,N_3945,N_2973);
or U4590 (N_4590,N_2425,N_2175);
nor U4591 (N_4591,N_3481,N_3482);
xor U4592 (N_4592,N_3287,N_3270);
or U4593 (N_4593,N_3909,N_2770);
nand U4594 (N_4594,N_2984,N_2790);
nor U4595 (N_4595,N_2690,N_2564);
or U4596 (N_4596,N_2106,N_3361);
and U4597 (N_4597,N_3229,N_3180);
nor U4598 (N_4598,N_2146,N_2523);
xor U4599 (N_4599,N_2726,N_3456);
nand U4600 (N_4600,N_2864,N_2894);
xnor U4601 (N_4601,N_2557,N_3950);
nor U4602 (N_4602,N_3240,N_2747);
nor U4603 (N_4603,N_2302,N_2397);
and U4604 (N_4604,N_2282,N_3618);
or U4605 (N_4605,N_2895,N_2277);
and U4606 (N_4606,N_3191,N_3124);
nand U4607 (N_4607,N_2428,N_3370);
and U4608 (N_4608,N_2709,N_3788);
or U4609 (N_4609,N_2940,N_3197);
or U4610 (N_4610,N_2420,N_3946);
nand U4611 (N_4611,N_2132,N_2707);
and U4612 (N_4612,N_2005,N_2960);
and U4613 (N_4613,N_2351,N_2446);
nand U4614 (N_4614,N_3092,N_2692);
or U4615 (N_4615,N_3828,N_3271);
nand U4616 (N_4616,N_2582,N_2184);
nor U4617 (N_4617,N_3108,N_3199);
nor U4618 (N_4618,N_2985,N_2470);
or U4619 (N_4619,N_3725,N_3042);
and U4620 (N_4620,N_2127,N_2171);
nor U4621 (N_4621,N_2739,N_3843);
and U4622 (N_4622,N_3794,N_3503);
and U4623 (N_4623,N_2206,N_3523);
nor U4624 (N_4624,N_3332,N_2970);
nand U4625 (N_4625,N_3930,N_3982);
nand U4626 (N_4626,N_3487,N_3739);
xor U4627 (N_4627,N_3410,N_3043);
or U4628 (N_4628,N_2657,N_2197);
nand U4629 (N_4629,N_3501,N_2744);
and U4630 (N_4630,N_2392,N_3385);
xor U4631 (N_4631,N_2526,N_3085);
or U4632 (N_4632,N_2994,N_3252);
and U4633 (N_4633,N_3855,N_2466);
nand U4634 (N_4634,N_2362,N_2459);
xnor U4635 (N_4635,N_2355,N_3175);
xor U4636 (N_4636,N_2000,N_2631);
nand U4637 (N_4637,N_3696,N_2886);
nor U4638 (N_4638,N_2733,N_2223);
nand U4639 (N_4639,N_2569,N_3239);
or U4640 (N_4640,N_2149,N_3989);
and U4641 (N_4641,N_3204,N_2265);
nand U4642 (N_4642,N_2695,N_2729);
or U4643 (N_4643,N_2848,N_2983);
nor U4644 (N_4644,N_3518,N_3202);
nor U4645 (N_4645,N_2957,N_3632);
or U4646 (N_4646,N_2457,N_2609);
nand U4647 (N_4647,N_3477,N_2203);
or U4648 (N_4648,N_2030,N_2419);
nor U4649 (N_4649,N_3067,N_3118);
nor U4650 (N_4650,N_2461,N_2333);
nor U4651 (N_4651,N_3884,N_3922);
xnor U4652 (N_4652,N_2501,N_3570);
and U4653 (N_4653,N_3789,N_2141);
nand U4654 (N_4654,N_2050,N_3294);
nand U4655 (N_4655,N_3777,N_2055);
and U4656 (N_4656,N_2089,N_3168);
nand U4657 (N_4657,N_3935,N_3673);
and U4658 (N_4658,N_3540,N_3870);
or U4659 (N_4659,N_2826,N_2071);
nand U4660 (N_4660,N_3597,N_3951);
nand U4661 (N_4661,N_2301,N_3203);
and U4662 (N_4662,N_3888,N_3863);
nand U4663 (N_4663,N_3906,N_3434);
and U4664 (N_4664,N_3925,N_3624);
nand U4665 (N_4665,N_3135,N_2636);
and U4666 (N_4666,N_3771,N_2492);
or U4667 (N_4667,N_3761,N_2832);
nand U4668 (N_4668,N_2436,N_2158);
nand U4669 (N_4669,N_3859,N_2531);
or U4670 (N_4670,N_2818,N_2165);
or U4671 (N_4671,N_2410,N_2650);
or U4672 (N_4672,N_3383,N_2687);
nor U4673 (N_4673,N_2900,N_3490);
nor U4674 (N_4674,N_2427,N_3349);
or U4675 (N_4675,N_3488,N_2947);
nor U4676 (N_4676,N_3542,N_3657);
and U4677 (N_4677,N_3337,N_2614);
or U4678 (N_4678,N_3917,N_3023);
xnor U4679 (N_4679,N_3808,N_3119);
and U4680 (N_4680,N_3757,N_3724);
nand U4681 (N_4681,N_3839,N_2367);
or U4682 (N_4682,N_2015,N_2365);
nand U4683 (N_4683,N_2395,N_2104);
nand U4684 (N_4684,N_3990,N_2768);
or U4685 (N_4685,N_3770,N_3494);
nand U4686 (N_4686,N_2921,N_2505);
and U4687 (N_4687,N_3151,N_2982);
and U4688 (N_4688,N_3378,N_3059);
or U4689 (N_4689,N_3167,N_3511);
nand U4690 (N_4690,N_2850,N_3279);
and U4691 (N_4691,N_3541,N_2225);
or U4692 (N_4692,N_2018,N_3628);
and U4693 (N_4693,N_3264,N_3606);
or U4694 (N_4694,N_3366,N_2212);
nor U4695 (N_4695,N_3562,N_2454);
and U4696 (N_4696,N_2228,N_2844);
nor U4697 (N_4697,N_3084,N_3323);
and U4698 (N_4698,N_3850,N_2721);
nor U4699 (N_4699,N_3804,N_3579);
and U4700 (N_4700,N_2524,N_2340);
nor U4701 (N_4701,N_2511,N_3129);
nand U4702 (N_4702,N_3559,N_3123);
xnor U4703 (N_4703,N_2078,N_2979);
nand U4704 (N_4704,N_2732,N_3921);
nand U4705 (N_4705,N_3053,N_2139);
nor U4706 (N_4706,N_2637,N_3637);
or U4707 (N_4707,N_3901,N_3320);
nor U4708 (N_4708,N_2396,N_2331);
or U4709 (N_4709,N_3354,N_2021);
nor U4710 (N_4710,N_2951,N_3316);
nor U4711 (N_4711,N_3675,N_3940);
or U4712 (N_4712,N_3061,N_2949);
nand U4713 (N_4713,N_2661,N_3717);
or U4714 (N_4714,N_3447,N_3409);
or U4715 (N_4715,N_3063,N_3276);
nand U4716 (N_4716,N_3473,N_2157);
and U4717 (N_4717,N_3443,N_2416);
nor U4718 (N_4718,N_2183,N_2271);
nor U4719 (N_4719,N_3210,N_3054);
xnor U4720 (N_4720,N_3089,N_3578);
or U4721 (N_4721,N_3033,N_2862);
or U4722 (N_4722,N_3120,N_2779);
nor U4723 (N_4723,N_2674,N_2389);
nor U4724 (N_4724,N_2497,N_2889);
and U4725 (N_4725,N_3220,N_2798);
nor U4726 (N_4726,N_3858,N_3357);
and U4727 (N_4727,N_3299,N_3340);
and U4728 (N_4728,N_2793,N_3232);
xnor U4729 (N_4729,N_2513,N_3534);
xnor U4730 (N_4730,N_3321,N_2907);
nand U4731 (N_4731,N_3766,N_2783);
nand U4732 (N_4732,N_3815,N_3031);
nand U4733 (N_4733,N_2456,N_2883);
xor U4734 (N_4734,N_3508,N_3721);
or U4735 (N_4735,N_2802,N_2934);
and U4736 (N_4736,N_2163,N_2838);
nand U4737 (N_4737,N_2746,N_2932);
or U4738 (N_4738,N_3772,N_3611);
nand U4739 (N_4739,N_3931,N_3952);
nand U4740 (N_4740,N_3069,N_2210);
nor U4741 (N_4741,N_2468,N_2002);
xor U4742 (N_4742,N_3010,N_2958);
nor U4743 (N_4743,N_2032,N_3251);
nand U4744 (N_4744,N_3249,N_2876);
or U4745 (N_4745,N_2182,N_2736);
nand U4746 (N_4746,N_2063,N_2353);
nand U4747 (N_4747,N_3652,N_2592);
nand U4748 (N_4748,N_2664,N_3169);
and U4749 (N_4749,N_2131,N_3726);
and U4750 (N_4750,N_2632,N_3759);
nor U4751 (N_4751,N_2136,N_2056);
nor U4752 (N_4752,N_2869,N_2579);
and U4753 (N_4753,N_2755,N_2688);
xor U4754 (N_4754,N_2606,N_2134);
and U4755 (N_4755,N_2245,N_3670);
or U4756 (N_4756,N_3530,N_3035);
nor U4757 (N_4757,N_3569,N_2437);
nand U4758 (N_4758,N_3834,N_2300);
nand U4759 (N_4759,N_2941,N_3041);
and U4760 (N_4760,N_2773,N_3215);
nand U4761 (N_4761,N_3148,N_2267);
nor U4762 (N_4762,N_3885,N_3791);
nand U4763 (N_4763,N_2538,N_2658);
nor U4764 (N_4764,N_2871,N_2045);
and U4765 (N_4765,N_3139,N_3633);
nand U4766 (N_4766,N_2589,N_2776);
nor U4767 (N_4767,N_2286,N_2194);
nand U4768 (N_4768,N_2058,N_2188);
or U4769 (N_4769,N_3592,N_2989);
or U4770 (N_4770,N_3902,N_2347);
or U4771 (N_4771,N_2293,N_2048);
and U4772 (N_4772,N_2666,N_3605);
or U4773 (N_4773,N_3094,N_3640);
and U4774 (N_4774,N_2029,N_3607);
nand U4775 (N_4775,N_3298,N_2160);
and U4776 (N_4776,N_2647,N_2231);
nand U4777 (N_4777,N_2791,N_2988);
nor U4778 (N_4778,N_2510,N_3261);
nand U4779 (N_4779,N_3493,N_2540);
nand U4780 (N_4780,N_2152,N_3132);
nand U4781 (N_4781,N_3549,N_3142);
and U4782 (N_4782,N_3750,N_3458);
xnor U4783 (N_4783,N_2074,N_3715);
nor U4784 (N_4784,N_3577,N_3849);
xor U4785 (N_4785,N_3341,N_3057);
and U4786 (N_4786,N_2119,N_3976);
and U4787 (N_4787,N_3088,N_3326);
or U4788 (N_4788,N_3143,N_2954);
or U4789 (N_4789,N_3176,N_3747);
or U4790 (N_4790,N_2491,N_2955);
nand U4791 (N_4791,N_2114,N_3021);
or U4792 (N_4792,N_2358,N_2939);
nor U4793 (N_4793,N_3114,N_2380);
xor U4794 (N_4794,N_2082,N_2547);
and U4795 (N_4795,N_3100,N_2243);
xnor U4796 (N_4796,N_3391,N_2884);
and U4797 (N_4797,N_3504,N_2113);
or U4798 (N_4798,N_2805,N_2449);
nor U4799 (N_4799,N_2042,N_3319);
and U4800 (N_4800,N_2006,N_2031);
nand U4801 (N_4801,N_3604,N_3188);
nand U4802 (N_4802,N_2234,N_2730);
or U4803 (N_4803,N_2275,N_2587);
nand U4804 (N_4804,N_3201,N_3079);
and U4805 (N_4805,N_3639,N_2912);
nor U4806 (N_4806,N_2120,N_3355);
nor U4807 (N_4807,N_2708,N_2147);
xnor U4808 (N_4808,N_3414,N_2997);
or U4809 (N_4809,N_2543,N_3623);
and U4810 (N_4810,N_3986,N_3853);
nor U4811 (N_4811,N_3165,N_3156);
and U4812 (N_4812,N_3194,N_2195);
xnor U4813 (N_4813,N_3006,N_3653);
or U4814 (N_4814,N_3645,N_3775);
and U4815 (N_4815,N_2216,N_3980);
and U4816 (N_4816,N_2972,N_3655);
or U4817 (N_4817,N_3992,N_3955);
and U4818 (N_4818,N_2986,N_3507);
nand U4819 (N_4819,N_3551,N_2929);
and U4820 (N_4820,N_3590,N_2345);
or U4821 (N_4821,N_2509,N_3567);
nor U4822 (N_4822,N_3491,N_2950);
nor U4823 (N_4823,N_3975,N_3285);
nor U4824 (N_4824,N_3368,N_2629);
or U4825 (N_4825,N_3073,N_3973);
nor U4826 (N_4826,N_3546,N_3778);
nand U4827 (N_4827,N_2897,N_3468);
or U4828 (N_4828,N_3941,N_3679);
or U4829 (N_4829,N_3407,N_3528);
and U4830 (N_4830,N_3598,N_2448);
and U4831 (N_4831,N_2699,N_3281);
xor U4832 (N_4832,N_3701,N_3720);
and U4833 (N_4833,N_2740,N_2408);
and U4834 (N_4834,N_2399,N_3363);
nand U4835 (N_4835,N_2101,N_3874);
nor U4836 (N_4836,N_3740,N_2851);
or U4837 (N_4837,N_3144,N_3466);
or U4838 (N_4838,N_2260,N_2057);
and U4839 (N_4839,N_2008,N_3733);
nand U4840 (N_4840,N_2800,N_2959);
xor U4841 (N_4841,N_3687,N_3278);
xor U4842 (N_4842,N_3768,N_2542);
or U4843 (N_4843,N_3506,N_3406);
nand U4844 (N_4844,N_2720,N_2338);
nand U4845 (N_4845,N_3086,N_2836);
nand U4846 (N_4846,N_2928,N_2544);
and U4847 (N_4847,N_2648,N_3656);
nor U4848 (N_4848,N_2936,N_3497);
or U4849 (N_4849,N_2041,N_2109);
nand U4850 (N_4850,N_3039,N_3798);
or U4851 (N_4851,N_3533,N_3743);
nor U4852 (N_4852,N_2308,N_3428);
and U4853 (N_4853,N_2602,N_3432);
nand U4854 (N_4854,N_3911,N_2701);
nand U4855 (N_4855,N_2227,N_3609);
or U4856 (N_4856,N_3425,N_2999);
nand U4857 (N_4857,N_2700,N_3565);
or U4858 (N_4858,N_2010,N_2718);
or U4859 (N_4859,N_3895,N_2600);
and U4860 (N_4860,N_3746,N_2593);
and U4861 (N_4861,N_3159,N_2169);
nand U4862 (N_4862,N_2431,N_2819);
nand U4863 (N_4863,N_2604,N_2099);
xor U4864 (N_4864,N_3550,N_2035);
or U4865 (N_4865,N_2445,N_3734);
or U4866 (N_4866,N_3997,N_2742);
and U4867 (N_4867,N_3585,N_2840);
nor U4868 (N_4868,N_3478,N_2017);
and U4869 (N_4869,N_3398,N_3649);
and U4870 (N_4870,N_2633,N_2976);
or U4871 (N_4871,N_3638,N_3422);
and U4872 (N_4872,N_2075,N_2076);
nand U4873 (N_4873,N_3492,N_3072);
nand U4874 (N_4874,N_2328,N_2574);
and U4875 (N_4875,N_2938,N_3525);
nand U4876 (N_4876,N_2578,N_3631);
nand U4877 (N_4877,N_2319,N_2244);
nor U4878 (N_4878,N_3659,N_2012);
nand U4879 (N_4879,N_2065,N_2386);
nand U4880 (N_4880,N_2181,N_2930);
nand U4881 (N_4881,N_3998,N_3972);
nor U4882 (N_4882,N_2823,N_3289);
and U4883 (N_4883,N_3526,N_2288);
nand U4884 (N_4884,N_3868,N_2676);
nand U4885 (N_4885,N_3439,N_2239);
or U4886 (N_4886,N_3241,N_2953);
nor U4887 (N_4887,N_3897,N_3651);
and U4888 (N_4888,N_2298,N_2110);
nand U4889 (N_4889,N_3548,N_3274);
nor U4890 (N_4890,N_2662,N_2176);
nor U4891 (N_4891,N_2778,N_2765);
nand U4892 (N_4892,N_3573,N_3438);
nand U4893 (N_4893,N_3745,N_3881);
and U4894 (N_4894,N_3128,N_3732);
nand U4895 (N_4895,N_2646,N_3744);
and U4896 (N_4896,N_3718,N_3790);
and U4897 (N_4897,N_2992,N_3595);
and U4898 (N_4898,N_3779,N_2259);
nor U4899 (N_4899,N_3697,N_3706);
or U4900 (N_4900,N_2276,N_3793);
and U4901 (N_4901,N_2294,N_3650);
nand U4902 (N_4902,N_3964,N_3646);
or U4903 (N_4903,N_2628,N_3296);
or U4904 (N_4904,N_2062,N_3613);
and U4905 (N_4905,N_3927,N_2843);
nand U4906 (N_4906,N_2096,N_3786);
and U4907 (N_4907,N_3237,N_3978);
nand U4908 (N_4908,N_2332,N_2363);
or U4909 (N_4909,N_3803,N_3509);
nor U4910 (N_4910,N_2024,N_3763);
or U4911 (N_4911,N_3773,N_3392);
nor U4912 (N_4912,N_3515,N_2379);
nor U4913 (N_4913,N_3024,N_2913);
nand U4914 (N_4914,N_2678,N_3949);
nand U4915 (N_4915,N_3026,N_3301);
nand U4916 (N_4916,N_3783,N_2977);
xnor U4917 (N_4917,N_3890,N_3695);
and U4918 (N_4918,N_3097,N_3729);
xnor U4919 (N_4919,N_3247,N_2352);
nor U4920 (N_4920,N_3753,N_3376);
or U4921 (N_4921,N_2144,N_3377);
and U4922 (N_4922,N_3702,N_3630);
or U4923 (N_4923,N_2155,N_3496);
or U4924 (N_4924,N_2344,N_3221);
or U4925 (N_4925,N_3133,N_2051);
nand U4926 (N_4926,N_2202,N_2215);
nor U4927 (N_4927,N_2861,N_3669);
nand U4928 (N_4928,N_3991,N_2506);
nor U4929 (N_4929,N_2879,N_3433);
and U4930 (N_4930,N_2821,N_2830);
or U4931 (N_4931,N_3146,N_2382);
nand U4932 (N_4932,N_2705,N_2539);
or U4933 (N_4933,N_3413,N_3217);
or U4934 (N_4934,N_3256,N_2124);
xnor U4935 (N_4935,N_3831,N_2809);
xor U4936 (N_4936,N_2262,N_2098);
or U4937 (N_4937,N_3913,N_2610);
nand U4938 (N_4938,N_3304,N_3027);
and U4939 (N_4939,N_2618,N_2607);
nand U4940 (N_4940,N_2684,N_3313);
xor U4941 (N_4941,N_2046,N_3943);
xor U4942 (N_4942,N_3399,N_2043);
nor U4943 (N_4943,N_2284,N_2882);
nor U4944 (N_4944,N_2023,N_3105);
or U4945 (N_4945,N_3580,N_2727);
and U4946 (N_4946,N_3712,N_3171);
or U4947 (N_4947,N_3703,N_2837);
xnor U4948 (N_4948,N_3861,N_2728);
or U4949 (N_4949,N_2201,N_3476);
nand U4950 (N_4950,N_3603,N_2638);
and U4951 (N_4951,N_3840,N_3004);
xor U4952 (N_4952,N_3082,N_3218);
nor U4953 (N_4953,N_2391,N_3062);
nand U4954 (N_4954,N_3040,N_2458);
nand U4955 (N_4955,N_2824,N_3774);
and U4956 (N_4956,N_3575,N_3813);
nand U4957 (N_4957,N_2488,N_3150);
nand U4958 (N_4958,N_3878,N_3185);
and U4959 (N_4959,N_3867,N_3622);
nand U4960 (N_4960,N_3643,N_2480);
or U4961 (N_4961,N_3822,N_3796);
and U4962 (N_4962,N_3347,N_3678);
nand U4963 (N_4963,N_3958,N_3216);
nor U4964 (N_4964,N_2128,N_2214);
nor U4965 (N_4965,N_2653,N_2278);
nor U4966 (N_4966,N_2310,N_2072);
and U4967 (N_4967,N_2651,N_3214);
nand U4968 (N_4968,N_2863,N_3686);
or U4969 (N_4969,N_3516,N_2525);
nor U4970 (N_4970,N_3939,N_2285);
nand U4971 (N_4971,N_2541,N_2471);
or U4972 (N_4972,N_2909,N_2917);
nand U4973 (N_4973,N_3371,N_2083);
or U4974 (N_4974,N_3610,N_2698);
or U4975 (N_4975,N_2112,N_2771);
or U4976 (N_4976,N_2624,N_2172);
xor U4977 (N_4977,N_3892,N_2080);
xor U4978 (N_4978,N_2548,N_3070);
nor U4979 (N_4979,N_2782,N_2027);
and U4980 (N_4980,N_2627,N_2537);
and U4981 (N_4981,N_3293,N_3352);
nor U4982 (N_4982,N_2028,N_2704);
and U4983 (N_4983,N_2902,N_3527);
nand U4984 (N_4984,N_2385,N_3865);
and U4985 (N_4985,N_3495,N_3166);
nand U4986 (N_4986,N_3253,N_2059);
or U4987 (N_4987,N_2519,N_3512);
nand U4988 (N_4988,N_2563,N_2335);
or U4989 (N_4989,N_3485,N_3236);
nand U4990 (N_4990,N_3904,N_3315);
nand U4991 (N_4991,N_3011,N_2133);
xor U4992 (N_4992,N_3514,N_3141);
xnor U4993 (N_4993,N_2715,N_2749);
nor U4994 (N_4994,N_2273,N_3052);
and U4995 (N_4995,N_3847,N_2775);
nand U4996 (N_4996,N_3353,N_2336);
nand U4997 (N_4997,N_3022,N_2795);
nand U4998 (N_4998,N_3076,N_3924);
nand U4999 (N_4999,N_3615,N_3521);
nor U5000 (N_5000,N_2488,N_3770);
nor U5001 (N_5001,N_2751,N_3074);
nor U5002 (N_5002,N_3702,N_2035);
or U5003 (N_5003,N_3515,N_3630);
or U5004 (N_5004,N_2757,N_3808);
xnor U5005 (N_5005,N_2541,N_2644);
and U5006 (N_5006,N_2326,N_2521);
nand U5007 (N_5007,N_3619,N_3836);
and U5008 (N_5008,N_2027,N_2866);
and U5009 (N_5009,N_3399,N_2249);
and U5010 (N_5010,N_3361,N_2703);
or U5011 (N_5011,N_3047,N_3387);
and U5012 (N_5012,N_3982,N_2044);
or U5013 (N_5013,N_2398,N_3037);
nand U5014 (N_5014,N_3835,N_3684);
nor U5015 (N_5015,N_3625,N_2287);
nor U5016 (N_5016,N_2741,N_2742);
nand U5017 (N_5017,N_2153,N_3386);
xor U5018 (N_5018,N_2792,N_2927);
and U5019 (N_5019,N_3984,N_2766);
nor U5020 (N_5020,N_2515,N_2029);
nor U5021 (N_5021,N_2667,N_2794);
nand U5022 (N_5022,N_3106,N_3287);
and U5023 (N_5023,N_2023,N_3012);
nand U5024 (N_5024,N_2662,N_2300);
or U5025 (N_5025,N_2168,N_3466);
nand U5026 (N_5026,N_2841,N_3112);
xor U5027 (N_5027,N_3065,N_2316);
and U5028 (N_5028,N_3947,N_2222);
and U5029 (N_5029,N_2683,N_3785);
and U5030 (N_5030,N_2372,N_3457);
nor U5031 (N_5031,N_2749,N_3837);
or U5032 (N_5032,N_3744,N_2722);
and U5033 (N_5033,N_3074,N_3683);
nand U5034 (N_5034,N_2068,N_2645);
nor U5035 (N_5035,N_3186,N_2631);
and U5036 (N_5036,N_2145,N_2092);
nand U5037 (N_5037,N_3377,N_2466);
xor U5038 (N_5038,N_2236,N_2532);
or U5039 (N_5039,N_2444,N_3168);
or U5040 (N_5040,N_2895,N_3433);
nor U5041 (N_5041,N_3429,N_2141);
nor U5042 (N_5042,N_2337,N_3209);
nor U5043 (N_5043,N_3300,N_3093);
nand U5044 (N_5044,N_2074,N_3342);
and U5045 (N_5045,N_2643,N_2723);
xor U5046 (N_5046,N_2138,N_3796);
nor U5047 (N_5047,N_2110,N_3939);
nand U5048 (N_5048,N_3295,N_2540);
nand U5049 (N_5049,N_2925,N_3286);
nand U5050 (N_5050,N_2117,N_3061);
or U5051 (N_5051,N_2375,N_3012);
nor U5052 (N_5052,N_2204,N_2872);
xnor U5053 (N_5053,N_3614,N_3461);
xor U5054 (N_5054,N_2213,N_2774);
xor U5055 (N_5055,N_3658,N_3124);
nor U5056 (N_5056,N_2114,N_3929);
xor U5057 (N_5057,N_2650,N_2500);
xor U5058 (N_5058,N_3429,N_2147);
or U5059 (N_5059,N_2503,N_3701);
and U5060 (N_5060,N_2270,N_2485);
nor U5061 (N_5061,N_3555,N_3792);
xor U5062 (N_5062,N_3483,N_2968);
and U5063 (N_5063,N_3291,N_3907);
nor U5064 (N_5064,N_2128,N_3193);
or U5065 (N_5065,N_3121,N_3866);
or U5066 (N_5066,N_3428,N_3075);
or U5067 (N_5067,N_3361,N_2429);
nand U5068 (N_5068,N_3047,N_3228);
nand U5069 (N_5069,N_3194,N_2541);
nor U5070 (N_5070,N_3410,N_2612);
or U5071 (N_5071,N_2270,N_3408);
or U5072 (N_5072,N_3639,N_2823);
nor U5073 (N_5073,N_3721,N_2620);
and U5074 (N_5074,N_3223,N_3311);
nand U5075 (N_5075,N_3582,N_3316);
and U5076 (N_5076,N_2689,N_3075);
and U5077 (N_5077,N_2226,N_2791);
and U5078 (N_5078,N_3369,N_3777);
and U5079 (N_5079,N_3982,N_2567);
xor U5080 (N_5080,N_2230,N_2850);
nand U5081 (N_5081,N_3304,N_3598);
nand U5082 (N_5082,N_3147,N_2517);
nor U5083 (N_5083,N_3542,N_2352);
nor U5084 (N_5084,N_2558,N_2253);
nor U5085 (N_5085,N_3497,N_2161);
nand U5086 (N_5086,N_3535,N_3575);
and U5087 (N_5087,N_3058,N_3215);
or U5088 (N_5088,N_3788,N_3024);
or U5089 (N_5089,N_3143,N_3679);
or U5090 (N_5090,N_2179,N_3443);
or U5091 (N_5091,N_3965,N_2067);
nand U5092 (N_5092,N_3064,N_2079);
or U5093 (N_5093,N_3084,N_3313);
nand U5094 (N_5094,N_2292,N_3778);
nand U5095 (N_5095,N_3293,N_3180);
and U5096 (N_5096,N_2287,N_3493);
nand U5097 (N_5097,N_3149,N_3953);
and U5098 (N_5098,N_3927,N_3442);
and U5099 (N_5099,N_3183,N_2035);
or U5100 (N_5100,N_2456,N_2378);
nor U5101 (N_5101,N_2231,N_2649);
and U5102 (N_5102,N_2955,N_3524);
nor U5103 (N_5103,N_2888,N_2102);
nor U5104 (N_5104,N_2826,N_2923);
or U5105 (N_5105,N_2923,N_3320);
and U5106 (N_5106,N_2740,N_2511);
nand U5107 (N_5107,N_2639,N_2410);
nor U5108 (N_5108,N_3750,N_3443);
xnor U5109 (N_5109,N_2710,N_2146);
and U5110 (N_5110,N_2486,N_2221);
nor U5111 (N_5111,N_2504,N_3903);
xnor U5112 (N_5112,N_3177,N_2733);
xnor U5113 (N_5113,N_3809,N_2801);
nor U5114 (N_5114,N_2783,N_2755);
and U5115 (N_5115,N_2795,N_3999);
nor U5116 (N_5116,N_3491,N_3000);
and U5117 (N_5117,N_2822,N_3760);
nand U5118 (N_5118,N_2973,N_2837);
xor U5119 (N_5119,N_2160,N_2500);
xnor U5120 (N_5120,N_2425,N_2508);
nor U5121 (N_5121,N_2020,N_2003);
xnor U5122 (N_5122,N_3810,N_3916);
nand U5123 (N_5123,N_3266,N_2307);
nand U5124 (N_5124,N_3166,N_2625);
nor U5125 (N_5125,N_2731,N_2436);
or U5126 (N_5126,N_2201,N_3138);
nand U5127 (N_5127,N_3539,N_3494);
or U5128 (N_5128,N_2946,N_2492);
or U5129 (N_5129,N_2710,N_3039);
nand U5130 (N_5130,N_3256,N_3251);
and U5131 (N_5131,N_3071,N_3847);
nor U5132 (N_5132,N_3082,N_2841);
nor U5133 (N_5133,N_2562,N_2852);
xnor U5134 (N_5134,N_2886,N_2956);
and U5135 (N_5135,N_3161,N_3916);
xnor U5136 (N_5136,N_2228,N_2414);
or U5137 (N_5137,N_3739,N_3201);
nor U5138 (N_5138,N_2362,N_2215);
xor U5139 (N_5139,N_3513,N_2552);
nand U5140 (N_5140,N_3813,N_2924);
nand U5141 (N_5141,N_3528,N_2699);
nand U5142 (N_5142,N_2716,N_3795);
nand U5143 (N_5143,N_3923,N_2780);
nor U5144 (N_5144,N_3347,N_3557);
nor U5145 (N_5145,N_3029,N_2016);
nor U5146 (N_5146,N_3188,N_2911);
nand U5147 (N_5147,N_3901,N_2747);
and U5148 (N_5148,N_2278,N_3916);
nor U5149 (N_5149,N_2078,N_3352);
nor U5150 (N_5150,N_2716,N_2002);
nand U5151 (N_5151,N_3631,N_2876);
nand U5152 (N_5152,N_2559,N_3083);
nand U5153 (N_5153,N_2701,N_2305);
nor U5154 (N_5154,N_3125,N_2559);
or U5155 (N_5155,N_2914,N_2537);
nor U5156 (N_5156,N_2252,N_2606);
or U5157 (N_5157,N_3421,N_2808);
nand U5158 (N_5158,N_2884,N_3086);
nor U5159 (N_5159,N_3826,N_3625);
nand U5160 (N_5160,N_2401,N_3715);
or U5161 (N_5161,N_2328,N_2652);
nor U5162 (N_5162,N_2664,N_2027);
nor U5163 (N_5163,N_3958,N_3399);
xnor U5164 (N_5164,N_3363,N_2715);
xnor U5165 (N_5165,N_3559,N_3726);
nand U5166 (N_5166,N_2418,N_3579);
nand U5167 (N_5167,N_3248,N_2397);
nand U5168 (N_5168,N_3628,N_3956);
and U5169 (N_5169,N_2135,N_2895);
nand U5170 (N_5170,N_2236,N_2717);
nand U5171 (N_5171,N_3207,N_3617);
and U5172 (N_5172,N_3814,N_3007);
or U5173 (N_5173,N_3731,N_3798);
nand U5174 (N_5174,N_2520,N_3717);
nor U5175 (N_5175,N_2318,N_2518);
nand U5176 (N_5176,N_3764,N_3607);
and U5177 (N_5177,N_2779,N_3704);
nor U5178 (N_5178,N_3819,N_2177);
xnor U5179 (N_5179,N_2526,N_2954);
and U5180 (N_5180,N_2898,N_3309);
or U5181 (N_5181,N_2858,N_3703);
and U5182 (N_5182,N_2576,N_2585);
nor U5183 (N_5183,N_3682,N_2551);
or U5184 (N_5184,N_3978,N_2558);
and U5185 (N_5185,N_2463,N_2410);
and U5186 (N_5186,N_3986,N_3007);
nor U5187 (N_5187,N_3558,N_2579);
and U5188 (N_5188,N_3293,N_2843);
nor U5189 (N_5189,N_2107,N_2828);
nor U5190 (N_5190,N_3067,N_3042);
nor U5191 (N_5191,N_2411,N_3923);
or U5192 (N_5192,N_3669,N_2572);
or U5193 (N_5193,N_2120,N_3584);
and U5194 (N_5194,N_2530,N_2095);
nand U5195 (N_5195,N_3720,N_2687);
or U5196 (N_5196,N_2400,N_2869);
nand U5197 (N_5197,N_3535,N_2000);
or U5198 (N_5198,N_2350,N_2150);
nor U5199 (N_5199,N_2193,N_3348);
nor U5200 (N_5200,N_2699,N_3316);
nand U5201 (N_5201,N_3999,N_2137);
nand U5202 (N_5202,N_2443,N_3402);
nor U5203 (N_5203,N_3886,N_2745);
and U5204 (N_5204,N_2226,N_3554);
nand U5205 (N_5205,N_3775,N_3633);
xor U5206 (N_5206,N_3393,N_2124);
nand U5207 (N_5207,N_3142,N_3483);
and U5208 (N_5208,N_2249,N_3241);
nand U5209 (N_5209,N_2186,N_3937);
or U5210 (N_5210,N_3814,N_2779);
xor U5211 (N_5211,N_3839,N_2103);
nand U5212 (N_5212,N_2654,N_3401);
nor U5213 (N_5213,N_3185,N_2383);
and U5214 (N_5214,N_3089,N_2015);
or U5215 (N_5215,N_2821,N_3989);
and U5216 (N_5216,N_3968,N_2367);
or U5217 (N_5217,N_3026,N_3470);
and U5218 (N_5218,N_3053,N_2213);
or U5219 (N_5219,N_2108,N_3279);
nor U5220 (N_5220,N_3343,N_2025);
nand U5221 (N_5221,N_3775,N_3479);
and U5222 (N_5222,N_3683,N_2337);
nor U5223 (N_5223,N_3677,N_3810);
nor U5224 (N_5224,N_2086,N_3504);
and U5225 (N_5225,N_2343,N_3677);
nand U5226 (N_5226,N_3277,N_3397);
nor U5227 (N_5227,N_2495,N_3746);
and U5228 (N_5228,N_3153,N_2154);
or U5229 (N_5229,N_2131,N_2716);
nor U5230 (N_5230,N_3028,N_2764);
xor U5231 (N_5231,N_2981,N_2888);
nand U5232 (N_5232,N_3383,N_3270);
and U5233 (N_5233,N_2956,N_2547);
or U5234 (N_5234,N_3990,N_2096);
and U5235 (N_5235,N_3294,N_3372);
and U5236 (N_5236,N_2702,N_2443);
or U5237 (N_5237,N_2476,N_3556);
nand U5238 (N_5238,N_2217,N_2719);
and U5239 (N_5239,N_3907,N_3322);
or U5240 (N_5240,N_2723,N_3869);
or U5241 (N_5241,N_2757,N_2200);
and U5242 (N_5242,N_2955,N_3011);
or U5243 (N_5243,N_3956,N_2959);
or U5244 (N_5244,N_3098,N_3353);
and U5245 (N_5245,N_2277,N_2534);
nor U5246 (N_5246,N_2751,N_2197);
nor U5247 (N_5247,N_3284,N_2324);
nor U5248 (N_5248,N_2486,N_3380);
and U5249 (N_5249,N_3321,N_3474);
nor U5250 (N_5250,N_2968,N_3006);
or U5251 (N_5251,N_2349,N_3744);
and U5252 (N_5252,N_3474,N_3074);
xnor U5253 (N_5253,N_2951,N_3872);
and U5254 (N_5254,N_2170,N_3615);
or U5255 (N_5255,N_2993,N_2034);
and U5256 (N_5256,N_2299,N_3411);
nor U5257 (N_5257,N_2166,N_3850);
and U5258 (N_5258,N_2652,N_2731);
or U5259 (N_5259,N_3851,N_2153);
nand U5260 (N_5260,N_3923,N_3227);
nand U5261 (N_5261,N_2075,N_3937);
or U5262 (N_5262,N_3651,N_2084);
and U5263 (N_5263,N_2634,N_3476);
or U5264 (N_5264,N_3852,N_2764);
or U5265 (N_5265,N_3528,N_3150);
nand U5266 (N_5266,N_3717,N_3777);
and U5267 (N_5267,N_3570,N_2298);
or U5268 (N_5268,N_3273,N_2358);
nand U5269 (N_5269,N_2484,N_2704);
nor U5270 (N_5270,N_2346,N_2564);
nor U5271 (N_5271,N_3696,N_2299);
nor U5272 (N_5272,N_3663,N_2576);
nor U5273 (N_5273,N_2260,N_2850);
xor U5274 (N_5274,N_3859,N_2114);
xnor U5275 (N_5275,N_3669,N_3021);
or U5276 (N_5276,N_2332,N_2485);
or U5277 (N_5277,N_3593,N_2567);
or U5278 (N_5278,N_3287,N_3991);
or U5279 (N_5279,N_3821,N_3584);
and U5280 (N_5280,N_2965,N_3010);
nand U5281 (N_5281,N_2807,N_2536);
nor U5282 (N_5282,N_3141,N_3575);
and U5283 (N_5283,N_3428,N_2134);
and U5284 (N_5284,N_3597,N_3084);
and U5285 (N_5285,N_2215,N_2653);
nor U5286 (N_5286,N_3867,N_2635);
or U5287 (N_5287,N_3507,N_2616);
nor U5288 (N_5288,N_3135,N_2524);
nor U5289 (N_5289,N_3775,N_2655);
and U5290 (N_5290,N_3029,N_2279);
nand U5291 (N_5291,N_3708,N_3325);
nor U5292 (N_5292,N_3663,N_2019);
or U5293 (N_5293,N_2145,N_3778);
nand U5294 (N_5294,N_2188,N_2595);
nor U5295 (N_5295,N_2062,N_3718);
nor U5296 (N_5296,N_2956,N_2629);
nand U5297 (N_5297,N_2978,N_2336);
nand U5298 (N_5298,N_3190,N_2472);
or U5299 (N_5299,N_3029,N_2040);
or U5300 (N_5300,N_3574,N_3995);
xnor U5301 (N_5301,N_3511,N_2033);
and U5302 (N_5302,N_2329,N_2034);
nand U5303 (N_5303,N_2847,N_3841);
or U5304 (N_5304,N_2560,N_3840);
nor U5305 (N_5305,N_3152,N_2243);
or U5306 (N_5306,N_3459,N_2670);
xnor U5307 (N_5307,N_3465,N_2012);
and U5308 (N_5308,N_3946,N_3192);
nand U5309 (N_5309,N_2992,N_3664);
and U5310 (N_5310,N_2765,N_2457);
and U5311 (N_5311,N_2030,N_3561);
and U5312 (N_5312,N_2011,N_2582);
xor U5313 (N_5313,N_3128,N_2850);
nand U5314 (N_5314,N_3581,N_2124);
and U5315 (N_5315,N_2052,N_2999);
and U5316 (N_5316,N_2007,N_2919);
nand U5317 (N_5317,N_2174,N_2443);
nor U5318 (N_5318,N_2877,N_2462);
or U5319 (N_5319,N_3245,N_3585);
or U5320 (N_5320,N_3547,N_3443);
nand U5321 (N_5321,N_3410,N_3554);
nand U5322 (N_5322,N_3628,N_3130);
and U5323 (N_5323,N_3043,N_2615);
nand U5324 (N_5324,N_3243,N_3888);
or U5325 (N_5325,N_3526,N_2529);
xor U5326 (N_5326,N_3704,N_3093);
nand U5327 (N_5327,N_2988,N_2817);
nor U5328 (N_5328,N_2977,N_3692);
or U5329 (N_5329,N_3401,N_3002);
nor U5330 (N_5330,N_2372,N_3790);
or U5331 (N_5331,N_2125,N_2087);
nor U5332 (N_5332,N_3326,N_3719);
or U5333 (N_5333,N_3416,N_3848);
and U5334 (N_5334,N_3740,N_3707);
and U5335 (N_5335,N_3809,N_3095);
or U5336 (N_5336,N_3581,N_3882);
or U5337 (N_5337,N_3923,N_3557);
and U5338 (N_5338,N_3075,N_3589);
or U5339 (N_5339,N_3636,N_2188);
nor U5340 (N_5340,N_3499,N_3595);
or U5341 (N_5341,N_2950,N_2574);
nor U5342 (N_5342,N_2619,N_3479);
nand U5343 (N_5343,N_2151,N_2968);
or U5344 (N_5344,N_2021,N_3213);
nor U5345 (N_5345,N_3041,N_3307);
nand U5346 (N_5346,N_3273,N_3227);
and U5347 (N_5347,N_3970,N_2290);
and U5348 (N_5348,N_2093,N_2179);
nand U5349 (N_5349,N_3792,N_3627);
nand U5350 (N_5350,N_3519,N_2213);
nor U5351 (N_5351,N_3316,N_2253);
and U5352 (N_5352,N_2660,N_3775);
nand U5353 (N_5353,N_3496,N_3396);
xor U5354 (N_5354,N_3553,N_3246);
or U5355 (N_5355,N_3799,N_2150);
and U5356 (N_5356,N_3851,N_2589);
and U5357 (N_5357,N_2433,N_2352);
nor U5358 (N_5358,N_3992,N_3601);
nand U5359 (N_5359,N_2457,N_2189);
nand U5360 (N_5360,N_2069,N_3152);
or U5361 (N_5361,N_3212,N_2411);
nand U5362 (N_5362,N_3069,N_2648);
nor U5363 (N_5363,N_2889,N_2228);
nand U5364 (N_5364,N_3738,N_3948);
and U5365 (N_5365,N_3603,N_2335);
nor U5366 (N_5366,N_3553,N_2806);
and U5367 (N_5367,N_3853,N_2407);
or U5368 (N_5368,N_2893,N_2493);
and U5369 (N_5369,N_2599,N_2685);
nand U5370 (N_5370,N_2856,N_2721);
nand U5371 (N_5371,N_2124,N_3675);
nand U5372 (N_5372,N_3856,N_3342);
nor U5373 (N_5373,N_2404,N_3525);
nand U5374 (N_5374,N_3432,N_3951);
nand U5375 (N_5375,N_3596,N_3766);
or U5376 (N_5376,N_3834,N_3697);
xor U5377 (N_5377,N_3902,N_2564);
and U5378 (N_5378,N_2111,N_3517);
nor U5379 (N_5379,N_2765,N_3168);
nor U5380 (N_5380,N_3025,N_3903);
nor U5381 (N_5381,N_3966,N_2663);
or U5382 (N_5382,N_2133,N_3081);
nor U5383 (N_5383,N_3415,N_2627);
nor U5384 (N_5384,N_2345,N_3497);
nor U5385 (N_5385,N_2128,N_3727);
and U5386 (N_5386,N_2891,N_2151);
xor U5387 (N_5387,N_3183,N_2350);
or U5388 (N_5388,N_3968,N_2807);
nand U5389 (N_5389,N_2155,N_2118);
or U5390 (N_5390,N_2436,N_2390);
and U5391 (N_5391,N_2946,N_3772);
nand U5392 (N_5392,N_2571,N_2093);
nor U5393 (N_5393,N_2684,N_3123);
nand U5394 (N_5394,N_3927,N_2894);
or U5395 (N_5395,N_2688,N_3536);
xor U5396 (N_5396,N_3200,N_2319);
or U5397 (N_5397,N_2614,N_2837);
nor U5398 (N_5398,N_3977,N_3133);
nor U5399 (N_5399,N_3607,N_3939);
and U5400 (N_5400,N_2711,N_2855);
nand U5401 (N_5401,N_3205,N_3229);
nor U5402 (N_5402,N_3576,N_2184);
xor U5403 (N_5403,N_2009,N_3511);
nor U5404 (N_5404,N_3180,N_2094);
nand U5405 (N_5405,N_2831,N_3749);
nand U5406 (N_5406,N_2649,N_2929);
and U5407 (N_5407,N_2431,N_2551);
or U5408 (N_5408,N_2101,N_3204);
xor U5409 (N_5409,N_3204,N_2352);
nor U5410 (N_5410,N_3646,N_2287);
or U5411 (N_5411,N_2075,N_3887);
xor U5412 (N_5412,N_2073,N_3018);
and U5413 (N_5413,N_2923,N_2395);
nor U5414 (N_5414,N_2570,N_2928);
nand U5415 (N_5415,N_3088,N_3448);
nand U5416 (N_5416,N_2341,N_2658);
nand U5417 (N_5417,N_3524,N_3189);
and U5418 (N_5418,N_2297,N_2950);
nor U5419 (N_5419,N_2891,N_3509);
nand U5420 (N_5420,N_3093,N_3588);
or U5421 (N_5421,N_2641,N_3201);
nor U5422 (N_5422,N_3225,N_3164);
and U5423 (N_5423,N_3000,N_2622);
xor U5424 (N_5424,N_3847,N_2520);
and U5425 (N_5425,N_3910,N_2663);
nor U5426 (N_5426,N_2735,N_3174);
nand U5427 (N_5427,N_3901,N_2655);
nor U5428 (N_5428,N_3504,N_2159);
and U5429 (N_5429,N_3255,N_3856);
xnor U5430 (N_5430,N_2323,N_2955);
xnor U5431 (N_5431,N_2053,N_2078);
nor U5432 (N_5432,N_2483,N_3502);
nor U5433 (N_5433,N_3135,N_2053);
or U5434 (N_5434,N_2655,N_3158);
nand U5435 (N_5435,N_3871,N_3164);
or U5436 (N_5436,N_3340,N_2926);
xnor U5437 (N_5437,N_3487,N_2284);
and U5438 (N_5438,N_3583,N_3074);
nor U5439 (N_5439,N_3014,N_3570);
nand U5440 (N_5440,N_3893,N_2742);
nand U5441 (N_5441,N_3454,N_2823);
xnor U5442 (N_5442,N_3725,N_2296);
nor U5443 (N_5443,N_2039,N_2007);
nand U5444 (N_5444,N_3998,N_3374);
or U5445 (N_5445,N_2135,N_2784);
nor U5446 (N_5446,N_2741,N_3303);
or U5447 (N_5447,N_3329,N_2851);
nor U5448 (N_5448,N_2795,N_2402);
nor U5449 (N_5449,N_3795,N_3942);
nor U5450 (N_5450,N_3607,N_2671);
nor U5451 (N_5451,N_3539,N_2207);
nor U5452 (N_5452,N_3040,N_3939);
or U5453 (N_5453,N_2742,N_3943);
and U5454 (N_5454,N_2237,N_3085);
and U5455 (N_5455,N_2445,N_2413);
nand U5456 (N_5456,N_2398,N_3096);
or U5457 (N_5457,N_2526,N_3793);
or U5458 (N_5458,N_2374,N_3317);
nor U5459 (N_5459,N_3021,N_2226);
xor U5460 (N_5460,N_3104,N_3546);
or U5461 (N_5461,N_3417,N_3369);
and U5462 (N_5462,N_3859,N_2907);
nand U5463 (N_5463,N_3986,N_2666);
nor U5464 (N_5464,N_3324,N_2968);
or U5465 (N_5465,N_2931,N_2382);
nand U5466 (N_5466,N_3985,N_2542);
nor U5467 (N_5467,N_3167,N_2079);
or U5468 (N_5468,N_2957,N_2422);
or U5469 (N_5469,N_2570,N_2006);
or U5470 (N_5470,N_3393,N_3506);
nor U5471 (N_5471,N_2091,N_3216);
or U5472 (N_5472,N_2407,N_3905);
xor U5473 (N_5473,N_2617,N_3073);
xor U5474 (N_5474,N_3743,N_2087);
nand U5475 (N_5475,N_2035,N_2691);
nand U5476 (N_5476,N_2920,N_3916);
and U5477 (N_5477,N_3968,N_3785);
xnor U5478 (N_5478,N_3739,N_2828);
nor U5479 (N_5479,N_3874,N_3274);
and U5480 (N_5480,N_2220,N_3129);
nor U5481 (N_5481,N_3669,N_2336);
and U5482 (N_5482,N_3931,N_2285);
and U5483 (N_5483,N_2874,N_3119);
nor U5484 (N_5484,N_2788,N_3571);
nand U5485 (N_5485,N_2347,N_3910);
or U5486 (N_5486,N_2797,N_3788);
nand U5487 (N_5487,N_2122,N_2020);
nor U5488 (N_5488,N_2220,N_3230);
nor U5489 (N_5489,N_2220,N_2678);
nor U5490 (N_5490,N_3593,N_3861);
or U5491 (N_5491,N_3721,N_3920);
nand U5492 (N_5492,N_3934,N_2712);
nand U5493 (N_5493,N_3687,N_3249);
and U5494 (N_5494,N_2516,N_2770);
or U5495 (N_5495,N_3187,N_2787);
nand U5496 (N_5496,N_3115,N_3601);
or U5497 (N_5497,N_3991,N_2054);
and U5498 (N_5498,N_2936,N_2670);
nand U5499 (N_5499,N_3176,N_2322);
and U5500 (N_5500,N_2920,N_3498);
nor U5501 (N_5501,N_2070,N_3604);
xor U5502 (N_5502,N_3930,N_2767);
nor U5503 (N_5503,N_2396,N_3971);
and U5504 (N_5504,N_2455,N_3174);
nor U5505 (N_5505,N_2993,N_3720);
and U5506 (N_5506,N_2836,N_3940);
or U5507 (N_5507,N_3929,N_2444);
or U5508 (N_5508,N_3227,N_2902);
and U5509 (N_5509,N_3313,N_2904);
or U5510 (N_5510,N_3523,N_2363);
nand U5511 (N_5511,N_2700,N_2093);
nor U5512 (N_5512,N_2199,N_3112);
xor U5513 (N_5513,N_2553,N_2715);
and U5514 (N_5514,N_3219,N_2223);
or U5515 (N_5515,N_3554,N_2718);
nand U5516 (N_5516,N_3800,N_2172);
and U5517 (N_5517,N_3987,N_2365);
nor U5518 (N_5518,N_3404,N_2976);
nand U5519 (N_5519,N_2538,N_3101);
nor U5520 (N_5520,N_2375,N_2797);
nand U5521 (N_5521,N_3863,N_3421);
and U5522 (N_5522,N_2573,N_2905);
xor U5523 (N_5523,N_3207,N_2777);
nor U5524 (N_5524,N_3155,N_3338);
or U5525 (N_5525,N_3192,N_2809);
nor U5526 (N_5526,N_2227,N_2550);
and U5527 (N_5527,N_2517,N_2385);
nor U5528 (N_5528,N_3038,N_2616);
nor U5529 (N_5529,N_2700,N_2298);
and U5530 (N_5530,N_3577,N_3297);
xor U5531 (N_5531,N_2546,N_3826);
or U5532 (N_5532,N_3856,N_3012);
nor U5533 (N_5533,N_3157,N_2299);
or U5534 (N_5534,N_2400,N_2657);
xor U5535 (N_5535,N_3260,N_3071);
or U5536 (N_5536,N_2010,N_3405);
nand U5537 (N_5537,N_2375,N_3704);
or U5538 (N_5538,N_2696,N_2115);
nand U5539 (N_5539,N_2946,N_2737);
xnor U5540 (N_5540,N_2932,N_3182);
or U5541 (N_5541,N_2442,N_2362);
or U5542 (N_5542,N_2922,N_3403);
or U5543 (N_5543,N_3722,N_3608);
and U5544 (N_5544,N_3120,N_2437);
nand U5545 (N_5545,N_3316,N_3042);
nor U5546 (N_5546,N_3354,N_3139);
xor U5547 (N_5547,N_3781,N_2003);
nand U5548 (N_5548,N_2596,N_3056);
or U5549 (N_5549,N_2713,N_3312);
nand U5550 (N_5550,N_2394,N_3859);
nand U5551 (N_5551,N_3557,N_2415);
nor U5552 (N_5552,N_2491,N_3996);
nand U5553 (N_5553,N_2559,N_2362);
xor U5554 (N_5554,N_3699,N_2893);
or U5555 (N_5555,N_3740,N_3971);
or U5556 (N_5556,N_2276,N_2381);
and U5557 (N_5557,N_2711,N_3938);
nor U5558 (N_5558,N_2925,N_3470);
nand U5559 (N_5559,N_2063,N_3349);
nor U5560 (N_5560,N_2287,N_3682);
or U5561 (N_5561,N_3915,N_2073);
nor U5562 (N_5562,N_3693,N_3830);
nor U5563 (N_5563,N_3990,N_3994);
and U5564 (N_5564,N_2515,N_2273);
and U5565 (N_5565,N_3994,N_3579);
nand U5566 (N_5566,N_2790,N_3994);
nor U5567 (N_5567,N_2336,N_2509);
and U5568 (N_5568,N_3342,N_3865);
nand U5569 (N_5569,N_2230,N_2851);
nor U5570 (N_5570,N_2431,N_3887);
nand U5571 (N_5571,N_2116,N_3715);
nor U5572 (N_5572,N_2234,N_2586);
nor U5573 (N_5573,N_3510,N_3354);
and U5574 (N_5574,N_2689,N_2804);
nand U5575 (N_5575,N_3580,N_3503);
nor U5576 (N_5576,N_2820,N_2476);
nand U5577 (N_5577,N_2949,N_3623);
and U5578 (N_5578,N_3808,N_3005);
and U5579 (N_5579,N_2570,N_3655);
or U5580 (N_5580,N_2264,N_3241);
nand U5581 (N_5581,N_2271,N_2182);
nor U5582 (N_5582,N_2875,N_2460);
nand U5583 (N_5583,N_3972,N_3380);
and U5584 (N_5584,N_3077,N_2947);
nand U5585 (N_5585,N_2464,N_3104);
nand U5586 (N_5586,N_3685,N_2103);
or U5587 (N_5587,N_2088,N_3537);
or U5588 (N_5588,N_3753,N_2736);
nor U5589 (N_5589,N_2890,N_3084);
nand U5590 (N_5590,N_3885,N_3954);
nor U5591 (N_5591,N_2212,N_3856);
or U5592 (N_5592,N_3073,N_2558);
or U5593 (N_5593,N_3983,N_2717);
or U5594 (N_5594,N_3571,N_2570);
or U5595 (N_5595,N_2211,N_3775);
nand U5596 (N_5596,N_3909,N_2357);
and U5597 (N_5597,N_2340,N_2740);
nand U5598 (N_5598,N_2675,N_3448);
or U5599 (N_5599,N_3179,N_3294);
nand U5600 (N_5600,N_2121,N_3039);
nand U5601 (N_5601,N_3306,N_2720);
nor U5602 (N_5602,N_3652,N_3930);
or U5603 (N_5603,N_2272,N_3106);
or U5604 (N_5604,N_2800,N_2696);
or U5605 (N_5605,N_3212,N_3935);
or U5606 (N_5606,N_2058,N_2432);
nor U5607 (N_5607,N_2176,N_3698);
and U5608 (N_5608,N_2006,N_3757);
nor U5609 (N_5609,N_3268,N_2445);
xnor U5610 (N_5610,N_3126,N_3830);
nor U5611 (N_5611,N_2177,N_2234);
or U5612 (N_5612,N_2378,N_3004);
nor U5613 (N_5613,N_3686,N_2318);
and U5614 (N_5614,N_2107,N_2065);
and U5615 (N_5615,N_2947,N_3643);
or U5616 (N_5616,N_2332,N_2138);
and U5617 (N_5617,N_3242,N_2582);
nor U5618 (N_5618,N_3330,N_2799);
nand U5619 (N_5619,N_2401,N_3742);
nand U5620 (N_5620,N_3643,N_3628);
or U5621 (N_5621,N_2832,N_3631);
and U5622 (N_5622,N_2218,N_2964);
nand U5623 (N_5623,N_2349,N_2727);
nor U5624 (N_5624,N_3247,N_3037);
xor U5625 (N_5625,N_2394,N_3934);
or U5626 (N_5626,N_3686,N_3504);
and U5627 (N_5627,N_3676,N_2482);
nor U5628 (N_5628,N_3947,N_3578);
nor U5629 (N_5629,N_3723,N_3933);
and U5630 (N_5630,N_2738,N_2376);
or U5631 (N_5631,N_3927,N_3391);
nor U5632 (N_5632,N_3496,N_2408);
nand U5633 (N_5633,N_3300,N_3042);
or U5634 (N_5634,N_2325,N_2910);
nor U5635 (N_5635,N_2249,N_3663);
nand U5636 (N_5636,N_3961,N_3419);
nand U5637 (N_5637,N_2813,N_3527);
nand U5638 (N_5638,N_2040,N_2536);
and U5639 (N_5639,N_2851,N_2658);
or U5640 (N_5640,N_3757,N_2311);
nor U5641 (N_5641,N_2608,N_2103);
or U5642 (N_5642,N_3542,N_3073);
nand U5643 (N_5643,N_2050,N_3462);
nor U5644 (N_5644,N_3915,N_2241);
nand U5645 (N_5645,N_3004,N_2236);
and U5646 (N_5646,N_2856,N_2114);
nor U5647 (N_5647,N_3403,N_3641);
and U5648 (N_5648,N_3471,N_3926);
nor U5649 (N_5649,N_2755,N_3894);
nand U5650 (N_5650,N_2187,N_2095);
or U5651 (N_5651,N_2490,N_3473);
xnor U5652 (N_5652,N_2536,N_3073);
xor U5653 (N_5653,N_2699,N_2037);
nand U5654 (N_5654,N_3100,N_2405);
and U5655 (N_5655,N_2799,N_2285);
nand U5656 (N_5656,N_2303,N_3652);
and U5657 (N_5657,N_2686,N_2459);
nor U5658 (N_5658,N_2507,N_3920);
or U5659 (N_5659,N_3227,N_2572);
or U5660 (N_5660,N_2978,N_2355);
nand U5661 (N_5661,N_2756,N_3391);
or U5662 (N_5662,N_2955,N_3573);
xnor U5663 (N_5663,N_2166,N_3884);
nor U5664 (N_5664,N_3351,N_3754);
xnor U5665 (N_5665,N_2042,N_2529);
nor U5666 (N_5666,N_3479,N_3884);
xnor U5667 (N_5667,N_2374,N_3557);
nand U5668 (N_5668,N_3036,N_3534);
and U5669 (N_5669,N_2447,N_3328);
nand U5670 (N_5670,N_2960,N_3429);
or U5671 (N_5671,N_3866,N_3657);
or U5672 (N_5672,N_2451,N_2923);
and U5673 (N_5673,N_3142,N_2645);
nor U5674 (N_5674,N_2588,N_2797);
or U5675 (N_5675,N_2479,N_2869);
and U5676 (N_5676,N_3972,N_2272);
nand U5677 (N_5677,N_2554,N_2393);
or U5678 (N_5678,N_3637,N_2133);
or U5679 (N_5679,N_2004,N_2425);
or U5680 (N_5680,N_2615,N_3822);
nand U5681 (N_5681,N_2456,N_2023);
nand U5682 (N_5682,N_3146,N_2946);
nor U5683 (N_5683,N_3341,N_2763);
nor U5684 (N_5684,N_2621,N_2294);
xnor U5685 (N_5685,N_2429,N_3266);
nand U5686 (N_5686,N_3947,N_2704);
nand U5687 (N_5687,N_2052,N_2731);
or U5688 (N_5688,N_2646,N_3709);
and U5689 (N_5689,N_3837,N_2377);
nand U5690 (N_5690,N_3929,N_2900);
and U5691 (N_5691,N_2989,N_2093);
and U5692 (N_5692,N_3882,N_3275);
nand U5693 (N_5693,N_3967,N_3170);
nand U5694 (N_5694,N_2373,N_3769);
nand U5695 (N_5695,N_2630,N_3682);
nand U5696 (N_5696,N_2439,N_2334);
nand U5697 (N_5697,N_3199,N_2438);
nand U5698 (N_5698,N_3364,N_2923);
xnor U5699 (N_5699,N_3903,N_2204);
nor U5700 (N_5700,N_2700,N_3851);
nand U5701 (N_5701,N_2600,N_3199);
or U5702 (N_5702,N_3352,N_3298);
and U5703 (N_5703,N_2585,N_2341);
nand U5704 (N_5704,N_3819,N_2396);
nor U5705 (N_5705,N_2601,N_2503);
and U5706 (N_5706,N_3954,N_3502);
nor U5707 (N_5707,N_3216,N_3227);
nand U5708 (N_5708,N_3383,N_2823);
nand U5709 (N_5709,N_3089,N_3239);
and U5710 (N_5710,N_2533,N_2498);
nor U5711 (N_5711,N_3813,N_3441);
xor U5712 (N_5712,N_2333,N_3874);
and U5713 (N_5713,N_2861,N_3324);
nand U5714 (N_5714,N_2838,N_3601);
nand U5715 (N_5715,N_3956,N_2893);
and U5716 (N_5716,N_3771,N_2709);
or U5717 (N_5717,N_3946,N_3991);
nor U5718 (N_5718,N_3770,N_2952);
nand U5719 (N_5719,N_3521,N_2063);
or U5720 (N_5720,N_3773,N_2721);
nand U5721 (N_5721,N_3200,N_2035);
nand U5722 (N_5722,N_3946,N_2535);
nand U5723 (N_5723,N_3785,N_2361);
nand U5724 (N_5724,N_3257,N_2660);
and U5725 (N_5725,N_3150,N_2281);
or U5726 (N_5726,N_3867,N_3272);
or U5727 (N_5727,N_3914,N_3212);
or U5728 (N_5728,N_2379,N_3424);
and U5729 (N_5729,N_2078,N_2654);
nand U5730 (N_5730,N_2780,N_2956);
or U5731 (N_5731,N_2696,N_3618);
nor U5732 (N_5732,N_2605,N_2392);
xor U5733 (N_5733,N_2015,N_3275);
nand U5734 (N_5734,N_3364,N_3743);
nand U5735 (N_5735,N_2156,N_2462);
nand U5736 (N_5736,N_2736,N_3686);
nor U5737 (N_5737,N_2021,N_3504);
and U5738 (N_5738,N_2008,N_3113);
and U5739 (N_5739,N_3441,N_2568);
or U5740 (N_5740,N_3554,N_3025);
nand U5741 (N_5741,N_3253,N_3360);
nor U5742 (N_5742,N_3567,N_3307);
xor U5743 (N_5743,N_2179,N_2097);
or U5744 (N_5744,N_3402,N_2961);
or U5745 (N_5745,N_2656,N_3305);
nor U5746 (N_5746,N_2711,N_3207);
nand U5747 (N_5747,N_3386,N_3588);
nand U5748 (N_5748,N_2582,N_2642);
or U5749 (N_5749,N_3475,N_2777);
nand U5750 (N_5750,N_2088,N_2527);
nor U5751 (N_5751,N_2159,N_2326);
nor U5752 (N_5752,N_2339,N_3875);
or U5753 (N_5753,N_2590,N_2603);
nand U5754 (N_5754,N_3644,N_3191);
nor U5755 (N_5755,N_3229,N_2876);
and U5756 (N_5756,N_3600,N_3639);
and U5757 (N_5757,N_3938,N_2763);
nor U5758 (N_5758,N_3487,N_3025);
xor U5759 (N_5759,N_3812,N_2456);
xnor U5760 (N_5760,N_3027,N_2458);
and U5761 (N_5761,N_2347,N_3815);
or U5762 (N_5762,N_2781,N_2390);
or U5763 (N_5763,N_2820,N_3511);
and U5764 (N_5764,N_2184,N_3524);
and U5765 (N_5765,N_3253,N_3910);
nor U5766 (N_5766,N_3122,N_3176);
nor U5767 (N_5767,N_3745,N_3593);
nor U5768 (N_5768,N_2156,N_2802);
and U5769 (N_5769,N_2694,N_2126);
or U5770 (N_5770,N_2377,N_2108);
xnor U5771 (N_5771,N_2709,N_3304);
xor U5772 (N_5772,N_3566,N_3093);
nor U5773 (N_5773,N_2078,N_2775);
nor U5774 (N_5774,N_3703,N_2153);
nor U5775 (N_5775,N_3012,N_2588);
nand U5776 (N_5776,N_3973,N_2167);
xor U5777 (N_5777,N_2833,N_2290);
nand U5778 (N_5778,N_3514,N_3336);
nor U5779 (N_5779,N_2118,N_2059);
xnor U5780 (N_5780,N_3274,N_2861);
or U5781 (N_5781,N_2765,N_3040);
and U5782 (N_5782,N_3868,N_3710);
nand U5783 (N_5783,N_3648,N_2762);
nand U5784 (N_5784,N_3233,N_2312);
nand U5785 (N_5785,N_2062,N_3180);
nand U5786 (N_5786,N_3114,N_2894);
and U5787 (N_5787,N_3770,N_2227);
nor U5788 (N_5788,N_2464,N_2936);
or U5789 (N_5789,N_2469,N_2325);
nand U5790 (N_5790,N_2964,N_2997);
nand U5791 (N_5791,N_2222,N_3426);
nor U5792 (N_5792,N_2055,N_3274);
and U5793 (N_5793,N_2734,N_3782);
nand U5794 (N_5794,N_2309,N_3003);
and U5795 (N_5795,N_3203,N_2924);
or U5796 (N_5796,N_2532,N_3853);
xor U5797 (N_5797,N_2745,N_3133);
and U5798 (N_5798,N_3124,N_2892);
and U5799 (N_5799,N_2391,N_2690);
nor U5800 (N_5800,N_2079,N_2182);
and U5801 (N_5801,N_2786,N_2738);
or U5802 (N_5802,N_3476,N_3866);
xor U5803 (N_5803,N_3417,N_3468);
and U5804 (N_5804,N_3097,N_3787);
and U5805 (N_5805,N_2763,N_3179);
or U5806 (N_5806,N_3957,N_3184);
xor U5807 (N_5807,N_2182,N_2939);
nor U5808 (N_5808,N_2678,N_3788);
nand U5809 (N_5809,N_2765,N_2280);
xnor U5810 (N_5810,N_3444,N_2700);
or U5811 (N_5811,N_2716,N_2729);
nand U5812 (N_5812,N_2488,N_2087);
xor U5813 (N_5813,N_3456,N_2738);
nor U5814 (N_5814,N_3501,N_3197);
nand U5815 (N_5815,N_2768,N_2322);
nand U5816 (N_5816,N_2341,N_3686);
or U5817 (N_5817,N_2577,N_3660);
or U5818 (N_5818,N_2780,N_2606);
and U5819 (N_5819,N_3377,N_3382);
and U5820 (N_5820,N_3202,N_2321);
nor U5821 (N_5821,N_3119,N_3446);
nand U5822 (N_5822,N_3571,N_2861);
nor U5823 (N_5823,N_2510,N_2808);
and U5824 (N_5824,N_2227,N_3870);
nand U5825 (N_5825,N_3416,N_3280);
nor U5826 (N_5826,N_3283,N_3660);
nor U5827 (N_5827,N_2367,N_2163);
nor U5828 (N_5828,N_2052,N_3371);
nand U5829 (N_5829,N_2371,N_3492);
nor U5830 (N_5830,N_3394,N_2737);
nand U5831 (N_5831,N_3965,N_3119);
nand U5832 (N_5832,N_3575,N_2144);
nor U5833 (N_5833,N_3590,N_3105);
nor U5834 (N_5834,N_3233,N_2970);
or U5835 (N_5835,N_2033,N_2798);
and U5836 (N_5836,N_3779,N_2807);
or U5837 (N_5837,N_3927,N_2668);
nand U5838 (N_5838,N_3570,N_2911);
and U5839 (N_5839,N_2431,N_2541);
xor U5840 (N_5840,N_3053,N_2461);
and U5841 (N_5841,N_3690,N_3347);
and U5842 (N_5842,N_2394,N_2320);
nor U5843 (N_5843,N_2441,N_2951);
nand U5844 (N_5844,N_2590,N_3741);
or U5845 (N_5845,N_3202,N_3809);
or U5846 (N_5846,N_2059,N_2421);
nand U5847 (N_5847,N_2888,N_3093);
or U5848 (N_5848,N_2452,N_3229);
nor U5849 (N_5849,N_3775,N_2886);
nand U5850 (N_5850,N_3546,N_3530);
nor U5851 (N_5851,N_2542,N_2816);
nor U5852 (N_5852,N_2993,N_3917);
and U5853 (N_5853,N_3264,N_3453);
nor U5854 (N_5854,N_3948,N_2776);
or U5855 (N_5855,N_3201,N_2605);
and U5856 (N_5856,N_2350,N_2792);
nand U5857 (N_5857,N_3363,N_2307);
nand U5858 (N_5858,N_3859,N_3717);
nand U5859 (N_5859,N_2233,N_3428);
nand U5860 (N_5860,N_3045,N_2954);
nor U5861 (N_5861,N_2260,N_2185);
or U5862 (N_5862,N_3751,N_3895);
nor U5863 (N_5863,N_2847,N_2170);
nand U5864 (N_5864,N_3490,N_3644);
and U5865 (N_5865,N_2010,N_3944);
and U5866 (N_5866,N_2976,N_3123);
and U5867 (N_5867,N_2478,N_2026);
nand U5868 (N_5868,N_3908,N_3913);
and U5869 (N_5869,N_2703,N_2550);
nand U5870 (N_5870,N_2592,N_2294);
and U5871 (N_5871,N_2233,N_2084);
or U5872 (N_5872,N_2828,N_3820);
or U5873 (N_5873,N_2042,N_3110);
xor U5874 (N_5874,N_3059,N_3458);
or U5875 (N_5875,N_2942,N_3326);
nor U5876 (N_5876,N_3882,N_3044);
and U5877 (N_5877,N_2701,N_3692);
nor U5878 (N_5878,N_2620,N_2997);
nor U5879 (N_5879,N_3230,N_3327);
or U5880 (N_5880,N_3838,N_2324);
or U5881 (N_5881,N_3988,N_2599);
and U5882 (N_5882,N_3828,N_3266);
xor U5883 (N_5883,N_3648,N_2816);
and U5884 (N_5884,N_2874,N_3598);
or U5885 (N_5885,N_3917,N_2402);
or U5886 (N_5886,N_3811,N_3450);
nor U5887 (N_5887,N_2580,N_3612);
xor U5888 (N_5888,N_3353,N_2687);
or U5889 (N_5889,N_2649,N_3243);
or U5890 (N_5890,N_3003,N_3785);
nand U5891 (N_5891,N_2008,N_3537);
and U5892 (N_5892,N_2933,N_2861);
nand U5893 (N_5893,N_3338,N_3417);
xnor U5894 (N_5894,N_3930,N_3696);
nor U5895 (N_5895,N_3495,N_3187);
or U5896 (N_5896,N_3852,N_3866);
and U5897 (N_5897,N_2268,N_3945);
nor U5898 (N_5898,N_3435,N_2315);
and U5899 (N_5899,N_2575,N_3832);
or U5900 (N_5900,N_2663,N_2399);
nor U5901 (N_5901,N_3356,N_2088);
xnor U5902 (N_5902,N_3710,N_3147);
and U5903 (N_5903,N_2445,N_3860);
nand U5904 (N_5904,N_2663,N_2981);
nand U5905 (N_5905,N_3289,N_3102);
or U5906 (N_5906,N_2111,N_2130);
or U5907 (N_5907,N_2828,N_3978);
nor U5908 (N_5908,N_3704,N_2776);
or U5909 (N_5909,N_3595,N_3987);
nand U5910 (N_5910,N_2218,N_3238);
or U5911 (N_5911,N_3252,N_3455);
nand U5912 (N_5912,N_2872,N_3733);
or U5913 (N_5913,N_2187,N_2018);
nand U5914 (N_5914,N_3941,N_3238);
and U5915 (N_5915,N_3603,N_2149);
or U5916 (N_5916,N_2133,N_2395);
xnor U5917 (N_5917,N_2837,N_2922);
and U5918 (N_5918,N_2850,N_2233);
nand U5919 (N_5919,N_3743,N_2852);
or U5920 (N_5920,N_2604,N_3966);
nand U5921 (N_5921,N_3828,N_3026);
and U5922 (N_5922,N_3160,N_2818);
or U5923 (N_5923,N_2947,N_2451);
xnor U5924 (N_5924,N_2029,N_2380);
nand U5925 (N_5925,N_2429,N_2332);
xor U5926 (N_5926,N_3444,N_2385);
nor U5927 (N_5927,N_3497,N_3243);
or U5928 (N_5928,N_2658,N_2800);
nand U5929 (N_5929,N_2725,N_3013);
nor U5930 (N_5930,N_3406,N_2999);
xnor U5931 (N_5931,N_3047,N_3176);
and U5932 (N_5932,N_2542,N_2710);
nor U5933 (N_5933,N_2685,N_2377);
nand U5934 (N_5934,N_2159,N_2862);
or U5935 (N_5935,N_2211,N_2944);
nor U5936 (N_5936,N_2938,N_2279);
nand U5937 (N_5937,N_2927,N_2081);
and U5938 (N_5938,N_2449,N_2365);
nor U5939 (N_5939,N_2689,N_2725);
nand U5940 (N_5940,N_3218,N_3901);
nor U5941 (N_5941,N_3659,N_2049);
or U5942 (N_5942,N_2826,N_2958);
nor U5943 (N_5943,N_3551,N_3999);
nand U5944 (N_5944,N_3870,N_3587);
nand U5945 (N_5945,N_2816,N_3908);
and U5946 (N_5946,N_3091,N_3305);
nor U5947 (N_5947,N_3079,N_3988);
nor U5948 (N_5948,N_3698,N_2291);
nand U5949 (N_5949,N_2846,N_2449);
nor U5950 (N_5950,N_2489,N_2182);
xor U5951 (N_5951,N_3991,N_2653);
or U5952 (N_5952,N_2981,N_3204);
and U5953 (N_5953,N_3599,N_2160);
or U5954 (N_5954,N_3076,N_2857);
xnor U5955 (N_5955,N_3314,N_3406);
nor U5956 (N_5956,N_3237,N_3521);
xnor U5957 (N_5957,N_2076,N_3665);
nand U5958 (N_5958,N_2719,N_3036);
xnor U5959 (N_5959,N_2615,N_3985);
and U5960 (N_5960,N_3954,N_2224);
and U5961 (N_5961,N_3333,N_3001);
nand U5962 (N_5962,N_2128,N_2144);
and U5963 (N_5963,N_2931,N_2626);
nor U5964 (N_5964,N_2620,N_2251);
xnor U5965 (N_5965,N_2970,N_3516);
nor U5966 (N_5966,N_3524,N_2082);
or U5967 (N_5967,N_3314,N_2385);
nor U5968 (N_5968,N_2811,N_2616);
nand U5969 (N_5969,N_3201,N_2783);
nor U5970 (N_5970,N_3364,N_3248);
and U5971 (N_5971,N_3810,N_3765);
or U5972 (N_5972,N_2936,N_3130);
nand U5973 (N_5973,N_3004,N_3183);
nor U5974 (N_5974,N_2502,N_2832);
nor U5975 (N_5975,N_3555,N_3324);
xnor U5976 (N_5976,N_3004,N_2879);
xnor U5977 (N_5977,N_3716,N_2068);
or U5978 (N_5978,N_2402,N_3358);
or U5979 (N_5979,N_3642,N_3056);
and U5980 (N_5980,N_3182,N_2313);
and U5981 (N_5981,N_2688,N_3527);
and U5982 (N_5982,N_3109,N_2850);
or U5983 (N_5983,N_3754,N_3418);
and U5984 (N_5984,N_2299,N_2221);
and U5985 (N_5985,N_3054,N_3362);
or U5986 (N_5986,N_3547,N_2114);
and U5987 (N_5987,N_2786,N_3074);
or U5988 (N_5988,N_2670,N_3085);
nor U5989 (N_5989,N_3123,N_2234);
nor U5990 (N_5990,N_2255,N_2684);
and U5991 (N_5991,N_2237,N_3388);
nor U5992 (N_5992,N_2493,N_3600);
or U5993 (N_5993,N_3323,N_3132);
xor U5994 (N_5994,N_3481,N_3242);
xnor U5995 (N_5995,N_3141,N_3488);
xor U5996 (N_5996,N_3534,N_2727);
nor U5997 (N_5997,N_2221,N_2939);
nor U5998 (N_5998,N_3767,N_2586);
or U5999 (N_5999,N_2034,N_2028);
and U6000 (N_6000,N_5426,N_5003);
and U6001 (N_6001,N_4296,N_5414);
nor U6002 (N_6002,N_5261,N_5918);
and U6003 (N_6003,N_4375,N_4225);
nor U6004 (N_6004,N_4095,N_4114);
or U6005 (N_6005,N_4731,N_4641);
and U6006 (N_6006,N_4917,N_5260);
xnor U6007 (N_6007,N_4297,N_4987);
and U6008 (N_6008,N_4629,N_5388);
nand U6009 (N_6009,N_4436,N_4285);
and U6010 (N_6010,N_5509,N_4312);
nand U6011 (N_6011,N_5544,N_5104);
or U6012 (N_6012,N_5617,N_4728);
and U6013 (N_6013,N_4486,N_5836);
or U6014 (N_6014,N_4730,N_5114);
nand U6015 (N_6015,N_4282,N_5208);
nand U6016 (N_6016,N_5341,N_4462);
nand U6017 (N_6017,N_4125,N_4997);
nor U6018 (N_6018,N_4549,N_4659);
and U6019 (N_6019,N_4678,N_5151);
nand U6020 (N_6020,N_5355,N_4603);
and U6021 (N_6021,N_4460,N_5259);
nand U6022 (N_6022,N_4372,N_5646);
nor U6023 (N_6023,N_4623,N_4769);
nor U6024 (N_6024,N_4409,N_5204);
and U6025 (N_6025,N_5771,N_5135);
or U6026 (N_6026,N_4216,N_5267);
and U6027 (N_6027,N_4976,N_5116);
nand U6028 (N_6028,N_5143,N_4373);
and U6029 (N_6029,N_5699,N_4410);
and U6030 (N_6030,N_4964,N_4100);
and U6031 (N_6031,N_4147,N_5438);
or U6032 (N_6032,N_5644,N_4653);
or U6033 (N_6033,N_5896,N_4136);
nand U6034 (N_6034,N_4990,N_5036);
nand U6035 (N_6035,N_5560,N_5867);
or U6036 (N_6036,N_4243,N_4040);
nor U6037 (N_6037,N_4760,N_4129);
or U6038 (N_6038,N_5307,N_5422);
and U6039 (N_6039,N_4039,N_4433);
and U6040 (N_6040,N_4308,N_5590);
nand U6041 (N_6041,N_4176,N_5684);
xor U6042 (N_6042,N_4566,N_5978);
nand U6043 (N_6043,N_5427,N_5323);
and U6044 (N_6044,N_5049,N_5753);
nor U6045 (N_6045,N_4933,N_5606);
nor U6046 (N_6046,N_4194,N_5374);
or U6047 (N_6047,N_5488,N_4657);
and U6048 (N_6048,N_4547,N_4891);
nor U6049 (N_6049,N_4610,N_5121);
nand U6050 (N_6050,N_5213,N_5304);
or U6051 (N_6051,N_4576,N_4041);
or U6052 (N_6052,N_5481,N_5639);
and U6053 (N_6053,N_4759,N_4271);
nor U6054 (N_6054,N_5976,N_5894);
and U6055 (N_6055,N_4071,N_5674);
nand U6056 (N_6056,N_5608,N_4713);
nor U6057 (N_6057,N_4890,N_4859);
nor U6058 (N_6058,N_4443,N_5957);
or U6059 (N_6059,N_5305,N_4908);
nand U6060 (N_6060,N_5769,N_4184);
nor U6061 (N_6061,N_5732,N_5265);
nor U6062 (N_6062,N_4833,N_4925);
nand U6063 (N_6063,N_4494,N_5453);
xor U6064 (N_6064,N_4801,N_4259);
and U6065 (N_6065,N_4051,N_4628);
nand U6066 (N_6066,N_4935,N_4854);
nor U6067 (N_6067,N_4821,N_4419);
xor U6068 (N_6068,N_4464,N_5413);
nor U6069 (N_6069,N_4168,N_4912);
and U6070 (N_6070,N_5417,N_5232);
or U6071 (N_6071,N_4614,N_5020);
or U6072 (N_6072,N_4452,N_5435);
nor U6073 (N_6073,N_5429,N_5471);
or U6074 (N_6074,N_5269,N_5447);
or U6075 (N_6075,N_4946,N_5773);
nand U6076 (N_6076,N_4257,N_4579);
nor U6077 (N_6077,N_5856,N_4171);
or U6078 (N_6078,N_4949,N_5369);
and U6079 (N_6079,N_4982,N_5946);
or U6080 (N_6080,N_4740,N_4188);
nand U6081 (N_6081,N_5525,N_4165);
nor U6082 (N_6082,N_4822,N_4586);
or U6083 (N_6083,N_4708,N_4699);
and U6084 (N_6084,N_5433,N_4468);
or U6085 (N_6085,N_5353,N_4989);
nor U6086 (N_6086,N_5925,N_5785);
nor U6087 (N_6087,N_4971,N_4128);
and U6088 (N_6088,N_5162,N_4685);
nand U6089 (N_6089,N_4220,N_4047);
xnor U6090 (N_6090,N_5398,N_5120);
nand U6091 (N_6091,N_4093,N_5950);
or U6092 (N_6092,N_5700,N_4567);
nand U6093 (N_6093,N_4848,N_4885);
nand U6094 (N_6094,N_5289,N_5790);
and U6095 (N_6095,N_5175,N_5981);
xnor U6096 (N_6096,N_4601,N_5264);
nor U6097 (N_6097,N_5371,N_4944);
and U6098 (N_6098,N_4178,N_5543);
xor U6099 (N_6099,N_4245,N_4741);
xnor U6100 (N_6100,N_5430,N_4219);
and U6101 (N_6101,N_4700,N_5028);
nor U6102 (N_6102,N_5713,N_5951);
nand U6103 (N_6103,N_4438,N_4439);
or U6104 (N_6104,N_4123,N_5165);
xnor U6105 (N_6105,N_4045,N_5804);
nor U6106 (N_6106,N_5279,N_4910);
and U6107 (N_6107,N_4830,N_4250);
xor U6108 (N_6108,N_5064,N_5830);
and U6109 (N_6109,N_4482,N_4354);
or U6110 (N_6110,N_4046,N_4351);
nand U6111 (N_6111,N_4384,N_4672);
and U6112 (N_6112,N_5451,N_5899);
and U6113 (N_6113,N_4961,N_5597);
nor U6114 (N_6114,N_5665,N_5642);
or U6115 (N_6115,N_5296,N_4200);
and U6116 (N_6116,N_4585,N_4578);
and U6117 (N_6117,N_5933,N_5069);
and U6118 (N_6118,N_5404,N_5102);
and U6119 (N_6119,N_4266,N_4077);
nand U6120 (N_6120,N_5484,N_4066);
nor U6121 (N_6121,N_4998,N_4319);
or U6122 (N_6122,N_5152,N_4248);
nor U6123 (N_6123,N_4902,N_5067);
nand U6124 (N_6124,N_5277,N_5295);
nor U6125 (N_6125,N_5916,N_4959);
xnor U6126 (N_6126,N_5994,N_5478);
and U6127 (N_6127,N_4309,N_5647);
nor U6128 (N_6128,N_4226,N_4009);
or U6129 (N_6129,N_5229,N_5637);
or U6130 (N_6130,N_5600,N_4876);
nand U6131 (N_6131,N_5599,N_4790);
nand U6132 (N_6132,N_4268,N_5672);
nand U6133 (N_6133,N_4274,N_4518);
or U6134 (N_6134,N_5616,N_4573);
xor U6135 (N_6135,N_5325,N_4166);
nor U6136 (N_6136,N_5380,N_5179);
and U6137 (N_6137,N_5888,N_5847);
and U6138 (N_6138,N_4059,N_5057);
or U6139 (N_6139,N_4318,N_5418);
nand U6140 (N_6140,N_5657,N_4926);
and U6141 (N_6141,N_4788,N_4378);
nand U6142 (N_6142,N_4014,N_4777);
or U6143 (N_6143,N_4088,N_5897);
xnor U6144 (N_6144,N_4362,N_4356);
nor U6145 (N_6145,N_4284,N_5788);
or U6146 (N_6146,N_4209,N_5147);
nand U6147 (N_6147,N_4995,N_5898);
nor U6148 (N_6148,N_4979,N_5680);
nor U6149 (N_6149,N_4520,N_5740);
nand U6150 (N_6150,N_4510,N_5923);
and U6151 (N_6151,N_5387,N_4787);
nand U6152 (N_6152,N_4934,N_4393);
or U6153 (N_6153,N_4893,N_4224);
or U6154 (N_6154,N_4135,N_5195);
nand U6155 (N_6155,N_4426,N_4306);
or U6156 (N_6156,N_5343,N_4488);
nand U6157 (N_6157,N_5335,N_4582);
nand U6158 (N_6158,N_4064,N_4919);
nor U6159 (N_6159,N_5207,N_4921);
or U6160 (N_6160,N_5389,N_5623);
xnor U6161 (N_6161,N_5768,N_5215);
nand U6162 (N_6162,N_5718,N_4806);
or U6163 (N_6163,N_4634,N_5604);
and U6164 (N_6164,N_4721,N_5051);
and U6165 (N_6165,N_5357,N_5891);
xnor U6166 (N_6166,N_5942,N_5123);
and U6167 (N_6167,N_4726,N_4481);
and U6168 (N_6168,N_5907,N_5566);
xnor U6169 (N_6169,N_4210,N_5912);
xor U6170 (N_6170,N_4619,N_4418);
and U6171 (N_6171,N_5071,N_5583);
and U6172 (N_6172,N_5586,N_4339);
nor U6173 (N_6173,N_5301,N_5448);
nand U6174 (N_6174,N_5626,N_5693);
nor U6175 (N_6175,N_4540,N_4931);
xnor U6176 (N_6176,N_5314,N_4115);
nand U6177 (N_6177,N_5446,N_5712);
xnor U6178 (N_6178,N_5866,N_5405);
and U6179 (N_6179,N_4705,N_4538);
nand U6180 (N_6180,N_4841,N_5799);
xnor U6181 (N_6181,N_5745,N_5520);
or U6182 (N_6182,N_4845,N_4630);
or U6183 (N_6183,N_4031,N_4571);
nand U6184 (N_6184,N_5233,N_5294);
or U6185 (N_6185,N_4483,N_4665);
or U6186 (N_6186,N_4214,N_4564);
nand U6187 (N_6187,N_4015,N_4996);
or U6188 (N_6188,N_4953,N_5262);
nand U6189 (N_6189,N_4011,N_4013);
or U6190 (N_6190,N_5052,N_5258);
nand U6191 (N_6191,N_4645,N_5584);
nand U6192 (N_6192,N_4457,N_5144);
or U6193 (N_6193,N_5021,N_4541);
nor U6194 (N_6194,N_4253,N_4043);
and U6195 (N_6195,N_5169,N_5075);
nand U6196 (N_6196,N_4974,N_4793);
nand U6197 (N_6197,N_5991,N_5044);
or U6198 (N_6198,N_4892,N_5352);
nand U6199 (N_6199,N_5053,N_5153);
nand U6200 (N_6200,N_5652,N_4414);
nand U6201 (N_6201,N_4267,N_4666);
xnor U6202 (N_6202,N_4679,N_5337);
or U6203 (N_6203,N_5875,N_4975);
nor U6204 (N_6204,N_5460,N_4580);
nand U6205 (N_6205,N_5961,N_4742);
or U6206 (N_6206,N_5932,N_4235);
xnor U6207 (N_6207,N_5748,N_4558);
nand U6208 (N_6208,N_4560,N_5701);
or U6209 (N_6209,N_5884,N_4170);
xnor U6210 (N_6210,N_4904,N_4794);
and U6211 (N_6211,N_4528,N_4237);
nand U6212 (N_6212,N_5242,N_4888);
and U6213 (N_6213,N_4747,N_5031);
nand U6214 (N_6214,N_5761,N_5485);
or U6215 (N_6215,N_4475,N_4085);
or U6216 (N_6216,N_5872,N_5146);
nor U6217 (N_6217,N_5299,N_5834);
nand U6218 (N_6218,N_4198,N_4526);
and U6219 (N_6219,N_5971,N_5529);
nand U6220 (N_6220,N_4005,N_5434);
or U6221 (N_6221,N_5588,N_4207);
nor U6222 (N_6222,N_4978,N_4349);
nand U6223 (N_6223,N_4492,N_5585);
nand U6224 (N_6224,N_4316,N_5473);
nand U6225 (N_6225,N_5320,N_5037);
and U6226 (N_6226,N_4771,N_4361);
or U6227 (N_6227,N_4090,N_5011);
nor U6228 (N_6228,N_4081,N_5411);
nor U6229 (N_6229,N_4613,N_5579);
nand U6230 (N_6230,N_5070,N_5627);
and U6231 (N_6231,N_4435,N_5182);
and U6232 (N_6232,N_5166,N_4167);
and U6233 (N_6233,N_4503,N_4727);
nand U6234 (N_6234,N_4911,N_4856);
or U6235 (N_6235,N_5582,N_4938);
nor U6236 (N_6236,N_5820,N_4172);
and U6237 (N_6237,N_4029,N_5306);
nor U6238 (N_6238,N_5881,N_4325);
and U6239 (N_6239,N_5904,N_5648);
or U6240 (N_6240,N_4627,N_5730);
and U6241 (N_6241,N_4706,N_5241);
xor U6242 (N_6242,N_4555,N_5308);
and U6243 (N_6243,N_4999,N_5278);
or U6244 (N_6244,N_5641,N_4247);
nor U6245 (N_6245,N_4550,N_4052);
nand U6246 (N_6246,N_5318,N_5935);
nand U6247 (N_6247,N_4524,N_4766);
nand U6248 (N_6248,N_4142,N_4592);
or U6249 (N_6249,N_4772,N_5198);
nand U6250 (N_6250,N_5766,N_5456);
nor U6251 (N_6251,N_4690,N_4607);
nor U6252 (N_6252,N_5734,N_5244);
or U6253 (N_6253,N_4927,N_4420);
nor U6254 (N_6254,N_5876,N_5977);
and U6255 (N_6255,N_4866,N_4824);
or U6256 (N_6256,N_4695,N_5495);
or U6257 (N_6257,N_4263,N_4651);
and U6258 (N_6258,N_4322,N_4183);
nor U6259 (N_6259,N_5186,N_5705);
or U6260 (N_6260,N_4012,N_5344);
and U6261 (N_6261,N_4391,N_4341);
or U6262 (N_6262,N_4254,N_5594);
and U6263 (N_6263,N_5362,N_5338);
nor U6264 (N_6264,N_5423,N_4265);
nand U6265 (N_6265,N_4395,N_4301);
nand U6266 (N_6266,N_4374,N_4857);
and U6267 (N_6267,N_4738,N_5721);
and U6268 (N_6268,N_5844,N_5303);
and U6269 (N_6269,N_5088,N_5330);
nand U6270 (N_6270,N_5124,N_5470);
nand U6271 (N_6271,N_4661,N_5765);
or U6272 (N_6272,N_5363,N_5671);
or U6273 (N_6273,N_4466,N_4155);
nor U6274 (N_6274,N_4846,N_5459);
or U6275 (N_6275,N_4956,N_5287);
nor U6276 (N_6276,N_4376,N_5539);
nand U6277 (N_6277,N_4213,N_4299);
or U6278 (N_6278,N_4835,N_5170);
xnor U6279 (N_6279,N_4828,N_4024);
xor U6280 (N_6280,N_4662,N_5200);
or U6281 (N_6281,N_4387,N_5777);
and U6282 (N_6282,N_5086,N_5611);
or U6283 (N_6283,N_5098,N_5516);
nand U6284 (N_6284,N_4969,N_4137);
nor U6285 (N_6285,N_5465,N_5635);
and U6286 (N_6286,N_5860,N_5365);
or U6287 (N_6287,N_5677,N_4400);
nand U6288 (N_6288,N_4054,N_4517);
or U6289 (N_6289,N_4293,N_5668);
or U6290 (N_6290,N_4269,N_5838);
nor U6291 (N_6291,N_5770,N_4480);
or U6292 (N_6292,N_4421,N_5297);
or U6293 (N_6293,N_4298,N_5587);
nand U6294 (N_6294,N_5393,N_5613);
nand U6295 (N_6295,N_4035,N_4749);
or U6296 (N_6296,N_5673,N_5944);
nor U6297 (N_6297,N_5755,N_4616);
xor U6298 (N_6298,N_5240,N_4753);
and U6299 (N_6299,N_4026,N_4968);
nor U6300 (N_6300,N_5692,N_4057);
nand U6301 (N_6301,N_5131,N_5257);
and U6302 (N_6302,N_4144,N_5062);
nand U6303 (N_6303,N_5634,N_5578);
nor U6304 (N_6304,N_4369,N_4217);
xor U6305 (N_6305,N_4083,N_4175);
nand U6306 (N_6306,N_5729,N_4313);
and U6307 (N_6307,N_4062,N_5112);
xor U6308 (N_6308,N_4470,N_4108);
nor U6309 (N_6309,N_4383,N_5503);
nand U6310 (N_6310,N_4668,N_4260);
nor U6311 (N_6311,N_4739,N_5253);
or U6312 (N_6312,N_5840,N_4004);
or U6313 (N_6313,N_4120,N_4050);
nand U6314 (N_6314,N_5220,N_4448);
nand U6315 (N_6315,N_4321,N_4798);
xor U6316 (N_6316,N_5246,N_5742);
nand U6317 (N_6317,N_4344,N_4951);
nand U6318 (N_6318,N_5022,N_5480);
and U6319 (N_6319,N_5567,N_4397);
nor U6320 (N_6320,N_4962,N_5819);
and U6321 (N_6321,N_5367,N_4303);
nor U6322 (N_6322,N_4782,N_5203);
or U6323 (N_6323,N_5980,N_4689);
or U6324 (N_6324,N_4880,N_4649);
or U6325 (N_6325,N_5354,N_5833);
nand U6326 (N_6326,N_4352,N_5082);
nand U6327 (N_6327,N_4055,N_5893);
nor U6328 (N_6328,N_5445,N_5801);
and U6329 (N_6329,N_5800,N_4636);
nor U6330 (N_6330,N_4291,N_4889);
and U6331 (N_6331,N_4156,N_4089);
and U6332 (N_6332,N_5749,N_5895);
nor U6333 (N_6333,N_5327,N_4992);
nor U6334 (N_6334,N_5005,N_5171);
or U6335 (N_6335,N_4103,N_5025);
and U6336 (N_6336,N_4149,N_4006);
and U6337 (N_6337,N_4021,N_4851);
and U6338 (N_6338,N_5424,N_5225);
or U6339 (N_6339,N_5093,N_5115);
nor U6340 (N_6340,N_5592,N_4385);
and U6341 (N_6341,N_5682,N_4684);
nand U6342 (N_6342,N_4329,N_4240);
nand U6343 (N_6343,N_5822,N_4791);
xor U6344 (N_6344,N_4537,N_5015);
or U6345 (N_6345,N_5141,N_5999);
xnor U6346 (N_6346,N_5855,N_4724);
xnor U6347 (N_6347,N_4957,N_5212);
or U6348 (N_6348,N_4551,N_5276);
nor U6349 (N_6349,N_4599,N_5688);
nor U6350 (N_6350,N_4584,N_4826);
nor U6351 (N_6351,N_5651,N_4796);
and U6352 (N_6352,N_5211,N_4447);
nand U6353 (N_6353,N_5081,N_5395);
nand U6354 (N_6354,N_5328,N_5873);
nor U6355 (N_6355,N_5879,N_5072);
or U6356 (N_6356,N_5349,N_4789);
xor U6357 (N_6357,N_5645,N_5038);
nor U6358 (N_6358,N_4141,N_5666);
or U6359 (N_6359,N_4898,N_5181);
nor U6360 (N_6360,N_4288,N_5967);
and U6361 (N_6361,N_5210,N_5640);
nor U6362 (N_6362,N_5145,N_5826);
nor U6363 (N_6363,N_5576,N_5511);
nor U6364 (N_6364,N_5119,N_4729);
nor U6365 (N_6365,N_5990,N_5457);
nor U6366 (N_6366,N_5789,N_5127);
or U6367 (N_6367,N_5676,N_4531);
nand U6368 (N_6368,N_4922,N_5530);
xor U6369 (N_6369,N_5919,N_5662);
and U6370 (N_6370,N_5467,N_5821);
or U6371 (N_6371,N_5285,N_4228);
nor U6372 (N_6372,N_5234,N_5291);
nor U6373 (N_6373,N_4370,N_4413);
nand U6374 (N_6374,N_4988,N_4942);
nand U6375 (N_6375,N_5373,N_4417);
xnor U6376 (N_6376,N_4587,N_5963);
nor U6377 (N_6377,N_4745,N_4648);
and U6378 (N_6378,N_5184,N_5400);
nor U6379 (N_6379,N_4950,N_5964);
nor U6380 (N_6380,N_5235,N_4022);
nor U6381 (N_6381,N_4027,N_4850);
nor U6382 (N_6382,N_5483,N_4838);
or U6383 (N_6383,N_5047,N_4229);
or U6384 (N_6384,N_4489,N_4818);
and U6385 (N_6385,N_4302,N_5746);
and U6386 (N_6386,N_4078,N_4513);
nor U6387 (N_6387,N_4314,N_5591);
and U6388 (N_6388,N_5636,N_5118);
and U6389 (N_6389,N_4870,N_4122);
nor U6390 (N_6390,N_4191,N_4915);
and U6391 (N_6391,N_4852,N_4652);
nand U6392 (N_6392,N_4121,N_4715);
and U6393 (N_6393,N_5440,N_4450);
or U6394 (N_6394,N_5625,N_5807);
xor U6395 (N_6395,N_5508,N_4675);
or U6396 (N_6396,N_4307,N_4458);
xnor U6397 (N_6397,N_5399,N_4602);
or U6398 (N_6398,N_4206,N_4686);
nand U6399 (N_6399,N_4203,N_4251);
and U6400 (N_6400,N_4823,N_5073);
or U6401 (N_6401,N_5218,N_4423);
nor U6402 (N_6402,N_5596,N_4776);
nor U6403 (N_6403,N_5368,N_5331);
xor U6404 (N_6404,N_4688,N_5784);
or U6405 (N_6405,N_5173,N_5199);
nand U6406 (N_6406,N_4283,N_5042);
or U6407 (N_6407,N_5035,N_5571);
nand U6408 (N_6408,N_5281,N_4767);
nand U6409 (N_6409,N_4473,N_5723);
or U6410 (N_6410,N_5908,N_4546);
xor U6411 (N_6411,N_4635,N_5943);
and U6412 (N_6412,N_4811,N_4491);
xor U6413 (N_6413,N_5886,N_4954);
and U6414 (N_6414,N_4591,N_4199);
and U6415 (N_6415,N_5489,N_4664);
nand U6416 (N_6416,N_5007,N_4201);
xor U6417 (N_6417,N_5778,N_4404);
and U6418 (N_6418,N_5346,N_4367);
nand U6419 (N_6419,N_4569,N_5926);
nand U6420 (N_6420,N_5966,N_5030);
or U6421 (N_6421,N_5581,N_4696);
nand U6422 (N_6422,N_4594,N_5139);
nor U6423 (N_6423,N_4941,N_5915);
or U6424 (N_6424,N_5969,N_5914);
and U6425 (N_6425,N_4807,N_5556);
xor U6426 (N_6426,N_4280,N_5206);
or U6427 (N_6427,N_4487,N_4246);
and U6428 (N_6428,N_5224,N_5928);
xnor U6429 (N_6429,N_5477,N_4348);
and U6430 (N_6430,N_5420,N_5189);
nor U6431 (N_6431,N_5412,N_5827);
nor U6432 (N_6432,N_5796,N_4028);
or U6433 (N_6433,N_5975,N_4381);
nor U6434 (N_6434,N_5386,N_4812);
nor U6435 (N_6435,N_5707,N_4757);
or U6436 (N_6436,N_4337,N_4112);
nor U6437 (N_6437,N_5602,N_5458);
nand U6438 (N_6438,N_5568,N_5217);
nor U6439 (N_6439,N_5402,N_5310);
xor U6440 (N_6440,N_4105,N_5687);
or U6441 (N_6441,N_4612,N_5226);
nor U6442 (N_6442,N_4087,N_4408);
and U6443 (N_6443,N_5383,N_4674);
and U6444 (N_6444,N_5290,N_5948);
nor U6445 (N_6445,N_5557,N_4252);
nor U6446 (N_6446,N_4836,N_4132);
nor U6447 (N_6447,N_5910,N_5762);
nand U6448 (N_6448,N_5462,N_4667);
nand U6449 (N_6449,N_5690,N_5128);
nand U6450 (N_6450,N_4151,N_5077);
xor U6451 (N_6451,N_5621,N_5720);
nor U6452 (N_6452,N_4446,N_5129);
and U6453 (N_6453,N_5786,N_5547);
nand U6454 (N_6454,N_4543,N_5922);
xnor U6455 (N_6455,N_4765,N_5580);
or U6456 (N_6456,N_4924,N_4825);
or U6457 (N_6457,N_5650,N_5095);
nand U6458 (N_6458,N_4804,N_5810);
nand U6459 (N_6459,N_4676,N_4991);
and U6460 (N_6460,N_5744,N_5837);
nor U6461 (N_6461,N_5227,N_5302);
or U6462 (N_6462,N_5027,N_4311);
and U6463 (N_6463,N_4478,N_5094);
xnor U6464 (N_6464,N_5286,N_5248);
nor U6465 (N_6465,N_5832,N_4879);
or U6466 (N_6466,N_5995,N_4671);
and U6467 (N_6467,N_5313,N_5300);
and U6468 (N_6468,N_4744,N_5083);
nor U6469 (N_6469,N_4901,N_5900);
nor U6470 (N_6470,N_5315,N_5573);
nand U6471 (N_6471,N_4444,N_5917);
nor U6472 (N_6472,N_4877,N_5178);
and U6473 (N_6473,N_5708,N_4815);
or U6474 (N_6474,N_5505,N_5521);
or U6475 (N_6475,N_5103,N_5336);
nor U6476 (N_6476,N_5487,N_4565);
or U6477 (N_6477,N_4764,N_5012);
nor U6478 (N_6478,N_5033,N_4272);
and U6479 (N_6479,N_5703,N_5298);
and U6480 (N_6480,N_5040,N_4440);
and U6481 (N_6481,N_5614,N_4113);
nand U6482 (N_6482,N_5979,N_5245);
and U6483 (N_6483,N_5089,N_5507);
nor U6484 (N_6484,N_4844,N_4347);
nor U6485 (N_6485,N_4179,N_5415);
nor U6486 (N_6486,N_4784,N_4186);
or U6487 (N_6487,N_4597,N_4958);
or U6488 (N_6488,N_5871,N_4521);
or U6489 (N_6489,N_5601,N_5795);
nand U6490 (N_6490,N_5542,N_4294);
nand U6491 (N_6491,N_5063,N_5846);
or U6492 (N_6492,N_5499,N_4003);
or U6493 (N_6493,N_4755,N_4032);
nand U6494 (N_6494,N_5527,N_4097);
and U6495 (N_6495,N_4802,N_4118);
and U6496 (N_6496,N_4020,N_5835);
or U6497 (N_6497,N_5486,N_5345);
or U6498 (N_6498,N_4986,N_4146);
nor U6499 (N_6499,N_4681,N_5554);
and U6500 (N_6500,N_4557,N_4262);
nand U6501 (N_6501,N_5076,N_4164);
and U6502 (N_6502,N_4909,N_5222);
nor U6503 (N_6503,N_5767,N_5538);
or U6504 (N_6504,N_4669,N_5552);
or U6505 (N_6505,N_4913,N_5660);
and U6506 (N_6506,N_5437,N_4377);
nand U6507 (N_6507,N_4799,N_4936);
or U6508 (N_6508,N_4270,N_5097);
nand U6509 (N_6509,N_5174,N_4637);
nand U6510 (N_6510,N_5441,N_4598);
nor U6511 (N_6511,N_5324,N_5883);
and U6512 (N_6512,N_5205,N_4677);
and U6513 (N_6513,N_4983,N_4223);
and U6514 (N_6514,N_4750,N_5983);
or U6515 (N_6515,N_4500,N_4434);
xor U6516 (N_6516,N_5779,N_4428);
or U6517 (N_6517,N_4278,N_4553);
nand U6518 (N_6518,N_5741,N_4816);
nand U6519 (N_6519,N_5284,N_5250);
xor U6520 (N_6520,N_4454,N_4873);
or U6521 (N_6521,N_4963,N_5513);
nand U6522 (N_6522,N_4350,N_4145);
nand U6523 (N_6523,N_4819,N_4548);
xnor U6524 (N_6524,N_5461,N_4887);
nand U6525 (N_6525,N_4697,N_5230);
and U6526 (N_6526,N_5754,N_5523);
nor U6527 (N_6527,N_5317,N_5612);
nor U6528 (N_6528,N_4190,N_5187);
nand U6529 (N_6529,N_4914,N_5940);
nand U6530 (N_6530,N_4394,N_5329);
nand U6531 (N_6531,N_4778,N_5661);
nand U6532 (N_6532,N_4104,N_5180);
xnor U6533 (N_6533,N_5023,N_5100);
nor U6534 (N_6534,N_5428,N_5726);
nand U6535 (N_6535,N_5709,N_4687);
nor U6536 (N_6536,N_5985,N_5564);
xor U6537 (N_6537,N_4281,N_5061);
or U6538 (N_6538,N_4642,N_5024);
nand U6539 (N_6539,N_4416,N_5263);
nand U6540 (N_6540,N_5501,N_4053);
and U6541 (N_6541,N_4831,N_4952);
or U6542 (N_6542,N_5493,N_5105);
and U6543 (N_6543,N_5679,N_5378);
nor U6544 (N_6544,N_5890,N_5464);
nor U6545 (N_6545,N_4019,N_5196);
xnor U6546 (N_6546,N_4539,N_4320);
nand U6547 (N_6547,N_5494,N_4977);
xor U6548 (N_6548,N_4182,N_4490);
nor U6549 (N_6549,N_5439,N_4894);
nand U6550 (N_6550,N_4710,N_5845);
and U6551 (N_6551,N_4930,N_4346);
nor U6552 (N_6552,N_4264,N_4530);
nand U6553 (N_6553,N_5359,N_5273);
nand U6554 (N_6554,N_4746,N_5603);
or U6555 (N_6555,N_4709,N_4572);
nand U6556 (N_6556,N_4016,N_5332);
nand U6557 (N_6557,N_4570,N_4754);
nand U6558 (N_6558,N_4343,N_4632);
and U6559 (N_6559,N_5517,N_5252);
nor U6560 (N_6560,N_5074,N_5512);
nor U6561 (N_6561,N_4160,N_5553);
nor U6562 (N_6562,N_4752,N_5750);
nand U6563 (N_6563,N_5361,N_5984);
nand U6564 (N_6564,N_4920,N_4355);
nand U6565 (N_6565,N_4633,N_4863);
nand U6566 (N_6566,N_5731,N_4069);
and U6567 (N_6567,N_4086,N_4918);
or U6568 (N_6568,N_5569,N_4897);
and U6569 (N_6569,N_4463,N_4624);
nor U6570 (N_6570,N_4159,N_5854);
xor U6571 (N_6571,N_5443,N_4379);
and U6572 (N_6572,N_4865,N_4304);
and U6573 (N_6573,N_4758,N_5060);
or U6574 (N_6574,N_5292,N_4133);
xnor U6575 (N_6575,N_5880,N_4717);
nor U6576 (N_6576,N_4670,N_5001);
nor U6577 (N_6577,N_5758,N_4785);
nand U6578 (N_6578,N_5432,N_4574);
nor U6579 (N_6579,N_5436,N_4084);
nor U6580 (N_6580,N_5048,N_4683);
or U6581 (N_6581,N_4639,N_4472);
or U6582 (N_6582,N_5998,N_4884);
or U6583 (N_6583,N_5939,N_4832);
or U6584 (N_6584,N_5805,N_5558);
or U6585 (N_6585,N_4363,N_4868);
and U6586 (N_6586,N_5813,N_4241);
xnor U6587 (N_6587,N_4427,N_5125);
or U6588 (N_6588,N_4000,N_4609);
xnor U6589 (N_6589,N_4625,N_4119);
nand U6590 (N_6590,N_4008,N_4732);
xnor U6591 (N_6591,N_5255,N_5638);
or U6592 (N_6592,N_5510,N_4534);
xnor U6593 (N_6593,N_4474,N_4092);
nor U6594 (N_6594,N_4631,N_4803);
nand U6595 (N_6595,N_4401,N_4353);
and U6596 (N_6596,N_4402,N_5649);
and U6597 (N_6597,N_4469,N_5113);
xnor U6598 (N_6598,N_5046,N_4720);
and U6599 (N_6599,N_4929,N_5733);
and U6600 (N_6600,N_5163,N_4817);
nand U6601 (N_6601,N_5231,N_5811);
nor U6602 (N_6602,N_5717,N_4258);
nor U6603 (N_6603,N_4716,N_5575);
nand U6604 (N_6604,N_5168,N_5955);
nor U6605 (N_6605,N_4124,N_5533);
xnor U6606 (N_6606,N_4554,N_5619);
nand U6607 (N_6607,N_5885,N_5970);
or U6608 (N_6608,N_4079,N_4981);
and U6609 (N_6609,N_4437,N_4869);
and U6610 (N_6610,N_5803,N_5137);
xor U6611 (N_6611,N_4324,N_5670);
nor U6612 (N_6612,N_4073,N_5376);
nor U6613 (N_6613,N_4127,N_4001);
or U6614 (N_6614,N_4508,N_4762);
or U6615 (N_6615,N_5823,N_4275);
and U6616 (N_6616,N_4875,N_4581);
nand U6617 (N_6617,N_5947,N_4076);
xnor U6618 (N_6618,N_4878,N_4152);
nand U6619 (N_6619,N_4196,N_5476);
and U6620 (N_6620,N_4357,N_5379);
and U6621 (N_6621,N_4140,N_4820);
and U6622 (N_6622,N_4082,N_4556);
nor U6623 (N_6623,N_5738,N_5524);
and U6624 (N_6624,N_5781,N_5039);
and U6625 (N_6625,N_4493,N_4660);
nor U6626 (N_6626,N_4038,N_4154);
and U6627 (N_6627,N_5696,N_4218);
and U6628 (N_6628,N_4358,N_4449);
nor U6629 (N_6629,N_4970,N_5534);
nand U6630 (N_6630,N_5236,N_4590);
nand U6631 (N_6631,N_4973,N_5954);
and U6632 (N_6632,N_5059,N_5117);
nand U6633 (N_6633,N_4036,N_4018);
xor U6634 (N_6634,N_4126,N_4023);
xnor U6635 (N_6635,N_5216,N_4568);
and U6636 (N_6636,N_5410,N_4947);
xor U6637 (N_6637,N_5535,N_4774);
and U6638 (N_6638,N_4972,N_5719);
nand U6639 (N_6639,N_4380,N_5202);
or U6640 (N_6640,N_5536,N_5056);
nor U6641 (N_6641,N_4456,N_5808);
and U6642 (N_6642,N_4663,N_5909);
xor U6643 (N_6643,N_5348,N_5249);
nand U6644 (N_6644,N_5710,N_4596);
nor U6645 (N_6645,N_4317,N_5058);
xnor U6646 (N_6646,N_4331,N_5794);
nor U6647 (N_6647,N_4808,N_5938);
and U6648 (N_6648,N_5358,N_4737);
xor U6649 (N_6649,N_4542,N_4010);
nor U6650 (N_6650,N_5722,N_5757);
nor U6651 (N_6651,N_5316,N_5798);
or U6652 (N_6652,N_4626,N_5859);
and U6653 (N_6653,N_4563,N_4405);
and U6654 (N_6654,N_5669,N_5191);
nand U6655 (N_6655,N_4163,N_5172);
or U6656 (N_6656,N_5605,N_5572);
nor U6657 (N_6657,N_4837,N_4338);
or U6658 (N_6658,N_4611,N_5004);
and U6659 (N_6659,N_5711,N_5450);
and U6660 (N_6660,N_4514,N_5403);
and U6661 (N_6661,N_4056,N_4327);
or U6662 (N_6662,N_4945,N_4748);
nor U6663 (N_6663,N_5628,N_4527);
and U6664 (N_6664,N_5667,N_5725);
nand U6665 (N_6665,N_5492,N_4916);
and U6666 (N_6666,N_4205,N_4496);
nand U6667 (N_6667,N_5282,N_4192);
or U6668 (N_6668,N_4230,N_4116);
xnor U6669 (N_6669,N_5853,N_4484);
or U6670 (N_6670,N_4432,N_5685);
and U6671 (N_6671,N_5992,N_5454);
or U6672 (N_6672,N_5797,N_5982);
or U6673 (N_6673,N_5084,N_5824);
or U6674 (N_6674,N_4360,N_4276);
nand U6675 (N_6675,N_4098,N_4583);
xnor U6676 (N_6676,N_5394,N_4621);
nand U6677 (N_6677,N_4905,N_4048);
nand U6678 (N_6678,N_4091,N_5197);
or U6679 (N_6679,N_4208,N_4903);
nor U6680 (N_6680,N_4234,N_4858);
nand U6681 (N_6681,N_5903,N_5130);
nor U6682 (N_6682,N_5392,N_4734);
or U6683 (N_6683,N_4177,N_4204);
nand U6684 (N_6684,N_4693,N_4588);
nand U6685 (N_6685,N_5201,N_5356);
nand U6686 (N_6686,N_4532,N_4273);
xor U6687 (N_6687,N_5268,N_5468);
and U6688 (N_6688,N_5514,N_4017);
xor U6689 (N_6689,N_4595,N_5351);
and U6690 (N_6690,N_5825,N_5929);
or U6691 (N_6691,N_4392,N_4511);
nand U6692 (N_6692,N_4600,N_5018);
xnor U6693 (N_6693,N_4861,N_5630);
nand U6694 (N_6694,N_5270,N_4512);
and U6695 (N_6695,N_5675,N_5691);
or U6696 (N_6696,N_4604,N_4827);
and U6697 (N_6697,N_5016,N_5391);
and U6698 (N_6698,N_4412,N_4340);
or U6699 (N_6699,N_4336,N_4364);
nor U6700 (N_6700,N_5193,N_4326);
nand U6701 (N_6701,N_5664,N_4173);
or U6702 (N_6702,N_5996,N_5851);
and U6703 (N_6703,N_5322,N_4650);
nor U6704 (N_6704,N_5122,N_4638);
and U6705 (N_6705,N_5952,N_5997);
or U6706 (N_6706,N_4723,N_4037);
and U6707 (N_6707,N_5877,N_5643);
nand U6708 (N_6708,N_4328,N_4030);
and U6709 (N_6709,N_4509,N_5079);
or U6710 (N_6710,N_5760,N_5455);
nand U6711 (N_6711,N_5772,N_5340);
nand U6712 (N_6712,N_5659,N_5663);
nor U6713 (N_6713,N_5973,N_4107);
nor U6714 (N_6714,N_5550,N_4522);
nand U6715 (N_6715,N_5841,N_5409);
nor U6716 (N_6716,N_5319,N_5541);
xor U6717 (N_6717,N_4150,N_5989);
and U6718 (N_6718,N_5228,N_5653);
or U6719 (N_6719,N_4158,N_4654);
xor U6720 (N_6720,N_4535,N_5096);
and U6721 (N_6721,N_4606,N_4244);
and U6722 (N_6722,N_4780,N_5190);
or U6723 (N_6723,N_5256,N_5549);
and U6724 (N_6724,N_5160,N_4781);
and U6725 (N_6725,N_4853,N_5157);
and U6726 (N_6726,N_5401,N_5366);
nand U6727 (N_6727,N_5561,N_5960);
and U6728 (N_6728,N_5333,N_5452);
or U6729 (N_6729,N_5006,N_4834);
nand U6730 (N_6730,N_4422,N_4775);
or U6731 (N_6731,N_5043,N_5384);
nor U6732 (N_6732,N_5150,N_5901);
and U6733 (N_6733,N_5406,N_4389);
nor U6734 (N_6734,N_5715,N_5479);
and U6735 (N_6735,N_5334,N_4025);
nor U6736 (N_6736,N_5140,N_4044);
xor U6737 (N_6737,N_4442,N_5188);
nand U6738 (N_6738,N_4967,N_4286);
nand U6739 (N_6739,N_4608,N_5111);
xor U6740 (N_6740,N_4215,N_4197);
nand U6741 (N_6741,N_4719,N_5828);
nand U6742 (N_6742,N_4965,N_5809);
nor U6743 (N_6743,N_5956,N_5463);
and U6744 (N_6744,N_5272,N_5655);
xnor U6745 (N_6745,N_4620,N_4809);
xnor U6746 (N_6746,N_4498,N_5629);
nand U6747 (N_6747,N_4536,N_5632);
or U6748 (N_6748,N_5090,N_4305);
nor U6749 (N_6749,N_4779,N_5055);
xor U6750 (N_6750,N_5091,N_5154);
nor U6751 (N_6751,N_4388,N_4864);
nand U6752 (N_6752,N_5782,N_5099);
and U6753 (N_6753,N_5372,N_5589);
and U6754 (N_6754,N_5593,N_4939);
nor U6755 (N_6755,N_4692,N_5142);
nor U6756 (N_6756,N_4227,N_5868);
nor U6757 (N_6757,N_5350,N_5686);
or U6758 (N_6758,N_4425,N_4399);
nor U6759 (N_6759,N_5831,N_5774);
nor U6760 (N_6760,N_4101,N_4768);
nand U6761 (N_6761,N_4680,N_4733);
or U6762 (N_6762,N_4505,N_4212);
and U6763 (N_6763,N_5624,N_4169);
or U6764 (N_6764,N_4396,N_5490);
and U6765 (N_6765,N_5014,N_4060);
xor U6766 (N_6766,N_5563,N_5953);
and U6767 (N_6767,N_4703,N_5607);
and U6768 (N_6768,N_4249,N_4415);
nand U6769 (N_6769,N_5274,N_5017);
xor U6770 (N_6770,N_5848,N_4211);
nor U6771 (N_6771,N_5958,N_5254);
and U6772 (N_6772,N_5008,N_5577);
and U6773 (N_6773,N_5370,N_5815);
nand U6774 (N_6774,N_5595,N_5321);
or U6775 (N_6775,N_5419,N_4430);
or U6776 (N_6776,N_4862,N_5381);
and U6777 (N_6777,N_4277,N_5878);
nand U6778 (N_6778,N_5756,N_4618);
or U6779 (N_6779,N_5987,N_5502);
and U6780 (N_6780,N_4643,N_4948);
nor U6781 (N_6781,N_5889,N_4403);
and U6782 (N_6782,N_4722,N_4761);
nand U6783 (N_6783,N_4499,N_5959);
xnor U6784 (N_6784,N_5874,N_5482);
and U6785 (N_6785,N_4533,N_5598);
xor U6786 (N_6786,N_4153,N_4342);
nor U6787 (N_6787,N_4424,N_4411);
xor U6788 (N_6788,N_5271,N_4736);
nand U6789 (N_6789,N_5737,N_5654);
and U6790 (N_6790,N_5633,N_4130);
nor U6791 (N_6791,N_5237,N_4507);
nand U6792 (N_6792,N_4398,N_5126);
nor U6793 (N_6793,N_5610,N_5293);
nand U6794 (N_6794,N_5850,N_4180);
nand U6795 (N_6795,N_5364,N_4646);
nand U6796 (N_6796,N_5026,N_5780);
nor U6797 (N_6797,N_5209,N_5045);
and U6798 (N_6798,N_5702,N_5689);
or U6799 (N_6799,N_5618,N_4332);
nor U6800 (N_6800,N_5962,N_4980);
and U6801 (N_6801,N_4042,N_5159);
and U6802 (N_6802,N_5858,N_4061);
nand U6803 (N_6803,N_4994,N_5239);
or U6804 (N_6804,N_4195,N_5728);
nand U6805 (N_6805,N_4955,N_5802);
nand U6806 (N_6806,N_4187,N_5739);
nand U6807 (N_6807,N_4068,N_5751);
xor U6808 (N_6808,N_5339,N_5132);
nand U6809 (N_6809,N_5390,N_5176);
nor U6810 (N_6810,N_5416,N_5283);
and U6811 (N_6811,N_5764,N_4406);
nor U6812 (N_6812,N_5425,N_5243);
and U6813 (N_6813,N_5148,N_4471);
nand U6814 (N_6814,N_4529,N_4368);
and U6815 (N_6815,N_4371,N_5545);
and U6816 (N_6816,N_5002,N_5656);
or U6817 (N_6817,N_4519,N_5972);
nor U6818 (N_6818,N_5275,N_5724);
or U6819 (N_6819,N_5763,N_4109);
xor U6820 (N_6820,N_4525,N_4842);
and U6821 (N_6821,N_4477,N_4174);
nand U6822 (N_6822,N_4725,N_4966);
nor U6823 (N_6823,N_4323,N_5407);
or U6824 (N_6824,N_5397,N_5442);
nor U6825 (N_6825,N_5526,N_5375);
or U6826 (N_6826,N_5546,N_4138);
and U6827 (N_6827,N_4810,N_4502);
nand U6828 (N_6828,N_5161,N_4382);
and U6829 (N_6829,N_5155,N_5683);
nand U6830 (N_6830,N_4847,N_4882);
xnor U6831 (N_6831,N_4289,N_4872);
xor U6832 (N_6832,N_5498,N_5408);
and U6833 (N_6833,N_5092,N_5522);
or U6834 (N_6834,N_4034,N_5783);
nor U6835 (N_6835,N_4111,N_4698);
nor U6836 (N_6836,N_4743,N_5506);
nor U6837 (N_6837,N_5622,N_5134);
nand U6838 (N_6838,N_4139,N_5158);
and U6839 (N_6839,N_4756,N_5156);
nand U6840 (N_6840,N_4007,N_5787);
nand U6841 (N_6841,N_4829,N_5078);
and U6842 (N_6842,N_5678,N_5968);
and U6843 (N_6843,N_4134,N_4763);
nor U6844 (N_6844,N_4233,N_5727);
or U6845 (N_6845,N_5219,N_4792);
nand U6846 (N_6846,N_4049,N_4504);
nor U6847 (N_6847,N_4162,N_4074);
or U6848 (N_6848,N_4840,N_5342);
nor U6849 (N_6849,N_5759,N_4102);
nor U6850 (N_6850,N_5177,N_4906);
and U6851 (N_6851,N_5869,N_4751);
or U6852 (N_6852,N_4315,N_5565);
or U6853 (N_6853,N_5863,N_5839);
or U6854 (N_6854,N_5396,N_5167);
or U6855 (N_6855,N_4658,N_5138);
nand U6856 (N_6856,N_4441,N_5931);
nor U6857 (N_6857,N_5698,N_4067);
nor U6858 (N_6858,N_5620,N_4682);
nor U6859 (N_6859,N_4896,N_5000);
or U6860 (N_6860,N_4390,N_5449);
nand U6861 (N_6861,N_4075,N_5531);
nor U6862 (N_6862,N_5326,N_4545);
or U6863 (N_6863,N_5347,N_5497);
and U6864 (N_6864,N_4559,N_4640);
nor U6865 (N_6865,N_5852,N_5185);
nor U6866 (N_6866,N_4255,N_5068);
nor U6867 (N_6867,N_4345,N_4932);
or U6868 (N_6868,N_4577,N_4786);
nor U6869 (N_6869,N_4937,N_5029);
and U6870 (N_6870,N_5528,N_5864);
nor U6871 (N_6871,N_4561,N_5816);
nand U6872 (N_6872,N_5551,N_5032);
nand U6873 (N_6873,N_5775,N_5631);
or U6874 (N_6874,N_4795,N_4928);
or U6875 (N_6875,N_5013,N_4287);
nand U6876 (N_6876,N_4445,N_5882);
and U6877 (N_6877,N_4704,N_5681);
or U6878 (N_6878,N_4148,N_4292);
or U6879 (N_6879,N_4453,N_5087);
nand U6880 (N_6880,N_4333,N_5791);
nand U6881 (N_6881,N_4479,N_5559);
nand U6882 (N_6882,N_4256,N_4805);
nand U6883 (N_6883,N_4874,N_4099);
and U6884 (N_6884,N_5934,N_4239);
nand U6885 (N_6885,N_4523,N_5192);
and U6886 (N_6886,N_4855,N_5736);
or U6887 (N_6887,N_4300,N_5247);
xnor U6888 (N_6888,N_5548,N_5496);
or U6889 (N_6889,N_4849,N_5309);
nand U6890 (N_6890,N_5164,N_4544);
or U6891 (N_6891,N_4515,N_4242);
nand U6892 (N_6892,N_5085,N_4261);
and U6893 (N_6893,N_5704,N_5949);
or U6894 (N_6894,N_5221,N_5472);
nand U6895 (N_6895,N_4310,N_4386);
nand U6896 (N_6896,N_5887,N_5054);
or U6897 (N_6897,N_5537,N_5469);
and U6898 (N_6898,N_5694,N_4497);
or U6899 (N_6899,N_4359,N_4647);
and U6900 (N_6900,N_4655,N_4295);
xnor U6901 (N_6901,N_5050,N_5108);
or U6902 (N_6902,N_4485,N_4161);
nand U6903 (N_6903,N_5986,N_5993);
xor U6904 (N_6904,N_5936,N_4238);
and U6905 (N_6905,N_4783,N_5518);
nand U6906 (N_6906,N_5924,N_4189);
nor U6907 (N_6907,N_5360,N_5945);
and U6908 (N_6908,N_5927,N_4096);
nor U6909 (N_6909,N_5776,N_4117);
nand U6910 (N_6910,N_5385,N_5066);
or U6911 (N_6911,N_5019,N_4800);
or U6912 (N_6912,N_4899,N_4702);
nand U6913 (N_6913,N_5792,N_4907);
and U6914 (N_6914,N_4735,N_4984);
nand U6915 (N_6915,N_4366,N_4002);
nor U6916 (N_6916,N_5818,N_5562);
nand U6917 (N_6917,N_5555,N_4222);
nand U6918 (N_6918,N_4718,N_4673);
and U6919 (N_6919,N_4923,N_5288);
or U6920 (N_6920,N_4714,N_5475);
and U6921 (N_6921,N_4843,N_5913);
nor U6922 (N_6922,N_5106,N_4467);
nor U6923 (N_6923,N_5110,N_5697);
or U6924 (N_6924,N_5695,N_5609);
nand U6925 (N_6925,N_4143,N_4431);
nand U6926 (N_6926,N_5466,N_5930);
or U6927 (N_6927,N_5857,N_4940);
or U6928 (N_6928,N_5920,N_5010);
nor U6929 (N_6929,N_5009,N_5806);
and U6930 (N_6930,N_5280,N_5519);
and U6931 (N_6931,N_4615,N_5311);
xor U6932 (N_6932,N_5377,N_4993);
and U6933 (N_6933,N_5658,N_5937);
nand U6934 (N_6934,N_4694,N_4985);
nor U6935 (N_6935,N_4593,N_4617);
and U6936 (N_6936,N_4813,N_4202);
xor U6937 (N_6937,N_5849,N_5133);
nor U6938 (N_6938,N_4707,N_4476);
nand U6939 (N_6939,N_4501,N_5735);
nor U6940 (N_6940,N_5865,N_5911);
nand U6941 (N_6941,N_5902,N_4797);
nand U6942 (N_6942,N_5842,N_4110);
nor U6943 (N_6943,N_5491,N_4131);
nor U6944 (N_6944,N_5574,N_4701);
nand U6945 (N_6945,N_5706,N_5238);
and U6946 (N_6946,N_5817,N_5570);
or U6947 (N_6947,N_4589,N_5515);
and U6948 (N_6948,N_4495,N_4070);
and U6949 (N_6949,N_4770,N_5251);
nor U6950 (N_6950,N_5892,N_5194);
or U6951 (N_6951,N_5540,N_4279);
or U6952 (N_6952,N_4883,N_5814);
and U6953 (N_6953,N_5431,N_5714);
xor U6954 (N_6954,N_5743,N_4065);
nand U6955 (N_6955,N_5747,N_5965);
nand U6956 (N_6956,N_5870,N_5382);
and U6957 (N_6957,N_4773,N_4451);
and U6958 (N_6958,N_4506,N_4605);
nor U6959 (N_6959,N_4459,N_4943);
nand U6960 (N_6960,N_5862,N_5906);
nor U6961 (N_6961,N_4960,N_4867);
and U6962 (N_6962,N_4656,N_5421);
nand U6963 (N_6963,N_5974,N_4465);
or U6964 (N_6964,N_5183,N_5752);
and U6965 (N_6965,N_4461,N_4871);
or U6966 (N_6966,N_5861,N_4711);
or U6967 (N_6967,N_5041,N_4886);
nand U6968 (N_6968,N_4236,N_5716);
or U6969 (N_6969,N_4334,N_4712);
nand U6970 (N_6970,N_5905,N_5101);
xnor U6971 (N_6971,N_4365,N_4033);
xor U6972 (N_6972,N_4181,N_5223);
and U6973 (N_6973,N_5843,N_5312);
and U6974 (N_6974,N_5532,N_4221);
or U6975 (N_6975,N_5107,N_5941);
or U6976 (N_6976,N_4881,N_5812);
xnor U6977 (N_6977,N_5921,N_5136);
and U6978 (N_6978,N_5080,N_5988);
and U6979 (N_6979,N_5214,N_4516);
and U6980 (N_6980,N_4335,N_4814);
or U6981 (N_6981,N_4691,N_5444);
and U6982 (N_6982,N_4330,N_4231);
nand U6983 (N_6983,N_5065,N_5500);
nand U6984 (N_6984,N_5109,N_4106);
xnor U6985 (N_6985,N_4860,N_4232);
nor U6986 (N_6986,N_4455,N_4290);
xor U6987 (N_6987,N_5504,N_4072);
nor U6988 (N_6988,N_5615,N_5034);
or U6989 (N_6989,N_5829,N_4429);
or U6990 (N_6990,N_4562,N_4185);
and U6991 (N_6991,N_4063,N_4193);
or U6992 (N_6992,N_4644,N_4839);
xor U6993 (N_6993,N_4575,N_5793);
xor U6994 (N_6994,N_4080,N_4900);
nor U6995 (N_6995,N_4094,N_4407);
nand U6996 (N_6996,N_5149,N_4157);
nand U6997 (N_6997,N_4622,N_4552);
or U6998 (N_6998,N_4895,N_5266);
nand U6999 (N_6999,N_4058,N_5474);
and U7000 (N_7000,N_5175,N_4134);
xor U7001 (N_7001,N_4814,N_4974);
nor U7002 (N_7002,N_4715,N_5560);
and U7003 (N_7003,N_5656,N_4688);
nor U7004 (N_7004,N_4450,N_5210);
and U7005 (N_7005,N_5884,N_5412);
xnor U7006 (N_7006,N_4821,N_5918);
and U7007 (N_7007,N_4787,N_4030);
nand U7008 (N_7008,N_5384,N_4902);
and U7009 (N_7009,N_4376,N_4126);
or U7010 (N_7010,N_4300,N_5934);
or U7011 (N_7011,N_4091,N_5882);
nand U7012 (N_7012,N_5167,N_4861);
nor U7013 (N_7013,N_5564,N_5688);
and U7014 (N_7014,N_4440,N_4286);
nand U7015 (N_7015,N_5901,N_5869);
and U7016 (N_7016,N_4208,N_5275);
nor U7017 (N_7017,N_5631,N_5366);
nor U7018 (N_7018,N_4673,N_4560);
nand U7019 (N_7019,N_4552,N_5382);
and U7020 (N_7020,N_4743,N_4872);
and U7021 (N_7021,N_4259,N_5959);
and U7022 (N_7022,N_4741,N_4266);
or U7023 (N_7023,N_4321,N_4033);
and U7024 (N_7024,N_4701,N_4619);
nand U7025 (N_7025,N_5392,N_4244);
or U7026 (N_7026,N_4026,N_5780);
nor U7027 (N_7027,N_5352,N_5949);
and U7028 (N_7028,N_4600,N_5811);
nand U7029 (N_7029,N_4920,N_4470);
nor U7030 (N_7030,N_4809,N_5809);
and U7031 (N_7031,N_5686,N_4081);
nor U7032 (N_7032,N_4656,N_5310);
nand U7033 (N_7033,N_5970,N_5094);
and U7034 (N_7034,N_4922,N_4080);
nand U7035 (N_7035,N_5876,N_5692);
nor U7036 (N_7036,N_4717,N_4961);
nand U7037 (N_7037,N_4956,N_4970);
nand U7038 (N_7038,N_4956,N_4537);
or U7039 (N_7039,N_4562,N_4532);
nand U7040 (N_7040,N_5110,N_5656);
nand U7041 (N_7041,N_5877,N_4839);
and U7042 (N_7042,N_4862,N_5985);
and U7043 (N_7043,N_5489,N_4953);
and U7044 (N_7044,N_5372,N_4309);
or U7045 (N_7045,N_4297,N_4694);
nand U7046 (N_7046,N_5722,N_4880);
and U7047 (N_7047,N_4118,N_4294);
xor U7048 (N_7048,N_5147,N_5198);
xnor U7049 (N_7049,N_4611,N_5053);
and U7050 (N_7050,N_4069,N_5262);
nand U7051 (N_7051,N_4936,N_4471);
nor U7052 (N_7052,N_5031,N_5560);
or U7053 (N_7053,N_5727,N_4941);
nor U7054 (N_7054,N_5697,N_5722);
nand U7055 (N_7055,N_4432,N_5566);
nor U7056 (N_7056,N_4120,N_5078);
or U7057 (N_7057,N_5519,N_4429);
and U7058 (N_7058,N_5946,N_5179);
or U7059 (N_7059,N_4057,N_4882);
nand U7060 (N_7060,N_5061,N_5578);
and U7061 (N_7061,N_5375,N_5592);
nand U7062 (N_7062,N_5903,N_5905);
or U7063 (N_7063,N_5610,N_4805);
or U7064 (N_7064,N_4330,N_5695);
or U7065 (N_7065,N_5461,N_5168);
or U7066 (N_7066,N_5143,N_4583);
or U7067 (N_7067,N_5938,N_4010);
or U7068 (N_7068,N_5187,N_4752);
and U7069 (N_7069,N_4703,N_4064);
and U7070 (N_7070,N_5954,N_5377);
nor U7071 (N_7071,N_5792,N_4314);
and U7072 (N_7072,N_4568,N_5981);
nand U7073 (N_7073,N_5767,N_5694);
or U7074 (N_7074,N_4443,N_5585);
and U7075 (N_7075,N_5772,N_4474);
or U7076 (N_7076,N_4308,N_4919);
xnor U7077 (N_7077,N_4924,N_5244);
nand U7078 (N_7078,N_4249,N_5978);
nor U7079 (N_7079,N_5070,N_4271);
and U7080 (N_7080,N_4953,N_5923);
and U7081 (N_7081,N_5265,N_4443);
nor U7082 (N_7082,N_4733,N_4210);
or U7083 (N_7083,N_4009,N_4983);
nand U7084 (N_7084,N_4979,N_5094);
nor U7085 (N_7085,N_4176,N_4876);
or U7086 (N_7086,N_4481,N_5172);
and U7087 (N_7087,N_5702,N_5561);
nor U7088 (N_7088,N_4880,N_4973);
or U7089 (N_7089,N_4815,N_4309);
nand U7090 (N_7090,N_4381,N_4671);
nand U7091 (N_7091,N_5928,N_4386);
and U7092 (N_7092,N_5288,N_4685);
nand U7093 (N_7093,N_5767,N_5713);
and U7094 (N_7094,N_4204,N_5741);
or U7095 (N_7095,N_5165,N_4789);
xor U7096 (N_7096,N_4917,N_4064);
and U7097 (N_7097,N_5582,N_4684);
nand U7098 (N_7098,N_5867,N_4014);
nor U7099 (N_7099,N_5721,N_4445);
nor U7100 (N_7100,N_5656,N_4304);
nor U7101 (N_7101,N_4186,N_5243);
nand U7102 (N_7102,N_4063,N_5024);
and U7103 (N_7103,N_4914,N_5606);
nor U7104 (N_7104,N_5278,N_5655);
nor U7105 (N_7105,N_4485,N_5898);
nor U7106 (N_7106,N_5153,N_5244);
and U7107 (N_7107,N_4698,N_5226);
or U7108 (N_7108,N_5172,N_4994);
nor U7109 (N_7109,N_4781,N_5962);
nor U7110 (N_7110,N_5195,N_5868);
or U7111 (N_7111,N_5875,N_4576);
xor U7112 (N_7112,N_4022,N_4303);
or U7113 (N_7113,N_5051,N_5264);
nand U7114 (N_7114,N_4892,N_4952);
nor U7115 (N_7115,N_4323,N_4026);
nand U7116 (N_7116,N_5914,N_4078);
and U7117 (N_7117,N_4109,N_5620);
or U7118 (N_7118,N_5560,N_5660);
xnor U7119 (N_7119,N_4118,N_4932);
and U7120 (N_7120,N_5063,N_5582);
or U7121 (N_7121,N_4197,N_5118);
xnor U7122 (N_7122,N_5406,N_5881);
xor U7123 (N_7123,N_5610,N_4252);
or U7124 (N_7124,N_4934,N_5754);
and U7125 (N_7125,N_4648,N_5534);
xnor U7126 (N_7126,N_4371,N_4247);
nand U7127 (N_7127,N_4799,N_4236);
nand U7128 (N_7128,N_5215,N_5194);
nor U7129 (N_7129,N_5370,N_5552);
xor U7130 (N_7130,N_4914,N_5051);
nor U7131 (N_7131,N_5867,N_5292);
nand U7132 (N_7132,N_4306,N_5913);
or U7133 (N_7133,N_5747,N_4991);
nor U7134 (N_7134,N_4665,N_5387);
or U7135 (N_7135,N_5560,N_4250);
and U7136 (N_7136,N_4449,N_5838);
or U7137 (N_7137,N_5119,N_5305);
or U7138 (N_7138,N_4043,N_4760);
nor U7139 (N_7139,N_5622,N_4325);
or U7140 (N_7140,N_4981,N_4679);
or U7141 (N_7141,N_4638,N_5658);
and U7142 (N_7142,N_5362,N_5840);
nand U7143 (N_7143,N_4939,N_5862);
and U7144 (N_7144,N_5005,N_5407);
or U7145 (N_7145,N_4254,N_4134);
nor U7146 (N_7146,N_4061,N_4796);
xor U7147 (N_7147,N_4490,N_4831);
and U7148 (N_7148,N_5574,N_4894);
and U7149 (N_7149,N_4339,N_4804);
and U7150 (N_7150,N_5842,N_5837);
and U7151 (N_7151,N_4768,N_5027);
and U7152 (N_7152,N_5867,N_4282);
or U7153 (N_7153,N_4567,N_5647);
nor U7154 (N_7154,N_4491,N_4298);
and U7155 (N_7155,N_5541,N_4196);
nor U7156 (N_7156,N_5916,N_4974);
nor U7157 (N_7157,N_4289,N_4561);
nor U7158 (N_7158,N_4773,N_4941);
and U7159 (N_7159,N_5503,N_5800);
xnor U7160 (N_7160,N_5533,N_4300);
nand U7161 (N_7161,N_4921,N_4627);
nor U7162 (N_7162,N_4979,N_5100);
nand U7163 (N_7163,N_4061,N_4625);
and U7164 (N_7164,N_4152,N_4439);
xor U7165 (N_7165,N_4648,N_4867);
nor U7166 (N_7166,N_4289,N_4269);
or U7167 (N_7167,N_4527,N_4500);
nor U7168 (N_7168,N_4633,N_4353);
and U7169 (N_7169,N_4330,N_5373);
nor U7170 (N_7170,N_4569,N_5255);
or U7171 (N_7171,N_5208,N_5281);
xnor U7172 (N_7172,N_5385,N_4850);
xnor U7173 (N_7173,N_4564,N_5652);
or U7174 (N_7174,N_5758,N_4604);
or U7175 (N_7175,N_5409,N_5597);
nand U7176 (N_7176,N_5804,N_5329);
nand U7177 (N_7177,N_4925,N_5762);
and U7178 (N_7178,N_4539,N_5852);
and U7179 (N_7179,N_5289,N_4095);
xnor U7180 (N_7180,N_4145,N_4252);
or U7181 (N_7181,N_5684,N_5847);
xor U7182 (N_7182,N_4317,N_4767);
or U7183 (N_7183,N_5295,N_5917);
or U7184 (N_7184,N_4612,N_5650);
nor U7185 (N_7185,N_4315,N_4014);
xor U7186 (N_7186,N_4193,N_5896);
or U7187 (N_7187,N_4636,N_5003);
nand U7188 (N_7188,N_4331,N_5730);
nand U7189 (N_7189,N_5251,N_4699);
or U7190 (N_7190,N_5710,N_4012);
nor U7191 (N_7191,N_5372,N_4923);
nor U7192 (N_7192,N_5519,N_5297);
nor U7193 (N_7193,N_5881,N_4433);
nor U7194 (N_7194,N_5266,N_4187);
xor U7195 (N_7195,N_5400,N_5133);
nor U7196 (N_7196,N_4160,N_5856);
xor U7197 (N_7197,N_4734,N_4801);
or U7198 (N_7198,N_4096,N_5596);
and U7199 (N_7199,N_4891,N_5548);
and U7200 (N_7200,N_5799,N_4850);
nand U7201 (N_7201,N_4298,N_4288);
xor U7202 (N_7202,N_5689,N_4093);
nor U7203 (N_7203,N_4614,N_4126);
and U7204 (N_7204,N_5455,N_5583);
or U7205 (N_7205,N_4714,N_5907);
and U7206 (N_7206,N_5344,N_5253);
or U7207 (N_7207,N_4179,N_4249);
or U7208 (N_7208,N_4280,N_4609);
nand U7209 (N_7209,N_5095,N_5162);
xor U7210 (N_7210,N_4287,N_4818);
nand U7211 (N_7211,N_4337,N_4771);
nand U7212 (N_7212,N_4508,N_5289);
nor U7213 (N_7213,N_5173,N_4774);
nand U7214 (N_7214,N_5982,N_4598);
nand U7215 (N_7215,N_5395,N_4826);
or U7216 (N_7216,N_5222,N_4946);
nand U7217 (N_7217,N_5495,N_5834);
nor U7218 (N_7218,N_5591,N_5598);
nand U7219 (N_7219,N_4944,N_5072);
or U7220 (N_7220,N_5273,N_4361);
nand U7221 (N_7221,N_4536,N_4617);
nor U7222 (N_7222,N_4080,N_4776);
nand U7223 (N_7223,N_4823,N_5484);
xnor U7224 (N_7224,N_4562,N_4257);
and U7225 (N_7225,N_5453,N_5084);
xnor U7226 (N_7226,N_5947,N_5530);
or U7227 (N_7227,N_5338,N_5779);
or U7228 (N_7228,N_4017,N_4734);
nor U7229 (N_7229,N_4476,N_5543);
and U7230 (N_7230,N_4018,N_5287);
nor U7231 (N_7231,N_4029,N_4225);
or U7232 (N_7232,N_5112,N_5782);
nor U7233 (N_7233,N_5873,N_4394);
and U7234 (N_7234,N_4540,N_5547);
nand U7235 (N_7235,N_4248,N_5630);
nand U7236 (N_7236,N_5025,N_4454);
and U7237 (N_7237,N_4615,N_5054);
and U7238 (N_7238,N_4738,N_4923);
nand U7239 (N_7239,N_5755,N_5268);
or U7240 (N_7240,N_4915,N_4162);
and U7241 (N_7241,N_5192,N_5565);
and U7242 (N_7242,N_5869,N_5666);
nor U7243 (N_7243,N_5043,N_4724);
nand U7244 (N_7244,N_4788,N_4688);
and U7245 (N_7245,N_4703,N_5204);
nor U7246 (N_7246,N_4397,N_5614);
or U7247 (N_7247,N_5040,N_4486);
or U7248 (N_7248,N_5719,N_4408);
nor U7249 (N_7249,N_5884,N_5565);
or U7250 (N_7250,N_4837,N_5521);
and U7251 (N_7251,N_5608,N_5343);
nor U7252 (N_7252,N_4591,N_5793);
and U7253 (N_7253,N_5510,N_4378);
nand U7254 (N_7254,N_5986,N_4939);
or U7255 (N_7255,N_5159,N_5271);
nand U7256 (N_7256,N_5857,N_4593);
nand U7257 (N_7257,N_4111,N_5479);
nor U7258 (N_7258,N_4684,N_4522);
and U7259 (N_7259,N_5300,N_5332);
or U7260 (N_7260,N_4788,N_5918);
nor U7261 (N_7261,N_5674,N_5226);
and U7262 (N_7262,N_4319,N_4261);
nand U7263 (N_7263,N_5870,N_4966);
and U7264 (N_7264,N_5609,N_5644);
or U7265 (N_7265,N_4859,N_4247);
nor U7266 (N_7266,N_4848,N_4520);
xor U7267 (N_7267,N_5818,N_5519);
or U7268 (N_7268,N_5429,N_4810);
and U7269 (N_7269,N_4758,N_4659);
xor U7270 (N_7270,N_4504,N_5599);
and U7271 (N_7271,N_4836,N_5805);
nor U7272 (N_7272,N_5139,N_5111);
xor U7273 (N_7273,N_4612,N_4508);
nand U7274 (N_7274,N_4532,N_5764);
nand U7275 (N_7275,N_4454,N_4262);
nor U7276 (N_7276,N_5884,N_4910);
xor U7277 (N_7277,N_4323,N_5307);
nor U7278 (N_7278,N_5115,N_5525);
nor U7279 (N_7279,N_5046,N_4363);
nor U7280 (N_7280,N_5874,N_4876);
and U7281 (N_7281,N_5146,N_4827);
and U7282 (N_7282,N_4143,N_5230);
and U7283 (N_7283,N_4702,N_5144);
and U7284 (N_7284,N_5390,N_5892);
nor U7285 (N_7285,N_4968,N_5139);
nor U7286 (N_7286,N_4838,N_5818);
or U7287 (N_7287,N_5662,N_4105);
and U7288 (N_7288,N_4603,N_5349);
nand U7289 (N_7289,N_4296,N_5327);
nor U7290 (N_7290,N_4408,N_4199);
nor U7291 (N_7291,N_5843,N_5610);
or U7292 (N_7292,N_5659,N_4423);
nand U7293 (N_7293,N_4738,N_4464);
nand U7294 (N_7294,N_4735,N_4468);
xnor U7295 (N_7295,N_4227,N_5007);
or U7296 (N_7296,N_4200,N_5485);
and U7297 (N_7297,N_5644,N_4507);
nand U7298 (N_7298,N_5918,N_4600);
nand U7299 (N_7299,N_4975,N_4619);
and U7300 (N_7300,N_5503,N_5854);
nor U7301 (N_7301,N_4890,N_5991);
nand U7302 (N_7302,N_4898,N_4750);
and U7303 (N_7303,N_4498,N_4529);
or U7304 (N_7304,N_4928,N_4335);
and U7305 (N_7305,N_5916,N_4910);
xnor U7306 (N_7306,N_5203,N_4128);
and U7307 (N_7307,N_5977,N_4780);
or U7308 (N_7308,N_5249,N_4296);
xnor U7309 (N_7309,N_4072,N_5244);
and U7310 (N_7310,N_5593,N_4936);
xnor U7311 (N_7311,N_5605,N_5995);
nand U7312 (N_7312,N_5453,N_5930);
xor U7313 (N_7313,N_4294,N_4023);
xor U7314 (N_7314,N_4496,N_5925);
or U7315 (N_7315,N_4969,N_5148);
and U7316 (N_7316,N_4330,N_4543);
nor U7317 (N_7317,N_5829,N_5610);
or U7318 (N_7318,N_5169,N_5870);
nand U7319 (N_7319,N_5459,N_4164);
or U7320 (N_7320,N_4693,N_4750);
nand U7321 (N_7321,N_4091,N_4925);
or U7322 (N_7322,N_5793,N_5731);
and U7323 (N_7323,N_5233,N_4442);
and U7324 (N_7324,N_5019,N_4774);
xor U7325 (N_7325,N_4797,N_4221);
or U7326 (N_7326,N_4647,N_5846);
xor U7327 (N_7327,N_5799,N_5913);
nor U7328 (N_7328,N_4611,N_5282);
nand U7329 (N_7329,N_5935,N_5113);
nand U7330 (N_7330,N_4284,N_5744);
nor U7331 (N_7331,N_5737,N_4818);
and U7332 (N_7332,N_5443,N_4264);
or U7333 (N_7333,N_5286,N_5742);
nor U7334 (N_7334,N_4693,N_5444);
and U7335 (N_7335,N_4227,N_5257);
nor U7336 (N_7336,N_5170,N_5096);
or U7337 (N_7337,N_5406,N_4990);
nor U7338 (N_7338,N_4322,N_5888);
and U7339 (N_7339,N_4959,N_5522);
nor U7340 (N_7340,N_5806,N_4306);
nor U7341 (N_7341,N_4160,N_4357);
nand U7342 (N_7342,N_5181,N_4709);
or U7343 (N_7343,N_5224,N_4899);
nor U7344 (N_7344,N_4587,N_4313);
nor U7345 (N_7345,N_4002,N_4669);
and U7346 (N_7346,N_4440,N_4754);
or U7347 (N_7347,N_4163,N_5732);
nand U7348 (N_7348,N_4895,N_4692);
or U7349 (N_7349,N_5618,N_4031);
xnor U7350 (N_7350,N_4079,N_5348);
nand U7351 (N_7351,N_5018,N_5133);
nor U7352 (N_7352,N_5020,N_5745);
nor U7353 (N_7353,N_5604,N_5750);
xnor U7354 (N_7354,N_4530,N_5174);
nor U7355 (N_7355,N_4813,N_5411);
and U7356 (N_7356,N_4361,N_4976);
nor U7357 (N_7357,N_5355,N_4892);
nand U7358 (N_7358,N_5229,N_4377);
nand U7359 (N_7359,N_5827,N_5859);
or U7360 (N_7360,N_5260,N_4610);
or U7361 (N_7361,N_4345,N_4962);
nand U7362 (N_7362,N_4856,N_4447);
or U7363 (N_7363,N_5671,N_4589);
nor U7364 (N_7364,N_4517,N_4057);
nand U7365 (N_7365,N_5729,N_4425);
xnor U7366 (N_7366,N_4386,N_4758);
and U7367 (N_7367,N_5572,N_5450);
and U7368 (N_7368,N_5682,N_4546);
nand U7369 (N_7369,N_5820,N_4906);
nand U7370 (N_7370,N_5094,N_4201);
and U7371 (N_7371,N_5353,N_4184);
nand U7372 (N_7372,N_4649,N_5672);
or U7373 (N_7373,N_5246,N_4326);
and U7374 (N_7374,N_4856,N_4112);
xor U7375 (N_7375,N_4826,N_5270);
and U7376 (N_7376,N_4957,N_4402);
and U7377 (N_7377,N_4759,N_4775);
xnor U7378 (N_7378,N_5905,N_4361);
nor U7379 (N_7379,N_4269,N_4750);
and U7380 (N_7380,N_4926,N_4193);
and U7381 (N_7381,N_4348,N_4806);
and U7382 (N_7382,N_5399,N_4884);
nor U7383 (N_7383,N_4283,N_5359);
nor U7384 (N_7384,N_5404,N_4390);
nor U7385 (N_7385,N_4554,N_4271);
nor U7386 (N_7386,N_5622,N_4598);
nor U7387 (N_7387,N_5126,N_5475);
and U7388 (N_7388,N_4635,N_5900);
nor U7389 (N_7389,N_5005,N_5934);
nor U7390 (N_7390,N_5950,N_5079);
nor U7391 (N_7391,N_5490,N_5005);
nand U7392 (N_7392,N_4061,N_4130);
nand U7393 (N_7393,N_4304,N_5124);
xnor U7394 (N_7394,N_5546,N_5489);
or U7395 (N_7395,N_5813,N_5651);
nand U7396 (N_7396,N_4710,N_5122);
or U7397 (N_7397,N_5371,N_4850);
nor U7398 (N_7398,N_5145,N_4587);
or U7399 (N_7399,N_5280,N_5183);
xor U7400 (N_7400,N_4242,N_5596);
xnor U7401 (N_7401,N_4120,N_5645);
nor U7402 (N_7402,N_5753,N_5814);
nor U7403 (N_7403,N_4409,N_4167);
nand U7404 (N_7404,N_4003,N_5227);
or U7405 (N_7405,N_4616,N_4612);
and U7406 (N_7406,N_4915,N_4861);
nor U7407 (N_7407,N_4491,N_5214);
xor U7408 (N_7408,N_5297,N_4737);
or U7409 (N_7409,N_4983,N_5664);
nand U7410 (N_7410,N_5076,N_4975);
nor U7411 (N_7411,N_4137,N_4463);
or U7412 (N_7412,N_5195,N_5877);
and U7413 (N_7413,N_5838,N_4495);
nand U7414 (N_7414,N_4934,N_4984);
nand U7415 (N_7415,N_5799,N_4752);
or U7416 (N_7416,N_5186,N_5191);
nor U7417 (N_7417,N_5440,N_5522);
nand U7418 (N_7418,N_5770,N_4398);
nor U7419 (N_7419,N_5728,N_4705);
or U7420 (N_7420,N_5647,N_4874);
or U7421 (N_7421,N_4678,N_5195);
and U7422 (N_7422,N_5560,N_5765);
or U7423 (N_7423,N_4374,N_5252);
nor U7424 (N_7424,N_5502,N_4210);
and U7425 (N_7425,N_5675,N_4923);
nor U7426 (N_7426,N_5616,N_5579);
nand U7427 (N_7427,N_5853,N_5197);
nor U7428 (N_7428,N_5252,N_5306);
nand U7429 (N_7429,N_4722,N_5022);
nor U7430 (N_7430,N_4067,N_4698);
nor U7431 (N_7431,N_4715,N_4018);
nor U7432 (N_7432,N_5994,N_4365);
and U7433 (N_7433,N_5805,N_5763);
nand U7434 (N_7434,N_4052,N_4613);
or U7435 (N_7435,N_5259,N_5324);
or U7436 (N_7436,N_4350,N_4783);
nand U7437 (N_7437,N_4151,N_5801);
and U7438 (N_7438,N_4685,N_5422);
nor U7439 (N_7439,N_5819,N_4024);
nand U7440 (N_7440,N_4083,N_4321);
or U7441 (N_7441,N_5003,N_4641);
and U7442 (N_7442,N_4204,N_4287);
nor U7443 (N_7443,N_4164,N_5011);
nor U7444 (N_7444,N_5493,N_5056);
xnor U7445 (N_7445,N_4686,N_4987);
or U7446 (N_7446,N_5235,N_4135);
nor U7447 (N_7447,N_5263,N_4831);
or U7448 (N_7448,N_5273,N_5358);
xnor U7449 (N_7449,N_5832,N_5124);
xnor U7450 (N_7450,N_5098,N_5965);
or U7451 (N_7451,N_5339,N_5194);
nor U7452 (N_7452,N_5601,N_5668);
nor U7453 (N_7453,N_5555,N_5441);
or U7454 (N_7454,N_4421,N_5954);
and U7455 (N_7455,N_5413,N_5023);
and U7456 (N_7456,N_5299,N_5730);
nor U7457 (N_7457,N_4467,N_5251);
nor U7458 (N_7458,N_5773,N_5427);
or U7459 (N_7459,N_5190,N_4687);
nand U7460 (N_7460,N_5503,N_4810);
or U7461 (N_7461,N_5962,N_4669);
or U7462 (N_7462,N_4033,N_4909);
nor U7463 (N_7463,N_4800,N_5464);
and U7464 (N_7464,N_4506,N_5586);
nor U7465 (N_7465,N_5662,N_5868);
or U7466 (N_7466,N_5528,N_5211);
nand U7467 (N_7467,N_5353,N_4419);
xor U7468 (N_7468,N_4446,N_4185);
xor U7469 (N_7469,N_4769,N_5688);
and U7470 (N_7470,N_5905,N_4887);
or U7471 (N_7471,N_5304,N_4291);
or U7472 (N_7472,N_5762,N_5724);
and U7473 (N_7473,N_5081,N_5380);
nand U7474 (N_7474,N_4920,N_4424);
nor U7475 (N_7475,N_5751,N_4315);
and U7476 (N_7476,N_5898,N_5084);
nand U7477 (N_7477,N_5437,N_5743);
and U7478 (N_7478,N_4854,N_5936);
or U7479 (N_7479,N_5590,N_5189);
and U7480 (N_7480,N_5209,N_5097);
nor U7481 (N_7481,N_5266,N_5655);
or U7482 (N_7482,N_5380,N_4886);
and U7483 (N_7483,N_5931,N_5770);
or U7484 (N_7484,N_4045,N_5625);
or U7485 (N_7485,N_5100,N_5942);
nand U7486 (N_7486,N_5705,N_5056);
or U7487 (N_7487,N_4577,N_4603);
or U7488 (N_7488,N_5627,N_4238);
and U7489 (N_7489,N_4453,N_5559);
nor U7490 (N_7490,N_5795,N_5060);
nor U7491 (N_7491,N_4806,N_4542);
xor U7492 (N_7492,N_4526,N_4884);
or U7493 (N_7493,N_4996,N_5695);
and U7494 (N_7494,N_4892,N_4152);
and U7495 (N_7495,N_4446,N_4218);
or U7496 (N_7496,N_5380,N_5460);
or U7497 (N_7497,N_4386,N_5882);
and U7498 (N_7498,N_5539,N_4975);
nor U7499 (N_7499,N_5034,N_4394);
nor U7500 (N_7500,N_4053,N_5007);
xnor U7501 (N_7501,N_5570,N_4292);
xnor U7502 (N_7502,N_4253,N_4992);
or U7503 (N_7503,N_4760,N_4796);
or U7504 (N_7504,N_5525,N_5523);
or U7505 (N_7505,N_5835,N_4902);
or U7506 (N_7506,N_5013,N_4284);
nor U7507 (N_7507,N_4356,N_5875);
nor U7508 (N_7508,N_4296,N_5651);
and U7509 (N_7509,N_5454,N_4117);
nor U7510 (N_7510,N_4943,N_5732);
nand U7511 (N_7511,N_4999,N_4610);
xor U7512 (N_7512,N_5903,N_5430);
or U7513 (N_7513,N_5673,N_4331);
nand U7514 (N_7514,N_4324,N_5808);
and U7515 (N_7515,N_4969,N_4674);
nand U7516 (N_7516,N_5689,N_5173);
nand U7517 (N_7517,N_5027,N_5294);
or U7518 (N_7518,N_4503,N_4262);
nor U7519 (N_7519,N_5377,N_5917);
nor U7520 (N_7520,N_5958,N_5737);
xnor U7521 (N_7521,N_5493,N_5059);
or U7522 (N_7522,N_4277,N_5991);
nor U7523 (N_7523,N_5771,N_4090);
xor U7524 (N_7524,N_5408,N_5562);
nand U7525 (N_7525,N_4571,N_4691);
xnor U7526 (N_7526,N_4307,N_4933);
or U7527 (N_7527,N_4179,N_4828);
or U7528 (N_7528,N_5351,N_5898);
nand U7529 (N_7529,N_4733,N_4217);
or U7530 (N_7530,N_4793,N_4774);
and U7531 (N_7531,N_5619,N_5594);
nor U7532 (N_7532,N_5555,N_5404);
nor U7533 (N_7533,N_4914,N_5530);
or U7534 (N_7534,N_4609,N_4706);
nor U7535 (N_7535,N_5596,N_5477);
nor U7536 (N_7536,N_5906,N_4334);
nor U7537 (N_7537,N_5212,N_5252);
or U7538 (N_7538,N_4402,N_4653);
or U7539 (N_7539,N_4870,N_4115);
and U7540 (N_7540,N_4241,N_5115);
nor U7541 (N_7541,N_5803,N_5463);
and U7542 (N_7542,N_4825,N_4131);
or U7543 (N_7543,N_5345,N_4450);
nor U7544 (N_7544,N_5748,N_4601);
or U7545 (N_7545,N_5073,N_5131);
and U7546 (N_7546,N_5108,N_4633);
nor U7547 (N_7547,N_5083,N_4255);
xor U7548 (N_7548,N_5453,N_5748);
or U7549 (N_7549,N_4266,N_5183);
nand U7550 (N_7550,N_4912,N_4058);
nor U7551 (N_7551,N_5663,N_4779);
nand U7552 (N_7552,N_4871,N_5420);
and U7553 (N_7553,N_4092,N_4598);
xor U7554 (N_7554,N_5275,N_5513);
or U7555 (N_7555,N_5825,N_4009);
xor U7556 (N_7556,N_5734,N_5308);
and U7557 (N_7557,N_4821,N_5249);
nor U7558 (N_7558,N_4599,N_4620);
nand U7559 (N_7559,N_4810,N_4870);
or U7560 (N_7560,N_4901,N_4210);
nor U7561 (N_7561,N_5542,N_5149);
or U7562 (N_7562,N_5629,N_4990);
and U7563 (N_7563,N_4106,N_5647);
xor U7564 (N_7564,N_5359,N_5728);
nor U7565 (N_7565,N_5356,N_5103);
xnor U7566 (N_7566,N_5902,N_4014);
nand U7567 (N_7567,N_4963,N_5663);
or U7568 (N_7568,N_5447,N_5533);
nand U7569 (N_7569,N_4243,N_5852);
nor U7570 (N_7570,N_4006,N_5491);
or U7571 (N_7571,N_4209,N_4294);
nand U7572 (N_7572,N_4838,N_4293);
nand U7573 (N_7573,N_5334,N_5500);
or U7574 (N_7574,N_4233,N_4822);
nand U7575 (N_7575,N_4223,N_4632);
or U7576 (N_7576,N_4909,N_4217);
or U7577 (N_7577,N_4382,N_4576);
and U7578 (N_7578,N_4981,N_4226);
nand U7579 (N_7579,N_5827,N_5544);
or U7580 (N_7580,N_4804,N_5184);
and U7581 (N_7581,N_5419,N_5172);
or U7582 (N_7582,N_5409,N_4157);
or U7583 (N_7583,N_5277,N_5616);
or U7584 (N_7584,N_5290,N_4524);
nor U7585 (N_7585,N_4625,N_4666);
nor U7586 (N_7586,N_5352,N_5140);
nor U7587 (N_7587,N_5379,N_5099);
and U7588 (N_7588,N_4762,N_4967);
or U7589 (N_7589,N_5951,N_5968);
nor U7590 (N_7590,N_4953,N_5201);
or U7591 (N_7591,N_5128,N_5653);
nand U7592 (N_7592,N_5662,N_4013);
nor U7593 (N_7593,N_4516,N_4450);
or U7594 (N_7594,N_5277,N_4789);
or U7595 (N_7595,N_5547,N_4692);
or U7596 (N_7596,N_5827,N_5161);
or U7597 (N_7597,N_5524,N_5631);
nor U7598 (N_7598,N_4450,N_4091);
and U7599 (N_7599,N_5434,N_4120);
and U7600 (N_7600,N_4770,N_4586);
nor U7601 (N_7601,N_5434,N_5565);
or U7602 (N_7602,N_4396,N_4851);
or U7603 (N_7603,N_4841,N_5893);
xor U7604 (N_7604,N_4537,N_4221);
nand U7605 (N_7605,N_5285,N_4552);
or U7606 (N_7606,N_5919,N_4264);
or U7607 (N_7607,N_4856,N_5401);
and U7608 (N_7608,N_4547,N_5442);
and U7609 (N_7609,N_5326,N_5799);
and U7610 (N_7610,N_5636,N_4538);
nor U7611 (N_7611,N_4770,N_5781);
nand U7612 (N_7612,N_5155,N_5801);
nor U7613 (N_7613,N_4664,N_4236);
and U7614 (N_7614,N_4932,N_4839);
nor U7615 (N_7615,N_4199,N_4828);
xor U7616 (N_7616,N_5759,N_4281);
and U7617 (N_7617,N_4046,N_5882);
nor U7618 (N_7618,N_5119,N_5744);
or U7619 (N_7619,N_5450,N_4814);
nor U7620 (N_7620,N_4704,N_4566);
nand U7621 (N_7621,N_4057,N_4205);
and U7622 (N_7622,N_5236,N_4444);
or U7623 (N_7623,N_4659,N_4262);
nor U7624 (N_7624,N_4991,N_5964);
nand U7625 (N_7625,N_5519,N_4386);
or U7626 (N_7626,N_4047,N_4314);
and U7627 (N_7627,N_4961,N_4732);
xor U7628 (N_7628,N_4301,N_4607);
nand U7629 (N_7629,N_5765,N_4266);
and U7630 (N_7630,N_5180,N_5437);
or U7631 (N_7631,N_4969,N_4823);
nand U7632 (N_7632,N_4215,N_4752);
and U7633 (N_7633,N_4573,N_5540);
xnor U7634 (N_7634,N_5789,N_5705);
and U7635 (N_7635,N_5319,N_4877);
or U7636 (N_7636,N_5032,N_5925);
nor U7637 (N_7637,N_4119,N_5542);
and U7638 (N_7638,N_4772,N_4260);
nand U7639 (N_7639,N_4400,N_4647);
xor U7640 (N_7640,N_4233,N_5860);
and U7641 (N_7641,N_5852,N_5887);
or U7642 (N_7642,N_4160,N_5986);
nand U7643 (N_7643,N_5199,N_5419);
and U7644 (N_7644,N_5739,N_4425);
or U7645 (N_7645,N_5744,N_5066);
and U7646 (N_7646,N_4681,N_5290);
or U7647 (N_7647,N_4850,N_5632);
and U7648 (N_7648,N_4962,N_4012);
and U7649 (N_7649,N_4133,N_4108);
or U7650 (N_7650,N_4505,N_4526);
nor U7651 (N_7651,N_5593,N_5654);
or U7652 (N_7652,N_4555,N_4986);
nor U7653 (N_7653,N_4306,N_4983);
or U7654 (N_7654,N_5389,N_5600);
and U7655 (N_7655,N_5661,N_4681);
nor U7656 (N_7656,N_4012,N_4137);
nand U7657 (N_7657,N_4145,N_4349);
and U7658 (N_7658,N_4926,N_5247);
nor U7659 (N_7659,N_5771,N_4197);
nand U7660 (N_7660,N_4090,N_5752);
nand U7661 (N_7661,N_4602,N_4528);
or U7662 (N_7662,N_5720,N_4692);
and U7663 (N_7663,N_5133,N_4598);
nand U7664 (N_7664,N_4252,N_5631);
nand U7665 (N_7665,N_5304,N_5521);
and U7666 (N_7666,N_5227,N_4711);
nor U7667 (N_7667,N_5004,N_5961);
or U7668 (N_7668,N_4519,N_4632);
or U7669 (N_7669,N_5949,N_5559);
nor U7670 (N_7670,N_5428,N_5492);
nand U7671 (N_7671,N_5118,N_5129);
or U7672 (N_7672,N_4969,N_4477);
nor U7673 (N_7673,N_5156,N_4379);
nor U7674 (N_7674,N_4853,N_5246);
nand U7675 (N_7675,N_5527,N_5599);
nand U7676 (N_7676,N_4832,N_5025);
and U7677 (N_7677,N_4902,N_5054);
or U7678 (N_7678,N_5388,N_5196);
and U7679 (N_7679,N_5818,N_5354);
nor U7680 (N_7680,N_4783,N_4577);
xor U7681 (N_7681,N_4278,N_5443);
nor U7682 (N_7682,N_5501,N_5756);
xnor U7683 (N_7683,N_4521,N_5776);
nor U7684 (N_7684,N_4665,N_4749);
nand U7685 (N_7685,N_5635,N_4368);
or U7686 (N_7686,N_4844,N_5653);
nor U7687 (N_7687,N_4987,N_5531);
and U7688 (N_7688,N_5330,N_5752);
nor U7689 (N_7689,N_4879,N_5824);
nand U7690 (N_7690,N_4761,N_5840);
and U7691 (N_7691,N_5413,N_5780);
nand U7692 (N_7692,N_5316,N_5390);
or U7693 (N_7693,N_5850,N_5896);
nor U7694 (N_7694,N_4539,N_4877);
nor U7695 (N_7695,N_5869,N_4885);
or U7696 (N_7696,N_5894,N_5288);
nor U7697 (N_7697,N_4130,N_5799);
or U7698 (N_7698,N_4097,N_5891);
nor U7699 (N_7699,N_4084,N_5714);
nand U7700 (N_7700,N_4226,N_4324);
and U7701 (N_7701,N_5794,N_4966);
nor U7702 (N_7702,N_4495,N_4746);
or U7703 (N_7703,N_5252,N_4423);
or U7704 (N_7704,N_5803,N_4685);
nand U7705 (N_7705,N_4422,N_4440);
nand U7706 (N_7706,N_4932,N_4527);
or U7707 (N_7707,N_4244,N_4691);
or U7708 (N_7708,N_5474,N_5602);
nor U7709 (N_7709,N_4058,N_5768);
xor U7710 (N_7710,N_4232,N_4080);
and U7711 (N_7711,N_4975,N_5346);
or U7712 (N_7712,N_4343,N_4760);
and U7713 (N_7713,N_4875,N_5954);
nand U7714 (N_7714,N_5740,N_5042);
and U7715 (N_7715,N_4877,N_5655);
nand U7716 (N_7716,N_5142,N_5158);
or U7717 (N_7717,N_4880,N_4827);
xnor U7718 (N_7718,N_5136,N_5491);
nand U7719 (N_7719,N_4921,N_4997);
and U7720 (N_7720,N_4645,N_4817);
and U7721 (N_7721,N_4680,N_5943);
or U7722 (N_7722,N_5778,N_5706);
and U7723 (N_7723,N_5092,N_5818);
or U7724 (N_7724,N_4738,N_5845);
nand U7725 (N_7725,N_4539,N_4439);
and U7726 (N_7726,N_4757,N_5679);
and U7727 (N_7727,N_4500,N_4493);
and U7728 (N_7728,N_5091,N_4550);
nor U7729 (N_7729,N_4468,N_4011);
and U7730 (N_7730,N_4111,N_4741);
or U7731 (N_7731,N_5730,N_4020);
nor U7732 (N_7732,N_4169,N_5719);
and U7733 (N_7733,N_5624,N_5786);
and U7734 (N_7734,N_5141,N_4175);
and U7735 (N_7735,N_4948,N_4615);
nor U7736 (N_7736,N_5565,N_5400);
nand U7737 (N_7737,N_5882,N_4258);
nor U7738 (N_7738,N_4522,N_4062);
nand U7739 (N_7739,N_5011,N_5662);
nor U7740 (N_7740,N_5993,N_5547);
nor U7741 (N_7741,N_4988,N_4355);
nor U7742 (N_7742,N_5632,N_4141);
xnor U7743 (N_7743,N_5290,N_5319);
nor U7744 (N_7744,N_4371,N_5564);
or U7745 (N_7745,N_4787,N_4143);
nand U7746 (N_7746,N_4666,N_4136);
and U7747 (N_7747,N_5625,N_5133);
nand U7748 (N_7748,N_5256,N_4844);
or U7749 (N_7749,N_5974,N_5115);
xnor U7750 (N_7750,N_5547,N_5299);
or U7751 (N_7751,N_4390,N_4393);
nand U7752 (N_7752,N_4534,N_5425);
nand U7753 (N_7753,N_5686,N_4149);
nor U7754 (N_7754,N_4242,N_4742);
nor U7755 (N_7755,N_5059,N_5750);
nand U7756 (N_7756,N_5104,N_5036);
xor U7757 (N_7757,N_5119,N_4360);
nor U7758 (N_7758,N_5203,N_5178);
or U7759 (N_7759,N_4710,N_5946);
nand U7760 (N_7760,N_4497,N_5225);
nand U7761 (N_7761,N_4807,N_4298);
nor U7762 (N_7762,N_5454,N_5698);
nand U7763 (N_7763,N_5079,N_5730);
or U7764 (N_7764,N_5886,N_5245);
nor U7765 (N_7765,N_5247,N_4116);
nor U7766 (N_7766,N_5373,N_5143);
and U7767 (N_7767,N_4310,N_5740);
or U7768 (N_7768,N_5862,N_4773);
and U7769 (N_7769,N_5896,N_5722);
nand U7770 (N_7770,N_5916,N_5124);
or U7771 (N_7771,N_5635,N_5942);
xnor U7772 (N_7772,N_5392,N_4912);
nand U7773 (N_7773,N_5798,N_5401);
nor U7774 (N_7774,N_5212,N_4793);
or U7775 (N_7775,N_4531,N_4675);
and U7776 (N_7776,N_4269,N_4671);
or U7777 (N_7777,N_4418,N_4848);
and U7778 (N_7778,N_5402,N_4222);
nor U7779 (N_7779,N_4439,N_4370);
nor U7780 (N_7780,N_4510,N_5991);
nor U7781 (N_7781,N_5144,N_4069);
nor U7782 (N_7782,N_4804,N_4430);
and U7783 (N_7783,N_4877,N_4546);
or U7784 (N_7784,N_5830,N_4677);
nand U7785 (N_7785,N_5882,N_5470);
and U7786 (N_7786,N_4357,N_4800);
or U7787 (N_7787,N_4521,N_4275);
nor U7788 (N_7788,N_4269,N_4831);
nor U7789 (N_7789,N_4127,N_4643);
nor U7790 (N_7790,N_5401,N_4217);
nand U7791 (N_7791,N_5989,N_5018);
nand U7792 (N_7792,N_5931,N_4329);
or U7793 (N_7793,N_5345,N_5459);
or U7794 (N_7794,N_5291,N_4650);
nor U7795 (N_7795,N_5276,N_5958);
nand U7796 (N_7796,N_4415,N_4391);
nor U7797 (N_7797,N_5522,N_4885);
or U7798 (N_7798,N_5483,N_4424);
and U7799 (N_7799,N_5737,N_4483);
nor U7800 (N_7800,N_4665,N_5695);
xor U7801 (N_7801,N_4121,N_5559);
nand U7802 (N_7802,N_5014,N_4704);
nor U7803 (N_7803,N_5834,N_5533);
nor U7804 (N_7804,N_4104,N_4667);
nor U7805 (N_7805,N_4372,N_4699);
or U7806 (N_7806,N_5686,N_5476);
or U7807 (N_7807,N_5313,N_4904);
nor U7808 (N_7808,N_4808,N_5570);
or U7809 (N_7809,N_5951,N_4085);
nor U7810 (N_7810,N_5978,N_5577);
nor U7811 (N_7811,N_5717,N_5956);
nand U7812 (N_7812,N_5787,N_4158);
and U7813 (N_7813,N_5212,N_5725);
nand U7814 (N_7814,N_5826,N_4678);
or U7815 (N_7815,N_5990,N_5216);
nand U7816 (N_7816,N_5740,N_5726);
nand U7817 (N_7817,N_4010,N_4762);
nor U7818 (N_7818,N_4779,N_5346);
nand U7819 (N_7819,N_5176,N_4063);
and U7820 (N_7820,N_5854,N_4314);
nor U7821 (N_7821,N_4112,N_5092);
nor U7822 (N_7822,N_4351,N_4022);
and U7823 (N_7823,N_5886,N_4151);
nand U7824 (N_7824,N_5516,N_5888);
or U7825 (N_7825,N_5001,N_4055);
nor U7826 (N_7826,N_5039,N_4951);
and U7827 (N_7827,N_5564,N_4588);
nor U7828 (N_7828,N_4184,N_5059);
nand U7829 (N_7829,N_5694,N_4950);
xnor U7830 (N_7830,N_4576,N_4675);
nor U7831 (N_7831,N_5924,N_5932);
nor U7832 (N_7832,N_4879,N_5730);
nand U7833 (N_7833,N_5971,N_5455);
nand U7834 (N_7834,N_4875,N_4595);
or U7835 (N_7835,N_4324,N_5944);
nor U7836 (N_7836,N_5829,N_5406);
or U7837 (N_7837,N_4778,N_5458);
and U7838 (N_7838,N_5462,N_5346);
and U7839 (N_7839,N_4807,N_5922);
or U7840 (N_7840,N_4872,N_5318);
nor U7841 (N_7841,N_5560,N_5195);
or U7842 (N_7842,N_4257,N_4894);
or U7843 (N_7843,N_5947,N_5642);
nor U7844 (N_7844,N_5595,N_5709);
nor U7845 (N_7845,N_4763,N_5281);
or U7846 (N_7846,N_4468,N_5576);
and U7847 (N_7847,N_4970,N_4622);
nor U7848 (N_7848,N_4965,N_5364);
nand U7849 (N_7849,N_4449,N_4532);
or U7850 (N_7850,N_4840,N_4943);
and U7851 (N_7851,N_5845,N_5683);
or U7852 (N_7852,N_5138,N_5629);
and U7853 (N_7853,N_5245,N_5023);
nor U7854 (N_7854,N_4522,N_4195);
xor U7855 (N_7855,N_5703,N_5732);
nor U7856 (N_7856,N_4268,N_4696);
and U7857 (N_7857,N_5070,N_4944);
xnor U7858 (N_7858,N_4838,N_4181);
and U7859 (N_7859,N_4647,N_4845);
and U7860 (N_7860,N_5102,N_5746);
nand U7861 (N_7861,N_5596,N_4998);
nor U7862 (N_7862,N_5543,N_5031);
nor U7863 (N_7863,N_4416,N_4664);
nand U7864 (N_7864,N_4946,N_4944);
xor U7865 (N_7865,N_5250,N_4261);
nor U7866 (N_7866,N_5823,N_4965);
or U7867 (N_7867,N_5498,N_4471);
or U7868 (N_7868,N_5682,N_5923);
xnor U7869 (N_7869,N_5162,N_5435);
nand U7870 (N_7870,N_5575,N_4270);
and U7871 (N_7871,N_4974,N_4254);
and U7872 (N_7872,N_5463,N_4962);
or U7873 (N_7873,N_4963,N_5747);
nor U7874 (N_7874,N_4733,N_4579);
nand U7875 (N_7875,N_4996,N_4446);
and U7876 (N_7876,N_5668,N_4953);
nand U7877 (N_7877,N_4380,N_4499);
nand U7878 (N_7878,N_5769,N_4939);
xnor U7879 (N_7879,N_4158,N_4581);
or U7880 (N_7880,N_4367,N_4231);
and U7881 (N_7881,N_5214,N_4854);
and U7882 (N_7882,N_5354,N_5583);
or U7883 (N_7883,N_4283,N_5126);
nor U7884 (N_7884,N_4279,N_4097);
nor U7885 (N_7885,N_5257,N_4751);
or U7886 (N_7886,N_4251,N_4548);
or U7887 (N_7887,N_4090,N_4305);
nor U7888 (N_7888,N_4753,N_5950);
nand U7889 (N_7889,N_5838,N_4028);
nor U7890 (N_7890,N_5695,N_4346);
nand U7891 (N_7891,N_4765,N_5657);
nor U7892 (N_7892,N_5337,N_4891);
and U7893 (N_7893,N_5856,N_4068);
and U7894 (N_7894,N_4594,N_4262);
nand U7895 (N_7895,N_4876,N_5913);
nor U7896 (N_7896,N_4079,N_5152);
nor U7897 (N_7897,N_4136,N_5356);
or U7898 (N_7898,N_5821,N_4400);
or U7899 (N_7899,N_5005,N_5563);
xnor U7900 (N_7900,N_4726,N_4045);
xor U7901 (N_7901,N_5516,N_5145);
nor U7902 (N_7902,N_5305,N_4753);
and U7903 (N_7903,N_5189,N_5609);
or U7904 (N_7904,N_5587,N_5796);
xnor U7905 (N_7905,N_5247,N_4099);
or U7906 (N_7906,N_5676,N_5120);
nand U7907 (N_7907,N_5315,N_5115);
nand U7908 (N_7908,N_4186,N_4741);
nor U7909 (N_7909,N_5554,N_4877);
or U7910 (N_7910,N_4192,N_4575);
and U7911 (N_7911,N_5901,N_4218);
nand U7912 (N_7912,N_5480,N_5425);
nand U7913 (N_7913,N_4355,N_5348);
nor U7914 (N_7914,N_5655,N_4206);
or U7915 (N_7915,N_5832,N_5793);
or U7916 (N_7916,N_4673,N_4705);
xor U7917 (N_7917,N_5423,N_5645);
xor U7918 (N_7918,N_5863,N_4271);
nor U7919 (N_7919,N_4795,N_5070);
xor U7920 (N_7920,N_4960,N_4458);
nor U7921 (N_7921,N_5646,N_5524);
or U7922 (N_7922,N_4561,N_4294);
nand U7923 (N_7923,N_5453,N_4653);
xor U7924 (N_7924,N_4717,N_5074);
nand U7925 (N_7925,N_4332,N_5360);
or U7926 (N_7926,N_4756,N_5239);
nor U7927 (N_7927,N_4146,N_4987);
or U7928 (N_7928,N_5907,N_4357);
and U7929 (N_7929,N_5137,N_4878);
and U7930 (N_7930,N_4401,N_4580);
nor U7931 (N_7931,N_4693,N_4169);
and U7932 (N_7932,N_5387,N_5546);
nor U7933 (N_7933,N_5232,N_4979);
nor U7934 (N_7934,N_4040,N_5557);
nor U7935 (N_7935,N_4176,N_5564);
nor U7936 (N_7936,N_4399,N_4395);
and U7937 (N_7937,N_5927,N_5046);
nor U7938 (N_7938,N_5986,N_5793);
nand U7939 (N_7939,N_4268,N_5360);
nor U7940 (N_7940,N_4053,N_5673);
and U7941 (N_7941,N_5963,N_4141);
xnor U7942 (N_7942,N_4095,N_4555);
xor U7943 (N_7943,N_4969,N_5913);
xnor U7944 (N_7944,N_4281,N_4421);
and U7945 (N_7945,N_5398,N_4895);
nand U7946 (N_7946,N_4229,N_4519);
nand U7947 (N_7947,N_5283,N_4761);
and U7948 (N_7948,N_5771,N_5822);
nand U7949 (N_7949,N_5870,N_5597);
nand U7950 (N_7950,N_4070,N_4137);
and U7951 (N_7951,N_4109,N_5106);
nand U7952 (N_7952,N_5694,N_4549);
nand U7953 (N_7953,N_4732,N_5302);
and U7954 (N_7954,N_5047,N_4181);
nand U7955 (N_7955,N_5435,N_4140);
and U7956 (N_7956,N_4169,N_4438);
or U7957 (N_7957,N_4629,N_4214);
and U7958 (N_7958,N_5769,N_5680);
and U7959 (N_7959,N_5424,N_5014);
or U7960 (N_7960,N_4844,N_5028);
nand U7961 (N_7961,N_4758,N_5167);
nand U7962 (N_7962,N_5884,N_4579);
and U7963 (N_7963,N_5938,N_5699);
nand U7964 (N_7964,N_5180,N_5664);
and U7965 (N_7965,N_5050,N_5017);
or U7966 (N_7966,N_4823,N_5043);
nor U7967 (N_7967,N_5685,N_5841);
and U7968 (N_7968,N_5864,N_4512);
nand U7969 (N_7969,N_4815,N_4551);
nand U7970 (N_7970,N_5314,N_4941);
or U7971 (N_7971,N_5596,N_5613);
and U7972 (N_7972,N_4481,N_4680);
and U7973 (N_7973,N_4933,N_5847);
and U7974 (N_7974,N_4783,N_4959);
nand U7975 (N_7975,N_4896,N_5964);
or U7976 (N_7976,N_4009,N_4886);
nor U7977 (N_7977,N_5048,N_5133);
and U7978 (N_7978,N_4220,N_4817);
and U7979 (N_7979,N_5793,N_4965);
xor U7980 (N_7980,N_4330,N_4756);
xnor U7981 (N_7981,N_4801,N_5531);
nor U7982 (N_7982,N_4549,N_5098);
nor U7983 (N_7983,N_4010,N_4308);
xnor U7984 (N_7984,N_4763,N_5076);
nand U7985 (N_7985,N_4739,N_4337);
and U7986 (N_7986,N_4977,N_5751);
nand U7987 (N_7987,N_5397,N_4633);
or U7988 (N_7988,N_5413,N_5271);
nand U7989 (N_7989,N_4290,N_5137);
nor U7990 (N_7990,N_4726,N_5747);
or U7991 (N_7991,N_5380,N_4285);
or U7992 (N_7992,N_5168,N_5060);
or U7993 (N_7993,N_5283,N_5750);
nor U7994 (N_7994,N_5101,N_4856);
and U7995 (N_7995,N_4804,N_4966);
xnor U7996 (N_7996,N_5162,N_5011);
or U7997 (N_7997,N_4521,N_5639);
nand U7998 (N_7998,N_4706,N_4588);
nor U7999 (N_7999,N_5956,N_4493);
nand U8000 (N_8000,N_6574,N_7434);
nor U8001 (N_8001,N_7637,N_7499);
and U8002 (N_8002,N_6261,N_6803);
xor U8003 (N_8003,N_6867,N_6071);
nor U8004 (N_8004,N_7986,N_7985);
and U8005 (N_8005,N_6094,N_7925);
or U8006 (N_8006,N_6570,N_7507);
nor U8007 (N_8007,N_7948,N_6181);
and U8008 (N_8008,N_6338,N_6645);
or U8009 (N_8009,N_7278,N_7223);
and U8010 (N_8010,N_6909,N_7182);
nor U8011 (N_8011,N_7658,N_7381);
nor U8012 (N_8012,N_7805,N_7685);
or U8013 (N_8013,N_7515,N_6706);
nand U8014 (N_8014,N_7933,N_6063);
or U8015 (N_8015,N_7075,N_7043);
nand U8016 (N_8016,N_7768,N_7409);
or U8017 (N_8017,N_6337,N_6179);
and U8018 (N_8018,N_7326,N_6908);
xor U8019 (N_8019,N_7599,N_7821);
or U8020 (N_8020,N_6992,N_7188);
nor U8021 (N_8021,N_6786,N_6457);
and U8022 (N_8022,N_7494,N_7401);
xor U8023 (N_8023,N_7708,N_7078);
nor U8024 (N_8024,N_7934,N_7905);
nor U8025 (N_8025,N_6498,N_7876);
nor U8026 (N_8026,N_7254,N_6150);
xor U8027 (N_8027,N_7879,N_7063);
and U8028 (N_8028,N_6630,N_7784);
and U8029 (N_8029,N_7842,N_7760);
or U8030 (N_8030,N_7815,N_7110);
or U8031 (N_8031,N_6636,N_7462);
nor U8032 (N_8032,N_6906,N_6823);
nor U8033 (N_8033,N_7915,N_7414);
nor U8034 (N_8034,N_6465,N_7102);
xor U8035 (N_8035,N_7984,N_7606);
xor U8036 (N_8036,N_6349,N_7686);
nand U8037 (N_8037,N_6155,N_7283);
or U8038 (N_8038,N_6217,N_7529);
nor U8039 (N_8039,N_6342,N_7631);
xor U8040 (N_8040,N_6006,N_6784);
nand U8041 (N_8041,N_7077,N_6933);
or U8042 (N_8042,N_6527,N_6348);
nor U8043 (N_8043,N_6715,N_7846);
and U8044 (N_8044,N_6259,N_6252);
or U8045 (N_8045,N_6792,N_6731);
nand U8046 (N_8046,N_6931,N_6542);
and U8047 (N_8047,N_6627,N_7580);
nor U8048 (N_8048,N_7410,N_6843);
and U8049 (N_8049,N_7699,N_7474);
nor U8050 (N_8050,N_7547,N_7539);
xnor U8051 (N_8051,N_6104,N_6969);
nand U8052 (N_8052,N_6318,N_7528);
and U8053 (N_8053,N_6932,N_6363);
nand U8054 (N_8054,N_6147,N_7097);
nand U8055 (N_8055,N_7333,N_6173);
or U8056 (N_8056,N_7183,N_7875);
nor U8057 (N_8057,N_7305,N_7327);
nand U8058 (N_8058,N_7368,N_7093);
nand U8059 (N_8059,N_7928,N_6226);
or U8060 (N_8060,N_6799,N_7313);
nor U8061 (N_8061,N_7859,N_7137);
xnor U8062 (N_8062,N_7593,N_6670);
nor U8063 (N_8063,N_7092,N_6689);
nand U8064 (N_8064,N_6501,N_6255);
nor U8065 (N_8065,N_7769,N_7651);
or U8066 (N_8066,N_6431,N_6978);
or U8067 (N_8067,N_7282,N_7908);
and U8068 (N_8068,N_6667,N_6145);
and U8069 (N_8069,N_6531,N_6166);
and U8070 (N_8070,N_6011,N_7475);
or U8071 (N_8071,N_6873,N_6671);
nor U8072 (N_8072,N_7892,N_7731);
nor U8073 (N_8073,N_6285,N_6118);
and U8074 (N_8074,N_7989,N_6437);
xnor U8075 (N_8075,N_7839,N_6276);
nor U8076 (N_8076,N_6354,N_6578);
and U8077 (N_8077,N_6123,N_6874);
and U8078 (N_8078,N_6185,N_6036);
nor U8079 (N_8079,N_6772,N_6162);
nor U8080 (N_8080,N_6002,N_6545);
and U8081 (N_8081,N_6499,N_7981);
or U8082 (N_8082,N_6129,N_6880);
and U8083 (N_8083,N_7049,N_6759);
nor U8084 (N_8084,N_6918,N_7490);
nand U8085 (N_8085,N_6331,N_6223);
and U8086 (N_8086,N_7729,N_6826);
nand U8087 (N_8087,N_6983,N_6827);
nor U8088 (N_8088,N_7689,N_7671);
nand U8089 (N_8089,N_6870,N_6359);
nand U8090 (N_8090,N_6642,N_7639);
nand U8091 (N_8091,N_7486,N_7952);
and U8092 (N_8092,N_6098,N_7324);
and U8093 (N_8093,N_6045,N_7429);
and U8094 (N_8094,N_6481,N_7527);
or U8095 (N_8095,N_6825,N_7123);
and U8096 (N_8096,N_6060,N_7229);
nor U8097 (N_8097,N_6709,N_6495);
xor U8098 (N_8098,N_7592,N_6494);
nor U8099 (N_8099,N_7430,N_6790);
or U8100 (N_8100,N_7248,N_7939);
and U8101 (N_8101,N_6973,N_6568);
nor U8102 (N_8102,N_7992,N_6262);
and U8103 (N_8103,N_7969,N_7317);
nand U8104 (N_8104,N_7762,N_7907);
and U8105 (N_8105,N_6442,N_6083);
xor U8106 (N_8106,N_6010,N_7961);
nand U8107 (N_8107,N_6284,N_6921);
nand U8108 (N_8108,N_6780,N_7346);
or U8109 (N_8109,N_7491,N_7041);
nand U8110 (N_8110,N_7433,N_7405);
nor U8111 (N_8111,N_7321,N_7504);
nand U8112 (N_8112,N_7163,N_7696);
nor U8113 (N_8113,N_7756,N_6444);
and U8114 (N_8114,N_7046,N_6315);
nor U8115 (N_8115,N_6916,N_6950);
nand U8116 (N_8116,N_6037,N_7392);
and U8117 (N_8117,N_6387,N_6143);
nor U8118 (N_8118,N_6369,N_7958);
nand U8119 (N_8119,N_6174,N_6206);
nand U8120 (N_8120,N_6726,N_7463);
nor U8121 (N_8121,N_6583,N_6378);
xor U8122 (N_8122,N_6801,N_6456);
nor U8123 (N_8123,N_6151,N_7067);
nand U8124 (N_8124,N_6633,N_6725);
or U8125 (N_8125,N_6681,N_7827);
xnor U8126 (N_8126,N_7465,N_6468);
nand U8127 (N_8127,N_7603,N_7295);
nand U8128 (N_8128,N_7752,N_6915);
nand U8129 (N_8129,N_7168,N_7705);
nand U8130 (N_8130,N_7664,N_7425);
nand U8131 (N_8131,N_6469,N_7226);
nor U8132 (N_8132,N_6240,N_7408);
nand U8133 (N_8133,N_6316,N_7798);
nor U8134 (N_8134,N_7776,N_6798);
nand U8135 (N_8135,N_6159,N_6941);
nand U8136 (N_8136,N_7822,N_7974);
nor U8137 (N_8137,N_7881,N_6040);
nor U8138 (N_8138,N_6686,N_7199);
or U8139 (N_8139,N_7079,N_7899);
nor U8140 (N_8140,N_6652,N_6530);
or U8141 (N_8141,N_6447,N_6735);
and U8142 (N_8142,N_7354,N_7398);
nand U8143 (N_8143,N_6515,N_6575);
nor U8144 (N_8144,N_6998,N_7745);
or U8145 (N_8145,N_7786,N_7143);
nor U8146 (N_8146,N_7763,N_6942);
nand U8147 (N_8147,N_6410,N_6334);
nor U8148 (N_8148,N_7116,N_6487);
nand U8149 (N_8149,N_7918,N_7645);
and U8150 (N_8150,N_7623,N_6220);
or U8151 (N_8151,N_6956,N_6329);
and U8152 (N_8152,N_7190,N_6379);
or U8153 (N_8153,N_6019,N_6899);
nor U8154 (N_8154,N_7205,N_7774);
xnor U8155 (N_8155,N_6260,N_7739);
nor U8156 (N_8156,N_6736,N_6120);
nand U8157 (N_8157,N_7121,N_6535);
and U8158 (N_8158,N_6061,N_6991);
nor U8159 (N_8159,N_7109,N_6388);
and U8160 (N_8160,N_6813,N_7903);
xor U8161 (N_8161,N_6312,N_7878);
nor U8162 (N_8162,N_7980,N_7251);
or U8163 (N_8163,N_6757,N_6866);
or U8164 (N_8164,N_6072,N_6520);
or U8165 (N_8165,N_6054,N_6018);
nand U8166 (N_8166,N_7877,N_7949);
nor U8167 (N_8167,N_7314,N_6326);
nor U8168 (N_8168,N_6987,N_7454);
or U8169 (N_8169,N_7341,N_7608);
nand U8170 (N_8170,N_7342,N_6139);
nor U8171 (N_8171,N_7135,N_7418);
xor U8172 (N_8172,N_7819,N_6835);
nand U8173 (N_8173,N_7450,N_7098);
nor U8174 (N_8174,N_7707,N_6131);
nor U8175 (N_8175,N_6043,N_7029);
nor U8176 (N_8176,N_7550,N_6272);
xnor U8177 (N_8177,N_7158,N_6382);
xnor U8178 (N_8178,N_6021,N_6113);
xnor U8179 (N_8179,N_6615,N_6576);
and U8180 (N_8180,N_6293,N_7087);
nor U8181 (N_8181,N_6848,N_6443);
and U8182 (N_8182,N_6197,N_7161);
and U8183 (N_8183,N_7460,N_7582);
nand U8184 (N_8184,N_7909,N_7924);
nor U8185 (N_8185,N_7035,N_6721);
and U8186 (N_8186,N_7432,N_7001);
nand U8187 (N_8187,N_7021,N_6056);
nand U8188 (N_8188,N_6218,N_6455);
nor U8189 (N_8189,N_6544,N_7204);
and U8190 (N_8190,N_6984,N_6788);
nand U8191 (N_8191,N_7120,N_7579);
nand U8192 (N_8192,N_7801,N_6925);
or U8193 (N_8193,N_6821,N_6092);
nand U8194 (N_8194,N_6279,N_6816);
nor U8195 (N_8195,N_7072,N_6288);
nor U8196 (N_8196,N_6264,N_7818);
and U8197 (N_8197,N_6560,N_7793);
xnor U8198 (N_8198,N_7853,N_7820);
nand U8199 (N_8199,N_6614,N_7173);
nor U8200 (N_8200,N_7096,N_6834);
nand U8201 (N_8201,N_6748,N_6394);
nor U8202 (N_8202,N_7562,N_6112);
nand U8203 (N_8203,N_6026,N_6882);
and U8204 (N_8204,N_6624,N_7510);
and U8205 (N_8205,N_6967,N_7068);
and U8206 (N_8206,N_6281,N_6532);
nand U8207 (N_8207,N_6851,N_6764);
and U8208 (N_8208,N_7322,N_7792);
nand U8209 (N_8209,N_7483,N_6879);
and U8210 (N_8210,N_7307,N_7139);
nand U8211 (N_8211,N_7581,N_6253);
nor U8212 (N_8212,N_7535,N_6791);
nand U8213 (N_8213,N_7480,N_6558);
and U8214 (N_8214,N_7570,N_6710);
nor U8215 (N_8215,N_6283,N_6646);
nand U8216 (N_8216,N_6345,N_7390);
xnor U8217 (N_8217,N_7607,N_6339);
nor U8218 (N_8218,N_7070,N_6859);
nor U8219 (N_8219,N_7447,N_6787);
nor U8220 (N_8220,N_6199,N_7247);
or U8221 (N_8221,N_7219,N_7703);
or U8222 (N_8222,N_7332,N_6015);
xnor U8223 (N_8223,N_6336,N_7840);
nand U8224 (N_8224,N_6588,N_7832);
and U8225 (N_8225,N_6023,N_7807);
nand U8226 (N_8226,N_6695,N_7904);
xnor U8227 (N_8227,N_7850,N_6745);
nand U8228 (N_8228,N_6108,N_7286);
or U8229 (N_8229,N_6486,N_7329);
nand U8230 (N_8230,N_6832,N_6522);
and U8231 (N_8231,N_7764,N_7973);
nand U8232 (N_8232,N_7265,N_6412);
nand U8233 (N_8233,N_6244,N_7289);
nand U8234 (N_8234,N_7222,N_6358);
and U8235 (N_8235,N_7027,N_7373);
or U8236 (N_8236,N_6599,N_7602);
nor U8237 (N_8237,N_6282,N_7383);
or U8238 (N_8238,N_7757,N_7681);
and U8239 (N_8239,N_6540,N_7466);
nor U8240 (N_8240,N_6078,N_6467);
or U8241 (N_8241,N_6739,N_7566);
or U8242 (N_8242,N_7207,N_7770);
xor U8243 (N_8243,N_6756,N_7153);
or U8244 (N_8244,N_6402,N_6032);
and U8245 (N_8245,N_7650,N_6067);
nor U8246 (N_8246,N_7202,N_6367);
and U8247 (N_8247,N_7310,N_6176);
and U8248 (N_8248,N_6038,N_6528);
xor U8249 (N_8249,N_6537,N_7013);
nor U8250 (N_8250,N_6724,N_7540);
nand U8251 (N_8251,N_7759,N_7748);
nand U8252 (N_8252,N_6595,N_7249);
nor U8253 (N_8253,N_7052,N_6556);
or U8254 (N_8254,N_6210,N_6153);
or U8255 (N_8255,N_6610,N_7175);
nand U8256 (N_8256,N_7628,N_7040);
and U8257 (N_8257,N_7937,N_7885);
nor U8258 (N_8258,N_6117,N_7356);
nand U8259 (N_8259,N_6413,N_7585);
nand U8260 (N_8260,N_7834,N_7979);
nand U8261 (N_8261,N_7099,N_6551);
nand U8262 (N_8262,N_6256,N_7297);
or U8263 (N_8263,N_6579,N_6052);
nand U8264 (N_8264,N_6003,N_6135);
and U8265 (N_8265,N_6783,N_7017);
or U8266 (N_8266,N_6035,N_6507);
nand U8267 (N_8267,N_6985,N_7843);
nor U8268 (N_8268,N_7308,N_6563);
or U8269 (N_8269,N_7053,N_7210);
nor U8270 (N_8270,N_6732,N_7836);
or U8271 (N_8271,N_7670,N_7825);
and U8272 (N_8272,N_6273,N_6140);
or U8273 (N_8273,N_6994,N_7988);
and U8274 (N_8274,N_7388,N_7635);
xnor U8275 (N_8275,N_7896,N_6789);
nand U8276 (N_8276,N_6049,N_7235);
or U8277 (N_8277,N_6124,N_7349);
or U8278 (N_8278,N_7054,N_7448);
or U8279 (N_8279,N_7868,N_6592);
nand U8280 (N_8280,N_7932,N_6656);
and U8281 (N_8281,N_7091,N_6510);
nor U8282 (N_8282,N_7133,N_7498);
nor U8283 (N_8283,N_6707,N_7468);
nor U8284 (N_8284,N_6611,N_7537);
nor U8285 (N_8285,N_7245,N_7415);
nor U8286 (N_8286,N_7794,N_7997);
and U8287 (N_8287,N_6426,N_7830);
and U8288 (N_8288,N_7755,N_7618);
and U8289 (N_8289,N_7028,N_7166);
and U8290 (N_8290,N_6418,N_6133);
nand U8291 (N_8291,N_6621,N_7085);
nand U8292 (N_8292,N_7370,N_6698);
xor U8293 (N_8293,N_7233,N_6893);
xnor U8294 (N_8294,N_7750,N_6436);
nand U8295 (N_8295,N_6251,N_7567);
or U8296 (N_8296,N_6355,N_7221);
nor U8297 (N_8297,N_7086,N_6694);
nor U8298 (N_8298,N_6257,N_6662);
and U8299 (N_8299,N_7338,N_7646);
and U8300 (N_8300,N_7488,N_7995);
nor U8301 (N_8301,N_7795,N_7838);
and U8302 (N_8302,N_6869,N_6910);
nand U8303 (N_8303,N_6650,N_6152);
or U8304 (N_8304,N_6314,N_7348);
or U8305 (N_8305,N_7037,N_6511);
nor U8306 (N_8306,N_7647,N_7831);
nand U8307 (N_8307,N_7501,N_6000);
and U8308 (N_8308,N_6683,N_7723);
xnor U8309 (N_8309,N_7604,N_6168);
nand U8310 (N_8310,N_6782,N_6594);
xor U8311 (N_8311,N_7747,N_7472);
nand U8312 (N_8312,N_7350,N_6659);
nand U8313 (N_8313,N_6237,N_6182);
and U8314 (N_8314,N_6684,N_6400);
nor U8315 (N_8315,N_6505,N_7142);
or U8316 (N_8316,N_6458,N_7309);
nor U8317 (N_8317,N_7880,N_7564);
nor U8318 (N_8318,N_6802,N_7125);
or U8319 (N_8319,N_6543,N_7452);
xor U8320 (N_8320,N_6366,N_7960);
or U8321 (N_8321,N_7165,N_6970);
and U8322 (N_8322,N_7039,N_7513);
and U8323 (N_8323,N_7653,N_7374);
or U8324 (N_8324,N_7789,N_7379);
nand U8325 (N_8325,N_7659,N_6863);
or U8326 (N_8326,N_7673,N_7187);
nand U8327 (N_8327,N_6857,N_7516);
xor U8328 (N_8328,N_7424,N_6972);
nand U8329 (N_8329,N_7471,N_7629);
or U8330 (N_8330,N_7935,N_6548);
nand U8331 (N_8331,N_6785,N_7551);
or U8332 (N_8332,N_6267,N_7002);
nor U8333 (N_8333,N_7443,N_6435);
and U8334 (N_8334,N_7999,N_6188);
and U8335 (N_8335,N_7023,N_6278);
and U8336 (N_8336,N_6503,N_6676);
or U8337 (N_8337,N_6343,N_6763);
nand U8338 (N_8338,N_6346,N_6902);
nand U8339 (N_8339,N_6471,N_6373);
nand U8340 (N_8340,N_7484,N_7697);
or U8341 (N_8341,N_7622,N_7787);
xnor U8342 (N_8342,N_6311,N_7519);
nor U8343 (N_8343,N_7375,N_7508);
xnor U8344 (N_8344,N_6327,N_6126);
nand U8345 (N_8345,N_7193,N_6042);
and U8346 (N_8346,N_7813,N_6473);
and U8347 (N_8347,N_7680,N_7082);
and U8348 (N_8348,N_6708,N_7612);
or U8349 (N_8349,N_6878,N_6623);
and U8350 (N_8350,N_6330,N_7791);
or U8351 (N_8351,N_7365,N_7923);
and U8352 (N_8352,N_6768,N_6463);
nand U8353 (N_8353,N_6231,N_7359);
and U8354 (N_8354,N_6172,N_6093);
and U8355 (N_8355,N_7117,N_7197);
and U8356 (N_8356,N_6765,N_7531);
xnor U8357 (N_8357,N_6233,N_6470);
nand U8358 (N_8358,N_7189,N_6989);
and U8359 (N_8359,N_6572,N_6945);
nand U8360 (N_8360,N_7674,N_6302);
nor U8361 (N_8361,N_6090,N_6858);
or U8362 (N_8362,N_6597,N_6952);
nor U8363 (N_8363,N_7011,N_7276);
or U8364 (N_8364,N_6215,N_7284);
nor U8365 (N_8365,N_7159,N_6957);
nor U8366 (N_8366,N_7944,N_6509);
xnor U8367 (N_8367,N_6479,N_6490);
or U8368 (N_8368,N_7571,N_7030);
and U8369 (N_8369,N_7240,N_6525);
or U8370 (N_8370,N_6690,N_6059);
nand U8371 (N_8371,N_7778,N_7845);
nor U8372 (N_8372,N_6640,N_7104);
or U8373 (N_8373,N_7352,N_6831);
nand U8374 (N_8374,N_6986,N_7965);
xnor U8375 (N_8375,N_6350,N_6344);
and U8376 (N_8376,N_7503,N_7682);
nand U8377 (N_8377,N_6777,N_6612);
nor U8378 (N_8378,N_6077,N_7266);
xnor U8379 (N_8379,N_6022,N_6491);
nor U8380 (N_8380,N_7917,N_7181);
or U8381 (N_8381,N_6300,N_6716);
or U8382 (N_8382,N_6850,N_7530);
or U8383 (N_8383,N_7594,N_6274);
and U8384 (N_8384,N_6796,N_6904);
nand U8385 (N_8385,N_6234,N_7019);
and U8386 (N_8386,N_7678,N_7237);
or U8387 (N_8387,N_6533,N_6075);
or U8388 (N_8388,N_6618,N_7521);
xor U8389 (N_8389,N_7672,N_6876);
nand U8390 (N_8390,N_7520,N_7626);
xnor U8391 (N_8391,N_7257,N_7084);
nor U8392 (N_8392,N_6017,N_7162);
xor U8393 (N_8393,N_6103,N_6306);
and U8394 (N_8394,N_7852,N_6247);
or U8395 (N_8395,N_6753,N_6929);
nand U8396 (N_8396,N_6622,N_6031);
nand U8397 (N_8397,N_7217,N_6585);
nor U8398 (N_8398,N_7496,N_6085);
nor U8399 (N_8399,N_6347,N_7945);
and U8400 (N_8400,N_6928,N_7476);
and U8401 (N_8401,N_7377,N_6406);
nand U8402 (N_8402,N_6089,N_6304);
or U8403 (N_8403,N_6613,N_7236);
and U8404 (N_8404,N_7611,N_7882);
or U8405 (N_8405,N_7929,N_6743);
and U8406 (N_8406,N_7200,N_6087);
nor U8407 (N_8407,N_6044,N_7620);
nand U8408 (N_8408,N_7887,N_6028);
or U8409 (N_8409,N_6500,N_6325);
nand U8410 (N_8410,N_7000,N_6958);
nand U8411 (N_8411,N_7625,N_6452);
and U8412 (N_8412,N_7584,N_7677);
and U8413 (N_8413,N_7344,N_7886);
xnor U8414 (N_8414,N_7347,N_6156);
or U8415 (N_8415,N_7242,N_6555);
nor U8416 (N_8416,N_6137,N_7300);
or U8417 (N_8417,N_6489,N_7721);
xor U8418 (N_8418,N_7244,N_6718);
and U8419 (N_8419,N_7492,N_7898);
nand U8420 (N_8420,N_6440,N_7642);
nand U8421 (N_8421,N_7728,N_7268);
nand U8422 (N_8422,N_6308,N_6534);
nor U8423 (N_8423,N_7652,N_7991);
and U8424 (N_8424,N_6474,N_7185);
nor U8425 (N_8425,N_7404,N_6229);
xor U8426 (N_8426,N_7090,N_7074);
or U8427 (N_8427,N_6566,N_7569);
xnor U8428 (N_8428,N_6324,N_7306);
or U8429 (N_8429,N_7275,N_7252);
nor U8430 (N_8430,N_6111,N_7155);
and U8431 (N_8431,N_7319,N_6573);
nor U8432 (N_8432,N_7088,N_7239);
and U8433 (N_8433,N_6186,N_6012);
and U8434 (N_8434,N_7218,N_6472);
or U8435 (N_8435,N_6496,N_7279);
or U8436 (N_8436,N_6896,N_7195);
nor U8437 (N_8437,N_7018,N_6964);
and U8438 (N_8438,N_6202,N_7045);
nand U8439 (N_8439,N_7411,N_7130);
xor U8440 (N_8440,N_7412,N_6008);
nand U8441 (N_8441,N_7753,N_6169);
nand U8442 (N_8442,N_6464,N_6951);
nand U8443 (N_8443,N_7495,N_7869);
nor U8444 (N_8444,N_7525,N_7089);
nand U8445 (N_8445,N_6034,N_6020);
nor U8446 (N_8446,N_7542,N_6136);
or U8447 (N_8447,N_7361,N_6371);
xor U8448 (N_8448,N_6432,N_7926);
and U8449 (N_8449,N_6328,N_6996);
or U8450 (N_8450,N_7613,N_6305);
or U8451 (N_8451,N_7816,N_7693);
nand U8452 (N_8452,N_7914,N_7005);
nand U8453 (N_8453,N_6122,N_6461);
xor U8454 (N_8454,N_6920,N_6871);
nand U8455 (N_8455,N_6191,N_6886);
and U8456 (N_8456,N_7698,N_7396);
or U8457 (N_8457,N_6250,N_6062);
nor U8458 (N_8458,N_7394,N_7777);
nand U8459 (N_8459,N_6762,N_6923);
and U8460 (N_8460,N_6198,N_6717);
nor U8461 (N_8461,N_6949,N_6287);
or U8462 (N_8462,N_6408,N_6521);
and U8463 (N_8463,N_6712,N_7294);
and U8464 (N_8464,N_6187,N_6905);
and U8465 (N_8465,N_7191,N_7506);
nand U8466 (N_8466,N_6541,N_6064);
nand U8467 (N_8467,N_6091,N_7006);
nand U8468 (N_8468,N_7993,N_6911);
nor U8469 (N_8469,N_7717,N_6438);
xor U8470 (N_8470,N_6794,N_7883);
and U8471 (N_8471,N_7641,N_7262);
and U8472 (N_8472,N_6211,N_6066);
and U8473 (N_8473,N_6881,N_7605);
nor U8474 (N_8474,N_7927,N_7632);
or U8475 (N_8475,N_6492,N_6653);
and U8476 (N_8476,N_7470,N_6506);
nand U8477 (N_8477,N_7738,N_6723);
nor U8478 (N_8478,N_6514,N_7453);
nor U8479 (N_8479,N_7982,N_7290);
and U8480 (N_8480,N_7873,N_7800);
and U8481 (N_8481,N_6362,N_6885);
or U8482 (N_8482,N_6760,N_7334);
nand U8483 (N_8483,N_6852,N_7048);
nor U8484 (N_8484,N_6552,N_7194);
or U8485 (N_8485,N_7676,N_6007);
nand U8486 (N_8486,N_6502,N_6232);
nor U8487 (N_8487,N_7780,N_6701);
or U8488 (N_8488,N_7154,N_6175);
nor U8489 (N_8489,N_6720,N_7395);
nand U8490 (N_8490,N_7292,N_7062);
nor U8491 (N_8491,N_6517,N_6476);
or U8492 (N_8492,N_6795,N_7720);
and U8493 (N_8493,N_6478,N_7725);
or U8494 (N_8494,N_6214,N_7482);
nor U8495 (N_8495,N_7802,N_6254);
nor U8496 (N_8496,N_7775,N_7277);
or U8497 (N_8497,N_7779,N_7847);
and U8498 (N_8498,N_6897,N_7380);
nand U8499 (N_8499,N_6849,N_6569);
and U8500 (N_8500,N_6102,N_7094);
or U8501 (N_8501,N_6699,N_7323);
or U8502 (N_8502,N_7083,N_6603);
xnor U8503 (N_8503,N_7114,N_6641);
nand U8504 (N_8504,N_6245,N_6046);
and U8505 (N_8505,N_7812,N_6892);
or U8506 (N_8506,N_7066,N_6230);
nand U8507 (N_8507,N_6353,N_6901);
nor U8508 (N_8508,N_6752,N_7666);
nand U8509 (N_8509,N_7862,N_6526);
nor U8510 (N_8510,N_6665,N_6411);
nor U8511 (N_8511,N_6451,N_7823);
nor U8512 (N_8512,N_7920,N_7473);
nor U8513 (N_8513,N_7568,N_6294);
or U8514 (N_8514,N_6968,N_6033);
nor U8515 (N_8515,N_7058,N_6536);
or U8516 (N_8516,N_7112,N_6811);
nor U8517 (N_8517,N_6405,N_7552);
or U8518 (N_8518,N_7848,N_7724);
nand U8519 (N_8519,N_7339,N_6146);
nand U8520 (N_8520,N_7440,N_6655);
nor U8521 (N_8521,N_7867,N_6894);
and U8522 (N_8522,N_7601,N_7170);
and U8523 (N_8523,N_6856,N_7711);
or U8524 (N_8524,N_7238,N_6271);
or U8525 (N_8525,N_7014,N_6940);
xor U8526 (N_8526,N_7435,N_6030);
nand U8527 (N_8527,N_6557,N_6212);
xnor U8528 (N_8528,N_7954,N_6982);
or U8529 (N_8529,N_6360,N_7164);
and U8530 (N_8530,N_6620,N_7272);
nand U8531 (N_8531,N_7174,N_6291);
or U8532 (N_8532,N_6519,N_6380);
nand U8533 (N_8533,N_6638,N_6914);
nor U8534 (N_8534,N_6883,N_6872);
nand U8535 (N_8535,N_7336,N_6127);
and U8536 (N_8536,N_6793,N_7716);
nor U8537 (N_8537,N_6403,N_6286);
and U8538 (N_8538,N_6778,N_7972);
nor U8539 (N_8539,N_6321,N_7841);
nor U8540 (N_8540,N_7071,N_7766);
nand U8541 (N_8541,N_7749,N_7095);
and U8542 (N_8542,N_6208,N_6948);
nor U8543 (N_8543,N_7132,N_6395);
or U8544 (N_8544,N_6453,N_6204);
and U8545 (N_8545,N_7754,N_7351);
nor U8546 (N_8546,N_7400,N_7541);
nand U8547 (N_8547,N_7107,N_7511);
nor U8548 (N_8548,N_7489,N_7576);
nor U8549 (N_8549,N_7493,N_7302);
nand U8550 (N_8550,N_6041,N_7971);
and U8551 (N_8551,N_7357,N_6577);
or U8552 (N_8552,N_7714,N_7597);
nor U8553 (N_8553,N_7888,N_6847);
or U8554 (N_8554,N_6677,N_6845);
or U8555 (N_8555,N_7146,N_6946);
nand U8556 (N_8556,N_7105,N_6356);
xnor U8557 (N_8557,N_6084,N_7243);
nor U8558 (N_8558,N_7872,N_6290);
nand U8559 (N_8559,N_6070,N_7718);
nor U8560 (N_8560,N_7128,N_7649);
and U8561 (N_8561,N_6074,N_6448);
nand U8562 (N_8562,N_7534,N_6390);
xnor U8563 (N_8563,N_6048,N_7061);
nor U8564 (N_8564,N_6483,N_6180);
or U8565 (N_8565,N_7627,N_6884);
nand U8566 (N_8566,N_6571,N_6109);
nor U8567 (N_8567,N_6009,N_6423);
and U8568 (N_8568,N_7555,N_7957);
xnor U8569 (N_8569,N_7367,N_7710);
nor U8570 (N_8570,N_7727,N_6589);
and U8571 (N_8571,N_6935,N_6959);
or U8572 (N_8572,N_6497,N_7285);
and U8573 (N_8573,N_7076,N_7771);
nor U8574 (N_8574,N_7421,N_7911);
nor U8575 (N_8575,N_7296,N_7171);
xor U8576 (N_8576,N_7340,N_7758);
nor U8577 (N_8577,N_6361,N_6297);
nor U8578 (N_8578,N_6351,N_6770);
xor U8579 (N_8579,N_6564,N_6961);
and U8580 (N_8580,N_7059,N_6606);
nor U8581 (N_8581,N_6565,N_6466);
nor U8582 (N_8582,N_6384,N_7108);
and U8583 (N_8583,N_6524,N_7860);
nand U8584 (N_8584,N_6738,N_7301);
nand U8585 (N_8585,N_6679,N_7811);
or U8586 (N_8586,N_6729,N_7316);
nor U8587 (N_8587,N_7732,N_7050);
and U8588 (N_8588,N_7938,N_7280);
nand U8589 (N_8589,N_6586,N_6680);
or U8590 (N_8590,N_6947,N_7797);
xnor U8591 (N_8591,N_6399,N_7514);
nand U8592 (N_8592,N_6263,N_6819);
nand U8593 (N_8593,N_6246,N_6974);
and U8594 (N_8594,N_7740,N_6106);
or U8595 (N_8595,N_7849,N_7976);
nand U8596 (N_8596,N_6320,N_7742);
or U8597 (N_8597,N_7364,N_6079);
or U8598 (N_8598,N_6449,N_7360);
nor U8599 (N_8599,N_7003,N_6392);
and U8600 (N_8600,N_6602,N_7149);
nand U8601 (N_8601,N_6421,N_7328);
nor U8602 (N_8602,N_7889,N_7669);
and U8603 (N_8603,N_6051,N_7312);
xor U8604 (N_8604,N_6898,N_7863);
nand U8605 (N_8605,N_7281,N_7457);
and U8606 (N_8606,N_7150,N_6868);
nand U8607 (N_8607,N_7808,N_7684);
xor U8608 (N_8608,N_6600,N_7804);
or U8609 (N_8609,N_7420,N_7687);
and U8610 (N_8610,N_6529,N_7782);
and U8611 (N_8611,N_7241,N_6841);
nor U8612 (N_8612,N_7902,N_7145);
and U8613 (N_8613,N_7180,N_7661);
and U8614 (N_8614,N_7919,N_6097);
or U8615 (N_8615,N_7624,N_7600);
nand U8616 (N_8616,N_7113,N_6682);
or U8617 (N_8617,N_6484,N_7656);
and U8618 (N_8618,N_7810,N_7975);
nor U8619 (N_8619,N_7436,N_6766);
nand U8620 (N_8620,N_7010,N_7943);
or U8621 (N_8621,N_7610,N_7695);
or U8622 (N_8622,N_6890,N_6073);
xor U8623 (N_8623,N_7100,N_6213);
or U8624 (N_8624,N_7055,N_6225);
nand U8625 (N_8625,N_7691,N_6236);
or U8626 (N_8626,N_7549,N_6134);
nand U8627 (N_8627,N_7022,N_6742);
nor U8628 (N_8628,N_7587,N_6962);
nor U8629 (N_8629,N_6057,N_7015);
xnor U8630 (N_8630,N_7232,N_6462);
xnor U8631 (N_8631,N_6165,N_7556);
or U8632 (N_8632,N_7131,N_6270);
or U8633 (N_8633,N_7391,N_7343);
nor U8634 (N_8634,N_6713,N_6854);
and U8635 (N_8635,N_7942,N_7269);
and U8636 (N_8636,N_6417,N_7331);
or U8637 (N_8637,N_7186,N_6660);
nor U8638 (N_8638,N_6995,N_6628);
or U8639 (N_8639,N_6685,N_6979);
or U8640 (N_8640,N_7455,N_7726);
or U8641 (N_8641,N_6875,N_6924);
nand U8642 (N_8642,N_6822,N_6157);
or U8643 (N_8643,N_7106,N_7209);
nor U8644 (N_8644,N_6446,N_6654);
nor U8645 (N_8645,N_6668,N_7212);
and U8646 (N_8646,N_7148,N_7406);
nor U8647 (N_8647,N_7366,N_7574);
and U8648 (N_8648,N_7246,N_6862);
and U8649 (N_8649,N_6280,N_6167);
xnor U8650 (N_8650,N_6383,N_6207);
nor U8651 (N_8651,N_6830,N_7184);
or U8652 (N_8652,N_7258,N_6887);
and U8653 (N_8653,N_7783,N_7543);
or U8654 (N_8654,N_7857,N_7505);
or U8655 (N_8655,N_6737,N_6058);
and U8656 (N_8656,N_6485,N_7213);
nor U8657 (N_8657,N_6357,N_6414);
nand U8658 (N_8658,N_6516,N_6553);
or U8659 (N_8659,N_7335,N_7835);
and U8660 (N_8660,N_7586,N_7304);
or U8661 (N_8661,N_7964,N_6714);
and U8662 (N_8662,N_6518,N_7073);
and U8663 (N_8663,N_6944,N_7057);
nand U8664 (N_8664,N_6222,N_7996);
xnor U8665 (N_8665,N_6809,N_6141);
xnor U8666 (N_8666,N_6550,N_6728);
nor U8667 (N_8667,N_6450,N_6249);
and U8668 (N_8668,N_7712,N_6697);
nor U8669 (N_8669,N_6733,N_6105);
nor U8670 (N_8670,N_7385,N_6661);
nor U8671 (N_8671,N_7419,N_6377);
or U8672 (N_8672,N_6195,N_7026);
xor U8673 (N_8673,N_7906,N_6971);
nand U8674 (N_8674,N_6663,N_6389);
xor U8675 (N_8675,N_6747,N_7273);
nand U8676 (N_8676,N_7318,N_6755);
nor U8677 (N_8677,N_6672,N_7038);
or U8678 (N_8678,N_7619,N_7417);
or U8679 (N_8679,N_7660,N_7416);
nor U8680 (N_8680,N_7561,N_6864);
and U8681 (N_8681,N_6333,N_6301);
xnor U8682 (N_8682,N_6598,N_6398);
and U8683 (N_8683,N_6903,N_6907);
xnor U8684 (N_8684,N_7871,N_6370);
xor U8685 (N_8685,N_6919,N_6076);
xnor U8686 (N_8686,N_7441,N_6319);
xnor U8687 (N_8687,N_7399,N_6607);
nor U8688 (N_8688,N_7824,N_7469);
nand U8689 (N_8689,N_7683,N_7376);
nand U8690 (N_8690,N_7634,N_6445);
or U8691 (N_8691,N_6427,N_6303);
and U8692 (N_8692,N_7256,N_7546);
or U8693 (N_8693,N_6673,N_6593);
nor U8694 (N_8694,N_7428,N_7734);
nor U8695 (N_8695,N_6425,N_6332);
and U8696 (N_8696,N_6258,N_7464);
and U8697 (N_8697,N_6554,N_6687);
and U8698 (N_8698,N_6797,N_6608);
and U8699 (N_8699,N_6016,N_6239);
nand U8700 (N_8700,N_7081,N_6913);
nand U8701 (N_8701,N_7178,N_7230);
nor U8702 (N_8702,N_6549,N_6295);
or U8703 (N_8703,N_7788,N_7829);
or U8704 (N_8704,N_6644,N_7544);
nand U8705 (N_8705,N_6634,N_6125);
nor U8706 (N_8706,N_7479,N_7378);
or U8707 (N_8707,N_7291,N_6298);
and U8708 (N_8708,N_7051,N_7451);
and U8709 (N_8709,N_7481,N_7227);
or U8710 (N_8710,N_7931,N_6808);
or U8711 (N_8711,N_6523,N_6025);
and U8712 (N_8712,N_7402,N_6095);
nor U8713 (N_8713,N_6053,N_7990);
or U8714 (N_8714,N_6853,N_6616);
and U8715 (N_8715,N_6990,N_7956);
or U8716 (N_8716,N_6088,N_6376);
or U8717 (N_8717,N_7438,N_6364);
or U8718 (N_8718,N_6508,N_7345);
xor U8719 (N_8719,N_6101,N_7355);
nand U8720 (N_8720,N_7557,N_7598);
and U8721 (N_8721,N_7456,N_7167);
nor U8722 (N_8722,N_6488,N_6538);
nor U8723 (N_8723,N_7577,N_7772);
xor U8724 (N_8724,N_6960,N_6704);
or U8725 (N_8725,N_7437,N_6119);
or U8726 (N_8726,N_7983,N_6861);
or U8727 (N_8727,N_7203,N_7069);
nand U8728 (N_8728,N_6454,N_7522);
or U8729 (N_8729,N_7129,N_6963);
nor U8730 (N_8730,N_7502,N_7809);
or U8731 (N_8731,N_6228,N_6480);
nand U8732 (N_8732,N_6374,N_6203);
nand U8733 (N_8733,N_6567,N_6648);
nor U8734 (N_8734,N_6895,N_7854);
nor U8735 (N_8735,N_6999,N_7930);
or U8736 (N_8736,N_6433,N_6754);
nand U8737 (N_8737,N_6401,N_7837);
nor U8738 (N_8738,N_6099,N_6219);
nor U8739 (N_8739,N_6773,N_7431);
nor U8740 (N_8740,N_6926,N_7103);
or U8741 (N_8741,N_6705,N_7220);
xnor U8742 (N_8742,N_7477,N_6817);
or U8743 (N_8743,N_7111,N_6004);
or U8744 (N_8744,N_7751,N_7311);
nand U8745 (N_8745,N_7234,N_6647);
nand U8746 (N_8746,N_7042,N_7337);
xnor U8747 (N_8747,N_7959,N_7016);
or U8748 (N_8748,N_6422,N_7371);
nor U8749 (N_8749,N_6241,N_7261);
nand U8750 (N_8750,N_6649,N_7950);
nor U8751 (N_8751,N_7864,N_7389);
nor U8752 (N_8752,N_6068,N_6368);
xor U8753 (N_8753,N_7897,N_6238);
and U8754 (N_8754,N_6065,N_6980);
xor U8755 (N_8755,N_6163,N_6619);
and U8756 (N_8756,N_7743,N_6144);
or U8757 (N_8757,N_7702,N_6820);
nand U8758 (N_8758,N_7138,N_7500);
or U8759 (N_8759,N_7449,N_7955);
and U8760 (N_8760,N_7147,N_7201);
nor U8761 (N_8761,N_6815,N_6183);
nor U8762 (N_8762,N_6375,N_7215);
and U8763 (N_8763,N_7706,N_6242);
and U8764 (N_8764,N_6936,N_6116);
nand U8765 (N_8765,N_6584,N_7701);
nor U8766 (N_8766,N_7912,N_7397);
and U8767 (N_8767,N_7179,N_7730);
or U8768 (N_8768,N_6658,N_6029);
nor U8769 (N_8769,N_7828,N_6993);
and U8770 (N_8770,N_6080,N_6703);
xor U8771 (N_8771,N_7894,N_7523);
nor U8772 (N_8772,N_7968,N_6289);
nand U8773 (N_8773,N_7047,N_6744);
nor U8774 (N_8774,N_6415,N_7330);
or U8775 (N_8775,N_7575,N_6939);
and U8776 (N_8776,N_7036,N_6419);
nor U8777 (N_8777,N_6248,N_6082);
or U8778 (N_8778,N_6130,N_7253);
nor U8779 (N_8779,N_7709,N_6877);
nand U8780 (N_8780,N_7636,N_7773);
and U8781 (N_8781,N_6024,N_7573);
nor U8782 (N_8782,N_6746,N_7690);
or U8783 (N_8783,N_6761,N_6741);
nor U8784 (N_8784,N_6055,N_6385);
xor U8785 (N_8785,N_7941,N_7386);
and U8786 (N_8786,N_7614,N_7994);
and U8787 (N_8787,N_7442,N_7152);
nor U8788 (N_8788,N_7861,N_7617);
nand U8789 (N_8789,N_7998,N_7444);
nor U8790 (N_8790,N_6775,N_6096);
or U8791 (N_8791,N_6702,N_7206);
and U8792 (N_8792,N_6424,N_7746);
and U8793 (N_8793,N_7590,N_6170);
and U8794 (N_8794,N_7298,N_6292);
nand U8795 (N_8795,N_7033,N_7169);
and U8796 (N_8796,N_7583,N_6562);
nor U8797 (N_8797,N_6275,N_6580);
xnor U8798 (N_8798,N_7719,N_6420);
nor U8799 (N_8799,N_6937,N_7891);
nand U8800 (N_8800,N_7497,N_6609);
and U8801 (N_8801,N_6148,N_7588);
xor U8802 (N_8802,N_6814,N_6475);
nor U8803 (N_8803,N_7536,N_6930);
and U8804 (N_8804,N_6027,N_7461);
nand U8805 (N_8805,N_6039,N_7101);
nor U8806 (N_8806,N_6981,N_6323);
nand U8807 (N_8807,N_6769,N_7288);
nand U8808 (N_8808,N_6193,N_7427);
and U8809 (N_8809,N_7910,N_7638);
nand U8810 (N_8810,N_7874,N_6734);
and U8811 (N_8811,N_7741,N_6459);
or U8812 (N_8812,N_6310,N_7407);
nand U8813 (N_8813,N_6265,N_6900);
xnor U8814 (N_8814,N_6397,N_7826);
and U8815 (N_8815,N_7478,N_6069);
nor U8816 (N_8816,N_7064,N_7198);
nor U8817 (N_8817,N_6121,N_6749);
or U8818 (N_8818,N_7817,N_6441);
and U8819 (N_8819,N_6190,N_7382);
and U8820 (N_8820,N_7532,N_6629);
nand U8821 (N_8821,N_7287,N_7426);
xnor U8822 (N_8822,N_6688,N_7216);
nor U8823 (N_8823,N_6632,N_6205);
and U8824 (N_8824,N_6781,N_7134);
nand U8825 (N_8825,N_6842,N_7124);
or U8826 (N_8826,N_7533,N_7267);
nor U8827 (N_8827,N_7458,N_6493);
and U8828 (N_8828,N_6269,N_7806);
nand U8829 (N_8829,N_6138,N_6977);
or U8830 (N_8830,N_7560,N_6428);
nand U8831 (N_8831,N_6340,N_7767);
nor U8832 (N_8832,N_7065,N_6975);
nand U8833 (N_8833,N_7034,N_7228);
or U8834 (N_8834,N_7591,N_7648);
or U8835 (N_8835,N_6386,N_6807);
and U8836 (N_8836,N_6806,N_6158);
nand U8837 (N_8837,N_6396,N_6604);
and U8838 (N_8838,N_6014,N_7260);
and U8839 (N_8839,N_6194,N_6966);
and U8840 (N_8840,N_7439,N_7722);
xor U8841 (N_8841,N_7796,N_7700);
nand U8842 (N_8842,N_6154,N_7032);
and U8843 (N_8843,N_7865,N_6513);
and U8844 (N_8844,N_6776,N_7866);
and U8845 (N_8845,N_6581,N_7855);
and U8846 (N_8846,N_6840,N_7122);
and U8847 (N_8847,N_7966,N_6322);
nand U8848 (N_8848,N_6674,N_6100);
nor U8849 (N_8849,N_6313,N_7487);
nand U8850 (N_8850,N_7485,N_6988);
nor U8851 (N_8851,N_6953,N_6635);
nand U8852 (N_8852,N_6976,N_6891);
or U8853 (N_8853,N_6812,N_7524);
and U8854 (N_8854,N_7231,N_7963);
or U8855 (N_8855,N_6184,N_7422);
nor U8856 (N_8856,N_6381,N_7553);
or U8857 (N_8857,N_6434,N_6546);
nand U8858 (N_8858,N_7446,N_7293);
and U8859 (N_8859,N_6013,N_7224);
and U8860 (N_8860,N_7978,N_7621);
or U8861 (N_8861,N_6482,N_7596);
and U8862 (N_8862,N_6299,N_6309);
or U8863 (N_8863,N_6818,N_7362);
nor U8864 (N_8864,N_7675,N_7136);
or U8865 (N_8865,N_6115,N_6429);
nor U8866 (N_8866,N_7665,N_7946);
nor U8867 (N_8867,N_6631,N_7141);
or U8868 (N_8868,N_7177,N_7208);
xnor U8869 (N_8869,N_6268,N_6625);
and U8870 (N_8870,N_6561,N_6504);
nand U8871 (N_8871,N_6722,N_7856);
or U8872 (N_8872,N_6439,N_7517);
nor U8873 (N_8873,N_6829,N_7578);
and U8874 (N_8874,N_6912,N_6954);
nand U8875 (N_8875,N_7255,N_7548);
or U8876 (N_8876,N_6675,N_6965);
or U8877 (N_8877,N_7140,N_6800);
nand U8878 (N_8878,N_7545,N_7657);
xor U8879 (N_8879,N_6142,N_7115);
or U8880 (N_8880,N_6601,N_6243);
nor U8881 (N_8881,N_7644,N_7056);
and U8882 (N_8882,N_7270,N_7951);
nor U8883 (N_8883,N_7118,N_7563);
nor U8884 (N_8884,N_7020,N_7160);
nor U8885 (N_8885,N_6833,N_7358);
or U8886 (N_8886,N_7372,N_7715);
nand U8887 (N_8887,N_7694,N_7844);
xor U8888 (N_8888,N_7953,N_7940);
and U8889 (N_8889,N_7643,N_7192);
nand U8890 (N_8890,N_7353,N_7080);
nand U8891 (N_8891,N_6001,N_7851);
nor U8892 (N_8892,N_7884,N_6643);
and U8893 (N_8893,N_6559,N_7060);
nor U8894 (N_8894,N_7833,N_6341);
and U8895 (N_8895,N_7692,N_6209);
nand U8896 (N_8896,N_7369,N_6774);
or U8897 (N_8897,N_7559,N_6477);
nor U8898 (N_8898,N_7467,N_7737);
nand U8899 (N_8899,N_7916,N_6596);
xor U8900 (N_8900,N_7922,N_7630);
and U8901 (N_8901,N_7913,N_7936);
nor U8902 (N_8902,N_7554,N_6178);
xnor U8903 (N_8903,N_6335,N_7538);
nand U8904 (N_8904,N_6352,N_6114);
nor U8905 (N_8905,N_7320,N_7662);
nor U8906 (N_8906,N_7509,N_7127);
and U8907 (N_8907,N_7393,N_6161);
nor U8908 (N_8908,N_7413,N_7790);
nor U8909 (N_8909,N_6086,N_6404);
or U8910 (N_8910,N_6810,N_7640);
nor U8911 (N_8911,N_6693,N_7947);
or U8912 (N_8912,N_6727,N_7176);
or U8913 (N_8913,N_6393,N_7572);
xor U8914 (N_8914,N_6221,N_6917);
nor U8915 (N_8915,N_7518,N_6692);
nand U8916 (N_8916,N_7615,N_6997);
xor U8917 (N_8917,N_7654,N_6587);
nor U8918 (N_8918,N_6617,N_6664);
or U8919 (N_8919,N_6865,N_6582);
nand U8920 (N_8920,N_6846,N_6460);
or U8921 (N_8921,N_6837,N_7012);
and U8922 (N_8922,N_7633,N_7044);
nor U8923 (N_8923,N_6224,N_7781);
nand U8924 (N_8924,N_6678,N_7259);
nand U8925 (N_8925,N_7870,N_6277);
nand U8926 (N_8926,N_7526,N_6669);
nand U8927 (N_8927,N_6651,N_6177);
and U8928 (N_8928,N_6637,N_7667);
or U8929 (N_8929,N_6047,N_7225);
and U8930 (N_8930,N_7299,N_7264);
nor U8931 (N_8931,N_7655,N_7901);
nor U8932 (N_8932,N_6266,N_6828);
or U8933 (N_8933,N_6767,N_6943);
and U8934 (N_8934,N_6771,N_6740);
and U8935 (N_8935,N_6200,N_7890);
nand U8936 (N_8936,N_6730,N_7387);
xnor U8937 (N_8937,N_6050,N_6171);
or U8938 (N_8938,N_6196,N_7156);
nand U8939 (N_8939,N_6888,N_6696);
nor U8940 (N_8940,N_7799,N_7007);
and U8941 (N_8941,N_7172,N_7403);
and U8942 (N_8942,N_7858,N_6409);
nor U8943 (N_8943,N_7423,N_6372);
and U8944 (N_8944,N_7679,N_7009);
nand U8945 (N_8945,N_7704,N_6132);
nor U8946 (N_8946,N_7895,N_6160);
nand U8947 (N_8947,N_7384,N_6081);
xor U8948 (N_8948,N_6430,N_7688);
nand U8949 (N_8949,N_7025,N_6889);
xnor U8950 (N_8950,N_7263,N_6149);
xor U8951 (N_8951,N_7445,N_7589);
nor U8952 (N_8952,N_6938,N_6751);
and U8953 (N_8953,N_7967,N_6591);
xnor U8954 (N_8954,N_6805,N_6539);
and U8955 (N_8955,N_7765,N_6128);
nand U8956 (N_8956,N_6750,N_7595);
or U8957 (N_8957,N_7250,N_7008);
nand U8958 (N_8958,N_7977,N_6804);
and U8959 (N_8959,N_6590,N_6416);
or U8960 (N_8960,N_7736,N_7211);
nor U8961 (N_8961,N_7609,N_7512);
and U8962 (N_8962,N_6657,N_7126);
xnor U8963 (N_8963,N_7893,N_6307);
and U8964 (N_8964,N_6407,N_7663);
nor U8965 (N_8965,N_7119,N_7803);
or U8966 (N_8966,N_6844,N_6824);
nor U8967 (N_8967,N_6927,N_7744);
nor U8968 (N_8968,N_7735,N_6639);
nand U8969 (N_8969,N_7962,N_7987);
nor U8970 (N_8970,N_6216,N_7031);
and U8971 (N_8971,N_6296,N_7814);
nor U8972 (N_8972,N_7144,N_6855);
nand U8973 (N_8973,N_7900,N_6860);
nand U8974 (N_8974,N_7004,N_6547);
nand U8975 (N_8975,N_6934,N_6626);
nand U8976 (N_8976,N_7325,N_7151);
xnor U8977 (N_8977,N_6955,N_7024);
nor U8978 (N_8978,N_7459,N_7196);
and U8979 (N_8979,N_6719,N_7565);
or U8980 (N_8980,N_6164,N_6107);
nand U8981 (N_8981,N_6201,N_6779);
xnor U8982 (N_8982,N_6700,N_6365);
or U8983 (N_8983,N_6838,N_6839);
nand U8984 (N_8984,N_6391,N_7558);
and U8985 (N_8985,N_6227,N_7363);
or U8986 (N_8986,N_7733,N_6005);
nor U8987 (N_8987,N_7616,N_7761);
nand U8988 (N_8988,N_6512,N_6235);
xnor U8989 (N_8989,N_6605,N_6836);
or U8990 (N_8990,N_7713,N_6666);
nor U8991 (N_8991,N_7315,N_7274);
nand U8992 (N_8992,N_6110,N_6691);
and U8993 (N_8993,N_7271,N_7785);
and U8994 (N_8994,N_6192,N_6711);
nor U8995 (N_8995,N_6189,N_7157);
xor U8996 (N_8996,N_7921,N_7668);
and U8997 (N_8997,N_7303,N_6922);
nor U8998 (N_8998,N_6758,N_7970);
or U8999 (N_8999,N_6317,N_7214);
or U9000 (N_9000,N_7406,N_7497);
nor U9001 (N_9001,N_6798,N_7338);
nor U9002 (N_9002,N_7127,N_6128);
and U9003 (N_9003,N_6232,N_6797);
xor U9004 (N_9004,N_6378,N_6626);
and U9005 (N_9005,N_7036,N_7275);
and U9006 (N_9006,N_7607,N_6681);
nor U9007 (N_9007,N_6453,N_6390);
nand U9008 (N_9008,N_6115,N_7840);
nor U9009 (N_9009,N_6842,N_7980);
and U9010 (N_9010,N_7820,N_7119);
nand U9011 (N_9011,N_6473,N_7716);
and U9012 (N_9012,N_6483,N_6835);
and U9013 (N_9013,N_7855,N_7417);
nor U9014 (N_9014,N_7553,N_7510);
nor U9015 (N_9015,N_6867,N_6094);
nor U9016 (N_9016,N_7676,N_7329);
nor U9017 (N_9017,N_6185,N_7833);
nand U9018 (N_9018,N_6240,N_6053);
and U9019 (N_9019,N_7031,N_7740);
or U9020 (N_9020,N_7054,N_6743);
nand U9021 (N_9021,N_6380,N_7625);
and U9022 (N_9022,N_7251,N_6062);
and U9023 (N_9023,N_6803,N_7242);
or U9024 (N_9024,N_6765,N_6016);
nand U9025 (N_9025,N_6721,N_6046);
or U9026 (N_9026,N_7845,N_7347);
nand U9027 (N_9027,N_6211,N_6181);
and U9028 (N_9028,N_7877,N_6994);
and U9029 (N_9029,N_7798,N_7546);
nand U9030 (N_9030,N_6669,N_6884);
or U9031 (N_9031,N_7622,N_6606);
nor U9032 (N_9032,N_7366,N_7485);
nand U9033 (N_9033,N_7490,N_6168);
nor U9034 (N_9034,N_6124,N_6856);
and U9035 (N_9035,N_7630,N_7356);
nor U9036 (N_9036,N_6552,N_6361);
or U9037 (N_9037,N_6772,N_7832);
nand U9038 (N_9038,N_6734,N_6753);
nor U9039 (N_9039,N_7313,N_6841);
nand U9040 (N_9040,N_7014,N_6819);
and U9041 (N_9041,N_6093,N_6120);
nand U9042 (N_9042,N_6301,N_6485);
nor U9043 (N_9043,N_6983,N_7415);
nor U9044 (N_9044,N_7309,N_6098);
or U9045 (N_9045,N_6439,N_7618);
nand U9046 (N_9046,N_7868,N_6368);
nor U9047 (N_9047,N_7953,N_7384);
and U9048 (N_9048,N_6931,N_7240);
nor U9049 (N_9049,N_7409,N_7699);
xnor U9050 (N_9050,N_6599,N_7244);
or U9051 (N_9051,N_6612,N_6978);
or U9052 (N_9052,N_7928,N_7409);
nor U9053 (N_9053,N_6411,N_6205);
and U9054 (N_9054,N_6873,N_7870);
nor U9055 (N_9055,N_7252,N_7407);
nand U9056 (N_9056,N_6259,N_6911);
nor U9057 (N_9057,N_6564,N_7025);
nand U9058 (N_9058,N_6813,N_6436);
or U9059 (N_9059,N_7774,N_6281);
and U9060 (N_9060,N_7565,N_6221);
nor U9061 (N_9061,N_6694,N_7554);
or U9062 (N_9062,N_6757,N_7687);
nand U9063 (N_9063,N_6548,N_7883);
or U9064 (N_9064,N_6603,N_7353);
and U9065 (N_9065,N_6820,N_7226);
nor U9066 (N_9066,N_6923,N_7460);
and U9067 (N_9067,N_6970,N_7048);
xor U9068 (N_9068,N_6611,N_6358);
xor U9069 (N_9069,N_6530,N_6730);
nand U9070 (N_9070,N_6425,N_6303);
nor U9071 (N_9071,N_7428,N_7993);
or U9072 (N_9072,N_6938,N_7296);
nand U9073 (N_9073,N_7578,N_6602);
or U9074 (N_9074,N_7082,N_7354);
and U9075 (N_9075,N_6338,N_6160);
nand U9076 (N_9076,N_6746,N_7977);
nor U9077 (N_9077,N_6225,N_6859);
nand U9078 (N_9078,N_7689,N_7026);
nor U9079 (N_9079,N_7663,N_6346);
xor U9080 (N_9080,N_7877,N_7972);
nand U9081 (N_9081,N_7390,N_6446);
or U9082 (N_9082,N_7586,N_6384);
or U9083 (N_9083,N_6727,N_6076);
nand U9084 (N_9084,N_7512,N_6456);
xnor U9085 (N_9085,N_6774,N_6113);
nand U9086 (N_9086,N_6831,N_6423);
nand U9087 (N_9087,N_6979,N_7761);
nand U9088 (N_9088,N_7054,N_6706);
and U9089 (N_9089,N_6793,N_6946);
nor U9090 (N_9090,N_6701,N_6343);
nor U9091 (N_9091,N_6549,N_7061);
or U9092 (N_9092,N_7065,N_6273);
nand U9093 (N_9093,N_6025,N_6227);
or U9094 (N_9094,N_7990,N_7581);
nor U9095 (N_9095,N_7890,N_7873);
or U9096 (N_9096,N_6206,N_7261);
nor U9097 (N_9097,N_6018,N_6329);
nor U9098 (N_9098,N_6275,N_7744);
nand U9099 (N_9099,N_7294,N_6447);
nand U9100 (N_9100,N_6318,N_6373);
or U9101 (N_9101,N_6244,N_6089);
or U9102 (N_9102,N_7779,N_6230);
xor U9103 (N_9103,N_7184,N_6612);
xor U9104 (N_9104,N_7894,N_6294);
nor U9105 (N_9105,N_7978,N_6683);
or U9106 (N_9106,N_7540,N_6772);
nand U9107 (N_9107,N_7154,N_7321);
nor U9108 (N_9108,N_7817,N_7435);
and U9109 (N_9109,N_7120,N_7436);
and U9110 (N_9110,N_6098,N_7842);
nand U9111 (N_9111,N_7453,N_7670);
xor U9112 (N_9112,N_7462,N_6676);
nand U9113 (N_9113,N_7130,N_7459);
xnor U9114 (N_9114,N_6513,N_7255);
nor U9115 (N_9115,N_6856,N_6936);
xor U9116 (N_9116,N_7333,N_7485);
nor U9117 (N_9117,N_6116,N_6450);
or U9118 (N_9118,N_7085,N_6004);
and U9119 (N_9119,N_7303,N_7098);
nor U9120 (N_9120,N_7898,N_6725);
nand U9121 (N_9121,N_7793,N_7006);
or U9122 (N_9122,N_6411,N_7525);
and U9123 (N_9123,N_7603,N_6312);
or U9124 (N_9124,N_6706,N_6104);
and U9125 (N_9125,N_6390,N_6194);
and U9126 (N_9126,N_7849,N_7984);
and U9127 (N_9127,N_7857,N_6709);
and U9128 (N_9128,N_6770,N_6184);
and U9129 (N_9129,N_7695,N_7479);
or U9130 (N_9130,N_7309,N_6159);
nor U9131 (N_9131,N_6388,N_6001);
nand U9132 (N_9132,N_6044,N_6796);
nand U9133 (N_9133,N_7384,N_7171);
nor U9134 (N_9134,N_6945,N_7409);
nor U9135 (N_9135,N_7529,N_7624);
nand U9136 (N_9136,N_6056,N_6269);
or U9137 (N_9137,N_7419,N_6008);
nor U9138 (N_9138,N_7901,N_6190);
and U9139 (N_9139,N_6422,N_6260);
nand U9140 (N_9140,N_6922,N_6040);
and U9141 (N_9141,N_7238,N_6304);
or U9142 (N_9142,N_7843,N_7045);
and U9143 (N_9143,N_7377,N_7936);
or U9144 (N_9144,N_6103,N_6992);
nor U9145 (N_9145,N_6609,N_7652);
nor U9146 (N_9146,N_6276,N_6954);
and U9147 (N_9147,N_7681,N_6715);
nor U9148 (N_9148,N_7220,N_7857);
and U9149 (N_9149,N_7811,N_6943);
nor U9150 (N_9150,N_7127,N_7986);
or U9151 (N_9151,N_7701,N_6764);
or U9152 (N_9152,N_6457,N_6097);
nor U9153 (N_9153,N_6067,N_6424);
nand U9154 (N_9154,N_7506,N_7650);
nor U9155 (N_9155,N_6296,N_6685);
or U9156 (N_9156,N_6777,N_6344);
xor U9157 (N_9157,N_6192,N_6586);
and U9158 (N_9158,N_6080,N_7189);
or U9159 (N_9159,N_6287,N_7242);
and U9160 (N_9160,N_6027,N_7582);
or U9161 (N_9161,N_6251,N_6810);
nor U9162 (N_9162,N_7154,N_6113);
nand U9163 (N_9163,N_6665,N_6436);
or U9164 (N_9164,N_7182,N_6420);
nor U9165 (N_9165,N_7348,N_7179);
nand U9166 (N_9166,N_6362,N_7112);
and U9167 (N_9167,N_7336,N_7902);
or U9168 (N_9168,N_6233,N_7299);
or U9169 (N_9169,N_7482,N_6847);
and U9170 (N_9170,N_7424,N_6772);
and U9171 (N_9171,N_7472,N_7851);
or U9172 (N_9172,N_6315,N_6369);
and U9173 (N_9173,N_7616,N_6133);
and U9174 (N_9174,N_7736,N_6106);
nor U9175 (N_9175,N_6441,N_6856);
nand U9176 (N_9176,N_7980,N_6493);
nand U9177 (N_9177,N_7685,N_7835);
nor U9178 (N_9178,N_7444,N_6446);
nand U9179 (N_9179,N_7672,N_7811);
nand U9180 (N_9180,N_7506,N_7915);
or U9181 (N_9181,N_6308,N_7047);
nor U9182 (N_9182,N_7669,N_7787);
nor U9183 (N_9183,N_7957,N_7946);
and U9184 (N_9184,N_7384,N_6201);
and U9185 (N_9185,N_6536,N_6033);
and U9186 (N_9186,N_7288,N_7981);
xor U9187 (N_9187,N_6703,N_6596);
and U9188 (N_9188,N_7320,N_7455);
nor U9189 (N_9189,N_6971,N_6106);
nor U9190 (N_9190,N_7716,N_7782);
nand U9191 (N_9191,N_6391,N_7634);
nand U9192 (N_9192,N_6943,N_6603);
xnor U9193 (N_9193,N_7906,N_6407);
nor U9194 (N_9194,N_7478,N_7902);
nand U9195 (N_9195,N_6502,N_6119);
nand U9196 (N_9196,N_6431,N_6208);
nand U9197 (N_9197,N_7133,N_7249);
nand U9198 (N_9198,N_7969,N_7398);
and U9199 (N_9199,N_7596,N_6717);
or U9200 (N_9200,N_7741,N_7270);
xor U9201 (N_9201,N_6981,N_6755);
and U9202 (N_9202,N_6442,N_7121);
and U9203 (N_9203,N_7786,N_7177);
and U9204 (N_9204,N_7690,N_6290);
nand U9205 (N_9205,N_6410,N_6468);
or U9206 (N_9206,N_7802,N_6518);
or U9207 (N_9207,N_7553,N_7550);
nor U9208 (N_9208,N_6309,N_6855);
and U9209 (N_9209,N_6574,N_6550);
nor U9210 (N_9210,N_6435,N_6394);
and U9211 (N_9211,N_7752,N_6459);
nor U9212 (N_9212,N_6736,N_7807);
or U9213 (N_9213,N_7201,N_7065);
nor U9214 (N_9214,N_6843,N_6259);
xor U9215 (N_9215,N_7482,N_6084);
or U9216 (N_9216,N_7232,N_7319);
and U9217 (N_9217,N_7382,N_6207);
and U9218 (N_9218,N_6143,N_7255);
nand U9219 (N_9219,N_6829,N_6409);
or U9220 (N_9220,N_7726,N_6141);
or U9221 (N_9221,N_6541,N_7174);
or U9222 (N_9222,N_6446,N_7440);
nand U9223 (N_9223,N_6034,N_7761);
nor U9224 (N_9224,N_6559,N_6930);
nand U9225 (N_9225,N_7438,N_6711);
nand U9226 (N_9226,N_7127,N_6262);
nand U9227 (N_9227,N_6586,N_7299);
or U9228 (N_9228,N_6093,N_6656);
nand U9229 (N_9229,N_6547,N_7401);
or U9230 (N_9230,N_6445,N_7165);
and U9231 (N_9231,N_7094,N_7463);
xnor U9232 (N_9232,N_6364,N_7756);
nand U9233 (N_9233,N_7470,N_6893);
and U9234 (N_9234,N_6241,N_7775);
xnor U9235 (N_9235,N_7028,N_7925);
and U9236 (N_9236,N_6276,N_7578);
or U9237 (N_9237,N_7097,N_6764);
or U9238 (N_9238,N_7383,N_7551);
nand U9239 (N_9239,N_6082,N_7330);
nand U9240 (N_9240,N_6853,N_7765);
nand U9241 (N_9241,N_7439,N_7867);
and U9242 (N_9242,N_6875,N_6371);
nor U9243 (N_9243,N_6861,N_7034);
nand U9244 (N_9244,N_7096,N_6671);
or U9245 (N_9245,N_7036,N_7713);
and U9246 (N_9246,N_7340,N_7204);
nand U9247 (N_9247,N_6317,N_7239);
nor U9248 (N_9248,N_7248,N_6269);
xor U9249 (N_9249,N_7981,N_7132);
nand U9250 (N_9250,N_7663,N_7821);
nor U9251 (N_9251,N_7957,N_7079);
nor U9252 (N_9252,N_6645,N_7333);
nor U9253 (N_9253,N_7271,N_7309);
nor U9254 (N_9254,N_7225,N_7097);
and U9255 (N_9255,N_7254,N_6056);
nor U9256 (N_9256,N_6357,N_6852);
nor U9257 (N_9257,N_6680,N_6879);
nand U9258 (N_9258,N_6576,N_7613);
nand U9259 (N_9259,N_7350,N_6151);
xnor U9260 (N_9260,N_6687,N_7161);
xnor U9261 (N_9261,N_6053,N_6088);
or U9262 (N_9262,N_6281,N_6852);
nand U9263 (N_9263,N_6173,N_6400);
nand U9264 (N_9264,N_7001,N_6507);
and U9265 (N_9265,N_6106,N_6698);
nor U9266 (N_9266,N_6886,N_6438);
or U9267 (N_9267,N_6085,N_6260);
nand U9268 (N_9268,N_6833,N_6402);
or U9269 (N_9269,N_6111,N_6395);
or U9270 (N_9270,N_7487,N_7819);
xnor U9271 (N_9271,N_7118,N_6805);
and U9272 (N_9272,N_6520,N_6414);
and U9273 (N_9273,N_6382,N_6114);
and U9274 (N_9274,N_6090,N_7255);
xor U9275 (N_9275,N_6300,N_6242);
nor U9276 (N_9276,N_6292,N_6518);
and U9277 (N_9277,N_7349,N_7337);
xor U9278 (N_9278,N_7921,N_7993);
nor U9279 (N_9279,N_7503,N_6850);
nor U9280 (N_9280,N_7058,N_7422);
nand U9281 (N_9281,N_6380,N_7553);
nor U9282 (N_9282,N_7267,N_7026);
and U9283 (N_9283,N_7755,N_7185);
or U9284 (N_9284,N_7195,N_7559);
nor U9285 (N_9285,N_6517,N_7168);
nand U9286 (N_9286,N_6323,N_6963);
nand U9287 (N_9287,N_7822,N_7552);
nor U9288 (N_9288,N_7432,N_7148);
or U9289 (N_9289,N_7751,N_6478);
and U9290 (N_9290,N_7097,N_6258);
and U9291 (N_9291,N_7411,N_7955);
or U9292 (N_9292,N_6718,N_7348);
nor U9293 (N_9293,N_6193,N_7888);
and U9294 (N_9294,N_6559,N_7484);
and U9295 (N_9295,N_7488,N_6186);
nand U9296 (N_9296,N_6336,N_6535);
nand U9297 (N_9297,N_7942,N_6181);
and U9298 (N_9298,N_6827,N_7160);
and U9299 (N_9299,N_6381,N_6252);
nand U9300 (N_9300,N_6710,N_6448);
or U9301 (N_9301,N_6383,N_6788);
nand U9302 (N_9302,N_7140,N_6224);
nor U9303 (N_9303,N_7429,N_6628);
xor U9304 (N_9304,N_7113,N_7784);
or U9305 (N_9305,N_6863,N_6163);
xnor U9306 (N_9306,N_6016,N_7358);
and U9307 (N_9307,N_7911,N_7629);
or U9308 (N_9308,N_7658,N_7906);
or U9309 (N_9309,N_7443,N_6213);
nand U9310 (N_9310,N_7850,N_6255);
nand U9311 (N_9311,N_6946,N_7166);
and U9312 (N_9312,N_6943,N_7709);
and U9313 (N_9313,N_6195,N_6292);
nor U9314 (N_9314,N_6967,N_7034);
or U9315 (N_9315,N_6978,N_6744);
nand U9316 (N_9316,N_6724,N_7126);
and U9317 (N_9317,N_7977,N_6259);
and U9318 (N_9318,N_6447,N_6458);
and U9319 (N_9319,N_6208,N_7381);
nor U9320 (N_9320,N_6496,N_6904);
or U9321 (N_9321,N_6027,N_7706);
and U9322 (N_9322,N_6305,N_7529);
nor U9323 (N_9323,N_7749,N_6336);
and U9324 (N_9324,N_6969,N_6610);
and U9325 (N_9325,N_7629,N_7939);
nand U9326 (N_9326,N_7201,N_7638);
or U9327 (N_9327,N_7110,N_6897);
nand U9328 (N_9328,N_6195,N_7686);
nor U9329 (N_9329,N_6013,N_7509);
nor U9330 (N_9330,N_7806,N_6926);
xnor U9331 (N_9331,N_7131,N_7421);
nor U9332 (N_9332,N_6473,N_6638);
nor U9333 (N_9333,N_7221,N_6136);
or U9334 (N_9334,N_6434,N_7213);
xor U9335 (N_9335,N_7293,N_6480);
nand U9336 (N_9336,N_6987,N_6630);
nor U9337 (N_9337,N_7260,N_6139);
nand U9338 (N_9338,N_6505,N_7727);
and U9339 (N_9339,N_7601,N_7869);
xnor U9340 (N_9340,N_7589,N_6270);
or U9341 (N_9341,N_6342,N_6337);
or U9342 (N_9342,N_6426,N_7810);
xnor U9343 (N_9343,N_7630,N_6457);
and U9344 (N_9344,N_7970,N_7439);
nand U9345 (N_9345,N_7612,N_7245);
nor U9346 (N_9346,N_6252,N_6998);
nand U9347 (N_9347,N_6317,N_6084);
nor U9348 (N_9348,N_7490,N_6722);
nor U9349 (N_9349,N_6901,N_7709);
nand U9350 (N_9350,N_7129,N_7910);
nor U9351 (N_9351,N_6818,N_6702);
nor U9352 (N_9352,N_7427,N_7191);
nand U9353 (N_9353,N_6262,N_6086);
and U9354 (N_9354,N_7281,N_7366);
nor U9355 (N_9355,N_7229,N_6427);
xor U9356 (N_9356,N_7191,N_7628);
and U9357 (N_9357,N_6050,N_7603);
and U9358 (N_9358,N_6193,N_6714);
xnor U9359 (N_9359,N_6249,N_7301);
or U9360 (N_9360,N_6023,N_6581);
or U9361 (N_9361,N_6728,N_6595);
or U9362 (N_9362,N_6175,N_7211);
nand U9363 (N_9363,N_7998,N_6293);
or U9364 (N_9364,N_7342,N_7420);
or U9365 (N_9365,N_6646,N_6334);
nor U9366 (N_9366,N_7605,N_7640);
nand U9367 (N_9367,N_6237,N_6804);
xnor U9368 (N_9368,N_7370,N_6442);
nand U9369 (N_9369,N_6279,N_6916);
xnor U9370 (N_9370,N_7767,N_7983);
xor U9371 (N_9371,N_7258,N_6778);
xor U9372 (N_9372,N_6936,N_7531);
nand U9373 (N_9373,N_7815,N_7972);
nor U9374 (N_9374,N_6431,N_7308);
or U9375 (N_9375,N_6198,N_7782);
nand U9376 (N_9376,N_7064,N_6288);
xnor U9377 (N_9377,N_6681,N_6935);
xor U9378 (N_9378,N_7064,N_7172);
xor U9379 (N_9379,N_7754,N_6955);
nand U9380 (N_9380,N_6768,N_7780);
xnor U9381 (N_9381,N_7497,N_7188);
or U9382 (N_9382,N_6077,N_7558);
nor U9383 (N_9383,N_6676,N_7687);
and U9384 (N_9384,N_6736,N_6262);
and U9385 (N_9385,N_7116,N_7311);
and U9386 (N_9386,N_6818,N_7049);
nor U9387 (N_9387,N_7902,N_7628);
or U9388 (N_9388,N_6315,N_7788);
or U9389 (N_9389,N_6994,N_7097);
or U9390 (N_9390,N_6861,N_7171);
nand U9391 (N_9391,N_7009,N_7858);
or U9392 (N_9392,N_6860,N_6189);
or U9393 (N_9393,N_7051,N_7630);
and U9394 (N_9394,N_7009,N_6826);
nor U9395 (N_9395,N_6380,N_6292);
nand U9396 (N_9396,N_7351,N_7415);
or U9397 (N_9397,N_7107,N_7374);
and U9398 (N_9398,N_6057,N_7887);
nand U9399 (N_9399,N_7899,N_6348);
nor U9400 (N_9400,N_6337,N_6825);
nand U9401 (N_9401,N_6980,N_7275);
and U9402 (N_9402,N_7706,N_7731);
or U9403 (N_9403,N_7968,N_7031);
nand U9404 (N_9404,N_7020,N_7794);
nand U9405 (N_9405,N_6603,N_7668);
and U9406 (N_9406,N_7125,N_6716);
and U9407 (N_9407,N_7410,N_7066);
or U9408 (N_9408,N_6453,N_7985);
and U9409 (N_9409,N_7305,N_6394);
nor U9410 (N_9410,N_6169,N_7828);
or U9411 (N_9411,N_7475,N_7139);
nand U9412 (N_9412,N_7437,N_7369);
or U9413 (N_9413,N_7303,N_6369);
or U9414 (N_9414,N_6158,N_6684);
nand U9415 (N_9415,N_6640,N_7500);
nor U9416 (N_9416,N_6783,N_7474);
and U9417 (N_9417,N_7234,N_6569);
and U9418 (N_9418,N_6123,N_6117);
or U9419 (N_9419,N_6654,N_6722);
and U9420 (N_9420,N_6662,N_6822);
nand U9421 (N_9421,N_6484,N_6690);
nand U9422 (N_9422,N_7813,N_6086);
or U9423 (N_9423,N_7699,N_7491);
nor U9424 (N_9424,N_6494,N_7324);
nor U9425 (N_9425,N_6868,N_6966);
nor U9426 (N_9426,N_6236,N_7775);
nor U9427 (N_9427,N_6983,N_6076);
or U9428 (N_9428,N_7769,N_6171);
nor U9429 (N_9429,N_7874,N_6458);
and U9430 (N_9430,N_6628,N_6120);
and U9431 (N_9431,N_7554,N_6255);
or U9432 (N_9432,N_6748,N_6195);
nand U9433 (N_9433,N_6735,N_7705);
nor U9434 (N_9434,N_6664,N_7871);
nand U9435 (N_9435,N_6976,N_7912);
nand U9436 (N_9436,N_7363,N_7825);
and U9437 (N_9437,N_7014,N_7822);
and U9438 (N_9438,N_7191,N_6415);
nor U9439 (N_9439,N_7086,N_7826);
or U9440 (N_9440,N_7854,N_6978);
nand U9441 (N_9441,N_6352,N_6835);
nor U9442 (N_9442,N_7730,N_6242);
or U9443 (N_9443,N_7947,N_6598);
xor U9444 (N_9444,N_6208,N_6775);
or U9445 (N_9445,N_7229,N_6544);
nor U9446 (N_9446,N_7574,N_7275);
and U9447 (N_9447,N_7957,N_7049);
and U9448 (N_9448,N_7006,N_7131);
xor U9449 (N_9449,N_6303,N_7601);
xnor U9450 (N_9450,N_7497,N_6180);
nor U9451 (N_9451,N_7987,N_7559);
or U9452 (N_9452,N_6908,N_7204);
nand U9453 (N_9453,N_7773,N_7007);
nand U9454 (N_9454,N_7808,N_6916);
xor U9455 (N_9455,N_7558,N_7633);
or U9456 (N_9456,N_7208,N_7233);
and U9457 (N_9457,N_6985,N_7260);
or U9458 (N_9458,N_7646,N_6305);
and U9459 (N_9459,N_7687,N_6513);
or U9460 (N_9460,N_7528,N_7860);
and U9461 (N_9461,N_7085,N_7369);
nand U9462 (N_9462,N_7578,N_6685);
and U9463 (N_9463,N_6325,N_6390);
nor U9464 (N_9464,N_7463,N_7219);
and U9465 (N_9465,N_7768,N_6538);
xor U9466 (N_9466,N_7604,N_7815);
nor U9467 (N_9467,N_7833,N_6834);
or U9468 (N_9468,N_6758,N_7662);
nor U9469 (N_9469,N_6648,N_6492);
and U9470 (N_9470,N_7695,N_6994);
xnor U9471 (N_9471,N_7026,N_7437);
or U9472 (N_9472,N_6877,N_7333);
or U9473 (N_9473,N_6183,N_6028);
nand U9474 (N_9474,N_7254,N_7452);
and U9475 (N_9475,N_7893,N_7831);
and U9476 (N_9476,N_7458,N_7173);
and U9477 (N_9477,N_7530,N_7551);
nand U9478 (N_9478,N_6018,N_6846);
nand U9479 (N_9479,N_7767,N_6718);
and U9480 (N_9480,N_6265,N_6133);
and U9481 (N_9481,N_7755,N_7637);
xor U9482 (N_9482,N_7334,N_7891);
and U9483 (N_9483,N_6278,N_7237);
and U9484 (N_9484,N_7563,N_7492);
nor U9485 (N_9485,N_7511,N_7553);
and U9486 (N_9486,N_7801,N_6387);
nor U9487 (N_9487,N_6715,N_7881);
nor U9488 (N_9488,N_7140,N_7739);
nand U9489 (N_9489,N_7323,N_6912);
and U9490 (N_9490,N_6283,N_7040);
nor U9491 (N_9491,N_6992,N_6168);
and U9492 (N_9492,N_7954,N_6239);
xor U9493 (N_9493,N_6280,N_6828);
and U9494 (N_9494,N_7895,N_7963);
nor U9495 (N_9495,N_7866,N_6386);
nor U9496 (N_9496,N_7275,N_7101);
or U9497 (N_9497,N_7344,N_6802);
xnor U9498 (N_9498,N_6332,N_7316);
or U9499 (N_9499,N_6451,N_6175);
and U9500 (N_9500,N_7444,N_7309);
or U9501 (N_9501,N_7329,N_6806);
nand U9502 (N_9502,N_6035,N_7325);
or U9503 (N_9503,N_7405,N_7779);
and U9504 (N_9504,N_7596,N_7479);
nand U9505 (N_9505,N_6986,N_6729);
nand U9506 (N_9506,N_7722,N_6654);
nor U9507 (N_9507,N_6637,N_6052);
nor U9508 (N_9508,N_6700,N_7713);
or U9509 (N_9509,N_7949,N_6332);
xor U9510 (N_9510,N_6999,N_7415);
and U9511 (N_9511,N_7514,N_7552);
or U9512 (N_9512,N_7628,N_7099);
or U9513 (N_9513,N_6460,N_7763);
and U9514 (N_9514,N_6582,N_6810);
nand U9515 (N_9515,N_6428,N_6954);
nor U9516 (N_9516,N_7498,N_6726);
nand U9517 (N_9517,N_7624,N_7725);
xor U9518 (N_9518,N_6452,N_6603);
or U9519 (N_9519,N_6489,N_6062);
or U9520 (N_9520,N_7483,N_6102);
and U9521 (N_9521,N_7536,N_6843);
or U9522 (N_9522,N_7684,N_7505);
nand U9523 (N_9523,N_6503,N_7402);
or U9524 (N_9524,N_7093,N_6493);
xor U9525 (N_9525,N_7823,N_7585);
nand U9526 (N_9526,N_6926,N_7282);
nor U9527 (N_9527,N_7329,N_6866);
nor U9528 (N_9528,N_7452,N_6300);
or U9529 (N_9529,N_7906,N_7572);
nor U9530 (N_9530,N_7606,N_6319);
and U9531 (N_9531,N_6461,N_6394);
or U9532 (N_9532,N_7050,N_6088);
or U9533 (N_9533,N_7198,N_6565);
nor U9534 (N_9534,N_6764,N_6664);
nand U9535 (N_9535,N_6241,N_6940);
or U9536 (N_9536,N_7612,N_6671);
or U9537 (N_9537,N_6869,N_6069);
or U9538 (N_9538,N_7634,N_7929);
nor U9539 (N_9539,N_7079,N_7141);
or U9540 (N_9540,N_6260,N_7093);
nor U9541 (N_9541,N_6563,N_6167);
and U9542 (N_9542,N_7360,N_7287);
xor U9543 (N_9543,N_6806,N_7948);
nand U9544 (N_9544,N_7598,N_7842);
or U9545 (N_9545,N_6167,N_7394);
or U9546 (N_9546,N_7213,N_6536);
nand U9547 (N_9547,N_7807,N_7241);
nor U9548 (N_9548,N_7611,N_7568);
and U9549 (N_9549,N_6616,N_6431);
nor U9550 (N_9550,N_6867,N_7023);
nor U9551 (N_9551,N_6421,N_6414);
or U9552 (N_9552,N_6620,N_6675);
nor U9553 (N_9553,N_7739,N_6398);
nand U9554 (N_9554,N_6005,N_7009);
or U9555 (N_9555,N_7492,N_7440);
nor U9556 (N_9556,N_6915,N_6814);
xor U9557 (N_9557,N_7663,N_7863);
xor U9558 (N_9558,N_7276,N_6966);
xor U9559 (N_9559,N_7992,N_6170);
or U9560 (N_9560,N_7759,N_6603);
or U9561 (N_9561,N_7151,N_6094);
and U9562 (N_9562,N_6898,N_6808);
nand U9563 (N_9563,N_6518,N_7479);
and U9564 (N_9564,N_6099,N_6340);
or U9565 (N_9565,N_7931,N_7061);
and U9566 (N_9566,N_6870,N_7252);
xor U9567 (N_9567,N_7050,N_7518);
nor U9568 (N_9568,N_7378,N_6650);
nor U9569 (N_9569,N_7186,N_7329);
and U9570 (N_9570,N_6441,N_7863);
nor U9571 (N_9571,N_7566,N_7829);
nor U9572 (N_9572,N_6770,N_7411);
or U9573 (N_9573,N_6752,N_7887);
nand U9574 (N_9574,N_7822,N_7203);
or U9575 (N_9575,N_7061,N_6455);
or U9576 (N_9576,N_7433,N_7208);
xnor U9577 (N_9577,N_6465,N_7581);
and U9578 (N_9578,N_6918,N_6806);
xnor U9579 (N_9579,N_7130,N_6652);
and U9580 (N_9580,N_6316,N_7577);
nand U9581 (N_9581,N_6950,N_7495);
and U9582 (N_9582,N_6555,N_7111);
xor U9583 (N_9583,N_7568,N_6217);
or U9584 (N_9584,N_6189,N_6195);
nor U9585 (N_9585,N_7870,N_7468);
nand U9586 (N_9586,N_6003,N_7002);
or U9587 (N_9587,N_6251,N_7328);
nor U9588 (N_9588,N_7365,N_6165);
or U9589 (N_9589,N_6466,N_7770);
or U9590 (N_9590,N_7595,N_7732);
nor U9591 (N_9591,N_6944,N_6832);
and U9592 (N_9592,N_6623,N_6647);
nor U9593 (N_9593,N_7337,N_7328);
and U9594 (N_9594,N_7557,N_6517);
or U9595 (N_9595,N_7084,N_7277);
nand U9596 (N_9596,N_7517,N_7216);
or U9597 (N_9597,N_7083,N_6337);
nand U9598 (N_9598,N_7201,N_6373);
and U9599 (N_9599,N_7398,N_7247);
nor U9600 (N_9600,N_6389,N_7357);
nand U9601 (N_9601,N_6021,N_7334);
and U9602 (N_9602,N_7164,N_6531);
nor U9603 (N_9603,N_6202,N_7437);
and U9604 (N_9604,N_6641,N_6633);
and U9605 (N_9605,N_7583,N_7910);
or U9606 (N_9606,N_6033,N_7737);
and U9607 (N_9607,N_6398,N_6533);
and U9608 (N_9608,N_7583,N_7469);
nand U9609 (N_9609,N_7439,N_6713);
or U9610 (N_9610,N_6020,N_7194);
nand U9611 (N_9611,N_7230,N_7837);
nor U9612 (N_9612,N_7834,N_6154);
nand U9613 (N_9613,N_7319,N_6720);
and U9614 (N_9614,N_6680,N_7714);
xor U9615 (N_9615,N_6385,N_7733);
xor U9616 (N_9616,N_6249,N_7436);
nor U9617 (N_9617,N_6392,N_6488);
xor U9618 (N_9618,N_6753,N_6510);
or U9619 (N_9619,N_6166,N_7444);
nand U9620 (N_9620,N_7766,N_7265);
nand U9621 (N_9621,N_6654,N_7053);
nand U9622 (N_9622,N_6138,N_7735);
nand U9623 (N_9623,N_7309,N_6901);
and U9624 (N_9624,N_6544,N_6413);
xor U9625 (N_9625,N_6066,N_6633);
or U9626 (N_9626,N_6729,N_7365);
nor U9627 (N_9627,N_7737,N_7485);
and U9628 (N_9628,N_7433,N_7601);
or U9629 (N_9629,N_7369,N_7838);
nor U9630 (N_9630,N_6729,N_6306);
nor U9631 (N_9631,N_7517,N_6653);
and U9632 (N_9632,N_7341,N_6338);
or U9633 (N_9633,N_6088,N_7774);
or U9634 (N_9634,N_6793,N_7707);
and U9635 (N_9635,N_7185,N_6620);
nand U9636 (N_9636,N_7470,N_7150);
nor U9637 (N_9637,N_7545,N_7994);
nor U9638 (N_9638,N_7911,N_7977);
nor U9639 (N_9639,N_6363,N_6174);
nor U9640 (N_9640,N_6109,N_7294);
nor U9641 (N_9641,N_6864,N_6708);
or U9642 (N_9642,N_6393,N_7557);
and U9643 (N_9643,N_7883,N_7591);
nor U9644 (N_9644,N_7331,N_7806);
and U9645 (N_9645,N_6234,N_7047);
nor U9646 (N_9646,N_7034,N_7862);
or U9647 (N_9647,N_6215,N_7397);
nand U9648 (N_9648,N_7505,N_6053);
or U9649 (N_9649,N_7904,N_6788);
and U9650 (N_9650,N_7798,N_7682);
nand U9651 (N_9651,N_7131,N_6634);
xor U9652 (N_9652,N_7034,N_7442);
nand U9653 (N_9653,N_6009,N_7003);
nor U9654 (N_9654,N_7877,N_6279);
nand U9655 (N_9655,N_6792,N_7581);
and U9656 (N_9656,N_7748,N_6317);
nor U9657 (N_9657,N_6995,N_6301);
nor U9658 (N_9658,N_7330,N_7270);
nor U9659 (N_9659,N_6321,N_7296);
and U9660 (N_9660,N_7633,N_7629);
nand U9661 (N_9661,N_7440,N_6592);
or U9662 (N_9662,N_7385,N_6472);
nor U9663 (N_9663,N_6419,N_6250);
or U9664 (N_9664,N_6791,N_7275);
or U9665 (N_9665,N_7483,N_7161);
xor U9666 (N_9666,N_7092,N_7320);
xor U9667 (N_9667,N_7418,N_6207);
or U9668 (N_9668,N_6192,N_7817);
or U9669 (N_9669,N_7447,N_7409);
and U9670 (N_9670,N_6791,N_7965);
nor U9671 (N_9671,N_6102,N_7386);
nor U9672 (N_9672,N_7907,N_7437);
nor U9673 (N_9673,N_6087,N_6386);
and U9674 (N_9674,N_6230,N_6028);
xnor U9675 (N_9675,N_7744,N_6568);
xnor U9676 (N_9676,N_6096,N_7483);
or U9677 (N_9677,N_7500,N_7145);
nor U9678 (N_9678,N_7720,N_6941);
or U9679 (N_9679,N_7951,N_6370);
nor U9680 (N_9680,N_6142,N_7408);
nor U9681 (N_9681,N_6922,N_6974);
or U9682 (N_9682,N_7718,N_6727);
xnor U9683 (N_9683,N_6250,N_6674);
or U9684 (N_9684,N_6660,N_7700);
nand U9685 (N_9685,N_7379,N_6042);
nor U9686 (N_9686,N_7528,N_6886);
or U9687 (N_9687,N_7542,N_7269);
and U9688 (N_9688,N_7731,N_6357);
and U9689 (N_9689,N_6274,N_6864);
nor U9690 (N_9690,N_6351,N_6793);
nor U9691 (N_9691,N_7585,N_7209);
nand U9692 (N_9692,N_7098,N_6168);
nand U9693 (N_9693,N_7735,N_6915);
or U9694 (N_9694,N_6900,N_7181);
or U9695 (N_9695,N_7920,N_7622);
or U9696 (N_9696,N_6855,N_7752);
and U9697 (N_9697,N_6746,N_7903);
nor U9698 (N_9698,N_7502,N_6617);
nand U9699 (N_9699,N_7165,N_7075);
nand U9700 (N_9700,N_7269,N_7083);
nand U9701 (N_9701,N_6182,N_6552);
and U9702 (N_9702,N_7613,N_7503);
or U9703 (N_9703,N_6400,N_7101);
or U9704 (N_9704,N_7962,N_6800);
nor U9705 (N_9705,N_6917,N_7432);
nor U9706 (N_9706,N_7111,N_6553);
or U9707 (N_9707,N_7727,N_7843);
xor U9708 (N_9708,N_6210,N_6747);
nand U9709 (N_9709,N_6372,N_6580);
nand U9710 (N_9710,N_7978,N_7146);
and U9711 (N_9711,N_7575,N_6347);
and U9712 (N_9712,N_6048,N_6067);
xor U9713 (N_9713,N_7713,N_6180);
or U9714 (N_9714,N_7534,N_7691);
nor U9715 (N_9715,N_7291,N_6486);
nand U9716 (N_9716,N_6038,N_7275);
nor U9717 (N_9717,N_6503,N_6918);
nor U9718 (N_9718,N_6034,N_7050);
nor U9719 (N_9719,N_7248,N_7151);
nor U9720 (N_9720,N_7847,N_6796);
and U9721 (N_9721,N_7808,N_6704);
nand U9722 (N_9722,N_6580,N_7940);
nor U9723 (N_9723,N_7139,N_7040);
xnor U9724 (N_9724,N_6211,N_7236);
nor U9725 (N_9725,N_7928,N_6277);
nand U9726 (N_9726,N_6723,N_6396);
and U9727 (N_9727,N_7844,N_6961);
nor U9728 (N_9728,N_7509,N_7347);
or U9729 (N_9729,N_7237,N_7106);
or U9730 (N_9730,N_6478,N_7774);
nand U9731 (N_9731,N_6022,N_6973);
or U9732 (N_9732,N_7378,N_7571);
nor U9733 (N_9733,N_6335,N_6912);
and U9734 (N_9734,N_6901,N_6161);
nand U9735 (N_9735,N_7574,N_7508);
nor U9736 (N_9736,N_6984,N_7164);
nand U9737 (N_9737,N_7832,N_7726);
nor U9738 (N_9738,N_6540,N_6555);
nor U9739 (N_9739,N_7736,N_6281);
and U9740 (N_9740,N_6771,N_6383);
or U9741 (N_9741,N_7361,N_7897);
and U9742 (N_9742,N_7772,N_7608);
or U9743 (N_9743,N_7659,N_7181);
or U9744 (N_9744,N_7552,N_6206);
nor U9745 (N_9745,N_7945,N_7268);
nor U9746 (N_9746,N_6000,N_6769);
nor U9747 (N_9747,N_6464,N_7257);
nand U9748 (N_9748,N_7112,N_6491);
nor U9749 (N_9749,N_7370,N_6384);
or U9750 (N_9750,N_7279,N_6305);
nor U9751 (N_9751,N_6203,N_6356);
nand U9752 (N_9752,N_6641,N_7425);
and U9753 (N_9753,N_6210,N_6946);
nor U9754 (N_9754,N_7798,N_6829);
or U9755 (N_9755,N_6364,N_6601);
and U9756 (N_9756,N_6874,N_6224);
nor U9757 (N_9757,N_6319,N_6581);
nor U9758 (N_9758,N_7468,N_6809);
nor U9759 (N_9759,N_6197,N_6383);
and U9760 (N_9760,N_6916,N_6105);
nor U9761 (N_9761,N_6696,N_6121);
or U9762 (N_9762,N_6747,N_6266);
nor U9763 (N_9763,N_7067,N_7629);
nand U9764 (N_9764,N_6000,N_7930);
or U9765 (N_9765,N_6877,N_6634);
or U9766 (N_9766,N_6962,N_7781);
nand U9767 (N_9767,N_6311,N_7870);
and U9768 (N_9768,N_6111,N_7773);
or U9769 (N_9769,N_6334,N_6374);
nor U9770 (N_9770,N_7249,N_7248);
nor U9771 (N_9771,N_7013,N_6119);
or U9772 (N_9772,N_7473,N_7853);
or U9773 (N_9773,N_6804,N_7720);
nand U9774 (N_9774,N_6626,N_7703);
nor U9775 (N_9775,N_6537,N_6769);
nor U9776 (N_9776,N_7510,N_7872);
or U9777 (N_9777,N_6165,N_6023);
nand U9778 (N_9778,N_7967,N_6392);
and U9779 (N_9779,N_7770,N_7117);
or U9780 (N_9780,N_6879,N_6442);
nand U9781 (N_9781,N_7403,N_6032);
nand U9782 (N_9782,N_7151,N_6044);
or U9783 (N_9783,N_7408,N_6169);
and U9784 (N_9784,N_6996,N_6796);
nand U9785 (N_9785,N_6183,N_6444);
or U9786 (N_9786,N_7311,N_7375);
or U9787 (N_9787,N_6345,N_7569);
nand U9788 (N_9788,N_6216,N_6331);
or U9789 (N_9789,N_6278,N_6459);
nor U9790 (N_9790,N_7797,N_7015);
nand U9791 (N_9791,N_7522,N_6665);
nor U9792 (N_9792,N_7151,N_7107);
nand U9793 (N_9793,N_6447,N_6903);
and U9794 (N_9794,N_7570,N_7986);
nand U9795 (N_9795,N_6475,N_6643);
or U9796 (N_9796,N_6331,N_7503);
and U9797 (N_9797,N_7374,N_7493);
and U9798 (N_9798,N_6475,N_7082);
and U9799 (N_9799,N_7668,N_6321);
and U9800 (N_9800,N_7390,N_6795);
xor U9801 (N_9801,N_7321,N_6202);
nor U9802 (N_9802,N_6705,N_6477);
or U9803 (N_9803,N_7847,N_6684);
nand U9804 (N_9804,N_6586,N_7314);
and U9805 (N_9805,N_6375,N_6660);
or U9806 (N_9806,N_6563,N_6661);
nor U9807 (N_9807,N_7963,N_7641);
nand U9808 (N_9808,N_6364,N_7022);
xnor U9809 (N_9809,N_6833,N_6571);
xor U9810 (N_9810,N_6529,N_7030);
nor U9811 (N_9811,N_6757,N_6833);
nand U9812 (N_9812,N_7026,N_7425);
nor U9813 (N_9813,N_6649,N_7974);
xnor U9814 (N_9814,N_7746,N_7254);
nor U9815 (N_9815,N_6494,N_7279);
and U9816 (N_9816,N_6567,N_7530);
and U9817 (N_9817,N_6862,N_7139);
nor U9818 (N_9818,N_6083,N_6177);
and U9819 (N_9819,N_6816,N_6261);
xnor U9820 (N_9820,N_6091,N_6148);
and U9821 (N_9821,N_6631,N_6108);
or U9822 (N_9822,N_7866,N_6660);
xor U9823 (N_9823,N_6873,N_6940);
nor U9824 (N_9824,N_6291,N_7678);
nor U9825 (N_9825,N_7627,N_7092);
nand U9826 (N_9826,N_6486,N_7524);
and U9827 (N_9827,N_7340,N_7886);
and U9828 (N_9828,N_6752,N_6509);
xnor U9829 (N_9829,N_6456,N_7877);
and U9830 (N_9830,N_7532,N_6883);
nor U9831 (N_9831,N_6743,N_6388);
nand U9832 (N_9832,N_7230,N_6452);
nand U9833 (N_9833,N_6833,N_6816);
or U9834 (N_9834,N_6454,N_6402);
and U9835 (N_9835,N_6760,N_6798);
nor U9836 (N_9836,N_6126,N_7751);
or U9837 (N_9837,N_7659,N_7945);
and U9838 (N_9838,N_6014,N_7457);
and U9839 (N_9839,N_6975,N_7946);
nand U9840 (N_9840,N_7065,N_7455);
nor U9841 (N_9841,N_7540,N_6043);
or U9842 (N_9842,N_7203,N_6744);
and U9843 (N_9843,N_6466,N_7288);
or U9844 (N_9844,N_6917,N_7292);
and U9845 (N_9845,N_7547,N_7306);
or U9846 (N_9846,N_6527,N_6583);
nor U9847 (N_9847,N_7910,N_6151);
xnor U9848 (N_9848,N_6648,N_6918);
and U9849 (N_9849,N_7783,N_7545);
or U9850 (N_9850,N_7313,N_6202);
xnor U9851 (N_9851,N_6577,N_6189);
nor U9852 (N_9852,N_7445,N_7211);
or U9853 (N_9853,N_6512,N_6296);
nand U9854 (N_9854,N_7398,N_7636);
nor U9855 (N_9855,N_7567,N_7559);
and U9856 (N_9856,N_7576,N_6247);
nand U9857 (N_9857,N_6993,N_6307);
xor U9858 (N_9858,N_7450,N_6317);
nor U9859 (N_9859,N_6184,N_6843);
xnor U9860 (N_9860,N_6051,N_6530);
and U9861 (N_9861,N_6298,N_6536);
nor U9862 (N_9862,N_7830,N_7946);
or U9863 (N_9863,N_6188,N_7866);
and U9864 (N_9864,N_7638,N_7780);
xnor U9865 (N_9865,N_6855,N_6815);
nand U9866 (N_9866,N_7977,N_6056);
or U9867 (N_9867,N_6544,N_6996);
or U9868 (N_9868,N_6248,N_6553);
xnor U9869 (N_9869,N_6740,N_6950);
or U9870 (N_9870,N_7992,N_6828);
nand U9871 (N_9871,N_7802,N_7539);
nor U9872 (N_9872,N_6570,N_7022);
nand U9873 (N_9873,N_7595,N_6964);
nand U9874 (N_9874,N_6106,N_6211);
and U9875 (N_9875,N_6290,N_6181);
or U9876 (N_9876,N_7770,N_7103);
nand U9877 (N_9877,N_6903,N_6258);
xor U9878 (N_9878,N_7895,N_7237);
nand U9879 (N_9879,N_6447,N_7975);
nor U9880 (N_9880,N_7698,N_7622);
nand U9881 (N_9881,N_7326,N_7407);
or U9882 (N_9882,N_6405,N_6872);
or U9883 (N_9883,N_7234,N_7571);
xor U9884 (N_9884,N_7860,N_6018);
nor U9885 (N_9885,N_6028,N_6721);
nand U9886 (N_9886,N_7292,N_7692);
nand U9887 (N_9887,N_7660,N_6776);
xnor U9888 (N_9888,N_7327,N_7489);
and U9889 (N_9889,N_6532,N_6609);
or U9890 (N_9890,N_7356,N_7990);
nor U9891 (N_9891,N_7941,N_7597);
nor U9892 (N_9892,N_6610,N_6963);
nor U9893 (N_9893,N_6645,N_7574);
nand U9894 (N_9894,N_7327,N_6240);
or U9895 (N_9895,N_6236,N_7117);
and U9896 (N_9896,N_7687,N_7658);
or U9897 (N_9897,N_6803,N_6353);
and U9898 (N_9898,N_6855,N_6279);
nand U9899 (N_9899,N_6774,N_7317);
nor U9900 (N_9900,N_7683,N_7612);
or U9901 (N_9901,N_7173,N_7393);
or U9902 (N_9902,N_6300,N_7713);
nand U9903 (N_9903,N_7932,N_6472);
nand U9904 (N_9904,N_6382,N_7922);
and U9905 (N_9905,N_7537,N_7045);
and U9906 (N_9906,N_7078,N_7549);
nor U9907 (N_9907,N_7552,N_6459);
or U9908 (N_9908,N_6597,N_6677);
xor U9909 (N_9909,N_7480,N_7939);
and U9910 (N_9910,N_7122,N_7371);
and U9911 (N_9911,N_7213,N_6031);
or U9912 (N_9912,N_7883,N_6740);
nor U9913 (N_9913,N_6589,N_7293);
or U9914 (N_9914,N_7560,N_6513);
or U9915 (N_9915,N_7575,N_6965);
nor U9916 (N_9916,N_7393,N_6448);
nand U9917 (N_9917,N_7603,N_6238);
or U9918 (N_9918,N_6538,N_6198);
nor U9919 (N_9919,N_7445,N_6470);
nand U9920 (N_9920,N_7071,N_7728);
nand U9921 (N_9921,N_7293,N_7941);
or U9922 (N_9922,N_6467,N_6679);
or U9923 (N_9923,N_6217,N_6488);
and U9924 (N_9924,N_6050,N_6068);
and U9925 (N_9925,N_6476,N_6639);
nand U9926 (N_9926,N_7646,N_6678);
and U9927 (N_9927,N_6261,N_6861);
and U9928 (N_9928,N_6544,N_7299);
nand U9929 (N_9929,N_6602,N_7887);
nand U9930 (N_9930,N_7328,N_6991);
or U9931 (N_9931,N_6205,N_6498);
and U9932 (N_9932,N_6082,N_6383);
nor U9933 (N_9933,N_7556,N_6204);
nor U9934 (N_9934,N_6526,N_6593);
nand U9935 (N_9935,N_7757,N_7282);
or U9936 (N_9936,N_6971,N_6006);
or U9937 (N_9937,N_6530,N_7940);
nand U9938 (N_9938,N_6671,N_7947);
and U9939 (N_9939,N_6478,N_7750);
and U9940 (N_9940,N_7257,N_6340);
or U9941 (N_9941,N_7584,N_6621);
nor U9942 (N_9942,N_7611,N_6104);
nand U9943 (N_9943,N_7868,N_6311);
or U9944 (N_9944,N_6179,N_6359);
nor U9945 (N_9945,N_6826,N_7177);
nand U9946 (N_9946,N_6652,N_6630);
and U9947 (N_9947,N_6745,N_6805);
nand U9948 (N_9948,N_6990,N_7197);
and U9949 (N_9949,N_6767,N_6594);
or U9950 (N_9950,N_7042,N_7896);
xnor U9951 (N_9951,N_7928,N_7805);
nor U9952 (N_9952,N_6881,N_7105);
or U9953 (N_9953,N_6822,N_6735);
nor U9954 (N_9954,N_6895,N_6272);
nand U9955 (N_9955,N_6740,N_6221);
or U9956 (N_9956,N_7771,N_7705);
or U9957 (N_9957,N_6502,N_6494);
or U9958 (N_9958,N_7937,N_6618);
and U9959 (N_9959,N_6653,N_6253);
nand U9960 (N_9960,N_6327,N_6158);
nand U9961 (N_9961,N_7106,N_7604);
or U9962 (N_9962,N_7629,N_7330);
xnor U9963 (N_9963,N_7657,N_7597);
or U9964 (N_9964,N_7718,N_7846);
xnor U9965 (N_9965,N_7330,N_7626);
and U9966 (N_9966,N_7947,N_6131);
nand U9967 (N_9967,N_7387,N_6217);
nand U9968 (N_9968,N_7372,N_7809);
and U9969 (N_9969,N_7617,N_6406);
nand U9970 (N_9970,N_7367,N_6377);
nor U9971 (N_9971,N_7268,N_7442);
nand U9972 (N_9972,N_7257,N_6714);
or U9973 (N_9973,N_6779,N_6328);
or U9974 (N_9974,N_6920,N_7601);
nor U9975 (N_9975,N_6650,N_7780);
nor U9976 (N_9976,N_6108,N_7596);
or U9977 (N_9977,N_7536,N_7511);
nand U9978 (N_9978,N_6038,N_6760);
nor U9979 (N_9979,N_6719,N_7553);
or U9980 (N_9980,N_6042,N_6331);
nor U9981 (N_9981,N_7077,N_6639);
nor U9982 (N_9982,N_6318,N_7486);
nand U9983 (N_9983,N_7922,N_7994);
or U9984 (N_9984,N_7419,N_6532);
xnor U9985 (N_9985,N_7741,N_6713);
or U9986 (N_9986,N_6141,N_7741);
nand U9987 (N_9987,N_6108,N_6468);
nor U9988 (N_9988,N_7893,N_7520);
or U9989 (N_9989,N_7893,N_7456);
nor U9990 (N_9990,N_6778,N_7014);
or U9991 (N_9991,N_7513,N_7659);
nand U9992 (N_9992,N_7341,N_7704);
nand U9993 (N_9993,N_7492,N_6494);
xnor U9994 (N_9994,N_6167,N_6646);
nand U9995 (N_9995,N_7064,N_7708);
nor U9996 (N_9996,N_7534,N_6864);
and U9997 (N_9997,N_7638,N_7544);
nor U9998 (N_9998,N_7510,N_7762);
nand U9999 (N_9999,N_6435,N_7530);
or UO_0 (O_0,N_9562,N_8086);
xnor UO_1 (O_1,N_9041,N_9643);
nor UO_2 (O_2,N_9935,N_9660);
nand UO_3 (O_3,N_9081,N_9474);
or UO_4 (O_4,N_9869,N_9141);
nand UO_5 (O_5,N_9342,N_9183);
and UO_6 (O_6,N_8011,N_9299);
nor UO_7 (O_7,N_9467,N_9149);
or UO_8 (O_8,N_9551,N_8314);
or UO_9 (O_9,N_9791,N_9675);
nand UO_10 (O_10,N_9876,N_9622);
nand UO_11 (O_11,N_8069,N_9086);
and UO_12 (O_12,N_9512,N_9497);
nor UO_13 (O_13,N_8167,N_8198);
and UO_14 (O_14,N_8413,N_9648);
nor UO_15 (O_15,N_9953,N_8348);
or UO_16 (O_16,N_8565,N_9872);
or UO_17 (O_17,N_9752,N_9559);
nand UO_18 (O_18,N_8634,N_8131);
nand UO_19 (O_19,N_8029,N_9504);
and UO_20 (O_20,N_9138,N_9315);
or UO_21 (O_21,N_9939,N_9679);
nor UO_22 (O_22,N_8951,N_8989);
nor UO_23 (O_23,N_9166,N_8145);
or UO_24 (O_24,N_8098,N_8187);
xnor UO_25 (O_25,N_9806,N_8068);
and UO_26 (O_26,N_8263,N_8383);
nand UO_27 (O_27,N_8447,N_9819);
nand UO_28 (O_28,N_9054,N_9764);
nand UO_29 (O_29,N_9451,N_9775);
or UO_30 (O_30,N_8518,N_9613);
nand UO_31 (O_31,N_8859,N_9453);
nand UO_32 (O_32,N_9347,N_9820);
or UO_33 (O_33,N_9947,N_8467);
nor UO_34 (O_34,N_9069,N_9962);
xnor UO_35 (O_35,N_8705,N_8328);
and UO_36 (O_36,N_9331,N_8508);
nor UO_37 (O_37,N_8577,N_9236);
nand UO_38 (O_38,N_8191,N_8762);
nor UO_39 (O_39,N_9080,N_9237);
and UO_40 (O_40,N_9986,N_8226);
nand UO_41 (O_41,N_8470,N_9289);
and UO_42 (O_42,N_9618,N_9416);
xor UO_43 (O_43,N_8689,N_8387);
nand UO_44 (O_44,N_9387,N_8775);
or UO_45 (O_45,N_9240,N_8540);
nor UO_46 (O_46,N_8400,N_9544);
xor UO_47 (O_47,N_8599,N_9473);
or UO_48 (O_48,N_8062,N_9824);
xor UO_49 (O_49,N_8290,N_9663);
xnor UO_50 (O_50,N_9298,N_8258);
nand UO_51 (O_51,N_9136,N_8351);
and UO_52 (O_52,N_8428,N_8305);
or UO_53 (O_53,N_8552,N_9659);
nand UO_54 (O_54,N_9634,N_9248);
nor UO_55 (O_55,N_9624,N_8378);
or UO_56 (O_56,N_8169,N_9513);
or UO_57 (O_57,N_9734,N_8390);
or UO_58 (O_58,N_8717,N_9501);
nand UO_59 (O_59,N_8287,N_9860);
and UO_60 (O_60,N_9528,N_9014);
nor UO_61 (O_61,N_8589,N_9281);
and UO_62 (O_62,N_8507,N_8255);
nor UO_63 (O_63,N_9181,N_8529);
and UO_64 (O_64,N_9162,N_8993);
and UO_65 (O_65,N_8481,N_9768);
and UO_66 (O_66,N_8528,N_8855);
or UO_67 (O_67,N_9914,N_9175);
or UO_68 (O_68,N_9150,N_9147);
nor UO_69 (O_69,N_9484,N_8054);
nor UO_70 (O_70,N_9977,N_9856);
nand UO_71 (O_71,N_9079,N_9524);
nor UO_72 (O_72,N_9087,N_8444);
nand UO_73 (O_73,N_9530,N_9950);
and UO_74 (O_74,N_8306,N_9182);
and UO_75 (O_75,N_8120,N_9034);
xnor UO_76 (O_76,N_9554,N_9038);
nand UO_77 (O_77,N_9793,N_9796);
nor UO_78 (O_78,N_9447,N_8064);
nand UO_79 (O_79,N_8431,N_9408);
and UO_80 (O_80,N_8190,N_9714);
nor UO_81 (O_81,N_9811,N_8141);
xnor UO_82 (O_82,N_8632,N_8071);
nand UO_83 (O_83,N_9572,N_9592);
nor UO_84 (O_84,N_8184,N_9144);
nor UO_85 (O_85,N_8964,N_8970);
and UO_86 (O_86,N_8417,N_9421);
or UO_87 (O_87,N_8566,N_9760);
nand UO_88 (O_88,N_9531,N_8690);
nor UO_89 (O_89,N_9328,N_9568);
or UO_90 (O_90,N_9871,N_8002);
and UO_91 (O_91,N_8580,N_8237);
or UO_92 (O_92,N_9085,N_9642);
xnor UO_93 (O_93,N_9156,N_9174);
and UO_94 (O_94,N_9365,N_9912);
nor UO_95 (O_95,N_9699,N_9410);
nand UO_96 (O_96,N_9353,N_8977);
nor UO_97 (O_97,N_8605,N_8683);
or UO_98 (O_98,N_9160,N_9225);
nand UO_99 (O_99,N_9946,N_9340);
and UO_100 (O_100,N_9930,N_8665);
xnor UO_101 (O_101,N_8020,N_9197);
and UO_102 (O_102,N_9461,N_8743);
nand UO_103 (O_103,N_9858,N_9841);
or UO_104 (O_104,N_8028,N_8721);
nor UO_105 (O_105,N_8979,N_9193);
or UO_106 (O_106,N_9435,N_8407);
or UO_107 (O_107,N_8077,N_9605);
nor UO_108 (O_108,N_8746,N_9620);
and UO_109 (O_109,N_9655,N_8199);
nor UO_110 (O_110,N_9252,N_8049);
and UO_111 (O_111,N_8525,N_8489);
and UO_112 (O_112,N_9534,N_9446);
xnor UO_113 (O_113,N_9688,N_9427);
nand UO_114 (O_114,N_9617,N_9722);
or UO_115 (O_115,N_9724,N_8543);
nor UO_116 (O_116,N_9619,N_9604);
and UO_117 (O_117,N_8569,N_8896);
nand UO_118 (O_118,N_8371,N_9867);
nand UO_119 (O_119,N_8202,N_8381);
nand UO_120 (O_120,N_9143,N_8241);
and UO_121 (O_121,N_8960,N_9486);
and UO_122 (O_122,N_9850,N_8596);
and UO_123 (O_123,N_9987,N_9165);
nor UO_124 (O_124,N_8653,N_8587);
nand UO_125 (O_125,N_9934,N_8445);
nand UO_126 (O_126,N_9809,N_8398);
xor UO_127 (O_127,N_9626,N_9201);
nand UO_128 (O_128,N_8253,N_9723);
xor UO_129 (O_129,N_8004,N_9703);
and UO_130 (O_130,N_9212,N_8695);
nand UO_131 (O_131,N_8363,N_8227);
or UO_132 (O_132,N_8629,N_9903);
and UO_133 (O_133,N_8396,N_8225);
nor UO_134 (O_134,N_9857,N_9433);
or UO_135 (O_135,N_9747,N_8078);
or UO_136 (O_136,N_9595,N_8531);
or UO_137 (O_137,N_8292,N_8358);
nand UO_138 (O_138,N_8910,N_8975);
nand UO_139 (O_139,N_9976,N_8076);
nand UO_140 (O_140,N_8795,N_9208);
nand UO_141 (O_141,N_8987,N_9273);
nor UO_142 (O_142,N_8493,N_9042);
nand UO_143 (O_143,N_9596,N_8035);
xnor UO_144 (O_144,N_9776,N_9475);
nor UO_145 (O_145,N_9682,N_8461);
nor UO_146 (O_146,N_9535,N_8161);
xnor UO_147 (O_147,N_9506,N_8872);
or UO_148 (O_148,N_9729,N_9279);
nor UO_149 (O_149,N_8688,N_8009);
nand UO_150 (O_150,N_9422,N_9394);
nor UO_151 (O_151,N_8155,N_8965);
xnor UO_152 (O_152,N_8585,N_9094);
nand UO_153 (O_153,N_9966,N_9419);
nand UO_154 (O_154,N_8121,N_8143);
and UO_155 (O_155,N_9509,N_9995);
nor UO_156 (O_156,N_8904,N_9311);
nor UO_157 (O_157,N_9526,N_8716);
nor UO_158 (O_158,N_9961,N_9630);
and UO_159 (O_159,N_9616,N_8671);
and UO_160 (O_160,N_8621,N_8511);
and UO_161 (O_161,N_9721,N_9099);
nand UO_162 (O_162,N_9495,N_9217);
nor UO_163 (O_163,N_8288,N_8276);
and UO_164 (O_164,N_9538,N_8794);
nor UO_165 (O_165,N_8127,N_9442);
or UO_166 (O_166,N_8564,N_8452);
and UO_167 (O_167,N_8070,N_8021);
xnor UO_168 (O_168,N_8442,N_9804);
nor UO_169 (O_169,N_9748,N_9275);
nor UO_170 (O_170,N_8079,N_8016);
and UO_171 (O_171,N_9564,N_9169);
xor UO_172 (O_172,N_8440,N_9058);
nor UO_173 (O_173,N_8033,N_9397);
or UO_174 (O_174,N_9753,N_9980);
nand UO_175 (O_175,N_9579,N_9061);
and UO_176 (O_176,N_8154,N_8425);
nand UO_177 (O_177,N_9478,N_8130);
and UO_178 (O_178,N_9805,N_9052);
nor UO_179 (O_179,N_9482,N_9125);
or UO_180 (O_180,N_9230,N_8483);
or UO_181 (O_181,N_9948,N_9113);
xnor UO_182 (O_182,N_8998,N_8630);
and UO_183 (O_183,N_9516,N_9392);
nand UO_184 (O_184,N_8401,N_8545);
or UO_185 (O_185,N_8034,N_8830);
and UO_186 (O_186,N_8601,N_9910);
and UO_187 (O_187,N_8533,N_9719);
or UO_188 (O_188,N_8860,N_9285);
nor UO_189 (O_189,N_8136,N_9154);
nand UO_190 (O_190,N_8232,N_9272);
or UO_191 (O_191,N_9001,N_8106);
or UO_192 (O_192,N_9098,N_8112);
nor UO_193 (O_193,N_9915,N_9514);
and UO_194 (O_194,N_8789,N_9250);
nor UO_195 (O_195,N_9897,N_8242);
and UO_196 (O_196,N_9778,N_8469);
and UO_197 (O_197,N_8080,N_8831);
and UO_198 (O_198,N_9917,N_8945);
nor UO_199 (O_199,N_9599,N_9018);
nor UO_200 (O_200,N_9883,N_9291);
nor UO_201 (O_201,N_8395,N_8323);
xor UO_202 (O_202,N_9908,N_8494);
and UO_203 (O_203,N_9712,N_8609);
and UO_204 (O_204,N_8419,N_8482);
nand UO_205 (O_205,N_8412,N_8604);
or UO_206 (O_206,N_8666,N_9556);
nand UO_207 (O_207,N_8727,N_9350);
or UO_208 (O_208,N_9194,N_9116);
nor UO_209 (O_209,N_8844,N_8884);
xnor UO_210 (O_210,N_8359,N_9670);
nand UO_211 (O_211,N_8879,N_9133);
and UO_212 (O_212,N_8886,N_8504);
nand UO_213 (O_213,N_9153,N_8012);
or UO_214 (O_214,N_9677,N_8667);
or UO_215 (O_215,N_8648,N_8075);
and UO_216 (O_216,N_8243,N_8066);
nor UO_217 (O_217,N_9800,N_9582);
nor UO_218 (O_218,N_9701,N_9911);
and UO_219 (O_219,N_8180,N_9294);
or UO_220 (O_220,N_8618,N_9384);
or UO_221 (O_221,N_8092,N_9100);
nor UO_222 (O_222,N_8973,N_9854);
or UO_223 (O_223,N_8228,N_8809);
nand UO_224 (O_224,N_8252,N_9945);
or UO_225 (O_225,N_9831,N_8703);
and UO_226 (O_226,N_9304,N_9577);
or UO_227 (O_227,N_9239,N_9882);
nor UO_228 (O_228,N_9011,N_8538);
nand UO_229 (O_229,N_8777,N_9439);
nand UO_230 (O_230,N_9828,N_9965);
and UO_231 (O_231,N_8072,N_8812);
or UO_232 (O_232,N_8386,N_9529);
nand UO_233 (O_233,N_9573,N_8159);
nor UO_234 (O_234,N_8790,N_8332);
nor UO_235 (O_235,N_8514,N_8819);
or UO_236 (O_236,N_8544,N_8403);
and UO_237 (O_237,N_8772,N_9555);
nor UO_238 (O_238,N_9146,N_9381);
and UO_239 (O_239,N_9647,N_8377);
and UO_240 (O_240,N_9093,N_9866);
or UO_241 (O_241,N_8894,N_8749);
nor UO_242 (O_242,N_9460,N_8600);
or UO_243 (O_243,N_9859,N_8825);
or UO_244 (O_244,N_9296,N_9135);
nor UO_245 (O_245,N_8608,N_8046);
nor UO_246 (O_246,N_9782,N_9810);
nand UO_247 (O_247,N_9881,N_9575);
nand UO_248 (O_248,N_8623,N_8739);
nand UO_249 (O_249,N_9329,N_9766);
xor UO_250 (O_250,N_9834,N_8822);
or UO_251 (O_251,N_8250,N_8279);
nand UO_252 (O_252,N_9375,N_9812);
xor UO_253 (O_253,N_9832,N_9825);
or UO_254 (O_254,N_8846,N_8561);
and UO_255 (O_255,N_8909,N_8924);
or UO_256 (O_256,N_9432,N_8267);
and UO_257 (O_257,N_9465,N_8861);
and UO_258 (O_258,N_8194,N_9145);
or UO_259 (O_259,N_9176,N_9349);
nor UO_260 (O_260,N_9817,N_9108);
xnor UO_261 (O_261,N_8091,N_8513);
or UO_262 (O_262,N_8804,N_9982);
nand UO_263 (O_263,N_9091,N_9785);
and UO_264 (O_264,N_8935,N_8856);
or UO_265 (O_265,N_8810,N_8347);
and UO_266 (O_266,N_8586,N_8327);
and UO_267 (O_267,N_8778,N_8015);
or UO_268 (O_268,N_8857,N_8976);
or UO_269 (O_269,N_8501,N_9971);
nand UO_270 (O_270,N_9887,N_9823);
or UO_271 (O_271,N_8918,N_9126);
or UO_272 (O_272,N_8465,N_9313);
or UO_273 (O_273,N_8952,N_8416);
nand UO_274 (O_274,N_8645,N_8268);
or UO_275 (O_275,N_8754,N_9814);
xnor UO_276 (O_276,N_8438,N_8882);
xnor UO_277 (O_277,N_9715,N_9200);
and UO_278 (O_278,N_8635,N_9813);
nand UO_279 (O_279,N_8492,N_8375);
nor UO_280 (O_280,N_8867,N_9507);
or UO_281 (O_281,N_9424,N_8466);
or UO_282 (O_282,N_9454,N_9082);
xnor UO_283 (O_283,N_9875,N_8298);
or UO_284 (O_284,N_8380,N_9808);
nand UO_285 (O_285,N_9550,N_9765);
or UO_286 (O_286,N_8156,N_8639);
nor UO_287 (O_287,N_8813,N_9491);
nor UO_288 (O_288,N_9187,N_8139);
or UO_289 (O_289,N_8737,N_8551);
nand UO_290 (O_290,N_9137,N_8354);
xor UO_291 (O_291,N_8764,N_9967);
nand UO_292 (O_292,N_9263,N_8474);
nand UO_293 (O_293,N_8738,N_9763);
nor UO_294 (O_294,N_9590,N_9180);
nor UO_295 (O_295,N_8724,N_8248);
nor UO_296 (O_296,N_9155,N_9646);
or UO_297 (O_297,N_9071,N_9282);
or UO_298 (O_298,N_8331,N_8574);
nand UO_299 (O_299,N_8588,N_8610);
and UO_300 (O_300,N_8176,N_9855);
nor UO_301 (O_301,N_9739,N_8388);
or UO_302 (O_302,N_9343,N_9653);
nor UO_303 (O_303,N_9031,N_9428);
or UO_304 (O_304,N_8740,N_9864);
nand UO_305 (O_305,N_8249,N_9319);
nor UO_306 (O_306,N_8758,N_9235);
nand UO_307 (O_307,N_8869,N_8207);
or UO_308 (O_308,N_8111,N_8725);
xor UO_309 (O_309,N_8990,N_9219);
nand UO_310 (O_310,N_8537,N_8369);
nor UO_311 (O_311,N_8256,N_8410);
nand UO_312 (O_312,N_8668,N_8319);
or UO_313 (O_313,N_8505,N_8937);
or UO_314 (O_314,N_8384,N_9131);
nor UO_315 (O_315,N_8573,N_8691);
nor UO_316 (O_316,N_8594,N_8968);
nor UO_317 (O_317,N_8670,N_9068);
nand UO_318 (O_318,N_8506,N_8490);
xor UO_319 (O_319,N_8966,N_8464);
nor UO_320 (O_320,N_9017,N_9731);
nor UO_321 (O_321,N_9493,N_8245);
xor UO_322 (O_322,N_8931,N_8718);
or UO_323 (O_323,N_9756,N_8179);
xnor UO_324 (O_324,N_8753,N_9111);
nand UO_325 (O_325,N_9826,N_9276);
nand UO_326 (O_326,N_9916,N_8863);
nor UO_327 (O_327,N_8972,N_8307);
and UO_328 (O_328,N_8119,N_9284);
xor UO_329 (O_329,N_9578,N_8709);
and UO_330 (O_330,N_9110,N_9413);
nand UO_331 (O_331,N_9633,N_9368);
or UO_332 (O_332,N_9759,N_8811);
or UO_333 (O_333,N_9702,N_8453);
and UO_334 (O_334,N_8415,N_9611);
nand UO_335 (O_335,N_8030,N_8660);
nand UO_336 (O_336,N_8026,N_9191);
nand UO_337 (O_337,N_9733,N_8603);
and UO_338 (O_338,N_8985,N_8956);
nand UO_339 (O_339,N_8353,N_8181);
xor UO_340 (O_340,N_9692,N_9398);
xnor UO_341 (O_341,N_9978,N_8559);
or UO_342 (O_342,N_8053,N_9121);
and UO_343 (O_343,N_9268,N_8949);
nor UO_344 (O_344,N_8224,N_8140);
nor UO_345 (O_345,N_9769,N_8117);
and UO_346 (O_346,N_8881,N_8941);
nor UO_347 (O_347,N_8231,N_9895);
nor UO_348 (O_348,N_8379,N_9015);
nand UO_349 (O_349,N_8424,N_8230);
nor UO_350 (O_350,N_8188,N_9128);
and UO_351 (O_351,N_8959,N_9742);
and UO_352 (O_352,N_8463,N_9401);
nand UO_353 (O_353,N_9520,N_9210);
nand UO_354 (O_354,N_8361,N_8498);
nor UO_355 (O_355,N_8920,N_8297);
nor UO_356 (O_356,N_9414,N_8067);
nand UO_357 (O_357,N_8741,N_9565);
xnor UO_358 (O_358,N_9779,N_8732);
or UO_359 (O_359,N_8244,N_9344);
nand UO_360 (O_360,N_8838,N_9852);
or UO_361 (O_361,N_9704,N_9399);
nand UO_362 (O_362,N_8346,N_9999);
nor UO_363 (O_363,N_9787,N_9332);
or UO_364 (O_364,N_8669,N_8549);
and UO_365 (O_365,N_8729,N_9849);
or UO_366 (O_366,N_8912,N_8938);
nor UO_367 (O_367,N_8850,N_8087);
nor UO_368 (O_368,N_9676,N_9989);
nand UO_369 (O_369,N_9185,N_8907);
nor UO_370 (O_370,N_9683,N_9218);
nand UO_371 (O_371,N_9802,N_8917);
or UO_372 (O_372,N_8783,N_8808);
xnor UO_373 (O_373,N_9735,N_8638);
nand UO_374 (O_374,N_8473,N_8100);
nor UO_375 (O_375,N_9879,N_8829);
nand UO_376 (O_376,N_8591,N_8982);
nand UO_377 (O_377,N_9940,N_8443);
and UO_378 (O_378,N_8969,N_8057);
nand UO_379 (O_379,N_8942,N_8930);
xor UO_380 (O_380,N_9587,N_9525);
nand UO_381 (O_381,N_9784,N_9256);
nand UO_382 (O_382,N_8302,N_9553);
or UO_383 (O_383,N_8271,N_9972);
nand UO_384 (O_384,N_8459,N_9621);
nor UO_385 (O_385,N_8402,N_8877);
or UO_386 (O_386,N_9586,N_9751);
nor UO_387 (O_387,N_8893,N_9593);
xnor UO_388 (O_388,N_8272,N_9990);
nand UO_389 (O_389,N_8044,N_8765);
and UO_390 (O_390,N_8038,N_9786);
nand UO_391 (O_391,N_8891,N_9533);
or UO_392 (O_392,N_9707,N_8643);
or UO_393 (O_393,N_8422,N_8455);
nor UO_394 (O_394,N_9560,N_8488);
or UO_395 (O_395,N_9815,N_9736);
nor UO_396 (O_396,N_9221,N_8160);
xor UO_397 (O_397,N_8771,N_9639);
or UO_398 (O_398,N_9868,N_8581);
or UO_399 (O_399,N_8895,N_9888);
nor UO_400 (O_400,N_8031,N_8368);
xnor UO_401 (O_401,N_9468,N_8206);
nand UO_402 (O_402,N_8868,N_8234);
nand UO_403 (O_403,N_9159,N_8747);
and UO_404 (O_404,N_9229,N_9963);
nor UO_405 (O_405,N_8301,N_8696);
nor UO_406 (O_406,N_8766,N_8278);
nor UO_407 (O_407,N_8595,N_9485);
nor UO_408 (O_408,N_8270,N_8682);
nand UO_409 (O_409,N_9297,N_9196);
nand UO_410 (O_410,N_9277,N_8661);
and UO_411 (O_411,N_8491,N_9244);
and UO_412 (O_412,N_9352,N_9637);
nor UO_413 (O_413,N_8680,N_9681);
nand UO_414 (O_414,N_9177,N_9519);
and UO_415 (O_415,N_8547,N_8730);
nor UO_416 (O_416,N_9696,N_8815);
nand UO_417 (O_417,N_8165,N_8008);
xnor UO_418 (O_418,N_8837,N_9023);
nand UO_419 (O_419,N_9380,N_9892);
or UO_420 (O_420,N_8125,N_9118);
or UO_421 (O_421,N_9089,N_8084);
nor UO_422 (O_422,N_9840,N_9077);
xnor UO_423 (O_423,N_8974,N_8532);
or UO_424 (O_424,N_8343,N_8785);
nand UO_425 (O_425,N_8217,N_9088);
and UO_426 (O_426,N_8720,N_8650);
or UO_427 (O_427,N_9129,N_8997);
nand UO_428 (O_428,N_9674,N_8953);
xor UO_429 (O_429,N_9124,N_8627);
xnor UO_430 (O_430,N_8655,N_8185);
or UO_431 (O_431,N_8572,N_9105);
or UO_432 (O_432,N_9449,N_9561);
and UO_433 (O_433,N_9245,N_8793);
and UO_434 (O_434,N_8592,N_8950);
and UO_435 (O_435,N_8871,N_9691);
nand UO_436 (O_436,N_9346,N_8006);
nand UO_437 (O_437,N_9835,N_8955);
nand UO_438 (O_438,N_9270,N_8657);
and UO_439 (O_439,N_8449,N_8392);
and UO_440 (O_440,N_9743,N_8013);
nor UO_441 (O_441,N_8579,N_8649);
xor UO_442 (O_442,N_9412,N_9207);
nand UO_443 (O_443,N_9374,N_8734);
nand UO_444 (O_444,N_9822,N_9066);
or UO_445 (O_445,N_9644,N_8768);
nor UO_446 (O_446,N_8742,N_8800);
or UO_447 (O_447,N_9333,N_8468);
or UO_448 (O_448,N_9532,N_8906);
or UO_449 (O_449,N_8560,N_8370);
nand UO_450 (O_450,N_9943,N_8750);
and UO_451 (O_451,N_9400,N_8852);
nand UO_452 (O_452,N_8576,N_8409);
nand UO_453 (O_453,N_8058,N_9407);
or UO_454 (O_454,N_8622,N_8770);
nor UO_455 (O_455,N_9157,N_9356);
and UO_456 (O_456,N_8612,N_8209);
or UO_457 (O_457,N_8324,N_9570);
or UO_458 (O_458,N_9580,N_8326);
nand UO_459 (O_459,N_8517,N_8063);
and UO_460 (O_460,N_9255,N_8876);
or UO_461 (O_461,N_9695,N_8752);
nand UO_462 (O_462,N_9838,N_8320);
or UO_463 (O_463,N_8152,N_8684);
and UO_464 (O_464,N_8503,N_8546);
and UO_465 (O_465,N_8858,N_9941);
or UO_466 (O_466,N_8172,N_9758);
and UO_467 (O_467,N_8457,N_8616);
and UO_468 (O_468,N_8122,N_8345);
nand UO_469 (O_469,N_8978,N_8277);
nor UO_470 (O_470,N_9318,N_8497);
and UO_471 (O_471,N_9293,N_8692);
nor UO_472 (O_472,N_9557,N_9777);
and UO_473 (O_473,N_9022,N_9152);
or UO_474 (O_474,N_9005,N_8487);
or UO_475 (O_475,N_9109,N_8052);
xor UO_476 (O_476,N_9689,N_9861);
nand UO_477 (O_477,N_9942,N_8423);
or UO_478 (O_478,N_9890,N_9012);
nand UO_479 (O_479,N_8555,N_9295);
nor UO_480 (O_480,N_8548,N_8512);
and UO_481 (O_481,N_9547,N_8048);
nor UO_482 (O_482,N_9690,N_9338);
nand UO_483 (O_483,N_9443,N_8878);
or UO_484 (O_484,N_9899,N_9900);
nor UO_485 (O_485,N_8699,N_9064);
nand UO_486 (O_486,N_9227,N_9669);
nand UO_487 (O_487,N_8223,N_8756);
nand UO_488 (O_488,N_8710,N_8744);
and UO_489 (O_489,N_8797,N_9862);
or UO_490 (O_490,N_8707,N_9843);
and UO_491 (O_491,N_8236,N_9558);
nand UO_492 (O_492,N_8814,N_8834);
nand UO_493 (O_493,N_8853,N_8939);
and UO_494 (O_494,N_9139,N_8839);
or UO_495 (O_495,N_9312,N_8408);
nand UO_496 (O_496,N_8628,N_9406);
and UO_497 (O_497,N_8128,N_9393);
and UO_498 (O_498,N_9013,N_8539);
nor UO_499 (O_499,N_9035,N_8807);
or UO_500 (O_500,N_8251,N_9923);
and UO_501 (O_501,N_9585,N_9873);
nor UO_502 (O_502,N_8926,N_8175);
nand UO_503 (O_503,N_8626,N_9163);
or UO_504 (O_504,N_9694,N_8065);
nand UO_505 (O_505,N_8748,N_8933);
and UO_506 (O_506,N_8921,N_8366);
and UO_507 (O_507,N_9213,N_9463);
or UO_508 (O_508,N_8568,N_8177);
xnor UO_509 (O_509,N_9974,N_9505);
nand UO_510 (O_510,N_9307,N_9095);
and UO_511 (O_511,N_8847,N_8733);
nand UO_512 (O_512,N_8421,N_9067);
nor UO_513 (O_513,N_9922,N_8673);
and UO_514 (O_514,N_9549,N_8104);
xor UO_515 (O_515,N_9078,N_8686);
nand UO_516 (O_516,N_9223,N_9377);
or UO_517 (O_517,N_9120,N_9002);
or UO_518 (O_518,N_8541,N_8702);
or UO_519 (O_519,N_8003,N_8848);
nand UO_520 (O_520,N_8963,N_8731);
nor UO_521 (O_521,N_9957,N_9395);
nor UO_522 (O_522,N_9258,N_8309);
nor UO_523 (O_523,N_8352,N_8567);
nand UO_524 (O_524,N_8640,N_8385);
and UO_525 (O_525,N_8471,N_9992);
and UO_526 (O_526,N_8597,N_8711);
and UO_527 (O_527,N_9189,N_9970);
or UO_528 (O_528,N_8706,N_8435);
nand UO_529 (O_529,N_8472,N_8123);
nor UO_530 (O_530,N_9671,N_9354);
or UO_531 (O_531,N_8791,N_9437);
or UO_532 (O_532,N_8178,N_9363);
nor UO_533 (O_533,N_9716,N_9203);
or UO_534 (O_534,N_9431,N_9684);
nand UO_535 (O_535,N_9324,N_8835);
or UO_536 (O_536,N_9790,N_8001);
nand UO_537 (O_537,N_8992,N_9305);
or UO_538 (O_538,N_8883,N_8784);
or UO_539 (O_539,N_9429,N_8414);
and UO_540 (O_540,N_8994,N_8674);
and UO_541 (O_541,N_9101,N_8903);
or UO_542 (O_542,N_8905,N_8542);
nand UO_543 (O_543,N_8329,N_8500);
xor UO_544 (O_544,N_9789,N_8041);
or UO_545 (O_545,N_9391,N_8023);
or UO_546 (O_546,N_9204,N_8763);
and UO_547 (O_547,N_9292,N_9511);
or UO_548 (O_548,N_9070,N_8018);
or UO_549 (O_549,N_9726,N_9508);
or UO_550 (O_550,N_9055,N_9405);
or UO_551 (O_551,N_8584,N_8832);
nand UO_552 (O_552,N_9233,N_9283);
and UO_553 (O_553,N_8451,N_9096);
or UO_554 (O_554,N_9322,N_9807);
and UO_555 (O_555,N_9846,N_9016);
or UO_556 (O_556,N_9865,N_9288);
and UO_557 (O_557,N_8318,N_8115);
and UO_558 (O_558,N_8841,N_9072);
nor UO_559 (O_559,N_8901,N_9249);
or UO_560 (O_560,N_9075,N_9678);
nor UO_561 (O_561,N_8947,N_9190);
nor UO_562 (O_562,N_8708,N_8295);
and UO_563 (O_563,N_8116,N_9337);
and UO_564 (O_564,N_8144,N_8129);
and UO_565 (O_565,N_9334,N_8874);
nor UO_566 (O_566,N_9851,N_8678);
and UO_567 (O_567,N_8722,N_9537);
nor UO_568 (O_568,N_9907,N_8336);
nor UO_569 (O_569,N_9316,N_9192);
or UO_570 (O_570,N_9600,N_9848);
or UO_571 (O_571,N_9896,N_8189);
nor UO_572 (O_572,N_9975,N_9541);
and UO_573 (O_573,N_8017,N_8842);
xor UO_574 (O_574,N_9452,N_8265);
and UO_575 (O_575,N_8036,N_8148);
xnor UO_576 (O_576,N_9902,N_9991);
and UO_577 (O_577,N_8282,N_8759);
and UO_578 (O_578,N_9996,N_9664);
nand UO_579 (O_579,N_9919,N_9385);
nand UO_580 (O_580,N_9818,N_9059);
nand UO_581 (O_581,N_8437,N_9998);
nor UO_582 (O_582,N_8496,N_9794);
nor UO_583 (O_583,N_9933,N_8315);
or UO_584 (O_584,N_8192,N_8995);
or UO_585 (O_585,N_9004,N_9837);
nor UO_586 (O_586,N_8254,N_8675);
nand UO_587 (O_587,N_9607,N_8096);
nor UO_588 (O_588,N_9436,N_9969);
xor UO_589 (O_589,N_8010,N_8698);
or UO_590 (O_590,N_9988,N_8355);
or UO_591 (O_591,N_8082,N_9877);
or UO_592 (O_592,N_8043,N_9628);
nor UO_593 (O_593,N_8625,N_8818);
nand UO_594 (O_594,N_9494,N_9909);
and UO_595 (O_595,N_9119,N_9629);
nor UO_596 (O_596,N_8880,N_9490);
nand UO_597 (O_597,N_9464,N_8149);
and UO_598 (O_598,N_9062,N_8168);
xor UO_599 (O_599,N_9030,N_8659);
nor UO_600 (O_600,N_8340,N_8286);
and UO_601 (O_601,N_8337,N_9336);
or UO_602 (O_602,N_8520,N_8114);
and UO_603 (O_603,N_8132,N_8499);
nor UO_604 (O_604,N_8840,N_8602);
or UO_605 (O_605,N_9750,N_8264);
nand UO_606 (O_606,N_9097,N_9545);
nand UO_607 (O_607,N_9112,N_9720);
nand UO_608 (O_608,N_8448,N_8475);
and UO_609 (O_609,N_8662,N_8575);
and UO_610 (O_610,N_8050,N_8875);
and UO_611 (O_611,N_9266,N_8238);
nand UO_612 (O_612,N_9198,N_9216);
nand UO_613 (O_613,N_9594,N_8059);
nor UO_614 (O_614,N_9889,N_8433);
nor UO_615 (O_615,N_9891,N_8356);
nor UO_616 (O_616,N_9386,N_9842);
or UO_617 (O_617,N_8458,N_8478);
xnor UO_618 (O_618,N_8047,N_8946);
or UO_619 (O_619,N_8137,N_9224);
and UO_620 (O_620,N_8658,N_9209);
nand UO_621 (O_621,N_9056,N_8892);
and UO_622 (O_622,N_9047,N_9364);
or UO_623 (O_623,N_9488,N_8317);
nand UO_624 (O_624,N_9323,N_9360);
and UO_625 (O_625,N_8485,N_8304);
nor UO_626 (O_626,N_9046,N_8936);
or UO_627 (O_627,N_9115,N_9717);
or UO_628 (O_628,N_8420,N_8787);
nand UO_629 (O_629,N_9361,N_8056);
or UO_630 (O_630,N_9521,N_9232);
nor UO_631 (O_631,N_9369,N_8193);
nand UO_632 (O_632,N_9003,N_9430);
or UO_633 (O_633,N_9029,N_9402);
or UO_634 (O_634,N_9636,N_8322);
nand UO_635 (O_635,N_8108,N_8019);
nor UO_636 (O_636,N_8103,N_9359);
and UO_637 (O_637,N_9259,N_9472);
xnor UO_638 (O_638,N_9024,N_9280);
and UO_639 (O_639,N_9027,N_9076);
or UO_640 (O_640,N_9130,N_8714);
and UO_641 (O_641,N_9672,N_8195);
or UO_642 (O_642,N_9797,N_8864);
nand UO_643 (O_643,N_8611,N_8646);
or UO_644 (O_644,N_8735,N_9205);
nand UO_645 (O_645,N_8299,N_8477);
or UO_646 (O_646,N_8205,N_9668);
xor UO_647 (O_647,N_8404,N_8827);
nor UO_648 (O_648,N_8303,N_8055);
nand UO_649 (O_649,N_8713,N_9993);
or UO_650 (O_650,N_9983,N_9510);
and UO_651 (O_651,N_8607,N_8590);
or UO_652 (O_652,N_8656,N_8239);
nor UO_653 (O_653,N_9662,N_9958);
and UO_654 (O_654,N_8981,N_8334);
nand UO_655 (O_655,N_8776,N_8045);
and UO_656 (O_656,N_8330,N_9161);
nand UO_657 (O_657,N_9566,N_8865);
nand UO_658 (O_658,N_8240,N_9265);
xor UO_659 (O_659,N_8961,N_8927);
and UO_660 (O_660,N_8786,N_8436);
and UO_661 (O_661,N_9920,N_9792);
or UO_662 (O_662,N_9028,N_8333);
or UO_663 (O_663,N_8073,N_9202);
and UO_664 (O_664,N_9262,N_8781);
and UO_665 (O_665,N_8454,N_8550);
nand UO_666 (O_666,N_9314,N_8996);
nand UO_667 (O_667,N_9774,N_8213);
or UO_668 (O_668,N_8849,N_8200);
nor UO_669 (O_669,N_9762,N_9261);
xor UO_670 (O_670,N_9608,N_9697);
nand UO_671 (O_671,N_9122,N_8958);
nor UO_672 (O_672,N_8074,N_9226);
or UO_673 (O_673,N_8911,N_8364);
nor UO_674 (O_674,N_9317,N_9214);
and UO_675 (O_675,N_8350,N_8767);
nor UO_676 (O_676,N_8983,N_9050);
and UO_677 (O_677,N_8024,N_9536);
xnor UO_678 (O_678,N_8007,N_8898);
xor UO_679 (O_679,N_9114,N_8957);
or UO_680 (O_680,N_9325,N_9839);
nand UO_681 (O_681,N_8430,N_8183);
xor UO_682 (O_682,N_9389,N_9434);
nand UO_683 (O_683,N_8218,N_9417);
nand UO_684 (O_684,N_9680,N_8147);
and UO_685 (O_685,N_9426,N_9745);
nor UO_686 (O_686,N_9376,N_9944);
or UO_687 (O_687,N_9773,N_8557);
nor UO_688 (O_688,N_9257,N_9597);
and UO_689 (O_689,N_8280,N_9656);
or UO_690 (O_690,N_9847,N_8845);
and UO_691 (O_691,N_9184,N_9287);
or UO_692 (O_692,N_9641,N_8556);
and UO_693 (O_693,N_9687,N_9798);
xor UO_694 (O_694,N_8570,N_9795);
or UO_695 (O_695,N_8944,N_8291);
and UO_696 (O_696,N_9327,N_8833);
nor UO_697 (O_697,N_9574,N_8266);
and UO_698 (O_698,N_8885,N_9552);
nand UO_699 (O_699,N_9614,N_8357);
xnor UO_700 (O_700,N_9222,N_8802);
nand UO_701 (O_701,N_8313,N_8633);
or UO_702 (O_702,N_8851,N_9341);
xor UO_703 (O_703,N_8197,N_8113);
or UO_704 (O_704,N_9476,N_8014);
and UO_705 (O_705,N_8900,N_8321);
or UO_706 (O_706,N_8269,N_8980);
and UO_707 (O_707,N_9772,N_9243);
and UO_708 (O_708,N_9780,N_9457);
or UO_709 (O_709,N_8521,N_8426);
and UO_710 (O_710,N_9744,N_8211);
nand UO_711 (O_711,N_9140,N_9043);
or UO_712 (O_712,N_9938,N_8126);
nor UO_713 (O_713,N_9388,N_8134);
nand UO_714 (O_714,N_8434,N_8967);
or UO_715 (O_715,N_9546,N_9517);
and UO_716 (O_716,N_8118,N_9044);
or UO_717 (O_717,N_8162,N_8509);
xor UO_718 (O_718,N_8142,N_8025);
or UO_719 (O_719,N_8817,N_8102);
or UO_720 (O_720,N_9650,N_8124);
and UO_721 (O_721,N_9543,N_8246);
and UO_722 (O_722,N_9496,N_8606);
nor UO_723 (O_723,N_9106,N_9423);
and UO_724 (O_724,N_8925,N_9886);
or UO_725 (O_725,N_8526,N_9799);
and UO_726 (O_726,N_8081,N_9770);
nor UO_727 (O_727,N_9379,N_9415);
nand UO_728 (O_728,N_8094,N_8991);
xnor UO_729 (O_729,N_9649,N_8005);
nand UO_730 (O_730,N_9527,N_9151);
or UO_731 (O_731,N_9026,N_8399);
and UO_732 (O_732,N_8247,N_8578);
nand UO_733 (O_733,N_8374,N_8367);
and UO_734 (O_734,N_9251,N_8151);
nor UO_735 (O_735,N_9480,N_9037);
and UO_736 (O_736,N_8637,N_8524);
or UO_737 (O_737,N_8296,N_8899);
nor UO_738 (O_738,N_9459,N_9658);
nor UO_739 (O_739,N_8365,N_8801);
or UO_740 (O_740,N_9382,N_8220);
or UO_741 (O_741,N_9954,N_8259);
or UO_742 (O_742,N_8971,N_8135);
and UO_743 (O_743,N_8755,N_9051);
nand UO_744 (O_744,N_8216,N_8479);
or UO_745 (O_745,N_8312,N_9215);
nor UO_746 (O_746,N_9477,N_9074);
nand UO_747 (O_747,N_9901,N_9396);
or UO_748 (O_748,N_9104,N_9123);
nand UO_749 (O_749,N_9803,N_9827);
and UO_750 (O_750,N_9878,N_8962);
and UO_751 (O_751,N_9567,N_9260);
xor UO_752 (O_752,N_8214,N_9627);
nor UO_753 (O_753,N_9709,N_9348);
or UO_754 (O_754,N_9968,N_9142);
and UO_755 (O_755,N_9727,N_9749);
nor UO_756 (O_756,N_9601,N_9829);
nand UO_757 (O_757,N_8215,N_8427);
nand UO_758 (O_758,N_9583,N_8429);
xor UO_759 (O_759,N_8663,N_9539);
nor UO_760 (O_760,N_9045,N_9959);
nor UO_761 (O_761,N_9450,N_9186);
nand UO_762 (O_762,N_8389,N_9732);
or UO_763 (O_763,N_9246,N_8923);
nor UO_764 (O_764,N_9373,N_8051);
nor UO_765 (O_765,N_9188,N_9606);
nor UO_766 (O_766,N_9542,N_8099);
or UO_767 (O_767,N_8308,N_8796);
or UO_768 (O_768,N_8338,N_8495);
or UO_769 (O_769,N_8816,N_9499);
nor UO_770 (O_770,N_8235,N_8173);
and UO_771 (O_771,N_8687,N_8300);
or UO_772 (O_772,N_8870,N_9926);
nand UO_773 (O_773,N_8311,N_8519);
xnor UO_774 (O_774,N_9498,N_9362);
nor UO_775 (O_775,N_9320,N_8536);
nand UO_776 (O_776,N_8283,N_9905);
nor UO_777 (O_777,N_9148,N_9730);
nand UO_778 (O_778,N_8257,N_9928);
nor UO_779 (O_779,N_8060,N_8562);
and UO_780 (O_780,N_9652,N_9700);
or UO_781 (O_781,N_8480,N_9053);
nand UO_782 (O_782,N_8164,N_9000);
xnor UO_783 (O_783,N_9403,N_8866);
nor UO_784 (O_784,N_9489,N_9040);
nand UO_785 (O_785,N_9741,N_8681);
or UO_786 (O_786,N_8516,N_8873);
and UO_787 (O_787,N_8676,N_9371);
or UO_788 (O_788,N_8954,N_8163);
and UO_789 (O_789,N_8914,N_8208);
nand UO_790 (O_790,N_9708,N_9358);
nand UO_791 (O_791,N_9836,N_9021);
or UO_792 (O_792,N_9673,N_9746);
and UO_793 (O_793,N_8613,N_9588);
and UO_794 (O_794,N_9894,N_8679);
nand UO_795 (O_795,N_8204,N_8212);
or UO_796 (O_796,N_9979,N_9893);
and UO_797 (O_797,N_8558,N_8462);
and UO_798 (O_798,N_8948,N_8677);
nand UO_799 (O_799,N_9321,N_8418);
or UO_800 (O_800,N_9718,N_9253);
and UO_801 (O_801,N_9060,N_9458);
nand UO_802 (O_802,N_9300,N_9456);
nor UO_803 (O_803,N_9602,N_9821);
or UO_804 (O_804,N_8527,N_8406);
nand UO_805 (O_805,N_9929,N_9009);
xor UO_806 (O_806,N_9880,N_8554);
and UO_807 (O_807,N_8788,N_8393);
nand UO_808 (O_808,N_9390,N_8203);
nand UO_809 (O_809,N_9898,N_9931);
or UO_810 (O_810,N_9960,N_8037);
or UO_811 (O_811,N_8405,N_9609);
or UO_812 (O_812,N_8325,N_8158);
or UO_813 (O_813,N_9994,N_9335);
and UO_814 (O_814,N_9483,N_9048);
nor UO_815 (O_815,N_8439,N_8774);
nor UO_816 (O_816,N_9084,N_9167);
or UO_817 (O_817,N_9132,N_9372);
or UO_818 (O_818,N_8940,N_8779);
or UO_819 (O_819,N_8095,N_9409);
and UO_820 (O_820,N_8854,N_9271);
nor UO_821 (O_821,N_9049,N_9469);
and UO_822 (O_822,N_9581,N_9661);
nor UO_823 (O_823,N_8373,N_9383);
and UO_824 (O_824,N_8598,N_9801);
xnor UO_825 (O_825,N_9303,N_9286);
and UO_826 (O_826,N_9301,N_8615);
and UO_827 (O_827,N_8712,N_9610);
nand UO_828 (O_828,N_9083,N_8943);
nand UO_829 (O_829,N_8523,N_9666);
nor UO_830 (O_830,N_9936,N_8376);
nand UO_831 (O_831,N_8736,N_9171);
nor UO_832 (O_832,N_9267,N_9952);
or UO_833 (O_833,N_8534,N_9569);
nand UO_834 (O_834,N_8262,N_8196);
and UO_835 (O_835,N_8486,N_8182);
nand UO_836 (O_836,N_9503,N_9006);
or UO_837 (O_837,N_9206,N_9170);
nor UO_838 (O_838,N_9710,N_9367);
nor UO_839 (O_839,N_8672,N_8294);
xor UO_840 (O_840,N_8799,N_8929);
nor UO_841 (O_841,N_9020,N_8723);
or UO_842 (O_842,N_9231,N_8110);
or UO_843 (O_843,N_8760,N_9757);
nor UO_844 (O_844,N_8274,N_8260);
nand UO_845 (O_845,N_9269,N_9767);
or UO_846 (O_846,N_9019,N_8715);
and UO_847 (O_847,N_9090,N_9178);
and UO_848 (O_848,N_8908,N_9438);
nor UO_849 (O_849,N_9645,N_9705);
xor UO_850 (O_850,N_8984,N_8888);
or UO_851 (O_851,N_9956,N_9584);
or UO_852 (O_852,N_9500,N_9117);
nand UO_853 (O_853,N_8040,N_9487);
and UO_854 (O_854,N_8685,N_8450);
or UO_855 (O_855,N_8222,N_8456);
and UO_856 (O_856,N_9065,N_9462);
xnor UO_857 (O_857,N_9540,N_8803);
or UO_858 (O_858,N_9092,N_9863);
nor UO_859 (O_859,N_9411,N_9103);
nand UO_860 (O_860,N_9492,N_8027);
or UO_861 (O_861,N_8316,N_9591);
nand UO_862 (O_862,N_8826,N_9563);
and UO_863 (O_863,N_9885,N_8090);
nand UO_864 (O_864,N_9951,N_9651);
nor UO_865 (O_865,N_9711,N_8664);
nand UO_866 (O_866,N_9640,N_8582);
nand UO_867 (O_867,N_8782,N_8484);
and UO_868 (O_868,N_9913,N_8170);
or UO_869 (O_869,N_8726,N_8617);
and UO_870 (O_870,N_9816,N_8843);
nand UO_871 (O_871,N_9625,N_9444);
and UO_872 (O_872,N_9238,N_8032);
xnor UO_873 (O_873,N_9949,N_9783);
nor UO_874 (O_874,N_8285,N_8915);
and UO_875 (O_875,N_9010,N_9698);
or UO_876 (O_876,N_9418,N_9728);
nand UO_877 (O_877,N_9713,N_9598);
nand UO_878 (O_878,N_8798,N_8913);
and UO_879 (O_879,N_8652,N_9632);
or UO_880 (O_880,N_9254,N_8928);
or UO_881 (O_881,N_8097,N_8773);
and UO_882 (O_882,N_8394,N_8109);
or UO_883 (O_883,N_8229,N_8889);
xor UO_884 (O_884,N_8293,N_8631);
and UO_885 (O_885,N_9845,N_8362);
nand UO_886 (O_886,N_8339,N_9172);
xor UO_887 (O_887,N_8583,N_9937);
or UO_888 (O_888,N_9471,N_8751);
nor UO_889 (O_889,N_8341,N_8042);
nand UO_890 (O_890,N_8728,N_9007);
nand UO_891 (O_891,N_9870,N_9844);
and UO_892 (O_892,N_8636,N_9310);
nor UO_893 (O_893,N_8210,N_9548);
or UO_894 (O_894,N_9635,N_9039);
or UO_895 (O_895,N_8289,N_9025);
or UO_896 (O_896,N_9522,N_8769);
and UO_897 (O_897,N_9073,N_8890);
xor UO_898 (O_898,N_9420,N_8806);
and UO_899 (O_899,N_9964,N_9761);
or UO_900 (O_900,N_9984,N_9274);
nor UO_901 (O_901,N_8828,N_8620);
nand UO_902 (O_902,N_8101,N_8563);
or UO_903 (O_903,N_9781,N_9884);
nand UO_904 (O_904,N_8171,N_8897);
xnor UO_905 (O_905,N_8441,N_9173);
and UO_906 (O_906,N_8647,N_9278);
nand UO_907 (O_907,N_9997,N_9440);
xor UO_908 (O_908,N_9370,N_8745);
nor UO_909 (O_909,N_9654,N_8823);
and UO_910 (O_910,N_9247,N_9771);
or UO_911 (O_911,N_9615,N_9033);
and UO_912 (O_912,N_9518,N_8887);
xnor UO_913 (O_913,N_9164,N_8261);
nor UO_914 (O_914,N_9242,N_8916);
nor UO_915 (O_915,N_9339,N_9904);
nand UO_916 (O_916,N_8372,N_8105);
nand UO_917 (O_917,N_9302,N_8061);
and UO_918 (O_918,N_8411,N_9107);
or UO_919 (O_919,N_8088,N_9455);
or UO_920 (O_920,N_8174,N_8644);
xor UO_921 (O_921,N_9754,N_9685);
nand UO_922 (O_922,N_9571,N_8166);
nor UO_923 (O_923,N_8641,N_8432);
nand UO_924 (O_924,N_9158,N_8701);
xor UO_925 (O_925,N_8614,N_9955);
nand UO_926 (O_926,N_8654,N_9925);
or UO_927 (O_927,N_9665,N_9623);
or UO_928 (O_928,N_9228,N_9725);
or UO_929 (O_929,N_8792,N_9366);
and UO_930 (O_930,N_8719,N_8476);
nor UO_931 (O_931,N_8000,N_9924);
or UO_932 (O_932,N_8281,N_8535);
and UO_933 (O_933,N_8934,N_9102);
nand UO_934 (O_934,N_8157,N_9345);
nor UO_935 (O_935,N_9179,N_9667);
or UO_936 (O_936,N_9932,N_8150);
nand UO_937 (O_937,N_9057,N_9330);
or UO_938 (O_938,N_9502,N_8382);
nand UO_939 (O_939,N_8153,N_8999);
or UO_940 (O_940,N_8986,N_8391);
nor UO_941 (O_941,N_9576,N_9351);
and UO_942 (O_942,N_9195,N_9264);
and UO_943 (O_943,N_8335,N_9706);
nor UO_944 (O_944,N_8083,N_9220);
nand UO_945 (O_945,N_8761,N_8530);
nor UO_946 (O_946,N_9985,N_9853);
nand UO_947 (O_947,N_8619,N_8522);
nand UO_948 (O_948,N_8201,N_8460);
and UO_949 (O_949,N_8138,N_8694);
or UO_950 (O_950,N_9355,N_8642);
nand UO_951 (O_951,N_8821,N_9738);
xnor UO_952 (O_952,N_9425,N_9445);
nor UO_953 (O_953,N_9448,N_8133);
nor UO_954 (O_954,N_9523,N_9657);
nand UO_955 (O_955,N_8219,N_9127);
or UO_956 (O_956,N_9479,N_9589);
and UO_957 (O_957,N_8922,N_9612);
nor UO_958 (O_958,N_8700,N_8704);
nand UO_959 (O_959,N_9466,N_8651);
nand UO_960 (O_960,N_8571,N_8902);
and UO_961 (O_961,N_9441,N_8284);
xor UO_962 (O_962,N_9032,N_8342);
and UO_963 (O_963,N_8275,N_9906);
nor UO_964 (O_964,N_9357,N_9788);
nor UO_965 (O_965,N_9740,N_9921);
nor UO_966 (O_966,N_8221,N_8360);
nand UO_967 (O_967,N_8780,N_8146);
xnor UO_968 (O_968,N_9168,N_8932);
nand UO_969 (O_969,N_8697,N_8022);
nor UO_970 (O_970,N_9241,N_8039);
nand UO_971 (O_971,N_9199,N_9211);
nand UO_972 (O_972,N_9638,N_9603);
or UO_973 (O_973,N_8502,N_9737);
nand UO_974 (O_974,N_9234,N_8089);
or UO_975 (O_975,N_8107,N_8510);
or UO_976 (O_976,N_8820,N_9693);
nor UO_977 (O_977,N_8273,N_9686);
nor UO_978 (O_978,N_9918,N_9481);
or UO_979 (O_979,N_9290,N_9326);
and UO_980 (O_980,N_9927,N_8553);
and UO_981 (O_981,N_8593,N_8446);
and UO_982 (O_982,N_8310,N_9470);
xor UO_983 (O_983,N_8862,N_8515);
or UO_984 (O_984,N_9755,N_8836);
nor UO_985 (O_985,N_8349,N_8824);
nor UO_986 (O_986,N_8397,N_8693);
nor UO_987 (O_987,N_8344,N_8085);
nand UO_988 (O_988,N_9874,N_8919);
nand UO_989 (O_989,N_9631,N_9404);
and UO_990 (O_990,N_9515,N_9008);
xor UO_991 (O_991,N_9309,N_8186);
and UO_992 (O_992,N_9830,N_8233);
xnor UO_993 (O_993,N_8093,N_9833);
and UO_994 (O_994,N_9378,N_8988);
nor UO_995 (O_995,N_9973,N_9308);
nand UO_996 (O_996,N_9306,N_9036);
and UO_997 (O_997,N_8624,N_9981);
nand UO_998 (O_998,N_8805,N_8757);
nand UO_999 (O_999,N_9063,N_9134);
or UO_1000 (O_1000,N_9524,N_9779);
or UO_1001 (O_1001,N_8885,N_8408);
xor UO_1002 (O_1002,N_9597,N_9167);
and UO_1003 (O_1003,N_9518,N_9503);
or UO_1004 (O_1004,N_9083,N_8103);
xor UO_1005 (O_1005,N_9851,N_9140);
or UO_1006 (O_1006,N_9173,N_9645);
nor UO_1007 (O_1007,N_9100,N_8611);
nand UO_1008 (O_1008,N_9826,N_9452);
and UO_1009 (O_1009,N_8211,N_9829);
xnor UO_1010 (O_1010,N_8124,N_9498);
and UO_1011 (O_1011,N_9245,N_9136);
nand UO_1012 (O_1012,N_9876,N_8017);
xnor UO_1013 (O_1013,N_8856,N_8933);
or UO_1014 (O_1014,N_8358,N_8108);
or UO_1015 (O_1015,N_9663,N_9667);
nor UO_1016 (O_1016,N_9223,N_8589);
or UO_1017 (O_1017,N_8528,N_8628);
and UO_1018 (O_1018,N_8488,N_8895);
nand UO_1019 (O_1019,N_9437,N_9900);
or UO_1020 (O_1020,N_9625,N_8967);
or UO_1021 (O_1021,N_9153,N_8357);
and UO_1022 (O_1022,N_9201,N_8961);
or UO_1023 (O_1023,N_9744,N_9105);
nand UO_1024 (O_1024,N_9133,N_8476);
nor UO_1025 (O_1025,N_9887,N_9338);
nand UO_1026 (O_1026,N_9320,N_8324);
nor UO_1027 (O_1027,N_8073,N_9675);
or UO_1028 (O_1028,N_8925,N_9162);
nor UO_1029 (O_1029,N_9104,N_9608);
and UO_1030 (O_1030,N_9579,N_9846);
nor UO_1031 (O_1031,N_8899,N_9944);
nor UO_1032 (O_1032,N_8452,N_9110);
or UO_1033 (O_1033,N_8358,N_8280);
or UO_1034 (O_1034,N_8432,N_8884);
nor UO_1035 (O_1035,N_8151,N_9474);
nand UO_1036 (O_1036,N_8045,N_9660);
and UO_1037 (O_1037,N_9156,N_9804);
nand UO_1038 (O_1038,N_8288,N_8373);
nand UO_1039 (O_1039,N_9087,N_9887);
and UO_1040 (O_1040,N_8482,N_8345);
nor UO_1041 (O_1041,N_9235,N_9012);
xnor UO_1042 (O_1042,N_9132,N_9019);
and UO_1043 (O_1043,N_9526,N_8588);
and UO_1044 (O_1044,N_9601,N_8321);
nand UO_1045 (O_1045,N_9826,N_9144);
nor UO_1046 (O_1046,N_9569,N_8197);
and UO_1047 (O_1047,N_8832,N_8978);
or UO_1048 (O_1048,N_8539,N_9499);
and UO_1049 (O_1049,N_9326,N_9730);
or UO_1050 (O_1050,N_8558,N_9885);
nand UO_1051 (O_1051,N_9810,N_9147);
or UO_1052 (O_1052,N_8934,N_9439);
or UO_1053 (O_1053,N_8208,N_9247);
or UO_1054 (O_1054,N_9190,N_9371);
xor UO_1055 (O_1055,N_8051,N_9052);
nand UO_1056 (O_1056,N_8601,N_8784);
and UO_1057 (O_1057,N_9178,N_9869);
nand UO_1058 (O_1058,N_9578,N_8890);
or UO_1059 (O_1059,N_8801,N_8787);
or UO_1060 (O_1060,N_8697,N_9732);
or UO_1061 (O_1061,N_8621,N_9040);
nand UO_1062 (O_1062,N_9107,N_9403);
nor UO_1063 (O_1063,N_8825,N_9951);
nand UO_1064 (O_1064,N_9557,N_8851);
nand UO_1065 (O_1065,N_9250,N_8532);
xnor UO_1066 (O_1066,N_9380,N_9972);
or UO_1067 (O_1067,N_9330,N_8628);
or UO_1068 (O_1068,N_9007,N_9663);
nand UO_1069 (O_1069,N_8458,N_9704);
nand UO_1070 (O_1070,N_9371,N_9078);
nand UO_1071 (O_1071,N_8402,N_9139);
xor UO_1072 (O_1072,N_9292,N_8766);
and UO_1073 (O_1073,N_8894,N_8156);
and UO_1074 (O_1074,N_8870,N_9655);
or UO_1075 (O_1075,N_8891,N_8687);
and UO_1076 (O_1076,N_9015,N_8325);
nand UO_1077 (O_1077,N_8809,N_9980);
xnor UO_1078 (O_1078,N_9558,N_9040);
nor UO_1079 (O_1079,N_8402,N_9815);
nor UO_1080 (O_1080,N_9339,N_9240);
nand UO_1081 (O_1081,N_9658,N_9137);
and UO_1082 (O_1082,N_9948,N_8242);
and UO_1083 (O_1083,N_8454,N_8539);
or UO_1084 (O_1084,N_9184,N_8312);
or UO_1085 (O_1085,N_9972,N_8269);
or UO_1086 (O_1086,N_8337,N_9491);
nor UO_1087 (O_1087,N_8690,N_8482);
or UO_1088 (O_1088,N_9620,N_9566);
nand UO_1089 (O_1089,N_9658,N_9657);
or UO_1090 (O_1090,N_8569,N_8338);
or UO_1091 (O_1091,N_9772,N_9653);
and UO_1092 (O_1092,N_9190,N_8121);
xnor UO_1093 (O_1093,N_8296,N_9150);
xnor UO_1094 (O_1094,N_8170,N_8391);
or UO_1095 (O_1095,N_8986,N_8958);
nor UO_1096 (O_1096,N_9585,N_9352);
or UO_1097 (O_1097,N_8919,N_8910);
and UO_1098 (O_1098,N_8560,N_8028);
and UO_1099 (O_1099,N_9585,N_9392);
or UO_1100 (O_1100,N_9600,N_8079);
nand UO_1101 (O_1101,N_8469,N_9372);
nor UO_1102 (O_1102,N_8965,N_8052);
nor UO_1103 (O_1103,N_9386,N_8570);
xnor UO_1104 (O_1104,N_9073,N_9346);
xor UO_1105 (O_1105,N_8714,N_9263);
nand UO_1106 (O_1106,N_8787,N_8611);
and UO_1107 (O_1107,N_8330,N_9835);
or UO_1108 (O_1108,N_9613,N_8081);
and UO_1109 (O_1109,N_8866,N_9793);
nand UO_1110 (O_1110,N_8353,N_9519);
or UO_1111 (O_1111,N_8295,N_8871);
nand UO_1112 (O_1112,N_9174,N_8820);
or UO_1113 (O_1113,N_9970,N_9956);
xnor UO_1114 (O_1114,N_9483,N_9841);
nand UO_1115 (O_1115,N_9437,N_9958);
nand UO_1116 (O_1116,N_8456,N_9787);
nor UO_1117 (O_1117,N_9486,N_9521);
nor UO_1118 (O_1118,N_9334,N_9553);
nor UO_1119 (O_1119,N_9421,N_8448);
and UO_1120 (O_1120,N_9217,N_8330);
and UO_1121 (O_1121,N_8271,N_9826);
nor UO_1122 (O_1122,N_9549,N_8904);
or UO_1123 (O_1123,N_9148,N_8432);
or UO_1124 (O_1124,N_9310,N_8593);
and UO_1125 (O_1125,N_8715,N_8694);
or UO_1126 (O_1126,N_8460,N_8090);
nor UO_1127 (O_1127,N_8210,N_8678);
and UO_1128 (O_1128,N_8382,N_9979);
and UO_1129 (O_1129,N_8446,N_8148);
xor UO_1130 (O_1130,N_9242,N_9037);
nor UO_1131 (O_1131,N_9512,N_8381);
and UO_1132 (O_1132,N_9113,N_8419);
or UO_1133 (O_1133,N_8501,N_8572);
nor UO_1134 (O_1134,N_9828,N_8794);
nand UO_1135 (O_1135,N_8039,N_8021);
nor UO_1136 (O_1136,N_8485,N_9431);
xnor UO_1137 (O_1137,N_9222,N_8708);
nand UO_1138 (O_1138,N_8043,N_9504);
and UO_1139 (O_1139,N_8272,N_8795);
and UO_1140 (O_1140,N_8027,N_9607);
nor UO_1141 (O_1141,N_8711,N_9821);
xor UO_1142 (O_1142,N_8462,N_8639);
nor UO_1143 (O_1143,N_9738,N_8973);
or UO_1144 (O_1144,N_9255,N_9605);
and UO_1145 (O_1145,N_8541,N_9296);
xor UO_1146 (O_1146,N_8980,N_8841);
nand UO_1147 (O_1147,N_9842,N_8655);
xor UO_1148 (O_1148,N_8530,N_8048);
and UO_1149 (O_1149,N_9368,N_8262);
or UO_1150 (O_1150,N_9461,N_9228);
nor UO_1151 (O_1151,N_9108,N_9578);
nand UO_1152 (O_1152,N_9599,N_9166);
nand UO_1153 (O_1153,N_8705,N_9895);
or UO_1154 (O_1154,N_9709,N_9927);
and UO_1155 (O_1155,N_9939,N_9284);
nand UO_1156 (O_1156,N_8430,N_8162);
nand UO_1157 (O_1157,N_9132,N_8796);
or UO_1158 (O_1158,N_9448,N_9628);
nand UO_1159 (O_1159,N_9330,N_9519);
nor UO_1160 (O_1160,N_9432,N_8459);
or UO_1161 (O_1161,N_8731,N_8055);
and UO_1162 (O_1162,N_9582,N_9356);
or UO_1163 (O_1163,N_8950,N_9776);
nor UO_1164 (O_1164,N_9939,N_8819);
and UO_1165 (O_1165,N_8659,N_8210);
xor UO_1166 (O_1166,N_8782,N_8774);
or UO_1167 (O_1167,N_9402,N_9692);
xnor UO_1168 (O_1168,N_9065,N_9296);
or UO_1169 (O_1169,N_9392,N_8229);
nand UO_1170 (O_1170,N_8710,N_9737);
nor UO_1171 (O_1171,N_9699,N_9407);
nand UO_1172 (O_1172,N_8824,N_8371);
nand UO_1173 (O_1173,N_8196,N_8708);
nand UO_1174 (O_1174,N_8785,N_8593);
nand UO_1175 (O_1175,N_8974,N_8748);
nor UO_1176 (O_1176,N_8203,N_9688);
nor UO_1177 (O_1177,N_8144,N_9801);
and UO_1178 (O_1178,N_8367,N_8199);
nand UO_1179 (O_1179,N_8998,N_9048);
xnor UO_1180 (O_1180,N_8984,N_8218);
nor UO_1181 (O_1181,N_8840,N_9325);
nand UO_1182 (O_1182,N_8105,N_9952);
xor UO_1183 (O_1183,N_8448,N_8495);
and UO_1184 (O_1184,N_8583,N_9749);
nor UO_1185 (O_1185,N_8266,N_9506);
and UO_1186 (O_1186,N_9258,N_8833);
and UO_1187 (O_1187,N_9166,N_8735);
xnor UO_1188 (O_1188,N_8266,N_9235);
nor UO_1189 (O_1189,N_9190,N_8807);
nor UO_1190 (O_1190,N_8410,N_9980);
or UO_1191 (O_1191,N_9951,N_9729);
nor UO_1192 (O_1192,N_8513,N_9605);
or UO_1193 (O_1193,N_8896,N_8409);
nor UO_1194 (O_1194,N_9716,N_9124);
or UO_1195 (O_1195,N_9291,N_8857);
or UO_1196 (O_1196,N_8691,N_8065);
or UO_1197 (O_1197,N_8223,N_8874);
xnor UO_1198 (O_1198,N_9859,N_8901);
or UO_1199 (O_1199,N_9669,N_8443);
nand UO_1200 (O_1200,N_9517,N_8561);
xor UO_1201 (O_1201,N_9856,N_9806);
or UO_1202 (O_1202,N_8364,N_9098);
or UO_1203 (O_1203,N_8923,N_8179);
nand UO_1204 (O_1204,N_8639,N_8654);
or UO_1205 (O_1205,N_9961,N_8398);
nor UO_1206 (O_1206,N_8727,N_9338);
xnor UO_1207 (O_1207,N_8571,N_8490);
and UO_1208 (O_1208,N_8188,N_9513);
or UO_1209 (O_1209,N_9814,N_9727);
and UO_1210 (O_1210,N_8670,N_8743);
xor UO_1211 (O_1211,N_9339,N_8313);
or UO_1212 (O_1212,N_8467,N_8705);
or UO_1213 (O_1213,N_8565,N_9228);
nor UO_1214 (O_1214,N_8637,N_8224);
xor UO_1215 (O_1215,N_8860,N_8843);
and UO_1216 (O_1216,N_9330,N_9347);
and UO_1217 (O_1217,N_8593,N_8515);
nor UO_1218 (O_1218,N_8464,N_8141);
nand UO_1219 (O_1219,N_9257,N_9625);
nand UO_1220 (O_1220,N_8967,N_9876);
and UO_1221 (O_1221,N_8951,N_9879);
or UO_1222 (O_1222,N_8257,N_8902);
or UO_1223 (O_1223,N_8778,N_8508);
or UO_1224 (O_1224,N_9998,N_8319);
nor UO_1225 (O_1225,N_8185,N_9946);
nor UO_1226 (O_1226,N_8157,N_9171);
or UO_1227 (O_1227,N_8895,N_9305);
nand UO_1228 (O_1228,N_9604,N_8300);
and UO_1229 (O_1229,N_9801,N_9531);
and UO_1230 (O_1230,N_9496,N_8888);
and UO_1231 (O_1231,N_8478,N_9064);
and UO_1232 (O_1232,N_8440,N_9189);
xor UO_1233 (O_1233,N_9366,N_8495);
or UO_1234 (O_1234,N_8832,N_8707);
and UO_1235 (O_1235,N_9400,N_8955);
nor UO_1236 (O_1236,N_9803,N_8289);
nand UO_1237 (O_1237,N_8455,N_8684);
and UO_1238 (O_1238,N_9924,N_8321);
or UO_1239 (O_1239,N_9517,N_9281);
nor UO_1240 (O_1240,N_8029,N_8552);
xor UO_1241 (O_1241,N_9522,N_8533);
nor UO_1242 (O_1242,N_8820,N_9793);
nor UO_1243 (O_1243,N_9296,N_9373);
and UO_1244 (O_1244,N_9796,N_8121);
and UO_1245 (O_1245,N_8007,N_8681);
nand UO_1246 (O_1246,N_8760,N_8271);
and UO_1247 (O_1247,N_9475,N_9144);
or UO_1248 (O_1248,N_9225,N_8795);
or UO_1249 (O_1249,N_8159,N_8250);
nand UO_1250 (O_1250,N_8228,N_9431);
nor UO_1251 (O_1251,N_8040,N_9000);
xnor UO_1252 (O_1252,N_9826,N_9215);
nand UO_1253 (O_1253,N_9699,N_8616);
nor UO_1254 (O_1254,N_8948,N_9646);
xor UO_1255 (O_1255,N_8868,N_8249);
or UO_1256 (O_1256,N_9678,N_8515);
nor UO_1257 (O_1257,N_9896,N_8092);
and UO_1258 (O_1258,N_9948,N_9953);
or UO_1259 (O_1259,N_9595,N_8875);
nand UO_1260 (O_1260,N_9806,N_9913);
and UO_1261 (O_1261,N_9505,N_9864);
nor UO_1262 (O_1262,N_9153,N_9957);
nor UO_1263 (O_1263,N_9365,N_9153);
or UO_1264 (O_1264,N_8007,N_9476);
nand UO_1265 (O_1265,N_8426,N_8776);
nand UO_1266 (O_1266,N_9217,N_9479);
or UO_1267 (O_1267,N_8630,N_9261);
nand UO_1268 (O_1268,N_8563,N_8986);
nand UO_1269 (O_1269,N_9365,N_9989);
nor UO_1270 (O_1270,N_8211,N_9012);
nor UO_1271 (O_1271,N_8085,N_8343);
nor UO_1272 (O_1272,N_8604,N_9981);
and UO_1273 (O_1273,N_9518,N_9895);
nand UO_1274 (O_1274,N_8887,N_8959);
xnor UO_1275 (O_1275,N_9301,N_9076);
nor UO_1276 (O_1276,N_9275,N_9060);
or UO_1277 (O_1277,N_9100,N_9272);
nor UO_1278 (O_1278,N_8859,N_9408);
nor UO_1279 (O_1279,N_8492,N_9966);
nand UO_1280 (O_1280,N_9429,N_8750);
nand UO_1281 (O_1281,N_8311,N_8474);
nor UO_1282 (O_1282,N_9470,N_8229);
nor UO_1283 (O_1283,N_9847,N_9291);
nand UO_1284 (O_1284,N_8246,N_8242);
nand UO_1285 (O_1285,N_8990,N_8958);
and UO_1286 (O_1286,N_8925,N_8166);
xnor UO_1287 (O_1287,N_8942,N_8511);
nand UO_1288 (O_1288,N_8374,N_9379);
nand UO_1289 (O_1289,N_9501,N_8703);
nand UO_1290 (O_1290,N_9583,N_9060);
nor UO_1291 (O_1291,N_8287,N_8508);
and UO_1292 (O_1292,N_8275,N_8309);
nor UO_1293 (O_1293,N_8655,N_8864);
or UO_1294 (O_1294,N_9891,N_8008);
nand UO_1295 (O_1295,N_9420,N_8286);
xor UO_1296 (O_1296,N_9043,N_9404);
nand UO_1297 (O_1297,N_9001,N_8580);
or UO_1298 (O_1298,N_9625,N_8182);
and UO_1299 (O_1299,N_9060,N_9065);
nor UO_1300 (O_1300,N_9298,N_9999);
xnor UO_1301 (O_1301,N_8927,N_8444);
and UO_1302 (O_1302,N_8917,N_8317);
nor UO_1303 (O_1303,N_8215,N_9269);
nor UO_1304 (O_1304,N_9549,N_9484);
nor UO_1305 (O_1305,N_8471,N_8578);
nor UO_1306 (O_1306,N_9158,N_9536);
and UO_1307 (O_1307,N_9168,N_8861);
nand UO_1308 (O_1308,N_9740,N_8616);
nand UO_1309 (O_1309,N_9825,N_8265);
nor UO_1310 (O_1310,N_8285,N_9616);
nand UO_1311 (O_1311,N_8208,N_9032);
nand UO_1312 (O_1312,N_9877,N_9463);
nor UO_1313 (O_1313,N_9787,N_8816);
xor UO_1314 (O_1314,N_8577,N_8174);
nor UO_1315 (O_1315,N_8286,N_9439);
and UO_1316 (O_1316,N_8225,N_9083);
nor UO_1317 (O_1317,N_8980,N_9094);
nand UO_1318 (O_1318,N_8885,N_9151);
and UO_1319 (O_1319,N_8829,N_8565);
nor UO_1320 (O_1320,N_8658,N_9643);
xor UO_1321 (O_1321,N_8524,N_8153);
nor UO_1322 (O_1322,N_8652,N_9624);
and UO_1323 (O_1323,N_9182,N_8649);
xor UO_1324 (O_1324,N_9299,N_8588);
nand UO_1325 (O_1325,N_9781,N_8399);
nor UO_1326 (O_1326,N_8769,N_8468);
or UO_1327 (O_1327,N_8352,N_8306);
xor UO_1328 (O_1328,N_9276,N_8075);
nand UO_1329 (O_1329,N_9760,N_9845);
nor UO_1330 (O_1330,N_8951,N_9817);
or UO_1331 (O_1331,N_8523,N_9572);
nor UO_1332 (O_1332,N_8770,N_8402);
or UO_1333 (O_1333,N_8385,N_8059);
and UO_1334 (O_1334,N_8396,N_9834);
and UO_1335 (O_1335,N_8099,N_8063);
nor UO_1336 (O_1336,N_8875,N_8729);
and UO_1337 (O_1337,N_9969,N_9730);
xnor UO_1338 (O_1338,N_9185,N_8152);
nor UO_1339 (O_1339,N_8328,N_8175);
nor UO_1340 (O_1340,N_8176,N_9904);
xor UO_1341 (O_1341,N_8288,N_9200);
or UO_1342 (O_1342,N_8901,N_8431);
and UO_1343 (O_1343,N_9158,N_9648);
and UO_1344 (O_1344,N_9611,N_9099);
nor UO_1345 (O_1345,N_8803,N_9928);
nand UO_1346 (O_1346,N_8039,N_9622);
nand UO_1347 (O_1347,N_9648,N_8728);
nor UO_1348 (O_1348,N_9683,N_8086);
and UO_1349 (O_1349,N_8057,N_9879);
and UO_1350 (O_1350,N_9890,N_8470);
or UO_1351 (O_1351,N_8726,N_8448);
or UO_1352 (O_1352,N_9875,N_8630);
nor UO_1353 (O_1353,N_9140,N_9991);
nor UO_1354 (O_1354,N_9209,N_9921);
or UO_1355 (O_1355,N_9371,N_9383);
and UO_1356 (O_1356,N_8196,N_9052);
or UO_1357 (O_1357,N_9875,N_9030);
nand UO_1358 (O_1358,N_9111,N_9829);
nand UO_1359 (O_1359,N_9116,N_8144);
and UO_1360 (O_1360,N_9227,N_8568);
nor UO_1361 (O_1361,N_8324,N_9822);
and UO_1362 (O_1362,N_9219,N_8736);
nand UO_1363 (O_1363,N_8178,N_9069);
or UO_1364 (O_1364,N_8111,N_8619);
xnor UO_1365 (O_1365,N_9532,N_8272);
and UO_1366 (O_1366,N_8656,N_8408);
nand UO_1367 (O_1367,N_8326,N_9393);
nor UO_1368 (O_1368,N_9135,N_9637);
and UO_1369 (O_1369,N_9031,N_9217);
xor UO_1370 (O_1370,N_8050,N_9603);
or UO_1371 (O_1371,N_8111,N_8476);
xnor UO_1372 (O_1372,N_8761,N_8378);
or UO_1373 (O_1373,N_9756,N_9387);
nand UO_1374 (O_1374,N_8645,N_9156);
or UO_1375 (O_1375,N_8154,N_8257);
and UO_1376 (O_1376,N_9139,N_8557);
and UO_1377 (O_1377,N_8763,N_9785);
nor UO_1378 (O_1378,N_9999,N_9688);
and UO_1379 (O_1379,N_9216,N_8044);
nand UO_1380 (O_1380,N_8677,N_9316);
xnor UO_1381 (O_1381,N_9846,N_8761);
or UO_1382 (O_1382,N_9813,N_9736);
nand UO_1383 (O_1383,N_8566,N_9185);
nand UO_1384 (O_1384,N_8610,N_9409);
and UO_1385 (O_1385,N_8249,N_8026);
and UO_1386 (O_1386,N_9065,N_9910);
and UO_1387 (O_1387,N_8924,N_8381);
and UO_1388 (O_1388,N_9608,N_8718);
xnor UO_1389 (O_1389,N_9343,N_8190);
xor UO_1390 (O_1390,N_8439,N_9114);
and UO_1391 (O_1391,N_9649,N_8365);
or UO_1392 (O_1392,N_8596,N_8445);
nand UO_1393 (O_1393,N_9021,N_9538);
xor UO_1394 (O_1394,N_9022,N_9822);
nand UO_1395 (O_1395,N_8356,N_8308);
nand UO_1396 (O_1396,N_8457,N_9338);
and UO_1397 (O_1397,N_9752,N_9853);
or UO_1398 (O_1398,N_9685,N_8105);
nand UO_1399 (O_1399,N_9880,N_9667);
or UO_1400 (O_1400,N_8176,N_9244);
or UO_1401 (O_1401,N_9619,N_8402);
nor UO_1402 (O_1402,N_8986,N_9400);
and UO_1403 (O_1403,N_9907,N_8065);
nand UO_1404 (O_1404,N_9445,N_8915);
nand UO_1405 (O_1405,N_9138,N_8878);
and UO_1406 (O_1406,N_9252,N_8411);
nor UO_1407 (O_1407,N_8884,N_9651);
and UO_1408 (O_1408,N_9740,N_8551);
or UO_1409 (O_1409,N_9360,N_9391);
or UO_1410 (O_1410,N_8795,N_9814);
and UO_1411 (O_1411,N_9412,N_9686);
nor UO_1412 (O_1412,N_8007,N_9304);
nor UO_1413 (O_1413,N_8158,N_9325);
nand UO_1414 (O_1414,N_9346,N_8854);
and UO_1415 (O_1415,N_8074,N_8225);
or UO_1416 (O_1416,N_9255,N_9580);
and UO_1417 (O_1417,N_9850,N_8644);
and UO_1418 (O_1418,N_9904,N_9913);
and UO_1419 (O_1419,N_9407,N_8768);
and UO_1420 (O_1420,N_8775,N_9291);
nand UO_1421 (O_1421,N_9260,N_9196);
and UO_1422 (O_1422,N_9346,N_8485);
nand UO_1423 (O_1423,N_9177,N_8301);
nor UO_1424 (O_1424,N_9824,N_8778);
xor UO_1425 (O_1425,N_8007,N_9105);
nor UO_1426 (O_1426,N_8849,N_9074);
or UO_1427 (O_1427,N_8882,N_9865);
nor UO_1428 (O_1428,N_8165,N_8064);
nor UO_1429 (O_1429,N_8429,N_8086);
nor UO_1430 (O_1430,N_8752,N_8472);
nand UO_1431 (O_1431,N_9649,N_8839);
xor UO_1432 (O_1432,N_9484,N_9726);
nand UO_1433 (O_1433,N_8663,N_9721);
nand UO_1434 (O_1434,N_9541,N_8382);
nand UO_1435 (O_1435,N_9432,N_9673);
xor UO_1436 (O_1436,N_8452,N_8111);
or UO_1437 (O_1437,N_8322,N_8604);
nor UO_1438 (O_1438,N_8870,N_9433);
or UO_1439 (O_1439,N_9848,N_9667);
nand UO_1440 (O_1440,N_9425,N_9159);
nor UO_1441 (O_1441,N_9544,N_8573);
or UO_1442 (O_1442,N_9896,N_8736);
or UO_1443 (O_1443,N_8671,N_8976);
and UO_1444 (O_1444,N_8857,N_8873);
and UO_1445 (O_1445,N_9222,N_8032);
nand UO_1446 (O_1446,N_9434,N_9678);
and UO_1447 (O_1447,N_9331,N_9819);
and UO_1448 (O_1448,N_9870,N_9292);
or UO_1449 (O_1449,N_8108,N_9790);
or UO_1450 (O_1450,N_9905,N_9504);
or UO_1451 (O_1451,N_9653,N_9337);
xnor UO_1452 (O_1452,N_9135,N_8984);
nor UO_1453 (O_1453,N_9117,N_9289);
nand UO_1454 (O_1454,N_9484,N_9308);
xor UO_1455 (O_1455,N_8898,N_8309);
or UO_1456 (O_1456,N_9461,N_9202);
xnor UO_1457 (O_1457,N_8859,N_9753);
nor UO_1458 (O_1458,N_9792,N_8343);
nor UO_1459 (O_1459,N_8653,N_8939);
or UO_1460 (O_1460,N_9557,N_9336);
and UO_1461 (O_1461,N_9422,N_8900);
nand UO_1462 (O_1462,N_9421,N_8357);
xor UO_1463 (O_1463,N_8866,N_9090);
nor UO_1464 (O_1464,N_8811,N_8665);
nand UO_1465 (O_1465,N_9895,N_8148);
nand UO_1466 (O_1466,N_9628,N_9502);
nand UO_1467 (O_1467,N_8849,N_9046);
and UO_1468 (O_1468,N_9940,N_8125);
and UO_1469 (O_1469,N_8065,N_9789);
or UO_1470 (O_1470,N_9363,N_9986);
nor UO_1471 (O_1471,N_9742,N_9094);
or UO_1472 (O_1472,N_9336,N_9586);
or UO_1473 (O_1473,N_8989,N_8139);
nand UO_1474 (O_1474,N_9070,N_8968);
nand UO_1475 (O_1475,N_8443,N_9744);
nand UO_1476 (O_1476,N_8839,N_9736);
and UO_1477 (O_1477,N_8629,N_9794);
or UO_1478 (O_1478,N_8890,N_8408);
xnor UO_1479 (O_1479,N_9185,N_8576);
nor UO_1480 (O_1480,N_9594,N_9474);
and UO_1481 (O_1481,N_9646,N_8342);
or UO_1482 (O_1482,N_9538,N_9817);
or UO_1483 (O_1483,N_9561,N_9343);
or UO_1484 (O_1484,N_9925,N_8409);
nand UO_1485 (O_1485,N_8638,N_8530);
nor UO_1486 (O_1486,N_8218,N_8828);
xnor UO_1487 (O_1487,N_8171,N_9456);
and UO_1488 (O_1488,N_8598,N_9034);
nand UO_1489 (O_1489,N_8742,N_8712);
and UO_1490 (O_1490,N_8196,N_8052);
and UO_1491 (O_1491,N_8765,N_9889);
and UO_1492 (O_1492,N_9340,N_9065);
or UO_1493 (O_1493,N_8720,N_9397);
nor UO_1494 (O_1494,N_8463,N_8298);
and UO_1495 (O_1495,N_8125,N_8034);
and UO_1496 (O_1496,N_9138,N_8593);
and UO_1497 (O_1497,N_8239,N_9913);
xnor UO_1498 (O_1498,N_8473,N_9736);
or UO_1499 (O_1499,N_9612,N_8224);
endmodule