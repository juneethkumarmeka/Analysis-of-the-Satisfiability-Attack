module basic_1000_10000_1500_2_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5006,N_5010,N_5012,N_5013,N_5014,N_5015,N_5017,N_5018,N_5019,N_5020,N_5022,N_5023,N_5024,N_5025,N_5026,N_5028,N_5029,N_5030,N_5031,N_5033,N_5034,N_5037,N_5038,N_5039,N_5040,N_5041,N_5043,N_5046,N_5048,N_5049,N_5050,N_5052,N_5053,N_5054,N_5055,N_5057,N_5058,N_5059,N_5061,N_5062,N_5065,N_5072,N_5083,N_5084,N_5085,N_5086,N_5087,N_5090,N_5091,N_5092,N_5094,N_5095,N_5103,N_5107,N_5108,N_5110,N_5112,N_5113,N_5114,N_5117,N_5119,N_5125,N_5126,N_5127,N_5129,N_5131,N_5133,N_5136,N_5137,N_5140,N_5145,N_5146,N_5147,N_5148,N_5149,N_5151,N_5153,N_5154,N_5155,N_5156,N_5158,N_5162,N_5163,N_5164,N_5167,N_5168,N_5169,N_5170,N_5171,N_5173,N_5174,N_5176,N_5178,N_5181,N_5183,N_5184,N_5185,N_5186,N_5187,N_5189,N_5191,N_5192,N_5193,N_5197,N_5199,N_5201,N_5203,N_5206,N_5207,N_5208,N_5209,N_5211,N_5213,N_5214,N_5215,N_5216,N_5219,N_5221,N_5222,N_5223,N_5224,N_5225,N_5228,N_5230,N_5231,N_5233,N_5235,N_5237,N_5238,N_5245,N_5246,N_5249,N_5250,N_5251,N_5254,N_5256,N_5258,N_5260,N_5261,N_5263,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5272,N_5273,N_5274,N_5275,N_5276,N_5278,N_5279,N_5281,N_5282,N_5283,N_5285,N_5289,N_5290,N_5291,N_5293,N_5295,N_5296,N_5300,N_5301,N_5302,N_5303,N_5304,N_5307,N_5308,N_5309,N_5310,N_5311,N_5313,N_5317,N_5319,N_5320,N_5321,N_5322,N_5323,N_5326,N_5327,N_5330,N_5335,N_5336,N_5338,N_5342,N_5343,N_5344,N_5346,N_5347,N_5348,N_5350,N_5351,N_5352,N_5356,N_5358,N_5359,N_5360,N_5361,N_5362,N_5364,N_5365,N_5366,N_5367,N_5370,N_5371,N_5374,N_5376,N_5379,N_5381,N_5385,N_5386,N_5387,N_5389,N_5390,N_5392,N_5393,N_5394,N_5396,N_5397,N_5398,N_5399,N_5402,N_5406,N_5407,N_5409,N_5410,N_5411,N_5412,N_5414,N_5415,N_5417,N_5418,N_5419,N_5422,N_5423,N_5424,N_5427,N_5429,N_5430,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5445,N_5446,N_5447,N_5448,N_5449,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5459,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5469,N_5470,N_5471,N_5472,N_5474,N_5475,N_5477,N_5478,N_5479,N_5481,N_5483,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5504,N_5506,N_5507,N_5508,N_5509,N_5512,N_5516,N_5517,N_5518,N_5519,N_5521,N_5522,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5537,N_5538,N_5540,N_5542,N_5543,N_5545,N_5548,N_5550,N_5552,N_5554,N_5557,N_5559,N_5560,N_5564,N_5565,N_5566,N_5568,N_5569,N_5570,N_5572,N_5573,N_5575,N_5579,N_5580,N_5581,N_5582,N_5586,N_5589,N_5591,N_5594,N_5596,N_5598,N_5599,N_5600,N_5601,N_5602,N_5604,N_5605,N_5607,N_5608,N_5610,N_5612,N_5614,N_5616,N_5618,N_5619,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5630,N_5631,N_5632,N_5633,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5642,N_5643,N_5645,N_5646,N_5649,N_5651,N_5653,N_5654,N_5655,N_5656,N_5658,N_5659,N_5660,N_5666,N_5669,N_5670,N_5671,N_5673,N_5678,N_5679,N_5680,N_5681,N_5683,N_5684,N_5685,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5695,N_5698,N_5699,N_5700,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5710,N_5713,N_5714,N_5715,N_5716,N_5717,N_5720,N_5721,N_5722,N_5727,N_5729,N_5731,N_5733,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5745,N_5749,N_5750,N_5751,N_5752,N_5753,N_5755,N_5756,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5767,N_5769,N_5771,N_5773,N_5774,N_5776,N_5779,N_5781,N_5782,N_5785,N_5786,N_5788,N_5791,N_5793,N_5794,N_5797,N_5798,N_5800,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5812,N_5813,N_5814,N_5816,N_5819,N_5820,N_5822,N_5823,N_5824,N_5826,N_5828,N_5830,N_5831,N_5832,N_5836,N_5837,N_5838,N_5839,N_5840,N_5842,N_5844,N_5845,N_5847,N_5848,N_5850,N_5851,N_5852,N_5859,N_5860,N_5861,N_5862,N_5864,N_5866,N_5867,N_5868,N_5869,N_5870,N_5872,N_5873,N_5874,N_5875,N_5876,N_5878,N_5881,N_5883,N_5886,N_5887,N_5889,N_5891,N_5895,N_5896,N_5897,N_5899,N_5900,N_5901,N_5903,N_5904,N_5905,N_5908,N_5909,N_5914,N_5915,N_5916,N_5920,N_5921,N_5924,N_5925,N_5926,N_5927,N_5933,N_5938,N_5940,N_5941,N_5942,N_5944,N_5947,N_5948,N_5949,N_5950,N_5952,N_5953,N_5954,N_5956,N_5957,N_5958,N_5959,N_5963,N_5964,N_5965,N_5967,N_5968,N_5969,N_5971,N_5972,N_5973,N_5976,N_5978,N_5980,N_5981,N_5982,N_5983,N_5984,N_5986,N_5988,N_5994,N_5996,N_5998,N_6000,N_6001,N_6002,N_6004,N_6005,N_6006,N_6007,N_6008,N_6010,N_6012,N_6015,N_6016,N_6018,N_6019,N_6020,N_6022,N_6025,N_6028,N_6029,N_6031,N_6032,N_6033,N_6035,N_6036,N_6039,N_6040,N_6042,N_6043,N_6044,N_6046,N_6049,N_6052,N_6053,N_6055,N_6057,N_6058,N_6060,N_6063,N_6064,N_6065,N_6068,N_6069,N_6070,N_6071,N_6073,N_6074,N_6075,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6086,N_6087,N_6092,N_6093,N_6094,N_6096,N_6097,N_6098,N_6100,N_6101,N_6102,N_6103,N_6106,N_6108,N_6109,N_6110,N_6113,N_6114,N_6115,N_6117,N_6119,N_6120,N_6123,N_6125,N_6127,N_6128,N_6130,N_6131,N_6133,N_6134,N_6135,N_6137,N_6138,N_6143,N_6145,N_6146,N_6148,N_6150,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6161,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6172,N_6173,N_6174,N_6176,N_6177,N_6178,N_6182,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6193,N_6194,N_6195,N_6200,N_6202,N_6203,N_6204,N_6207,N_6208,N_6209,N_6210,N_6212,N_6213,N_6217,N_6218,N_6219,N_6220,N_6222,N_6224,N_6225,N_6226,N_6227,N_6228,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6239,N_6243,N_6244,N_6245,N_6246,N_6249,N_6251,N_6252,N_6253,N_6254,N_6259,N_6260,N_6261,N_6262,N_6265,N_6266,N_6268,N_6269,N_6272,N_6276,N_6277,N_6279,N_6280,N_6283,N_6284,N_6285,N_6286,N_6289,N_6292,N_6293,N_6295,N_6297,N_6298,N_6300,N_6301,N_6302,N_6304,N_6307,N_6312,N_6313,N_6314,N_6318,N_6320,N_6321,N_6324,N_6325,N_6326,N_6331,N_6332,N_6333,N_6334,N_6336,N_6337,N_6338,N_6341,N_6342,N_6343,N_6345,N_6346,N_6348,N_6349,N_6351,N_6352,N_6353,N_6355,N_6360,N_6361,N_6362,N_6363,N_6366,N_6367,N_6368,N_6369,N_6373,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6387,N_6389,N_6392,N_6393,N_6394,N_6397,N_6398,N_6400,N_6401,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6411,N_6412,N_6413,N_6416,N_6418,N_6421,N_6422,N_6423,N_6427,N_6429,N_6430,N_6432,N_6435,N_6436,N_6437,N_6443,N_6444,N_6445,N_6446,N_6447,N_6451,N_6452,N_6453,N_6454,N_6455,N_6458,N_6459,N_6460,N_6464,N_6465,N_6466,N_6467,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6477,N_6478,N_6483,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6494,N_6496,N_6497,N_6500,N_6501,N_6504,N_6505,N_6506,N_6510,N_6512,N_6514,N_6515,N_6517,N_6518,N_6519,N_6520,N_6521,N_6523,N_6524,N_6526,N_6527,N_6529,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6552,N_6553,N_6554,N_6557,N_6560,N_6564,N_6565,N_6571,N_6574,N_6575,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6586,N_6588,N_6589,N_6590,N_6592,N_6594,N_6595,N_6597,N_6598,N_6600,N_6604,N_6605,N_6607,N_6608,N_6609,N_6613,N_6615,N_6616,N_6617,N_6619,N_6620,N_6621,N_6622,N_6624,N_6626,N_6628,N_6632,N_6633,N_6638,N_6639,N_6641,N_6646,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6658,N_6659,N_6660,N_6662,N_6666,N_6668,N_6671,N_6674,N_6675,N_6676,N_6678,N_6679,N_6681,N_6683,N_6684,N_6687,N_6690,N_6691,N_6694,N_6696,N_6697,N_6700,N_6702,N_6704,N_6706,N_6707,N_6709,N_6710,N_6714,N_6716,N_6718,N_6719,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6752,N_6753,N_6755,N_6757,N_6759,N_6760,N_6762,N_6763,N_6764,N_6765,N_6768,N_6769,N_6770,N_6772,N_6774,N_6777,N_6778,N_6780,N_6781,N_6782,N_6785,N_6787,N_6789,N_6790,N_6791,N_6792,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6803,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6813,N_6814,N_6815,N_6816,N_6818,N_6819,N_6823,N_6824,N_6827,N_6828,N_6829,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6855,N_6858,N_6860,N_6862,N_6864,N_6865,N_6866,N_6867,N_6868,N_6870,N_6872,N_6873,N_6875,N_6878,N_6879,N_6882,N_6885,N_6889,N_6891,N_6892,N_6893,N_6895,N_6897,N_6899,N_6901,N_6902,N_6903,N_6904,N_6906,N_6907,N_6908,N_6909,N_6910,N_6913,N_6915,N_6919,N_6920,N_6921,N_6922,N_6925,N_6927,N_6930,N_6933,N_6936,N_6940,N_6942,N_6943,N_6947,N_6948,N_6951,N_6952,N_6953,N_6956,N_6960,N_6961,N_6963,N_6964,N_6965,N_6967,N_6969,N_6971,N_6972,N_6973,N_6975,N_6977,N_6978,N_6979,N_6980,N_6981,N_6985,N_6986,N_6987,N_6989,N_6991,N_6992,N_6993,N_6995,N_6996,N_6997,N_6998,N_7002,N_7004,N_7006,N_7007,N_7008,N_7011,N_7014,N_7015,N_7017,N_7020,N_7021,N_7022,N_7025,N_7026,N_7028,N_7029,N_7030,N_7031,N_7032,N_7034,N_7039,N_7041,N_7042,N_7044,N_7045,N_7046,N_7050,N_7051,N_7053,N_7054,N_7057,N_7058,N_7059,N_7061,N_7062,N_7063,N_7064,N_7065,N_7067,N_7069,N_7070,N_7072,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7082,N_7084,N_7085,N_7086,N_7087,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7106,N_7110,N_7112,N_7114,N_7115,N_7117,N_7123,N_7125,N_7126,N_7131,N_7132,N_7133,N_7135,N_7137,N_7138,N_7140,N_7141,N_7142,N_7143,N_7146,N_7147,N_7151,N_7153,N_7155,N_7156,N_7157,N_7158,N_7159,N_7163,N_7164,N_7165,N_7167,N_7168,N_7170,N_7172,N_7174,N_7175,N_7176,N_7182,N_7184,N_7185,N_7187,N_7188,N_7190,N_7192,N_7193,N_7196,N_7197,N_7199,N_7200,N_7204,N_7205,N_7206,N_7211,N_7217,N_7218,N_7219,N_7220,N_7223,N_7224,N_7225,N_7226,N_7227,N_7230,N_7231,N_7233,N_7234,N_7235,N_7237,N_7239,N_7241,N_7242,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7264,N_7265,N_7269,N_7270,N_7271,N_7272,N_7274,N_7276,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7285,N_7286,N_7289,N_7291,N_7292,N_7293,N_7294,N_7297,N_7298,N_7299,N_7302,N_7303,N_7305,N_7309,N_7311,N_7312,N_7313,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7329,N_7331,N_7334,N_7337,N_7338,N_7339,N_7342,N_7343,N_7344,N_7347,N_7349,N_7351,N_7352,N_7354,N_7355,N_7356,N_7358,N_7359,N_7363,N_7364,N_7365,N_7366,N_7369,N_7370,N_7371,N_7376,N_7378,N_7379,N_7380,N_7381,N_7385,N_7389,N_7391,N_7392,N_7394,N_7396,N_7400,N_7401,N_7402,N_7403,N_7405,N_7408,N_7409,N_7411,N_7412,N_7413,N_7414,N_7415,N_7417,N_7419,N_7420,N_7421,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7433,N_7435,N_7436,N_7440,N_7441,N_7442,N_7444,N_7445,N_7448,N_7450,N_7451,N_7452,N_7453,N_7455,N_7459,N_7460,N_7464,N_7465,N_7466,N_7467,N_7468,N_7471,N_7472,N_7473,N_7475,N_7477,N_7479,N_7480,N_7482,N_7483,N_7484,N_7485,N_7486,N_7488,N_7491,N_7494,N_7496,N_7497,N_7499,N_7502,N_7503,N_7504,N_7508,N_7509,N_7511,N_7514,N_7515,N_7516,N_7517,N_7519,N_7522,N_7524,N_7525,N_7526,N_7527,N_7528,N_7530,N_7534,N_7535,N_7536,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7548,N_7549,N_7550,N_7551,N_7552,N_7554,N_7555,N_7559,N_7560,N_7561,N_7562,N_7564,N_7566,N_7567,N_7570,N_7572,N_7574,N_7580,N_7582,N_7585,N_7586,N_7587,N_7588,N_7589,N_7593,N_7597,N_7598,N_7599,N_7602,N_7604,N_7605,N_7606,N_7608,N_7612,N_7613,N_7614,N_7615,N_7617,N_7618,N_7619,N_7621,N_7622,N_7623,N_7626,N_7627,N_7628,N_7631,N_7633,N_7634,N_7636,N_7638,N_7639,N_7641,N_7642,N_7643,N_7645,N_7649,N_7650,N_7652,N_7653,N_7655,N_7659,N_7662,N_7663,N_7664,N_7666,N_7667,N_7670,N_7671,N_7672,N_7673,N_7676,N_7677,N_7679,N_7681,N_7682,N_7683,N_7684,N_7685,N_7687,N_7688,N_7689,N_7690,N_7692,N_7693,N_7695,N_7696,N_7697,N_7698,N_7700,N_7701,N_7702,N_7703,N_7705,N_7706,N_7708,N_7709,N_7710,N_7714,N_7716,N_7717,N_7718,N_7719,N_7720,N_7722,N_7723,N_7728,N_7729,N_7733,N_7734,N_7735,N_7738,N_7739,N_7740,N_7742,N_7743,N_7744,N_7746,N_7747,N_7748,N_7750,N_7753,N_7755,N_7756,N_7757,N_7760,N_7761,N_7764,N_7765,N_7766,N_7767,N_7771,N_7772,N_7774,N_7775,N_7776,N_7777,N_7779,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7794,N_7795,N_7796,N_7797,N_7801,N_7802,N_7803,N_7804,N_7806,N_7807,N_7809,N_7810,N_7811,N_7813,N_7814,N_7815,N_7816,N_7818,N_7821,N_7822,N_7823,N_7827,N_7828,N_7829,N_7833,N_7834,N_7835,N_7837,N_7838,N_7840,N_7841,N_7843,N_7844,N_7846,N_7847,N_7849,N_7853,N_7854,N_7855,N_7857,N_7859,N_7860,N_7861,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7872,N_7873,N_7877,N_7878,N_7879,N_7880,N_7883,N_7884,N_7888,N_7889,N_7891,N_7892,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7906,N_7908,N_7909,N_7910,N_7912,N_7915,N_7916,N_7917,N_7920,N_7922,N_7923,N_7924,N_7926,N_7927,N_7928,N_7930,N_7931,N_7933,N_7935,N_7936,N_7939,N_7940,N_7941,N_7942,N_7948,N_7949,N_7950,N_7951,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7967,N_7968,N_7969,N_7970,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7983,N_7986,N_7987,N_7988,N_7989,N_7991,N_7992,N_7993,N_7994,N_7995,N_7997,N_7998,N_7999,N_8000,N_8001,N_8003,N_8004,N_8007,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8017,N_8018,N_8019,N_8020,N_8022,N_8026,N_8031,N_8034,N_8035,N_8038,N_8039,N_8040,N_8044,N_8045,N_8046,N_8048,N_8050,N_8054,N_8055,N_8058,N_8059,N_8060,N_8061,N_8062,N_8066,N_8067,N_8070,N_8071,N_8074,N_8077,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8088,N_8089,N_8092,N_8093,N_8095,N_8099,N_8101,N_8102,N_8105,N_8107,N_8108,N_8109,N_8114,N_8115,N_8118,N_8119,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8131,N_8135,N_8136,N_8138,N_8142,N_8143,N_8145,N_8146,N_8148,N_8150,N_8151,N_8152,N_8153,N_8157,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8170,N_8171,N_8172,N_8173,N_8176,N_8178,N_8180,N_8182,N_8184,N_8185,N_8187,N_8188,N_8189,N_8190,N_8191,N_8193,N_8194,N_8196,N_8198,N_8199,N_8201,N_8202,N_8204,N_8206,N_8207,N_8209,N_8211,N_8213,N_8214,N_8216,N_8217,N_8220,N_8221,N_8222,N_8226,N_8229,N_8230,N_8231,N_8232,N_8233,N_8235,N_8236,N_8238,N_8244,N_8248,N_8249,N_8250,N_8252,N_8253,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8265,N_8266,N_8267,N_8268,N_8271,N_8272,N_8273,N_8274,N_8275,N_8277,N_8278,N_8280,N_8281,N_8282,N_8284,N_8285,N_8287,N_8288,N_8289,N_8292,N_8295,N_8296,N_8297,N_8298,N_8299,N_8301,N_8302,N_8304,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8314,N_8315,N_8317,N_8321,N_8322,N_8325,N_8326,N_8329,N_8330,N_8333,N_8335,N_8337,N_8339,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8354,N_8356,N_8357,N_8359,N_8361,N_8362,N_8363,N_8364,N_8366,N_8368,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8391,N_8393,N_8395,N_8397,N_8398,N_8400,N_8401,N_8402,N_8403,N_8404,N_8406,N_8409,N_8411,N_8414,N_8416,N_8418,N_8419,N_8420,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8433,N_8434,N_8435,N_8436,N_8437,N_8441,N_8442,N_8443,N_8444,N_8448,N_8449,N_8455,N_8458,N_8460,N_8463,N_8464,N_8465,N_8467,N_8468,N_8471,N_8472,N_8473,N_8474,N_8475,N_8477,N_8478,N_8479,N_8481,N_8482,N_8485,N_8486,N_8487,N_8490,N_8491,N_8492,N_8493,N_8494,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8503,N_8504,N_8505,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8524,N_8525,N_8526,N_8529,N_8530,N_8531,N_8533,N_8534,N_8536,N_8538,N_8539,N_8540,N_8544,N_8545,N_8549,N_8551,N_8552,N_8554,N_8558,N_8561,N_8563,N_8564,N_8565,N_8566,N_8568,N_8571,N_8572,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8583,N_8584,N_8586,N_8587,N_8588,N_8591,N_8594,N_8596,N_8597,N_8598,N_8599,N_8600,N_8603,N_8604,N_8606,N_8608,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8617,N_8618,N_8619,N_8623,N_8625,N_8626,N_8628,N_8629,N_8630,N_8631,N_8632,N_8635,N_8636,N_8637,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8649,N_8652,N_8654,N_8655,N_8657,N_8658,N_8662,N_8664,N_8665,N_8667,N_8669,N_8672,N_8675,N_8676,N_8680,N_8681,N_8684,N_8686,N_8691,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8705,N_8707,N_8710,N_8711,N_8712,N_8715,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8736,N_8737,N_8738,N_8739,N_8743,N_8744,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8754,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8767,N_8768,N_8769,N_8770,N_8771,N_8773,N_8774,N_8777,N_8778,N_8780,N_8781,N_8784,N_8785,N_8786,N_8787,N_8789,N_8790,N_8791,N_8792,N_8794,N_8797,N_8799,N_8800,N_8801,N_8803,N_8804,N_8807,N_8810,N_8812,N_8814,N_8815,N_8816,N_8817,N_8819,N_8820,N_8821,N_8824,N_8825,N_8829,N_8831,N_8832,N_8833,N_8834,N_8836,N_8838,N_8840,N_8841,N_8842,N_8844,N_8845,N_8846,N_8850,N_8852,N_8854,N_8855,N_8856,N_8858,N_8859,N_8860,N_8862,N_8863,N_8864,N_8865,N_8868,N_8869,N_8870,N_8872,N_8874,N_8875,N_8876,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8885,N_8886,N_8887,N_8889,N_8890,N_8892,N_8894,N_8895,N_8896,N_8897,N_8899,N_8900,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8909,N_8910,N_8911,N_8912,N_8915,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8935,N_8936,N_8939,N_8940,N_8941,N_8943,N_8944,N_8946,N_8947,N_8948,N_8950,N_8952,N_8953,N_8955,N_8956,N_8957,N_8958,N_8959,N_8962,N_8963,N_8964,N_8965,N_8966,N_8968,N_8971,N_8975,N_8977,N_8979,N_8982,N_8983,N_8984,N_8985,N_8987,N_8992,N_8993,N_8994,N_8995,N_9000,N_9005,N_9007,N_9008,N_9010,N_9011,N_9012,N_9013,N_9015,N_9017,N_9018,N_9019,N_9023,N_9024,N_9025,N_9026,N_9027,N_9029,N_9031,N_9033,N_9035,N_9036,N_9037,N_9039,N_9041,N_9043,N_9045,N_9046,N_9047,N_9051,N_9052,N_9053,N_9054,N_9056,N_9057,N_9058,N_9059,N_9064,N_9065,N_9067,N_9069,N_9072,N_9074,N_9075,N_9076,N_9079,N_9080,N_9081,N_9084,N_9086,N_9087,N_9089,N_9090,N_9092,N_9094,N_9095,N_9099,N_9100,N_9104,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9113,N_9119,N_9120,N_9124,N_9125,N_9127,N_9133,N_9135,N_9136,N_9139,N_9140,N_9144,N_9146,N_9147,N_9148,N_9149,N_9150,N_9152,N_9154,N_9155,N_9157,N_9159,N_9160,N_9161,N_9163,N_9164,N_9165,N_9169,N_9171,N_9173,N_9174,N_9176,N_9177,N_9180,N_9181,N_9182,N_9184,N_9185,N_9187,N_9188,N_9189,N_9190,N_9192,N_9193,N_9195,N_9197,N_9199,N_9200,N_9202,N_9203,N_9205,N_9206,N_9209,N_9212,N_9214,N_9215,N_9216,N_9218,N_9219,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9233,N_9234,N_9235,N_9236,N_9239,N_9240,N_9241,N_9243,N_9249,N_9250,N_9252,N_9253,N_9256,N_9258,N_9261,N_9262,N_9264,N_9265,N_9266,N_9267,N_9272,N_9274,N_9275,N_9276,N_9281,N_9282,N_9283,N_9284,N_9286,N_9287,N_9290,N_9295,N_9296,N_9298,N_9300,N_9303,N_9304,N_9305,N_9308,N_9310,N_9311,N_9315,N_9317,N_9319,N_9320,N_9321,N_9323,N_9324,N_9325,N_9326,N_9327,N_9330,N_9331,N_9332,N_9333,N_9334,N_9336,N_9337,N_9338,N_9339,N_9341,N_9342,N_9343,N_9344,N_9345,N_9348,N_9351,N_9356,N_9357,N_9358,N_9359,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9369,N_9370,N_9371,N_9372,N_9374,N_9379,N_9382,N_9383,N_9385,N_9386,N_9388,N_9391,N_9392,N_9393,N_9394,N_9395,N_9399,N_9400,N_9401,N_9404,N_9408,N_9412,N_9413,N_9414,N_9415,N_9417,N_9418,N_9420,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9433,N_9434,N_9436,N_9437,N_9438,N_9439,N_9444,N_9445,N_9446,N_9447,N_9450,N_9451,N_9453,N_9454,N_9455,N_9457,N_9458,N_9461,N_9462,N_9463,N_9464,N_9469,N_9470,N_9471,N_9472,N_9475,N_9476,N_9478,N_9480,N_9481,N_9482,N_9483,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9494,N_9495,N_9496,N_9499,N_9503,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9515,N_9516,N_9517,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9536,N_9538,N_9540,N_9542,N_9543,N_9544,N_9546,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9557,N_9558,N_9559,N_9560,N_9562,N_9568,N_9569,N_9571,N_9572,N_9574,N_9575,N_9579,N_9583,N_9584,N_9586,N_9587,N_9591,N_9592,N_9593,N_9595,N_9596,N_9597,N_9601,N_9603,N_9605,N_9608,N_9612,N_9613,N_9614,N_9616,N_9618,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9629,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9640,N_9641,N_9642,N_9646,N_9647,N_9648,N_9649,N_9651,N_9653,N_9655,N_9656,N_9657,N_9659,N_9661,N_9666,N_9668,N_9669,N_9671,N_9672,N_9673,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9683,N_9685,N_9686,N_9688,N_9689,N_9690,N_9691,N_9693,N_9694,N_9695,N_9699,N_9700,N_9701,N_9702,N_9705,N_9706,N_9708,N_9711,N_9713,N_9714,N_9715,N_9716,N_9717,N_9719,N_9721,N_9722,N_9724,N_9726,N_9729,N_9734,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9745,N_9746,N_9747,N_9748,N_9749,N_9751,N_9752,N_9754,N_9755,N_9759,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9768,N_9770,N_9771,N_9774,N_9777,N_9778,N_9779,N_9780,N_9782,N_9783,N_9785,N_9786,N_9788,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9798,N_9799,N_9800,N_9803,N_9804,N_9806,N_9807,N_9808,N_9809,N_9811,N_9813,N_9814,N_9815,N_9817,N_9818,N_9819,N_9820,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9833,N_9834,N_9836,N_9837,N_9839,N_9840,N_9842,N_9844,N_9847,N_9848,N_9850,N_9853,N_9854,N_9855,N_9857,N_9859,N_9862,N_9863,N_9864,N_9867,N_9869,N_9871,N_9872,N_9874,N_9878,N_9879,N_9880,N_9881,N_9882,N_9884,N_9886,N_9888,N_9889,N_9890,N_9892,N_9895,N_9897,N_9898,N_9899,N_9902,N_9903,N_9906,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9916,N_9918,N_9919,N_9921,N_9922,N_9924,N_9925,N_9926,N_9927,N_9928,N_9930,N_9931,N_9932,N_9934,N_9935,N_9936,N_9938,N_9939,N_9940,N_9941,N_9942,N_9946,N_9947,N_9949,N_9950,N_9951,N_9952,N_9953,N_9956,N_9957,N_9960,N_9961,N_9963,N_9964,N_9967,N_9968,N_9969,N_9971,N_9972,N_9973,N_9977,N_9978,N_9979,N_9983,N_9984,N_9985,N_9986,N_9990,N_9992,N_9993,N_9994,N_9995,N_9998,N_9999;
or U0 (N_0,In_266,In_167);
nor U1 (N_1,In_446,In_525);
or U2 (N_2,In_540,In_919);
and U3 (N_3,In_715,In_500);
nand U4 (N_4,In_469,In_428);
or U5 (N_5,In_275,In_961);
or U6 (N_6,In_641,In_753);
and U7 (N_7,In_203,In_455);
and U8 (N_8,In_567,In_64);
and U9 (N_9,In_402,In_856);
nor U10 (N_10,In_981,In_707);
nor U11 (N_11,In_538,In_30);
nand U12 (N_12,In_68,In_116);
or U13 (N_13,In_725,In_899);
or U14 (N_14,In_957,In_118);
nor U15 (N_15,In_733,In_443);
nor U16 (N_16,In_996,In_143);
and U17 (N_17,In_794,In_530);
nand U18 (N_18,In_59,In_234);
nand U19 (N_19,In_965,In_461);
nand U20 (N_20,In_32,In_375);
nand U21 (N_21,In_233,In_687);
nand U22 (N_22,In_44,In_781);
nand U23 (N_23,In_175,In_762);
nand U24 (N_24,In_183,In_204);
and U25 (N_25,In_142,In_328);
nor U26 (N_26,In_975,In_580);
nor U27 (N_27,In_172,In_63);
and U28 (N_28,In_246,In_703);
or U29 (N_29,In_0,In_739);
nor U30 (N_30,In_813,In_437);
xor U31 (N_31,In_836,In_651);
and U32 (N_32,In_290,In_481);
and U33 (N_33,In_216,In_646);
and U34 (N_34,In_863,In_51);
and U35 (N_35,In_156,In_327);
xnor U36 (N_36,In_70,In_135);
and U37 (N_37,In_879,In_405);
nand U38 (N_38,In_11,In_946);
nor U39 (N_39,In_810,In_48);
and U40 (N_40,In_952,In_858);
or U41 (N_41,In_416,In_657);
and U42 (N_42,In_241,In_303);
nor U43 (N_43,In_129,In_441);
nor U44 (N_44,In_320,In_690);
and U45 (N_45,In_360,In_171);
or U46 (N_46,In_424,In_34);
and U47 (N_47,In_133,In_238);
nor U48 (N_48,In_72,In_341);
or U49 (N_49,In_754,In_471);
nand U50 (N_50,In_199,In_205);
or U51 (N_51,In_683,In_491);
or U52 (N_52,In_230,In_224);
or U53 (N_53,In_12,In_406);
and U54 (N_54,In_571,In_463);
nand U55 (N_55,In_928,In_758);
and U56 (N_56,In_512,In_779);
and U57 (N_57,In_716,In_583);
or U58 (N_58,In_589,In_608);
nand U59 (N_59,In_296,In_252);
nand U60 (N_60,In_990,In_955);
nor U61 (N_61,In_594,In_737);
or U62 (N_62,In_977,In_237);
or U63 (N_63,In_679,In_647);
nand U64 (N_64,In_901,In_968);
or U65 (N_65,In_759,In_126);
nand U66 (N_66,In_165,In_862);
xor U67 (N_67,In_848,In_526);
or U68 (N_68,In_89,In_113);
and U69 (N_69,In_736,In_6);
nand U70 (N_70,In_685,In_676);
or U71 (N_71,In_950,In_780);
nor U72 (N_72,In_342,In_556);
and U73 (N_73,In_192,In_381);
nand U74 (N_74,In_382,In_144);
and U75 (N_75,In_395,In_778);
nand U76 (N_76,In_131,In_728);
nor U77 (N_77,In_174,In_958);
or U78 (N_78,In_91,In_558);
and U79 (N_79,In_939,In_574);
nor U80 (N_80,In_591,In_811);
xnor U81 (N_81,In_371,In_206);
nor U82 (N_82,In_564,In_934);
and U83 (N_83,In_547,In_849);
or U84 (N_84,In_403,In_756);
nor U85 (N_85,In_527,In_450);
xor U86 (N_86,In_136,In_384);
nor U87 (N_87,In_912,In_55);
or U88 (N_88,In_937,In_807);
or U89 (N_89,In_141,In_378);
nand U90 (N_90,In_677,In_642);
or U91 (N_91,In_221,In_742);
and U92 (N_92,In_495,In_826);
nand U93 (N_93,In_573,In_622);
nand U94 (N_94,In_837,In_768);
nor U95 (N_95,In_845,In_684);
nand U96 (N_96,In_488,In_81);
and U97 (N_97,In_2,In_308);
and U98 (N_98,In_732,In_734);
nor U99 (N_99,In_309,In_138);
nor U100 (N_100,In_741,In_701);
nor U101 (N_101,In_812,In_503);
nor U102 (N_102,In_602,In_370);
nor U103 (N_103,In_694,In_897);
nand U104 (N_104,In_572,In_902);
nor U105 (N_105,In_379,In_470);
and U106 (N_106,In_232,In_688);
and U107 (N_107,In_648,In_933);
nor U108 (N_108,In_3,In_343);
nand U109 (N_109,In_692,In_255);
nor U110 (N_110,In_835,In_605);
nand U111 (N_111,In_562,In_14);
nor U112 (N_112,In_289,In_760);
and U113 (N_113,In_58,In_537);
nor U114 (N_114,In_804,In_531);
nand U115 (N_115,In_757,In_13);
nor U116 (N_116,In_367,In_740);
and U117 (N_117,In_417,In_41);
nand U118 (N_118,In_168,In_498);
nor U119 (N_119,In_595,In_501);
or U120 (N_120,In_42,In_351);
or U121 (N_121,In_823,In_253);
nand U122 (N_122,In_465,In_774);
or U123 (N_123,In_288,In_776);
nand U124 (N_124,In_421,In_28);
or U125 (N_125,In_816,In_904);
nor U126 (N_126,In_997,In_551);
and U127 (N_127,In_795,In_453);
and U128 (N_128,In_793,In_448);
or U129 (N_129,In_82,In_159);
nor U130 (N_130,In_999,In_160);
and U131 (N_131,In_185,In_814);
or U132 (N_132,In_248,In_483);
nand U133 (N_133,In_983,In_980);
or U134 (N_134,In_400,In_978);
nor U135 (N_135,In_743,In_154);
or U136 (N_136,In_299,In_818);
nand U137 (N_137,In_960,In_103);
and U138 (N_138,In_350,In_456);
xor U139 (N_139,In_936,In_691);
nor U140 (N_140,In_261,In_827);
and U141 (N_141,In_738,In_47);
or U142 (N_142,In_967,In_607);
and U143 (N_143,In_669,In_429);
or U144 (N_144,In_969,In_932);
and U145 (N_145,In_713,In_336);
nand U146 (N_146,In_60,In_942);
and U147 (N_147,In_925,In_891);
nand U148 (N_148,In_390,In_998);
nor U149 (N_149,In_730,In_26);
or U150 (N_150,In_392,In_831);
nand U151 (N_151,In_473,In_765);
or U152 (N_152,In_560,In_166);
or U153 (N_153,In_553,In_844);
nand U154 (N_154,In_412,In_783);
xor U155 (N_155,In_766,In_930);
nor U156 (N_156,In_374,In_22);
nand U157 (N_157,In_949,In_90);
and U158 (N_158,In_581,In_764);
or U159 (N_159,In_621,In_763);
nand U160 (N_160,In_660,In_52);
and U161 (N_161,In_365,In_18);
or U162 (N_162,In_331,In_888);
or U163 (N_163,In_102,In_236);
or U164 (N_164,In_941,In_935);
nor U165 (N_165,In_427,In_654);
nor U166 (N_166,In_312,In_127);
or U167 (N_167,In_563,In_419);
and U168 (N_168,In_130,In_228);
or U169 (N_169,In_723,In_265);
nor U170 (N_170,In_182,In_330);
nand U171 (N_171,In_627,In_666);
or U172 (N_172,In_566,In_115);
nand U173 (N_173,In_750,In_956);
and U174 (N_174,In_854,In_636);
or U175 (N_175,In_549,In_74);
nor U176 (N_176,In_69,In_77);
nand U177 (N_177,In_578,In_601);
nor U178 (N_178,In_119,In_46);
nand U179 (N_179,In_974,In_62);
nor U180 (N_180,In_954,In_575);
and U181 (N_181,In_515,In_88);
nand U182 (N_182,In_179,In_96);
nand U183 (N_183,In_297,In_434);
and U184 (N_184,In_339,In_287);
nor U185 (N_185,In_366,In_245);
nor U186 (N_186,In_803,In_132);
nand U187 (N_187,In_259,In_482);
and U188 (N_188,In_440,In_842);
and U189 (N_189,In_302,In_7);
and U190 (N_190,In_623,In_786);
nand U191 (N_191,In_445,In_630);
nor U192 (N_192,In_632,In_430);
nor U193 (N_193,In_714,In_383);
or U194 (N_194,In_466,In_273);
nand U195 (N_195,In_755,In_239);
or U196 (N_196,In_634,In_993);
nor U197 (N_197,In_529,In_436);
or U198 (N_198,In_208,In_924);
or U199 (N_199,In_250,In_86);
and U200 (N_200,In_535,In_256);
nand U201 (N_201,In_301,In_678);
nor U202 (N_202,In_663,In_513);
and U203 (N_203,In_358,In_114);
nor U204 (N_204,In_94,In_661);
or U205 (N_205,In_886,In_45);
nand U206 (N_206,In_354,In_702);
or U207 (N_207,In_212,In_561);
or U208 (N_208,In_307,In_598);
nand U209 (N_209,In_536,In_911);
nand U210 (N_210,In_909,In_181);
nor U211 (N_211,In_217,In_699);
nand U212 (N_212,In_866,In_511);
nor U213 (N_213,In_979,In_986);
or U214 (N_214,In_545,In_347);
or U215 (N_215,In_170,In_505);
xor U216 (N_216,In_926,In_889);
or U217 (N_217,In_244,In_388);
or U218 (N_218,In_78,In_251);
nor U219 (N_219,In_134,In_921);
and U220 (N_220,In_884,In_846);
nand U221 (N_221,In_31,In_709);
nor U222 (N_222,In_396,In_294);
and U223 (N_223,In_973,In_518);
nor U224 (N_224,In_479,In_480);
nor U225 (N_225,In_721,In_914);
and U226 (N_226,In_617,In_502);
and U227 (N_227,In_704,In_729);
nor U228 (N_228,In_944,In_872);
nand U229 (N_229,In_752,In_337);
nor U230 (N_230,In_346,In_868);
or U231 (N_231,In_585,In_325);
nand U232 (N_232,In_368,In_910);
nand U233 (N_233,In_613,In_857);
nand U234 (N_234,In_670,In_590);
and U235 (N_235,In_293,In_711);
and U236 (N_236,In_604,In_992);
or U237 (N_237,In_484,In_146);
nor U238 (N_238,In_913,In_705);
and U239 (N_239,In_976,In_398);
or U240 (N_240,In_927,In_528);
nand U241 (N_241,In_782,In_163);
and U242 (N_242,In_861,In_798);
or U243 (N_243,In_649,In_603);
nand U244 (N_244,In_317,In_260);
xor U245 (N_245,In_283,In_698);
nor U246 (N_246,In_270,In_800);
or U247 (N_247,In_139,In_464);
nand U248 (N_248,In_458,In_292);
nand U249 (N_249,In_322,In_363);
nand U250 (N_250,In_544,In_348);
or U251 (N_251,In_614,In_539);
nor U252 (N_252,In_258,In_681);
nand U253 (N_253,In_903,In_124);
or U254 (N_254,In_945,In_148);
and U255 (N_255,In_724,In_71);
or U256 (N_256,In_407,In_971);
or U257 (N_257,In_907,In_867);
nand U258 (N_258,In_696,In_271);
nand U259 (N_259,In_247,In_67);
and U260 (N_260,In_616,In_353);
and U261 (N_261,In_791,In_467);
and U262 (N_262,In_435,In_321);
or U263 (N_263,In_125,In_664);
nor U264 (N_264,In_225,In_584);
and U265 (N_265,In_821,In_279);
nand U266 (N_266,In_414,In_213);
nand U267 (N_267,In_319,In_655);
nand U268 (N_268,In_460,In_109);
nand U269 (N_269,In_376,In_316);
and U270 (N_270,In_372,In_85);
or U271 (N_271,In_659,In_878);
nand U272 (N_272,In_896,In_882);
nor U273 (N_273,In_408,In_462);
and U274 (N_274,In_508,In_95);
nand U275 (N_275,In_789,In_313);
and U276 (N_276,In_291,In_682);
and U277 (N_277,In_227,In_905);
nor U278 (N_278,In_140,In_853);
or U279 (N_279,In_17,In_689);
and U280 (N_280,In_894,In_653);
and U281 (N_281,In_357,In_425);
nor U282 (N_282,In_100,In_625);
nand U283 (N_283,In_223,In_311);
and U284 (N_284,In_117,In_523);
nor U285 (N_285,In_439,In_329);
or U286 (N_286,In_438,In_306);
nand U287 (N_287,In_860,In_272);
and U288 (N_288,In_817,In_300);
and U289 (N_289,In_596,In_497);
or U290 (N_290,In_184,In_507);
nand U291 (N_291,In_727,In_243);
nor U292 (N_292,In_477,In_988);
and U293 (N_293,In_147,In_33);
and U294 (N_294,In_592,In_447);
nor U295 (N_295,In_269,In_305);
and U296 (N_296,In_284,In_37);
nand U297 (N_297,In_478,In_304);
xor U298 (N_298,In_839,In_394);
nand U299 (N_299,In_35,In_50);
or U300 (N_300,In_788,In_611);
nand U301 (N_301,In_644,In_674);
or U302 (N_302,In_514,In_619);
nand U303 (N_303,In_559,In_20);
nand U304 (N_304,In_640,In_808);
nor U305 (N_305,In_310,In_8);
nand U306 (N_306,In_966,In_801);
nor U307 (N_307,In_542,In_87);
nand U308 (N_308,In_264,In_496);
and U309 (N_309,In_624,In_486);
or U310 (N_310,In_274,In_240);
nand U311 (N_311,In_770,In_105);
or U312 (N_312,In_54,In_599);
nor U313 (N_313,In_892,In_187);
nand U314 (N_314,In_324,In_972);
and U315 (N_315,In_151,In_25);
and U316 (N_316,In_610,In_635);
xor U317 (N_317,In_833,In_377);
or U318 (N_318,In_333,In_53);
nand U319 (N_319,In_799,In_873);
nand U320 (N_320,In_790,In_796);
nand U321 (N_321,In_176,In_207);
nand U322 (N_322,In_104,In_819);
nor U323 (N_323,In_340,In_586);
or U324 (N_324,In_620,In_57);
or U325 (N_325,In_66,In_459);
nand U326 (N_326,In_735,In_422);
and U327 (N_327,In_838,In_19);
nor U328 (N_328,In_832,In_169);
nand U329 (N_329,In_364,In_633);
nor U330 (N_330,In_829,In_286);
nand U331 (N_331,In_665,In_541);
xnor U332 (N_332,In_432,In_215);
or U333 (N_333,In_864,In_219);
nor U334 (N_334,In_587,In_579);
and U335 (N_335,In_76,In_220);
or U336 (N_336,In_697,In_9);
nand U337 (N_337,In_629,In_420);
nand U338 (N_338,In_29,In_546);
and U339 (N_339,In_5,In_344);
nand U340 (N_340,In_851,In_451);
or U341 (N_341,In_533,In_982);
or U342 (N_342,In_943,In_906);
nor U343 (N_343,In_161,In_667);
and U344 (N_344,In_652,In_509);
and U345 (N_345,In_680,In_970);
nand U346 (N_346,In_893,In_638);
nor U347 (N_347,In_922,In_843);
xnor U348 (N_348,In_235,In_675);
nor U349 (N_349,In_281,In_908);
or U350 (N_350,In_285,In_771);
or U351 (N_351,In_410,In_257);
and U352 (N_352,In_524,In_92);
and U353 (N_353,In_23,In_373);
and U354 (N_354,In_226,In_457);
nor U355 (N_355,In_280,In_210);
xor U356 (N_356,In_195,In_385);
or U357 (N_357,In_194,In_994);
and U358 (N_358,In_506,In_947);
nand U359 (N_359,In_984,In_431);
or U360 (N_360,In_569,In_211);
or U361 (N_361,In_612,In_577);
nand U362 (N_362,In_49,In_21);
and U363 (N_363,In_214,In_820);
and U364 (N_364,In_494,In_731);
and U365 (N_365,In_850,In_887);
or U366 (N_366,In_401,In_744);
nand U367 (N_367,In_885,In_995);
or U368 (N_368,In_834,In_387);
and U369 (N_369,In_315,In_80);
nand U370 (N_370,In_399,In_209);
xnor U371 (N_371,In_359,In_606);
or U372 (N_372,In_111,In_940);
or U373 (N_373,In_875,In_468);
nor U374 (N_374,In_474,In_487);
nand U375 (N_375,In_915,In_177);
or U376 (N_376,In_609,In_769);
and U377 (N_377,In_189,In_852);
and U378 (N_378,In_485,In_706);
or U379 (N_379,In_686,In_106);
nor U380 (N_380,In_39,In_881);
nor U381 (N_381,In_231,In_668);
xnor U382 (N_382,In_393,In_155);
nand U383 (N_383,In_369,In_61);
nor U384 (N_384,In_36,In_122);
nand U385 (N_385,In_520,In_145);
or U386 (N_386,In_631,In_726);
nor U387 (N_387,In_865,In_552);
nand U388 (N_388,In_582,In_200);
nand U389 (N_389,In_84,In_229);
nor U390 (N_390,In_157,In_792);
nand U391 (N_391,In_824,In_99);
nor U392 (N_392,In_27,In_362);
or U393 (N_393,In_841,In_600);
or U394 (N_394,In_948,In_671);
nor U395 (N_395,In_355,In_871);
or U396 (N_396,In_639,In_923);
nor U397 (N_397,In_991,In_123);
nand U398 (N_398,In_475,In_521);
nor U399 (N_399,In_717,In_415);
and U400 (N_400,In_918,In_626);
nor U401 (N_401,In_107,In_645);
nor U402 (N_402,In_916,In_550);
and U403 (N_403,In_880,In_75);
or U404 (N_404,In_890,In_314);
or U405 (N_405,In_883,In_489);
and U406 (N_406,In_73,In_158);
or U407 (N_407,In_748,In_178);
and U408 (N_408,In_806,In_449);
nand U409 (N_409,In_191,In_65);
and U410 (N_410,In_672,In_874);
or U411 (N_411,In_938,In_38);
nor U412 (N_412,In_504,In_352);
or U413 (N_413,In_193,In_444);
nand U414 (N_414,In_276,In_43);
nand U415 (N_415,In_332,In_548);
nor U416 (N_416,In_121,In_345);
and U417 (N_417,In_476,In_749);
or U418 (N_418,In_137,In_855);
or U419 (N_419,In_534,In_202);
or U420 (N_420,In_775,In_628);
xnor U421 (N_421,In_597,In_719);
nand U422 (N_422,In_454,In_423);
and U423 (N_423,In_802,In_93);
nand U424 (N_424,In_951,In_565);
nor U425 (N_425,In_593,In_576);
nand U426 (N_426,In_334,In_840);
and U427 (N_427,In_805,In_356);
nand U428 (N_428,In_746,In_267);
nand U429 (N_429,In_693,In_254);
or U430 (N_430,In_847,In_149);
and U431 (N_431,In_249,In_809);
nand U432 (N_432,In_712,In_859);
or U433 (N_433,In_110,In_785);
and U434 (N_434,In_877,In_277);
nor U435 (N_435,In_637,In_335);
or U436 (N_436,In_298,In_391);
nand U437 (N_437,In_128,In_15);
nor U438 (N_438,In_747,In_499);
nor U439 (N_439,In_673,In_188);
nand U440 (N_440,In_761,In_97);
or U441 (N_441,In_797,In_718);
or U442 (N_442,In_222,In_318);
and U443 (N_443,In_108,In_898);
and U444 (N_444,In_323,In_876);
and U445 (N_445,In_380,In_197);
or U446 (N_446,In_413,In_869);
or U447 (N_447,In_150,In_101);
and U448 (N_448,In_263,In_557);
nor U449 (N_449,In_777,In_650);
or U450 (N_450,In_787,In_418);
nand U451 (N_451,In_722,In_326);
xnor U452 (N_452,In_282,In_409);
or U453 (N_453,In_218,In_555);
or U454 (N_454,In_570,In_618);
nand U455 (N_455,In_773,In_700);
nand U456 (N_456,In_917,In_190);
nand U457 (N_457,In_426,In_615);
nand U458 (N_458,In_987,In_186);
nand U459 (N_459,In_268,In_338);
nor U460 (N_460,In_643,In_920);
or U461 (N_461,In_83,In_201);
nand U462 (N_462,In_953,In_900);
or U463 (N_463,In_490,In_815);
or U464 (N_464,In_162,In_656);
nor U465 (N_465,In_695,In_895);
and U466 (N_466,In_4,In_822);
or U467 (N_467,In_767,In_112);
and U468 (N_468,In_98,In_510);
nor U469 (N_469,In_472,In_532);
nor U470 (N_470,In_442,In_588);
and U471 (N_471,In_784,In_242);
nand U472 (N_472,In_710,In_16);
or U473 (N_473,In_397,In_452);
or U474 (N_474,In_708,In_152);
or U475 (N_475,In_180,In_543);
nand U476 (N_476,In_10,In_720);
nand U477 (N_477,In_262,In_963);
nor U478 (N_478,In_870,In_568);
or U479 (N_479,In_554,In_493);
and U480 (N_480,In_79,In_56);
and U481 (N_481,In_198,In_745);
or U482 (N_482,In_164,In_989);
or U483 (N_483,In_929,In_1);
nor U484 (N_484,In_522,In_962);
and U485 (N_485,In_517,In_931);
and U486 (N_486,In_662,In_24);
nand U487 (N_487,In_120,In_404);
nand U488 (N_488,In_389,In_173);
and U489 (N_489,In_519,In_964);
or U490 (N_490,In_40,In_825);
or U491 (N_491,In_516,In_196);
nand U492 (N_492,In_278,In_386);
or U493 (N_493,In_959,In_830);
nand U494 (N_494,In_349,In_828);
nand U495 (N_495,In_772,In_411);
and U496 (N_496,In_492,In_433);
nand U497 (N_497,In_153,In_985);
or U498 (N_498,In_361,In_751);
nand U499 (N_499,In_658,In_295);
nand U500 (N_500,In_912,In_194);
or U501 (N_501,In_759,In_780);
nand U502 (N_502,In_266,In_241);
or U503 (N_503,In_232,In_356);
and U504 (N_504,In_463,In_734);
and U505 (N_505,In_315,In_180);
or U506 (N_506,In_582,In_724);
nor U507 (N_507,In_520,In_829);
nor U508 (N_508,In_246,In_55);
xor U509 (N_509,In_813,In_714);
and U510 (N_510,In_258,In_856);
nand U511 (N_511,In_992,In_244);
or U512 (N_512,In_652,In_241);
nor U513 (N_513,In_595,In_860);
and U514 (N_514,In_346,In_260);
nor U515 (N_515,In_810,In_764);
nand U516 (N_516,In_352,In_523);
nor U517 (N_517,In_892,In_241);
nor U518 (N_518,In_476,In_518);
nand U519 (N_519,In_372,In_569);
nor U520 (N_520,In_384,In_884);
nand U521 (N_521,In_517,In_24);
nand U522 (N_522,In_179,In_308);
nand U523 (N_523,In_507,In_414);
nand U524 (N_524,In_135,In_468);
nor U525 (N_525,In_145,In_381);
nor U526 (N_526,In_616,In_311);
and U527 (N_527,In_195,In_952);
nand U528 (N_528,In_17,In_296);
or U529 (N_529,In_936,In_892);
nand U530 (N_530,In_343,In_402);
and U531 (N_531,In_289,In_51);
nand U532 (N_532,In_556,In_294);
and U533 (N_533,In_830,In_989);
and U534 (N_534,In_249,In_993);
and U535 (N_535,In_387,In_613);
and U536 (N_536,In_224,In_34);
nand U537 (N_537,In_566,In_210);
and U538 (N_538,In_107,In_471);
nor U539 (N_539,In_942,In_263);
and U540 (N_540,In_454,In_745);
or U541 (N_541,In_381,In_424);
and U542 (N_542,In_825,In_358);
or U543 (N_543,In_168,In_817);
and U544 (N_544,In_788,In_974);
or U545 (N_545,In_816,In_67);
nor U546 (N_546,In_521,In_656);
nor U547 (N_547,In_435,In_411);
or U548 (N_548,In_791,In_192);
nor U549 (N_549,In_91,In_955);
or U550 (N_550,In_822,In_845);
and U551 (N_551,In_72,In_903);
or U552 (N_552,In_860,In_767);
and U553 (N_553,In_147,In_716);
nand U554 (N_554,In_303,In_970);
and U555 (N_555,In_646,In_817);
or U556 (N_556,In_660,In_568);
and U557 (N_557,In_121,In_365);
or U558 (N_558,In_80,In_931);
nand U559 (N_559,In_777,In_821);
nor U560 (N_560,In_742,In_338);
and U561 (N_561,In_605,In_123);
nand U562 (N_562,In_641,In_529);
and U563 (N_563,In_688,In_295);
or U564 (N_564,In_186,In_485);
or U565 (N_565,In_295,In_522);
or U566 (N_566,In_845,In_759);
or U567 (N_567,In_208,In_824);
and U568 (N_568,In_267,In_239);
nand U569 (N_569,In_8,In_303);
and U570 (N_570,In_735,In_425);
and U571 (N_571,In_258,In_943);
or U572 (N_572,In_317,In_571);
nand U573 (N_573,In_832,In_70);
nand U574 (N_574,In_42,In_2);
or U575 (N_575,In_993,In_501);
and U576 (N_576,In_629,In_727);
nand U577 (N_577,In_838,In_54);
nand U578 (N_578,In_140,In_251);
nand U579 (N_579,In_406,In_618);
nand U580 (N_580,In_970,In_435);
and U581 (N_581,In_781,In_734);
or U582 (N_582,In_928,In_300);
or U583 (N_583,In_337,In_332);
and U584 (N_584,In_673,In_81);
nand U585 (N_585,In_629,In_198);
or U586 (N_586,In_362,In_482);
nor U587 (N_587,In_510,In_172);
nand U588 (N_588,In_582,In_805);
or U589 (N_589,In_537,In_495);
nor U590 (N_590,In_10,In_771);
nor U591 (N_591,In_852,In_962);
nor U592 (N_592,In_479,In_306);
nor U593 (N_593,In_675,In_216);
and U594 (N_594,In_102,In_974);
or U595 (N_595,In_703,In_515);
nand U596 (N_596,In_896,In_235);
nor U597 (N_597,In_689,In_105);
and U598 (N_598,In_200,In_125);
nand U599 (N_599,In_415,In_753);
nand U600 (N_600,In_752,In_387);
nor U601 (N_601,In_624,In_800);
and U602 (N_602,In_484,In_214);
nor U603 (N_603,In_685,In_312);
and U604 (N_604,In_763,In_421);
or U605 (N_605,In_959,In_533);
and U606 (N_606,In_53,In_248);
nand U607 (N_607,In_594,In_784);
nand U608 (N_608,In_397,In_245);
nand U609 (N_609,In_367,In_505);
or U610 (N_610,In_982,In_372);
nor U611 (N_611,In_903,In_974);
nor U612 (N_612,In_693,In_972);
or U613 (N_613,In_286,In_916);
nand U614 (N_614,In_368,In_141);
nand U615 (N_615,In_801,In_821);
nand U616 (N_616,In_319,In_972);
and U617 (N_617,In_979,In_721);
nand U618 (N_618,In_289,In_38);
nand U619 (N_619,In_83,In_378);
nor U620 (N_620,In_882,In_39);
and U621 (N_621,In_729,In_580);
nor U622 (N_622,In_274,In_187);
nand U623 (N_623,In_205,In_686);
nor U624 (N_624,In_671,In_944);
or U625 (N_625,In_218,In_957);
nor U626 (N_626,In_397,In_653);
nor U627 (N_627,In_621,In_307);
and U628 (N_628,In_882,In_843);
or U629 (N_629,In_363,In_395);
or U630 (N_630,In_727,In_535);
or U631 (N_631,In_333,In_866);
and U632 (N_632,In_49,In_379);
and U633 (N_633,In_323,In_429);
nor U634 (N_634,In_892,In_196);
nor U635 (N_635,In_57,In_841);
or U636 (N_636,In_516,In_811);
and U637 (N_637,In_311,In_715);
nor U638 (N_638,In_357,In_812);
nor U639 (N_639,In_549,In_28);
or U640 (N_640,In_450,In_509);
nor U641 (N_641,In_321,In_893);
nor U642 (N_642,In_599,In_387);
or U643 (N_643,In_423,In_205);
or U644 (N_644,In_286,In_593);
nand U645 (N_645,In_19,In_74);
nand U646 (N_646,In_609,In_743);
and U647 (N_647,In_227,In_383);
and U648 (N_648,In_211,In_329);
nand U649 (N_649,In_961,In_331);
nor U650 (N_650,In_983,In_342);
and U651 (N_651,In_53,In_24);
and U652 (N_652,In_669,In_78);
nand U653 (N_653,In_318,In_565);
nand U654 (N_654,In_335,In_317);
and U655 (N_655,In_101,In_690);
nand U656 (N_656,In_944,In_780);
nor U657 (N_657,In_841,In_157);
or U658 (N_658,In_436,In_40);
or U659 (N_659,In_437,In_355);
and U660 (N_660,In_396,In_384);
or U661 (N_661,In_157,In_685);
nor U662 (N_662,In_705,In_163);
and U663 (N_663,In_355,In_711);
or U664 (N_664,In_528,In_646);
or U665 (N_665,In_429,In_437);
and U666 (N_666,In_595,In_858);
nor U667 (N_667,In_804,In_559);
and U668 (N_668,In_472,In_937);
and U669 (N_669,In_442,In_90);
nand U670 (N_670,In_546,In_84);
nand U671 (N_671,In_937,In_449);
or U672 (N_672,In_624,In_466);
and U673 (N_673,In_738,In_812);
nand U674 (N_674,In_73,In_518);
nand U675 (N_675,In_742,In_50);
nand U676 (N_676,In_937,In_304);
or U677 (N_677,In_371,In_45);
and U678 (N_678,In_684,In_765);
nor U679 (N_679,In_997,In_358);
nand U680 (N_680,In_743,In_473);
nor U681 (N_681,In_751,In_556);
nand U682 (N_682,In_219,In_972);
nand U683 (N_683,In_631,In_542);
and U684 (N_684,In_340,In_956);
and U685 (N_685,In_808,In_194);
nand U686 (N_686,In_64,In_864);
or U687 (N_687,In_193,In_126);
nor U688 (N_688,In_188,In_585);
or U689 (N_689,In_264,In_772);
and U690 (N_690,In_174,In_27);
and U691 (N_691,In_598,In_21);
nor U692 (N_692,In_862,In_995);
nand U693 (N_693,In_164,In_880);
and U694 (N_694,In_912,In_181);
and U695 (N_695,In_536,In_241);
and U696 (N_696,In_568,In_156);
and U697 (N_697,In_470,In_505);
nand U698 (N_698,In_870,In_865);
or U699 (N_699,In_471,In_741);
nand U700 (N_700,In_561,In_614);
nand U701 (N_701,In_21,In_393);
nand U702 (N_702,In_469,In_256);
and U703 (N_703,In_563,In_927);
nor U704 (N_704,In_510,In_307);
nand U705 (N_705,In_929,In_192);
or U706 (N_706,In_487,In_984);
nor U707 (N_707,In_695,In_405);
or U708 (N_708,In_663,In_956);
or U709 (N_709,In_898,In_261);
xor U710 (N_710,In_274,In_941);
or U711 (N_711,In_999,In_910);
nand U712 (N_712,In_885,In_834);
and U713 (N_713,In_280,In_375);
or U714 (N_714,In_479,In_663);
nand U715 (N_715,In_457,In_5);
nand U716 (N_716,In_779,In_273);
nand U717 (N_717,In_155,In_90);
and U718 (N_718,In_543,In_996);
nor U719 (N_719,In_364,In_609);
nor U720 (N_720,In_54,In_349);
nor U721 (N_721,In_425,In_171);
and U722 (N_722,In_610,In_910);
or U723 (N_723,In_780,In_96);
or U724 (N_724,In_139,In_393);
nand U725 (N_725,In_862,In_321);
and U726 (N_726,In_161,In_471);
nand U727 (N_727,In_91,In_456);
or U728 (N_728,In_202,In_998);
nor U729 (N_729,In_483,In_134);
and U730 (N_730,In_964,In_925);
and U731 (N_731,In_416,In_474);
or U732 (N_732,In_953,In_248);
nor U733 (N_733,In_991,In_249);
nor U734 (N_734,In_933,In_312);
nor U735 (N_735,In_761,In_17);
and U736 (N_736,In_768,In_415);
nor U737 (N_737,In_461,In_510);
and U738 (N_738,In_334,In_81);
and U739 (N_739,In_160,In_464);
nor U740 (N_740,In_792,In_89);
and U741 (N_741,In_628,In_786);
nand U742 (N_742,In_74,In_270);
nand U743 (N_743,In_924,In_955);
or U744 (N_744,In_968,In_749);
and U745 (N_745,In_34,In_637);
nor U746 (N_746,In_386,In_102);
and U747 (N_747,In_126,In_826);
and U748 (N_748,In_331,In_412);
and U749 (N_749,In_531,In_117);
and U750 (N_750,In_841,In_955);
and U751 (N_751,In_35,In_581);
and U752 (N_752,In_257,In_470);
nor U753 (N_753,In_5,In_587);
nand U754 (N_754,In_394,In_183);
and U755 (N_755,In_265,In_532);
nor U756 (N_756,In_24,In_302);
and U757 (N_757,In_578,In_885);
and U758 (N_758,In_953,In_351);
and U759 (N_759,In_857,In_779);
nand U760 (N_760,In_938,In_341);
nor U761 (N_761,In_897,In_75);
nand U762 (N_762,In_867,In_701);
or U763 (N_763,In_631,In_891);
and U764 (N_764,In_270,In_792);
and U765 (N_765,In_437,In_955);
and U766 (N_766,In_800,In_108);
nand U767 (N_767,In_212,In_245);
nand U768 (N_768,In_240,In_752);
nor U769 (N_769,In_991,In_143);
or U770 (N_770,In_375,In_212);
or U771 (N_771,In_438,In_103);
nor U772 (N_772,In_189,In_588);
nand U773 (N_773,In_795,In_57);
nor U774 (N_774,In_679,In_944);
or U775 (N_775,In_798,In_727);
or U776 (N_776,In_273,In_910);
nor U777 (N_777,In_487,In_334);
nor U778 (N_778,In_263,In_230);
or U779 (N_779,In_492,In_455);
or U780 (N_780,In_941,In_318);
or U781 (N_781,In_689,In_200);
nor U782 (N_782,In_76,In_563);
or U783 (N_783,In_956,In_247);
or U784 (N_784,In_0,In_531);
and U785 (N_785,In_355,In_997);
and U786 (N_786,In_944,In_711);
nor U787 (N_787,In_908,In_78);
and U788 (N_788,In_124,In_714);
nand U789 (N_789,In_2,In_917);
and U790 (N_790,In_466,In_135);
or U791 (N_791,In_409,In_981);
nor U792 (N_792,In_469,In_87);
and U793 (N_793,In_700,In_982);
nor U794 (N_794,In_142,In_806);
xnor U795 (N_795,In_643,In_963);
and U796 (N_796,In_93,In_823);
or U797 (N_797,In_832,In_126);
nand U798 (N_798,In_476,In_633);
and U799 (N_799,In_507,In_178);
nor U800 (N_800,In_612,In_245);
nand U801 (N_801,In_237,In_920);
and U802 (N_802,In_964,In_581);
nor U803 (N_803,In_536,In_378);
or U804 (N_804,In_765,In_525);
nand U805 (N_805,In_116,In_215);
nand U806 (N_806,In_646,In_402);
nor U807 (N_807,In_502,In_931);
nand U808 (N_808,In_29,In_195);
nor U809 (N_809,In_23,In_826);
and U810 (N_810,In_340,In_439);
or U811 (N_811,In_290,In_321);
nor U812 (N_812,In_508,In_956);
and U813 (N_813,In_867,In_451);
nor U814 (N_814,In_786,In_739);
or U815 (N_815,In_321,In_416);
or U816 (N_816,In_592,In_20);
nor U817 (N_817,In_295,In_422);
or U818 (N_818,In_223,In_292);
or U819 (N_819,In_105,In_86);
nand U820 (N_820,In_413,In_222);
or U821 (N_821,In_266,In_327);
nand U822 (N_822,In_773,In_887);
or U823 (N_823,In_833,In_341);
and U824 (N_824,In_0,In_260);
nor U825 (N_825,In_569,In_662);
xnor U826 (N_826,In_869,In_376);
or U827 (N_827,In_997,In_67);
or U828 (N_828,In_692,In_828);
nand U829 (N_829,In_407,In_394);
nand U830 (N_830,In_604,In_141);
nor U831 (N_831,In_411,In_961);
nand U832 (N_832,In_694,In_700);
nor U833 (N_833,In_676,In_226);
nand U834 (N_834,In_657,In_526);
nor U835 (N_835,In_724,In_906);
nand U836 (N_836,In_839,In_524);
or U837 (N_837,In_762,In_772);
or U838 (N_838,In_500,In_357);
or U839 (N_839,In_123,In_400);
nand U840 (N_840,In_3,In_612);
nor U841 (N_841,In_31,In_184);
or U842 (N_842,In_575,In_543);
nor U843 (N_843,In_131,In_606);
and U844 (N_844,In_24,In_359);
nand U845 (N_845,In_218,In_277);
and U846 (N_846,In_205,In_292);
nor U847 (N_847,In_678,In_54);
nor U848 (N_848,In_967,In_253);
nand U849 (N_849,In_415,In_982);
and U850 (N_850,In_914,In_783);
or U851 (N_851,In_332,In_53);
xnor U852 (N_852,In_927,In_727);
and U853 (N_853,In_191,In_246);
or U854 (N_854,In_270,In_357);
and U855 (N_855,In_585,In_762);
nand U856 (N_856,In_530,In_392);
or U857 (N_857,In_594,In_564);
nor U858 (N_858,In_389,In_159);
nor U859 (N_859,In_878,In_351);
and U860 (N_860,In_222,In_898);
nor U861 (N_861,In_729,In_500);
nand U862 (N_862,In_433,In_135);
or U863 (N_863,In_493,In_5);
or U864 (N_864,In_129,In_406);
or U865 (N_865,In_658,In_147);
or U866 (N_866,In_780,In_88);
nor U867 (N_867,In_940,In_172);
and U868 (N_868,In_563,In_277);
and U869 (N_869,In_862,In_481);
or U870 (N_870,In_37,In_858);
nand U871 (N_871,In_13,In_145);
or U872 (N_872,In_836,In_373);
nor U873 (N_873,In_913,In_280);
or U874 (N_874,In_888,In_681);
or U875 (N_875,In_151,In_666);
or U876 (N_876,In_767,In_986);
or U877 (N_877,In_924,In_638);
nor U878 (N_878,In_637,In_23);
and U879 (N_879,In_648,In_423);
and U880 (N_880,In_689,In_67);
nor U881 (N_881,In_986,In_821);
and U882 (N_882,In_519,In_677);
nor U883 (N_883,In_526,In_820);
nand U884 (N_884,In_598,In_658);
or U885 (N_885,In_191,In_879);
nand U886 (N_886,In_417,In_365);
or U887 (N_887,In_338,In_283);
or U888 (N_888,In_25,In_338);
nor U889 (N_889,In_667,In_92);
nor U890 (N_890,In_442,In_145);
and U891 (N_891,In_219,In_952);
nor U892 (N_892,In_458,In_880);
or U893 (N_893,In_792,In_435);
and U894 (N_894,In_667,In_242);
and U895 (N_895,In_931,In_671);
and U896 (N_896,In_249,In_81);
nor U897 (N_897,In_432,In_966);
or U898 (N_898,In_963,In_841);
or U899 (N_899,In_213,In_156);
or U900 (N_900,In_87,In_136);
and U901 (N_901,In_470,In_939);
and U902 (N_902,In_270,In_718);
and U903 (N_903,In_704,In_843);
and U904 (N_904,In_143,In_63);
and U905 (N_905,In_759,In_321);
nand U906 (N_906,In_403,In_265);
nor U907 (N_907,In_837,In_782);
or U908 (N_908,In_895,In_885);
and U909 (N_909,In_820,In_564);
and U910 (N_910,In_974,In_546);
or U911 (N_911,In_526,In_943);
nand U912 (N_912,In_628,In_892);
or U913 (N_913,In_766,In_713);
nand U914 (N_914,In_909,In_9);
or U915 (N_915,In_226,In_533);
nand U916 (N_916,In_237,In_468);
and U917 (N_917,In_565,In_69);
nor U918 (N_918,In_285,In_176);
or U919 (N_919,In_731,In_233);
or U920 (N_920,In_471,In_381);
or U921 (N_921,In_255,In_106);
or U922 (N_922,In_773,In_12);
nand U923 (N_923,In_957,In_952);
and U924 (N_924,In_274,In_455);
nand U925 (N_925,In_640,In_805);
and U926 (N_926,In_531,In_400);
nor U927 (N_927,In_434,In_905);
or U928 (N_928,In_445,In_127);
nand U929 (N_929,In_811,In_789);
nand U930 (N_930,In_555,In_938);
xor U931 (N_931,In_406,In_613);
nor U932 (N_932,In_247,In_755);
and U933 (N_933,In_326,In_905);
nand U934 (N_934,In_777,In_144);
nand U935 (N_935,In_658,In_142);
nor U936 (N_936,In_755,In_84);
and U937 (N_937,In_802,In_264);
and U938 (N_938,In_731,In_80);
nor U939 (N_939,In_905,In_324);
nor U940 (N_940,In_864,In_109);
nor U941 (N_941,In_538,In_122);
or U942 (N_942,In_567,In_297);
and U943 (N_943,In_963,In_857);
nand U944 (N_944,In_121,In_785);
xor U945 (N_945,In_20,In_706);
and U946 (N_946,In_507,In_113);
and U947 (N_947,In_563,In_687);
or U948 (N_948,In_310,In_404);
or U949 (N_949,In_691,In_209);
and U950 (N_950,In_674,In_66);
nor U951 (N_951,In_827,In_929);
nor U952 (N_952,In_824,In_381);
xor U953 (N_953,In_982,In_611);
or U954 (N_954,In_492,In_932);
and U955 (N_955,In_604,In_528);
nor U956 (N_956,In_981,In_421);
or U957 (N_957,In_681,In_81);
nand U958 (N_958,In_885,In_255);
and U959 (N_959,In_421,In_692);
or U960 (N_960,In_583,In_44);
or U961 (N_961,In_47,In_453);
xor U962 (N_962,In_482,In_760);
nand U963 (N_963,In_523,In_607);
nand U964 (N_964,In_995,In_633);
nor U965 (N_965,In_226,In_297);
xnor U966 (N_966,In_2,In_738);
nand U967 (N_967,In_88,In_308);
or U968 (N_968,In_970,In_137);
xor U969 (N_969,In_78,In_789);
and U970 (N_970,In_16,In_749);
and U971 (N_971,In_987,In_754);
or U972 (N_972,In_240,In_783);
nor U973 (N_973,In_665,In_427);
and U974 (N_974,In_376,In_291);
or U975 (N_975,In_697,In_408);
xnor U976 (N_976,In_507,In_177);
and U977 (N_977,In_538,In_425);
nor U978 (N_978,In_829,In_103);
and U979 (N_979,In_399,In_744);
or U980 (N_980,In_963,In_373);
and U981 (N_981,In_673,In_378);
nand U982 (N_982,In_836,In_974);
nor U983 (N_983,In_363,In_150);
nand U984 (N_984,In_811,In_775);
nand U985 (N_985,In_911,In_79);
or U986 (N_986,In_151,In_692);
nand U987 (N_987,In_366,In_643);
nand U988 (N_988,In_125,In_803);
xnor U989 (N_989,In_199,In_368);
or U990 (N_990,In_477,In_780);
nor U991 (N_991,In_67,In_910);
xor U992 (N_992,In_287,In_35);
and U993 (N_993,In_973,In_179);
xor U994 (N_994,In_914,In_708);
xor U995 (N_995,In_415,In_36);
or U996 (N_996,In_126,In_250);
and U997 (N_997,In_617,In_683);
or U998 (N_998,In_971,In_17);
and U999 (N_999,In_975,In_539);
nor U1000 (N_1000,In_23,In_591);
or U1001 (N_1001,In_947,In_816);
and U1002 (N_1002,In_246,In_20);
and U1003 (N_1003,In_105,In_121);
nand U1004 (N_1004,In_666,In_453);
and U1005 (N_1005,In_733,In_538);
or U1006 (N_1006,In_122,In_950);
and U1007 (N_1007,In_607,In_516);
and U1008 (N_1008,In_835,In_756);
or U1009 (N_1009,In_535,In_791);
nand U1010 (N_1010,In_372,In_850);
and U1011 (N_1011,In_38,In_478);
or U1012 (N_1012,In_459,In_288);
xnor U1013 (N_1013,In_428,In_791);
nand U1014 (N_1014,In_888,In_483);
nor U1015 (N_1015,In_731,In_14);
or U1016 (N_1016,In_4,In_3);
or U1017 (N_1017,In_905,In_47);
or U1018 (N_1018,In_765,In_287);
and U1019 (N_1019,In_247,In_42);
or U1020 (N_1020,In_193,In_888);
and U1021 (N_1021,In_723,In_721);
nor U1022 (N_1022,In_336,In_273);
or U1023 (N_1023,In_589,In_58);
xnor U1024 (N_1024,In_548,In_979);
nor U1025 (N_1025,In_367,In_744);
nor U1026 (N_1026,In_965,In_518);
and U1027 (N_1027,In_265,In_481);
or U1028 (N_1028,In_202,In_70);
nand U1029 (N_1029,In_749,In_156);
nor U1030 (N_1030,In_174,In_340);
and U1031 (N_1031,In_910,In_662);
xnor U1032 (N_1032,In_958,In_140);
xor U1033 (N_1033,In_694,In_56);
nand U1034 (N_1034,In_388,In_622);
and U1035 (N_1035,In_808,In_774);
xnor U1036 (N_1036,In_445,In_805);
and U1037 (N_1037,In_444,In_597);
nand U1038 (N_1038,In_405,In_297);
nand U1039 (N_1039,In_31,In_290);
nor U1040 (N_1040,In_274,In_302);
and U1041 (N_1041,In_334,In_310);
and U1042 (N_1042,In_20,In_629);
or U1043 (N_1043,In_389,In_965);
nand U1044 (N_1044,In_377,In_240);
or U1045 (N_1045,In_98,In_921);
nand U1046 (N_1046,In_642,In_577);
and U1047 (N_1047,In_153,In_576);
or U1048 (N_1048,In_726,In_968);
and U1049 (N_1049,In_239,In_899);
and U1050 (N_1050,In_33,In_763);
and U1051 (N_1051,In_436,In_910);
and U1052 (N_1052,In_417,In_420);
and U1053 (N_1053,In_120,In_496);
or U1054 (N_1054,In_574,In_325);
and U1055 (N_1055,In_416,In_494);
or U1056 (N_1056,In_242,In_431);
nand U1057 (N_1057,In_170,In_676);
nand U1058 (N_1058,In_338,In_633);
nor U1059 (N_1059,In_841,In_644);
or U1060 (N_1060,In_841,In_742);
nand U1061 (N_1061,In_920,In_805);
xnor U1062 (N_1062,In_512,In_865);
and U1063 (N_1063,In_169,In_5);
nor U1064 (N_1064,In_4,In_760);
and U1065 (N_1065,In_177,In_142);
and U1066 (N_1066,In_277,In_541);
or U1067 (N_1067,In_447,In_159);
nand U1068 (N_1068,In_549,In_215);
or U1069 (N_1069,In_567,In_244);
nand U1070 (N_1070,In_118,In_399);
nor U1071 (N_1071,In_135,In_790);
and U1072 (N_1072,In_620,In_572);
or U1073 (N_1073,In_957,In_688);
and U1074 (N_1074,In_281,In_117);
or U1075 (N_1075,In_514,In_747);
and U1076 (N_1076,In_468,In_209);
xnor U1077 (N_1077,In_439,In_289);
and U1078 (N_1078,In_826,In_783);
or U1079 (N_1079,In_761,In_207);
nor U1080 (N_1080,In_544,In_345);
and U1081 (N_1081,In_113,In_265);
nand U1082 (N_1082,In_468,In_357);
and U1083 (N_1083,In_652,In_497);
nand U1084 (N_1084,In_136,In_980);
nor U1085 (N_1085,In_467,In_880);
nor U1086 (N_1086,In_990,In_151);
nand U1087 (N_1087,In_379,In_230);
nand U1088 (N_1088,In_745,In_278);
nor U1089 (N_1089,In_369,In_737);
nand U1090 (N_1090,In_261,In_913);
nor U1091 (N_1091,In_649,In_431);
nand U1092 (N_1092,In_733,In_157);
nand U1093 (N_1093,In_27,In_622);
nor U1094 (N_1094,In_478,In_708);
nor U1095 (N_1095,In_215,In_117);
and U1096 (N_1096,In_816,In_346);
xor U1097 (N_1097,In_85,In_360);
nor U1098 (N_1098,In_281,In_343);
nor U1099 (N_1099,In_981,In_802);
and U1100 (N_1100,In_354,In_667);
nor U1101 (N_1101,In_296,In_134);
nand U1102 (N_1102,In_616,In_908);
nor U1103 (N_1103,In_272,In_803);
nand U1104 (N_1104,In_423,In_978);
nand U1105 (N_1105,In_735,In_338);
or U1106 (N_1106,In_165,In_763);
nor U1107 (N_1107,In_0,In_650);
and U1108 (N_1108,In_590,In_20);
and U1109 (N_1109,In_415,In_617);
nor U1110 (N_1110,In_338,In_883);
nand U1111 (N_1111,In_324,In_774);
nor U1112 (N_1112,In_221,In_426);
nor U1113 (N_1113,In_334,In_513);
nor U1114 (N_1114,In_194,In_17);
nor U1115 (N_1115,In_583,In_182);
nor U1116 (N_1116,In_334,In_403);
or U1117 (N_1117,In_770,In_805);
nor U1118 (N_1118,In_580,In_849);
and U1119 (N_1119,In_712,In_382);
and U1120 (N_1120,In_165,In_314);
or U1121 (N_1121,In_203,In_747);
nand U1122 (N_1122,In_167,In_216);
or U1123 (N_1123,In_285,In_777);
nand U1124 (N_1124,In_923,In_938);
nor U1125 (N_1125,In_714,In_250);
nand U1126 (N_1126,In_581,In_592);
nand U1127 (N_1127,In_512,In_325);
nand U1128 (N_1128,In_842,In_159);
nor U1129 (N_1129,In_820,In_160);
nor U1130 (N_1130,In_913,In_0);
nor U1131 (N_1131,In_868,In_598);
and U1132 (N_1132,In_413,In_509);
and U1133 (N_1133,In_46,In_959);
nand U1134 (N_1134,In_782,In_513);
and U1135 (N_1135,In_494,In_866);
nand U1136 (N_1136,In_834,In_205);
nand U1137 (N_1137,In_173,In_355);
nand U1138 (N_1138,In_586,In_459);
nor U1139 (N_1139,In_878,In_355);
or U1140 (N_1140,In_913,In_890);
nor U1141 (N_1141,In_419,In_797);
nor U1142 (N_1142,In_355,In_162);
nand U1143 (N_1143,In_505,In_710);
nor U1144 (N_1144,In_401,In_906);
nand U1145 (N_1145,In_407,In_148);
nor U1146 (N_1146,In_781,In_692);
nor U1147 (N_1147,In_223,In_240);
or U1148 (N_1148,In_943,In_795);
nand U1149 (N_1149,In_132,In_853);
and U1150 (N_1150,In_208,In_934);
nor U1151 (N_1151,In_332,In_481);
nor U1152 (N_1152,In_853,In_600);
nand U1153 (N_1153,In_601,In_102);
or U1154 (N_1154,In_60,In_190);
or U1155 (N_1155,In_453,In_207);
nor U1156 (N_1156,In_792,In_370);
and U1157 (N_1157,In_376,In_565);
nand U1158 (N_1158,In_779,In_399);
or U1159 (N_1159,In_658,In_251);
or U1160 (N_1160,In_266,In_245);
nor U1161 (N_1161,In_184,In_220);
or U1162 (N_1162,In_66,In_553);
nor U1163 (N_1163,In_766,In_413);
and U1164 (N_1164,In_564,In_266);
or U1165 (N_1165,In_330,In_78);
xnor U1166 (N_1166,In_543,In_797);
nand U1167 (N_1167,In_667,In_56);
nor U1168 (N_1168,In_760,In_981);
and U1169 (N_1169,In_496,In_4);
or U1170 (N_1170,In_489,In_607);
or U1171 (N_1171,In_405,In_301);
or U1172 (N_1172,In_725,In_135);
nand U1173 (N_1173,In_407,In_194);
or U1174 (N_1174,In_843,In_72);
or U1175 (N_1175,In_876,In_906);
and U1176 (N_1176,In_322,In_607);
and U1177 (N_1177,In_509,In_647);
and U1178 (N_1178,In_893,In_527);
nor U1179 (N_1179,In_300,In_272);
and U1180 (N_1180,In_441,In_448);
and U1181 (N_1181,In_483,In_225);
nor U1182 (N_1182,In_633,In_616);
or U1183 (N_1183,In_493,In_160);
or U1184 (N_1184,In_185,In_587);
or U1185 (N_1185,In_84,In_651);
nor U1186 (N_1186,In_30,In_475);
and U1187 (N_1187,In_570,In_26);
nor U1188 (N_1188,In_598,In_794);
nor U1189 (N_1189,In_702,In_946);
and U1190 (N_1190,In_975,In_558);
nand U1191 (N_1191,In_485,In_170);
and U1192 (N_1192,In_536,In_740);
nor U1193 (N_1193,In_430,In_108);
nor U1194 (N_1194,In_712,In_750);
nand U1195 (N_1195,In_166,In_3);
nand U1196 (N_1196,In_111,In_375);
or U1197 (N_1197,In_27,In_118);
or U1198 (N_1198,In_496,In_864);
nand U1199 (N_1199,In_537,In_95);
and U1200 (N_1200,In_548,In_725);
nor U1201 (N_1201,In_998,In_562);
nor U1202 (N_1202,In_869,In_499);
and U1203 (N_1203,In_205,In_273);
or U1204 (N_1204,In_559,In_994);
or U1205 (N_1205,In_909,In_961);
or U1206 (N_1206,In_282,In_336);
or U1207 (N_1207,In_257,In_589);
and U1208 (N_1208,In_43,In_650);
and U1209 (N_1209,In_30,In_724);
or U1210 (N_1210,In_967,In_152);
or U1211 (N_1211,In_754,In_677);
nor U1212 (N_1212,In_697,In_632);
nand U1213 (N_1213,In_559,In_8);
and U1214 (N_1214,In_989,In_104);
or U1215 (N_1215,In_515,In_805);
nand U1216 (N_1216,In_764,In_249);
nor U1217 (N_1217,In_839,In_611);
nor U1218 (N_1218,In_229,In_963);
nand U1219 (N_1219,In_528,In_231);
and U1220 (N_1220,In_597,In_996);
or U1221 (N_1221,In_451,In_594);
and U1222 (N_1222,In_915,In_990);
nor U1223 (N_1223,In_42,In_774);
and U1224 (N_1224,In_292,In_198);
and U1225 (N_1225,In_521,In_279);
or U1226 (N_1226,In_95,In_397);
and U1227 (N_1227,In_54,In_761);
nor U1228 (N_1228,In_596,In_685);
and U1229 (N_1229,In_242,In_903);
and U1230 (N_1230,In_807,In_716);
and U1231 (N_1231,In_193,In_337);
nand U1232 (N_1232,In_675,In_748);
or U1233 (N_1233,In_780,In_699);
nand U1234 (N_1234,In_85,In_111);
and U1235 (N_1235,In_81,In_696);
nor U1236 (N_1236,In_848,In_742);
nand U1237 (N_1237,In_63,In_829);
nor U1238 (N_1238,In_62,In_380);
and U1239 (N_1239,In_728,In_933);
and U1240 (N_1240,In_776,In_55);
and U1241 (N_1241,In_113,In_549);
or U1242 (N_1242,In_248,In_360);
nor U1243 (N_1243,In_63,In_476);
nor U1244 (N_1244,In_477,In_485);
and U1245 (N_1245,In_302,In_595);
or U1246 (N_1246,In_261,In_576);
or U1247 (N_1247,In_427,In_60);
nand U1248 (N_1248,In_591,In_553);
nand U1249 (N_1249,In_84,In_334);
nand U1250 (N_1250,In_914,In_460);
and U1251 (N_1251,In_626,In_439);
nand U1252 (N_1252,In_358,In_247);
nor U1253 (N_1253,In_46,In_161);
and U1254 (N_1254,In_621,In_650);
and U1255 (N_1255,In_758,In_417);
nor U1256 (N_1256,In_301,In_294);
nand U1257 (N_1257,In_838,In_86);
or U1258 (N_1258,In_867,In_956);
nor U1259 (N_1259,In_876,In_648);
or U1260 (N_1260,In_600,In_413);
nand U1261 (N_1261,In_322,In_112);
nand U1262 (N_1262,In_27,In_138);
or U1263 (N_1263,In_483,In_957);
or U1264 (N_1264,In_961,In_50);
or U1265 (N_1265,In_476,In_472);
nor U1266 (N_1266,In_535,In_5);
nor U1267 (N_1267,In_915,In_674);
nand U1268 (N_1268,In_762,In_492);
or U1269 (N_1269,In_281,In_888);
and U1270 (N_1270,In_920,In_360);
nor U1271 (N_1271,In_533,In_69);
or U1272 (N_1272,In_536,In_686);
and U1273 (N_1273,In_80,In_846);
nor U1274 (N_1274,In_321,In_438);
or U1275 (N_1275,In_357,In_874);
nor U1276 (N_1276,In_666,In_714);
nand U1277 (N_1277,In_978,In_770);
or U1278 (N_1278,In_171,In_386);
nand U1279 (N_1279,In_944,In_401);
nand U1280 (N_1280,In_533,In_54);
and U1281 (N_1281,In_537,In_801);
or U1282 (N_1282,In_364,In_411);
xor U1283 (N_1283,In_947,In_135);
nand U1284 (N_1284,In_842,In_690);
nor U1285 (N_1285,In_559,In_678);
nor U1286 (N_1286,In_252,In_796);
and U1287 (N_1287,In_484,In_323);
nor U1288 (N_1288,In_601,In_157);
nor U1289 (N_1289,In_34,In_126);
nor U1290 (N_1290,In_749,In_570);
and U1291 (N_1291,In_826,In_730);
nor U1292 (N_1292,In_806,In_472);
nand U1293 (N_1293,In_857,In_474);
nor U1294 (N_1294,In_968,In_623);
and U1295 (N_1295,In_775,In_306);
or U1296 (N_1296,In_581,In_633);
nand U1297 (N_1297,In_336,In_874);
nor U1298 (N_1298,In_75,In_566);
and U1299 (N_1299,In_290,In_956);
and U1300 (N_1300,In_774,In_197);
or U1301 (N_1301,In_595,In_428);
nor U1302 (N_1302,In_255,In_520);
nor U1303 (N_1303,In_223,In_941);
and U1304 (N_1304,In_848,In_418);
and U1305 (N_1305,In_826,In_403);
and U1306 (N_1306,In_815,In_586);
nor U1307 (N_1307,In_759,In_312);
nor U1308 (N_1308,In_238,In_246);
nor U1309 (N_1309,In_959,In_491);
nand U1310 (N_1310,In_417,In_430);
nor U1311 (N_1311,In_161,In_652);
nor U1312 (N_1312,In_209,In_25);
nand U1313 (N_1313,In_804,In_197);
and U1314 (N_1314,In_781,In_21);
and U1315 (N_1315,In_202,In_225);
xnor U1316 (N_1316,In_727,In_769);
nand U1317 (N_1317,In_749,In_245);
nor U1318 (N_1318,In_724,In_979);
nand U1319 (N_1319,In_407,In_451);
or U1320 (N_1320,In_968,In_846);
nor U1321 (N_1321,In_176,In_283);
nor U1322 (N_1322,In_55,In_894);
nand U1323 (N_1323,In_691,In_801);
and U1324 (N_1324,In_804,In_823);
or U1325 (N_1325,In_708,In_712);
nand U1326 (N_1326,In_694,In_954);
or U1327 (N_1327,In_368,In_110);
nand U1328 (N_1328,In_656,In_849);
or U1329 (N_1329,In_891,In_857);
nand U1330 (N_1330,In_667,In_723);
nor U1331 (N_1331,In_715,In_678);
or U1332 (N_1332,In_749,In_368);
and U1333 (N_1333,In_750,In_29);
nand U1334 (N_1334,In_251,In_297);
nor U1335 (N_1335,In_289,In_21);
or U1336 (N_1336,In_446,In_307);
nor U1337 (N_1337,In_802,In_154);
nor U1338 (N_1338,In_784,In_482);
nand U1339 (N_1339,In_290,In_944);
and U1340 (N_1340,In_656,In_187);
or U1341 (N_1341,In_685,In_887);
or U1342 (N_1342,In_385,In_519);
or U1343 (N_1343,In_2,In_504);
or U1344 (N_1344,In_167,In_483);
nor U1345 (N_1345,In_37,In_115);
nand U1346 (N_1346,In_300,In_259);
nand U1347 (N_1347,In_277,In_726);
and U1348 (N_1348,In_932,In_772);
and U1349 (N_1349,In_573,In_123);
and U1350 (N_1350,In_907,In_178);
and U1351 (N_1351,In_918,In_527);
and U1352 (N_1352,In_899,In_990);
or U1353 (N_1353,In_26,In_467);
and U1354 (N_1354,In_923,In_836);
nor U1355 (N_1355,In_210,In_48);
or U1356 (N_1356,In_95,In_820);
or U1357 (N_1357,In_52,In_502);
and U1358 (N_1358,In_801,In_328);
nor U1359 (N_1359,In_481,In_498);
or U1360 (N_1360,In_716,In_829);
nor U1361 (N_1361,In_916,In_165);
nand U1362 (N_1362,In_508,In_612);
and U1363 (N_1363,In_338,In_661);
nand U1364 (N_1364,In_681,In_874);
nand U1365 (N_1365,In_337,In_284);
nor U1366 (N_1366,In_35,In_576);
nor U1367 (N_1367,In_617,In_920);
or U1368 (N_1368,In_980,In_270);
xor U1369 (N_1369,In_869,In_63);
nor U1370 (N_1370,In_707,In_775);
nand U1371 (N_1371,In_682,In_136);
nand U1372 (N_1372,In_778,In_74);
and U1373 (N_1373,In_47,In_345);
nor U1374 (N_1374,In_579,In_760);
nand U1375 (N_1375,In_907,In_373);
or U1376 (N_1376,In_781,In_680);
or U1377 (N_1377,In_294,In_629);
or U1378 (N_1378,In_150,In_759);
or U1379 (N_1379,In_360,In_108);
and U1380 (N_1380,In_10,In_545);
nor U1381 (N_1381,In_642,In_52);
nor U1382 (N_1382,In_920,In_506);
or U1383 (N_1383,In_334,In_198);
nand U1384 (N_1384,In_277,In_443);
and U1385 (N_1385,In_435,In_423);
nand U1386 (N_1386,In_759,In_325);
nor U1387 (N_1387,In_318,In_958);
nand U1388 (N_1388,In_316,In_535);
and U1389 (N_1389,In_933,In_433);
nor U1390 (N_1390,In_813,In_645);
and U1391 (N_1391,In_53,In_396);
and U1392 (N_1392,In_125,In_975);
and U1393 (N_1393,In_494,In_317);
nor U1394 (N_1394,In_703,In_983);
or U1395 (N_1395,In_281,In_15);
nand U1396 (N_1396,In_825,In_174);
nand U1397 (N_1397,In_981,In_235);
nor U1398 (N_1398,In_420,In_413);
and U1399 (N_1399,In_66,In_383);
nand U1400 (N_1400,In_812,In_95);
and U1401 (N_1401,In_697,In_472);
nand U1402 (N_1402,In_457,In_876);
nand U1403 (N_1403,In_776,In_298);
nand U1404 (N_1404,In_663,In_731);
nand U1405 (N_1405,In_169,In_254);
and U1406 (N_1406,In_857,In_588);
and U1407 (N_1407,In_573,In_527);
and U1408 (N_1408,In_81,In_711);
and U1409 (N_1409,In_743,In_449);
and U1410 (N_1410,In_50,In_960);
and U1411 (N_1411,In_717,In_898);
or U1412 (N_1412,In_668,In_359);
or U1413 (N_1413,In_640,In_517);
and U1414 (N_1414,In_905,In_583);
nand U1415 (N_1415,In_466,In_61);
nor U1416 (N_1416,In_716,In_338);
and U1417 (N_1417,In_546,In_321);
or U1418 (N_1418,In_911,In_26);
xor U1419 (N_1419,In_750,In_141);
nand U1420 (N_1420,In_362,In_987);
or U1421 (N_1421,In_162,In_159);
nor U1422 (N_1422,In_107,In_426);
and U1423 (N_1423,In_94,In_171);
nand U1424 (N_1424,In_832,In_864);
nand U1425 (N_1425,In_85,In_108);
nor U1426 (N_1426,In_762,In_349);
and U1427 (N_1427,In_206,In_461);
and U1428 (N_1428,In_897,In_54);
xnor U1429 (N_1429,In_890,In_184);
or U1430 (N_1430,In_101,In_469);
and U1431 (N_1431,In_583,In_422);
or U1432 (N_1432,In_442,In_277);
nor U1433 (N_1433,In_357,In_20);
nor U1434 (N_1434,In_855,In_378);
or U1435 (N_1435,In_773,In_537);
and U1436 (N_1436,In_470,In_858);
nand U1437 (N_1437,In_580,In_677);
and U1438 (N_1438,In_325,In_145);
and U1439 (N_1439,In_545,In_788);
or U1440 (N_1440,In_526,In_19);
nor U1441 (N_1441,In_135,In_457);
or U1442 (N_1442,In_939,In_131);
nor U1443 (N_1443,In_429,In_591);
or U1444 (N_1444,In_10,In_736);
nand U1445 (N_1445,In_903,In_788);
or U1446 (N_1446,In_505,In_180);
nand U1447 (N_1447,In_822,In_132);
or U1448 (N_1448,In_860,In_711);
and U1449 (N_1449,In_344,In_40);
xnor U1450 (N_1450,In_837,In_17);
or U1451 (N_1451,In_964,In_10);
nor U1452 (N_1452,In_624,In_910);
and U1453 (N_1453,In_446,In_47);
and U1454 (N_1454,In_146,In_891);
or U1455 (N_1455,In_206,In_551);
nor U1456 (N_1456,In_245,In_872);
or U1457 (N_1457,In_23,In_998);
and U1458 (N_1458,In_623,In_708);
and U1459 (N_1459,In_185,In_775);
and U1460 (N_1460,In_236,In_26);
nor U1461 (N_1461,In_831,In_197);
or U1462 (N_1462,In_719,In_114);
and U1463 (N_1463,In_239,In_990);
nand U1464 (N_1464,In_618,In_688);
nand U1465 (N_1465,In_430,In_73);
xnor U1466 (N_1466,In_582,In_295);
and U1467 (N_1467,In_772,In_543);
or U1468 (N_1468,In_176,In_406);
xor U1469 (N_1469,In_910,In_286);
or U1470 (N_1470,In_790,In_585);
and U1471 (N_1471,In_288,In_760);
and U1472 (N_1472,In_463,In_338);
nand U1473 (N_1473,In_761,In_620);
nor U1474 (N_1474,In_302,In_368);
nor U1475 (N_1475,In_27,In_318);
and U1476 (N_1476,In_975,In_178);
and U1477 (N_1477,In_166,In_129);
nor U1478 (N_1478,In_83,In_619);
nand U1479 (N_1479,In_993,In_894);
and U1480 (N_1480,In_978,In_82);
nand U1481 (N_1481,In_187,In_739);
or U1482 (N_1482,In_728,In_868);
nor U1483 (N_1483,In_271,In_285);
nand U1484 (N_1484,In_394,In_584);
or U1485 (N_1485,In_27,In_767);
or U1486 (N_1486,In_133,In_910);
nand U1487 (N_1487,In_702,In_696);
nor U1488 (N_1488,In_438,In_423);
nand U1489 (N_1489,In_16,In_680);
nor U1490 (N_1490,In_63,In_929);
nor U1491 (N_1491,In_105,In_415);
or U1492 (N_1492,In_740,In_178);
nor U1493 (N_1493,In_185,In_849);
nor U1494 (N_1494,In_948,In_175);
and U1495 (N_1495,In_742,In_405);
and U1496 (N_1496,In_680,In_368);
nor U1497 (N_1497,In_630,In_290);
and U1498 (N_1498,In_555,In_345);
nor U1499 (N_1499,In_61,In_672);
nor U1500 (N_1500,In_166,In_965);
or U1501 (N_1501,In_984,In_323);
or U1502 (N_1502,In_555,In_647);
and U1503 (N_1503,In_799,In_366);
nor U1504 (N_1504,In_618,In_881);
nand U1505 (N_1505,In_51,In_404);
and U1506 (N_1506,In_415,In_637);
or U1507 (N_1507,In_246,In_781);
and U1508 (N_1508,In_930,In_422);
and U1509 (N_1509,In_699,In_611);
and U1510 (N_1510,In_679,In_142);
nor U1511 (N_1511,In_203,In_562);
nor U1512 (N_1512,In_801,In_297);
or U1513 (N_1513,In_743,In_61);
nand U1514 (N_1514,In_248,In_739);
and U1515 (N_1515,In_547,In_376);
xnor U1516 (N_1516,In_83,In_992);
and U1517 (N_1517,In_510,In_938);
or U1518 (N_1518,In_604,In_755);
and U1519 (N_1519,In_901,In_942);
nor U1520 (N_1520,In_846,In_370);
and U1521 (N_1521,In_902,In_530);
nor U1522 (N_1522,In_673,In_421);
xor U1523 (N_1523,In_679,In_1);
nand U1524 (N_1524,In_62,In_723);
or U1525 (N_1525,In_206,In_833);
or U1526 (N_1526,In_855,In_140);
and U1527 (N_1527,In_856,In_631);
or U1528 (N_1528,In_604,In_981);
xnor U1529 (N_1529,In_229,In_350);
or U1530 (N_1530,In_558,In_503);
nand U1531 (N_1531,In_73,In_521);
or U1532 (N_1532,In_384,In_996);
or U1533 (N_1533,In_337,In_849);
nor U1534 (N_1534,In_79,In_108);
and U1535 (N_1535,In_543,In_707);
nand U1536 (N_1536,In_108,In_178);
and U1537 (N_1537,In_615,In_381);
or U1538 (N_1538,In_869,In_693);
and U1539 (N_1539,In_928,In_201);
or U1540 (N_1540,In_220,In_557);
or U1541 (N_1541,In_189,In_517);
and U1542 (N_1542,In_604,In_252);
or U1543 (N_1543,In_973,In_661);
and U1544 (N_1544,In_999,In_360);
nand U1545 (N_1545,In_888,In_807);
nor U1546 (N_1546,In_64,In_682);
and U1547 (N_1547,In_972,In_495);
and U1548 (N_1548,In_957,In_11);
nor U1549 (N_1549,In_455,In_572);
nand U1550 (N_1550,In_638,In_85);
or U1551 (N_1551,In_403,In_16);
and U1552 (N_1552,In_547,In_453);
and U1553 (N_1553,In_327,In_373);
nand U1554 (N_1554,In_296,In_594);
and U1555 (N_1555,In_283,In_686);
nand U1556 (N_1556,In_948,In_936);
or U1557 (N_1557,In_904,In_868);
nand U1558 (N_1558,In_785,In_476);
nor U1559 (N_1559,In_829,In_89);
and U1560 (N_1560,In_463,In_731);
or U1561 (N_1561,In_547,In_84);
or U1562 (N_1562,In_434,In_956);
nor U1563 (N_1563,In_392,In_114);
or U1564 (N_1564,In_465,In_552);
nand U1565 (N_1565,In_815,In_719);
nor U1566 (N_1566,In_772,In_841);
nor U1567 (N_1567,In_43,In_11);
or U1568 (N_1568,In_282,In_728);
or U1569 (N_1569,In_323,In_465);
and U1570 (N_1570,In_36,In_480);
and U1571 (N_1571,In_686,In_633);
or U1572 (N_1572,In_77,In_868);
or U1573 (N_1573,In_303,In_283);
nor U1574 (N_1574,In_922,In_283);
and U1575 (N_1575,In_564,In_915);
nor U1576 (N_1576,In_395,In_801);
nand U1577 (N_1577,In_691,In_958);
nor U1578 (N_1578,In_880,In_345);
nor U1579 (N_1579,In_738,In_253);
nand U1580 (N_1580,In_402,In_955);
nor U1581 (N_1581,In_722,In_350);
nand U1582 (N_1582,In_107,In_814);
or U1583 (N_1583,In_93,In_997);
and U1584 (N_1584,In_673,In_269);
nand U1585 (N_1585,In_179,In_26);
nor U1586 (N_1586,In_356,In_52);
xnor U1587 (N_1587,In_801,In_996);
and U1588 (N_1588,In_399,In_935);
nor U1589 (N_1589,In_888,In_173);
and U1590 (N_1590,In_629,In_861);
nor U1591 (N_1591,In_392,In_304);
and U1592 (N_1592,In_118,In_780);
and U1593 (N_1593,In_709,In_871);
xnor U1594 (N_1594,In_324,In_21);
and U1595 (N_1595,In_486,In_292);
and U1596 (N_1596,In_565,In_726);
nor U1597 (N_1597,In_289,In_344);
nor U1598 (N_1598,In_775,In_262);
and U1599 (N_1599,In_706,In_905);
and U1600 (N_1600,In_305,In_700);
or U1601 (N_1601,In_371,In_265);
or U1602 (N_1602,In_404,In_694);
nand U1603 (N_1603,In_652,In_653);
nor U1604 (N_1604,In_815,In_883);
nor U1605 (N_1605,In_63,In_955);
and U1606 (N_1606,In_747,In_998);
xnor U1607 (N_1607,In_882,In_381);
and U1608 (N_1608,In_449,In_721);
or U1609 (N_1609,In_314,In_746);
and U1610 (N_1610,In_133,In_586);
and U1611 (N_1611,In_619,In_67);
nor U1612 (N_1612,In_447,In_680);
nand U1613 (N_1613,In_247,In_397);
nor U1614 (N_1614,In_484,In_912);
and U1615 (N_1615,In_950,In_322);
nor U1616 (N_1616,In_388,In_640);
and U1617 (N_1617,In_499,In_12);
or U1618 (N_1618,In_468,In_321);
and U1619 (N_1619,In_848,In_468);
nand U1620 (N_1620,In_194,In_465);
or U1621 (N_1621,In_755,In_147);
and U1622 (N_1622,In_638,In_391);
and U1623 (N_1623,In_629,In_126);
nor U1624 (N_1624,In_389,In_850);
and U1625 (N_1625,In_244,In_34);
and U1626 (N_1626,In_401,In_597);
and U1627 (N_1627,In_727,In_638);
nor U1628 (N_1628,In_427,In_84);
and U1629 (N_1629,In_642,In_879);
nand U1630 (N_1630,In_717,In_854);
and U1631 (N_1631,In_407,In_260);
nor U1632 (N_1632,In_384,In_180);
and U1633 (N_1633,In_256,In_563);
nor U1634 (N_1634,In_208,In_476);
nor U1635 (N_1635,In_375,In_853);
and U1636 (N_1636,In_430,In_814);
or U1637 (N_1637,In_554,In_681);
nor U1638 (N_1638,In_746,In_332);
nand U1639 (N_1639,In_492,In_630);
nand U1640 (N_1640,In_338,In_422);
nor U1641 (N_1641,In_71,In_281);
nand U1642 (N_1642,In_228,In_71);
or U1643 (N_1643,In_998,In_599);
xnor U1644 (N_1644,In_36,In_190);
nand U1645 (N_1645,In_25,In_110);
and U1646 (N_1646,In_153,In_354);
or U1647 (N_1647,In_115,In_405);
xnor U1648 (N_1648,In_887,In_176);
and U1649 (N_1649,In_942,In_151);
and U1650 (N_1650,In_452,In_80);
nor U1651 (N_1651,In_832,In_232);
and U1652 (N_1652,In_524,In_569);
nor U1653 (N_1653,In_203,In_8);
nand U1654 (N_1654,In_216,In_70);
nand U1655 (N_1655,In_834,In_764);
or U1656 (N_1656,In_521,In_837);
nor U1657 (N_1657,In_526,In_125);
and U1658 (N_1658,In_903,In_504);
or U1659 (N_1659,In_784,In_478);
nor U1660 (N_1660,In_28,In_890);
nor U1661 (N_1661,In_969,In_253);
nor U1662 (N_1662,In_485,In_309);
or U1663 (N_1663,In_311,In_767);
nand U1664 (N_1664,In_35,In_375);
nor U1665 (N_1665,In_137,In_57);
or U1666 (N_1666,In_123,In_919);
nor U1667 (N_1667,In_483,In_157);
nand U1668 (N_1668,In_446,In_318);
or U1669 (N_1669,In_488,In_410);
nor U1670 (N_1670,In_867,In_102);
nor U1671 (N_1671,In_320,In_695);
and U1672 (N_1672,In_117,In_838);
nor U1673 (N_1673,In_420,In_756);
nand U1674 (N_1674,In_411,In_529);
nor U1675 (N_1675,In_74,In_602);
and U1676 (N_1676,In_127,In_520);
or U1677 (N_1677,In_292,In_233);
and U1678 (N_1678,In_800,In_192);
and U1679 (N_1679,In_456,In_135);
nor U1680 (N_1680,In_31,In_908);
and U1681 (N_1681,In_287,In_526);
and U1682 (N_1682,In_985,In_129);
and U1683 (N_1683,In_129,In_226);
and U1684 (N_1684,In_916,In_527);
nor U1685 (N_1685,In_918,In_806);
nor U1686 (N_1686,In_948,In_191);
nor U1687 (N_1687,In_181,In_174);
nand U1688 (N_1688,In_484,In_833);
or U1689 (N_1689,In_594,In_189);
or U1690 (N_1690,In_431,In_371);
or U1691 (N_1691,In_490,In_394);
nor U1692 (N_1692,In_620,In_531);
nand U1693 (N_1693,In_619,In_666);
and U1694 (N_1694,In_891,In_848);
nor U1695 (N_1695,In_874,In_523);
nor U1696 (N_1696,In_484,In_989);
nand U1697 (N_1697,In_5,In_198);
or U1698 (N_1698,In_404,In_748);
nor U1699 (N_1699,In_861,In_747);
and U1700 (N_1700,In_404,In_132);
nand U1701 (N_1701,In_849,In_77);
and U1702 (N_1702,In_41,In_104);
nand U1703 (N_1703,In_676,In_192);
nor U1704 (N_1704,In_136,In_914);
nor U1705 (N_1705,In_337,In_860);
nand U1706 (N_1706,In_380,In_18);
nand U1707 (N_1707,In_447,In_516);
or U1708 (N_1708,In_774,In_921);
and U1709 (N_1709,In_401,In_764);
or U1710 (N_1710,In_968,In_228);
nand U1711 (N_1711,In_399,In_354);
xor U1712 (N_1712,In_814,In_569);
xnor U1713 (N_1713,In_114,In_331);
and U1714 (N_1714,In_857,In_68);
or U1715 (N_1715,In_154,In_966);
nand U1716 (N_1716,In_618,In_229);
nor U1717 (N_1717,In_547,In_788);
or U1718 (N_1718,In_184,In_266);
xor U1719 (N_1719,In_320,In_58);
and U1720 (N_1720,In_962,In_513);
and U1721 (N_1721,In_879,In_115);
nor U1722 (N_1722,In_888,In_870);
nor U1723 (N_1723,In_741,In_859);
nor U1724 (N_1724,In_886,In_95);
or U1725 (N_1725,In_655,In_283);
nor U1726 (N_1726,In_146,In_665);
nor U1727 (N_1727,In_965,In_130);
or U1728 (N_1728,In_401,In_591);
and U1729 (N_1729,In_259,In_274);
nor U1730 (N_1730,In_641,In_971);
and U1731 (N_1731,In_514,In_815);
or U1732 (N_1732,In_174,In_886);
nor U1733 (N_1733,In_558,In_591);
nand U1734 (N_1734,In_355,In_420);
and U1735 (N_1735,In_524,In_407);
and U1736 (N_1736,In_929,In_75);
and U1737 (N_1737,In_695,In_995);
nand U1738 (N_1738,In_625,In_297);
nand U1739 (N_1739,In_204,In_671);
or U1740 (N_1740,In_743,In_630);
nand U1741 (N_1741,In_759,In_756);
and U1742 (N_1742,In_696,In_155);
and U1743 (N_1743,In_990,In_783);
nor U1744 (N_1744,In_824,In_403);
nor U1745 (N_1745,In_918,In_444);
nor U1746 (N_1746,In_781,In_173);
nor U1747 (N_1747,In_513,In_698);
and U1748 (N_1748,In_293,In_722);
nor U1749 (N_1749,In_299,In_426);
nor U1750 (N_1750,In_458,In_582);
xnor U1751 (N_1751,In_227,In_222);
nand U1752 (N_1752,In_938,In_89);
xnor U1753 (N_1753,In_391,In_791);
nand U1754 (N_1754,In_333,In_630);
nor U1755 (N_1755,In_933,In_601);
nor U1756 (N_1756,In_819,In_396);
or U1757 (N_1757,In_369,In_515);
or U1758 (N_1758,In_189,In_531);
nor U1759 (N_1759,In_419,In_47);
nand U1760 (N_1760,In_464,In_20);
and U1761 (N_1761,In_925,In_978);
nor U1762 (N_1762,In_936,In_946);
nand U1763 (N_1763,In_31,In_447);
or U1764 (N_1764,In_637,In_405);
and U1765 (N_1765,In_109,In_601);
nand U1766 (N_1766,In_759,In_226);
nor U1767 (N_1767,In_669,In_218);
nor U1768 (N_1768,In_909,In_452);
nand U1769 (N_1769,In_170,In_796);
nor U1770 (N_1770,In_674,In_914);
nor U1771 (N_1771,In_70,In_666);
and U1772 (N_1772,In_95,In_903);
and U1773 (N_1773,In_158,In_567);
and U1774 (N_1774,In_231,In_120);
or U1775 (N_1775,In_487,In_813);
nor U1776 (N_1776,In_617,In_726);
nor U1777 (N_1777,In_342,In_588);
and U1778 (N_1778,In_168,In_51);
and U1779 (N_1779,In_74,In_673);
or U1780 (N_1780,In_428,In_739);
and U1781 (N_1781,In_623,In_489);
nand U1782 (N_1782,In_948,In_411);
or U1783 (N_1783,In_635,In_771);
or U1784 (N_1784,In_853,In_539);
nand U1785 (N_1785,In_321,In_800);
nor U1786 (N_1786,In_908,In_559);
and U1787 (N_1787,In_258,In_465);
and U1788 (N_1788,In_781,In_502);
nand U1789 (N_1789,In_644,In_918);
nand U1790 (N_1790,In_150,In_866);
nor U1791 (N_1791,In_58,In_540);
or U1792 (N_1792,In_849,In_482);
nand U1793 (N_1793,In_158,In_3);
nand U1794 (N_1794,In_108,In_318);
nor U1795 (N_1795,In_894,In_308);
nor U1796 (N_1796,In_11,In_542);
nor U1797 (N_1797,In_209,In_893);
nor U1798 (N_1798,In_796,In_852);
or U1799 (N_1799,In_148,In_402);
or U1800 (N_1800,In_378,In_875);
and U1801 (N_1801,In_182,In_729);
nor U1802 (N_1802,In_230,In_619);
or U1803 (N_1803,In_280,In_116);
nor U1804 (N_1804,In_591,In_285);
nand U1805 (N_1805,In_422,In_89);
nand U1806 (N_1806,In_272,In_155);
nor U1807 (N_1807,In_706,In_3);
nand U1808 (N_1808,In_388,In_201);
and U1809 (N_1809,In_750,In_379);
or U1810 (N_1810,In_436,In_682);
nand U1811 (N_1811,In_224,In_398);
and U1812 (N_1812,In_553,In_255);
nor U1813 (N_1813,In_863,In_586);
nor U1814 (N_1814,In_911,In_696);
nand U1815 (N_1815,In_658,In_249);
nand U1816 (N_1816,In_953,In_580);
nor U1817 (N_1817,In_184,In_215);
xnor U1818 (N_1818,In_678,In_681);
nand U1819 (N_1819,In_691,In_969);
xor U1820 (N_1820,In_455,In_399);
nor U1821 (N_1821,In_389,In_537);
nor U1822 (N_1822,In_565,In_64);
or U1823 (N_1823,In_648,In_871);
and U1824 (N_1824,In_570,In_411);
and U1825 (N_1825,In_941,In_565);
or U1826 (N_1826,In_699,In_954);
and U1827 (N_1827,In_149,In_205);
and U1828 (N_1828,In_15,In_333);
and U1829 (N_1829,In_439,In_234);
or U1830 (N_1830,In_389,In_556);
and U1831 (N_1831,In_916,In_927);
nand U1832 (N_1832,In_76,In_641);
xnor U1833 (N_1833,In_83,In_697);
and U1834 (N_1834,In_475,In_800);
nor U1835 (N_1835,In_700,In_202);
nand U1836 (N_1836,In_722,In_98);
nand U1837 (N_1837,In_325,In_224);
nand U1838 (N_1838,In_287,In_15);
or U1839 (N_1839,In_387,In_133);
nand U1840 (N_1840,In_235,In_110);
and U1841 (N_1841,In_349,In_587);
and U1842 (N_1842,In_338,In_551);
or U1843 (N_1843,In_869,In_615);
and U1844 (N_1844,In_780,In_739);
nand U1845 (N_1845,In_716,In_450);
or U1846 (N_1846,In_192,In_820);
or U1847 (N_1847,In_144,In_451);
xor U1848 (N_1848,In_343,In_766);
and U1849 (N_1849,In_794,In_764);
or U1850 (N_1850,In_527,In_912);
or U1851 (N_1851,In_138,In_213);
nand U1852 (N_1852,In_563,In_470);
and U1853 (N_1853,In_600,In_508);
or U1854 (N_1854,In_447,In_517);
nor U1855 (N_1855,In_231,In_563);
nor U1856 (N_1856,In_46,In_662);
nor U1857 (N_1857,In_624,In_756);
or U1858 (N_1858,In_885,In_596);
and U1859 (N_1859,In_276,In_715);
and U1860 (N_1860,In_595,In_149);
or U1861 (N_1861,In_496,In_292);
xor U1862 (N_1862,In_843,In_376);
nand U1863 (N_1863,In_666,In_665);
and U1864 (N_1864,In_34,In_603);
or U1865 (N_1865,In_696,In_346);
and U1866 (N_1866,In_982,In_754);
nor U1867 (N_1867,In_289,In_685);
nand U1868 (N_1868,In_820,In_133);
nor U1869 (N_1869,In_871,In_876);
and U1870 (N_1870,In_80,In_23);
nand U1871 (N_1871,In_62,In_253);
nand U1872 (N_1872,In_651,In_358);
nor U1873 (N_1873,In_709,In_384);
nand U1874 (N_1874,In_244,In_371);
and U1875 (N_1875,In_245,In_753);
and U1876 (N_1876,In_427,In_314);
and U1877 (N_1877,In_893,In_309);
or U1878 (N_1878,In_902,In_331);
nand U1879 (N_1879,In_742,In_508);
or U1880 (N_1880,In_287,In_996);
nor U1881 (N_1881,In_67,In_408);
nand U1882 (N_1882,In_254,In_43);
and U1883 (N_1883,In_11,In_969);
and U1884 (N_1884,In_783,In_687);
nand U1885 (N_1885,In_713,In_353);
and U1886 (N_1886,In_653,In_695);
and U1887 (N_1887,In_412,In_281);
and U1888 (N_1888,In_649,In_730);
nor U1889 (N_1889,In_720,In_890);
or U1890 (N_1890,In_448,In_664);
nand U1891 (N_1891,In_510,In_949);
nand U1892 (N_1892,In_856,In_87);
nand U1893 (N_1893,In_934,In_440);
nor U1894 (N_1894,In_585,In_670);
and U1895 (N_1895,In_1,In_942);
nand U1896 (N_1896,In_160,In_871);
nand U1897 (N_1897,In_734,In_205);
and U1898 (N_1898,In_701,In_342);
nor U1899 (N_1899,In_684,In_310);
nor U1900 (N_1900,In_721,In_374);
xor U1901 (N_1901,In_911,In_77);
nand U1902 (N_1902,In_219,In_127);
nor U1903 (N_1903,In_736,In_834);
or U1904 (N_1904,In_431,In_773);
or U1905 (N_1905,In_458,In_229);
or U1906 (N_1906,In_11,In_891);
nor U1907 (N_1907,In_561,In_90);
and U1908 (N_1908,In_701,In_809);
and U1909 (N_1909,In_625,In_342);
nand U1910 (N_1910,In_917,In_180);
and U1911 (N_1911,In_447,In_20);
nand U1912 (N_1912,In_969,In_80);
and U1913 (N_1913,In_55,In_181);
or U1914 (N_1914,In_935,In_243);
nand U1915 (N_1915,In_835,In_904);
or U1916 (N_1916,In_618,In_401);
nand U1917 (N_1917,In_854,In_334);
nand U1918 (N_1918,In_71,In_845);
nand U1919 (N_1919,In_257,In_531);
or U1920 (N_1920,In_196,In_776);
or U1921 (N_1921,In_475,In_481);
nor U1922 (N_1922,In_92,In_458);
or U1923 (N_1923,In_894,In_256);
and U1924 (N_1924,In_990,In_76);
nor U1925 (N_1925,In_20,In_654);
or U1926 (N_1926,In_861,In_379);
nand U1927 (N_1927,In_289,In_527);
nand U1928 (N_1928,In_800,In_538);
nand U1929 (N_1929,In_104,In_845);
nor U1930 (N_1930,In_508,In_136);
or U1931 (N_1931,In_886,In_770);
xor U1932 (N_1932,In_910,In_384);
and U1933 (N_1933,In_388,In_61);
or U1934 (N_1934,In_97,In_752);
or U1935 (N_1935,In_859,In_395);
nand U1936 (N_1936,In_142,In_297);
nor U1937 (N_1937,In_539,In_794);
or U1938 (N_1938,In_330,In_560);
nand U1939 (N_1939,In_940,In_191);
nand U1940 (N_1940,In_321,In_748);
nand U1941 (N_1941,In_707,In_477);
and U1942 (N_1942,In_196,In_252);
nand U1943 (N_1943,In_338,In_872);
or U1944 (N_1944,In_665,In_437);
nand U1945 (N_1945,In_840,In_810);
or U1946 (N_1946,In_537,In_228);
and U1947 (N_1947,In_958,In_482);
or U1948 (N_1948,In_612,In_435);
xor U1949 (N_1949,In_710,In_752);
or U1950 (N_1950,In_158,In_219);
nor U1951 (N_1951,In_184,In_153);
nor U1952 (N_1952,In_566,In_156);
or U1953 (N_1953,In_717,In_351);
nor U1954 (N_1954,In_810,In_248);
nor U1955 (N_1955,In_567,In_800);
and U1956 (N_1956,In_898,In_95);
and U1957 (N_1957,In_690,In_112);
or U1958 (N_1958,In_232,In_543);
nand U1959 (N_1959,In_928,In_246);
nand U1960 (N_1960,In_773,In_528);
nand U1961 (N_1961,In_218,In_677);
nand U1962 (N_1962,In_560,In_747);
or U1963 (N_1963,In_746,In_892);
nor U1964 (N_1964,In_582,In_402);
or U1965 (N_1965,In_811,In_575);
and U1966 (N_1966,In_213,In_93);
nor U1967 (N_1967,In_227,In_457);
nor U1968 (N_1968,In_982,In_133);
xor U1969 (N_1969,In_330,In_523);
nand U1970 (N_1970,In_290,In_396);
and U1971 (N_1971,In_206,In_395);
nor U1972 (N_1972,In_434,In_123);
xor U1973 (N_1973,In_678,In_569);
nor U1974 (N_1974,In_175,In_870);
nand U1975 (N_1975,In_155,In_79);
nand U1976 (N_1976,In_658,In_185);
or U1977 (N_1977,In_852,In_966);
nand U1978 (N_1978,In_756,In_75);
or U1979 (N_1979,In_735,In_707);
nand U1980 (N_1980,In_135,In_284);
nand U1981 (N_1981,In_528,In_26);
or U1982 (N_1982,In_109,In_222);
nor U1983 (N_1983,In_502,In_923);
xnor U1984 (N_1984,In_324,In_828);
nand U1985 (N_1985,In_335,In_357);
or U1986 (N_1986,In_1,In_976);
and U1987 (N_1987,In_366,In_820);
nand U1988 (N_1988,In_889,In_751);
and U1989 (N_1989,In_818,In_687);
nor U1990 (N_1990,In_93,In_990);
or U1991 (N_1991,In_314,In_867);
xor U1992 (N_1992,In_834,In_488);
xor U1993 (N_1993,In_865,In_254);
and U1994 (N_1994,In_780,In_75);
xnor U1995 (N_1995,In_35,In_986);
nor U1996 (N_1996,In_854,In_111);
or U1997 (N_1997,In_865,In_26);
or U1998 (N_1998,In_445,In_362);
nand U1999 (N_1999,In_198,In_840);
nor U2000 (N_2000,In_741,In_37);
xor U2001 (N_2001,In_521,In_69);
and U2002 (N_2002,In_390,In_19);
or U2003 (N_2003,In_693,In_460);
nand U2004 (N_2004,In_590,In_823);
and U2005 (N_2005,In_770,In_710);
and U2006 (N_2006,In_149,In_722);
or U2007 (N_2007,In_130,In_816);
and U2008 (N_2008,In_535,In_607);
or U2009 (N_2009,In_117,In_271);
nand U2010 (N_2010,In_376,In_850);
or U2011 (N_2011,In_3,In_291);
and U2012 (N_2012,In_435,In_585);
or U2013 (N_2013,In_674,In_797);
and U2014 (N_2014,In_401,In_893);
nand U2015 (N_2015,In_652,In_725);
or U2016 (N_2016,In_144,In_377);
nand U2017 (N_2017,In_502,In_10);
nor U2018 (N_2018,In_369,In_611);
or U2019 (N_2019,In_200,In_778);
and U2020 (N_2020,In_937,In_705);
nor U2021 (N_2021,In_250,In_927);
or U2022 (N_2022,In_772,In_936);
or U2023 (N_2023,In_855,In_188);
xnor U2024 (N_2024,In_286,In_130);
or U2025 (N_2025,In_302,In_35);
nor U2026 (N_2026,In_331,In_895);
and U2027 (N_2027,In_770,In_481);
or U2028 (N_2028,In_542,In_574);
or U2029 (N_2029,In_646,In_292);
nand U2030 (N_2030,In_160,In_135);
and U2031 (N_2031,In_679,In_166);
and U2032 (N_2032,In_56,In_72);
or U2033 (N_2033,In_433,In_512);
and U2034 (N_2034,In_949,In_486);
nor U2035 (N_2035,In_187,In_23);
and U2036 (N_2036,In_518,In_328);
nor U2037 (N_2037,In_360,In_780);
nand U2038 (N_2038,In_646,In_120);
nor U2039 (N_2039,In_283,In_714);
or U2040 (N_2040,In_30,In_827);
and U2041 (N_2041,In_951,In_171);
or U2042 (N_2042,In_885,In_131);
and U2043 (N_2043,In_925,In_923);
nand U2044 (N_2044,In_182,In_361);
nor U2045 (N_2045,In_167,In_777);
or U2046 (N_2046,In_423,In_867);
nand U2047 (N_2047,In_294,In_940);
nor U2048 (N_2048,In_665,In_172);
and U2049 (N_2049,In_713,In_586);
nor U2050 (N_2050,In_954,In_550);
nor U2051 (N_2051,In_865,In_18);
nor U2052 (N_2052,In_644,In_491);
nand U2053 (N_2053,In_576,In_964);
or U2054 (N_2054,In_599,In_285);
and U2055 (N_2055,In_360,In_853);
nor U2056 (N_2056,In_241,In_185);
nand U2057 (N_2057,In_979,In_148);
nand U2058 (N_2058,In_246,In_551);
nand U2059 (N_2059,In_632,In_951);
or U2060 (N_2060,In_647,In_692);
nand U2061 (N_2061,In_608,In_300);
and U2062 (N_2062,In_297,In_433);
nand U2063 (N_2063,In_671,In_541);
or U2064 (N_2064,In_250,In_993);
nand U2065 (N_2065,In_826,In_113);
nand U2066 (N_2066,In_987,In_369);
and U2067 (N_2067,In_570,In_610);
nand U2068 (N_2068,In_322,In_612);
nand U2069 (N_2069,In_125,In_100);
nand U2070 (N_2070,In_726,In_381);
or U2071 (N_2071,In_170,In_108);
nand U2072 (N_2072,In_865,In_379);
or U2073 (N_2073,In_743,In_994);
nor U2074 (N_2074,In_998,In_917);
or U2075 (N_2075,In_409,In_246);
or U2076 (N_2076,In_311,In_163);
nor U2077 (N_2077,In_304,In_384);
nand U2078 (N_2078,In_632,In_917);
nor U2079 (N_2079,In_770,In_702);
nor U2080 (N_2080,In_618,In_9);
nor U2081 (N_2081,In_134,In_963);
nand U2082 (N_2082,In_498,In_133);
nor U2083 (N_2083,In_681,In_819);
or U2084 (N_2084,In_323,In_887);
or U2085 (N_2085,In_911,In_155);
nor U2086 (N_2086,In_930,In_330);
or U2087 (N_2087,In_952,In_715);
nor U2088 (N_2088,In_397,In_339);
nor U2089 (N_2089,In_408,In_609);
nor U2090 (N_2090,In_369,In_138);
and U2091 (N_2091,In_730,In_575);
nor U2092 (N_2092,In_707,In_343);
nand U2093 (N_2093,In_366,In_500);
nor U2094 (N_2094,In_45,In_973);
nor U2095 (N_2095,In_813,In_31);
nand U2096 (N_2096,In_8,In_180);
xor U2097 (N_2097,In_149,In_894);
nand U2098 (N_2098,In_657,In_634);
nor U2099 (N_2099,In_218,In_383);
or U2100 (N_2100,In_337,In_113);
nor U2101 (N_2101,In_403,In_165);
and U2102 (N_2102,In_889,In_626);
or U2103 (N_2103,In_593,In_852);
nand U2104 (N_2104,In_879,In_898);
and U2105 (N_2105,In_381,In_370);
and U2106 (N_2106,In_704,In_998);
or U2107 (N_2107,In_130,In_867);
and U2108 (N_2108,In_775,In_93);
or U2109 (N_2109,In_573,In_787);
and U2110 (N_2110,In_370,In_929);
and U2111 (N_2111,In_522,In_344);
or U2112 (N_2112,In_330,In_574);
or U2113 (N_2113,In_236,In_248);
or U2114 (N_2114,In_493,In_865);
and U2115 (N_2115,In_183,In_532);
nand U2116 (N_2116,In_697,In_191);
nor U2117 (N_2117,In_806,In_287);
nor U2118 (N_2118,In_225,In_923);
nand U2119 (N_2119,In_66,In_585);
or U2120 (N_2120,In_878,In_556);
nor U2121 (N_2121,In_923,In_833);
nand U2122 (N_2122,In_102,In_592);
nor U2123 (N_2123,In_904,In_930);
nand U2124 (N_2124,In_500,In_650);
nor U2125 (N_2125,In_980,In_745);
and U2126 (N_2126,In_832,In_482);
nand U2127 (N_2127,In_921,In_785);
xnor U2128 (N_2128,In_601,In_99);
xor U2129 (N_2129,In_959,In_149);
or U2130 (N_2130,In_328,In_511);
nand U2131 (N_2131,In_963,In_475);
nand U2132 (N_2132,In_471,In_308);
and U2133 (N_2133,In_988,In_267);
or U2134 (N_2134,In_30,In_545);
xnor U2135 (N_2135,In_609,In_612);
and U2136 (N_2136,In_542,In_433);
and U2137 (N_2137,In_824,In_571);
and U2138 (N_2138,In_83,In_291);
or U2139 (N_2139,In_161,In_203);
and U2140 (N_2140,In_532,In_694);
nor U2141 (N_2141,In_28,In_120);
nor U2142 (N_2142,In_597,In_341);
xnor U2143 (N_2143,In_507,In_70);
nand U2144 (N_2144,In_857,In_25);
and U2145 (N_2145,In_633,In_646);
and U2146 (N_2146,In_51,In_279);
nor U2147 (N_2147,In_23,In_805);
nor U2148 (N_2148,In_825,In_742);
nand U2149 (N_2149,In_261,In_201);
nand U2150 (N_2150,In_571,In_8);
or U2151 (N_2151,In_613,In_881);
or U2152 (N_2152,In_942,In_167);
nor U2153 (N_2153,In_265,In_570);
nand U2154 (N_2154,In_705,In_852);
and U2155 (N_2155,In_977,In_188);
nor U2156 (N_2156,In_35,In_98);
nor U2157 (N_2157,In_388,In_460);
nand U2158 (N_2158,In_848,In_71);
or U2159 (N_2159,In_727,In_828);
and U2160 (N_2160,In_182,In_564);
nand U2161 (N_2161,In_797,In_698);
nand U2162 (N_2162,In_877,In_832);
or U2163 (N_2163,In_243,In_94);
nor U2164 (N_2164,In_798,In_875);
nor U2165 (N_2165,In_621,In_758);
nand U2166 (N_2166,In_756,In_469);
nand U2167 (N_2167,In_699,In_141);
nand U2168 (N_2168,In_273,In_236);
or U2169 (N_2169,In_763,In_284);
and U2170 (N_2170,In_232,In_753);
nand U2171 (N_2171,In_472,In_196);
nor U2172 (N_2172,In_681,In_18);
or U2173 (N_2173,In_707,In_113);
nor U2174 (N_2174,In_173,In_833);
xnor U2175 (N_2175,In_672,In_864);
and U2176 (N_2176,In_974,In_357);
and U2177 (N_2177,In_613,In_982);
nor U2178 (N_2178,In_996,In_6);
nor U2179 (N_2179,In_581,In_202);
or U2180 (N_2180,In_308,In_53);
and U2181 (N_2181,In_727,In_79);
nand U2182 (N_2182,In_485,In_205);
and U2183 (N_2183,In_796,In_463);
or U2184 (N_2184,In_869,In_209);
nor U2185 (N_2185,In_942,In_741);
or U2186 (N_2186,In_322,In_54);
and U2187 (N_2187,In_40,In_315);
nor U2188 (N_2188,In_722,In_813);
nand U2189 (N_2189,In_103,In_603);
nor U2190 (N_2190,In_60,In_524);
and U2191 (N_2191,In_579,In_170);
nand U2192 (N_2192,In_695,In_161);
nand U2193 (N_2193,In_143,In_108);
and U2194 (N_2194,In_671,In_366);
or U2195 (N_2195,In_44,In_190);
nand U2196 (N_2196,In_298,In_489);
nor U2197 (N_2197,In_360,In_707);
nand U2198 (N_2198,In_551,In_778);
or U2199 (N_2199,In_863,In_57);
and U2200 (N_2200,In_978,In_206);
nand U2201 (N_2201,In_561,In_903);
nor U2202 (N_2202,In_834,In_579);
and U2203 (N_2203,In_911,In_577);
or U2204 (N_2204,In_575,In_700);
nor U2205 (N_2205,In_456,In_856);
and U2206 (N_2206,In_407,In_259);
and U2207 (N_2207,In_592,In_662);
and U2208 (N_2208,In_866,In_425);
nand U2209 (N_2209,In_852,In_893);
nand U2210 (N_2210,In_551,In_496);
and U2211 (N_2211,In_721,In_881);
or U2212 (N_2212,In_839,In_981);
and U2213 (N_2213,In_563,In_190);
nor U2214 (N_2214,In_282,In_911);
nand U2215 (N_2215,In_369,In_373);
nand U2216 (N_2216,In_536,In_844);
nor U2217 (N_2217,In_278,In_306);
and U2218 (N_2218,In_689,In_679);
nand U2219 (N_2219,In_788,In_350);
or U2220 (N_2220,In_429,In_236);
or U2221 (N_2221,In_459,In_20);
or U2222 (N_2222,In_67,In_473);
or U2223 (N_2223,In_265,In_768);
and U2224 (N_2224,In_786,In_451);
or U2225 (N_2225,In_479,In_816);
and U2226 (N_2226,In_745,In_825);
nand U2227 (N_2227,In_852,In_769);
and U2228 (N_2228,In_744,In_864);
and U2229 (N_2229,In_952,In_935);
or U2230 (N_2230,In_165,In_661);
nand U2231 (N_2231,In_649,In_81);
nand U2232 (N_2232,In_724,In_450);
and U2233 (N_2233,In_838,In_726);
or U2234 (N_2234,In_540,In_761);
and U2235 (N_2235,In_593,In_757);
and U2236 (N_2236,In_462,In_918);
or U2237 (N_2237,In_577,In_704);
and U2238 (N_2238,In_690,In_185);
xor U2239 (N_2239,In_62,In_404);
and U2240 (N_2240,In_39,In_211);
and U2241 (N_2241,In_979,In_335);
nor U2242 (N_2242,In_789,In_12);
nand U2243 (N_2243,In_346,In_496);
nand U2244 (N_2244,In_607,In_415);
and U2245 (N_2245,In_757,In_717);
and U2246 (N_2246,In_59,In_427);
nand U2247 (N_2247,In_713,In_781);
or U2248 (N_2248,In_781,In_524);
and U2249 (N_2249,In_379,In_587);
nand U2250 (N_2250,In_814,In_825);
nand U2251 (N_2251,In_815,In_362);
nand U2252 (N_2252,In_227,In_962);
or U2253 (N_2253,In_485,In_491);
and U2254 (N_2254,In_18,In_423);
nor U2255 (N_2255,In_289,In_462);
or U2256 (N_2256,In_576,In_95);
xor U2257 (N_2257,In_976,In_759);
nand U2258 (N_2258,In_663,In_565);
nor U2259 (N_2259,In_75,In_294);
and U2260 (N_2260,In_260,In_454);
and U2261 (N_2261,In_552,In_932);
and U2262 (N_2262,In_47,In_985);
or U2263 (N_2263,In_613,In_896);
nor U2264 (N_2264,In_683,In_225);
or U2265 (N_2265,In_530,In_64);
or U2266 (N_2266,In_887,In_416);
and U2267 (N_2267,In_185,In_266);
nor U2268 (N_2268,In_746,In_379);
nor U2269 (N_2269,In_560,In_45);
nor U2270 (N_2270,In_133,In_331);
or U2271 (N_2271,In_217,In_178);
nor U2272 (N_2272,In_479,In_655);
nor U2273 (N_2273,In_398,In_761);
and U2274 (N_2274,In_778,In_690);
nand U2275 (N_2275,In_224,In_183);
nor U2276 (N_2276,In_300,In_152);
xor U2277 (N_2277,In_258,In_47);
or U2278 (N_2278,In_280,In_601);
or U2279 (N_2279,In_8,In_275);
nand U2280 (N_2280,In_646,In_248);
or U2281 (N_2281,In_580,In_762);
or U2282 (N_2282,In_448,In_369);
nor U2283 (N_2283,In_942,In_278);
or U2284 (N_2284,In_537,In_890);
nand U2285 (N_2285,In_667,In_118);
nand U2286 (N_2286,In_855,In_865);
nand U2287 (N_2287,In_340,In_849);
and U2288 (N_2288,In_132,In_508);
or U2289 (N_2289,In_709,In_549);
xnor U2290 (N_2290,In_78,In_123);
nand U2291 (N_2291,In_471,In_980);
nor U2292 (N_2292,In_708,In_303);
or U2293 (N_2293,In_298,In_571);
or U2294 (N_2294,In_953,In_616);
nand U2295 (N_2295,In_206,In_994);
nor U2296 (N_2296,In_169,In_341);
nor U2297 (N_2297,In_705,In_225);
nor U2298 (N_2298,In_927,In_123);
nor U2299 (N_2299,In_116,In_276);
and U2300 (N_2300,In_58,In_343);
and U2301 (N_2301,In_726,In_949);
nand U2302 (N_2302,In_617,In_529);
or U2303 (N_2303,In_543,In_715);
nand U2304 (N_2304,In_323,In_104);
and U2305 (N_2305,In_385,In_559);
nand U2306 (N_2306,In_933,In_305);
or U2307 (N_2307,In_687,In_883);
and U2308 (N_2308,In_716,In_432);
and U2309 (N_2309,In_215,In_782);
and U2310 (N_2310,In_555,In_774);
and U2311 (N_2311,In_467,In_388);
and U2312 (N_2312,In_514,In_732);
nand U2313 (N_2313,In_225,In_476);
nand U2314 (N_2314,In_745,In_104);
nand U2315 (N_2315,In_451,In_318);
and U2316 (N_2316,In_649,In_523);
nor U2317 (N_2317,In_185,In_868);
or U2318 (N_2318,In_281,In_144);
nor U2319 (N_2319,In_870,In_937);
and U2320 (N_2320,In_692,In_901);
or U2321 (N_2321,In_282,In_831);
nand U2322 (N_2322,In_404,In_573);
or U2323 (N_2323,In_444,In_339);
nand U2324 (N_2324,In_149,In_612);
nor U2325 (N_2325,In_420,In_166);
nand U2326 (N_2326,In_765,In_406);
nand U2327 (N_2327,In_786,In_135);
nor U2328 (N_2328,In_157,In_892);
nand U2329 (N_2329,In_558,In_568);
and U2330 (N_2330,In_746,In_733);
or U2331 (N_2331,In_843,In_131);
nor U2332 (N_2332,In_257,In_614);
and U2333 (N_2333,In_298,In_497);
and U2334 (N_2334,In_515,In_409);
and U2335 (N_2335,In_31,In_617);
and U2336 (N_2336,In_915,In_489);
nand U2337 (N_2337,In_400,In_571);
nor U2338 (N_2338,In_44,In_987);
nand U2339 (N_2339,In_59,In_614);
or U2340 (N_2340,In_464,In_109);
nor U2341 (N_2341,In_727,In_628);
nor U2342 (N_2342,In_814,In_551);
or U2343 (N_2343,In_279,In_225);
nor U2344 (N_2344,In_353,In_228);
nand U2345 (N_2345,In_35,In_226);
nand U2346 (N_2346,In_279,In_131);
or U2347 (N_2347,In_930,In_863);
xor U2348 (N_2348,In_543,In_563);
nand U2349 (N_2349,In_396,In_681);
and U2350 (N_2350,In_814,In_473);
and U2351 (N_2351,In_720,In_961);
nor U2352 (N_2352,In_351,In_492);
nor U2353 (N_2353,In_188,In_310);
nor U2354 (N_2354,In_855,In_130);
nand U2355 (N_2355,In_574,In_94);
and U2356 (N_2356,In_930,In_698);
nand U2357 (N_2357,In_315,In_238);
nor U2358 (N_2358,In_111,In_120);
nor U2359 (N_2359,In_403,In_731);
nor U2360 (N_2360,In_975,In_449);
xor U2361 (N_2361,In_656,In_360);
nor U2362 (N_2362,In_221,In_736);
and U2363 (N_2363,In_304,In_5);
nand U2364 (N_2364,In_926,In_574);
and U2365 (N_2365,In_893,In_661);
nor U2366 (N_2366,In_538,In_598);
or U2367 (N_2367,In_35,In_660);
nor U2368 (N_2368,In_14,In_721);
nor U2369 (N_2369,In_199,In_554);
or U2370 (N_2370,In_247,In_376);
and U2371 (N_2371,In_699,In_105);
nor U2372 (N_2372,In_709,In_961);
nor U2373 (N_2373,In_81,In_214);
nand U2374 (N_2374,In_468,In_271);
nor U2375 (N_2375,In_650,In_72);
or U2376 (N_2376,In_805,In_651);
nor U2377 (N_2377,In_196,In_537);
or U2378 (N_2378,In_453,In_990);
nand U2379 (N_2379,In_28,In_813);
nor U2380 (N_2380,In_17,In_751);
and U2381 (N_2381,In_499,In_111);
nor U2382 (N_2382,In_486,In_914);
nand U2383 (N_2383,In_50,In_552);
or U2384 (N_2384,In_151,In_208);
nor U2385 (N_2385,In_154,In_474);
nor U2386 (N_2386,In_399,In_34);
or U2387 (N_2387,In_108,In_945);
and U2388 (N_2388,In_396,In_386);
nand U2389 (N_2389,In_151,In_436);
and U2390 (N_2390,In_271,In_957);
or U2391 (N_2391,In_578,In_722);
or U2392 (N_2392,In_504,In_522);
or U2393 (N_2393,In_105,In_429);
nand U2394 (N_2394,In_723,In_830);
or U2395 (N_2395,In_724,In_20);
nor U2396 (N_2396,In_513,In_112);
nor U2397 (N_2397,In_760,In_114);
nor U2398 (N_2398,In_353,In_201);
and U2399 (N_2399,In_965,In_798);
or U2400 (N_2400,In_380,In_344);
and U2401 (N_2401,In_487,In_898);
nor U2402 (N_2402,In_266,In_598);
nor U2403 (N_2403,In_803,In_158);
and U2404 (N_2404,In_344,In_213);
nand U2405 (N_2405,In_260,In_605);
nand U2406 (N_2406,In_830,In_171);
nor U2407 (N_2407,In_65,In_248);
nor U2408 (N_2408,In_573,In_59);
and U2409 (N_2409,In_19,In_519);
or U2410 (N_2410,In_671,In_816);
nor U2411 (N_2411,In_601,In_93);
nor U2412 (N_2412,In_224,In_874);
nand U2413 (N_2413,In_21,In_164);
nor U2414 (N_2414,In_479,In_275);
and U2415 (N_2415,In_23,In_684);
nor U2416 (N_2416,In_60,In_202);
nor U2417 (N_2417,In_192,In_683);
nor U2418 (N_2418,In_855,In_159);
nor U2419 (N_2419,In_961,In_334);
nand U2420 (N_2420,In_560,In_579);
and U2421 (N_2421,In_449,In_191);
nor U2422 (N_2422,In_418,In_688);
or U2423 (N_2423,In_587,In_948);
nand U2424 (N_2424,In_586,In_21);
and U2425 (N_2425,In_32,In_395);
or U2426 (N_2426,In_158,In_162);
xnor U2427 (N_2427,In_927,In_292);
nor U2428 (N_2428,In_603,In_762);
nand U2429 (N_2429,In_890,In_304);
nor U2430 (N_2430,In_725,In_735);
and U2431 (N_2431,In_665,In_104);
or U2432 (N_2432,In_826,In_997);
nor U2433 (N_2433,In_100,In_601);
and U2434 (N_2434,In_100,In_603);
and U2435 (N_2435,In_54,In_272);
nor U2436 (N_2436,In_658,In_376);
nand U2437 (N_2437,In_450,In_398);
nand U2438 (N_2438,In_703,In_103);
and U2439 (N_2439,In_500,In_709);
and U2440 (N_2440,In_784,In_231);
and U2441 (N_2441,In_646,In_461);
or U2442 (N_2442,In_673,In_442);
and U2443 (N_2443,In_412,In_490);
and U2444 (N_2444,In_583,In_218);
and U2445 (N_2445,In_769,In_643);
nand U2446 (N_2446,In_866,In_276);
nand U2447 (N_2447,In_607,In_429);
nor U2448 (N_2448,In_584,In_564);
nor U2449 (N_2449,In_813,In_682);
nand U2450 (N_2450,In_237,In_834);
nor U2451 (N_2451,In_713,In_862);
nand U2452 (N_2452,In_879,In_449);
or U2453 (N_2453,In_81,In_4);
nand U2454 (N_2454,In_231,In_949);
nor U2455 (N_2455,In_488,In_918);
and U2456 (N_2456,In_207,In_109);
or U2457 (N_2457,In_416,In_179);
and U2458 (N_2458,In_485,In_403);
and U2459 (N_2459,In_601,In_780);
nor U2460 (N_2460,In_154,In_394);
or U2461 (N_2461,In_314,In_626);
and U2462 (N_2462,In_116,In_97);
nand U2463 (N_2463,In_141,In_958);
nand U2464 (N_2464,In_403,In_424);
nand U2465 (N_2465,In_414,In_917);
and U2466 (N_2466,In_788,In_169);
or U2467 (N_2467,In_706,In_59);
and U2468 (N_2468,In_401,In_253);
nand U2469 (N_2469,In_421,In_213);
nand U2470 (N_2470,In_347,In_465);
or U2471 (N_2471,In_738,In_517);
and U2472 (N_2472,In_689,In_94);
nand U2473 (N_2473,In_427,In_594);
nand U2474 (N_2474,In_282,In_580);
nand U2475 (N_2475,In_873,In_433);
and U2476 (N_2476,In_564,In_218);
nor U2477 (N_2477,In_599,In_754);
nor U2478 (N_2478,In_35,In_603);
and U2479 (N_2479,In_106,In_879);
nor U2480 (N_2480,In_406,In_55);
and U2481 (N_2481,In_214,In_508);
nand U2482 (N_2482,In_312,In_863);
nand U2483 (N_2483,In_672,In_313);
or U2484 (N_2484,In_740,In_27);
and U2485 (N_2485,In_393,In_352);
nand U2486 (N_2486,In_85,In_434);
nand U2487 (N_2487,In_777,In_519);
and U2488 (N_2488,In_117,In_46);
nor U2489 (N_2489,In_669,In_388);
or U2490 (N_2490,In_304,In_319);
and U2491 (N_2491,In_603,In_243);
and U2492 (N_2492,In_958,In_576);
and U2493 (N_2493,In_923,In_51);
nand U2494 (N_2494,In_873,In_941);
and U2495 (N_2495,In_968,In_874);
nor U2496 (N_2496,In_897,In_353);
and U2497 (N_2497,In_621,In_762);
or U2498 (N_2498,In_792,In_159);
nand U2499 (N_2499,In_804,In_582);
or U2500 (N_2500,In_835,In_155);
and U2501 (N_2501,In_44,In_571);
nand U2502 (N_2502,In_853,In_977);
nand U2503 (N_2503,In_351,In_584);
nor U2504 (N_2504,In_899,In_462);
nor U2505 (N_2505,In_620,In_499);
or U2506 (N_2506,In_166,In_161);
and U2507 (N_2507,In_652,In_388);
xor U2508 (N_2508,In_516,In_562);
nand U2509 (N_2509,In_936,In_659);
or U2510 (N_2510,In_797,In_265);
nand U2511 (N_2511,In_671,In_172);
nand U2512 (N_2512,In_216,In_438);
nand U2513 (N_2513,In_102,In_207);
or U2514 (N_2514,In_787,In_768);
nor U2515 (N_2515,In_281,In_135);
nand U2516 (N_2516,In_638,In_3);
and U2517 (N_2517,In_274,In_181);
nand U2518 (N_2518,In_879,In_674);
or U2519 (N_2519,In_183,In_85);
and U2520 (N_2520,In_764,In_49);
or U2521 (N_2521,In_402,In_941);
nand U2522 (N_2522,In_154,In_89);
nor U2523 (N_2523,In_528,In_851);
nand U2524 (N_2524,In_651,In_160);
nand U2525 (N_2525,In_191,In_368);
nand U2526 (N_2526,In_112,In_407);
nand U2527 (N_2527,In_60,In_331);
and U2528 (N_2528,In_2,In_855);
nand U2529 (N_2529,In_59,In_28);
and U2530 (N_2530,In_621,In_548);
nand U2531 (N_2531,In_872,In_250);
xor U2532 (N_2532,In_881,In_142);
nor U2533 (N_2533,In_941,In_790);
nor U2534 (N_2534,In_1,In_431);
nand U2535 (N_2535,In_758,In_481);
or U2536 (N_2536,In_843,In_637);
nand U2537 (N_2537,In_250,In_857);
nand U2538 (N_2538,In_334,In_685);
and U2539 (N_2539,In_490,In_71);
nand U2540 (N_2540,In_680,In_132);
and U2541 (N_2541,In_648,In_203);
and U2542 (N_2542,In_279,In_498);
nand U2543 (N_2543,In_556,In_929);
or U2544 (N_2544,In_510,In_759);
and U2545 (N_2545,In_543,In_580);
nor U2546 (N_2546,In_288,In_931);
or U2547 (N_2547,In_577,In_574);
and U2548 (N_2548,In_518,In_179);
or U2549 (N_2549,In_349,In_389);
nor U2550 (N_2550,In_713,In_764);
xor U2551 (N_2551,In_236,In_904);
nor U2552 (N_2552,In_798,In_938);
and U2553 (N_2553,In_710,In_99);
or U2554 (N_2554,In_613,In_582);
nor U2555 (N_2555,In_957,In_858);
and U2556 (N_2556,In_293,In_25);
and U2557 (N_2557,In_829,In_372);
nand U2558 (N_2558,In_526,In_650);
and U2559 (N_2559,In_582,In_179);
and U2560 (N_2560,In_509,In_728);
or U2561 (N_2561,In_759,In_745);
or U2562 (N_2562,In_374,In_264);
and U2563 (N_2563,In_702,In_725);
and U2564 (N_2564,In_166,In_402);
nor U2565 (N_2565,In_873,In_47);
and U2566 (N_2566,In_745,In_84);
or U2567 (N_2567,In_936,In_581);
and U2568 (N_2568,In_954,In_49);
nand U2569 (N_2569,In_251,In_448);
or U2570 (N_2570,In_832,In_615);
nor U2571 (N_2571,In_377,In_988);
nor U2572 (N_2572,In_330,In_916);
nand U2573 (N_2573,In_830,In_86);
nor U2574 (N_2574,In_374,In_315);
nand U2575 (N_2575,In_405,In_172);
nand U2576 (N_2576,In_842,In_200);
or U2577 (N_2577,In_556,In_425);
and U2578 (N_2578,In_856,In_376);
xor U2579 (N_2579,In_458,In_558);
xor U2580 (N_2580,In_393,In_905);
and U2581 (N_2581,In_300,In_82);
or U2582 (N_2582,In_622,In_767);
or U2583 (N_2583,In_820,In_869);
nor U2584 (N_2584,In_785,In_383);
nor U2585 (N_2585,In_791,In_909);
and U2586 (N_2586,In_318,In_57);
nand U2587 (N_2587,In_672,In_907);
and U2588 (N_2588,In_695,In_856);
nand U2589 (N_2589,In_655,In_326);
or U2590 (N_2590,In_297,In_936);
nand U2591 (N_2591,In_426,In_970);
or U2592 (N_2592,In_247,In_875);
or U2593 (N_2593,In_844,In_487);
and U2594 (N_2594,In_636,In_398);
and U2595 (N_2595,In_963,In_574);
nor U2596 (N_2596,In_51,In_529);
nand U2597 (N_2597,In_527,In_93);
nor U2598 (N_2598,In_448,In_841);
and U2599 (N_2599,In_772,In_218);
nor U2600 (N_2600,In_276,In_65);
nand U2601 (N_2601,In_784,In_287);
xnor U2602 (N_2602,In_881,In_188);
or U2603 (N_2603,In_656,In_615);
and U2604 (N_2604,In_491,In_55);
and U2605 (N_2605,In_958,In_403);
nand U2606 (N_2606,In_288,In_350);
nand U2607 (N_2607,In_182,In_693);
and U2608 (N_2608,In_341,In_551);
or U2609 (N_2609,In_522,In_680);
or U2610 (N_2610,In_897,In_217);
nor U2611 (N_2611,In_360,In_117);
xor U2612 (N_2612,In_918,In_17);
nand U2613 (N_2613,In_300,In_935);
or U2614 (N_2614,In_178,In_271);
nor U2615 (N_2615,In_635,In_461);
nand U2616 (N_2616,In_816,In_414);
nor U2617 (N_2617,In_757,In_867);
nand U2618 (N_2618,In_702,In_114);
nand U2619 (N_2619,In_323,In_967);
and U2620 (N_2620,In_407,In_197);
and U2621 (N_2621,In_664,In_334);
or U2622 (N_2622,In_265,In_172);
or U2623 (N_2623,In_176,In_693);
or U2624 (N_2624,In_905,In_794);
nand U2625 (N_2625,In_443,In_338);
nand U2626 (N_2626,In_686,In_101);
or U2627 (N_2627,In_139,In_551);
nor U2628 (N_2628,In_953,In_829);
or U2629 (N_2629,In_633,In_460);
nor U2630 (N_2630,In_6,In_292);
nor U2631 (N_2631,In_163,In_329);
nor U2632 (N_2632,In_520,In_113);
nand U2633 (N_2633,In_721,In_201);
nor U2634 (N_2634,In_680,In_832);
nor U2635 (N_2635,In_934,In_783);
nor U2636 (N_2636,In_246,In_749);
nand U2637 (N_2637,In_479,In_772);
and U2638 (N_2638,In_259,In_534);
nand U2639 (N_2639,In_187,In_459);
or U2640 (N_2640,In_834,In_852);
nand U2641 (N_2641,In_446,In_596);
nor U2642 (N_2642,In_688,In_566);
nand U2643 (N_2643,In_536,In_64);
or U2644 (N_2644,In_726,In_456);
and U2645 (N_2645,In_294,In_959);
nand U2646 (N_2646,In_383,In_475);
and U2647 (N_2647,In_712,In_503);
or U2648 (N_2648,In_524,In_819);
and U2649 (N_2649,In_531,In_165);
and U2650 (N_2650,In_983,In_799);
nor U2651 (N_2651,In_37,In_827);
nand U2652 (N_2652,In_27,In_704);
nor U2653 (N_2653,In_275,In_57);
or U2654 (N_2654,In_224,In_975);
nand U2655 (N_2655,In_82,In_651);
and U2656 (N_2656,In_551,In_513);
and U2657 (N_2657,In_657,In_676);
nor U2658 (N_2658,In_506,In_263);
or U2659 (N_2659,In_618,In_443);
and U2660 (N_2660,In_109,In_794);
and U2661 (N_2661,In_317,In_498);
and U2662 (N_2662,In_602,In_921);
nor U2663 (N_2663,In_929,In_967);
or U2664 (N_2664,In_492,In_196);
nand U2665 (N_2665,In_91,In_509);
nand U2666 (N_2666,In_791,In_142);
and U2667 (N_2667,In_527,In_843);
nand U2668 (N_2668,In_59,In_431);
nor U2669 (N_2669,In_10,In_207);
nand U2670 (N_2670,In_872,In_503);
xnor U2671 (N_2671,In_675,In_159);
nor U2672 (N_2672,In_405,In_600);
nand U2673 (N_2673,In_769,In_375);
or U2674 (N_2674,In_876,In_46);
nand U2675 (N_2675,In_971,In_277);
and U2676 (N_2676,In_72,In_495);
xor U2677 (N_2677,In_888,In_43);
nand U2678 (N_2678,In_571,In_383);
nor U2679 (N_2679,In_870,In_579);
nand U2680 (N_2680,In_697,In_966);
or U2681 (N_2681,In_376,In_516);
nand U2682 (N_2682,In_336,In_964);
and U2683 (N_2683,In_230,In_481);
or U2684 (N_2684,In_366,In_559);
and U2685 (N_2685,In_204,In_132);
nor U2686 (N_2686,In_143,In_39);
nand U2687 (N_2687,In_603,In_231);
nor U2688 (N_2688,In_50,In_906);
or U2689 (N_2689,In_523,In_722);
nand U2690 (N_2690,In_917,In_553);
and U2691 (N_2691,In_47,In_550);
nand U2692 (N_2692,In_747,In_453);
and U2693 (N_2693,In_365,In_297);
xnor U2694 (N_2694,In_996,In_976);
xor U2695 (N_2695,In_173,In_969);
and U2696 (N_2696,In_493,In_103);
and U2697 (N_2697,In_308,In_581);
or U2698 (N_2698,In_229,In_896);
nand U2699 (N_2699,In_737,In_363);
nand U2700 (N_2700,In_723,In_524);
nand U2701 (N_2701,In_551,In_519);
nand U2702 (N_2702,In_127,In_501);
and U2703 (N_2703,In_686,In_333);
nand U2704 (N_2704,In_557,In_136);
nand U2705 (N_2705,In_26,In_852);
or U2706 (N_2706,In_208,In_350);
and U2707 (N_2707,In_128,In_998);
nor U2708 (N_2708,In_717,In_989);
nand U2709 (N_2709,In_743,In_374);
and U2710 (N_2710,In_827,In_994);
nand U2711 (N_2711,In_915,In_652);
and U2712 (N_2712,In_656,In_943);
or U2713 (N_2713,In_135,In_842);
nor U2714 (N_2714,In_102,In_969);
nand U2715 (N_2715,In_756,In_794);
nor U2716 (N_2716,In_323,In_929);
and U2717 (N_2717,In_424,In_188);
and U2718 (N_2718,In_86,In_682);
and U2719 (N_2719,In_204,In_114);
or U2720 (N_2720,In_579,In_482);
or U2721 (N_2721,In_891,In_127);
and U2722 (N_2722,In_434,In_855);
and U2723 (N_2723,In_911,In_170);
nand U2724 (N_2724,In_648,In_455);
and U2725 (N_2725,In_14,In_247);
xnor U2726 (N_2726,In_82,In_464);
and U2727 (N_2727,In_577,In_7);
and U2728 (N_2728,In_54,In_953);
or U2729 (N_2729,In_951,In_492);
xnor U2730 (N_2730,In_305,In_740);
nor U2731 (N_2731,In_890,In_268);
and U2732 (N_2732,In_340,In_733);
or U2733 (N_2733,In_541,In_749);
nand U2734 (N_2734,In_223,In_105);
nor U2735 (N_2735,In_573,In_589);
and U2736 (N_2736,In_258,In_652);
or U2737 (N_2737,In_682,In_63);
nand U2738 (N_2738,In_172,In_429);
or U2739 (N_2739,In_821,In_729);
or U2740 (N_2740,In_842,In_553);
nand U2741 (N_2741,In_352,In_513);
nand U2742 (N_2742,In_844,In_964);
nand U2743 (N_2743,In_128,In_821);
nor U2744 (N_2744,In_232,In_441);
or U2745 (N_2745,In_488,In_80);
or U2746 (N_2746,In_311,In_881);
nand U2747 (N_2747,In_87,In_889);
and U2748 (N_2748,In_814,In_494);
nor U2749 (N_2749,In_861,In_633);
and U2750 (N_2750,In_540,In_147);
and U2751 (N_2751,In_132,In_709);
nor U2752 (N_2752,In_239,In_280);
nor U2753 (N_2753,In_152,In_374);
nand U2754 (N_2754,In_922,In_396);
and U2755 (N_2755,In_52,In_636);
nor U2756 (N_2756,In_993,In_573);
or U2757 (N_2757,In_268,In_26);
nand U2758 (N_2758,In_469,In_598);
nor U2759 (N_2759,In_511,In_870);
xnor U2760 (N_2760,In_752,In_769);
nand U2761 (N_2761,In_840,In_102);
nor U2762 (N_2762,In_747,In_798);
and U2763 (N_2763,In_795,In_704);
or U2764 (N_2764,In_689,In_335);
and U2765 (N_2765,In_508,In_621);
nand U2766 (N_2766,In_984,In_290);
or U2767 (N_2767,In_383,In_984);
nor U2768 (N_2768,In_823,In_691);
or U2769 (N_2769,In_109,In_90);
nor U2770 (N_2770,In_909,In_721);
nand U2771 (N_2771,In_813,In_304);
nor U2772 (N_2772,In_776,In_654);
or U2773 (N_2773,In_806,In_11);
nand U2774 (N_2774,In_237,In_318);
nor U2775 (N_2775,In_879,In_133);
nand U2776 (N_2776,In_901,In_882);
or U2777 (N_2777,In_577,In_380);
or U2778 (N_2778,In_225,In_604);
or U2779 (N_2779,In_717,In_545);
nand U2780 (N_2780,In_411,In_41);
nand U2781 (N_2781,In_990,In_908);
nand U2782 (N_2782,In_422,In_621);
and U2783 (N_2783,In_998,In_982);
nand U2784 (N_2784,In_118,In_739);
or U2785 (N_2785,In_536,In_577);
or U2786 (N_2786,In_358,In_425);
xor U2787 (N_2787,In_40,In_651);
and U2788 (N_2788,In_385,In_279);
and U2789 (N_2789,In_994,In_924);
xnor U2790 (N_2790,In_302,In_130);
nand U2791 (N_2791,In_62,In_505);
or U2792 (N_2792,In_913,In_98);
xor U2793 (N_2793,In_658,In_312);
and U2794 (N_2794,In_928,In_16);
xor U2795 (N_2795,In_182,In_467);
nand U2796 (N_2796,In_863,In_970);
or U2797 (N_2797,In_32,In_526);
and U2798 (N_2798,In_202,In_43);
or U2799 (N_2799,In_965,In_238);
and U2800 (N_2800,In_520,In_177);
or U2801 (N_2801,In_615,In_334);
nor U2802 (N_2802,In_208,In_817);
nor U2803 (N_2803,In_504,In_137);
and U2804 (N_2804,In_9,In_962);
nor U2805 (N_2805,In_545,In_785);
and U2806 (N_2806,In_270,In_819);
or U2807 (N_2807,In_271,In_805);
and U2808 (N_2808,In_29,In_591);
nand U2809 (N_2809,In_498,In_756);
nor U2810 (N_2810,In_871,In_257);
or U2811 (N_2811,In_937,In_923);
nor U2812 (N_2812,In_229,In_637);
nand U2813 (N_2813,In_673,In_14);
or U2814 (N_2814,In_867,In_920);
nand U2815 (N_2815,In_317,In_741);
nor U2816 (N_2816,In_655,In_359);
nand U2817 (N_2817,In_752,In_661);
nand U2818 (N_2818,In_821,In_130);
or U2819 (N_2819,In_670,In_958);
xor U2820 (N_2820,In_1,In_225);
and U2821 (N_2821,In_712,In_903);
and U2822 (N_2822,In_995,In_35);
nor U2823 (N_2823,In_429,In_443);
nand U2824 (N_2824,In_405,In_962);
and U2825 (N_2825,In_673,In_619);
nor U2826 (N_2826,In_565,In_466);
or U2827 (N_2827,In_233,In_875);
xnor U2828 (N_2828,In_816,In_169);
nor U2829 (N_2829,In_887,In_641);
and U2830 (N_2830,In_923,In_307);
and U2831 (N_2831,In_409,In_801);
and U2832 (N_2832,In_641,In_212);
nor U2833 (N_2833,In_743,In_244);
nand U2834 (N_2834,In_172,In_33);
or U2835 (N_2835,In_166,In_792);
nand U2836 (N_2836,In_789,In_75);
or U2837 (N_2837,In_755,In_923);
and U2838 (N_2838,In_414,In_809);
or U2839 (N_2839,In_672,In_283);
nor U2840 (N_2840,In_494,In_840);
nand U2841 (N_2841,In_852,In_753);
or U2842 (N_2842,In_775,In_590);
or U2843 (N_2843,In_551,In_72);
nand U2844 (N_2844,In_44,In_876);
nand U2845 (N_2845,In_282,In_192);
or U2846 (N_2846,In_989,In_668);
or U2847 (N_2847,In_424,In_272);
and U2848 (N_2848,In_992,In_499);
or U2849 (N_2849,In_449,In_763);
and U2850 (N_2850,In_976,In_936);
xor U2851 (N_2851,In_648,In_800);
and U2852 (N_2852,In_516,In_232);
or U2853 (N_2853,In_180,In_535);
nand U2854 (N_2854,In_525,In_317);
nor U2855 (N_2855,In_162,In_575);
nand U2856 (N_2856,In_749,In_102);
nor U2857 (N_2857,In_849,In_502);
nor U2858 (N_2858,In_619,In_501);
and U2859 (N_2859,In_460,In_671);
and U2860 (N_2860,In_269,In_485);
nor U2861 (N_2861,In_327,In_346);
nor U2862 (N_2862,In_4,In_459);
or U2863 (N_2863,In_203,In_413);
nor U2864 (N_2864,In_914,In_782);
xor U2865 (N_2865,In_510,In_647);
nor U2866 (N_2866,In_438,In_612);
nand U2867 (N_2867,In_18,In_684);
and U2868 (N_2868,In_368,In_182);
and U2869 (N_2869,In_639,In_622);
or U2870 (N_2870,In_879,In_122);
nor U2871 (N_2871,In_209,In_654);
or U2872 (N_2872,In_522,In_648);
nand U2873 (N_2873,In_927,In_693);
or U2874 (N_2874,In_658,In_284);
nand U2875 (N_2875,In_693,In_85);
and U2876 (N_2876,In_681,In_299);
nor U2877 (N_2877,In_566,In_407);
nand U2878 (N_2878,In_125,In_301);
nand U2879 (N_2879,In_63,In_781);
nor U2880 (N_2880,In_937,In_607);
or U2881 (N_2881,In_32,In_704);
or U2882 (N_2882,In_374,In_324);
and U2883 (N_2883,In_272,In_212);
and U2884 (N_2884,In_130,In_124);
and U2885 (N_2885,In_221,In_687);
nand U2886 (N_2886,In_488,In_176);
or U2887 (N_2887,In_791,In_926);
nand U2888 (N_2888,In_46,In_985);
or U2889 (N_2889,In_122,In_521);
or U2890 (N_2890,In_423,In_647);
xnor U2891 (N_2891,In_515,In_969);
and U2892 (N_2892,In_395,In_77);
nor U2893 (N_2893,In_569,In_448);
nand U2894 (N_2894,In_644,In_892);
and U2895 (N_2895,In_37,In_428);
or U2896 (N_2896,In_89,In_841);
or U2897 (N_2897,In_426,In_517);
nor U2898 (N_2898,In_845,In_652);
and U2899 (N_2899,In_107,In_494);
nor U2900 (N_2900,In_431,In_999);
and U2901 (N_2901,In_511,In_700);
nand U2902 (N_2902,In_157,In_824);
nor U2903 (N_2903,In_546,In_12);
and U2904 (N_2904,In_120,In_177);
xnor U2905 (N_2905,In_323,In_217);
nor U2906 (N_2906,In_323,In_648);
nand U2907 (N_2907,In_416,In_244);
nand U2908 (N_2908,In_967,In_863);
nor U2909 (N_2909,In_459,In_71);
nand U2910 (N_2910,In_185,In_148);
nand U2911 (N_2911,In_638,In_536);
or U2912 (N_2912,In_29,In_780);
or U2913 (N_2913,In_447,In_709);
nand U2914 (N_2914,In_710,In_668);
nor U2915 (N_2915,In_232,In_769);
xnor U2916 (N_2916,In_6,In_535);
nand U2917 (N_2917,In_730,In_623);
nand U2918 (N_2918,In_674,In_365);
nor U2919 (N_2919,In_297,In_647);
or U2920 (N_2920,In_603,In_743);
or U2921 (N_2921,In_319,In_849);
nor U2922 (N_2922,In_930,In_143);
or U2923 (N_2923,In_34,In_444);
nand U2924 (N_2924,In_433,In_407);
nor U2925 (N_2925,In_639,In_318);
and U2926 (N_2926,In_745,In_329);
nor U2927 (N_2927,In_7,In_297);
or U2928 (N_2928,In_265,In_690);
or U2929 (N_2929,In_269,In_204);
nand U2930 (N_2930,In_285,In_680);
nand U2931 (N_2931,In_543,In_237);
or U2932 (N_2932,In_947,In_963);
and U2933 (N_2933,In_655,In_764);
xor U2934 (N_2934,In_171,In_531);
nor U2935 (N_2935,In_918,In_520);
nor U2936 (N_2936,In_298,In_85);
nand U2937 (N_2937,In_671,In_667);
and U2938 (N_2938,In_558,In_319);
and U2939 (N_2939,In_69,In_690);
and U2940 (N_2940,In_154,In_632);
nand U2941 (N_2941,In_163,In_752);
nand U2942 (N_2942,In_97,In_660);
or U2943 (N_2943,In_578,In_315);
nand U2944 (N_2944,In_421,In_428);
nand U2945 (N_2945,In_189,In_190);
nand U2946 (N_2946,In_307,In_475);
or U2947 (N_2947,In_394,In_758);
nand U2948 (N_2948,In_470,In_22);
and U2949 (N_2949,In_145,In_415);
and U2950 (N_2950,In_892,In_691);
and U2951 (N_2951,In_795,In_857);
nand U2952 (N_2952,In_225,In_257);
xnor U2953 (N_2953,In_327,In_722);
and U2954 (N_2954,In_251,In_284);
nor U2955 (N_2955,In_561,In_580);
nand U2956 (N_2956,In_761,In_879);
nor U2957 (N_2957,In_953,In_477);
nand U2958 (N_2958,In_481,In_890);
or U2959 (N_2959,In_575,In_152);
and U2960 (N_2960,In_773,In_238);
nor U2961 (N_2961,In_832,In_87);
nand U2962 (N_2962,In_782,In_841);
nor U2963 (N_2963,In_594,In_935);
or U2964 (N_2964,In_637,In_853);
or U2965 (N_2965,In_958,In_423);
or U2966 (N_2966,In_794,In_812);
nand U2967 (N_2967,In_972,In_949);
and U2968 (N_2968,In_680,In_716);
and U2969 (N_2969,In_824,In_195);
nand U2970 (N_2970,In_152,In_788);
xor U2971 (N_2971,In_808,In_494);
nand U2972 (N_2972,In_935,In_375);
nor U2973 (N_2973,In_846,In_387);
nor U2974 (N_2974,In_472,In_547);
and U2975 (N_2975,In_600,In_528);
or U2976 (N_2976,In_36,In_307);
or U2977 (N_2977,In_714,In_589);
nor U2978 (N_2978,In_162,In_772);
or U2979 (N_2979,In_920,In_372);
nand U2980 (N_2980,In_701,In_719);
and U2981 (N_2981,In_493,In_451);
and U2982 (N_2982,In_903,In_379);
nand U2983 (N_2983,In_859,In_700);
nor U2984 (N_2984,In_161,In_774);
or U2985 (N_2985,In_155,In_966);
nor U2986 (N_2986,In_171,In_44);
and U2987 (N_2987,In_811,In_921);
nor U2988 (N_2988,In_339,In_101);
nor U2989 (N_2989,In_721,In_821);
or U2990 (N_2990,In_37,In_388);
nand U2991 (N_2991,In_944,In_605);
and U2992 (N_2992,In_314,In_829);
and U2993 (N_2993,In_4,In_382);
or U2994 (N_2994,In_444,In_145);
nor U2995 (N_2995,In_757,In_390);
or U2996 (N_2996,In_268,In_151);
nor U2997 (N_2997,In_586,In_538);
nor U2998 (N_2998,In_848,In_321);
nand U2999 (N_2999,In_624,In_377);
or U3000 (N_3000,In_789,In_523);
nand U3001 (N_3001,In_304,In_265);
or U3002 (N_3002,In_890,In_794);
and U3003 (N_3003,In_784,In_508);
and U3004 (N_3004,In_554,In_300);
nand U3005 (N_3005,In_45,In_310);
or U3006 (N_3006,In_533,In_573);
nand U3007 (N_3007,In_322,In_785);
nor U3008 (N_3008,In_375,In_126);
and U3009 (N_3009,In_239,In_685);
nor U3010 (N_3010,In_537,In_233);
nor U3011 (N_3011,In_727,In_824);
and U3012 (N_3012,In_666,In_536);
nand U3013 (N_3013,In_335,In_692);
or U3014 (N_3014,In_555,In_527);
xor U3015 (N_3015,In_309,In_715);
or U3016 (N_3016,In_676,In_176);
and U3017 (N_3017,In_424,In_390);
and U3018 (N_3018,In_9,In_127);
nand U3019 (N_3019,In_425,In_86);
nor U3020 (N_3020,In_569,In_468);
or U3021 (N_3021,In_479,In_425);
nand U3022 (N_3022,In_785,In_434);
nand U3023 (N_3023,In_274,In_619);
and U3024 (N_3024,In_596,In_232);
or U3025 (N_3025,In_63,In_644);
and U3026 (N_3026,In_251,In_517);
and U3027 (N_3027,In_73,In_979);
and U3028 (N_3028,In_327,In_398);
nand U3029 (N_3029,In_334,In_733);
nand U3030 (N_3030,In_733,In_546);
nor U3031 (N_3031,In_275,In_514);
nand U3032 (N_3032,In_831,In_185);
and U3033 (N_3033,In_20,In_159);
nand U3034 (N_3034,In_332,In_282);
and U3035 (N_3035,In_564,In_625);
or U3036 (N_3036,In_743,In_16);
and U3037 (N_3037,In_795,In_12);
or U3038 (N_3038,In_648,In_830);
and U3039 (N_3039,In_503,In_587);
nand U3040 (N_3040,In_920,In_918);
nand U3041 (N_3041,In_107,In_244);
nand U3042 (N_3042,In_379,In_894);
nor U3043 (N_3043,In_345,In_943);
and U3044 (N_3044,In_34,In_662);
and U3045 (N_3045,In_821,In_203);
and U3046 (N_3046,In_904,In_19);
nand U3047 (N_3047,In_111,In_905);
and U3048 (N_3048,In_309,In_25);
and U3049 (N_3049,In_713,In_745);
nor U3050 (N_3050,In_712,In_932);
nor U3051 (N_3051,In_387,In_41);
and U3052 (N_3052,In_880,In_376);
or U3053 (N_3053,In_694,In_309);
nor U3054 (N_3054,In_58,In_76);
xor U3055 (N_3055,In_686,In_740);
and U3056 (N_3056,In_568,In_161);
nand U3057 (N_3057,In_335,In_948);
and U3058 (N_3058,In_802,In_742);
nor U3059 (N_3059,In_900,In_528);
and U3060 (N_3060,In_697,In_680);
nor U3061 (N_3061,In_249,In_640);
or U3062 (N_3062,In_43,In_281);
nor U3063 (N_3063,In_468,In_873);
and U3064 (N_3064,In_374,In_878);
nor U3065 (N_3065,In_927,In_543);
nor U3066 (N_3066,In_572,In_997);
nand U3067 (N_3067,In_919,In_65);
nor U3068 (N_3068,In_223,In_918);
and U3069 (N_3069,In_929,In_919);
xor U3070 (N_3070,In_916,In_428);
nand U3071 (N_3071,In_15,In_262);
nand U3072 (N_3072,In_541,In_144);
nand U3073 (N_3073,In_46,In_51);
xor U3074 (N_3074,In_533,In_203);
nand U3075 (N_3075,In_74,In_308);
or U3076 (N_3076,In_369,In_944);
nand U3077 (N_3077,In_693,In_124);
nand U3078 (N_3078,In_903,In_874);
or U3079 (N_3079,In_569,In_383);
or U3080 (N_3080,In_582,In_7);
nor U3081 (N_3081,In_983,In_498);
or U3082 (N_3082,In_5,In_909);
nor U3083 (N_3083,In_134,In_703);
nand U3084 (N_3084,In_643,In_362);
or U3085 (N_3085,In_116,In_636);
nor U3086 (N_3086,In_33,In_735);
and U3087 (N_3087,In_642,In_345);
nand U3088 (N_3088,In_952,In_969);
and U3089 (N_3089,In_409,In_495);
or U3090 (N_3090,In_517,In_246);
nor U3091 (N_3091,In_370,In_689);
nor U3092 (N_3092,In_739,In_275);
nand U3093 (N_3093,In_798,In_951);
or U3094 (N_3094,In_939,In_51);
or U3095 (N_3095,In_915,In_591);
and U3096 (N_3096,In_312,In_71);
nand U3097 (N_3097,In_991,In_388);
nor U3098 (N_3098,In_33,In_525);
or U3099 (N_3099,In_198,In_102);
nand U3100 (N_3100,In_100,In_252);
nand U3101 (N_3101,In_643,In_323);
nor U3102 (N_3102,In_39,In_958);
nor U3103 (N_3103,In_691,In_103);
or U3104 (N_3104,In_730,In_287);
and U3105 (N_3105,In_706,In_356);
nand U3106 (N_3106,In_802,In_235);
nand U3107 (N_3107,In_339,In_462);
and U3108 (N_3108,In_550,In_289);
or U3109 (N_3109,In_33,In_663);
and U3110 (N_3110,In_739,In_508);
or U3111 (N_3111,In_144,In_298);
nand U3112 (N_3112,In_790,In_546);
nor U3113 (N_3113,In_610,In_75);
or U3114 (N_3114,In_320,In_198);
or U3115 (N_3115,In_760,In_42);
and U3116 (N_3116,In_334,In_361);
or U3117 (N_3117,In_685,In_415);
nand U3118 (N_3118,In_687,In_995);
nand U3119 (N_3119,In_668,In_143);
nor U3120 (N_3120,In_490,In_359);
nand U3121 (N_3121,In_862,In_382);
or U3122 (N_3122,In_908,In_951);
or U3123 (N_3123,In_552,In_103);
nand U3124 (N_3124,In_531,In_827);
and U3125 (N_3125,In_222,In_700);
or U3126 (N_3126,In_935,In_475);
nand U3127 (N_3127,In_765,In_931);
nand U3128 (N_3128,In_217,In_138);
nor U3129 (N_3129,In_797,In_725);
nand U3130 (N_3130,In_412,In_62);
nand U3131 (N_3131,In_189,In_100);
nand U3132 (N_3132,In_803,In_398);
xor U3133 (N_3133,In_559,In_189);
and U3134 (N_3134,In_812,In_39);
and U3135 (N_3135,In_628,In_796);
nor U3136 (N_3136,In_505,In_308);
nand U3137 (N_3137,In_406,In_954);
nor U3138 (N_3138,In_944,In_273);
or U3139 (N_3139,In_458,In_150);
nor U3140 (N_3140,In_872,In_783);
or U3141 (N_3141,In_30,In_358);
nor U3142 (N_3142,In_496,In_490);
and U3143 (N_3143,In_611,In_406);
nor U3144 (N_3144,In_760,In_459);
or U3145 (N_3145,In_18,In_759);
and U3146 (N_3146,In_978,In_325);
nand U3147 (N_3147,In_67,In_670);
nand U3148 (N_3148,In_296,In_922);
nor U3149 (N_3149,In_949,In_292);
and U3150 (N_3150,In_75,In_543);
nand U3151 (N_3151,In_592,In_277);
xnor U3152 (N_3152,In_209,In_457);
nor U3153 (N_3153,In_506,In_593);
nand U3154 (N_3154,In_897,In_689);
or U3155 (N_3155,In_947,In_680);
and U3156 (N_3156,In_89,In_347);
nor U3157 (N_3157,In_777,In_53);
nand U3158 (N_3158,In_235,In_310);
nor U3159 (N_3159,In_824,In_337);
and U3160 (N_3160,In_480,In_989);
and U3161 (N_3161,In_475,In_245);
and U3162 (N_3162,In_743,In_872);
nand U3163 (N_3163,In_661,In_225);
or U3164 (N_3164,In_991,In_609);
nor U3165 (N_3165,In_988,In_791);
and U3166 (N_3166,In_79,In_247);
nand U3167 (N_3167,In_828,In_546);
or U3168 (N_3168,In_837,In_446);
and U3169 (N_3169,In_351,In_424);
or U3170 (N_3170,In_206,In_716);
or U3171 (N_3171,In_726,In_309);
or U3172 (N_3172,In_283,In_745);
nand U3173 (N_3173,In_95,In_198);
nor U3174 (N_3174,In_60,In_486);
nor U3175 (N_3175,In_179,In_501);
and U3176 (N_3176,In_168,In_629);
nand U3177 (N_3177,In_101,In_738);
nand U3178 (N_3178,In_508,In_232);
or U3179 (N_3179,In_75,In_148);
and U3180 (N_3180,In_148,In_563);
nand U3181 (N_3181,In_568,In_457);
or U3182 (N_3182,In_37,In_189);
and U3183 (N_3183,In_744,In_5);
nor U3184 (N_3184,In_118,In_498);
nand U3185 (N_3185,In_482,In_281);
nor U3186 (N_3186,In_2,In_204);
or U3187 (N_3187,In_77,In_587);
or U3188 (N_3188,In_425,In_843);
or U3189 (N_3189,In_573,In_208);
and U3190 (N_3190,In_817,In_898);
or U3191 (N_3191,In_699,In_766);
and U3192 (N_3192,In_541,In_16);
or U3193 (N_3193,In_106,In_550);
or U3194 (N_3194,In_43,In_708);
nand U3195 (N_3195,In_579,In_858);
or U3196 (N_3196,In_186,In_753);
and U3197 (N_3197,In_941,In_273);
nor U3198 (N_3198,In_692,In_998);
nand U3199 (N_3199,In_539,In_17);
and U3200 (N_3200,In_992,In_441);
or U3201 (N_3201,In_246,In_715);
nor U3202 (N_3202,In_745,In_170);
nand U3203 (N_3203,In_707,In_45);
nor U3204 (N_3204,In_135,In_883);
or U3205 (N_3205,In_464,In_894);
nor U3206 (N_3206,In_268,In_4);
nor U3207 (N_3207,In_904,In_138);
nand U3208 (N_3208,In_834,In_998);
and U3209 (N_3209,In_705,In_44);
nand U3210 (N_3210,In_795,In_44);
and U3211 (N_3211,In_919,In_601);
and U3212 (N_3212,In_871,In_760);
nor U3213 (N_3213,In_981,In_164);
nor U3214 (N_3214,In_650,In_670);
nor U3215 (N_3215,In_747,In_316);
and U3216 (N_3216,In_247,In_170);
or U3217 (N_3217,In_858,In_234);
and U3218 (N_3218,In_221,In_954);
or U3219 (N_3219,In_893,In_882);
or U3220 (N_3220,In_39,In_387);
and U3221 (N_3221,In_581,In_882);
nand U3222 (N_3222,In_466,In_728);
nor U3223 (N_3223,In_666,In_318);
or U3224 (N_3224,In_730,In_884);
or U3225 (N_3225,In_230,In_432);
nor U3226 (N_3226,In_839,In_690);
or U3227 (N_3227,In_245,In_64);
or U3228 (N_3228,In_736,In_279);
nand U3229 (N_3229,In_426,In_611);
and U3230 (N_3230,In_808,In_80);
nor U3231 (N_3231,In_199,In_510);
nand U3232 (N_3232,In_235,In_429);
or U3233 (N_3233,In_485,In_417);
xnor U3234 (N_3234,In_328,In_913);
nand U3235 (N_3235,In_657,In_546);
or U3236 (N_3236,In_349,In_23);
or U3237 (N_3237,In_885,In_197);
nor U3238 (N_3238,In_147,In_924);
nor U3239 (N_3239,In_855,In_568);
or U3240 (N_3240,In_989,In_35);
and U3241 (N_3241,In_887,In_976);
nor U3242 (N_3242,In_985,In_801);
or U3243 (N_3243,In_994,In_135);
nand U3244 (N_3244,In_170,In_634);
or U3245 (N_3245,In_642,In_951);
and U3246 (N_3246,In_974,In_40);
nor U3247 (N_3247,In_35,In_14);
nand U3248 (N_3248,In_799,In_523);
nand U3249 (N_3249,In_416,In_753);
and U3250 (N_3250,In_518,In_735);
nand U3251 (N_3251,In_242,In_944);
or U3252 (N_3252,In_172,In_904);
and U3253 (N_3253,In_979,In_447);
and U3254 (N_3254,In_767,In_835);
xor U3255 (N_3255,In_533,In_951);
or U3256 (N_3256,In_911,In_641);
xor U3257 (N_3257,In_704,In_658);
or U3258 (N_3258,In_632,In_273);
nor U3259 (N_3259,In_73,In_733);
and U3260 (N_3260,In_531,In_307);
or U3261 (N_3261,In_618,In_892);
xor U3262 (N_3262,In_363,In_350);
nor U3263 (N_3263,In_834,In_127);
and U3264 (N_3264,In_823,In_57);
and U3265 (N_3265,In_428,In_807);
nand U3266 (N_3266,In_238,In_850);
or U3267 (N_3267,In_422,In_618);
nor U3268 (N_3268,In_623,In_702);
or U3269 (N_3269,In_111,In_509);
or U3270 (N_3270,In_844,In_78);
or U3271 (N_3271,In_500,In_976);
and U3272 (N_3272,In_957,In_643);
nand U3273 (N_3273,In_239,In_64);
or U3274 (N_3274,In_798,In_683);
and U3275 (N_3275,In_222,In_281);
or U3276 (N_3276,In_818,In_441);
and U3277 (N_3277,In_411,In_166);
nor U3278 (N_3278,In_721,In_524);
and U3279 (N_3279,In_686,In_684);
or U3280 (N_3280,In_679,In_715);
and U3281 (N_3281,In_96,In_719);
nand U3282 (N_3282,In_441,In_632);
nand U3283 (N_3283,In_561,In_639);
nor U3284 (N_3284,In_790,In_79);
or U3285 (N_3285,In_542,In_706);
and U3286 (N_3286,In_592,In_141);
and U3287 (N_3287,In_94,In_694);
xor U3288 (N_3288,In_941,In_200);
nand U3289 (N_3289,In_410,In_310);
and U3290 (N_3290,In_851,In_540);
nor U3291 (N_3291,In_755,In_970);
nand U3292 (N_3292,In_714,In_509);
nand U3293 (N_3293,In_388,In_134);
nor U3294 (N_3294,In_730,In_782);
nand U3295 (N_3295,In_666,In_592);
and U3296 (N_3296,In_788,In_22);
or U3297 (N_3297,In_765,In_70);
or U3298 (N_3298,In_591,In_227);
and U3299 (N_3299,In_350,In_374);
or U3300 (N_3300,In_784,In_494);
nor U3301 (N_3301,In_493,In_686);
nand U3302 (N_3302,In_449,In_208);
nor U3303 (N_3303,In_338,In_408);
xor U3304 (N_3304,In_303,In_793);
or U3305 (N_3305,In_381,In_474);
and U3306 (N_3306,In_796,In_352);
nor U3307 (N_3307,In_201,In_601);
and U3308 (N_3308,In_305,In_714);
or U3309 (N_3309,In_44,In_541);
nand U3310 (N_3310,In_944,In_666);
nor U3311 (N_3311,In_821,In_499);
or U3312 (N_3312,In_502,In_233);
nand U3313 (N_3313,In_469,In_359);
nor U3314 (N_3314,In_825,In_158);
and U3315 (N_3315,In_687,In_47);
xor U3316 (N_3316,In_862,In_969);
and U3317 (N_3317,In_634,In_433);
nand U3318 (N_3318,In_858,In_860);
xnor U3319 (N_3319,In_60,In_67);
nand U3320 (N_3320,In_659,In_698);
or U3321 (N_3321,In_484,In_288);
nand U3322 (N_3322,In_886,In_845);
nor U3323 (N_3323,In_470,In_620);
or U3324 (N_3324,In_327,In_651);
and U3325 (N_3325,In_42,In_306);
or U3326 (N_3326,In_927,In_345);
or U3327 (N_3327,In_426,In_30);
nand U3328 (N_3328,In_32,In_822);
or U3329 (N_3329,In_102,In_617);
and U3330 (N_3330,In_482,In_835);
nand U3331 (N_3331,In_14,In_352);
nor U3332 (N_3332,In_653,In_377);
nand U3333 (N_3333,In_739,In_183);
nor U3334 (N_3334,In_942,In_313);
nor U3335 (N_3335,In_448,In_159);
nand U3336 (N_3336,In_992,In_849);
nand U3337 (N_3337,In_540,In_703);
nand U3338 (N_3338,In_152,In_740);
and U3339 (N_3339,In_576,In_368);
or U3340 (N_3340,In_978,In_630);
nor U3341 (N_3341,In_495,In_197);
or U3342 (N_3342,In_681,In_643);
or U3343 (N_3343,In_288,In_374);
or U3344 (N_3344,In_667,In_573);
nand U3345 (N_3345,In_278,In_103);
or U3346 (N_3346,In_394,In_478);
nand U3347 (N_3347,In_773,In_444);
and U3348 (N_3348,In_982,In_470);
nor U3349 (N_3349,In_375,In_841);
xnor U3350 (N_3350,In_362,In_64);
and U3351 (N_3351,In_127,In_495);
or U3352 (N_3352,In_232,In_471);
nor U3353 (N_3353,In_820,In_271);
or U3354 (N_3354,In_876,In_858);
or U3355 (N_3355,In_173,In_332);
nand U3356 (N_3356,In_195,In_80);
nand U3357 (N_3357,In_665,In_960);
and U3358 (N_3358,In_611,In_702);
or U3359 (N_3359,In_696,In_772);
nor U3360 (N_3360,In_518,In_538);
or U3361 (N_3361,In_165,In_526);
nand U3362 (N_3362,In_964,In_954);
or U3363 (N_3363,In_891,In_766);
nand U3364 (N_3364,In_311,In_899);
and U3365 (N_3365,In_491,In_532);
or U3366 (N_3366,In_558,In_187);
nor U3367 (N_3367,In_440,In_245);
and U3368 (N_3368,In_276,In_437);
or U3369 (N_3369,In_412,In_120);
or U3370 (N_3370,In_386,In_27);
nand U3371 (N_3371,In_429,In_762);
and U3372 (N_3372,In_45,In_376);
nand U3373 (N_3373,In_937,In_983);
nand U3374 (N_3374,In_191,In_917);
and U3375 (N_3375,In_924,In_704);
or U3376 (N_3376,In_889,In_284);
nand U3377 (N_3377,In_570,In_105);
nor U3378 (N_3378,In_308,In_267);
and U3379 (N_3379,In_152,In_579);
or U3380 (N_3380,In_988,In_196);
and U3381 (N_3381,In_635,In_776);
or U3382 (N_3382,In_117,In_274);
and U3383 (N_3383,In_701,In_936);
nand U3384 (N_3384,In_529,In_2);
nor U3385 (N_3385,In_193,In_970);
and U3386 (N_3386,In_183,In_652);
and U3387 (N_3387,In_44,In_990);
and U3388 (N_3388,In_709,In_116);
or U3389 (N_3389,In_252,In_241);
nand U3390 (N_3390,In_515,In_866);
nand U3391 (N_3391,In_680,In_198);
and U3392 (N_3392,In_903,In_592);
nor U3393 (N_3393,In_525,In_51);
or U3394 (N_3394,In_791,In_874);
nand U3395 (N_3395,In_819,In_414);
or U3396 (N_3396,In_462,In_291);
nand U3397 (N_3397,In_220,In_6);
nand U3398 (N_3398,In_344,In_200);
nand U3399 (N_3399,In_201,In_466);
or U3400 (N_3400,In_807,In_743);
nor U3401 (N_3401,In_766,In_34);
and U3402 (N_3402,In_465,In_132);
nor U3403 (N_3403,In_707,In_362);
nand U3404 (N_3404,In_250,In_100);
or U3405 (N_3405,In_969,In_263);
nor U3406 (N_3406,In_123,In_97);
nor U3407 (N_3407,In_235,In_30);
xor U3408 (N_3408,In_409,In_416);
xor U3409 (N_3409,In_28,In_318);
and U3410 (N_3410,In_140,In_57);
nor U3411 (N_3411,In_953,In_841);
and U3412 (N_3412,In_839,In_726);
nand U3413 (N_3413,In_893,In_892);
or U3414 (N_3414,In_299,In_312);
or U3415 (N_3415,In_962,In_449);
or U3416 (N_3416,In_783,In_486);
nand U3417 (N_3417,In_52,In_684);
and U3418 (N_3418,In_220,In_760);
nor U3419 (N_3419,In_778,In_73);
or U3420 (N_3420,In_611,In_180);
nor U3421 (N_3421,In_90,In_521);
xor U3422 (N_3422,In_311,In_528);
and U3423 (N_3423,In_378,In_896);
nor U3424 (N_3424,In_4,In_213);
or U3425 (N_3425,In_8,In_121);
nor U3426 (N_3426,In_625,In_492);
or U3427 (N_3427,In_79,In_118);
nor U3428 (N_3428,In_73,In_252);
and U3429 (N_3429,In_448,In_411);
nor U3430 (N_3430,In_94,In_366);
nand U3431 (N_3431,In_287,In_138);
nor U3432 (N_3432,In_475,In_149);
nand U3433 (N_3433,In_699,In_407);
and U3434 (N_3434,In_965,In_930);
and U3435 (N_3435,In_782,In_467);
or U3436 (N_3436,In_95,In_998);
nand U3437 (N_3437,In_119,In_461);
and U3438 (N_3438,In_360,In_644);
and U3439 (N_3439,In_811,In_23);
or U3440 (N_3440,In_753,In_548);
nand U3441 (N_3441,In_360,In_635);
or U3442 (N_3442,In_788,In_127);
and U3443 (N_3443,In_705,In_513);
nor U3444 (N_3444,In_576,In_147);
and U3445 (N_3445,In_602,In_899);
nor U3446 (N_3446,In_976,In_834);
or U3447 (N_3447,In_433,In_184);
or U3448 (N_3448,In_145,In_216);
or U3449 (N_3449,In_683,In_795);
nand U3450 (N_3450,In_592,In_268);
or U3451 (N_3451,In_979,In_490);
and U3452 (N_3452,In_965,In_791);
or U3453 (N_3453,In_283,In_81);
nor U3454 (N_3454,In_664,In_885);
and U3455 (N_3455,In_775,In_302);
nand U3456 (N_3456,In_378,In_594);
nor U3457 (N_3457,In_420,In_11);
nand U3458 (N_3458,In_446,In_707);
or U3459 (N_3459,In_322,In_871);
nand U3460 (N_3460,In_865,In_63);
nor U3461 (N_3461,In_913,In_183);
nand U3462 (N_3462,In_377,In_726);
or U3463 (N_3463,In_874,In_302);
nor U3464 (N_3464,In_85,In_376);
nor U3465 (N_3465,In_529,In_787);
or U3466 (N_3466,In_176,In_960);
nand U3467 (N_3467,In_650,In_195);
or U3468 (N_3468,In_920,In_50);
nor U3469 (N_3469,In_180,In_502);
or U3470 (N_3470,In_995,In_629);
and U3471 (N_3471,In_791,In_623);
nand U3472 (N_3472,In_982,In_398);
nor U3473 (N_3473,In_162,In_129);
nor U3474 (N_3474,In_391,In_89);
nand U3475 (N_3475,In_429,In_694);
and U3476 (N_3476,In_973,In_914);
and U3477 (N_3477,In_142,In_945);
or U3478 (N_3478,In_96,In_674);
nor U3479 (N_3479,In_322,In_981);
or U3480 (N_3480,In_613,In_374);
nand U3481 (N_3481,In_582,In_374);
nor U3482 (N_3482,In_602,In_606);
nor U3483 (N_3483,In_942,In_10);
nor U3484 (N_3484,In_331,In_898);
nor U3485 (N_3485,In_315,In_322);
nor U3486 (N_3486,In_966,In_639);
nand U3487 (N_3487,In_284,In_461);
nand U3488 (N_3488,In_364,In_954);
nor U3489 (N_3489,In_372,In_753);
nor U3490 (N_3490,In_59,In_739);
nor U3491 (N_3491,In_3,In_594);
or U3492 (N_3492,In_84,In_800);
and U3493 (N_3493,In_795,In_422);
or U3494 (N_3494,In_324,In_286);
nor U3495 (N_3495,In_882,In_937);
or U3496 (N_3496,In_35,In_588);
xnor U3497 (N_3497,In_230,In_730);
nor U3498 (N_3498,In_9,In_778);
nand U3499 (N_3499,In_519,In_381);
or U3500 (N_3500,In_912,In_24);
nor U3501 (N_3501,In_416,In_529);
nand U3502 (N_3502,In_57,In_102);
nand U3503 (N_3503,In_115,In_159);
nor U3504 (N_3504,In_927,In_465);
and U3505 (N_3505,In_378,In_13);
nand U3506 (N_3506,In_322,In_77);
or U3507 (N_3507,In_638,In_738);
and U3508 (N_3508,In_147,In_11);
and U3509 (N_3509,In_859,In_905);
nand U3510 (N_3510,In_585,In_363);
or U3511 (N_3511,In_495,In_684);
nand U3512 (N_3512,In_235,In_489);
nor U3513 (N_3513,In_239,In_65);
nand U3514 (N_3514,In_31,In_613);
or U3515 (N_3515,In_552,In_344);
or U3516 (N_3516,In_593,In_325);
and U3517 (N_3517,In_450,In_879);
nand U3518 (N_3518,In_574,In_494);
nand U3519 (N_3519,In_194,In_392);
nor U3520 (N_3520,In_554,In_636);
and U3521 (N_3521,In_946,In_581);
or U3522 (N_3522,In_282,In_413);
and U3523 (N_3523,In_636,In_92);
nor U3524 (N_3524,In_277,In_596);
or U3525 (N_3525,In_69,In_856);
nor U3526 (N_3526,In_742,In_292);
nor U3527 (N_3527,In_517,In_532);
or U3528 (N_3528,In_784,In_987);
nor U3529 (N_3529,In_248,In_256);
nor U3530 (N_3530,In_527,In_956);
or U3531 (N_3531,In_644,In_992);
and U3532 (N_3532,In_738,In_923);
and U3533 (N_3533,In_59,In_321);
nor U3534 (N_3534,In_560,In_618);
nand U3535 (N_3535,In_153,In_31);
nand U3536 (N_3536,In_197,In_255);
and U3537 (N_3537,In_877,In_54);
xnor U3538 (N_3538,In_825,In_333);
nand U3539 (N_3539,In_977,In_465);
and U3540 (N_3540,In_825,In_563);
and U3541 (N_3541,In_326,In_543);
or U3542 (N_3542,In_897,In_681);
nand U3543 (N_3543,In_498,In_907);
or U3544 (N_3544,In_28,In_306);
or U3545 (N_3545,In_281,In_956);
nor U3546 (N_3546,In_168,In_607);
or U3547 (N_3547,In_907,In_104);
xor U3548 (N_3548,In_595,In_147);
nor U3549 (N_3549,In_422,In_532);
nand U3550 (N_3550,In_986,In_830);
nor U3551 (N_3551,In_105,In_271);
and U3552 (N_3552,In_938,In_314);
or U3553 (N_3553,In_615,In_960);
or U3554 (N_3554,In_179,In_836);
nor U3555 (N_3555,In_940,In_803);
nor U3556 (N_3556,In_169,In_223);
or U3557 (N_3557,In_994,In_126);
or U3558 (N_3558,In_7,In_613);
or U3559 (N_3559,In_602,In_297);
or U3560 (N_3560,In_61,In_116);
and U3561 (N_3561,In_422,In_500);
and U3562 (N_3562,In_34,In_896);
or U3563 (N_3563,In_270,In_856);
nor U3564 (N_3564,In_23,In_305);
and U3565 (N_3565,In_405,In_539);
nand U3566 (N_3566,In_343,In_200);
and U3567 (N_3567,In_647,In_140);
nand U3568 (N_3568,In_321,In_923);
xor U3569 (N_3569,In_252,In_471);
nor U3570 (N_3570,In_46,In_53);
and U3571 (N_3571,In_602,In_675);
nor U3572 (N_3572,In_900,In_227);
nand U3573 (N_3573,In_914,In_436);
or U3574 (N_3574,In_201,In_772);
nor U3575 (N_3575,In_337,In_997);
nand U3576 (N_3576,In_950,In_934);
nand U3577 (N_3577,In_775,In_987);
xnor U3578 (N_3578,In_377,In_313);
nor U3579 (N_3579,In_930,In_624);
and U3580 (N_3580,In_886,In_131);
nor U3581 (N_3581,In_864,In_424);
and U3582 (N_3582,In_517,In_708);
nor U3583 (N_3583,In_318,In_124);
or U3584 (N_3584,In_712,In_665);
nand U3585 (N_3585,In_621,In_413);
nor U3586 (N_3586,In_425,In_200);
nand U3587 (N_3587,In_360,In_467);
nand U3588 (N_3588,In_664,In_112);
and U3589 (N_3589,In_979,In_503);
and U3590 (N_3590,In_507,In_396);
and U3591 (N_3591,In_135,In_715);
or U3592 (N_3592,In_331,In_633);
and U3593 (N_3593,In_412,In_204);
or U3594 (N_3594,In_234,In_309);
and U3595 (N_3595,In_361,In_22);
nand U3596 (N_3596,In_738,In_876);
and U3597 (N_3597,In_557,In_707);
or U3598 (N_3598,In_634,In_774);
or U3599 (N_3599,In_796,In_417);
and U3600 (N_3600,In_148,In_38);
nor U3601 (N_3601,In_510,In_153);
and U3602 (N_3602,In_6,In_62);
nor U3603 (N_3603,In_951,In_690);
nand U3604 (N_3604,In_534,In_303);
or U3605 (N_3605,In_513,In_231);
or U3606 (N_3606,In_440,In_740);
or U3607 (N_3607,In_604,In_731);
or U3608 (N_3608,In_900,In_949);
and U3609 (N_3609,In_920,In_230);
and U3610 (N_3610,In_114,In_160);
nor U3611 (N_3611,In_221,In_558);
nor U3612 (N_3612,In_108,In_186);
or U3613 (N_3613,In_593,In_903);
or U3614 (N_3614,In_91,In_560);
nor U3615 (N_3615,In_373,In_892);
or U3616 (N_3616,In_973,In_30);
nor U3617 (N_3617,In_161,In_354);
nand U3618 (N_3618,In_95,In_363);
nor U3619 (N_3619,In_78,In_145);
and U3620 (N_3620,In_779,In_148);
and U3621 (N_3621,In_154,In_124);
nor U3622 (N_3622,In_61,In_848);
nor U3623 (N_3623,In_504,In_647);
nor U3624 (N_3624,In_636,In_879);
nand U3625 (N_3625,In_612,In_361);
or U3626 (N_3626,In_23,In_460);
and U3627 (N_3627,In_991,In_723);
or U3628 (N_3628,In_225,In_342);
or U3629 (N_3629,In_14,In_283);
and U3630 (N_3630,In_637,In_486);
nor U3631 (N_3631,In_989,In_852);
and U3632 (N_3632,In_308,In_737);
nand U3633 (N_3633,In_382,In_299);
xor U3634 (N_3634,In_825,In_933);
and U3635 (N_3635,In_174,In_367);
nand U3636 (N_3636,In_40,In_553);
nand U3637 (N_3637,In_571,In_964);
and U3638 (N_3638,In_208,In_683);
or U3639 (N_3639,In_157,In_421);
and U3640 (N_3640,In_577,In_107);
nand U3641 (N_3641,In_318,In_500);
or U3642 (N_3642,In_562,In_618);
and U3643 (N_3643,In_74,In_479);
or U3644 (N_3644,In_499,In_17);
xor U3645 (N_3645,In_540,In_50);
nand U3646 (N_3646,In_753,In_731);
nor U3647 (N_3647,In_940,In_217);
or U3648 (N_3648,In_130,In_776);
xor U3649 (N_3649,In_126,In_528);
nand U3650 (N_3650,In_451,In_488);
and U3651 (N_3651,In_807,In_900);
or U3652 (N_3652,In_964,In_191);
or U3653 (N_3653,In_428,In_274);
and U3654 (N_3654,In_645,In_103);
or U3655 (N_3655,In_352,In_272);
nand U3656 (N_3656,In_857,In_434);
or U3657 (N_3657,In_670,In_852);
nor U3658 (N_3658,In_335,In_148);
nand U3659 (N_3659,In_895,In_125);
and U3660 (N_3660,In_847,In_134);
or U3661 (N_3661,In_623,In_29);
nand U3662 (N_3662,In_800,In_968);
and U3663 (N_3663,In_614,In_779);
and U3664 (N_3664,In_341,In_811);
nor U3665 (N_3665,In_794,In_191);
or U3666 (N_3666,In_890,In_588);
and U3667 (N_3667,In_22,In_832);
xor U3668 (N_3668,In_839,In_306);
xnor U3669 (N_3669,In_156,In_683);
nor U3670 (N_3670,In_379,In_272);
and U3671 (N_3671,In_906,In_406);
and U3672 (N_3672,In_34,In_451);
or U3673 (N_3673,In_81,In_362);
nand U3674 (N_3674,In_847,In_155);
nor U3675 (N_3675,In_7,In_623);
or U3676 (N_3676,In_228,In_243);
nor U3677 (N_3677,In_397,In_757);
and U3678 (N_3678,In_199,In_668);
nand U3679 (N_3679,In_584,In_903);
and U3680 (N_3680,In_573,In_688);
and U3681 (N_3681,In_62,In_19);
nor U3682 (N_3682,In_538,In_310);
nor U3683 (N_3683,In_870,In_368);
nand U3684 (N_3684,In_560,In_753);
nand U3685 (N_3685,In_935,In_244);
and U3686 (N_3686,In_427,In_821);
and U3687 (N_3687,In_428,In_494);
nand U3688 (N_3688,In_136,In_593);
or U3689 (N_3689,In_679,In_34);
nor U3690 (N_3690,In_289,In_780);
and U3691 (N_3691,In_502,In_776);
and U3692 (N_3692,In_212,In_483);
nand U3693 (N_3693,In_962,In_757);
nand U3694 (N_3694,In_508,In_969);
or U3695 (N_3695,In_262,In_161);
or U3696 (N_3696,In_468,In_417);
and U3697 (N_3697,In_618,In_324);
nand U3698 (N_3698,In_75,In_971);
and U3699 (N_3699,In_948,In_633);
or U3700 (N_3700,In_915,In_174);
nor U3701 (N_3701,In_640,In_374);
nor U3702 (N_3702,In_49,In_731);
nor U3703 (N_3703,In_858,In_3);
and U3704 (N_3704,In_408,In_984);
or U3705 (N_3705,In_245,In_695);
or U3706 (N_3706,In_164,In_770);
or U3707 (N_3707,In_378,In_524);
nor U3708 (N_3708,In_834,In_896);
nand U3709 (N_3709,In_406,In_286);
nor U3710 (N_3710,In_73,In_678);
nor U3711 (N_3711,In_876,In_312);
or U3712 (N_3712,In_764,In_337);
and U3713 (N_3713,In_698,In_694);
nor U3714 (N_3714,In_744,In_863);
xor U3715 (N_3715,In_490,In_660);
nand U3716 (N_3716,In_880,In_948);
nand U3717 (N_3717,In_911,In_421);
nor U3718 (N_3718,In_684,In_999);
or U3719 (N_3719,In_776,In_927);
nor U3720 (N_3720,In_692,In_569);
or U3721 (N_3721,In_546,In_331);
and U3722 (N_3722,In_721,In_439);
or U3723 (N_3723,In_789,In_136);
nor U3724 (N_3724,In_20,In_456);
or U3725 (N_3725,In_695,In_349);
nand U3726 (N_3726,In_392,In_43);
nor U3727 (N_3727,In_359,In_505);
xor U3728 (N_3728,In_116,In_180);
and U3729 (N_3729,In_122,In_656);
and U3730 (N_3730,In_736,In_391);
and U3731 (N_3731,In_604,In_417);
or U3732 (N_3732,In_710,In_988);
and U3733 (N_3733,In_121,In_493);
nor U3734 (N_3734,In_656,In_662);
nor U3735 (N_3735,In_399,In_560);
nand U3736 (N_3736,In_946,In_3);
nor U3737 (N_3737,In_330,In_797);
nand U3738 (N_3738,In_498,In_159);
and U3739 (N_3739,In_695,In_626);
and U3740 (N_3740,In_846,In_208);
nand U3741 (N_3741,In_924,In_618);
nand U3742 (N_3742,In_429,In_551);
nand U3743 (N_3743,In_302,In_30);
nand U3744 (N_3744,In_675,In_727);
or U3745 (N_3745,In_520,In_719);
and U3746 (N_3746,In_87,In_577);
and U3747 (N_3747,In_551,In_306);
and U3748 (N_3748,In_536,In_240);
and U3749 (N_3749,In_319,In_697);
nor U3750 (N_3750,In_816,In_686);
and U3751 (N_3751,In_116,In_487);
and U3752 (N_3752,In_649,In_106);
or U3753 (N_3753,In_314,In_575);
and U3754 (N_3754,In_19,In_432);
nor U3755 (N_3755,In_44,In_552);
or U3756 (N_3756,In_334,In_594);
nor U3757 (N_3757,In_809,In_834);
or U3758 (N_3758,In_440,In_42);
nand U3759 (N_3759,In_682,In_9);
nor U3760 (N_3760,In_490,In_420);
and U3761 (N_3761,In_770,In_143);
nand U3762 (N_3762,In_727,In_454);
nor U3763 (N_3763,In_381,In_335);
nand U3764 (N_3764,In_838,In_315);
xnor U3765 (N_3765,In_734,In_970);
and U3766 (N_3766,In_154,In_694);
nand U3767 (N_3767,In_118,In_878);
or U3768 (N_3768,In_49,In_537);
nor U3769 (N_3769,In_127,In_854);
and U3770 (N_3770,In_723,In_746);
nor U3771 (N_3771,In_384,In_339);
nor U3772 (N_3772,In_301,In_503);
nor U3773 (N_3773,In_164,In_379);
and U3774 (N_3774,In_268,In_38);
and U3775 (N_3775,In_545,In_174);
nand U3776 (N_3776,In_904,In_388);
or U3777 (N_3777,In_563,In_518);
nand U3778 (N_3778,In_649,In_979);
or U3779 (N_3779,In_496,In_466);
nor U3780 (N_3780,In_542,In_710);
nand U3781 (N_3781,In_33,In_404);
or U3782 (N_3782,In_605,In_544);
nor U3783 (N_3783,In_405,In_532);
and U3784 (N_3784,In_310,In_67);
and U3785 (N_3785,In_926,In_565);
nand U3786 (N_3786,In_441,In_913);
and U3787 (N_3787,In_412,In_517);
and U3788 (N_3788,In_62,In_665);
nor U3789 (N_3789,In_887,In_415);
nor U3790 (N_3790,In_55,In_140);
nor U3791 (N_3791,In_997,In_522);
xor U3792 (N_3792,In_515,In_41);
nor U3793 (N_3793,In_878,In_779);
nor U3794 (N_3794,In_291,In_386);
nor U3795 (N_3795,In_573,In_559);
and U3796 (N_3796,In_687,In_466);
nand U3797 (N_3797,In_322,In_649);
nor U3798 (N_3798,In_246,In_189);
nor U3799 (N_3799,In_947,In_779);
xnor U3800 (N_3800,In_198,In_928);
nand U3801 (N_3801,In_79,In_545);
or U3802 (N_3802,In_572,In_36);
and U3803 (N_3803,In_975,In_850);
nor U3804 (N_3804,In_31,In_315);
nor U3805 (N_3805,In_443,In_10);
nand U3806 (N_3806,In_943,In_315);
or U3807 (N_3807,In_920,In_597);
nor U3808 (N_3808,In_243,In_550);
nand U3809 (N_3809,In_546,In_94);
and U3810 (N_3810,In_338,In_681);
nand U3811 (N_3811,In_758,In_11);
or U3812 (N_3812,In_741,In_344);
or U3813 (N_3813,In_827,In_371);
and U3814 (N_3814,In_90,In_541);
nor U3815 (N_3815,In_457,In_936);
or U3816 (N_3816,In_155,In_19);
or U3817 (N_3817,In_857,In_724);
or U3818 (N_3818,In_719,In_995);
nand U3819 (N_3819,In_548,In_861);
or U3820 (N_3820,In_21,In_300);
nor U3821 (N_3821,In_699,In_710);
and U3822 (N_3822,In_966,In_637);
and U3823 (N_3823,In_634,In_571);
and U3824 (N_3824,In_899,In_815);
nand U3825 (N_3825,In_406,In_654);
or U3826 (N_3826,In_183,In_283);
or U3827 (N_3827,In_260,In_975);
and U3828 (N_3828,In_544,In_51);
nor U3829 (N_3829,In_421,In_91);
and U3830 (N_3830,In_899,In_30);
or U3831 (N_3831,In_822,In_984);
or U3832 (N_3832,In_716,In_749);
nor U3833 (N_3833,In_546,In_236);
nor U3834 (N_3834,In_109,In_106);
and U3835 (N_3835,In_346,In_369);
nor U3836 (N_3836,In_588,In_296);
nor U3837 (N_3837,In_140,In_158);
or U3838 (N_3838,In_163,In_862);
xor U3839 (N_3839,In_487,In_7);
and U3840 (N_3840,In_476,In_55);
or U3841 (N_3841,In_746,In_989);
and U3842 (N_3842,In_751,In_51);
nor U3843 (N_3843,In_939,In_778);
nor U3844 (N_3844,In_52,In_665);
or U3845 (N_3845,In_521,In_43);
nand U3846 (N_3846,In_571,In_632);
and U3847 (N_3847,In_743,In_980);
nand U3848 (N_3848,In_885,In_673);
or U3849 (N_3849,In_363,In_464);
or U3850 (N_3850,In_593,In_382);
and U3851 (N_3851,In_428,In_803);
xor U3852 (N_3852,In_980,In_245);
nor U3853 (N_3853,In_569,In_983);
xor U3854 (N_3854,In_494,In_635);
nor U3855 (N_3855,In_311,In_417);
or U3856 (N_3856,In_363,In_918);
nand U3857 (N_3857,In_668,In_332);
or U3858 (N_3858,In_472,In_517);
or U3859 (N_3859,In_469,In_947);
or U3860 (N_3860,In_683,In_354);
nor U3861 (N_3861,In_236,In_606);
nor U3862 (N_3862,In_730,In_685);
nor U3863 (N_3863,In_876,In_985);
nand U3864 (N_3864,In_123,In_494);
and U3865 (N_3865,In_527,In_247);
nor U3866 (N_3866,In_505,In_542);
and U3867 (N_3867,In_865,In_326);
and U3868 (N_3868,In_544,In_273);
and U3869 (N_3869,In_22,In_448);
nand U3870 (N_3870,In_619,In_545);
nand U3871 (N_3871,In_337,In_817);
nand U3872 (N_3872,In_452,In_81);
nand U3873 (N_3873,In_762,In_401);
nor U3874 (N_3874,In_255,In_547);
and U3875 (N_3875,In_965,In_50);
or U3876 (N_3876,In_558,In_302);
and U3877 (N_3877,In_963,In_346);
or U3878 (N_3878,In_199,In_320);
and U3879 (N_3879,In_707,In_703);
and U3880 (N_3880,In_625,In_60);
or U3881 (N_3881,In_46,In_84);
xor U3882 (N_3882,In_43,In_324);
nor U3883 (N_3883,In_30,In_352);
and U3884 (N_3884,In_106,In_884);
or U3885 (N_3885,In_170,In_106);
and U3886 (N_3886,In_27,In_641);
or U3887 (N_3887,In_808,In_290);
nor U3888 (N_3888,In_171,In_652);
nand U3889 (N_3889,In_120,In_652);
and U3890 (N_3890,In_466,In_792);
nor U3891 (N_3891,In_489,In_650);
nand U3892 (N_3892,In_417,In_33);
nand U3893 (N_3893,In_407,In_668);
and U3894 (N_3894,In_519,In_722);
or U3895 (N_3895,In_255,In_839);
nand U3896 (N_3896,In_241,In_118);
nand U3897 (N_3897,In_501,In_756);
or U3898 (N_3898,In_990,In_383);
or U3899 (N_3899,In_471,In_896);
and U3900 (N_3900,In_396,In_98);
nand U3901 (N_3901,In_845,In_691);
nor U3902 (N_3902,In_956,In_425);
nor U3903 (N_3903,In_260,In_575);
nand U3904 (N_3904,In_684,In_381);
nand U3905 (N_3905,In_4,In_502);
nor U3906 (N_3906,In_512,In_75);
and U3907 (N_3907,In_858,In_523);
or U3908 (N_3908,In_153,In_138);
and U3909 (N_3909,In_914,In_365);
or U3910 (N_3910,In_134,In_221);
nor U3911 (N_3911,In_759,In_406);
nor U3912 (N_3912,In_98,In_335);
nand U3913 (N_3913,In_494,In_158);
nor U3914 (N_3914,In_660,In_895);
nand U3915 (N_3915,In_508,In_559);
nand U3916 (N_3916,In_18,In_908);
and U3917 (N_3917,In_800,In_979);
or U3918 (N_3918,In_703,In_656);
nand U3919 (N_3919,In_105,In_454);
or U3920 (N_3920,In_824,In_969);
nand U3921 (N_3921,In_649,In_96);
or U3922 (N_3922,In_639,In_96);
or U3923 (N_3923,In_636,In_361);
nor U3924 (N_3924,In_92,In_949);
and U3925 (N_3925,In_208,In_629);
nor U3926 (N_3926,In_604,In_860);
nand U3927 (N_3927,In_868,In_812);
or U3928 (N_3928,In_270,In_468);
and U3929 (N_3929,In_317,In_658);
nor U3930 (N_3930,In_251,In_664);
xor U3931 (N_3931,In_401,In_658);
nor U3932 (N_3932,In_1,In_338);
and U3933 (N_3933,In_598,In_637);
nand U3934 (N_3934,In_519,In_706);
nand U3935 (N_3935,In_600,In_554);
nor U3936 (N_3936,In_182,In_436);
nand U3937 (N_3937,In_781,In_545);
or U3938 (N_3938,In_680,In_165);
xor U3939 (N_3939,In_195,In_592);
nand U3940 (N_3940,In_61,In_586);
or U3941 (N_3941,In_332,In_839);
nand U3942 (N_3942,In_430,In_697);
or U3943 (N_3943,In_818,In_760);
xnor U3944 (N_3944,In_689,In_962);
or U3945 (N_3945,In_433,In_619);
and U3946 (N_3946,In_322,In_738);
nor U3947 (N_3947,In_765,In_502);
or U3948 (N_3948,In_871,In_972);
or U3949 (N_3949,In_454,In_784);
nand U3950 (N_3950,In_276,In_847);
nand U3951 (N_3951,In_155,In_286);
or U3952 (N_3952,In_735,In_58);
xnor U3953 (N_3953,In_579,In_10);
nand U3954 (N_3954,In_580,In_347);
and U3955 (N_3955,In_826,In_232);
nor U3956 (N_3956,In_369,In_893);
nor U3957 (N_3957,In_612,In_364);
or U3958 (N_3958,In_198,In_799);
nand U3959 (N_3959,In_201,In_129);
or U3960 (N_3960,In_162,In_763);
nor U3961 (N_3961,In_502,In_823);
or U3962 (N_3962,In_459,In_447);
nand U3963 (N_3963,In_844,In_388);
and U3964 (N_3964,In_270,In_42);
xnor U3965 (N_3965,In_466,In_500);
and U3966 (N_3966,In_8,In_218);
nand U3967 (N_3967,In_186,In_189);
nand U3968 (N_3968,In_710,In_406);
and U3969 (N_3969,In_353,In_635);
nand U3970 (N_3970,In_185,In_272);
and U3971 (N_3971,In_762,In_379);
and U3972 (N_3972,In_112,In_698);
and U3973 (N_3973,In_816,In_582);
nand U3974 (N_3974,In_520,In_52);
or U3975 (N_3975,In_72,In_607);
xnor U3976 (N_3976,In_486,In_669);
and U3977 (N_3977,In_510,In_802);
xor U3978 (N_3978,In_11,In_156);
and U3979 (N_3979,In_706,In_371);
or U3980 (N_3980,In_556,In_724);
and U3981 (N_3981,In_3,In_794);
and U3982 (N_3982,In_640,In_256);
and U3983 (N_3983,In_416,In_645);
or U3984 (N_3984,In_681,In_675);
and U3985 (N_3985,In_234,In_586);
and U3986 (N_3986,In_808,In_964);
or U3987 (N_3987,In_528,In_575);
nor U3988 (N_3988,In_926,In_605);
nand U3989 (N_3989,In_354,In_293);
and U3990 (N_3990,In_503,In_642);
and U3991 (N_3991,In_874,In_651);
or U3992 (N_3992,In_970,In_156);
and U3993 (N_3993,In_766,In_448);
and U3994 (N_3994,In_709,In_103);
and U3995 (N_3995,In_504,In_817);
nor U3996 (N_3996,In_430,In_901);
and U3997 (N_3997,In_829,In_583);
nand U3998 (N_3998,In_749,In_292);
and U3999 (N_3999,In_578,In_21);
and U4000 (N_4000,In_271,In_527);
and U4001 (N_4001,In_10,In_482);
or U4002 (N_4002,In_618,In_274);
or U4003 (N_4003,In_718,In_973);
and U4004 (N_4004,In_790,In_160);
nor U4005 (N_4005,In_108,In_673);
and U4006 (N_4006,In_166,In_405);
and U4007 (N_4007,In_379,In_963);
nor U4008 (N_4008,In_80,In_989);
nor U4009 (N_4009,In_138,In_407);
and U4010 (N_4010,In_244,In_311);
or U4011 (N_4011,In_42,In_786);
nor U4012 (N_4012,In_644,In_754);
and U4013 (N_4013,In_421,In_679);
nor U4014 (N_4014,In_933,In_210);
nor U4015 (N_4015,In_109,In_395);
and U4016 (N_4016,In_426,In_126);
or U4017 (N_4017,In_188,In_257);
or U4018 (N_4018,In_919,In_846);
nand U4019 (N_4019,In_971,In_920);
nand U4020 (N_4020,In_291,In_469);
nor U4021 (N_4021,In_765,In_760);
nand U4022 (N_4022,In_593,In_232);
nand U4023 (N_4023,In_707,In_826);
or U4024 (N_4024,In_225,In_183);
or U4025 (N_4025,In_953,In_864);
or U4026 (N_4026,In_389,In_302);
and U4027 (N_4027,In_32,In_131);
nor U4028 (N_4028,In_766,In_815);
or U4029 (N_4029,In_420,In_957);
nand U4030 (N_4030,In_36,In_86);
nor U4031 (N_4031,In_792,In_727);
or U4032 (N_4032,In_966,In_955);
nor U4033 (N_4033,In_463,In_868);
or U4034 (N_4034,In_200,In_236);
and U4035 (N_4035,In_139,In_617);
nor U4036 (N_4036,In_128,In_956);
nor U4037 (N_4037,In_68,In_28);
or U4038 (N_4038,In_8,In_817);
nor U4039 (N_4039,In_336,In_421);
or U4040 (N_4040,In_875,In_326);
or U4041 (N_4041,In_746,In_167);
and U4042 (N_4042,In_209,In_1);
or U4043 (N_4043,In_45,In_151);
and U4044 (N_4044,In_564,In_151);
nand U4045 (N_4045,In_60,In_240);
or U4046 (N_4046,In_919,In_856);
or U4047 (N_4047,In_478,In_588);
and U4048 (N_4048,In_263,In_864);
or U4049 (N_4049,In_197,In_15);
nand U4050 (N_4050,In_993,In_15);
nand U4051 (N_4051,In_585,In_115);
nand U4052 (N_4052,In_494,In_329);
or U4053 (N_4053,In_76,In_799);
or U4054 (N_4054,In_300,In_683);
and U4055 (N_4055,In_30,In_895);
xor U4056 (N_4056,In_559,In_917);
nor U4057 (N_4057,In_379,In_859);
nand U4058 (N_4058,In_537,In_726);
or U4059 (N_4059,In_323,In_953);
or U4060 (N_4060,In_379,In_717);
nor U4061 (N_4061,In_453,In_467);
or U4062 (N_4062,In_847,In_974);
nand U4063 (N_4063,In_420,In_707);
or U4064 (N_4064,In_9,In_985);
nor U4065 (N_4065,In_941,In_517);
and U4066 (N_4066,In_154,In_937);
and U4067 (N_4067,In_774,In_503);
nor U4068 (N_4068,In_616,In_447);
or U4069 (N_4069,In_134,In_530);
nor U4070 (N_4070,In_877,In_170);
nor U4071 (N_4071,In_508,In_26);
nand U4072 (N_4072,In_836,In_645);
nor U4073 (N_4073,In_707,In_667);
and U4074 (N_4074,In_319,In_68);
and U4075 (N_4075,In_924,In_999);
and U4076 (N_4076,In_453,In_981);
nor U4077 (N_4077,In_285,In_553);
and U4078 (N_4078,In_204,In_904);
nand U4079 (N_4079,In_525,In_185);
nand U4080 (N_4080,In_541,In_493);
or U4081 (N_4081,In_69,In_873);
nor U4082 (N_4082,In_628,In_936);
nand U4083 (N_4083,In_899,In_662);
nor U4084 (N_4084,In_813,In_430);
nor U4085 (N_4085,In_888,In_889);
xor U4086 (N_4086,In_630,In_815);
and U4087 (N_4087,In_896,In_780);
nand U4088 (N_4088,In_926,In_156);
nand U4089 (N_4089,In_548,In_35);
or U4090 (N_4090,In_836,In_105);
xor U4091 (N_4091,In_307,In_286);
nor U4092 (N_4092,In_352,In_875);
and U4093 (N_4093,In_279,In_193);
or U4094 (N_4094,In_996,In_542);
or U4095 (N_4095,In_407,In_345);
or U4096 (N_4096,In_164,In_252);
xnor U4097 (N_4097,In_727,In_223);
or U4098 (N_4098,In_761,In_870);
or U4099 (N_4099,In_663,In_673);
nand U4100 (N_4100,In_436,In_809);
or U4101 (N_4101,In_907,In_838);
nand U4102 (N_4102,In_595,In_490);
or U4103 (N_4103,In_228,In_185);
or U4104 (N_4104,In_536,In_786);
and U4105 (N_4105,In_989,In_474);
or U4106 (N_4106,In_579,In_51);
nor U4107 (N_4107,In_731,In_766);
or U4108 (N_4108,In_496,In_640);
nor U4109 (N_4109,In_182,In_597);
nand U4110 (N_4110,In_508,In_236);
or U4111 (N_4111,In_724,In_587);
or U4112 (N_4112,In_828,In_128);
or U4113 (N_4113,In_25,In_343);
nand U4114 (N_4114,In_509,In_98);
and U4115 (N_4115,In_694,In_755);
nand U4116 (N_4116,In_13,In_219);
nand U4117 (N_4117,In_587,In_167);
and U4118 (N_4118,In_698,In_982);
or U4119 (N_4119,In_273,In_489);
or U4120 (N_4120,In_683,In_148);
and U4121 (N_4121,In_893,In_611);
and U4122 (N_4122,In_260,In_140);
nor U4123 (N_4123,In_727,In_687);
nor U4124 (N_4124,In_445,In_781);
or U4125 (N_4125,In_53,In_627);
nand U4126 (N_4126,In_609,In_435);
or U4127 (N_4127,In_290,In_440);
nand U4128 (N_4128,In_325,In_14);
xor U4129 (N_4129,In_126,In_879);
or U4130 (N_4130,In_835,In_545);
and U4131 (N_4131,In_271,In_792);
and U4132 (N_4132,In_219,In_596);
and U4133 (N_4133,In_72,In_201);
nand U4134 (N_4134,In_146,In_969);
and U4135 (N_4135,In_713,In_122);
or U4136 (N_4136,In_853,In_146);
nand U4137 (N_4137,In_600,In_670);
or U4138 (N_4138,In_934,In_448);
or U4139 (N_4139,In_809,In_916);
or U4140 (N_4140,In_218,In_456);
and U4141 (N_4141,In_417,In_665);
or U4142 (N_4142,In_62,In_837);
nor U4143 (N_4143,In_67,In_342);
nor U4144 (N_4144,In_336,In_401);
nand U4145 (N_4145,In_198,In_682);
or U4146 (N_4146,In_915,In_954);
and U4147 (N_4147,In_486,In_224);
nand U4148 (N_4148,In_678,In_865);
nor U4149 (N_4149,In_475,In_868);
or U4150 (N_4150,In_259,In_800);
nor U4151 (N_4151,In_482,In_818);
nor U4152 (N_4152,In_369,In_49);
nor U4153 (N_4153,In_473,In_85);
and U4154 (N_4154,In_655,In_157);
nor U4155 (N_4155,In_541,In_135);
nor U4156 (N_4156,In_781,In_293);
or U4157 (N_4157,In_166,In_25);
and U4158 (N_4158,In_935,In_558);
or U4159 (N_4159,In_560,In_265);
and U4160 (N_4160,In_662,In_804);
nor U4161 (N_4161,In_427,In_516);
nor U4162 (N_4162,In_606,In_444);
or U4163 (N_4163,In_743,In_887);
or U4164 (N_4164,In_936,In_578);
xor U4165 (N_4165,In_734,In_301);
nor U4166 (N_4166,In_47,In_918);
or U4167 (N_4167,In_226,In_843);
and U4168 (N_4168,In_15,In_626);
nor U4169 (N_4169,In_93,In_671);
xnor U4170 (N_4170,In_817,In_557);
nand U4171 (N_4171,In_485,In_206);
nand U4172 (N_4172,In_856,In_603);
nand U4173 (N_4173,In_509,In_883);
xor U4174 (N_4174,In_812,In_71);
and U4175 (N_4175,In_720,In_153);
nor U4176 (N_4176,In_513,In_673);
nand U4177 (N_4177,In_275,In_30);
nor U4178 (N_4178,In_136,In_986);
and U4179 (N_4179,In_137,In_984);
and U4180 (N_4180,In_368,In_978);
nand U4181 (N_4181,In_651,In_966);
nor U4182 (N_4182,In_59,In_564);
nor U4183 (N_4183,In_225,In_461);
or U4184 (N_4184,In_88,In_450);
or U4185 (N_4185,In_601,In_514);
xor U4186 (N_4186,In_230,In_457);
nand U4187 (N_4187,In_522,In_59);
and U4188 (N_4188,In_464,In_704);
nand U4189 (N_4189,In_538,In_503);
or U4190 (N_4190,In_145,In_528);
nor U4191 (N_4191,In_133,In_291);
nor U4192 (N_4192,In_844,In_975);
and U4193 (N_4193,In_733,In_300);
and U4194 (N_4194,In_143,In_442);
or U4195 (N_4195,In_670,In_229);
nor U4196 (N_4196,In_515,In_455);
nor U4197 (N_4197,In_747,In_934);
nand U4198 (N_4198,In_52,In_934);
or U4199 (N_4199,In_730,In_510);
nand U4200 (N_4200,In_442,In_648);
and U4201 (N_4201,In_617,In_27);
or U4202 (N_4202,In_537,In_349);
and U4203 (N_4203,In_418,In_659);
or U4204 (N_4204,In_482,In_213);
nor U4205 (N_4205,In_730,In_856);
nor U4206 (N_4206,In_175,In_477);
xnor U4207 (N_4207,In_450,In_873);
and U4208 (N_4208,In_485,In_5);
and U4209 (N_4209,In_159,In_50);
and U4210 (N_4210,In_898,In_236);
or U4211 (N_4211,In_877,In_858);
or U4212 (N_4212,In_471,In_506);
nor U4213 (N_4213,In_213,In_292);
and U4214 (N_4214,In_138,In_955);
nor U4215 (N_4215,In_805,In_186);
and U4216 (N_4216,In_813,In_231);
nand U4217 (N_4217,In_239,In_238);
and U4218 (N_4218,In_826,In_716);
nor U4219 (N_4219,In_296,In_983);
and U4220 (N_4220,In_104,In_495);
and U4221 (N_4221,In_135,In_413);
nand U4222 (N_4222,In_38,In_517);
nor U4223 (N_4223,In_318,In_526);
and U4224 (N_4224,In_195,In_33);
or U4225 (N_4225,In_54,In_631);
and U4226 (N_4226,In_875,In_797);
or U4227 (N_4227,In_475,In_337);
and U4228 (N_4228,In_158,In_502);
nor U4229 (N_4229,In_424,In_643);
or U4230 (N_4230,In_545,In_839);
or U4231 (N_4231,In_95,In_166);
and U4232 (N_4232,In_763,In_861);
nor U4233 (N_4233,In_839,In_758);
and U4234 (N_4234,In_25,In_769);
or U4235 (N_4235,In_96,In_133);
and U4236 (N_4236,In_515,In_785);
or U4237 (N_4237,In_538,In_115);
and U4238 (N_4238,In_175,In_545);
and U4239 (N_4239,In_168,In_279);
or U4240 (N_4240,In_253,In_886);
or U4241 (N_4241,In_789,In_363);
nand U4242 (N_4242,In_471,In_519);
or U4243 (N_4243,In_667,In_939);
xor U4244 (N_4244,In_418,In_539);
nor U4245 (N_4245,In_21,In_983);
and U4246 (N_4246,In_216,In_139);
or U4247 (N_4247,In_319,In_87);
and U4248 (N_4248,In_331,In_238);
nor U4249 (N_4249,In_98,In_612);
or U4250 (N_4250,In_124,In_277);
and U4251 (N_4251,In_609,In_414);
nor U4252 (N_4252,In_484,In_685);
or U4253 (N_4253,In_688,In_93);
and U4254 (N_4254,In_266,In_340);
or U4255 (N_4255,In_598,In_655);
nand U4256 (N_4256,In_40,In_712);
nand U4257 (N_4257,In_598,In_587);
or U4258 (N_4258,In_750,In_557);
nor U4259 (N_4259,In_878,In_796);
nor U4260 (N_4260,In_689,In_169);
nor U4261 (N_4261,In_184,In_742);
and U4262 (N_4262,In_17,In_742);
nand U4263 (N_4263,In_737,In_930);
nor U4264 (N_4264,In_164,In_592);
nor U4265 (N_4265,In_528,In_784);
xnor U4266 (N_4266,In_16,In_922);
or U4267 (N_4267,In_203,In_698);
and U4268 (N_4268,In_729,In_936);
nand U4269 (N_4269,In_206,In_470);
xor U4270 (N_4270,In_573,In_314);
nand U4271 (N_4271,In_443,In_361);
and U4272 (N_4272,In_405,In_978);
nand U4273 (N_4273,In_130,In_544);
or U4274 (N_4274,In_576,In_103);
or U4275 (N_4275,In_483,In_506);
and U4276 (N_4276,In_448,In_555);
or U4277 (N_4277,In_61,In_551);
and U4278 (N_4278,In_623,In_159);
and U4279 (N_4279,In_34,In_247);
and U4280 (N_4280,In_877,In_514);
or U4281 (N_4281,In_360,In_344);
and U4282 (N_4282,In_195,In_763);
and U4283 (N_4283,In_105,In_692);
and U4284 (N_4284,In_81,In_507);
nor U4285 (N_4285,In_393,In_239);
nor U4286 (N_4286,In_86,In_273);
nor U4287 (N_4287,In_123,In_596);
and U4288 (N_4288,In_310,In_795);
nor U4289 (N_4289,In_546,In_461);
or U4290 (N_4290,In_645,In_611);
or U4291 (N_4291,In_924,In_953);
nand U4292 (N_4292,In_352,In_600);
nand U4293 (N_4293,In_104,In_651);
xnor U4294 (N_4294,In_964,In_80);
or U4295 (N_4295,In_310,In_619);
nand U4296 (N_4296,In_819,In_626);
and U4297 (N_4297,In_438,In_439);
and U4298 (N_4298,In_472,In_153);
nand U4299 (N_4299,In_531,In_404);
and U4300 (N_4300,In_414,In_30);
and U4301 (N_4301,In_895,In_274);
or U4302 (N_4302,In_60,In_802);
and U4303 (N_4303,In_829,In_182);
or U4304 (N_4304,In_240,In_311);
nor U4305 (N_4305,In_99,In_860);
nor U4306 (N_4306,In_962,In_876);
or U4307 (N_4307,In_22,In_531);
or U4308 (N_4308,In_942,In_280);
nand U4309 (N_4309,In_733,In_61);
nand U4310 (N_4310,In_664,In_662);
or U4311 (N_4311,In_283,In_831);
or U4312 (N_4312,In_574,In_530);
nor U4313 (N_4313,In_132,In_113);
and U4314 (N_4314,In_75,In_775);
nor U4315 (N_4315,In_204,In_556);
and U4316 (N_4316,In_602,In_629);
nor U4317 (N_4317,In_360,In_599);
and U4318 (N_4318,In_146,In_464);
nand U4319 (N_4319,In_778,In_744);
and U4320 (N_4320,In_570,In_231);
nand U4321 (N_4321,In_5,In_62);
and U4322 (N_4322,In_319,In_857);
or U4323 (N_4323,In_212,In_918);
or U4324 (N_4324,In_371,In_640);
xor U4325 (N_4325,In_836,In_986);
or U4326 (N_4326,In_486,In_938);
nor U4327 (N_4327,In_683,In_950);
and U4328 (N_4328,In_3,In_30);
nand U4329 (N_4329,In_670,In_776);
nand U4330 (N_4330,In_388,In_77);
and U4331 (N_4331,In_572,In_462);
nand U4332 (N_4332,In_685,In_705);
nor U4333 (N_4333,In_243,In_975);
nand U4334 (N_4334,In_776,In_679);
nand U4335 (N_4335,In_575,In_376);
or U4336 (N_4336,In_643,In_755);
or U4337 (N_4337,In_624,In_918);
nor U4338 (N_4338,In_657,In_114);
or U4339 (N_4339,In_323,In_346);
or U4340 (N_4340,In_922,In_910);
nand U4341 (N_4341,In_826,In_249);
or U4342 (N_4342,In_311,In_298);
nor U4343 (N_4343,In_215,In_768);
and U4344 (N_4344,In_341,In_982);
or U4345 (N_4345,In_779,In_446);
or U4346 (N_4346,In_925,In_942);
or U4347 (N_4347,In_509,In_40);
nor U4348 (N_4348,In_903,In_243);
and U4349 (N_4349,In_32,In_240);
nand U4350 (N_4350,In_39,In_675);
nand U4351 (N_4351,In_887,In_934);
or U4352 (N_4352,In_691,In_33);
and U4353 (N_4353,In_166,In_768);
or U4354 (N_4354,In_974,In_786);
and U4355 (N_4355,In_989,In_502);
or U4356 (N_4356,In_247,In_131);
nor U4357 (N_4357,In_628,In_198);
and U4358 (N_4358,In_729,In_625);
and U4359 (N_4359,In_597,In_963);
nand U4360 (N_4360,In_505,In_790);
nor U4361 (N_4361,In_445,In_363);
and U4362 (N_4362,In_244,In_179);
and U4363 (N_4363,In_341,In_259);
nand U4364 (N_4364,In_462,In_701);
nand U4365 (N_4365,In_964,In_723);
nand U4366 (N_4366,In_731,In_672);
and U4367 (N_4367,In_952,In_144);
or U4368 (N_4368,In_857,In_110);
or U4369 (N_4369,In_247,In_36);
nor U4370 (N_4370,In_697,In_293);
or U4371 (N_4371,In_701,In_469);
nor U4372 (N_4372,In_836,In_995);
nand U4373 (N_4373,In_772,In_553);
nand U4374 (N_4374,In_926,In_685);
nand U4375 (N_4375,In_812,In_192);
and U4376 (N_4376,In_105,In_168);
nor U4377 (N_4377,In_180,In_350);
nand U4378 (N_4378,In_477,In_258);
or U4379 (N_4379,In_383,In_347);
and U4380 (N_4380,In_580,In_455);
and U4381 (N_4381,In_139,In_443);
and U4382 (N_4382,In_729,In_134);
nor U4383 (N_4383,In_732,In_600);
nor U4384 (N_4384,In_894,In_554);
or U4385 (N_4385,In_692,In_562);
xor U4386 (N_4386,In_3,In_358);
nand U4387 (N_4387,In_383,In_240);
nor U4388 (N_4388,In_6,In_612);
nand U4389 (N_4389,In_369,In_822);
or U4390 (N_4390,In_561,In_352);
nor U4391 (N_4391,In_576,In_536);
or U4392 (N_4392,In_987,In_37);
and U4393 (N_4393,In_857,In_701);
nand U4394 (N_4394,In_916,In_332);
or U4395 (N_4395,In_73,In_972);
nand U4396 (N_4396,In_986,In_636);
nor U4397 (N_4397,In_163,In_869);
or U4398 (N_4398,In_59,In_924);
nand U4399 (N_4399,In_934,In_611);
and U4400 (N_4400,In_191,In_166);
nor U4401 (N_4401,In_518,In_338);
and U4402 (N_4402,In_131,In_842);
and U4403 (N_4403,In_266,In_253);
and U4404 (N_4404,In_984,In_643);
nand U4405 (N_4405,In_618,In_71);
nor U4406 (N_4406,In_998,In_367);
nand U4407 (N_4407,In_905,In_429);
or U4408 (N_4408,In_85,In_481);
nor U4409 (N_4409,In_61,In_624);
nand U4410 (N_4410,In_96,In_37);
nand U4411 (N_4411,In_629,In_65);
or U4412 (N_4412,In_941,In_246);
nor U4413 (N_4413,In_115,In_862);
or U4414 (N_4414,In_894,In_162);
nand U4415 (N_4415,In_194,In_570);
nor U4416 (N_4416,In_945,In_279);
nor U4417 (N_4417,In_914,In_207);
and U4418 (N_4418,In_668,In_116);
or U4419 (N_4419,In_988,In_493);
or U4420 (N_4420,In_509,In_439);
nand U4421 (N_4421,In_870,In_879);
and U4422 (N_4422,In_909,In_182);
and U4423 (N_4423,In_590,In_772);
nand U4424 (N_4424,In_794,In_527);
and U4425 (N_4425,In_783,In_508);
and U4426 (N_4426,In_694,In_188);
or U4427 (N_4427,In_234,In_682);
and U4428 (N_4428,In_843,In_349);
and U4429 (N_4429,In_437,In_202);
nor U4430 (N_4430,In_399,In_510);
nand U4431 (N_4431,In_514,In_869);
nand U4432 (N_4432,In_1,In_703);
and U4433 (N_4433,In_595,In_271);
nand U4434 (N_4434,In_231,In_255);
or U4435 (N_4435,In_278,In_644);
and U4436 (N_4436,In_627,In_473);
or U4437 (N_4437,In_613,In_351);
and U4438 (N_4438,In_614,In_40);
and U4439 (N_4439,In_141,In_309);
nor U4440 (N_4440,In_324,In_72);
and U4441 (N_4441,In_82,In_102);
nand U4442 (N_4442,In_902,In_231);
nor U4443 (N_4443,In_909,In_126);
and U4444 (N_4444,In_67,In_375);
and U4445 (N_4445,In_378,In_701);
or U4446 (N_4446,In_226,In_505);
or U4447 (N_4447,In_355,In_90);
nor U4448 (N_4448,In_582,In_233);
nand U4449 (N_4449,In_241,In_637);
and U4450 (N_4450,In_481,In_777);
xnor U4451 (N_4451,In_656,In_927);
and U4452 (N_4452,In_384,In_168);
nor U4453 (N_4453,In_891,In_479);
or U4454 (N_4454,In_293,In_190);
xnor U4455 (N_4455,In_151,In_135);
or U4456 (N_4456,In_121,In_922);
and U4457 (N_4457,In_640,In_677);
or U4458 (N_4458,In_621,In_667);
and U4459 (N_4459,In_878,In_900);
nor U4460 (N_4460,In_531,In_90);
or U4461 (N_4461,In_449,In_999);
and U4462 (N_4462,In_155,In_790);
or U4463 (N_4463,In_656,In_585);
nor U4464 (N_4464,In_658,In_220);
nor U4465 (N_4465,In_914,In_242);
or U4466 (N_4466,In_633,In_21);
or U4467 (N_4467,In_622,In_760);
nand U4468 (N_4468,In_187,In_682);
nor U4469 (N_4469,In_693,In_206);
nand U4470 (N_4470,In_842,In_443);
or U4471 (N_4471,In_374,In_3);
or U4472 (N_4472,In_830,In_948);
nand U4473 (N_4473,In_776,In_474);
and U4474 (N_4474,In_68,In_91);
nand U4475 (N_4475,In_912,In_151);
nand U4476 (N_4476,In_896,In_920);
nor U4477 (N_4477,In_333,In_48);
nand U4478 (N_4478,In_269,In_769);
nand U4479 (N_4479,In_767,In_263);
nor U4480 (N_4480,In_580,In_287);
or U4481 (N_4481,In_702,In_481);
nand U4482 (N_4482,In_267,In_964);
nor U4483 (N_4483,In_888,In_458);
and U4484 (N_4484,In_359,In_612);
and U4485 (N_4485,In_454,In_910);
nor U4486 (N_4486,In_770,In_542);
or U4487 (N_4487,In_476,In_276);
nor U4488 (N_4488,In_530,In_292);
or U4489 (N_4489,In_742,In_151);
and U4490 (N_4490,In_821,In_377);
nand U4491 (N_4491,In_683,In_51);
or U4492 (N_4492,In_766,In_225);
and U4493 (N_4493,In_405,In_263);
nor U4494 (N_4494,In_273,In_788);
nand U4495 (N_4495,In_807,In_637);
and U4496 (N_4496,In_352,In_350);
or U4497 (N_4497,In_240,In_156);
and U4498 (N_4498,In_388,In_93);
nor U4499 (N_4499,In_744,In_850);
or U4500 (N_4500,In_843,In_259);
nor U4501 (N_4501,In_736,In_305);
and U4502 (N_4502,In_622,In_83);
nor U4503 (N_4503,In_348,In_673);
and U4504 (N_4504,In_999,In_270);
xor U4505 (N_4505,In_898,In_574);
nor U4506 (N_4506,In_748,In_796);
and U4507 (N_4507,In_288,In_110);
nand U4508 (N_4508,In_593,In_395);
and U4509 (N_4509,In_315,In_30);
nor U4510 (N_4510,In_843,In_952);
nand U4511 (N_4511,In_201,In_547);
or U4512 (N_4512,In_660,In_917);
nor U4513 (N_4513,In_881,In_775);
nor U4514 (N_4514,In_570,In_877);
nand U4515 (N_4515,In_786,In_721);
and U4516 (N_4516,In_191,In_729);
and U4517 (N_4517,In_835,In_96);
or U4518 (N_4518,In_119,In_430);
nand U4519 (N_4519,In_149,In_219);
nor U4520 (N_4520,In_565,In_98);
and U4521 (N_4521,In_660,In_693);
nor U4522 (N_4522,In_192,In_90);
and U4523 (N_4523,In_916,In_465);
and U4524 (N_4524,In_980,In_194);
xor U4525 (N_4525,In_135,In_971);
nand U4526 (N_4526,In_169,In_143);
and U4527 (N_4527,In_82,In_481);
or U4528 (N_4528,In_439,In_495);
or U4529 (N_4529,In_38,In_424);
nand U4530 (N_4530,In_354,In_498);
nor U4531 (N_4531,In_513,In_944);
or U4532 (N_4532,In_634,In_246);
and U4533 (N_4533,In_83,In_14);
nor U4534 (N_4534,In_640,In_989);
and U4535 (N_4535,In_415,In_458);
nor U4536 (N_4536,In_37,In_866);
nor U4537 (N_4537,In_197,In_330);
nand U4538 (N_4538,In_696,In_898);
or U4539 (N_4539,In_169,In_571);
and U4540 (N_4540,In_25,In_436);
or U4541 (N_4541,In_55,In_984);
and U4542 (N_4542,In_988,In_980);
and U4543 (N_4543,In_374,In_104);
and U4544 (N_4544,In_623,In_78);
nor U4545 (N_4545,In_133,In_281);
or U4546 (N_4546,In_665,In_63);
nand U4547 (N_4547,In_321,In_736);
nor U4548 (N_4548,In_431,In_990);
or U4549 (N_4549,In_37,In_380);
or U4550 (N_4550,In_172,In_169);
and U4551 (N_4551,In_152,In_574);
and U4552 (N_4552,In_434,In_75);
nand U4553 (N_4553,In_962,In_703);
nor U4554 (N_4554,In_695,In_296);
nand U4555 (N_4555,In_187,In_674);
nor U4556 (N_4556,In_313,In_708);
nor U4557 (N_4557,In_525,In_132);
and U4558 (N_4558,In_926,In_692);
nand U4559 (N_4559,In_986,In_430);
nand U4560 (N_4560,In_254,In_181);
and U4561 (N_4561,In_583,In_141);
or U4562 (N_4562,In_805,In_119);
nor U4563 (N_4563,In_142,In_875);
or U4564 (N_4564,In_766,In_374);
and U4565 (N_4565,In_52,In_587);
or U4566 (N_4566,In_256,In_850);
nor U4567 (N_4567,In_133,In_413);
or U4568 (N_4568,In_501,In_963);
or U4569 (N_4569,In_850,In_200);
nor U4570 (N_4570,In_873,In_488);
nand U4571 (N_4571,In_133,In_252);
or U4572 (N_4572,In_971,In_475);
nor U4573 (N_4573,In_294,In_485);
nand U4574 (N_4574,In_589,In_594);
nor U4575 (N_4575,In_976,In_864);
or U4576 (N_4576,In_995,In_989);
nand U4577 (N_4577,In_305,In_179);
nand U4578 (N_4578,In_960,In_458);
nor U4579 (N_4579,In_671,In_966);
nor U4580 (N_4580,In_493,In_226);
or U4581 (N_4581,In_775,In_517);
and U4582 (N_4582,In_691,In_36);
nor U4583 (N_4583,In_150,In_701);
and U4584 (N_4584,In_771,In_920);
nor U4585 (N_4585,In_11,In_201);
and U4586 (N_4586,In_130,In_100);
nor U4587 (N_4587,In_407,In_660);
nor U4588 (N_4588,In_330,In_550);
or U4589 (N_4589,In_616,In_664);
nand U4590 (N_4590,In_912,In_979);
or U4591 (N_4591,In_321,In_397);
nor U4592 (N_4592,In_741,In_813);
or U4593 (N_4593,In_235,In_330);
nor U4594 (N_4594,In_487,In_746);
nand U4595 (N_4595,In_437,In_232);
or U4596 (N_4596,In_782,In_345);
nand U4597 (N_4597,In_981,In_582);
or U4598 (N_4598,In_762,In_622);
and U4599 (N_4599,In_121,In_640);
and U4600 (N_4600,In_895,In_57);
or U4601 (N_4601,In_952,In_312);
and U4602 (N_4602,In_986,In_930);
or U4603 (N_4603,In_350,In_162);
nand U4604 (N_4604,In_406,In_78);
and U4605 (N_4605,In_790,In_373);
or U4606 (N_4606,In_41,In_564);
nand U4607 (N_4607,In_955,In_193);
nand U4608 (N_4608,In_828,In_445);
nor U4609 (N_4609,In_311,In_619);
nand U4610 (N_4610,In_195,In_309);
nand U4611 (N_4611,In_103,In_651);
nand U4612 (N_4612,In_987,In_148);
nand U4613 (N_4613,In_797,In_787);
nand U4614 (N_4614,In_750,In_277);
and U4615 (N_4615,In_181,In_227);
nor U4616 (N_4616,In_687,In_3);
nor U4617 (N_4617,In_368,In_348);
and U4618 (N_4618,In_558,In_860);
nor U4619 (N_4619,In_640,In_385);
or U4620 (N_4620,In_160,In_165);
nor U4621 (N_4621,In_398,In_165);
nor U4622 (N_4622,In_880,In_981);
or U4623 (N_4623,In_55,In_871);
nor U4624 (N_4624,In_39,In_489);
nand U4625 (N_4625,In_313,In_443);
nand U4626 (N_4626,In_895,In_130);
or U4627 (N_4627,In_187,In_118);
nor U4628 (N_4628,In_866,In_561);
nand U4629 (N_4629,In_479,In_327);
nor U4630 (N_4630,In_866,In_960);
nor U4631 (N_4631,In_853,In_884);
nor U4632 (N_4632,In_997,In_660);
and U4633 (N_4633,In_58,In_831);
or U4634 (N_4634,In_965,In_573);
nand U4635 (N_4635,In_96,In_697);
xor U4636 (N_4636,In_280,In_34);
and U4637 (N_4637,In_594,In_144);
and U4638 (N_4638,In_406,In_896);
nor U4639 (N_4639,In_84,In_612);
nor U4640 (N_4640,In_51,In_644);
nand U4641 (N_4641,In_197,In_697);
or U4642 (N_4642,In_515,In_116);
nor U4643 (N_4643,In_575,In_214);
or U4644 (N_4644,In_455,In_5);
or U4645 (N_4645,In_898,In_932);
nor U4646 (N_4646,In_68,In_166);
and U4647 (N_4647,In_187,In_128);
nor U4648 (N_4648,In_982,In_385);
nand U4649 (N_4649,In_8,In_777);
nor U4650 (N_4650,In_99,In_709);
and U4651 (N_4651,In_543,In_355);
or U4652 (N_4652,In_176,In_452);
or U4653 (N_4653,In_226,In_488);
and U4654 (N_4654,In_586,In_715);
and U4655 (N_4655,In_227,In_441);
xor U4656 (N_4656,In_888,In_527);
and U4657 (N_4657,In_681,In_996);
or U4658 (N_4658,In_391,In_18);
xnor U4659 (N_4659,In_838,In_333);
nor U4660 (N_4660,In_151,In_793);
nand U4661 (N_4661,In_653,In_25);
and U4662 (N_4662,In_835,In_815);
and U4663 (N_4663,In_779,In_252);
nand U4664 (N_4664,In_518,In_625);
and U4665 (N_4665,In_86,In_642);
nand U4666 (N_4666,In_137,In_77);
or U4667 (N_4667,In_901,In_831);
nand U4668 (N_4668,In_385,In_751);
nor U4669 (N_4669,In_360,In_974);
nor U4670 (N_4670,In_149,In_949);
and U4671 (N_4671,In_5,In_105);
nand U4672 (N_4672,In_483,In_927);
nand U4673 (N_4673,In_126,In_743);
nor U4674 (N_4674,In_723,In_897);
nand U4675 (N_4675,In_943,In_532);
xnor U4676 (N_4676,In_349,In_923);
and U4677 (N_4677,In_90,In_391);
nand U4678 (N_4678,In_484,In_120);
nor U4679 (N_4679,In_757,In_22);
or U4680 (N_4680,In_952,In_686);
and U4681 (N_4681,In_533,In_963);
nor U4682 (N_4682,In_104,In_840);
nor U4683 (N_4683,In_132,In_257);
and U4684 (N_4684,In_769,In_109);
or U4685 (N_4685,In_596,In_422);
or U4686 (N_4686,In_815,In_459);
nand U4687 (N_4687,In_926,In_799);
and U4688 (N_4688,In_927,In_172);
or U4689 (N_4689,In_561,In_776);
nand U4690 (N_4690,In_266,In_776);
and U4691 (N_4691,In_296,In_718);
nand U4692 (N_4692,In_499,In_51);
or U4693 (N_4693,In_37,In_693);
or U4694 (N_4694,In_104,In_269);
or U4695 (N_4695,In_280,In_474);
and U4696 (N_4696,In_595,In_760);
nor U4697 (N_4697,In_289,In_130);
nand U4698 (N_4698,In_803,In_56);
nand U4699 (N_4699,In_569,In_584);
xor U4700 (N_4700,In_532,In_733);
nand U4701 (N_4701,In_503,In_101);
or U4702 (N_4702,In_218,In_949);
or U4703 (N_4703,In_427,In_749);
nor U4704 (N_4704,In_578,In_694);
nand U4705 (N_4705,In_107,In_781);
and U4706 (N_4706,In_594,In_127);
or U4707 (N_4707,In_102,In_318);
nor U4708 (N_4708,In_946,In_117);
nor U4709 (N_4709,In_989,In_67);
and U4710 (N_4710,In_118,In_711);
nor U4711 (N_4711,In_749,In_599);
and U4712 (N_4712,In_622,In_400);
nand U4713 (N_4713,In_495,In_421);
or U4714 (N_4714,In_189,In_736);
nand U4715 (N_4715,In_462,In_926);
nor U4716 (N_4716,In_910,In_553);
or U4717 (N_4717,In_25,In_277);
nor U4718 (N_4718,In_779,In_515);
or U4719 (N_4719,In_819,In_553);
or U4720 (N_4720,In_35,In_534);
nor U4721 (N_4721,In_892,In_228);
nand U4722 (N_4722,In_467,In_376);
nor U4723 (N_4723,In_123,In_800);
and U4724 (N_4724,In_403,In_91);
and U4725 (N_4725,In_488,In_696);
or U4726 (N_4726,In_824,In_837);
and U4727 (N_4727,In_810,In_842);
nor U4728 (N_4728,In_384,In_974);
nor U4729 (N_4729,In_78,In_481);
or U4730 (N_4730,In_870,In_231);
nor U4731 (N_4731,In_233,In_470);
and U4732 (N_4732,In_30,In_355);
and U4733 (N_4733,In_587,In_800);
nand U4734 (N_4734,In_635,In_298);
nor U4735 (N_4735,In_387,In_781);
or U4736 (N_4736,In_641,In_71);
and U4737 (N_4737,In_259,In_302);
or U4738 (N_4738,In_226,In_724);
and U4739 (N_4739,In_849,In_182);
nand U4740 (N_4740,In_3,In_970);
nand U4741 (N_4741,In_191,In_394);
nand U4742 (N_4742,In_596,In_452);
nand U4743 (N_4743,In_338,In_65);
nand U4744 (N_4744,In_73,In_190);
or U4745 (N_4745,In_667,In_315);
nor U4746 (N_4746,In_410,In_672);
and U4747 (N_4747,In_952,In_307);
nor U4748 (N_4748,In_354,In_593);
nand U4749 (N_4749,In_301,In_160);
nand U4750 (N_4750,In_788,In_595);
or U4751 (N_4751,In_437,In_198);
or U4752 (N_4752,In_106,In_149);
and U4753 (N_4753,In_419,In_947);
or U4754 (N_4754,In_72,In_493);
nor U4755 (N_4755,In_818,In_948);
nand U4756 (N_4756,In_240,In_288);
nand U4757 (N_4757,In_196,In_554);
nor U4758 (N_4758,In_383,In_214);
or U4759 (N_4759,In_592,In_995);
and U4760 (N_4760,In_213,In_846);
xnor U4761 (N_4761,In_187,In_745);
nor U4762 (N_4762,In_144,In_703);
nand U4763 (N_4763,In_944,In_579);
and U4764 (N_4764,In_958,In_244);
or U4765 (N_4765,In_869,In_285);
nor U4766 (N_4766,In_700,In_619);
and U4767 (N_4767,In_508,In_395);
or U4768 (N_4768,In_970,In_512);
or U4769 (N_4769,In_35,In_697);
nor U4770 (N_4770,In_904,In_206);
and U4771 (N_4771,In_514,In_980);
or U4772 (N_4772,In_323,In_373);
and U4773 (N_4773,In_544,In_33);
nor U4774 (N_4774,In_25,In_380);
nor U4775 (N_4775,In_735,In_695);
nand U4776 (N_4776,In_42,In_609);
nor U4777 (N_4777,In_660,In_901);
nand U4778 (N_4778,In_435,In_146);
nor U4779 (N_4779,In_911,In_683);
nor U4780 (N_4780,In_122,In_126);
and U4781 (N_4781,In_406,In_762);
nand U4782 (N_4782,In_907,In_372);
nor U4783 (N_4783,In_918,In_950);
nand U4784 (N_4784,In_790,In_138);
or U4785 (N_4785,In_380,In_595);
nor U4786 (N_4786,In_207,In_27);
or U4787 (N_4787,In_282,In_247);
nor U4788 (N_4788,In_274,In_89);
or U4789 (N_4789,In_299,In_97);
and U4790 (N_4790,In_766,In_809);
or U4791 (N_4791,In_714,In_678);
or U4792 (N_4792,In_586,In_925);
or U4793 (N_4793,In_754,In_40);
nor U4794 (N_4794,In_676,In_279);
nor U4795 (N_4795,In_892,In_199);
or U4796 (N_4796,In_192,In_13);
nand U4797 (N_4797,In_984,In_129);
nand U4798 (N_4798,In_610,In_638);
xnor U4799 (N_4799,In_378,In_571);
nand U4800 (N_4800,In_971,In_976);
nor U4801 (N_4801,In_985,In_53);
xor U4802 (N_4802,In_160,In_962);
and U4803 (N_4803,In_637,In_628);
nor U4804 (N_4804,In_138,In_789);
xor U4805 (N_4805,In_598,In_13);
nand U4806 (N_4806,In_32,In_74);
or U4807 (N_4807,In_887,In_795);
or U4808 (N_4808,In_102,In_715);
nor U4809 (N_4809,In_909,In_782);
nor U4810 (N_4810,In_651,In_634);
or U4811 (N_4811,In_952,In_571);
and U4812 (N_4812,In_761,In_101);
nand U4813 (N_4813,In_474,In_933);
and U4814 (N_4814,In_613,In_820);
nand U4815 (N_4815,In_529,In_331);
nand U4816 (N_4816,In_591,In_513);
or U4817 (N_4817,In_378,In_830);
nand U4818 (N_4818,In_905,In_216);
nor U4819 (N_4819,In_75,In_250);
and U4820 (N_4820,In_225,In_618);
nor U4821 (N_4821,In_318,In_811);
nor U4822 (N_4822,In_746,In_958);
nand U4823 (N_4823,In_577,In_786);
nand U4824 (N_4824,In_688,In_247);
nor U4825 (N_4825,In_962,In_879);
nor U4826 (N_4826,In_893,In_141);
xor U4827 (N_4827,In_875,In_878);
or U4828 (N_4828,In_957,In_12);
nand U4829 (N_4829,In_171,In_910);
and U4830 (N_4830,In_451,In_899);
and U4831 (N_4831,In_805,In_375);
nor U4832 (N_4832,In_545,In_27);
nand U4833 (N_4833,In_831,In_987);
and U4834 (N_4834,In_973,In_706);
and U4835 (N_4835,In_22,In_116);
nand U4836 (N_4836,In_529,In_472);
or U4837 (N_4837,In_726,In_433);
nand U4838 (N_4838,In_951,In_762);
and U4839 (N_4839,In_825,In_799);
or U4840 (N_4840,In_85,In_93);
nor U4841 (N_4841,In_20,In_216);
or U4842 (N_4842,In_114,In_934);
and U4843 (N_4843,In_618,In_793);
or U4844 (N_4844,In_256,In_632);
or U4845 (N_4845,In_992,In_240);
nor U4846 (N_4846,In_204,In_746);
nand U4847 (N_4847,In_560,In_7);
nand U4848 (N_4848,In_554,In_743);
or U4849 (N_4849,In_939,In_37);
nand U4850 (N_4850,In_530,In_364);
and U4851 (N_4851,In_432,In_789);
or U4852 (N_4852,In_443,In_305);
nor U4853 (N_4853,In_136,In_300);
and U4854 (N_4854,In_62,In_68);
nand U4855 (N_4855,In_454,In_547);
nand U4856 (N_4856,In_879,In_426);
and U4857 (N_4857,In_691,In_262);
nor U4858 (N_4858,In_185,In_647);
or U4859 (N_4859,In_574,In_44);
nand U4860 (N_4860,In_172,In_491);
and U4861 (N_4861,In_664,In_651);
and U4862 (N_4862,In_484,In_325);
nor U4863 (N_4863,In_350,In_616);
nand U4864 (N_4864,In_581,In_91);
and U4865 (N_4865,In_413,In_278);
nor U4866 (N_4866,In_598,In_908);
nor U4867 (N_4867,In_827,In_625);
nand U4868 (N_4868,In_3,In_781);
or U4869 (N_4869,In_190,In_872);
and U4870 (N_4870,In_532,In_736);
or U4871 (N_4871,In_843,In_825);
nand U4872 (N_4872,In_402,In_724);
nor U4873 (N_4873,In_929,In_637);
nor U4874 (N_4874,In_412,In_531);
nand U4875 (N_4875,In_639,In_667);
nor U4876 (N_4876,In_955,In_700);
or U4877 (N_4877,In_883,In_662);
nand U4878 (N_4878,In_471,In_554);
and U4879 (N_4879,In_521,In_22);
nand U4880 (N_4880,In_103,In_366);
or U4881 (N_4881,In_537,In_665);
nor U4882 (N_4882,In_67,In_174);
or U4883 (N_4883,In_116,In_833);
nor U4884 (N_4884,In_948,In_166);
nand U4885 (N_4885,In_964,In_832);
or U4886 (N_4886,In_214,In_928);
nor U4887 (N_4887,In_349,In_902);
nor U4888 (N_4888,In_406,In_413);
nand U4889 (N_4889,In_95,In_193);
nor U4890 (N_4890,In_84,In_828);
nand U4891 (N_4891,In_119,In_725);
nand U4892 (N_4892,In_800,In_863);
nand U4893 (N_4893,In_945,In_381);
or U4894 (N_4894,In_790,In_911);
nand U4895 (N_4895,In_560,In_792);
or U4896 (N_4896,In_684,In_690);
nand U4897 (N_4897,In_611,In_891);
nand U4898 (N_4898,In_160,In_604);
nor U4899 (N_4899,In_56,In_105);
and U4900 (N_4900,In_21,In_298);
and U4901 (N_4901,In_90,In_248);
or U4902 (N_4902,In_293,In_175);
nand U4903 (N_4903,In_701,In_894);
nor U4904 (N_4904,In_552,In_132);
nor U4905 (N_4905,In_609,In_692);
nand U4906 (N_4906,In_747,In_113);
nand U4907 (N_4907,In_673,In_75);
nand U4908 (N_4908,In_59,In_341);
or U4909 (N_4909,In_992,In_881);
nor U4910 (N_4910,In_542,In_181);
or U4911 (N_4911,In_294,In_668);
and U4912 (N_4912,In_579,In_84);
and U4913 (N_4913,In_906,In_335);
and U4914 (N_4914,In_327,In_401);
and U4915 (N_4915,In_841,In_850);
nor U4916 (N_4916,In_34,In_633);
or U4917 (N_4917,In_157,In_375);
nand U4918 (N_4918,In_518,In_299);
xnor U4919 (N_4919,In_760,In_528);
and U4920 (N_4920,In_736,In_222);
nor U4921 (N_4921,In_138,In_37);
nand U4922 (N_4922,In_489,In_302);
nand U4923 (N_4923,In_924,In_608);
nor U4924 (N_4924,In_118,In_502);
nand U4925 (N_4925,In_42,In_172);
nor U4926 (N_4926,In_21,In_538);
and U4927 (N_4927,In_913,In_878);
and U4928 (N_4928,In_727,In_813);
nand U4929 (N_4929,In_678,In_385);
nand U4930 (N_4930,In_479,In_499);
and U4931 (N_4931,In_175,In_568);
and U4932 (N_4932,In_101,In_650);
nand U4933 (N_4933,In_142,In_305);
or U4934 (N_4934,In_809,In_600);
and U4935 (N_4935,In_324,In_469);
nand U4936 (N_4936,In_852,In_887);
nor U4937 (N_4937,In_489,In_36);
or U4938 (N_4938,In_44,In_263);
and U4939 (N_4939,In_301,In_731);
nor U4940 (N_4940,In_579,In_90);
or U4941 (N_4941,In_685,In_911);
or U4942 (N_4942,In_679,In_253);
xnor U4943 (N_4943,In_239,In_4);
or U4944 (N_4944,In_340,In_487);
nand U4945 (N_4945,In_412,In_714);
and U4946 (N_4946,In_135,In_87);
nand U4947 (N_4947,In_33,In_499);
and U4948 (N_4948,In_610,In_395);
and U4949 (N_4949,In_37,In_834);
xnor U4950 (N_4950,In_324,In_356);
nand U4951 (N_4951,In_274,In_48);
nand U4952 (N_4952,In_84,In_267);
and U4953 (N_4953,In_532,In_381);
xor U4954 (N_4954,In_442,In_773);
nor U4955 (N_4955,In_217,In_758);
nand U4956 (N_4956,In_149,In_502);
or U4957 (N_4957,In_360,In_605);
nand U4958 (N_4958,In_867,In_526);
or U4959 (N_4959,In_484,In_816);
nor U4960 (N_4960,In_569,In_259);
or U4961 (N_4961,In_194,In_154);
xnor U4962 (N_4962,In_979,In_400);
xor U4963 (N_4963,In_631,In_426);
xnor U4964 (N_4964,In_125,In_414);
and U4965 (N_4965,In_560,In_749);
nand U4966 (N_4966,In_982,In_445);
and U4967 (N_4967,In_460,In_84);
xnor U4968 (N_4968,In_408,In_93);
or U4969 (N_4969,In_681,In_955);
or U4970 (N_4970,In_533,In_906);
or U4971 (N_4971,In_5,In_353);
and U4972 (N_4972,In_773,In_342);
or U4973 (N_4973,In_808,In_409);
or U4974 (N_4974,In_988,In_91);
and U4975 (N_4975,In_589,In_247);
nand U4976 (N_4976,In_996,In_315);
and U4977 (N_4977,In_459,In_262);
or U4978 (N_4978,In_95,In_343);
nand U4979 (N_4979,In_907,In_926);
or U4980 (N_4980,In_39,In_374);
nor U4981 (N_4981,In_499,In_467);
nor U4982 (N_4982,In_680,In_305);
nor U4983 (N_4983,In_132,In_941);
and U4984 (N_4984,In_414,In_728);
or U4985 (N_4985,In_105,In_437);
and U4986 (N_4986,In_424,In_774);
and U4987 (N_4987,In_302,In_702);
nand U4988 (N_4988,In_75,In_398);
nand U4989 (N_4989,In_261,In_963);
nand U4990 (N_4990,In_357,In_791);
or U4991 (N_4991,In_427,In_712);
and U4992 (N_4992,In_197,In_630);
and U4993 (N_4993,In_141,In_411);
nor U4994 (N_4994,In_412,In_550);
nand U4995 (N_4995,In_986,In_746);
nor U4996 (N_4996,In_31,In_538);
nand U4997 (N_4997,In_257,In_0);
or U4998 (N_4998,In_311,In_676);
nand U4999 (N_4999,In_366,In_318);
nand U5000 (N_5000,N_3531,N_4407);
nand U5001 (N_5001,N_1370,N_3929);
nor U5002 (N_5002,N_4743,N_3984);
and U5003 (N_5003,N_706,N_4389);
or U5004 (N_5004,N_2656,N_4817);
nor U5005 (N_5005,N_4781,N_4511);
nand U5006 (N_5006,N_2694,N_3343);
nor U5007 (N_5007,N_4212,N_60);
or U5008 (N_5008,N_1512,N_3637);
nor U5009 (N_5009,N_4284,N_4094);
and U5010 (N_5010,N_619,N_2236);
or U5011 (N_5011,N_2814,N_304);
nor U5012 (N_5012,N_2040,N_3155);
nor U5013 (N_5013,N_4206,N_1909);
and U5014 (N_5014,N_2840,N_3028);
nand U5015 (N_5015,N_2316,N_1928);
nor U5016 (N_5016,N_1742,N_3474);
nor U5017 (N_5017,N_2618,N_51);
nor U5018 (N_5018,N_3649,N_1622);
and U5019 (N_5019,N_3255,N_1991);
nand U5020 (N_5020,N_169,N_2621);
nand U5021 (N_5021,N_4967,N_4381);
or U5022 (N_5022,N_3983,N_1365);
or U5023 (N_5023,N_2965,N_830);
nand U5024 (N_5024,N_111,N_4509);
or U5025 (N_5025,N_703,N_3257);
and U5026 (N_5026,N_2189,N_3612);
and U5027 (N_5027,N_4494,N_1193);
nand U5028 (N_5028,N_4460,N_4376);
and U5029 (N_5029,N_810,N_1732);
nand U5030 (N_5030,N_289,N_3442);
nor U5031 (N_5031,N_4708,N_3089);
nor U5032 (N_5032,N_517,N_635);
nand U5033 (N_5033,N_3213,N_2384);
and U5034 (N_5034,N_3045,N_3437);
nand U5035 (N_5035,N_2799,N_4770);
and U5036 (N_5036,N_2169,N_1879);
or U5037 (N_5037,N_2155,N_3628);
or U5038 (N_5038,N_312,N_1472);
nand U5039 (N_5039,N_1848,N_2176);
and U5040 (N_5040,N_1215,N_1858);
nand U5041 (N_5041,N_3116,N_2749);
nor U5042 (N_5042,N_2178,N_698);
or U5043 (N_5043,N_4912,N_1632);
nor U5044 (N_5044,N_2826,N_2370);
and U5045 (N_5045,N_1953,N_2545);
nand U5046 (N_5046,N_4391,N_751);
or U5047 (N_5047,N_3183,N_4790);
and U5048 (N_5048,N_3796,N_1190);
nand U5049 (N_5049,N_1672,N_2372);
and U5050 (N_5050,N_1976,N_4792);
or U5051 (N_5051,N_1534,N_3026);
nand U5052 (N_5052,N_4754,N_2868);
nor U5053 (N_5053,N_1123,N_2308);
or U5054 (N_5054,N_4691,N_4645);
or U5055 (N_5055,N_1683,N_3550);
nor U5056 (N_5056,N_2875,N_4347);
and U5057 (N_5057,N_1001,N_303);
and U5058 (N_5058,N_4066,N_2200);
nand U5059 (N_5059,N_1917,N_3149);
nor U5060 (N_5060,N_753,N_641);
nand U5061 (N_5061,N_1444,N_2170);
or U5062 (N_5062,N_1453,N_1181);
or U5063 (N_5063,N_2100,N_559);
nand U5064 (N_5064,N_2785,N_4906);
nand U5065 (N_5065,N_1091,N_3783);
xor U5066 (N_5066,N_3332,N_4523);
nand U5067 (N_5067,N_1075,N_3635);
and U5068 (N_5068,N_1639,N_904);
nand U5069 (N_5069,N_2118,N_64);
nand U5070 (N_5070,N_3763,N_4749);
nor U5071 (N_5071,N_3173,N_1762);
and U5072 (N_5072,N_3319,N_22);
or U5073 (N_5073,N_3259,N_250);
nor U5074 (N_5074,N_3393,N_4363);
nor U5075 (N_5075,N_808,N_3911);
and U5076 (N_5076,N_3695,N_1097);
nand U5077 (N_5077,N_3373,N_1542);
nor U5078 (N_5078,N_280,N_158);
nand U5079 (N_5079,N_4197,N_2376);
nor U5080 (N_5080,N_2452,N_4163);
nand U5081 (N_5081,N_293,N_3608);
and U5082 (N_5082,N_3340,N_3267);
or U5083 (N_5083,N_3044,N_1127);
or U5084 (N_5084,N_2080,N_759);
nand U5085 (N_5085,N_2904,N_763);
or U5086 (N_5086,N_3392,N_3816);
nor U5087 (N_5087,N_3665,N_1358);
nor U5088 (N_5088,N_3323,N_3966);
nand U5089 (N_5089,N_4510,N_4941);
or U5090 (N_5090,N_1681,N_1495);
or U5091 (N_5091,N_551,N_914);
nor U5092 (N_5092,N_3648,N_649);
nand U5093 (N_5093,N_518,N_1382);
nand U5094 (N_5094,N_4902,N_388);
nand U5095 (N_5095,N_1862,N_574);
and U5096 (N_5096,N_2086,N_2903);
and U5097 (N_5097,N_4151,N_3645);
and U5098 (N_5098,N_2792,N_1043);
nor U5099 (N_5099,N_1188,N_2834);
nor U5100 (N_5100,N_1685,N_29);
nand U5101 (N_5101,N_3072,N_4172);
and U5102 (N_5102,N_2259,N_1787);
nand U5103 (N_5103,N_966,N_3438);
nand U5104 (N_5104,N_2480,N_2944);
or U5105 (N_5105,N_831,N_335);
nor U5106 (N_5106,N_2207,N_3135);
and U5107 (N_5107,N_2960,N_2306);
nor U5108 (N_5108,N_2996,N_3584);
nand U5109 (N_5109,N_4964,N_2024);
nor U5110 (N_5110,N_2326,N_1993);
and U5111 (N_5111,N_2011,N_2349);
and U5112 (N_5112,N_1446,N_2629);
and U5113 (N_5113,N_2289,N_1575);
nor U5114 (N_5114,N_4255,N_836);
nor U5115 (N_5115,N_4506,N_4542);
nand U5116 (N_5116,N_4532,N_1836);
or U5117 (N_5117,N_2988,N_1291);
or U5118 (N_5118,N_389,N_3894);
or U5119 (N_5119,N_2241,N_718);
nor U5120 (N_5120,N_3052,N_4360);
and U5121 (N_5121,N_2194,N_4271);
nor U5122 (N_5122,N_1157,N_936);
xnor U5123 (N_5123,N_410,N_4503);
and U5124 (N_5124,N_3999,N_4880);
nor U5125 (N_5125,N_356,N_3889);
and U5126 (N_5126,N_4348,N_3965);
or U5127 (N_5127,N_3575,N_3679);
nand U5128 (N_5128,N_2589,N_138);
nor U5129 (N_5129,N_3282,N_286);
nand U5130 (N_5130,N_4179,N_1158);
and U5131 (N_5131,N_1202,N_2613);
or U5132 (N_5132,N_2731,N_1037);
or U5133 (N_5133,N_1630,N_870);
nor U5134 (N_5134,N_2757,N_3540);
and U5135 (N_5135,N_3915,N_3959);
nand U5136 (N_5136,N_3095,N_2872);
or U5137 (N_5137,N_1970,N_2899);
and U5138 (N_5138,N_4372,N_1329);
or U5139 (N_5139,N_827,N_1173);
and U5140 (N_5140,N_1261,N_2237);
nor U5141 (N_5141,N_3322,N_4927);
or U5142 (N_5142,N_3779,N_581);
nor U5143 (N_5143,N_3850,N_2935);
nand U5144 (N_5144,N_2524,N_3579);
nor U5145 (N_5145,N_2257,N_4154);
nor U5146 (N_5146,N_2685,N_373);
nor U5147 (N_5147,N_4375,N_903);
nor U5148 (N_5148,N_4125,N_3020);
or U5149 (N_5149,N_2897,N_3450);
nand U5150 (N_5150,N_2739,N_4809);
nand U5151 (N_5151,N_3893,N_3103);
nand U5152 (N_5152,N_3696,N_2560);
nor U5153 (N_5153,N_144,N_4855);
or U5154 (N_5154,N_3892,N_465);
and U5155 (N_5155,N_3593,N_167);
xnor U5156 (N_5156,N_603,N_3444);
nand U5157 (N_5157,N_1416,N_3472);
or U5158 (N_5158,N_3843,N_4400);
nor U5159 (N_5159,N_157,N_917);
or U5160 (N_5160,N_4972,N_1164);
nand U5161 (N_5161,N_4289,N_4742);
nand U5162 (N_5162,N_1564,N_3327);
nor U5163 (N_5163,N_4362,N_909);
nand U5164 (N_5164,N_1341,N_80);
and U5165 (N_5165,N_3204,N_721);
nor U5166 (N_5166,N_196,N_1204);
nand U5167 (N_5167,N_1020,N_1899);
and U5168 (N_5168,N_3449,N_3006);
xnor U5169 (N_5169,N_2361,N_991);
or U5170 (N_5170,N_2993,N_2410);
or U5171 (N_5171,N_2926,N_4968);
nand U5172 (N_5172,N_1196,N_4808);
and U5173 (N_5173,N_1892,N_1840);
nor U5174 (N_5174,N_4890,N_568);
nor U5175 (N_5175,N_4468,N_2555);
and U5176 (N_5176,N_1894,N_2981);
nand U5177 (N_5177,N_3462,N_2715);
nor U5178 (N_5178,N_933,N_376);
nand U5179 (N_5179,N_888,N_4042);
nor U5180 (N_5180,N_1684,N_781);
nor U5181 (N_5181,N_118,N_1999);
nor U5182 (N_5182,N_425,N_3754);
nor U5183 (N_5183,N_2832,N_3195);
and U5184 (N_5184,N_3201,N_4866);
or U5185 (N_5185,N_3709,N_2923);
and U5186 (N_5186,N_955,N_3954);
and U5187 (N_5187,N_4989,N_2846);
nor U5188 (N_5188,N_610,N_287);
nand U5189 (N_5189,N_4692,N_1150);
or U5190 (N_5190,N_4822,N_4061);
and U5191 (N_5191,N_214,N_165);
nor U5192 (N_5192,N_3300,N_3231);
nor U5193 (N_5193,N_4262,N_3249);
or U5194 (N_5194,N_2267,N_2367);
xor U5195 (N_5195,N_2668,N_1465);
and U5196 (N_5196,N_4432,N_3192);
or U5197 (N_5197,N_3566,N_2706);
and U5198 (N_5198,N_1413,N_2862);
xor U5199 (N_5199,N_3368,N_4044);
nor U5200 (N_5200,N_3599,N_826);
nor U5201 (N_5201,N_2424,N_4148);
nand U5202 (N_5202,N_3684,N_1825);
or U5203 (N_5203,N_2640,N_2538);
nand U5204 (N_5204,N_1207,N_4614);
nor U5205 (N_5205,N_3363,N_2609);
and U5206 (N_5206,N_4353,N_1764);
nor U5207 (N_5207,N_3756,N_2340);
nor U5208 (N_5208,N_3944,N_2845);
nand U5209 (N_5209,N_1303,N_2332);
and U5210 (N_5210,N_2117,N_4853);
and U5211 (N_5211,N_2447,N_1431);
nor U5212 (N_5212,N_873,N_4415);
nor U5213 (N_5213,N_4352,N_4040);
nand U5214 (N_5214,N_4938,N_3074);
and U5215 (N_5215,N_3633,N_2321);
nand U5216 (N_5216,N_1708,N_780);
nand U5217 (N_5217,N_3264,N_1344);
nand U5218 (N_5218,N_3718,N_4937);
and U5219 (N_5219,N_3009,N_4520);
nand U5220 (N_5220,N_2179,N_3682);
nand U5221 (N_5221,N_785,N_2743);
nand U5222 (N_5222,N_3036,N_3832);
nor U5223 (N_5223,N_1350,N_1080);
and U5224 (N_5224,N_1113,N_2145);
or U5225 (N_5225,N_2437,N_160);
nand U5226 (N_5226,N_3917,N_37);
and U5227 (N_5227,N_4886,N_3350);
or U5228 (N_5228,N_466,N_2697);
nand U5229 (N_5229,N_3224,N_609);
nor U5230 (N_5230,N_3168,N_4609);
nor U5231 (N_5231,N_747,N_4696);
nor U5232 (N_5232,N_3413,N_4615);
or U5233 (N_5233,N_1323,N_1005);
nor U5234 (N_5234,N_44,N_3023);
and U5235 (N_5235,N_4339,N_3147);
and U5236 (N_5236,N_2659,N_4203);
and U5237 (N_5237,N_1768,N_3172);
or U5238 (N_5238,N_3214,N_1086);
and U5239 (N_5239,N_852,N_219);
nand U5240 (N_5240,N_2476,N_3958);
nor U5241 (N_5241,N_1038,N_3939);
or U5242 (N_5242,N_3736,N_2658);
or U5243 (N_5243,N_2210,N_1015);
or U5244 (N_5244,N_1570,N_876);
and U5245 (N_5245,N_3215,N_883);
nand U5246 (N_5246,N_2772,N_2356);
xnor U5247 (N_5247,N_3537,N_1229);
xnor U5248 (N_5248,N_4297,N_2307);
or U5249 (N_5249,N_3818,N_4078);
and U5250 (N_5250,N_3144,N_4729);
nand U5251 (N_5251,N_1295,N_3650);
nor U5252 (N_5252,N_1849,N_2624);
and U5253 (N_5253,N_947,N_4820);
and U5254 (N_5254,N_1761,N_3447);
and U5255 (N_5255,N_2521,N_4204);
nand U5256 (N_5256,N_2997,N_95);
or U5257 (N_5257,N_1064,N_1);
nand U5258 (N_5258,N_2443,N_3312);
nor U5259 (N_5259,N_2101,N_3957);
and U5260 (N_5260,N_3996,N_1264);
nand U5261 (N_5261,N_4256,N_400);
and U5262 (N_5262,N_2085,N_2603);
and U5263 (N_5263,N_271,N_192);
nand U5264 (N_5264,N_3079,N_151);
or U5265 (N_5265,N_4643,N_1403);
nor U5266 (N_5266,N_916,N_1588);
or U5267 (N_5267,N_2774,N_1275);
and U5268 (N_5268,N_365,N_1581);
nor U5269 (N_5269,N_1304,N_3309);
and U5270 (N_5270,N_3871,N_3466);
and U5271 (N_5271,N_2245,N_4112);
or U5272 (N_5272,N_4785,N_3406);
and U5273 (N_5273,N_1851,N_4192);
nand U5274 (N_5274,N_3184,N_4607);
nor U5275 (N_5275,N_1060,N_2627);
nor U5276 (N_5276,N_795,N_4547);
or U5277 (N_5277,N_1285,N_4246);
nor U5278 (N_5278,N_2346,N_85);
or U5279 (N_5279,N_4208,N_3033);
or U5280 (N_5280,N_3233,N_417);
nor U5281 (N_5281,N_2266,N_409);
or U5282 (N_5282,N_3395,N_1070);
nand U5283 (N_5283,N_3625,N_1900);
nand U5284 (N_5284,N_2453,N_3778);
or U5285 (N_5285,N_490,N_2345);
or U5286 (N_5286,N_3921,N_1362);
nand U5287 (N_5287,N_1852,N_4807);
nand U5288 (N_5288,N_220,N_4756);
and U5289 (N_5289,N_4174,N_1646);
or U5290 (N_5290,N_3586,N_3101);
nor U5291 (N_5291,N_4933,N_1540);
nand U5292 (N_5292,N_3118,N_4776);
nor U5293 (N_5293,N_4536,N_4435);
nor U5294 (N_5294,N_453,N_2277);
or U5295 (N_5295,N_4991,N_1461);
and U5296 (N_5296,N_2752,N_688);
nand U5297 (N_5297,N_1167,N_1593);
nor U5298 (N_5298,N_369,N_4637);
or U5299 (N_5299,N_2272,N_3240);
and U5300 (N_5300,N_4164,N_4568);
and U5301 (N_5301,N_4988,N_2781);
or U5302 (N_5302,N_803,N_1242);
and U5303 (N_5303,N_3037,N_1033);
nand U5304 (N_5304,N_3199,N_403);
nor U5305 (N_5305,N_2371,N_2957);
nor U5306 (N_5306,N_2898,N_4093);
nand U5307 (N_5307,N_4675,N_68);
and U5308 (N_5308,N_2917,N_205);
and U5309 (N_5309,N_4069,N_1738);
or U5310 (N_5310,N_671,N_43);
and U5311 (N_5311,N_1419,N_106);
and U5312 (N_5312,N_4121,N_1192);
and U5313 (N_5313,N_1284,N_2248);
nor U5314 (N_5314,N_1914,N_4513);
nor U5315 (N_5315,N_252,N_4538);
nor U5316 (N_5316,N_1220,N_2279);
or U5317 (N_5317,N_777,N_421);
nor U5318 (N_5318,N_352,N_4089);
nor U5319 (N_5319,N_2830,N_2280);
or U5320 (N_5320,N_4784,N_3286);
or U5321 (N_5321,N_1605,N_3698);
and U5322 (N_5322,N_4404,N_1659);
and U5323 (N_5323,N_2680,N_1682);
and U5324 (N_5324,N_2362,N_3397);
nand U5325 (N_5325,N_1145,N_4916);
and U5326 (N_5326,N_3021,N_2575);
nor U5327 (N_5327,N_1558,N_4814);
nor U5328 (N_5328,N_2554,N_3529);
and U5329 (N_5329,N_4149,N_2761);
and U5330 (N_5330,N_3131,N_2095);
and U5331 (N_5331,N_198,N_3471);
and U5332 (N_5332,N_330,N_3266);
and U5333 (N_5333,N_4438,N_2450);
nor U5334 (N_5334,N_3632,N_912);
nand U5335 (N_5335,N_431,N_2123);
or U5336 (N_5336,N_2696,N_2914);
nand U5337 (N_5337,N_2510,N_4175);
nand U5338 (N_5338,N_1548,N_4947);
nand U5339 (N_5339,N_4114,N_4589);
and U5340 (N_5340,N_710,N_1538);
xor U5341 (N_5341,N_1808,N_1458);
nor U5342 (N_5342,N_272,N_2990);
nand U5343 (N_5343,N_2499,N_4481);
and U5344 (N_5344,N_476,N_2247);
or U5345 (N_5345,N_657,N_1343);
nor U5346 (N_5346,N_2223,N_1779);
nor U5347 (N_5347,N_2835,N_4705);
and U5348 (N_5348,N_1868,N_2771);
nand U5349 (N_5349,N_851,N_1116);
and U5350 (N_5350,N_1478,N_1281);
nand U5351 (N_5351,N_2592,N_2065);
and U5352 (N_5352,N_41,N_997);
xnor U5353 (N_5353,N_392,N_4838);
and U5354 (N_5354,N_1474,N_3247);
xnor U5355 (N_5355,N_3030,N_4434);
nor U5356 (N_5356,N_2181,N_4649);
nor U5357 (N_5357,N_302,N_4054);
nand U5358 (N_5358,N_1788,N_1981);
nand U5359 (N_5359,N_723,N_3658);
or U5360 (N_5360,N_3422,N_1300);
nor U5361 (N_5361,N_174,N_229);
nand U5362 (N_5362,N_3865,N_3459);
or U5363 (N_5363,N_3515,N_4219);
or U5364 (N_5364,N_1009,N_1552);
and U5365 (N_5365,N_2734,N_4448);
and U5366 (N_5366,N_2261,N_4470);
nor U5367 (N_5367,N_199,N_1081);
nor U5368 (N_5368,N_4097,N_3942);
or U5369 (N_5369,N_2166,N_1318);
and U5370 (N_5370,N_1126,N_4118);
nor U5371 (N_5371,N_2577,N_1781);
xor U5372 (N_5372,N_4427,N_3874);
and U5373 (N_5373,N_3069,N_2671);
or U5374 (N_5374,N_3032,N_2754);
nand U5375 (N_5375,N_2355,N_1067);
nor U5376 (N_5376,N_4288,N_3491);
and U5377 (N_5377,N_1835,N_4128);
nor U5378 (N_5378,N_4747,N_3339);
nor U5379 (N_5379,N_4828,N_3949);
and U5380 (N_5380,N_4340,N_2374);
nor U5381 (N_5381,N_3425,N_4270);
or U5382 (N_5382,N_1765,N_2968);
nor U5383 (N_5383,N_3140,N_1147);
or U5384 (N_5384,N_800,N_864);
or U5385 (N_5385,N_3697,N_877);
nor U5386 (N_5386,N_314,N_694);
or U5387 (N_5387,N_4898,N_1120);
and U5388 (N_5388,N_982,N_1813);
nand U5389 (N_5389,N_40,N_2704);
and U5390 (N_5390,N_2707,N_2662);
nor U5391 (N_5391,N_2728,N_1287);
nor U5392 (N_5392,N_481,N_2162);
nand U5393 (N_5393,N_3473,N_3848);
nor U5394 (N_5394,N_3539,N_2796);
nor U5395 (N_5395,N_4981,N_2691);
or U5396 (N_5396,N_2863,N_2420);
and U5397 (N_5397,N_1470,N_2880);
xor U5398 (N_5398,N_4605,N_1490);
nand U5399 (N_5399,N_2687,N_562);
nor U5400 (N_5400,N_1471,N_4628);
and U5401 (N_5401,N_2635,N_2253);
nand U5402 (N_5402,N_1557,N_4582);
nor U5403 (N_5403,N_4337,N_806);
nor U5404 (N_5404,N_4721,N_1774);
and U5405 (N_5405,N_1462,N_646);
or U5406 (N_5406,N_3007,N_998);
nand U5407 (N_5407,N_2809,N_1506);
nand U5408 (N_5408,N_4447,N_4669);
nor U5409 (N_5409,N_1947,N_2164);
or U5410 (N_5410,N_1089,N_4826);
nand U5411 (N_5411,N_2736,N_1078);
and U5412 (N_5412,N_1696,N_1541);
nor U5413 (N_5413,N_918,N_1895);
and U5414 (N_5414,N_1885,N_3071);
nor U5415 (N_5415,N_2719,N_2989);
and U5416 (N_5416,N_404,N_345);
and U5417 (N_5417,N_3511,N_3513);
nand U5418 (N_5418,N_1109,N_4567);
nor U5419 (N_5419,N_3411,N_879);
nor U5420 (N_5420,N_3156,N_3798);
or U5421 (N_5421,N_31,N_3245);
nand U5422 (N_5422,N_1930,N_2583);
nor U5423 (N_5423,N_3553,N_3533);
or U5424 (N_5424,N_2571,N_4515);
xor U5425 (N_5425,N_3930,N_2354);
nand U5426 (N_5426,N_3976,N_832);
and U5427 (N_5427,N_637,N_3617);
or U5428 (N_5428,N_4728,N_4730);
or U5429 (N_5429,N_942,N_3905);
or U5430 (N_5430,N_891,N_3349);
nand U5431 (N_5431,N_4298,N_1767);
or U5432 (N_5432,N_3752,N_605);
nand U5433 (N_5433,N_2877,N_1636);
nor U5434 (N_5434,N_3295,N_3112);
xor U5435 (N_5435,N_3817,N_3918);
and U5436 (N_5436,N_306,N_739);
nor U5437 (N_5437,N_1122,N_2490);
nand U5438 (N_5438,N_3968,N_62);
nor U5439 (N_5439,N_915,N_3497);
or U5440 (N_5440,N_4188,N_1971);
or U5441 (N_5441,N_3283,N_1460);
nor U5442 (N_5442,N_770,N_310);
and U5443 (N_5443,N_3613,N_1189);
and U5444 (N_5444,N_1503,N_1853);
and U5445 (N_5445,N_1386,N_679);
and U5446 (N_5446,N_4904,N_658);
nand U5447 (N_5447,N_3912,N_2018);
nand U5448 (N_5448,N_2353,N_3807);
nor U5449 (N_5449,N_572,N_2278);
nor U5450 (N_5450,N_1907,N_1002);
nand U5451 (N_5451,N_3429,N_4940);
or U5452 (N_5452,N_3256,N_1749);
nand U5453 (N_5453,N_4016,N_3435);
and U5454 (N_5454,N_2646,N_4797);
or U5455 (N_5455,N_372,N_4517);
or U5456 (N_5456,N_3624,N_4757);
or U5457 (N_5457,N_83,N_4959);
nand U5458 (N_5458,N_2422,N_4578);
and U5459 (N_5459,N_2888,N_3707);
and U5460 (N_5460,N_1141,N_341);
nor U5461 (N_5461,N_1421,N_597);
or U5462 (N_5462,N_57,N_3081);
or U5463 (N_5463,N_2458,N_1838);
and U5464 (N_5464,N_4346,N_4952);
or U5465 (N_5465,N_2188,N_1714);
and U5466 (N_5466,N_13,N_3995);
or U5467 (N_5467,N_1850,N_604);
and U5468 (N_5468,N_3065,N_2434);
nand U5469 (N_5469,N_4722,N_2240);
nor U5470 (N_5470,N_1338,N_1912);
and U5471 (N_5471,N_4020,N_1227);
and U5472 (N_5472,N_1000,N_3152);
xor U5473 (N_5473,N_73,N_1448);
nor U5474 (N_5474,N_101,N_3787);
and U5475 (N_5475,N_2869,N_1745);
or U5476 (N_5476,N_543,N_2206);
nor U5477 (N_5477,N_321,N_2400);
xnor U5478 (N_5478,N_3879,N_3062);
or U5479 (N_5479,N_3451,N_1315);
nor U5480 (N_5480,N_1870,N_2462);
and U5481 (N_5481,N_821,N_1452);
nand U5482 (N_5482,N_2740,N_450);
or U5483 (N_5483,N_4131,N_4584);
xor U5484 (N_5484,N_4882,N_889);
and U5485 (N_5485,N_3924,N_15);
nand U5486 (N_5486,N_849,N_4323);
and U5487 (N_5487,N_1496,N_4127);
or U5488 (N_5488,N_980,N_1677);
nor U5489 (N_5489,N_4133,N_2408);
or U5490 (N_5490,N_4571,N_4107);
nor U5491 (N_5491,N_2758,N_1637);
nor U5492 (N_5492,N_2182,N_2587);
nor U5493 (N_5493,N_4058,N_1039);
nor U5494 (N_5494,N_4413,N_3269);
and U5495 (N_5495,N_4563,N_2448);
and U5496 (N_5496,N_3860,N_4878);
nor U5497 (N_5497,N_4587,N_4081);
and U5498 (N_5498,N_3133,N_4630);
and U5499 (N_5499,N_2947,N_1601);
nor U5500 (N_5500,N_3086,N_4593);
and U5501 (N_5501,N_4580,N_4034);
and U5502 (N_5502,N_4220,N_3986);
nor U5503 (N_5503,N_4970,N_754);
and U5504 (N_5504,N_1255,N_4358);
and U5505 (N_5505,N_789,N_2165);
nand U5506 (N_5506,N_3382,N_4313);
nand U5507 (N_5507,N_2218,N_259);
and U5508 (N_5508,N_4813,N_612);
nand U5509 (N_5509,N_3398,N_262);
nand U5510 (N_5510,N_1212,N_268);
or U5511 (N_5511,N_4244,N_4857);
nand U5512 (N_5512,N_1022,N_422);
nand U5513 (N_5513,N_1582,N_1877);
nor U5514 (N_5514,N_2813,N_3815);
or U5515 (N_5515,N_794,N_1201);
and U5516 (N_5516,N_3381,N_1004);
or U5517 (N_5517,N_2336,N_1290);
nand U5518 (N_5518,N_1594,N_2631);
nor U5519 (N_5519,N_4555,N_2481);
nor U5520 (N_5520,N_1138,N_1501);
nor U5521 (N_5521,N_2233,N_3002);
nand U5522 (N_5522,N_2526,N_617);
and U5523 (N_5523,N_2397,N_4960);
nand U5524 (N_5524,N_344,N_626);
nand U5525 (N_5525,N_588,N_4268);
and U5526 (N_5526,N_4726,N_2216);
nor U5527 (N_5527,N_1248,N_3080);
and U5528 (N_5528,N_1463,N_4803);
and U5529 (N_5529,N_320,N_872);
or U5530 (N_5530,N_1741,N_2652);
and U5531 (N_5531,N_2660,N_1938);
xnor U5532 (N_5532,N_491,N_1871);
and U5533 (N_5533,N_3318,N_2377);
or U5534 (N_5534,N_3262,N_4486);
or U5535 (N_5535,N_3853,N_4746);
or U5536 (N_5536,N_4039,N_1385);
or U5537 (N_5537,N_1923,N_2075);
or U5538 (N_5538,N_2887,N_2387);
and U5539 (N_5539,N_3278,N_482);
nor U5540 (N_5540,N_2031,N_501);
nand U5541 (N_5541,N_4939,N_2578);
nand U5542 (N_5542,N_1572,N_1922);
nand U5543 (N_5543,N_3847,N_4601);
nand U5544 (N_5544,N_2630,N_3059);
nor U5545 (N_5545,N_2003,N_2405);
or U5546 (N_5546,N_11,N_3358);
nor U5547 (N_5547,N_2022,N_3055);
nand U5548 (N_5548,N_69,N_1962);
or U5549 (N_5549,N_4209,N_1296);
or U5550 (N_5550,N_4146,N_2654);
nand U5551 (N_5551,N_3580,N_3724);
or U5552 (N_5552,N_4059,N_179);
or U5553 (N_5553,N_1066,N_4693);
nand U5554 (N_5554,N_495,N_3132);
or U5555 (N_5555,N_4177,N_1802);
nand U5556 (N_5556,N_840,N_494);
nand U5557 (N_5557,N_1530,N_2185);
and U5558 (N_5558,N_815,N_4390);
or U5559 (N_5559,N_3070,N_1368);
and U5560 (N_5560,N_2128,N_1104);
nand U5561 (N_5561,N_816,N_3610);
nor U5562 (N_5562,N_1620,N_1292);
nor U5563 (N_5563,N_3506,N_1252);
nor U5564 (N_5564,N_2763,N_768);
nand U5565 (N_5565,N_2726,N_4852);
nand U5566 (N_5566,N_4731,N_2946);
nor U5567 (N_5567,N_3297,N_3559);
and U5568 (N_5568,N_3730,N_3621);
nor U5569 (N_5569,N_3468,N_88);
nor U5570 (N_5570,N_3234,N_2812);
and U5571 (N_5571,N_2665,N_659);
nor U5572 (N_5572,N_4865,N_4030);
or U5573 (N_5573,N_758,N_274);
nor U5574 (N_5574,N_714,N_4987);
nor U5575 (N_5575,N_393,N_2135);
nor U5576 (N_5576,N_4779,N_1746);
and U5577 (N_5577,N_467,N_2058);
and U5578 (N_5578,N_1467,N_3565);
or U5579 (N_5579,N_1532,N_2108);
nand U5580 (N_5580,N_4153,N_416);
nor U5581 (N_5581,N_654,N_1239);
or U5582 (N_5582,N_2843,N_4440);
nor U5583 (N_5583,N_822,N_2784);
and U5584 (N_5584,N_3913,N_1951);
and U5585 (N_5585,N_3352,N_4545);
or U5586 (N_5586,N_1535,N_1380);
nor U5587 (N_5587,N_3744,N_2504);
or U5588 (N_5588,N_2663,N_4342);
nor U5589 (N_5589,N_197,N_3602);
or U5590 (N_5590,N_2674,N_4260);
and U5591 (N_5591,N_1363,N_2493);
nand U5592 (N_5592,N_3713,N_4805);
nor U5593 (N_5593,N_2442,N_3833);
and U5594 (N_5594,N_19,N_4178);
nor U5595 (N_5595,N_2722,N_2385);
nand U5596 (N_5596,N_4664,N_3680);
and U5597 (N_5597,N_3826,N_4672);
or U5598 (N_5598,N_673,N_4889);
or U5599 (N_5599,N_2150,N_136);
and U5600 (N_5600,N_30,N_4974);
or U5601 (N_5601,N_1356,N_950);
and U5602 (N_5602,N_277,N_724);
or U5603 (N_5603,N_1182,N_2357);
and U5604 (N_5604,N_672,N_1502);
or U5605 (N_5605,N_1168,N_722);
nand U5606 (N_5606,N_1719,N_4325);
nand U5607 (N_5607,N_56,N_4479);
nor U5608 (N_5608,N_2298,N_2548);
or U5609 (N_5609,N_3043,N_552);
nand U5610 (N_5610,N_1505,N_1199);
or U5611 (N_5611,N_3235,N_4102);
nand U5612 (N_5612,N_2431,N_2684);
nor U5613 (N_5613,N_1750,N_2829);
nand U5614 (N_5614,N_2334,N_4526);
or U5615 (N_5615,N_3606,N_503);
or U5616 (N_5616,N_492,N_4228);
and U5617 (N_5617,N_2622,N_2036);
nand U5618 (N_5618,N_1891,N_2816);
nor U5619 (N_5619,N_1528,N_4702);
nand U5620 (N_5620,N_3308,N_1687);
and U5621 (N_5621,N_582,N_49);
or U5622 (N_5622,N_4648,N_596);
nor U5623 (N_5623,N_1011,N_1616);
nand U5624 (N_5624,N_3909,N_4695);
nor U5625 (N_5625,N_173,N_2632);
nand U5626 (N_5626,N_3414,N_4798);
or U5627 (N_5627,N_3167,N_3012);
and U5628 (N_5628,N_1982,N_2789);
nor U5629 (N_5629,N_3501,N_550);
and U5630 (N_5630,N_1758,N_3683);
and U5631 (N_5631,N_4918,N_4045);
nand U5632 (N_5632,N_4195,N_1125);
and U5633 (N_5633,N_3225,N_2274);
or U5634 (N_5634,N_206,N_2131);
nor U5635 (N_5635,N_224,N_3872);
or U5636 (N_5636,N_4639,N_3864);
nand U5637 (N_5637,N_4429,N_3379);
or U5638 (N_5638,N_969,N_1845);
or U5639 (N_5639,N_4401,N_4529);
nand U5640 (N_5640,N_546,N_3973);
and U5641 (N_5641,N_801,N_3547);
or U5642 (N_5642,N_1366,N_2760);
nor U5643 (N_5643,N_523,N_1556);
nor U5644 (N_5644,N_4380,N_2963);
and U5645 (N_5645,N_1469,N_3465);
nand U5646 (N_5646,N_4258,N_2797);
nor U5647 (N_5647,N_23,N_1367);
or U5648 (N_5648,N_2655,N_3542);
or U5649 (N_5649,N_2417,N_4296);
and U5650 (N_5650,N_2767,N_3955);
or U5651 (N_5651,N_2876,N_1966);
or U5652 (N_5652,N_2305,N_4160);
or U5653 (N_5653,N_1863,N_1235);
nor U5654 (N_5654,N_765,N_1222);
or U5655 (N_5655,N_1832,N_4387);
and U5656 (N_5656,N_504,N_1092);
nor U5657 (N_5657,N_1280,N_2879);
and U5658 (N_5658,N_4367,N_730);
and U5659 (N_5659,N_1887,N_1625);
nand U5660 (N_5660,N_3596,N_1324);
and U5661 (N_5661,N_1645,N_4856);
or U5662 (N_5662,N_1153,N_3115);
or U5663 (N_5663,N_2154,N_2120);
and U5664 (N_5664,N_2874,N_4329);
and U5665 (N_5665,N_707,N_2099);
nand U5666 (N_5666,N_4189,N_1137);
or U5667 (N_5667,N_4285,N_1468);
and U5668 (N_5668,N_1526,N_1939);
nor U5669 (N_5669,N_1019,N_3508);
and U5670 (N_5670,N_2536,N_325);
nor U5671 (N_5671,N_3799,N_368);
or U5672 (N_5672,N_3664,N_2885);
and U5673 (N_5673,N_1456,N_2045);
nor U5674 (N_5674,N_4026,N_1615);
nand U5675 (N_5675,N_2498,N_38);
or U5676 (N_5676,N_1241,N_2337);
or U5677 (N_5677,N_2992,N_4671);
nand U5678 (N_5678,N_2005,N_4800);
nor U5679 (N_5679,N_1057,N_1664);
nand U5680 (N_5680,N_835,N_4074);
or U5681 (N_5681,N_4444,N_2803);
or U5682 (N_5682,N_828,N_4963);
or U5683 (N_5683,N_1800,N_3162);
nor U5684 (N_5684,N_536,N_4677);
and U5685 (N_5685,N_2225,N_2148);
nand U5686 (N_5686,N_1434,N_4504);
and U5687 (N_5687,N_2016,N_4858);
and U5688 (N_5688,N_2678,N_509);
or U5689 (N_5689,N_2124,N_4821);
nor U5690 (N_5690,N_3216,N_2837);
and U5691 (N_5691,N_3385,N_2343);
and U5692 (N_5692,N_3927,N_560);
nand U5693 (N_5693,N_329,N_1319);
or U5694 (N_5694,N_2235,N_825);
nor U5695 (N_5695,N_618,N_3767);
xnor U5696 (N_5696,N_3761,N_1059);
or U5697 (N_5697,N_2986,N_33);
and U5698 (N_5698,N_2730,N_343);
xor U5699 (N_5699,N_3509,N_305);
nor U5700 (N_5700,N_4090,N_3803);
nand U5701 (N_5701,N_2636,N_3375);
nor U5702 (N_5702,N_3150,N_4759);
nor U5703 (N_5703,N_4793,N_267);
nor U5704 (N_5704,N_1258,N_899);
or U5705 (N_5705,N_4752,N_4281);
nand U5706 (N_5706,N_3212,N_2394);
and U5707 (N_5707,N_4579,N_163);
or U5708 (N_5708,N_638,N_4765);
or U5709 (N_5709,N_371,N_2076);
nor U5710 (N_5710,N_4392,N_4948);
or U5711 (N_5711,N_3090,N_2461);
or U5712 (N_5712,N_4287,N_1712);
nor U5713 (N_5713,N_4911,N_248);
nor U5714 (N_5714,N_2964,N_3503);
and U5715 (N_5715,N_3177,N_592);
nor U5716 (N_5716,N_4023,N_82);
and U5717 (N_5717,N_1673,N_2407);
and U5718 (N_5718,N_4119,N_4319);
and U5719 (N_5719,N_258,N_775);
or U5720 (N_5720,N_2328,N_420);
nor U5721 (N_5721,N_1805,N_1427);
nor U5722 (N_5722,N_2029,N_3523);
and U5723 (N_5723,N_3861,N_1376);
nand U5724 (N_5724,N_4561,N_4229);
or U5725 (N_5725,N_4185,N_3326);
and U5726 (N_5726,N_1806,N_1210);
nor U5727 (N_5727,N_1119,N_4958);
nor U5728 (N_5728,N_1908,N_3415);
nor U5729 (N_5729,N_200,N_432);
and U5730 (N_5730,N_2717,N_4426);
nor U5731 (N_5731,N_2535,N_216);
and U5732 (N_5732,N_4859,N_2167);
nand U5733 (N_5733,N_2313,N_945);
and U5734 (N_5734,N_2047,N_4100);
or U5735 (N_5735,N_3194,N_4231);
and U5736 (N_5736,N_699,N_3142);
nand U5737 (N_5737,N_4184,N_3281);
and U5738 (N_5738,N_2995,N_4531);
or U5739 (N_5739,N_1406,N_4461);
and U5740 (N_5740,N_4328,N_2637);
nand U5741 (N_5741,N_3925,N_284);
xnor U5742 (N_5742,N_238,N_2574);
nor U5743 (N_5743,N_3384,N_3717);
or U5744 (N_5744,N_748,N_1834);
and U5745 (N_5745,N_241,N_2657);
and U5746 (N_5746,N_4462,N_3200);
and U5747 (N_5747,N_2351,N_3388);
nand U5748 (N_5748,N_4453,N_3792);
and U5749 (N_5749,N_2870,N_4070);
and U5750 (N_5750,N_978,N_1975);
nor U5751 (N_5751,N_150,N_4971);
or U5752 (N_5752,N_3590,N_379);
nor U5753 (N_5753,N_3022,N_772);
or U5754 (N_5754,N_2956,N_257);
and U5755 (N_5755,N_1166,N_4221);
or U5756 (N_5756,N_3087,N_1035);
nor U5757 (N_5757,N_1392,N_3337);
nor U5758 (N_5758,N_3175,N_2692);
and U5759 (N_5759,N_2470,N_4572);
nand U5760 (N_5760,N_1509,N_1180);
nand U5761 (N_5761,N_2317,N_119);
or U5762 (N_5762,N_1933,N_2133);
or U5763 (N_5763,N_1320,N_2038);
nand U5764 (N_5764,N_1786,N_294);
or U5765 (N_5765,N_1650,N_3299);
nand U5766 (N_5766,N_2455,N_2441);
nand U5767 (N_5767,N_2161,N_1432);
or U5768 (N_5768,N_397,N_741);
or U5769 (N_5769,N_1797,N_4825);
and U5770 (N_5770,N_4488,N_1108);
nor U5771 (N_5771,N_2054,N_4657);
nor U5772 (N_5772,N_2712,N_3524);
and U5773 (N_5773,N_26,N_693);
nand U5774 (N_5774,N_182,N_391);
or U5775 (N_5775,N_1629,N_1203);
nand U5776 (N_5776,N_3127,N_4245);
nor U5777 (N_5777,N_1114,N_3181);
and U5778 (N_5778,N_4576,N_2020);
nor U5779 (N_5779,N_292,N_2163);
or U5780 (N_5780,N_1734,N_3841);
and U5781 (N_5781,N_3475,N_488);
or U5782 (N_5782,N_1163,N_3545);
nor U5783 (N_5783,N_3124,N_3171);
and U5784 (N_5784,N_4611,N_2679);
or U5785 (N_5785,N_1995,N_442);
or U5786 (N_5786,N_4559,N_3364);
nand U5787 (N_5787,N_4935,N_1003);
or U5788 (N_5788,N_1511,N_1045);
nand U5789 (N_5789,N_2388,N_731);
and U5790 (N_5790,N_2810,N_3700);
nor U5791 (N_5791,N_127,N_1510);
and U5792 (N_5792,N_652,N_1165);
nand U5793 (N_5793,N_4084,N_4627);
nand U5794 (N_5794,N_4129,N_2765);
and U5795 (N_5795,N_3421,N_2406);
and U5796 (N_5796,N_4211,N_113);
and U5797 (N_5797,N_102,N_510);
or U5798 (N_5798,N_2186,N_3239);
nand U5799 (N_5799,N_3538,N_3722);
nand U5800 (N_5800,N_4439,N_67);
nor U5801 (N_5801,N_3246,N_1579);
or U5802 (N_5802,N_1860,N_3076);
nand U5803 (N_5803,N_2382,N_2667);
nand U5804 (N_5804,N_4783,N_318);
nand U5805 (N_5805,N_4320,N_745);
nor U5806 (N_5806,N_4198,N_210);
and U5807 (N_5807,N_611,N_902);
nor U5808 (N_5808,N_4408,N_4333);
or U5809 (N_5809,N_3950,N_2202);
or U5810 (N_5810,N_3035,N_2239);
nor U5811 (N_5811,N_3389,N_4796);
xnor U5812 (N_5812,N_181,N_3003);
and U5813 (N_5813,N_4945,N_3528);
nor U5814 (N_5814,N_2841,N_3794);
or U5815 (N_5815,N_4965,N_4895);
xnor U5816 (N_5816,N_3616,N_4299);
and U5817 (N_5817,N_211,N_1896);
and U5818 (N_5818,N_434,N_2488);
nor U5819 (N_5819,N_3187,N_2927);
nand U5820 (N_5820,N_4629,N_4951);
nand U5821 (N_5821,N_3254,N_4004);
nand U5822 (N_5822,N_4080,N_989);
nand U5823 (N_5823,N_4143,N_1929);
or U5824 (N_5824,N_1507,N_1387);
or U5825 (N_5825,N_2070,N_2283);
or U5826 (N_5826,N_3998,N_1283);
and U5827 (N_5827,N_1179,N_4324);
and U5828 (N_5828,N_4193,N_3734);
or U5829 (N_5829,N_1671,N_734);
nor U5830 (N_5830,N_406,N_4524);
nor U5831 (N_5831,N_2484,N_3834);
nand U5832 (N_5832,N_905,N_162);
xnor U5833 (N_5833,N_4962,N_4837);
nor U5834 (N_5834,N_4183,N_4101);
or U5835 (N_5835,N_1230,N_935);
and U5836 (N_5836,N_4845,N_2358);
and U5837 (N_5837,N_3250,N_1331);
nor U5838 (N_5838,N_4064,N_1935);
and U5839 (N_5839,N_4412,N_2197);
and U5840 (N_5840,N_2865,N_115);
and U5841 (N_5841,N_3849,N_1657);
and U5842 (N_5842,N_4003,N_2010);
and U5843 (N_5843,N_1099,N_3750);
or U5844 (N_5844,N_1942,N_1216);
and U5845 (N_5845,N_4920,N_2119);
or U5846 (N_5846,N_1977,N_650);
and U5847 (N_5847,N_4010,N_477);
or U5848 (N_5848,N_732,N_3814);
or U5849 (N_5849,N_437,N_3604);
nand U5850 (N_5850,N_3926,N_4418);
nand U5851 (N_5851,N_3952,N_705);
nor U5852 (N_5852,N_4684,N_4405);
nand U5853 (N_5853,N_848,N_4786);
nor U5854 (N_5854,N_4286,N_3298);
and U5855 (N_5855,N_613,N_1430);
nor U5856 (N_5856,N_1451,N_3788);
nor U5857 (N_5857,N_3370,N_1964);
nor U5858 (N_5858,N_21,N_2090);
and U5859 (N_5859,N_4588,N_956);
or U5860 (N_5860,N_3705,N_4103);
nand U5861 (N_5861,N_2824,N_2572);
and U5862 (N_5862,N_4884,N_786);
and U5863 (N_5863,N_3587,N_4969);
nand U5864 (N_5864,N_2955,N_2616);
and U5865 (N_5865,N_2485,N_377);
or U5866 (N_5866,N_4306,N_1859);
nor U5867 (N_5867,N_995,N_4507);
or U5868 (N_5868,N_1335,N_1748);
or U5869 (N_5869,N_4500,N_4303);
nand U5870 (N_5870,N_339,N_823);
nor U5871 (N_5871,N_4758,N_3399);
nand U5872 (N_5872,N_3771,N_3898);
nor U5873 (N_5873,N_4723,N_2729);
nor U5874 (N_5874,N_3313,N_4946);
nand U5875 (N_5875,N_2294,N_4550);
or U5876 (N_5876,N_455,N_941);
or U5877 (N_5877,N_2111,N_4626);
nor U5878 (N_5878,N_1647,N_4586);
or U5879 (N_5879,N_4158,N_3077);
nor U5880 (N_5880,N_418,N_541);
nand U5881 (N_5881,N_773,N_4982);
nor U5882 (N_5882,N_3431,N_3242);
nand U5883 (N_5883,N_3117,N_4369);
or U5884 (N_5884,N_4768,N_2140);
and U5885 (N_5885,N_2177,N_4022);
or U5886 (N_5886,N_3108,N_3922);
nand U5887 (N_5887,N_1151,N_528);
and U5888 (N_5888,N_4295,N_3934);
nor U5889 (N_5889,N_4766,N_736);
or U5890 (N_5890,N_4242,N_4508);
nor U5891 (N_5891,N_616,N_2860);
nand U5892 (N_5892,N_4464,N_3857);
and U5893 (N_5893,N_4983,N_3806);
nor U5894 (N_5894,N_704,N_63);
nand U5895 (N_5895,N_2605,N_1606);
and U5896 (N_5896,N_2501,N_3663);
nand U5897 (N_5897,N_361,N_3039);
and U5898 (N_5898,N_2171,N_529);
and U5899 (N_5899,N_975,N_2060);
nor U5900 (N_5900,N_2762,N_2092);
nor U5901 (N_5901,N_3279,N_1724);
and U5902 (N_5902,N_4232,N_1607);
and U5903 (N_5903,N_1198,N_2976);
or U5904 (N_5904,N_1653,N_2445);
nor U5905 (N_5905,N_2744,N_4840);
and U5906 (N_5906,N_4733,N_4724);
nand U5907 (N_5907,N_1438,N_486);
and U5908 (N_5908,N_2910,N_1381);
nor U5909 (N_5909,N_3193,N_4548);
nor U5910 (N_5910,N_4062,N_729);
nand U5911 (N_5911,N_3726,N_1518);
nor U5912 (N_5912,N_3430,N_2500);
nand U5913 (N_5913,N_1263,N_3176);
nor U5914 (N_5914,N_3302,N_4949);
nor U5915 (N_5915,N_3452,N_2325);
or U5916 (N_5916,N_4818,N_817);
or U5917 (N_5917,N_2908,N_863);
or U5918 (N_5918,N_3829,N_265);
nor U5919 (N_5919,N_3441,N_3305);
nand U5920 (N_5920,N_2056,N_3688);
nor U5921 (N_5921,N_2949,N_4265);
nand U5922 (N_5922,N_4167,N_4909);
nor U5923 (N_5923,N_686,N_3346);
or U5924 (N_5924,N_2074,N_4761);
and U5925 (N_5925,N_4922,N_4632);
xnor U5926 (N_5926,N_919,N_132);
nor U5927 (N_5927,N_3978,N_86);
and U5928 (N_5928,N_1048,N_842);
and U5929 (N_5929,N_4711,N_2347);
or U5930 (N_5930,N_925,N_4162);
nand U5931 (N_5931,N_2438,N_2742);
or U5932 (N_5932,N_1905,N_3519);
nand U5933 (N_5933,N_533,N_2429);
nor U5934 (N_5934,N_2411,N_2804);
nand U5935 (N_5935,N_720,N_4592);
and U5936 (N_5936,N_3093,N_149);
and U5937 (N_5937,N_3631,N_2855);
nor U5938 (N_5938,N_1213,N_485);
nor U5939 (N_5939,N_1699,N_3710);
nand U5940 (N_5940,N_2428,N_1889);
nor U5941 (N_5941,N_2071,N_4833);
or U5942 (N_5942,N_2187,N_993);
or U5943 (N_5943,N_424,N_2051);
nor U5944 (N_5944,N_3178,N_45);
nor U5945 (N_5945,N_4466,N_275);
or U5946 (N_5946,N_3292,N_3897);
nor U5947 (N_5947,N_3082,N_2748);
or U5948 (N_5948,N_890,N_2175);
or U5949 (N_5949,N_3094,N_4311);
or U5950 (N_5950,N_3743,N_4126);
and U5951 (N_5951,N_2217,N_244);
or U5952 (N_5952,N_1360,N_1631);
nand U5953 (N_5953,N_2421,N_1547);
nand U5954 (N_5954,N_4273,N_662);
and U5955 (N_5955,N_1990,N_3643);
nor U5956 (N_5956,N_2295,N_208);
nand U5957 (N_5957,N_1585,N_636);
nor U5958 (N_5958,N_3291,N_1154);
nand U5959 (N_5959,N_1332,N_2392);
or U5960 (N_5960,N_1706,N_1691);
nor U5961 (N_5961,N_3598,N_4738);
or U5962 (N_5962,N_3223,N_3813);
and U5963 (N_5963,N_1946,N_1265);
and U5964 (N_5964,N_2620,N_764);
xor U5965 (N_5965,N_3303,N_315);
and U5966 (N_5966,N_1635,N_532);
and U5967 (N_5967,N_1816,N_796);
nand U5968 (N_5968,N_2800,N_3008);
nor U5969 (N_5969,N_2537,N_3764);
or U5970 (N_5970,N_1162,N_2801);
and U5971 (N_5971,N_2666,N_3835);
nor U5972 (N_5972,N_4104,N_4516);
and U5973 (N_5973,N_4098,N_2793);
and U5974 (N_5974,N_4476,N_3969);
xnor U5975 (N_5975,N_3198,N_4355);
nand U5976 (N_5976,N_1455,N_147);
or U5977 (N_5977,N_2254,N_2718);
or U5978 (N_5978,N_4300,N_2534);
or U5979 (N_5979,N_1232,N_1445);
and U5980 (N_5980,N_2063,N_2505);
or U5981 (N_5981,N_3106,N_1112);
xor U5982 (N_5982,N_2853,N_4556);
and U5983 (N_5983,N_2889,N_1954);
nand U5984 (N_5984,N_4421,N_4309);
or U5985 (N_5985,N_4868,N_61);
nand U5986 (N_5986,N_2068,N_4552);
and U5987 (N_5987,N_1084,N_116);
and U5988 (N_5988,N_920,N_3723);
nand U5989 (N_5989,N_430,N_50);
nand U5990 (N_5990,N_143,N_3251);
nand U5991 (N_5991,N_1983,N_155);
nand U5992 (N_5992,N_3609,N_3433);
nand U5993 (N_5993,N_4458,N_516);
and U5994 (N_5994,N_4688,N_813);
and U5995 (N_5995,N_296,N_2543);
or U5996 (N_5996,N_2836,N_2737);
xnor U5997 (N_5997,N_4544,N_4546);
and U5998 (N_5998,N_2759,N_4409);
or U5999 (N_5999,N_3458,N_3536);
nor U6000 (N_6000,N_1527,N_2414);
nand U6001 (N_6001,N_4321,N_2827);
nor U6002 (N_6002,N_923,N_1561);
nand U6003 (N_6003,N_1234,N_2966);
nor U6004 (N_6004,N_4823,N_2341);
nand U6005 (N_6005,N_6,N_1487);
nand U6006 (N_6006,N_2607,N_3160);
nor U6007 (N_6007,N_222,N_1778);
nor U6008 (N_6008,N_2818,N_665);
nor U6009 (N_6009,N_2581,N_2599);
nor U6010 (N_6010,N_2023,N_949);
and U6011 (N_6011,N_4452,N_1783);
and U6012 (N_6012,N_3809,N_1238);
and U6013 (N_6013,N_4280,N_3549);
nor U6014 (N_6014,N_4603,N_3427);
nand U6015 (N_6015,N_3360,N_3810);
and U6016 (N_6016,N_4652,N_1422);
nor U6017 (N_6017,N_4618,N_4553);
and U6018 (N_6018,N_4,N_3642);
nand U6019 (N_6019,N_3412,N_4087);
nand U6020 (N_6020,N_3936,N_1342);
and U6021 (N_6021,N_399,N_1424);
nand U6022 (N_6022,N_1058,N_3488);
and U6023 (N_6023,N_4368,N_433);
and U6024 (N_6024,N_4338,N_3500);
or U6025 (N_6025,N_3355,N_663);
and U6026 (N_6026,N_4925,N_4254);
nand U6027 (N_6027,N_2331,N_3970);
and U6028 (N_6028,N_653,N_3289);
nor U6029 (N_6029,N_1197,N_3402);
or U6030 (N_6030,N_3469,N_2055);
nand U6031 (N_6031,N_1623,N_2601);
nor U6032 (N_6032,N_3268,N_2412);
or U6033 (N_6033,N_3887,N_3974);
nor U6034 (N_6034,N_273,N_4788);
nand U6035 (N_6035,N_209,N_3158);
or U6036 (N_6036,N_3640,N_122);
or U6037 (N_6037,N_3423,N_2713);
and U6038 (N_6038,N_71,N_3938);
and U6039 (N_6039,N_3541,N_4598);
or U6040 (N_6040,N_687,N_240);
nand U6041 (N_6041,N_2103,N_322);
nand U6042 (N_6042,N_1313,N_2508);
nor U6043 (N_6043,N_4484,N_1589);
nand U6044 (N_6044,N_1880,N_1595);
nand U6045 (N_6045,N_2971,N_2302);
or U6046 (N_6046,N_3972,N_2639);
nor U6047 (N_6047,N_586,N_3366);
nor U6048 (N_6048,N_1618,N_4085);
nand U6049 (N_6049,N_1395,N_4000);
and U6050 (N_6050,N_4157,N_4931);
nand U6051 (N_6051,N_2214,N_2751);
and U6052 (N_6052,N_4442,N_1571);
xor U6053 (N_6053,N_2211,N_3811);
or U6054 (N_6054,N_4678,N_3380);
nor U6055 (N_6055,N_1398,N_1642);
and U6056 (N_6056,N_4953,N_3348);
nor U6057 (N_6057,N_502,N_2828);
or U6058 (N_6058,N_4065,N_4816);
nor U6059 (N_6059,N_255,N_2852);
and U6060 (N_6060,N_2440,N_2961);
xnor U6061 (N_6061,N_3229,N_2444);
nand U6062 (N_6062,N_2109,N_1726);
nand U6063 (N_6063,N_3749,N_3626);
nand U6064 (N_6064,N_524,N_4312);
nand U6065 (N_6065,N_2492,N_784);
nand U6066 (N_6066,N_2854,N_2348);
nor U6067 (N_6067,N_4076,N_18);
nor U6068 (N_6068,N_1831,N_1379);
nor U6069 (N_6069,N_3573,N_1186);
and U6070 (N_6070,N_684,N_2146);
xor U6071 (N_6071,N_347,N_2391);
and U6072 (N_6072,N_2882,N_2519);
and U6073 (N_6073,N_1247,N_1425);
or U6074 (N_6074,N_3827,N_2515);
or U6075 (N_6075,N_2847,N_3603);
and U6076 (N_6076,N_4541,N_1345);
and U6077 (N_6077,N_2457,N_3038);
and U6078 (N_6078,N_1149,N_1259);
nand U6079 (N_6079,N_2638,N_3306);
or U6080 (N_6080,N_472,N_886);
nand U6081 (N_6081,N_1823,N_1897);
and U6082 (N_6082,N_4041,N_2061);
nand U6083 (N_6083,N_58,N_1309);
nand U6084 (N_6084,N_2770,N_2582);
and U6085 (N_6085,N_2208,N_4686);
nand U6086 (N_6086,N_563,N_2541);
nor U6087 (N_6087,N_1437,N_807);
and U6088 (N_6088,N_4224,N_1272);
nor U6089 (N_6089,N_2561,N_4775);
or U6090 (N_6090,N_1115,N_4214);
xor U6091 (N_6091,N_4923,N_2378);
nand U6092 (N_6092,N_629,N_125);
and U6093 (N_6093,N_676,N_3507);
and U6094 (N_6094,N_3205,N_4872);
and U6095 (N_6095,N_2183,N_4769);
or U6096 (N_6096,N_1121,N_3903);
or U6097 (N_6097,N_1441,N_549);
and U6098 (N_6098,N_1812,N_2614);
nand U6099 (N_6099,N_168,N_2393);
or U6100 (N_6100,N_4917,N_1396);
nor U6101 (N_6101,N_2172,N_1837);
nand U6102 (N_6102,N_457,N_4654);
nor U6103 (N_6103,N_4804,N_263);
nand U6104 (N_6104,N_1132,N_2293);
nor U6105 (N_6105,N_4864,N_4378);
nand U6106 (N_6106,N_4944,N_4147);
nand U6107 (N_6107,N_1494,N_3945);
nor U6108 (N_6108,N_3651,N_3378);
nor U6109 (N_6109,N_4700,N_2025);
or U6110 (N_6110,N_4490,N_1128);
nor U6111 (N_6111,N_2398,N_1757);
nor U6112 (N_6112,N_774,N_2838);
nor U6113 (N_6113,N_3789,N_4888);
nand U6114 (N_6114,N_78,N_3066);
nor U6115 (N_6115,N_2383,N_3714);
nor U6116 (N_6116,N_1226,N_225);
or U6117 (N_6117,N_4424,N_1325);
nor U6118 (N_6118,N_3823,N_2483);
or U6119 (N_6119,N_2711,N_1529);
and U6120 (N_6120,N_4156,N_2242);
nand U6121 (N_6121,N_2088,N_931);
nor U6122 (N_6122,N_2322,N_2894);
and U6123 (N_6123,N_1118,N_4498);
nand U6124 (N_6124,N_3031,N_120);
nor U6125 (N_6125,N_1649,N_3356);
nand U6126 (N_6126,N_1031,N_402);
and U6127 (N_6127,N_987,N_2822);
nand U6128 (N_6128,N_1610,N_1079);
or U6129 (N_6129,N_716,N_1591);
and U6130 (N_6130,N_2234,N_3457);
or U6131 (N_6131,N_3731,N_2580);
nor U6132 (N_6132,N_4108,N_1674);
xnor U6133 (N_6133,N_1989,N_2610);
and U6134 (N_6134,N_4875,N_28);
nand U6135 (N_6135,N_1018,N_2143);
nor U6136 (N_6136,N_548,N_3895);
and U6137 (N_6137,N_4999,N_2831);
nand U6138 (N_6138,N_4382,N_346);
nor U6139 (N_6139,N_121,N_190);
or U6140 (N_6140,N_4894,N_3948);
or U6141 (N_6141,N_869,N_4570);
and U6142 (N_6142,N_313,N_3657);
nand U6143 (N_6143,N_185,N_2756);
nor U6144 (N_6144,N_4365,N_2494);
or U6145 (N_6145,N_1279,N_4717);
or U6146 (N_6146,N_3739,N_2970);
or U6147 (N_6147,N_3595,N_8);
or U6148 (N_6148,N_3900,N_3681);
nor U6149 (N_6149,N_1393,N_2746);
nand U6150 (N_6150,N_4425,N_4079);
and U6151 (N_6151,N_396,N_3362);
nor U6152 (N_6152,N_2013,N_55);
and U6153 (N_6153,N_4533,N_187);
nand U6154 (N_6154,N_4926,N_4841);
nand U6155 (N_6155,N_2127,N_4327);
or U6156 (N_6156,N_2951,N_3769);
and U6157 (N_6157,N_3301,N_4573);
or U6158 (N_6158,N_2556,N_1144);
and U6159 (N_6159,N_3129,N_2608);
nor U6160 (N_6160,N_1940,N_1731);
nor U6161 (N_6161,N_2475,N_4334);
nand U6162 (N_6162,N_3314,N_3703);
nor U6163 (N_6163,N_1107,N_3546);
and U6164 (N_6164,N_3812,N_3446);
nand U6165 (N_6165,N_2634,N_251);
nand U6166 (N_6166,N_2551,N_408);
nand U6167 (N_6167,N_3480,N_3088);
nand U6168 (N_6168,N_2474,N_593);
nand U6169 (N_6169,N_3690,N_3975);
and U6170 (N_6170,N_1617,N_1049);
nand U6171 (N_6171,N_1328,N_2725);
nor U6172 (N_6172,N_4799,N_276);
nor U6173 (N_6173,N_4848,N_2942);
and U6174 (N_6174,N_1567,N_1793);
nor U6175 (N_6175,N_4335,N_1025);
nor U6176 (N_6176,N_395,N_233);
or U6177 (N_6177,N_3971,N_608);
nor U6178 (N_6178,N_1236,N_1555);
or U6179 (N_6179,N_180,N_3581);
and U6180 (N_6180,N_844,N_2943);
nor U6181 (N_6181,N_967,N_2419);
nor U6182 (N_6182,N_4013,N_1794);
nand U6183 (N_6183,N_324,N_4497);
nand U6184 (N_6184,N_3667,N_962);
or U6185 (N_6185,N_4994,N_4123);
or U6186 (N_6186,N_4697,N_2919);
and U6187 (N_6187,N_123,N_798);
or U6188 (N_6188,N_2945,N_1394);
and U6189 (N_6189,N_853,N_1662);
nand U6190 (N_6190,N_1298,N_4763);
nand U6191 (N_6191,N_3845,N_1842);
and U6192 (N_6192,N_2686,N_1776);
nand U6193 (N_6193,N_3287,N_2569);
nand U6194 (N_6194,N_4874,N_2229);
or U6195 (N_6195,N_3219,N_3189);
nand U6196 (N_6196,N_2651,N_3585);
nor U6197 (N_6197,N_4292,N_4892);
or U6198 (N_6198,N_4812,N_1841);
nand U6199 (N_6199,N_4554,N_2901);
nor U6200 (N_6200,N_3820,N_2699);
and U6201 (N_6201,N_667,N_4111);
and U6202 (N_6202,N_498,N_3010);
or U6203 (N_6203,N_3552,N_301);
nor U6204 (N_6204,N_3357,N_985);
and U6205 (N_6205,N_627,N_2503);
and U6206 (N_6206,N_3725,N_2925);
and U6207 (N_6207,N_4810,N_1919);
and U6208 (N_6208,N_3182,N_1927);
and U6209 (N_6209,N_2290,N_4036);
xor U6210 (N_6210,N_2977,N_4689);
and U6211 (N_6211,N_602,N_3980);
and U6212 (N_6212,N_2250,N_1777);
nand U6213 (N_6213,N_1973,N_691);
and U6214 (N_6214,N_459,N_4687);
nand U6215 (N_6215,N_299,N_2330);
nand U6216 (N_6216,N_4891,N_4616);
or U6217 (N_6217,N_1233,N_4236);
nand U6218 (N_6218,N_1735,N_3757);
and U6219 (N_6219,N_154,N_134);
nand U6220 (N_6220,N_1882,N_2886);
and U6221 (N_6221,N_1910,N_1613);
nand U6222 (N_6222,N_3024,N_3487);
nor U6223 (N_6223,N_2820,N_1911);
nand U6224 (N_6224,N_3005,N_283);
nand U6225 (N_6225,N_4773,N_201);
xnor U6226 (N_6226,N_4740,N_937);
and U6227 (N_6227,N_94,N_3956);
or U6228 (N_6228,N_3685,N_2817);
and U6229 (N_6229,N_4736,N_2994);
nor U6230 (N_6230,N_226,N_4634);
and U6231 (N_6231,N_537,N_4794);
nand U6232 (N_6232,N_802,N_2389);
or U6233 (N_6233,N_1056,N_234);
or U6234 (N_6234,N_2795,N_580);
or U6235 (N_6235,N_153,N_971);
nand U6236 (N_6236,N_2125,N_195);
nand U6237 (N_6237,N_589,N_3085);
or U6238 (N_6238,N_3526,N_1586);
nor U6239 (N_6239,N_3456,N_4617);
nor U6240 (N_6240,N_2451,N_1883);
nand U6241 (N_6241,N_2611,N_3206);
or U6242 (N_6242,N_859,N_439);
nor U6243 (N_6243,N_1827,N_867);
nand U6244 (N_6244,N_1596,N_1815);
and U6245 (N_6245,N_4326,N_661);
nand U6246 (N_6246,N_590,N_4207);
or U6247 (N_6247,N_1219,N_2773);
nand U6248 (N_6248,N_793,N_2791);
nand U6249 (N_6249,N_4216,N_438);
or U6250 (N_6250,N_4396,N_448);
or U6251 (N_6251,N_4446,N_2213);
or U6252 (N_6252,N_1924,N_1551);
nand U6253 (N_6253,N_0,N_3672);
nand U6254 (N_6254,N_2168,N_4558);
or U6255 (N_6255,N_4176,N_1562);
nor U6256 (N_6256,N_4997,N_1218);
nand U6257 (N_6257,N_3785,N_1355);
or U6258 (N_6258,N_2602,N_48);
nand U6259 (N_6259,N_245,N_740);
nor U6260 (N_6260,N_3891,N_1297);
nand U6261 (N_6261,N_3493,N_1041);
and U6262 (N_6262,N_4530,N_778);
or U6263 (N_6263,N_1177,N_3190);
nor U6264 (N_6264,N_2693,N_2918);
or U6265 (N_6265,N_3467,N_2227);
xor U6266 (N_6266,N_493,N_3693);
nor U6267 (N_6267,N_1314,N_4420);
and U6268 (N_6268,N_713,N_4008);
xor U6269 (N_6269,N_2850,N_2907);
nand U6270 (N_6270,N_4613,N_1378);
nor U6271 (N_6271,N_309,N_1349);
nor U6272 (N_6272,N_2710,N_3407);
and U6273 (N_6273,N_647,N_1306);
or U6274 (N_6274,N_471,N_3354);
nand U6275 (N_6275,N_824,N_1979);
and U6276 (N_6276,N_4082,N_1969);
and U6277 (N_6277,N_1251,N_2032);
nor U6278 (N_6278,N_2549,N_1828);
or U6279 (N_6279,N_2559,N_4795);
and U6280 (N_6280,N_630,N_76);
xor U6281 (N_6281,N_3460,N_2219);
and U6282 (N_6282,N_3227,N_3804);
or U6283 (N_6283,N_25,N_749);
or U6284 (N_6284,N_279,N_4359);
nor U6285 (N_6285,N_4144,N_540);
and U6286 (N_6286,N_2733,N_1491);
nor U6287 (N_6287,N_1784,N_3692);
and U6288 (N_6288,N_1435,N_2807);
or U6289 (N_6289,N_1553,N_2766);
or U6290 (N_6290,N_2482,N_1521);
or U6291 (N_6291,N_4033,N_42);
or U6292 (N_6292,N_2291,N_2815);
or U6293 (N_6293,N_4293,N_2764);
or U6294 (N_6294,N_137,N_14);
nand U6295 (N_6295,N_3320,N_3445);
nor U6296 (N_6296,N_401,N_640);
or U6297 (N_6297,N_4354,N_4581);
xnor U6298 (N_6298,N_761,N_2900);
and U6299 (N_6299,N_3992,N_3525);
nand U6300 (N_6300,N_634,N_606);
or U6301 (N_6301,N_782,N_2867);
or U6302 (N_6302,N_3272,N_3808);
nor U6303 (N_6303,N_4995,N_1135);
and U6304 (N_6304,N_4264,N_1807);
and U6305 (N_6305,N_3935,N_685);
nor U6306 (N_6306,N_1516,N_3828);
or U6307 (N_6307,N_1464,N_1273);
nand U6308 (N_6308,N_2335,N_2174);
and U6309 (N_6309,N_4068,N_2805);
nor U6310 (N_6310,N_1587,N_2157);
xnor U6311 (N_6311,N_893,N_2369);
nand U6312 (N_6312,N_1072,N_2079);
nand U6313 (N_6313,N_1968,N_3994);
or U6314 (N_6314,N_527,N_1693);
nor U6315 (N_6315,N_4600,N_4134);
nand U6316 (N_6316,N_628,N_3821);
nand U6317 (N_6317,N_1856,N_3521);
or U6318 (N_6318,N_951,N_4240);
or U6319 (N_6319,N_1893,N_3011);
nand U6320 (N_6320,N_2430,N_4491);
nand U6321 (N_6321,N_2723,N_1544);
nand U6322 (N_6322,N_3856,N_4341);
or U6323 (N_6323,N_2623,N_1755);
and U6324 (N_6324,N_3963,N_2612);
nor U6325 (N_6325,N_327,N_1752);
or U6326 (N_6326,N_787,N_2682);
and U6327 (N_6327,N_3293,N_4591);
nor U6328 (N_6328,N_1369,N_4330);
nand U6329 (N_6329,N_4673,N_475);
and U6330 (N_6330,N_3504,N_2579);
and U6331 (N_6331,N_3426,N_4665);
and U6332 (N_6332,N_2312,N_2427);
nand U6333 (N_6333,N_3737,N_3572);
or U6334 (N_6334,N_1874,N_4394);
nor U6335 (N_6335,N_4205,N_862);
nor U6336 (N_6336,N_3409,N_4067);
and U6337 (N_6337,N_4660,N_1987);
nor U6338 (N_6338,N_462,N_3179);
nand U6339 (N_6339,N_1663,N_3768);
nor U6340 (N_6340,N_2902,N_1327);
nand U6341 (N_6341,N_3766,N_1093);
nand U6342 (N_6342,N_878,N_3015);
xnor U6343 (N_6343,N_3047,N_2594);
or U6344 (N_6344,N_2147,N_4455);
nand U6345 (N_6345,N_1680,N_1101);
or U6346 (N_6346,N_2352,N_4318);
nand U6347 (N_6347,N_719,N_683);
or U6348 (N_6348,N_1095,N_4834);
and U6349 (N_6349,N_2833,N_3387);
nand U6350 (N_6350,N_3078,N_2848);
and U6351 (N_6351,N_3638,N_1941);
or U6352 (N_6352,N_2884,N_1791);
nand U6353 (N_6353,N_108,N_1262);
or U6354 (N_6354,N_986,N_4237);
or U6355 (N_6355,N_2890,N_2256);
nand U6356 (N_6356,N_4612,N_4896);
nor U6357 (N_6357,N_2562,N_4908);
nand U6358 (N_6358,N_515,N_4252);
nand U6359 (N_6359,N_2300,N_354);
or U6360 (N_6360,N_573,N_4764);
nand U6361 (N_6361,N_3647,N_2525);
nand U6362 (N_6362,N_3600,N_1903);
or U6363 (N_6363,N_3989,N_1881);
nand U6364 (N_6364,N_4867,N_141);
or U6365 (N_6365,N_413,N_3576);
and U6366 (N_6366,N_3428,N_1321);
nand U6367 (N_6367,N_2905,N_3404);
nor U6368 (N_6368,N_2489,N_3053);
and U6369 (N_6369,N_644,N_1520);
or U6370 (N_6370,N_2296,N_2386);
and U6371 (N_6371,N_1440,N_2934);
nand U6372 (N_6372,N_3919,N_2282);
nand U6373 (N_6373,N_3502,N_3376);
nor U6374 (N_6374,N_202,N_695);
or U6375 (N_6375,N_755,N_3304);
nand U6376 (N_6376,N_4720,N_3675);
and U6377 (N_6377,N_3244,N_3770);
or U6378 (N_6378,N_690,N_4356);
nand U6379 (N_6379,N_3345,N_928);
and U6380 (N_6380,N_3489,N_566);
nand U6381 (N_6381,N_1223,N_2780);
or U6382 (N_6382,N_1390,N_1094);
xor U6383 (N_6383,N_1330,N_4710);
and U6384 (N_6384,N_20,N_2415);
nor U6385 (N_6385,N_152,N_1228);
nand U6386 (N_6386,N_2228,N_981);
nor U6387 (N_6387,N_4709,N_3732);
and U6388 (N_6388,N_727,N_943);
nand U6389 (N_6389,N_2465,N_4043);
or U6390 (N_6390,N_583,N_2586);
nand U6391 (N_6391,N_4035,N_4171);
nor U6392 (N_6392,N_756,N_4714);
and U6393 (N_6393,N_3554,N_2019);
and U6394 (N_6394,N_3786,N_394);
or U6395 (N_6395,N_4986,N_184);
and U6396 (N_6396,N_288,N_874);
nor U6397 (N_6397,N_3719,N_1271);
and U6398 (N_6398,N_2091,N_4651);
and U6399 (N_6399,N_601,N_2180);
or U6400 (N_6400,N_584,N_1514);
or U6401 (N_6401,N_4315,N_3977);
and U6402 (N_6402,N_2404,N_236);
nand U6403 (N_6403,N_651,N_3863);
and U6404 (N_6404,N_243,N_4138);
nand U6405 (N_6405,N_2844,N_3775);
and U6406 (N_6406,N_2913,N_2509);
or U6407 (N_6407,N_934,N_316);
nor U6408 (N_6408,N_3275,N_535);
and U6409 (N_6409,N_46,N_4966);
and U6410 (N_6410,N_3270,N_4734);
or U6411 (N_6411,N_2191,N_24);
nor U6412 (N_6412,N_429,N_1169);
and U6413 (N_6413,N_2619,N_4913);
and U6414 (N_6414,N_1442,N_4829);
and U6415 (N_6415,N_1568,N_2708);
and U6416 (N_6416,N_3490,N_2891);
and U6417 (N_6417,N_4393,N_2539);
or U6418 (N_6418,N_1065,N_2552);
nand U6419 (N_6419,N_2883,N_4930);
or U6420 (N_6420,N_3230,N_451);
xnor U6421 (N_6421,N_1243,N_4210);
nor U6422 (N_6422,N_1068,N_4215);
or U6423 (N_6423,N_3207,N_992);
or U6424 (N_6424,N_4806,N_454);
and U6425 (N_6425,N_473,N_3759);
and U6426 (N_6426,N_3671,N_2251);
nand U6427 (N_6427,N_762,N_4445);
nor U6428 (N_6428,N_4011,N_3494);
nand U6429 (N_6429,N_3797,N_172);
or U6430 (N_6430,N_709,N_2857);
nand U6431 (N_6431,N_4247,N_2606);
nor U6432 (N_6432,N_2390,N_350);
nor U6433 (N_6433,N_2978,N_1082);
and U6434 (N_6434,N_2192,N_2932);
nor U6435 (N_6435,N_411,N_2413);
nor U6436 (N_6436,N_188,N_4155);
and U6437 (N_6437,N_3068,N_3290);
nor U6438 (N_6438,N_1021,N_670);
nand U6439 (N_6439,N_1017,N_2318);
nor U6440 (N_6440,N_2873,N_2625);
nor U6441 (N_6441,N_1566,N_2363);
and U6442 (N_6442,N_733,N_207);
nor U6443 (N_6443,N_383,N_3534);
xor U6444 (N_6444,N_4835,N_326);
or U6445 (N_6445,N_3589,N_328);
nor U6446 (N_6446,N_3211,N_3910);
or U6447 (N_6447,N_1054,N_3568);
nand U6448 (N_6448,N_2878,N_2700);
and U6449 (N_6449,N_1276,N_1374);
nand U6450 (N_6450,N_1864,N_3146);
or U6451 (N_6451,N_974,N_464);
and U6452 (N_6452,N_4535,N_3405);
or U6453 (N_6453,N_1409,N_4973);
nor U6454 (N_6454,N_3708,N_2959);
and U6455 (N_6455,N_2220,N_4921);
and U6456 (N_6456,N_896,N_2514);
nand U6457 (N_6457,N_4900,N_1131);
or U6458 (N_6458,N_374,N_1948);
or U6459 (N_6459,N_3060,N_990);
or U6460 (N_6460,N_3801,N_1308);
or U6461 (N_6461,N_3851,N_964);
nor U6462 (N_6462,N_897,N_4881);
or U6463 (N_6463,N_84,N_1694);
or U6464 (N_6464,N_972,N_1477);
nor U6465 (N_6465,N_1322,N_871);
xor U6466 (N_6466,N_979,N_1936);
or U6467 (N_6467,N_1692,N_2615);
and U6468 (N_6468,N_1713,N_4787);
nand U6469 (N_6469,N_419,N_4239);
nand U6470 (N_6470,N_164,N_4658);
nor U6471 (N_6471,N_4739,N_4399);
or U6472 (N_6472,N_2093,N_3484);
or U6473 (N_6473,N_512,N_2464);
nand U6474 (N_6474,N_2096,N_3673);
nor U6475 (N_6475,N_4152,N_3163);
and U6476 (N_6476,N_217,N_4815);
and U6477 (N_6477,N_1161,N_1600);
nor U6478 (N_6478,N_2339,N_4887);
or U6479 (N_6479,N_2984,N_2778);
nand U6480 (N_6480,N_4602,N_3353);
nand U6481 (N_6481,N_4428,N_1814);
and U6482 (N_6482,N_2895,N_1921);
nor U6483 (N_6483,N_2077,N_114);
or U6484 (N_6484,N_2292,N_4377);
nand U6485 (N_6485,N_3041,N_689);
or U6486 (N_6486,N_4302,N_3512);
or U6487 (N_6487,N_3260,N_2496);
nor U6488 (N_6488,N_3611,N_4849);
and U6489 (N_6489,N_1485,N_171);
or U6490 (N_6490,N_4072,N_2911);
nand U6491 (N_6491,N_3188,N_3885);
or U6492 (N_6492,N_814,N_1130);
nand U6493 (N_6493,N_1352,N_4051);
nand U6494 (N_6494,N_2232,N_4899);
or U6495 (N_6495,N_166,N_1359);
and U6496 (N_6496,N_264,N_4005);
and U6497 (N_6497,N_1772,N_1820);
nand U6498 (N_6498,N_2104,N_3130);
nand U6499 (N_6499,N_2753,N_2974);
or U6500 (N_6500,N_1792,N_3904);
and U6501 (N_6501,N_4012,N_1013);
or U6502 (N_6502,N_2021,N_1221);
and U6503 (N_6503,N_1537,N_3369);
or U6504 (N_6504,N_367,N_79);
or U6505 (N_6505,N_2553,N_954);
xor U6506 (N_6506,N_1008,N_4622);
or U6507 (N_6507,N_3582,N_2395);
and U6508 (N_6508,N_336,N_452);
nor U6509 (N_6509,N_3148,N_4006);
nand U6510 (N_6510,N_4483,N_3166);
nand U6511 (N_6511,N_4778,N_4539);
or U6512 (N_6512,N_4200,N_247);
nand U6513 (N_6513,N_1986,N_1715);
or U6514 (N_6514,N_4345,N_1702);
nor U6515 (N_6515,N_2301,N_3870);
and U6516 (N_6516,N_2931,N_4979);
nor U6517 (N_6517,N_4519,N_752);
or U6518 (N_6518,N_4620,N_3126);
and U6519 (N_6519,N_3884,N_4767);
nand U6520 (N_6520,N_4487,N_3738);
nor U6521 (N_6521,N_2924,N_1389);
nor U6522 (N_6522,N_3061,N_2595);
and U6523 (N_6523,N_1996,N_2082);
nor U6524 (N_6524,N_4955,N_1071);
or U6525 (N_6525,N_3634,N_4903);
xnor U6526 (N_6526,N_522,N_939);
or U6527 (N_6527,N_3601,N_1171);
nor U6528 (N_6528,N_788,N_1450);
xnor U6529 (N_6529,N_2948,N_4275);
or U6530 (N_6530,N_4636,N_3386);
and U6531 (N_6531,N_881,N_4233);
nor U6532 (N_6532,N_3099,N_3271);
nand U6533 (N_6533,N_4077,N_1826);
and U6534 (N_6534,N_97,N_2842);
or U6535 (N_6535,N_297,N_1420);
and U6536 (N_6536,N_1727,N_1088);
and U6537 (N_6537,N_2439,N_3960);
and U6538 (N_6538,N_1208,N_4430);
xnor U6539 (N_6539,N_2705,N_3715);
or U6540 (N_6540,N_2650,N_4674);
and U6541 (N_6541,N_3417,N_1052);
nand U6542 (N_6542,N_3461,N_3854);
and U6543 (N_6543,N_2059,N_1133);
or U6544 (N_6544,N_1334,N_3967);
nand U6545 (N_6545,N_4844,N_1244);
or U6546 (N_6546,N_1106,N_3867);
nand U6547 (N_6547,N_4135,N_496);
or U6548 (N_6548,N_579,N_513);
and U6549 (N_6549,N_4165,N_3334);
nor U6550 (N_6550,N_3561,N_2513);
nor U6551 (N_6551,N_1209,N_2546);
and U6552 (N_6552,N_1231,N_2052);
and U6553 (N_6553,N_4383,N_3325);
nand U6554 (N_6554,N_2958,N_1974);
or U6555 (N_6555,N_1955,N_1665);
or U6556 (N_6556,N_866,N_1211);
nor U6557 (N_6557,N_1299,N_2381);
nor U6558 (N_6558,N_4869,N_547);
and U6559 (N_6559,N_2156,N_4499);
nand U6560 (N_6560,N_973,N_3560);
nor U6561 (N_6561,N_2626,N_4877);
nand U6562 (N_6562,N_715,N_3916);
nand U6563 (N_6563,N_2738,N_3746);
nand U6564 (N_6564,N_3877,N_3210);
or U6565 (N_6565,N_2664,N_4474);
or U6566 (N_6566,N_2014,N_129);
or U6567 (N_6567,N_1388,N_1311);
nor U6568 (N_6568,N_1373,N_1270);
or U6569 (N_6569,N_530,N_2015);
or U6570 (N_6570,N_2000,N_3990);
nor U6571 (N_6571,N_146,N_426);
and U6572 (N_6572,N_1743,N_2364);
and U6573 (N_6573,N_4492,N_4501);
or U6574 (N_6574,N_3842,N_1191);
nor U6575 (N_6575,N_3486,N_845);
nand U6576 (N_6576,N_571,N_4712);
nor U6577 (N_6577,N_1961,N_3453);
nor U6578 (N_6578,N_3742,N_1429);
nand U6579 (N_6579,N_4621,N_497);
or U6580 (N_6580,N_3518,N_308);
or U6581 (N_6581,N_3476,N_1245);
nand U6582 (N_6582,N_4496,N_4406);
nand U6583 (N_6583,N_4469,N_3114);
xnor U6584 (N_6584,N_3464,N_697);
and U6585 (N_6585,N_1711,N_2507);
nor U6586 (N_6586,N_3876,N_4279);
or U6587 (N_6587,N_2745,N_2732);
nor U6588 (N_6588,N_1846,N_3222);
or U6589 (N_6589,N_1855,N_625);
nor U6590 (N_6590,N_3556,N_334);
nor U6591 (N_6591,N_1029,N_2196);
or U6592 (N_6592,N_4001,N_744);
nor U6593 (N_6593,N_4261,N_2999);
and U6594 (N_6594,N_1533,N_381);
or U6595 (N_6595,N_4109,N_4655);
nand U6596 (N_6596,N_2670,N_3805);
or U6597 (N_6597,N_478,N_3197);
and U6598 (N_6598,N_633,N_1096);
xor U6599 (N_6599,N_4518,N_3499);
and U6600 (N_6600,N_2001,N_3064);
and U6601 (N_6601,N_577,N_3961);
nor U6602 (N_6602,N_3029,N_1178);
nor U6603 (N_6603,N_837,N_3336);
nand U6604 (N_6604,N_363,N_1690);
nor U6605 (N_6605,N_2246,N_7);
nor U6606 (N_6606,N_2596,N_3169);
or U6607 (N_6607,N_4950,N_460);
nand U6608 (N_6608,N_4631,N_3505);
nor U6609 (N_6609,N_66,N_525);
nand U6610 (N_6610,N_1483,N_2304);
nand U6611 (N_6611,N_4096,N_1803);
nor U6612 (N_6612,N_3396,N_3);
or U6613 (N_6613,N_1312,N_4830);
and U6614 (N_6614,N_1958,N_2375);
nand U6615 (N_6615,N_4608,N_1172);
nand U6616 (N_6616,N_2669,N_3931);
xnor U6617 (N_6617,N_3646,N_3191);
and U6618 (N_6618,N_792,N_2230);
nor U6619 (N_6619,N_1200,N_2849);
or U6620 (N_6620,N_728,N_2497);
nor U6621 (N_6621,N_1492,N_246);
nand U6622 (N_6622,N_4398,N_4566);
nor U6623 (N_6623,N_3120,N_2647);
or U6624 (N_6624,N_117,N_3882);
and U6625 (N_6625,N_4351,N_4493);
nand U6626 (N_6626,N_1668,N_3777);
nor U6627 (N_6627,N_600,N_677);
and U6628 (N_6628,N_3890,N_2264);
or U6629 (N_6629,N_3263,N_3878);
or U6630 (N_6630,N_77,N_1771);
nor U6631 (N_6631,N_2144,N_295);
nor U6632 (N_6632,N_545,N_3716);
or U6633 (N_6633,N_4653,N_2566);
or U6634 (N_6634,N_4436,N_3331);
nor U6635 (N_6635,N_189,N_771);
nor U6636 (N_6636,N_1187,N_4633);
and U6637 (N_6637,N_2271,N_441);
nand U6638 (N_6638,N_3669,N_2641);
nor U6639 (N_6639,N_1619,N_17);
nor U6640 (N_6640,N_534,N_1688);
and U6641 (N_6641,N_186,N_3623);
nand U6642 (N_6642,N_1972,N_2936);
or U6643 (N_6643,N_4402,N_4647);
nor U6644 (N_6644,N_4610,N_337);
and U6645 (N_6645,N_1006,N_242);
nand U6646 (N_6646,N_4083,N_4117);
and U6647 (N_6647,N_2677,N_1994);
nor U6648 (N_6648,N_1945,N_390);
nand U6649 (N_6649,N_2426,N_4182);
and U6650 (N_6650,N_1739,N_4650);
nor U6651 (N_6651,N_4173,N_443);
nor U6652 (N_6652,N_2132,N_558);
nor U6653 (N_6653,N_4371,N_2033);
or U6654 (N_6654,N_1926,N_4238);
or U6655 (N_6655,N_1014,N_3335);
or U6656 (N_6656,N_4467,N_682);
nand U6657 (N_6657,N_1484,N_3668);
nor U6658 (N_6658,N_3050,N_1775);
nor U6659 (N_6659,N_4985,N_1493);
and U6660 (N_6660,N_2962,N_819);
nor U6661 (N_6661,N_1543,N_260);
and U6662 (N_6662,N_1709,N_3034);
and U6663 (N_6663,N_183,N_1869);
or U6664 (N_6664,N_378,N_1217);
nand U6665 (N_6665,N_2286,N_3274);
nand U6666 (N_6666,N_2379,N_3258);
or U6667 (N_6667,N_4928,N_2138);
nand U6668 (N_6668,N_1155,N_1050);
nor U6669 (N_6669,N_2043,N_133);
and U6670 (N_6670,N_1997,N_567);
nand U6671 (N_6671,N_1624,N_3243);
and U6672 (N_6672,N_2653,N_4063);
nor U6673 (N_6673,N_1418,N_526);
and U6674 (N_6674,N_3943,N_2568);
xor U6675 (N_6675,N_2303,N_458);
or U6676 (N_6676,N_2201,N_2645);
xor U6677 (N_6677,N_3394,N_323);
and U6678 (N_6678,N_2081,N_3084);
nor U6679 (N_6679,N_3372,N_34);
and U6680 (N_6680,N_696,N_2072);
and U6681 (N_6681,N_1010,N_487);
nand U6682 (N_6682,N_746,N_3727);
nand U6683 (N_6683,N_4019,N_1766);
or U6684 (N_6684,N_3920,N_3277);
or U6685 (N_6685,N_2698,N_2802);
nand U6686 (N_6686,N_2042,N_3139);
nor U6687 (N_6687,N_2469,N_1590);
or U6688 (N_6688,N_1799,N_3741);
nand U6689 (N_6689,N_1839,N_578);
nor U6690 (N_6690,N_1525,N_1269);
nor U6691 (N_6691,N_2297,N_2477);
or U6692 (N_6692,N_4073,N_2026);
nand U6693 (N_6693,N_3220,N_456);
or U6694 (N_6694,N_307,N_2598);
or U6695 (N_6695,N_3592,N_4259);
nand U6696 (N_6696,N_4596,N_700);
nand U6697 (N_6697,N_3416,N_213);
or U6698 (N_6698,N_239,N_3615);
xnor U6699 (N_6699,N_4873,N_382);
or U6700 (N_6700,N_3470,N_3704);
and U6701 (N_6701,N_317,N_743);
xnor U6702 (N_6702,N_2466,N_4057);
nand U6703 (N_6703,N_4679,N_3677);
nor U6704 (N_6704,N_2786,N_4762);
and U6705 (N_6705,N_3054,N_4161);
nand U6706 (N_6706,N_655,N_2073);
or U6707 (N_6707,N_3252,N_2806);
or U6708 (N_6708,N_940,N_1148);
and U6709 (N_6709,N_1539,N_557);
or U6710 (N_6710,N_2436,N_4595);
nand U6711 (N_6711,N_3873,N_926);
or U6712 (N_6712,N_712,N_4038);
and U6713 (N_6713,N_2952,N_3838);
nand U6714 (N_6714,N_428,N_2460);
or U6715 (N_6715,N_737,N_360);
nor U6716 (N_6716,N_865,N_2991);
nor U6717 (N_6717,N_3670,N_3875);
or U6718 (N_6718,N_4514,N_1194);
and U6719 (N_6719,N_553,N_362);
and U6720 (N_6720,N_3765,N_4159);
nor U6721 (N_6721,N_3100,N_922);
or U6722 (N_6722,N_4190,N_4534);
nor U6723 (N_6723,N_4780,N_3740);
nand U6724 (N_6724,N_3164,N_3822);
and U6725 (N_6725,N_3001,N_1867);
and U6726 (N_6726,N_4278,N_598);
nor U6727 (N_6727,N_468,N_2198);
nand U6728 (N_6728,N_4106,N_2735);
nand U6729 (N_6729,N_4225,N_4870);
nand U6730 (N_6730,N_2506,N_338);
nand U6731 (N_6731,N_3151,N_1302);
nand U6732 (N_6732,N_4640,N_1475);
or U6733 (N_6733,N_4021,N_4569);
and U6734 (N_6734,N_1876,N_678);
nor U6735 (N_6735,N_4277,N_4836);
and U6736 (N_6736,N_4819,N_3896);
nand U6737 (N_6737,N_544,N_4624);
nand U6738 (N_6738,N_1433,N_1656);
xor U6739 (N_6739,N_2523,N_366);
nor U6740 (N_6740,N_999,N_340);
and U6741 (N_6741,N_230,N_2938);
nor U6742 (N_6742,N_4707,N_4644);
or U6743 (N_6743,N_1574,N_834);
nand U6744 (N_6744,N_2858,N_4017);
or U6745 (N_6745,N_4145,N_3906);
nand U6746 (N_6746,N_4984,N_2209);
and U6747 (N_6747,N_1407,N_1873);
xnor U6748 (N_6748,N_2856,N_839);
nand U6749 (N_6749,N_436,N_4276);
and U6750 (N_6750,N_3288,N_3782);
and U6751 (N_6751,N_3824,N_32);
xor U6752 (N_6752,N_1560,N_4802);
nand U6753 (N_6753,N_483,N_4662);
xnor U6754 (N_6754,N_1898,N_2121);
or U6755 (N_6755,N_1040,N_820);
or U6756 (N_6756,N_215,N_2224);
and U6757 (N_6757,N_3745,N_2004);
or U6758 (N_6758,N_887,N_2255);
nand U6759 (N_6759,N_2528,N_1844);
and U6760 (N_6760,N_996,N_4527);
and U6761 (N_6761,N_3228,N_1597);
or U6762 (N_6762,N_2520,N_576);
nand U6763 (N_6763,N_3901,N_2329);
and U6764 (N_6764,N_2714,N_2930);
nand U6765 (N_6765,N_4454,N_2920);
nor U6766 (N_6766,N_2724,N_4977);
and U6767 (N_6767,N_3753,N_1134);
nand U6768 (N_6768,N_1449,N_2231);
nand U6769 (N_6769,N_3659,N_1866);
or U6770 (N_6770,N_1760,N_3443);
nand U6771 (N_6771,N_4364,N_1129);
or U6772 (N_6772,N_1810,N_4489);
and U6773 (N_6773,N_1293,N_4124);
or U6774 (N_6774,N_1124,N_3202);
nor U6775 (N_6775,N_4919,N_1980);
and U6776 (N_6776,N_3735,N_929);
nor U6777 (N_6777,N_1254,N_3712);
nor U6778 (N_6778,N_769,N_2741);
nor U6779 (N_6779,N_4676,N_104);
and U6780 (N_6780,N_591,N_52);
or U6781 (N_6781,N_3793,N_725);
and U6782 (N_6782,N_2338,N_1670);
xnor U6783 (N_6783,N_2649,N_2839);
and U6784 (N_6784,N_3418,N_2747);
or U6785 (N_6785,N_4314,N_3597);
nor U6786 (N_6786,N_2775,N_2141);
nor U6787 (N_6787,N_4525,N_2041);
nand U6788 (N_6788,N_1723,N_4560);
nor U6789 (N_6789,N_4956,N_3532);
nor U6790 (N_6790,N_1950,N_953);
nor U6791 (N_6791,N_98,N_110);
nor U6792 (N_6792,N_2969,N_2937);
and U6793 (N_6793,N_4715,N_3420);
and U6794 (N_6794,N_3180,N_3729);
and U6795 (N_6795,N_3342,N_3361);
and U6796 (N_6796,N_4170,N_1016);
xor U6797 (N_6797,N_2522,N_2558);
nand U6798 (N_6798,N_2798,N_2479);
nor U6799 (N_6799,N_4824,N_1884);
and U6800 (N_6800,N_1829,N_177);
nor U6801 (N_6801,N_3940,N_1621);
xnor U6802 (N_6802,N_961,N_1282);
or U6803 (N_6803,N_3997,N_4557);
or U6804 (N_6804,N_648,N_1780);
and U6805 (N_6805,N_3953,N_3562);
nor U6806 (N_6806,N_2881,N_735);
nand U6807 (N_6807,N_3839,N_3436);
and U6808 (N_6808,N_1770,N_3157);
and U6809 (N_6809,N_212,N_2512);
and U6810 (N_6810,N_565,N_3852);
and U6811 (N_6811,N_1744,N_2380);
and U6812 (N_6812,N_3614,N_2701);
and U6813 (N_6813,N_2193,N_2716);
and U6814 (N_6814,N_3666,N_4049);
nand U6815 (N_6815,N_1949,N_3097);
or U6816 (N_6816,N_911,N_3639);
nor U6817 (N_6817,N_1288,N_2967);
nor U6818 (N_6818,N_1545,N_3057);
and U6819 (N_6819,N_3516,N_1383);
nor U6820 (N_6820,N_2790,N_3025);
nor U6821 (N_6821,N_2473,N_3795);
nor U6822 (N_6822,N_3711,N_3121);
and U6823 (N_6823,N_3186,N_1804);
and U6824 (N_6824,N_1098,N_1952);
and U6825 (N_6825,N_4929,N_1012);
and U6826 (N_6826,N_1654,N_3557);
and U6827 (N_6827,N_4863,N_1076);
nand U6828 (N_6828,N_194,N_3866);
nand U6829 (N_6829,N_1703,N_4443);
nand U6830 (N_6830,N_1069,N_4241);
nand U6831 (N_6831,N_4086,N_3802);
and U6832 (N_6832,N_2084,N_757);
nor U6833 (N_6833,N_783,N_2987);
nor U6834 (N_6834,N_4317,N_489);
or U6835 (N_6835,N_2633,N_3694);
nand U6836 (N_6836,N_161,N_614);
nand U6837 (N_6837,N_3067,N_4257);
nand U6838 (N_6838,N_4386,N_4871);
or U6839 (N_6839,N_3620,N_1256);
and U6840 (N_6840,N_4832,N_4071);
nor U6841 (N_6841,N_2982,N_1489);
or U6842 (N_6842,N_4349,N_4597);
nand U6843 (N_6843,N_3941,N_2344);
nor U6844 (N_6844,N_1722,N_2950);
and U6845 (N_6845,N_965,N_3153);
nor U6846 (N_6846,N_4235,N_2591);
and U6847 (N_6847,N_461,N_1733);
nand U6848 (N_6848,N_4137,N_4471);
or U6849 (N_6849,N_4774,N_2106);
or U6850 (N_6850,N_2083,N_3543);
and U6851 (N_6851,N_333,N_880);
nand U6852 (N_6852,N_1436,N_621);
and U6853 (N_6853,N_2314,N_3774);
and U6854 (N_6854,N_708,N_2681);
and U6855 (N_6855,N_1611,N_3662);
nand U6856 (N_6856,N_2249,N_3170);
and U6857 (N_6857,N_2034,N_3296);
or U6858 (N_6858,N_3676,N_1034);
or U6859 (N_6859,N_957,N_1549);
or U6860 (N_6860,N_4186,N_3899);
nor U6861 (N_6861,N_976,N_4992);
nor U6862 (N_6862,N_2113,N_561);
and U6863 (N_6863,N_2327,N_3908);
or U6864 (N_6864,N_2643,N_145);
or U6865 (N_6865,N_2896,N_1988);
or U6866 (N_6866,N_1087,N_2972);
nor U6867 (N_6867,N_4139,N_2769);
and U6868 (N_6868,N_599,N_3933);
or U6869 (N_6869,N_3165,N_1913);
or U6870 (N_6870,N_818,N_4451);
nor U6871 (N_6871,N_3791,N_227);
nor U6872 (N_6872,N_913,N_2563);
and U6873 (N_6873,N_1224,N_469);
and U6874 (N_6874,N_2275,N_2998);
and U6875 (N_6875,N_2776,N_4294);
nand U6876 (N_6876,N_615,N_556);
and U6877 (N_6877,N_1183,N_3310);
nor U6878 (N_6878,N_3825,N_1364);
nand U6879 (N_6879,N_1289,N_3019);
and U6880 (N_6880,N_3347,N_4115);
or U6881 (N_6881,N_1051,N_126);
nand U6882 (N_6882,N_3311,N_4577);
nand U6883 (N_6883,N_4901,N_1257);
nor U6884 (N_6884,N_1666,N_128);
and U6885 (N_6885,N_74,N_1998);
or U6886 (N_6886,N_505,N_1759);
nand U6887 (N_6887,N_4748,N_282);
nor U6888 (N_6888,N_3040,N_3748);
or U6889 (N_6889,N_500,N_776);
and U6890 (N_6890,N_1414,N_1577);
nand U6891 (N_6891,N_3558,N_3154);
and U6892 (N_6892,N_412,N_4191);
nand U6893 (N_6893,N_2463,N_4562);
nor U6894 (N_6894,N_3273,N_348);
or U6895 (N_6895,N_3946,N_3419);
xnor U6896 (N_6896,N_1707,N_2859);
and U6897 (N_6897,N_331,N_1697);
nand U6898 (N_6898,N_2263,N_2648);
nor U6899 (N_6899,N_948,N_4485);
and U6900 (N_6900,N_4827,N_4366);
or U6901 (N_6901,N_3136,N_2755);
or U6902 (N_6902,N_1821,N_484);
and U6903 (N_6903,N_4942,N_1073);
or U6904 (N_6904,N_4505,N_4706);
nand U6905 (N_6905,N_3844,N_1978);
nor U6906 (N_6906,N_70,N_1920);
and U6907 (N_6907,N_1676,N_1655);
or U6908 (N_6908,N_3982,N_4343);
nand U6909 (N_6909,N_963,N_4932);
xnor U6910 (N_6910,N_4854,N_4048);
nor U6911 (N_6911,N_3410,N_2532);
nor U6912 (N_6912,N_12,N_3514);
or U6913 (N_6913,N_4732,N_1584);
nand U6914 (N_6914,N_2768,N_3594);
or U6915 (N_6915,N_1347,N_3018);
or U6916 (N_6916,N_1102,N_3241);
and U6917 (N_6917,N_1698,N_2940);
nor U6918 (N_6918,N_1756,N_332);
nand U6919 (N_6919,N_3141,N_4635);
nor U6920 (N_6920,N_3914,N_4332);
and U6921 (N_6921,N_4893,N_2709);
or U6922 (N_6922,N_1253,N_300);
or U6923 (N_6923,N_799,N_2319);
nand U6924 (N_6924,N_4482,N_4423);
or U6925 (N_6925,N_112,N_447);
or U6926 (N_6926,N_2573,N_632);
nand U6927 (N_6927,N_4801,N_2675);
and U6928 (N_6928,N_39,N_1310);
or U6929 (N_6929,N_278,N_3781);
and U6930 (N_6930,N_3161,N_2459);
and U6931 (N_6931,N_1411,N_4473);
nand U6932 (N_6932,N_4846,N_3862);
xor U6933 (N_6933,N_910,N_4027);
or U6934 (N_6934,N_4661,N_4194);
or U6935 (N_6935,N_833,N_3321);
nand U6936 (N_6936,N_1457,N_254);
or U6937 (N_6937,N_3583,N_415);
or U6938 (N_6938,N_2983,N_1796);
or U6939 (N_6939,N_1785,N_2007);
nand U6940 (N_6940,N_4659,N_4521);
nor U6941 (N_6941,N_1578,N_2320);
or U6942 (N_6942,N_1790,N_4522);
nor U6943 (N_6943,N_1497,N_3629);
nand U6944 (N_6944,N_3951,N_1423);
and U6945 (N_6945,N_960,N_1563);
or U6946 (N_6946,N_2787,N_4199);
nor U6947 (N_6947,N_3881,N_178);
nand U6948 (N_6948,N_988,N_938);
nor U6949 (N_6949,N_4344,N_2779);
and U6950 (N_6950,N_4046,N_3138);
nor U6951 (N_6951,N_3137,N_2359);
and U6952 (N_6952,N_3075,N_3627);
and U6953 (N_6953,N_4331,N_4075);
nand U6954 (N_6954,N_3840,N_1159);
nand U6955 (N_6955,N_3869,N_3485);
nor U6956 (N_6956,N_2087,N_1301);
nor U6957 (N_6957,N_1294,N_1956);
and U6958 (N_6958,N_3706,N_203);
nor U6959 (N_6959,N_1348,N_1488);
nand U6960 (N_6960,N_423,N_385);
or U6961 (N_6961,N_1660,N_1439);
and U6962 (N_6962,N_351,N_2310);
and U6963 (N_6963,N_2066,N_2576);
nor U6964 (N_6964,N_3091,N_4670);
and U6965 (N_6965,N_2270,N_664);
or U6966 (N_6966,N_2454,N_2350);
nor U6967 (N_6967,N_2039,N_4417);
or U6968 (N_6968,N_4978,N_884);
nor U6969 (N_6969,N_4745,N_4047);
xor U6970 (N_6970,N_542,N_4403);
and U6971 (N_6971,N_2002,N_2028);
or U6972 (N_6972,N_711,N_3328);
nor U6973 (N_6973,N_3159,N_4565);
nor U6974 (N_6974,N_474,N_1353);
nor U6975 (N_6975,N_1918,N_2287);
and U6976 (N_6976,N_2396,N_1638);
nor U6977 (N_6977,N_3107,N_4267);
nand U6978 (N_6978,N_2585,N_4642);
and U6979 (N_6979,N_1397,N_2821);
and U6980 (N_6980,N_4477,N_405);
and U6981 (N_6981,N_2782,N_856);
nand U6982 (N_6982,N_223,N_2035);
nor U6983 (N_6983,N_3571,N_2067);
or U6984 (N_6984,N_3535,N_87);
nand U6985 (N_6985,N_1136,N_4885);
and U6986 (N_6986,N_4907,N_4976);
nand U6987 (N_6987,N_1346,N_3687);
or U6988 (N_6988,N_2916,N_2517);
nand U6989 (N_6989,N_738,N_3051);
or U6990 (N_6990,N_1736,N_1160);
or U6991 (N_6991,N_2939,N_2153);
and U6992 (N_6992,N_3988,N_1747);
or U6993 (N_6993,N_2628,N_4370);
and U6994 (N_6994,N_4180,N_4411);
or U6995 (N_6995,N_1667,N_3285);
nand U6996 (N_6996,N_2921,N_3294);
or U6997 (N_6997,N_4379,N_1481);
nand U6998 (N_6998,N_3185,N_175);
nor U6999 (N_6999,N_1372,N_1906);
nand U7000 (N_7000,N_2557,N_1103);
xnor U7001 (N_7001,N_9,N_2954);
nor U7002 (N_7002,N_4060,N_3880);
nand U7003 (N_7003,N_1679,N_4450);
or U7004 (N_7004,N_353,N_1857);
or U7005 (N_7005,N_2160,N_3017);
nand U7006 (N_7006,N_3481,N_701);
nor U7007 (N_7007,N_4272,N_281);
nor U7008 (N_7008,N_1710,N_3134);
nor U7009 (N_7009,N_4053,N_3439);
or U7010 (N_7010,N_1268,N_2570);
nor U7011 (N_7011,N_1686,N_2819);
and U7012 (N_7012,N_2702,N_1336);
nor U7013 (N_7013,N_1305,N_1721);
nand U7014 (N_7014,N_2531,N_970);
and U7015 (N_7015,N_3656,N_868);
and U7016 (N_7016,N_1769,N_3660);
nor U7017 (N_7017,N_2062,N_3316);
xor U7018 (N_7018,N_4032,N_1651);
xnor U7019 (N_7019,N_2102,N_4385);
nand U7020 (N_7020,N_156,N_1061);
nor U7021 (N_7021,N_660,N_4480);
nand U7022 (N_7022,N_4512,N_4594);
nand U7023 (N_7023,N_1402,N_946);
nor U7024 (N_7024,N_3102,N_4851);
or U7025 (N_7025,N_4936,N_2299);
and U7026 (N_7026,N_3232,N_3284);
nand U7027 (N_7027,N_2644,N_1963);
nand U7028 (N_7028,N_1454,N_2720);
and U7029 (N_7029,N_4760,N_3836);
or U7030 (N_7030,N_2721,N_4132);
and U7031 (N_7031,N_564,N_1384);
or U7032 (N_7032,N_3408,N_4680);
and U7033 (N_7033,N_1626,N_3762);
nand U7034 (N_7034,N_2107,N_3577);
nand U7035 (N_7035,N_4744,N_204);
and U7036 (N_7036,N_3253,N_470);
nor U7037 (N_7037,N_4910,N_1062);
or U7038 (N_7038,N_4847,N_2449);
or U7039 (N_7039,N_2495,N_2516);
and U7040 (N_7040,N_4422,N_2285);
or U7041 (N_7041,N_1753,N_1515);
nand U7042 (N_7042,N_3937,N_36);
xor U7043 (N_7043,N_4099,N_1573);
nand U7044 (N_7044,N_3564,N_290);
and U7045 (N_7045,N_2044,N_620);
nor U7046 (N_7046,N_861,N_89);
nand U7047 (N_7047,N_2204,N_3492);
nor U7048 (N_7048,N_4791,N_2975);
or U7049 (N_7049,N_3341,N_2456);
nor U7050 (N_7050,N_2142,N_3548);
nor U7051 (N_7051,N_4996,N_594);
or U7052 (N_7052,N_2544,N_4361);
and U7053 (N_7053,N_1901,N_2478);
nor U7054 (N_7054,N_4831,N_4266);
nor U7055 (N_7055,N_4861,N_3119);
nor U7056 (N_7056,N_4025,N_3401);
or U7057 (N_7057,N_3196,N_256);
nor U7058 (N_7058,N_4449,N_2425);
nor U7059 (N_7059,N_4113,N_3654);
or U7060 (N_7060,N_958,N_3962);
and U7061 (N_7061,N_1214,N_3338);
nor U7062 (N_7062,N_414,N_1801);
nand U7063 (N_7063,N_2009,N_3123);
or U7064 (N_7064,N_1249,N_355);
or U7065 (N_7065,N_3544,N_1140);
or U7066 (N_7066,N_4666,N_642);
or U7067 (N_7067,N_3868,N_1517);
or U7068 (N_7068,N_2689,N_2050);
xnor U7069 (N_7069,N_1716,N_4248);
nand U7070 (N_7070,N_1412,N_4990);
or U7071 (N_7071,N_4187,N_480);
nand U7072 (N_7072,N_2695,N_4472);
xnor U7073 (N_7073,N_1599,N_1960);
and U7074 (N_7074,N_105,N_984);
and U7075 (N_7075,N_1583,N_2288);
and U7076 (N_7076,N_2906,N_3440);
nor U7077 (N_7077,N_1658,N_4263);
and U7078 (N_7078,N_1550,N_4218);
or U7079 (N_7079,N_3374,N_1026);
and U7080 (N_7080,N_3886,N_1524);
nand U7081 (N_7081,N_4540,N_3226);
nor U7082 (N_7082,N_3477,N_2750);
xnor U7083 (N_7083,N_2866,N_1206);
or U7084 (N_7084,N_3758,N_2683);
nor U7085 (N_7085,N_1608,N_860);
or U7086 (N_7086,N_2511,N_3496);
nor U7087 (N_7087,N_3434,N_4604);
nor U7088 (N_7088,N_1417,N_53);
and U7089 (N_7089,N_3619,N_1546);
and U7090 (N_7090,N_4914,N_3498);
nand U7091 (N_7091,N_96,N_674);
and U7092 (N_7092,N_4703,N_750);
nor U7093 (N_7093,N_444,N_4663);
and U7094 (N_7094,N_1598,N_968);
and U7095 (N_7095,N_4993,N_4668);
nand U7096 (N_7096,N_675,N_159);
nor U7097 (N_7097,N_4110,N_4122);
nand U7098 (N_7098,N_1357,N_2468);
nand U7099 (N_7099,N_2252,N_3048);
or U7100 (N_7100,N_921,N_92);
nor U7101 (N_7101,N_2215,N_2333);
nand U7102 (N_7102,N_440,N_2151);
nor U7103 (N_7103,N_858,N_4169);
or U7104 (N_7104,N_3831,N_1943);
nand U7105 (N_7105,N_1700,N_1117);
nor U7106 (N_7106,N_4253,N_2642);
and U7107 (N_7107,N_285,N_4646);
and U7108 (N_7108,N_2190,N_3359);
and U7109 (N_7109,N_3907,N_4860);
nand U7110 (N_7110,N_4713,N_2281);
nor U7111 (N_7111,N_3981,N_1763);
nor U7112 (N_7112,N_692,N_2126);
or U7113 (N_7113,N_4431,N_1728);
and U7114 (N_7114,N_932,N_3448);
and U7115 (N_7115,N_1175,N_2584);
nand U7116 (N_7116,N_2418,N_2922);
or U7117 (N_7117,N_1508,N_231);
nand U7118 (N_7118,N_3330,N_3902);
or U7119 (N_7119,N_4282,N_791);
or U7120 (N_7120,N_4384,N_767);
nand U7121 (N_7121,N_1878,N_4599);
and U7122 (N_7122,N_261,N_4249);
and U7123 (N_7123,N_1499,N_3678);
nor U7124 (N_7124,N_669,N_3527);
or U7125 (N_7125,N_1830,N_1843);
and U7126 (N_7126,N_1822,N_4876);
nand U7127 (N_7127,N_4772,N_1717);
nand U7128 (N_7128,N_4410,N_2184);
and U7129 (N_7129,N_3691,N_2527);
nand U7130 (N_7130,N_1185,N_1146);
or U7131 (N_7131,N_1957,N_3883);
and U7132 (N_7132,N_2399,N_4537);
nor U7133 (N_7133,N_3985,N_1522);
nor U7134 (N_7134,N_3495,N_1326);
or U7135 (N_7135,N_1944,N_1902);
nand U7136 (N_7136,N_2661,N_4419);
and U7137 (N_7137,N_91,N_4350);
nand U7138 (N_7138,N_4463,N_1701);
nand U7139 (N_7139,N_3772,N_4897);
nor U7140 (N_7140,N_4641,N_959);
nor U7141 (N_7141,N_927,N_3784);
or U7142 (N_7142,N_906,N_131);
nand U7143 (N_7143,N_1937,N_3390);
and U7144 (N_7144,N_3027,N_2871);
nand U7145 (N_7145,N_1737,N_1443);
nor U7146 (N_7146,N_1720,N_4055);
nor U7147 (N_7147,N_407,N_1340);
nor U7148 (N_7148,N_4502,N_3776);
nor U7149 (N_7149,N_3517,N_2588);
nand U7150 (N_7150,N_4725,N_4575);
nand U7151 (N_7151,N_2212,N_4719);
nand U7152 (N_7152,N_1266,N_100);
nor U7153 (N_7153,N_511,N_2173);
nor U7154 (N_7154,N_3104,N_4009);
nand U7155 (N_7155,N_375,N_742);
and U7156 (N_7156,N_2435,N_4226);
or U7157 (N_7157,N_983,N_4623);
nand U7158 (N_7158,N_1142,N_4397);
and U7159 (N_7159,N_3569,N_668);
nor U7160 (N_7160,N_1675,N_47);
or U7161 (N_7161,N_2078,N_1404);
and U7162 (N_7162,N_4015,N_4029);
xor U7163 (N_7163,N_1351,N_4437);
and U7164 (N_7164,N_4181,N_838);
xor U7165 (N_7165,N_2098,N_2953);
and U7166 (N_7166,N_124,N_130);
nor U7167 (N_7167,N_1695,N_427);
nor U7168 (N_7168,N_3383,N_2017);
nand U7169 (N_7169,N_1824,N_3720);
nor U7170 (N_7170,N_1773,N_717);
or U7171 (N_7171,N_2432,N_4735);
or U7172 (N_7172,N_2825,N_2851);
and U7173 (N_7173,N_4656,N_1798);
and U7174 (N_7174,N_2097,N_2309);
nand U7175 (N_7175,N_2547,N_3377);
nand U7176 (N_7176,N_4305,N_944);
or U7177 (N_7177,N_4007,N_4223);
and U7178 (N_7178,N_2467,N_3721);
or U7179 (N_7179,N_1074,N_311);
nand U7180 (N_7180,N_1817,N_4002);
nand U7181 (N_7181,N_3128,N_3317);
or U7182 (N_7182,N_1139,N_3728);
nor U7183 (N_7183,N_1634,N_4230);
or U7184 (N_7184,N_2360,N_4879);
and U7185 (N_7185,N_81,N_1250);
or U7186 (N_7186,N_2260,N_2195);
or U7187 (N_7187,N_4998,N_2159);
and U7188 (N_7188,N_3574,N_900);
nor U7189 (N_7189,N_952,N_3551);
or U7190 (N_7190,N_2094,N_3991);
or U7191 (N_7191,N_2811,N_2929);
and U7192 (N_7192,N_3209,N_1225);
and U7193 (N_7193,N_4142,N_4980);
xor U7194 (N_7194,N_4789,N_1377);
or U7195 (N_7195,N_1847,N_3888);
nor U7196 (N_7196,N_4130,N_508);
or U7197 (N_7197,N_4701,N_3837);
or U7198 (N_7198,N_1498,N_4373);
and U7199 (N_7199,N_4883,N_2403);
or U7200 (N_7200,N_2673,N_4682);
or U7201 (N_7201,N_1143,N_16);
or U7202 (N_7202,N_994,N_1751);
or U7203 (N_7203,N_555,N_1317);
nand U7204 (N_7204,N_3391,N_1063);
and U7205 (N_7205,N_790,N_4092);
and U7206 (N_7206,N_1337,N_4606);
nor U7207 (N_7207,N_656,N_1641);
nor U7208 (N_7208,N_4475,N_1931);
and U7209 (N_7209,N_622,N_3928);
xor U7210 (N_7210,N_3858,N_463);
nor U7211 (N_7211,N_4304,N_1100);
or U7212 (N_7212,N_1985,N_1519);
or U7213 (N_7213,N_2941,N_2238);
nor U7214 (N_7214,N_3686,N_2315);
and U7215 (N_7215,N_2401,N_1077);
or U7216 (N_7216,N_2590,N_1504);
nand U7217 (N_7217,N_3482,N_3307);
or U7218 (N_7218,N_2433,N_1278);
xor U7219 (N_7219,N_4018,N_1565);
nor U7220 (N_7220,N_1333,N_3747);
or U7221 (N_7221,N_1669,N_3478);
nand U7222 (N_7222,N_1959,N_2487);
nor U7223 (N_7223,N_228,N_3455);
and U7224 (N_7224,N_1408,N_140);
or U7225 (N_7225,N_3367,N_3351);
xor U7226 (N_7226,N_4905,N_506);
nand U7227 (N_7227,N_1023,N_1391);
nor U7228 (N_7228,N_3125,N_3520);
or U7229 (N_7229,N_2262,N_291);
or U7230 (N_7230,N_4737,N_3329);
and U7231 (N_7231,N_1915,N_631);
or U7232 (N_7232,N_398,N_1361);
or U7233 (N_7233,N_3333,N_4954);
nand U7234 (N_7234,N_4862,N_2008);
nor U7235 (N_7235,N_4308,N_2672);
and U7236 (N_7236,N_4091,N_4843);
nand U7237 (N_7237,N_3979,N_4250);
or U7238 (N_7238,N_2137,N_587);
and U7239 (N_7239,N_2973,N_4811);
or U7240 (N_7240,N_1890,N_270);
nor U7241 (N_7241,N_1904,N_3365);
nor U7242 (N_7242,N_519,N_249);
nor U7243 (N_7243,N_1036,N_4683);
or U7244 (N_7244,N_1609,N_2533);
and U7245 (N_7245,N_364,N_1277);
or U7246 (N_7246,N_1246,N_2030);
or U7247 (N_7247,N_1085,N_2788);
nand U7248 (N_7248,N_269,N_3016);
nand U7249 (N_7249,N_4301,N_4549);
and U7250 (N_7250,N_3591,N_4690);
or U7251 (N_7251,N_3013,N_2892);
and U7252 (N_7252,N_1447,N_4050);
and U7253 (N_7253,N_3400,N_4957);
and U7254 (N_7254,N_4718,N_2129);
and U7255 (N_7255,N_193,N_266);
or U7256 (N_7256,N_253,N_103);
nand U7257 (N_7257,N_3463,N_1604);
nand U7258 (N_7258,N_4751,N_857);
nor U7259 (N_7259,N_3238,N_349);
nand U7260 (N_7260,N_2110,N_2564);
or U7261 (N_7261,N_1536,N_4088);
or U7262 (N_7262,N_4201,N_3122);
or U7263 (N_7263,N_2423,N_3315);
nand U7264 (N_7264,N_1476,N_575);
nand U7265 (N_7265,N_2823,N_4357);
and U7266 (N_7266,N_1267,N_2518);
nand U7267 (N_7267,N_1967,N_2893);
nor U7268 (N_7268,N_148,N_3923);
nor U7269 (N_7269,N_3578,N_1888);
and U7270 (N_7270,N_2416,N_4374);
nor U7271 (N_7271,N_109,N_2727);
and U7272 (N_7272,N_1809,N_10);
or U7273 (N_7273,N_4459,N_59);
xnor U7274 (N_7274,N_3661,N_3699);
nor U7275 (N_7275,N_1111,N_1984);
nor U7276 (N_7276,N_2864,N_2530);
or U7277 (N_7277,N_643,N_3261);
or U7278 (N_7278,N_3280,N_1410);
nand U7279 (N_7279,N_2366,N_4136);
or U7280 (N_7280,N_894,N_2909);
nand U7281 (N_7281,N_1090,N_3042);
or U7282 (N_7282,N_5,N_855);
nand U7283 (N_7283,N_841,N_1205);
and U7284 (N_7284,N_3993,N_1833);
and U7285 (N_7285,N_3110,N_142);
nor U7286 (N_7286,N_2491,N_2053);
and U7287 (N_7287,N_4457,N_531);
and U7288 (N_7288,N_875,N_1399);
or U7289 (N_7289,N_4141,N_4056);
nor U7290 (N_7290,N_2409,N_1531);
or U7291 (N_7291,N_3208,N_2134);
nor U7292 (N_7292,N_895,N_2006);
or U7293 (N_7293,N_4777,N_1925);
nand U7294 (N_7294,N_4583,N_538);
or U7295 (N_7295,N_804,N_3248);
nand U7296 (N_7296,N_218,N_4150);
nand U7297 (N_7297,N_1042,N_135);
or U7298 (N_7298,N_1730,N_3237);
nor U7299 (N_7299,N_4771,N_812);
and U7300 (N_7300,N_4961,N_3058);
or U7301 (N_7301,N_2012,N_2471);
nand U7302 (N_7302,N_2258,N_90);
or U7303 (N_7303,N_1704,N_3947);
nand U7304 (N_7304,N_4543,N_4943);
nor U7305 (N_7305,N_1260,N_4934);
or U7306 (N_7306,N_75,N_4716);
nand U7307 (N_7307,N_1652,N_3760);
or U7308 (N_7308,N_2324,N_1375);
nand U7309 (N_7309,N_1316,N_232);
or U7310 (N_7310,N_2593,N_930);
or U7311 (N_7311,N_2130,N_3674);
nor U7312 (N_7312,N_3644,N_1110);
and U7313 (N_7313,N_3522,N_1083);
nand U7314 (N_7314,N_1689,N_1030);
nand U7315 (N_7315,N_4028,N_3096);
nor U7316 (N_7316,N_2540,N_1633);
nand U7317 (N_7317,N_766,N_2808);
and U7318 (N_7318,N_1592,N_2565);
or U7319 (N_7319,N_1500,N_2783);
and U7320 (N_7320,N_4416,N_4694);
or U7321 (N_7321,N_1795,N_3932);
and U7322 (N_7322,N_4478,N_1028);
nand U7323 (N_7323,N_623,N_3113);
and U7324 (N_7324,N_726,N_2269);
or U7325 (N_7325,N_4685,N_1916);
nand U7326 (N_7326,N_521,N_1614);
nor U7327 (N_7327,N_4095,N_1627);
and U7328 (N_7328,N_2112,N_1576);
and U7329 (N_7329,N_681,N_4014);
or U7330 (N_7330,N_607,N_4217);
and U7331 (N_7331,N_3092,N_4310);
or U7332 (N_7332,N_2676,N_3630);
or U7333 (N_7333,N_1480,N_554);
or U7334 (N_7334,N_4551,N_3098);
or U7335 (N_7335,N_811,N_1648);
or U7336 (N_7336,N_72,N_3483);
nand U7337 (N_7337,N_1554,N_1861);
nor U7338 (N_7338,N_2057,N_892);
and U7339 (N_7339,N_2152,N_1643);
nand U7340 (N_7340,N_4753,N_1718);
nand U7341 (N_7341,N_2158,N_1872);
or U7342 (N_7342,N_2276,N_2064);
or U7343 (N_7343,N_585,N_3203);
nand U7344 (N_7344,N_843,N_3479);
nor U7345 (N_7345,N_1754,N_809);
nor U7346 (N_7346,N_4116,N_3751);
and U7347 (N_7347,N_4251,N_1640);
and U7348 (N_7348,N_1740,N_924);
or U7349 (N_7349,N_4564,N_4850);
or U7350 (N_7350,N_359,N_3046);
or U7351 (N_7351,N_384,N_2980);
nor U7352 (N_7352,N_4140,N_386);
and U7353 (N_7353,N_3652,N_2199);
and U7354 (N_7354,N_4322,N_3236);
nor U7355 (N_7355,N_1782,N_2567);
and U7356 (N_7356,N_1705,N_3733);
and U7357 (N_7357,N_479,N_3570);
or U7358 (N_7358,N_3567,N_1482);
nor U7359 (N_7359,N_2446,N_4441);
nand U7360 (N_7360,N_107,N_2027);
nor U7361 (N_7361,N_4698,N_2265);
or U7362 (N_7362,N_298,N_1152);
or U7363 (N_7363,N_3830,N_1479);
nand U7364 (N_7364,N_779,N_908);
nor U7365 (N_7365,N_3555,N_1426);
nand U7366 (N_7366,N_2049,N_4316);
or U7367 (N_7367,N_1176,N_3855);
and U7368 (N_7368,N_1354,N_666);
and U7369 (N_7369,N_847,N_850);
nor U7370 (N_7370,N_237,N_1339);
nor U7371 (N_7371,N_1428,N_2402);
nor U7372 (N_7372,N_1473,N_4213);
or U7373 (N_7373,N_3004,N_760);
nor U7374 (N_7374,N_1105,N_139);
or U7375 (N_7375,N_2542,N_221);
nor U7376 (N_7376,N_2502,N_2600);
or U7377 (N_7377,N_3403,N_1274);
or U7378 (N_7378,N_2794,N_1580);
nor U7379 (N_7379,N_514,N_1371);
or U7380 (N_7380,N_370,N_4574);
nand U7381 (N_7381,N_3371,N_4782);
nand U7382 (N_7382,N_1401,N_2114);
nand U7383 (N_7383,N_4227,N_797);
and U7384 (N_7384,N_3563,N_3324);
nor U7385 (N_7385,N_1486,N_2);
and U7386 (N_7386,N_2323,N_1046);
or U7387 (N_7387,N_2089,N_1729);
nand U7388 (N_7388,N_639,N_1854);
nor U7389 (N_7389,N_4590,N_4495);
nand U7390 (N_7390,N_3622,N_1612);
nor U7391 (N_7391,N_4681,N_3221);
or U7392 (N_7392,N_176,N_3701);
or U7393 (N_7393,N_3819,N_3056);
or U7394 (N_7394,N_507,N_2472);
or U7395 (N_7395,N_2597,N_854);
or U7396 (N_7396,N_4196,N_387);
xnor U7397 (N_7397,N_1240,N_380);
nor U7398 (N_7398,N_235,N_4031);
or U7399 (N_7399,N_4307,N_702);
nor U7400 (N_7400,N_4839,N_27);
nor U7401 (N_7401,N_4120,N_1932);
nand U7402 (N_7402,N_1559,N_1184);
or U7403 (N_7403,N_99,N_3780);
and U7404 (N_7404,N_4667,N_1628);
and U7405 (N_7405,N_358,N_1170);
and U7406 (N_7406,N_1047,N_1415);
and U7407 (N_7407,N_3217,N_3424);
or U7408 (N_7408,N_1569,N_1875);
and U7409 (N_7409,N_2037,N_2069);
or U7410 (N_7410,N_4433,N_4456);
nand U7411 (N_7411,N_1818,N_3174);
or U7412 (N_7412,N_4915,N_4283);
nor U7413 (N_7413,N_3653,N_449);
nand U7414 (N_7414,N_445,N_3265);
xor U7415 (N_7415,N_2046,N_4388);
nor U7416 (N_7416,N_191,N_3111);
and U7417 (N_7417,N_2205,N_1459);
or U7418 (N_7418,N_977,N_520);
nor U7419 (N_7419,N_2933,N_1819);
and U7420 (N_7420,N_1286,N_4975);
nor U7421 (N_7421,N_1044,N_624);
and U7422 (N_7422,N_1865,N_901);
nor U7423 (N_7423,N_1466,N_1405);
nor U7424 (N_7424,N_2226,N_1789);
or U7425 (N_7425,N_2690,N_2221);
or U7426 (N_7426,N_2529,N_3083);
or U7427 (N_7427,N_4528,N_4625);
nand U7428 (N_7428,N_4037,N_2928);
and U7429 (N_7429,N_4638,N_1603);
nor U7430 (N_7430,N_2550,N_3049);
and U7431 (N_7431,N_2115,N_1992);
and U7432 (N_7432,N_2912,N_3145);
and U7433 (N_7433,N_3109,N_4105);
nor U7434 (N_7434,N_3530,N_2985);
or U7435 (N_7435,N_4222,N_2617);
nand U7436 (N_7436,N_4924,N_4585);
or U7437 (N_7437,N_65,N_1053);
and U7438 (N_7438,N_4234,N_1174);
nand U7439 (N_7439,N_3344,N_2688);
or U7440 (N_7440,N_569,N_2368);
or U7441 (N_7441,N_3218,N_2486);
nand U7442 (N_7442,N_4291,N_4202);
nor U7443 (N_7443,N_1644,N_1523);
xor U7444 (N_7444,N_885,N_1195);
nand U7445 (N_7445,N_2273,N_805);
or U7446 (N_7446,N_1661,N_4465);
nand U7447 (N_7447,N_2105,N_2915);
and U7448 (N_7448,N_3655,N_3800);
or U7449 (N_7449,N_3143,N_2373);
nand U7450 (N_7450,N_882,N_3063);
or U7451 (N_7451,N_539,N_3432);
and U7452 (N_7452,N_3755,N_2136);
nand U7453 (N_7453,N_3964,N_2365);
and U7454 (N_7454,N_4395,N_1027);
or U7455 (N_7455,N_3636,N_4741);
and U7456 (N_7456,N_2243,N_3702);
nand U7457 (N_7457,N_54,N_570);
nor U7458 (N_7458,N_2604,N_2268);
nand U7459 (N_7459,N_4414,N_2122);
or U7460 (N_7460,N_595,N_1602);
or U7461 (N_7461,N_342,N_2244);
or U7462 (N_7462,N_3607,N_357);
or U7463 (N_7463,N_829,N_4168);
nand U7464 (N_7464,N_898,N_4704);
and U7465 (N_7465,N_3859,N_3276);
and U7466 (N_7466,N_3641,N_1513);
or U7467 (N_7467,N_2703,N_4842);
nand U7468 (N_7468,N_3105,N_4243);
or U7469 (N_7469,N_1965,N_3073);
or U7470 (N_7470,N_2342,N_846);
nor U7471 (N_7471,N_1237,N_1725);
nand U7472 (N_7472,N_2048,N_1307);
or U7473 (N_7473,N_1811,N_1007);
and U7474 (N_7474,N_4727,N_4699);
nand U7475 (N_7475,N_3000,N_2139);
nor U7476 (N_7476,N_1024,N_2203);
nand U7477 (N_7477,N_645,N_2222);
and U7478 (N_7478,N_3987,N_3605);
or U7479 (N_7479,N_1886,N_4024);
and U7480 (N_7480,N_907,N_2311);
nand U7481 (N_7481,N_3014,N_1032);
and U7482 (N_7482,N_435,N_4052);
and U7483 (N_7483,N_35,N_1156);
nor U7484 (N_7484,N_499,N_4274);
nand U7485 (N_7485,N_3773,N_2979);
nor U7486 (N_7486,N_3510,N_4336);
nand U7487 (N_7487,N_446,N_170);
nor U7488 (N_7488,N_3689,N_1934);
nand U7489 (N_7489,N_2777,N_2149);
nor U7490 (N_7490,N_1055,N_2861);
or U7491 (N_7491,N_3618,N_4750);
nand U7492 (N_7492,N_3588,N_2116);
nand U7493 (N_7493,N_1400,N_2284);
nor U7494 (N_7494,N_4619,N_4290);
nand U7495 (N_7495,N_1678,N_3846);
nor U7496 (N_7496,N_319,N_4166);
and U7497 (N_7497,N_93,N_4755);
and U7498 (N_7498,N_680,N_4269);
nor U7499 (N_7499,N_3454,N_3790);
and U7500 (N_7500,N_1436,N_3714);
nand U7501 (N_7501,N_4096,N_3907);
nand U7502 (N_7502,N_4996,N_4868);
and U7503 (N_7503,N_3968,N_4019);
nand U7504 (N_7504,N_4224,N_369);
or U7505 (N_7505,N_1643,N_1649);
nand U7506 (N_7506,N_3906,N_4701);
nand U7507 (N_7507,N_2659,N_3910);
nor U7508 (N_7508,N_4002,N_1584);
or U7509 (N_7509,N_2273,N_1841);
nand U7510 (N_7510,N_1083,N_3844);
and U7511 (N_7511,N_1800,N_4454);
nor U7512 (N_7512,N_1606,N_2801);
and U7513 (N_7513,N_2294,N_2476);
nor U7514 (N_7514,N_141,N_2797);
nor U7515 (N_7515,N_1228,N_608);
nor U7516 (N_7516,N_3432,N_2587);
nor U7517 (N_7517,N_3707,N_3243);
nand U7518 (N_7518,N_3359,N_2939);
nand U7519 (N_7519,N_3939,N_4942);
and U7520 (N_7520,N_2366,N_771);
and U7521 (N_7521,N_456,N_3394);
nand U7522 (N_7522,N_4348,N_794);
nor U7523 (N_7523,N_1447,N_4763);
and U7524 (N_7524,N_3634,N_304);
and U7525 (N_7525,N_1957,N_2953);
or U7526 (N_7526,N_2242,N_94);
nor U7527 (N_7527,N_4918,N_2481);
nand U7528 (N_7528,N_3666,N_1599);
and U7529 (N_7529,N_1085,N_2936);
nor U7530 (N_7530,N_3886,N_385);
nand U7531 (N_7531,N_2708,N_3695);
nor U7532 (N_7532,N_2364,N_4734);
nor U7533 (N_7533,N_2262,N_4495);
or U7534 (N_7534,N_3954,N_3396);
or U7535 (N_7535,N_225,N_2711);
nand U7536 (N_7536,N_625,N_2222);
or U7537 (N_7537,N_2349,N_188);
and U7538 (N_7538,N_1320,N_4988);
nor U7539 (N_7539,N_4960,N_4863);
and U7540 (N_7540,N_558,N_4578);
nand U7541 (N_7541,N_2934,N_2903);
nor U7542 (N_7542,N_1753,N_2745);
or U7543 (N_7543,N_2947,N_1953);
xnor U7544 (N_7544,N_4358,N_4952);
and U7545 (N_7545,N_4344,N_754);
or U7546 (N_7546,N_897,N_3583);
nor U7547 (N_7547,N_2740,N_1625);
nor U7548 (N_7548,N_4598,N_1997);
nor U7549 (N_7549,N_1340,N_2668);
nand U7550 (N_7550,N_2706,N_1432);
nor U7551 (N_7551,N_1315,N_2943);
nand U7552 (N_7552,N_404,N_1654);
or U7553 (N_7553,N_2641,N_3549);
and U7554 (N_7554,N_831,N_1204);
nor U7555 (N_7555,N_260,N_1528);
nor U7556 (N_7556,N_1953,N_4823);
and U7557 (N_7557,N_4442,N_4600);
or U7558 (N_7558,N_4234,N_4531);
and U7559 (N_7559,N_3289,N_1419);
or U7560 (N_7560,N_4414,N_1073);
nand U7561 (N_7561,N_4123,N_3671);
and U7562 (N_7562,N_834,N_3892);
and U7563 (N_7563,N_2769,N_4761);
and U7564 (N_7564,N_3585,N_4969);
and U7565 (N_7565,N_3343,N_2772);
or U7566 (N_7566,N_531,N_143);
nand U7567 (N_7567,N_2474,N_2235);
nor U7568 (N_7568,N_3641,N_1579);
or U7569 (N_7569,N_1472,N_197);
xnor U7570 (N_7570,N_3285,N_1767);
nor U7571 (N_7571,N_1916,N_1465);
nand U7572 (N_7572,N_4173,N_3987);
or U7573 (N_7573,N_3959,N_1318);
or U7574 (N_7574,N_2906,N_3102);
or U7575 (N_7575,N_2406,N_3088);
or U7576 (N_7576,N_2648,N_1357);
and U7577 (N_7577,N_1863,N_2332);
or U7578 (N_7578,N_4979,N_3107);
and U7579 (N_7579,N_1901,N_239);
nor U7580 (N_7580,N_1319,N_288);
or U7581 (N_7581,N_3988,N_2535);
nand U7582 (N_7582,N_538,N_3062);
nand U7583 (N_7583,N_3734,N_2797);
nand U7584 (N_7584,N_3268,N_1344);
nand U7585 (N_7585,N_175,N_785);
nand U7586 (N_7586,N_1413,N_965);
and U7587 (N_7587,N_1839,N_1202);
and U7588 (N_7588,N_1479,N_2248);
or U7589 (N_7589,N_1690,N_1719);
or U7590 (N_7590,N_324,N_3479);
nand U7591 (N_7591,N_2085,N_3891);
xnor U7592 (N_7592,N_1880,N_1929);
and U7593 (N_7593,N_582,N_4425);
nand U7594 (N_7594,N_626,N_4985);
and U7595 (N_7595,N_4372,N_3773);
or U7596 (N_7596,N_310,N_176);
nor U7597 (N_7597,N_2809,N_2595);
nor U7598 (N_7598,N_1782,N_3182);
nand U7599 (N_7599,N_1080,N_2133);
nor U7600 (N_7600,N_316,N_3860);
or U7601 (N_7601,N_776,N_2917);
nor U7602 (N_7602,N_1020,N_945);
and U7603 (N_7603,N_3368,N_2036);
and U7604 (N_7604,N_1092,N_3602);
nand U7605 (N_7605,N_4872,N_2720);
xor U7606 (N_7606,N_1125,N_3553);
and U7607 (N_7607,N_4966,N_894);
nand U7608 (N_7608,N_554,N_92);
nor U7609 (N_7609,N_747,N_4909);
nor U7610 (N_7610,N_1973,N_4185);
and U7611 (N_7611,N_2792,N_722);
nand U7612 (N_7612,N_2099,N_2871);
nor U7613 (N_7613,N_4041,N_4730);
or U7614 (N_7614,N_2766,N_1089);
nor U7615 (N_7615,N_1325,N_1699);
and U7616 (N_7616,N_423,N_1608);
nand U7617 (N_7617,N_4114,N_4889);
nand U7618 (N_7618,N_1282,N_114);
nor U7619 (N_7619,N_2502,N_1432);
and U7620 (N_7620,N_4530,N_2184);
nor U7621 (N_7621,N_4033,N_806);
nor U7622 (N_7622,N_2073,N_1658);
nor U7623 (N_7623,N_2702,N_1145);
or U7624 (N_7624,N_2946,N_925);
and U7625 (N_7625,N_27,N_4884);
nor U7626 (N_7626,N_2114,N_2590);
nor U7627 (N_7627,N_3346,N_4989);
or U7628 (N_7628,N_1515,N_2555);
nor U7629 (N_7629,N_1903,N_2728);
or U7630 (N_7630,N_3656,N_1373);
nand U7631 (N_7631,N_2375,N_2148);
nand U7632 (N_7632,N_2166,N_4502);
nor U7633 (N_7633,N_4038,N_1305);
and U7634 (N_7634,N_4884,N_3792);
or U7635 (N_7635,N_2251,N_3521);
or U7636 (N_7636,N_2754,N_2509);
or U7637 (N_7637,N_4789,N_4803);
xor U7638 (N_7638,N_1957,N_1899);
or U7639 (N_7639,N_3317,N_4992);
nor U7640 (N_7640,N_752,N_3536);
nor U7641 (N_7641,N_2794,N_3333);
nand U7642 (N_7642,N_4369,N_1777);
or U7643 (N_7643,N_4686,N_2213);
and U7644 (N_7644,N_3493,N_2831);
or U7645 (N_7645,N_4882,N_246);
nand U7646 (N_7646,N_4371,N_3185);
nand U7647 (N_7647,N_118,N_543);
nand U7648 (N_7648,N_1383,N_1837);
nor U7649 (N_7649,N_2525,N_3236);
and U7650 (N_7650,N_2359,N_138);
or U7651 (N_7651,N_4713,N_375);
nand U7652 (N_7652,N_556,N_414);
and U7653 (N_7653,N_1826,N_4289);
nand U7654 (N_7654,N_1419,N_317);
nand U7655 (N_7655,N_817,N_2862);
or U7656 (N_7656,N_1219,N_872);
or U7657 (N_7657,N_4522,N_2983);
nand U7658 (N_7658,N_3959,N_1217);
nor U7659 (N_7659,N_3689,N_1704);
nand U7660 (N_7660,N_161,N_1803);
and U7661 (N_7661,N_1808,N_911);
nor U7662 (N_7662,N_2891,N_1259);
and U7663 (N_7663,N_13,N_3842);
nand U7664 (N_7664,N_3923,N_1597);
nor U7665 (N_7665,N_3199,N_3027);
nand U7666 (N_7666,N_4439,N_2048);
or U7667 (N_7667,N_1179,N_2793);
nand U7668 (N_7668,N_4616,N_1918);
and U7669 (N_7669,N_4640,N_4538);
or U7670 (N_7670,N_3613,N_1412);
nand U7671 (N_7671,N_2170,N_2696);
and U7672 (N_7672,N_1110,N_1757);
and U7673 (N_7673,N_4687,N_1116);
xor U7674 (N_7674,N_1325,N_4408);
xnor U7675 (N_7675,N_1738,N_4485);
nor U7676 (N_7676,N_466,N_2007);
nor U7677 (N_7677,N_3745,N_3848);
xor U7678 (N_7678,N_8,N_3427);
nand U7679 (N_7679,N_2096,N_3890);
nand U7680 (N_7680,N_2666,N_3555);
nor U7681 (N_7681,N_3437,N_4658);
nand U7682 (N_7682,N_1266,N_2545);
and U7683 (N_7683,N_4432,N_1383);
nand U7684 (N_7684,N_636,N_1801);
nor U7685 (N_7685,N_4465,N_4340);
nand U7686 (N_7686,N_868,N_4129);
nand U7687 (N_7687,N_1877,N_1485);
nor U7688 (N_7688,N_3528,N_3389);
or U7689 (N_7689,N_1424,N_4624);
nand U7690 (N_7690,N_2384,N_671);
and U7691 (N_7691,N_4855,N_4427);
nand U7692 (N_7692,N_4089,N_1696);
nand U7693 (N_7693,N_3668,N_2931);
or U7694 (N_7694,N_2695,N_593);
and U7695 (N_7695,N_495,N_3066);
nor U7696 (N_7696,N_3379,N_4694);
nor U7697 (N_7697,N_3049,N_4532);
and U7698 (N_7698,N_922,N_3639);
nand U7699 (N_7699,N_1101,N_54);
nor U7700 (N_7700,N_3335,N_2083);
nand U7701 (N_7701,N_3900,N_1728);
nor U7702 (N_7702,N_124,N_954);
nor U7703 (N_7703,N_3622,N_1222);
nand U7704 (N_7704,N_4000,N_3848);
and U7705 (N_7705,N_314,N_3121);
or U7706 (N_7706,N_4387,N_2701);
and U7707 (N_7707,N_1230,N_666);
or U7708 (N_7708,N_628,N_3361);
nor U7709 (N_7709,N_192,N_3474);
and U7710 (N_7710,N_4476,N_1391);
nand U7711 (N_7711,N_4247,N_3304);
or U7712 (N_7712,N_1814,N_3664);
or U7713 (N_7713,N_4138,N_4559);
nor U7714 (N_7714,N_1245,N_139);
nor U7715 (N_7715,N_2611,N_2692);
or U7716 (N_7716,N_2633,N_1521);
or U7717 (N_7717,N_680,N_4559);
nor U7718 (N_7718,N_3152,N_4564);
and U7719 (N_7719,N_266,N_2589);
or U7720 (N_7720,N_1375,N_2076);
or U7721 (N_7721,N_4512,N_48);
and U7722 (N_7722,N_248,N_4387);
and U7723 (N_7723,N_4652,N_4751);
and U7724 (N_7724,N_1178,N_2892);
or U7725 (N_7725,N_1006,N_4947);
and U7726 (N_7726,N_4953,N_80);
and U7727 (N_7727,N_1794,N_4198);
and U7728 (N_7728,N_857,N_2643);
nor U7729 (N_7729,N_3315,N_4063);
or U7730 (N_7730,N_91,N_2997);
and U7731 (N_7731,N_1142,N_4301);
nand U7732 (N_7732,N_3049,N_4475);
or U7733 (N_7733,N_34,N_445);
or U7734 (N_7734,N_3046,N_864);
or U7735 (N_7735,N_4752,N_772);
and U7736 (N_7736,N_3222,N_683);
nand U7737 (N_7737,N_844,N_3871);
or U7738 (N_7738,N_3135,N_2016);
and U7739 (N_7739,N_3724,N_1210);
or U7740 (N_7740,N_3330,N_4212);
or U7741 (N_7741,N_1675,N_1301);
nand U7742 (N_7742,N_1706,N_2759);
or U7743 (N_7743,N_4946,N_2889);
or U7744 (N_7744,N_2280,N_4343);
nand U7745 (N_7745,N_4182,N_4808);
and U7746 (N_7746,N_4283,N_3497);
nand U7747 (N_7747,N_427,N_3765);
and U7748 (N_7748,N_684,N_4887);
nand U7749 (N_7749,N_1021,N_3733);
nand U7750 (N_7750,N_881,N_186);
or U7751 (N_7751,N_2397,N_3415);
nor U7752 (N_7752,N_1446,N_3369);
or U7753 (N_7753,N_1764,N_1564);
nor U7754 (N_7754,N_2511,N_1688);
or U7755 (N_7755,N_4919,N_2869);
and U7756 (N_7756,N_302,N_293);
nand U7757 (N_7757,N_4802,N_534);
nand U7758 (N_7758,N_2166,N_1642);
or U7759 (N_7759,N_4782,N_3794);
nor U7760 (N_7760,N_3,N_2002);
and U7761 (N_7761,N_2434,N_1357);
nor U7762 (N_7762,N_458,N_2469);
nand U7763 (N_7763,N_3170,N_4652);
nor U7764 (N_7764,N_357,N_1118);
or U7765 (N_7765,N_3115,N_2420);
nand U7766 (N_7766,N_1473,N_2111);
nand U7767 (N_7767,N_3080,N_2104);
xor U7768 (N_7768,N_2512,N_2134);
or U7769 (N_7769,N_1823,N_642);
and U7770 (N_7770,N_961,N_3586);
nand U7771 (N_7771,N_4087,N_653);
or U7772 (N_7772,N_4355,N_662);
nand U7773 (N_7773,N_188,N_475);
xnor U7774 (N_7774,N_133,N_4407);
nor U7775 (N_7775,N_1208,N_4876);
nand U7776 (N_7776,N_1229,N_196);
nor U7777 (N_7777,N_272,N_3452);
nor U7778 (N_7778,N_3008,N_4111);
nand U7779 (N_7779,N_1148,N_1328);
nor U7780 (N_7780,N_564,N_1294);
nor U7781 (N_7781,N_3309,N_611);
nand U7782 (N_7782,N_1943,N_1975);
nand U7783 (N_7783,N_2927,N_4718);
or U7784 (N_7784,N_1602,N_4978);
nor U7785 (N_7785,N_1747,N_3669);
nor U7786 (N_7786,N_2474,N_664);
nor U7787 (N_7787,N_3502,N_1394);
nor U7788 (N_7788,N_1389,N_4066);
nand U7789 (N_7789,N_3352,N_1116);
nand U7790 (N_7790,N_1235,N_653);
nor U7791 (N_7791,N_4216,N_4009);
xor U7792 (N_7792,N_1607,N_860);
or U7793 (N_7793,N_3200,N_1633);
or U7794 (N_7794,N_3915,N_4906);
and U7795 (N_7795,N_1013,N_2190);
or U7796 (N_7796,N_4621,N_4430);
or U7797 (N_7797,N_1518,N_718);
and U7798 (N_7798,N_4412,N_4432);
nand U7799 (N_7799,N_4294,N_812);
or U7800 (N_7800,N_4105,N_1520);
and U7801 (N_7801,N_1283,N_4307);
nor U7802 (N_7802,N_1244,N_1387);
nand U7803 (N_7803,N_1135,N_1389);
and U7804 (N_7804,N_1822,N_4521);
nand U7805 (N_7805,N_1051,N_4511);
and U7806 (N_7806,N_2396,N_3806);
and U7807 (N_7807,N_634,N_2199);
or U7808 (N_7808,N_1397,N_108);
nor U7809 (N_7809,N_1688,N_2703);
and U7810 (N_7810,N_2898,N_3943);
nor U7811 (N_7811,N_3514,N_2541);
or U7812 (N_7812,N_1824,N_4204);
nand U7813 (N_7813,N_3946,N_3224);
nor U7814 (N_7814,N_634,N_1137);
nand U7815 (N_7815,N_4604,N_1710);
and U7816 (N_7816,N_2561,N_312);
and U7817 (N_7817,N_2273,N_3536);
or U7818 (N_7818,N_1913,N_3764);
nand U7819 (N_7819,N_4594,N_2048);
xor U7820 (N_7820,N_237,N_2441);
nand U7821 (N_7821,N_3069,N_3122);
nor U7822 (N_7822,N_3388,N_4151);
or U7823 (N_7823,N_4792,N_2780);
or U7824 (N_7824,N_4416,N_3626);
and U7825 (N_7825,N_541,N_539);
nand U7826 (N_7826,N_328,N_1187);
or U7827 (N_7827,N_1251,N_137);
and U7828 (N_7828,N_2364,N_3738);
nor U7829 (N_7829,N_707,N_1330);
and U7830 (N_7830,N_1844,N_1763);
nor U7831 (N_7831,N_373,N_4187);
or U7832 (N_7832,N_336,N_4811);
nand U7833 (N_7833,N_3587,N_1214);
nand U7834 (N_7834,N_2580,N_3687);
nor U7835 (N_7835,N_4376,N_1521);
and U7836 (N_7836,N_4065,N_3681);
and U7837 (N_7837,N_438,N_3077);
and U7838 (N_7838,N_141,N_4501);
nand U7839 (N_7839,N_875,N_1541);
nor U7840 (N_7840,N_1284,N_3624);
and U7841 (N_7841,N_4104,N_3785);
or U7842 (N_7842,N_1454,N_1681);
and U7843 (N_7843,N_4730,N_1081);
nor U7844 (N_7844,N_3553,N_2233);
nand U7845 (N_7845,N_2959,N_698);
and U7846 (N_7846,N_62,N_496);
nor U7847 (N_7847,N_2801,N_1466);
nor U7848 (N_7848,N_1121,N_4986);
nand U7849 (N_7849,N_2939,N_973);
and U7850 (N_7850,N_4472,N_4342);
and U7851 (N_7851,N_4035,N_4022);
nand U7852 (N_7852,N_1547,N_756);
nor U7853 (N_7853,N_888,N_2116);
nand U7854 (N_7854,N_3447,N_3375);
xnor U7855 (N_7855,N_2838,N_2791);
or U7856 (N_7856,N_1624,N_1070);
or U7857 (N_7857,N_2208,N_248);
and U7858 (N_7858,N_1302,N_4244);
nand U7859 (N_7859,N_53,N_3748);
and U7860 (N_7860,N_4963,N_1437);
xnor U7861 (N_7861,N_4906,N_3640);
nor U7862 (N_7862,N_2932,N_1944);
nor U7863 (N_7863,N_3712,N_3547);
nor U7864 (N_7864,N_3014,N_3548);
nor U7865 (N_7865,N_83,N_1072);
nor U7866 (N_7866,N_1882,N_948);
nor U7867 (N_7867,N_4669,N_901);
nand U7868 (N_7868,N_1805,N_3221);
and U7869 (N_7869,N_497,N_3556);
nor U7870 (N_7870,N_2093,N_798);
nand U7871 (N_7871,N_77,N_3592);
xor U7872 (N_7872,N_2766,N_3751);
or U7873 (N_7873,N_2887,N_1283);
or U7874 (N_7874,N_323,N_696);
nand U7875 (N_7875,N_196,N_2095);
xor U7876 (N_7876,N_2864,N_2300);
nor U7877 (N_7877,N_4553,N_954);
nor U7878 (N_7878,N_891,N_3896);
or U7879 (N_7879,N_1819,N_246);
and U7880 (N_7880,N_232,N_695);
nand U7881 (N_7881,N_3033,N_3749);
nor U7882 (N_7882,N_1307,N_3974);
nor U7883 (N_7883,N_2130,N_2255);
or U7884 (N_7884,N_3172,N_4203);
nor U7885 (N_7885,N_1644,N_3357);
nor U7886 (N_7886,N_1900,N_2664);
nor U7887 (N_7887,N_3226,N_4788);
nand U7888 (N_7888,N_1207,N_1820);
or U7889 (N_7889,N_4231,N_3048);
or U7890 (N_7890,N_2969,N_2852);
or U7891 (N_7891,N_4968,N_4090);
xor U7892 (N_7892,N_1363,N_2593);
or U7893 (N_7893,N_779,N_3431);
nor U7894 (N_7894,N_4443,N_394);
or U7895 (N_7895,N_3456,N_2162);
nand U7896 (N_7896,N_1576,N_546);
and U7897 (N_7897,N_3796,N_948);
or U7898 (N_7898,N_247,N_2597);
and U7899 (N_7899,N_583,N_2466);
xor U7900 (N_7900,N_4898,N_158);
nor U7901 (N_7901,N_4653,N_1125);
and U7902 (N_7902,N_3589,N_295);
nor U7903 (N_7903,N_3125,N_4722);
nor U7904 (N_7904,N_2622,N_1352);
nand U7905 (N_7905,N_1896,N_3762);
or U7906 (N_7906,N_1593,N_3631);
and U7907 (N_7907,N_3020,N_1563);
and U7908 (N_7908,N_441,N_3611);
nor U7909 (N_7909,N_4683,N_2970);
or U7910 (N_7910,N_3778,N_387);
or U7911 (N_7911,N_3722,N_308);
nand U7912 (N_7912,N_3077,N_840);
nor U7913 (N_7913,N_992,N_2210);
or U7914 (N_7914,N_2843,N_3006);
nor U7915 (N_7915,N_1543,N_3955);
nor U7916 (N_7916,N_4777,N_2001);
nor U7917 (N_7917,N_1429,N_3074);
nor U7918 (N_7918,N_1751,N_4497);
nand U7919 (N_7919,N_2197,N_157);
xor U7920 (N_7920,N_839,N_96);
or U7921 (N_7921,N_3364,N_3842);
nand U7922 (N_7922,N_1358,N_2037);
or U7923 (N_7923,N_408,N_246);
nor U7924 (N_7924,N_4862,N_3334);
or U7925 (N_7925,N_279,N_985);
and U7926 (N_7926,N_2714,N_4819);
nor U7927 (N_7927,N_2734,N_297);
nor U7928 (N_7928,N_1474,N_2678);
or U7929 (N_7929,N_1585,N_200);
or U7930 (N_7930,N_513,N_1212);
and U7931 (N_7931,N_4053,N_3470);
xnor U7932 (N_7932,N_44,N_2169);
and U7933 (N_7933,N_4104,N_2960);
or U7934 (N_7934,N_1036,N_1192);
or U7935 (N_7935,N_2813,N_4394);
nand U7936 (N_7936,N_954,N_3299);
nand U7937 (N_7937,N_2672,N_4717);
nor U7938 (N_7938,N_2423,N_1185);
and U7939 (N_7939,N_243,N_4063);
or U7940 (N_7940,N_658,N_2058);
nor U7941 (N_7941,N_3138,N_2524);
and U7942 (N_7942,N_2796,N_4574);
or U7943 (N_7943,N_4151,N_2346);
nor U7944 (N_7944,N_3885,N_2136);
or U7945 (N_7945,N_1749,N_4876);
nor U7946 (N_7946,N_2607,N_1775);
nor U7947 (N_7947,N_507,N_1362);
xor U7948 (N_7948,N_3409,N_1272);
nand U7949 (N_7949,N_325,N_4443);
nand U7950 (N_7950,N_3689,N_2992);
nand U7951 (N_7951,N_2864,N_192);
nor U7952 (N_7952,N_1010,N_2512);
nand U7953 (N_7953,N_3133,N_744);
nand U7954 (N_7954,N_3455,N_4362);
and U7955 (N_7955,N_4745,N_2866);
or U7956 (N_7956,N_4299,N_483);
and U7957 (N_7957,N_636,N_1080);
or U7958 (N_7958,N_742,N_3560);
and U7959 (N_7959,N_1239,N_3134);
nand U7960 (N_7960,N_2061,N_3147);
or U7961 (N_7961,N_2363,N_284);
nand U7962 (N_7962,N_4106,N_1185);
and U7963 (N_7963,N_987,N_3107);
or U7964 (N_7964,N_3750,N_4273);
and U7965 (N_7965,N_919,N_1145);
or U7966 (N_7966,N_4933,N_1914);
nor U7967 (N_7967,N_2553,N_2530);
and U7968 (N_7968,N_3369,N_4699);
or U7969 (N_7969,N_3514,N_2721);
and U7970 (N_7970,N_2159,N_674);
or U7971 (N_7971,N_3465,N_2682);
or U7972 (N_7972,N_3066,N_4788);
nand U7973 (N_7973,N_1634,N_1268);
and U7974 (N_7974,N_158,N_4885);
and U7975 (N_7975,N_3114,N_2925);
and U7976 (N_7976,N_1442,N_533);
and U7977 (N_7977,N_1013,N_3916);
nand U7978 (N_7978,N_4631,N_1574);
and U7979 (N_7979,N_3671,N_540);
nand U7980 (N_7980,N_4559,N_685);
and U7981 (N_7981,N_4964,N_2148);
nand U7982 (N_7982,N_4065,N_2276);
nand U7983 (N_7983,N_4168,N_3790);
and U7984 (N_7984,N_1860,N_1378);
or U7985 (N_7985,N_606,N_680);
or U7986 (N_7986,N_848,N_4276);
or U7987 (N_7987,N_2321,N_4932);
nand U7988 (N_7988,N_973,N_1230);
nand U7989 (N_7989,N_726,N_3872);
nor U7990 (N_7990,N_2719,N_3378);
nor U7991 (N_7991,N_2379,N_1738);
nor U7992 (N_7992,N_4727,N_1010);
and U7993 (N_7993,N_3538,N_1236);
nand U7994 (N_7994,N_3487,N_427);
nand U7995 (N_7995,N_4788,N_1796);
xor U7996 (N_7996,N_558,N_4816);
xor U7997 (N_7997,N_2306,N_3325);
nand U7998 (N_7998,N_3943,N_3181);
nor U7999 (N_7999,N_3763,N_3684);
nand U8000 (N_8000,N_2947,N_4646);
nand U8001 (N_8001,N_2624,N_2810);
and U8002 (N_8002,N_1811,N_3605);
nor U8003 (N_8003,N_603,N_4585);
and U8004 (N_8004,N_1127,N_2588);
or U8005 (N_8005,N_1620,N_4388);
nor U8006 (N_8006,N_3353,N_657);
and U8007 (N_8007,N_512,N_4154);
and U8008 (N_8008,N_1648,N_3742);
nand U8009 (N_8009,N_4942,N_3053);
nor U8010 (N_8010,N_1544,N_453);
nand U8011 (N_8011,N_284,N_1160);
and U8012 (N_8012,N_4823,N_3891);
nor U8013 (N_8013,N_4454,N_468);
nor U8014 (N_8014,N_4036,N_3585);
and U8015 (N_8015,N_3555,N_1532);
nand U8016 (N_8016,N_2705,N_4199);
or U8017 (N_8017,N_1682,N_242);
and U8018 (N_8018,N_2524,N_3622);
and U8019 (N_8019,N_1566,N_3467);
nor U8020 (N_8020,N_3558,N_4674);
nand U8021 (N_8021,N_1608,N_3070);
nor U8022 (N_8022,N_1824,N_2641);
nand U8023 (N_8023,N_833,N_262);
nand U8024 (N_8024,N_4827,N_62);
and U8025 (N_8025,N_728,N_609);
nor U8026 (N_8026,N_3219,N_4201);
nand U8027 (N_8027,N_4855,N_1327);
and U8028 (N_8028,N_1822,N_2923);
nand U8029 (N_8029,N_3012,N_3818);
and U8030 (N_8030,N_1511,N_94);
and U8031 (N_8031,N_4539,N_2387);
or U8032 (N_8032,N_1974,N_3169);
nor U8033 (N_8033,N_3577,N_4099);
nand U8034 (N_8034,N_1803,N_457);
nor U8035 (N_8035,N_301,N_3792);
nor U8036 (N_8036,N_2327,N_4164);
or U8037 (N_8037,N_1300,N_3081);
nor U8038 (N_8038,N_2553,N_4377);
nand U8039 (N_8039,N_2323,N_4895);
nand U8040 (N_8040,N_2615,N_2725);
or U8041 (N_8041,N_2664,N_3332);
nor U8042 (N_8042,N_1076,N_2558);
or U8043 (N_8043,N_4939,N_3701);
nor U8044 (N_8044,N_1460,N_3439);
nand U8045 (N_8045,N_4957,N_2772);
or U8046 (N_8046,N_4021,N_1627);
nand U8047 (N_8047,N_4841,N_2850);
nor U8048 (N_8048,N_299,N_758);
nand U8049 (N_8049,N_2761,N_1616);
or U8050 (N_8050,N_2454,N_3101);
nand U8051 (N_8051,N_644,N_4086);
and U8052 (N_8052,N_3206,N_2686);
nand U8053 (N_8053,N_940,N_346);
nand U8054 (N_8054,N_4174,N_2208);
nand U8055 (N_8055,N_2580,N_4724);
or U8056 (N_8056,N_1107,N_2598);
or U8057 (N_8057,N_415,N_3031);
or U8058 (N_8058,N_1247,N_4682);
and U8059 (N_8059,N_2347,N_2994);
nand U8060 (N_8060,N_3424,N_1789);
nor U8061 (N_8061,N_1546,N_1016);
or U8062 (N_8062,N_1013,N_1698);
and U8063 (N_8063,N_4424,N_1405);
nand U8064 (N_8064,N_2611,N_344);
or U8065 (N_8065,N_2930,N_4552);
nor U8066 (N_8066,N_3610,N_4286);
and U8067 (N_8067,N_1591,N_1587);
nand U8068 (N_8068,N_818,N_3798);
nor U8069 (N_8069,N_4154,N_2074);
and U8070 (N_8070,N_3274,N_2753);
or U8071 (N_8071,N_4582,N_1515);
or U8072 (N_8072,N_4353,N_4238);
nor U8073 (N_8073,N_1499,N_2286);
nor U8074 (N_8074,N_3847,N_3575);
and U8075 (N_8075,N_1676,N_267);
and U8076 (N_8076,N_486,N_2023);
nor U8077 (N_8077,N_3969,N_2706);
and U8078 (N_8078,N_1767,N_4421);
nand U8079 (N_8079,N_2060,N_4315);
nand U8080 (N_8080,N_2555,N_1708);
nand U8081 (N_8081,N_661,N_3339);
and U8082 (N_8082,N_4284,N_3501);
nor U8083 (N_8083,N_2039,N_2779);
or U8084 (N_8084,N_1613,N_3399);
nand U8085 (N_8085,N_2392,N_3775);
nor U8086 (N_8086,N_2038,N_2990);
or U8087 (N_8087,N_1614,N_875);
nor U8088 (N_8088,N_2970,N_4492);
and U8089 (N_8089,N_4600,N_1622);
xor U8090 (N_8090,N_1053,N_2254);
nand U8091 (N_8091,N_1349,N_1035);
or U8092 (N_8092,N_777,N_3853);
or U8093 (N_8093,N_1905,N_4043);
nor U8094 (N_8094,N_4441,N_459);
nor U8095 (N_8095,N_2726,N_2551);
nand U8096 (N_8096,N_3383,N_4008);
or U8097 (N_8097,N_2721,N_4479);
nor U8098 (N_8098,N_3679,N_1023);
nand U8099 (N_8099,N_3615,N_4158);
or U8100 (N_8100,N_4253,N_4189);
or U8101 (N_8101,N_2297,N_2889);
nor U8102 (N_8102,N_2952,N_4531);
and U8103 (N_8103,N_3260,N_2178);
or U8104 (N_8104,N_1298,N_3015);
nor U8105 (N_8105,N_3020,N_4128);
or U8106 (N_8106,N_827,N_2367);
nand U8107 (N_8107,N_3908,N_2199);
and U8108 (N_8108,N_4156,N_3603);
nor U8109 (N_8109,N_1967,N_1746);
nand U8110 (N_8110,N_1951,N_1693);
or U8111 (N_8111,N_3794,N_4026);
nor U8112 (N_8112,N_2672,N_4654);
or U8113 (N_8113,N_249,N_925);
nor U8114 (N_8114,N_864,N_1161);
or U8115 (N_8115,N_4481,N_3754);
or U8116 (N_8116,N_3182,N_204);
nand U8117 (N_8117,N_2573,N_4903);
nand U8118 (N_8118,N_579,N_170);
or U8119 (N_8119,N_1279,N_2801);
nand U8120 (N_8120,N_1778,N_4515);
or U8121 (N_8121,N_1209,N_2585);
and U8122 (N_8122,N_4624,N_1215);
and U8123 (N_8123,N_2795,N_2001);
nand U8124 (N_8124,N_487,N_506);
nor U8125 (N_8125,N_4666,N_3128);
and U8126 (N_8126,N_4933,N_1207);
or U8127 (N_8127,N_716,N_4706);
nor U8128 (N_8128,N_2739,N_1740);
nand U8129 (N_8129,N_4068,N_3887);
and U8130 (N_8130,N_1532,N_2163);
and U8131 (N_8131,N_4332,N_2913);
nor U8132 (N_8132,N_4171,N_2306);
nor U8133 (N_8133,N_65,N_1957);
nor U8134 (N_8134,N_1399,N_1778);
and U8135 (N_8135,N_3835,N_2021);
nand U8136 (N_8136,N_3159,N_1867);
or U8137 (N_8137,N_2858,N_2370);
or U8138 (N_8138,N_2071,N_3946);
and U8139 (N_8139,N_4766,N_1784);
and U8140 (N_8140,N_3726,N_2708);
nor U8141 (N_8141,N_1724,N_309);
nor U8142 (N_8142,N_2549,N_718);
nand U8143 (N_8143,N_1783,N_1217);
nor U8144 (N_8144,N_4359,N_4736);
nor U8145 (N_8145,N_742,N_1649);
nand U8146 (N_8146,N_3779,N_321);
and U8147 (N_8147,N_3242,N_3474);
or U8148 (N_8148,N_4009,N_31);
nor U8149 (N_8149,N_1212,N_929);
or U8150 (N_8150,N_4849,N_1236);
or U8151 (N_8151,N_837,N_4304);
nor U8152 (N_8152,N_2648,N_4866);
or U8153 (N_8153,N_9,N_4223);
nand U8154 (N_8154,N_2988,N_4527);
or U8155 (N_8155,N_2178,N_3737);
or U8156 (N_8156,N_149,N_3660);
xor U8157 (N_8157,N_440,N_1491);
nor U8158 (N_8158,N_4577,N_3181);
and U8159 (N_8159,N_4574,N_95);
nor U8160 (N_8160,N_2961,N_1141);
or U8161 (N_8161,N_4528,N_369);
and U8162 (N_8162,N_2119,N_235);
or U8163 (N_8163,N_2872,N_2156);
and U8164 (N_8164,N_3181,N_4165);
nand U8165 (N_8165,N_2697,N_2885);
or U8166 (N_8166,N_2955,N_1968);
nand U8167 (N_8167,N_3411,N_1191);
nor U8168 (N_8168,N_950,N_2243);
nand U8169 (N_8169,N_2340,N_2409);
nand U8170 (N_8170,N_575,N_1535);
nor U8171 (N_8171,N_1774,N_4405);
and U8172 (N_8172,N_52,N_3952);
or U8173 (N_8173,N_4454,N_4916);
or U8174 (N_8174,N_3242,N_752);
and U8175 (N_8175,N_109,N_650);
and U8176 (N_8176,N_285,N_428);
or U8177 (N_8177,N_3097,N_3752);
nand U8178 (N_8178,N_150,N_3743);
or U8179 (N_8179,N_1916,N_750);
nor U8180 (N_8180,N_4506,N_2840);
nand U8181 (N_8181,N_3569,N_4608);
nor U8182 (N_8182,N_3886,N_4595);
or U8183 (N_8183,N_3800,N_4298);
and U8184 (N_8184,N_3058,N_298);
or U8185 (N_8185,N_3752,N_4703);
nand U8186 (N_8186,N_4632,N_2269);
nor U8187 (N_8187,N_204,N_2028);
or U8188 (N_8188,N_1472,N_2123);
and U8189 (N_8189,N_2912,N_4756);
nor U8190 (N_8190,N_2020,N_1312);
nor U8191 (N_8191,N_1212,N_1702);
or U8192 (N_8192,N_4865,N_1178);
nor U8193 (N_8193,N_3352,N_3696);
nor U8194 (N_8194,N_4396,N_4266);
nand U8195 (N_8195,N_2099,N_1452);
or U8196 (N_8196,N_283,N_217);
nand U8197 (N_8197,N_4364,N_3266);
nor U8198 (N_8198,N_1961,N_3524);
nand U8199 (N_8199,N_1526,N_1901);
and U8200 (N_8200,N_4406,N_1495);
or U8201 (N_8201,N_3296,N_2654);
or U8202 (N_8202,N_541,N_2071);
and U8203 (N_8203,N_2474,N_1211);
nand U8204 (N_8204,N_3753,N_694);
and U8205 (N_8205,N_673,N_686);
nand U8206 (N_8206,N_4358,N_4444);
xor U8207 (N_8207,N_967,N_3181);
nor U8208 (N_8208,N_2588,N_1277);
nor U8209 (N_8209,N_4066,N_4030);
nor U8210 (N_8210,N_560,N_2411);
xor U8211 (N_8211,N_1144,N_1621);
and U8212 (N_8212,N_1013,N_1507);
or U8213 (N_8213,N_1230,N_757);
or U8214 (N_8214,N_3824,N_1519);
nor U8215 (N_8215,N_4936,N_1246);
or U8216 (N_8216,N_2543,N_2650);
or U8217 (N_8217,N_4568,N_2095);
nor U8218 (N_8218,N_3845,N_2824);
nand U8219 (N_8219,N_984,N_436);
nand U8220 (N_8220,N_4488,N_3868);
and U8221 (N_8221,N_3516,N_849);
nor U8222 (N_8222,N_1217,N_1880);
nand U8223 (N_8223,N_2085,N_1636);
or U8224 (N_8224,N_4631,N_3151);
nand U8225 (N_8225,N_2419,N_3901);
or U8226 (N_8226,N_3096,N_775);
and U8227 (N_8227,N_2352,N_2319);
or U8228 (N_8228,N_579,N_3289);
nor U8229 (N_8229,N_131,N_3408);
nand U8230 (N_8230,N_2025,N_3853);
nor U8231 (N_8231,N_4939,N_281);
or U8232 (N_8232,N_2347,N_4884);
nor U8233 (N_8233,N_4970,N_513);
nand U8234 (N_8234,N_1441,N_3975);
nor U8235 (N_8235,N_1247,N_4061);
nand U8236 (N_8236,N_3512,N_2631);
or U8237 (N_8237,N_3302,N_3769);
or U8238 (N_8238,N_402,N_4165);
or U8239 (N_8239,N_4129,N_2755);
nand U8240 (N_8240,N_4451,N_2734);
or U8241 (N_8241,N_3807,N_518);
nand U8242 (N_8242,N_704,N_438);
nand U8243 (N_8243,N_2429,N_2111);
and U8244 (N_8244,N_1786,N_145);
nand U8245 (N_8245,N_2959,N_3877);
or U8246 (N_8246,N_2746,N_2502);
nor U8247 (N_8247,N_2226,N_4423);
and U8248 (N_8248,N_4873,N_4609);
xnor U8249 (N_8249,N_4934,N_3857);
nor U8250 (N_8250,N_4347,N_47);
nor U8251 (N_8251,N_211,N_4233);
or U8252 (N_8252,N_2356,N_100);
xor U8253 (N_8253,N_960,N_170);
and U8254 (N_8254,N_4434,N_230);
and U8255 (N_8255,N_3665,N_1129);
or U8256 (N_8256,N_1536,N_740);
and U8257 (N_8257,N_203,N_1092);
nand U8258 (N_8258,N_3314,N_4598);
nor U8259 (N_8259,N_1678,N_759);
nor U8260 (N_8260,N_1278,N_934);
nor U8261 (N_8261,N_3687,N_362);
nand U8262 (N_8262,N_4545,N_4712);
and U8263 (N_8263,N_1854,N_4290);
and U8264 (N_8264,N_3678,N_4109);
nor U8265 (N_8265,N_4257,N_3720);
and U8266 (N_8266,N_2678,N_2889);
and U8267 (N_8267,N_4967,N_2909);
nand U8268 (N_8268,N_1153,N_3772);
nor U8269 (N_8269,N_2877,N_1933);
nand U8270 (N_8270,N_1730,N_1254);
or U8271 (N_8271,N_340,N_3988);
xnor U8272 (N_8272,N_1908,N_4122);
and U8273 (N_8273,N_4630,N_1757);
and U8274 (N_8274,N_3948,N_921);
or U8275 (N_8275,N_4820,N_3323);
nor U8276 (N_8276,N_3967,N_579);
or U8277 (N_8277,N_2436,N_2934);
or U8278 (N_8278,N_1174,N_2532);
nand U8279 (N_8279,N_2657,N_3437);
nor U8280 (N_8280,N_3197,N_3092);
nor U8281 (N_8281,N_3573,N_2986);
nor U8282 (N_8282,N_201,N_3613);
nand U8283 (N_8283,N_3952,N_1306);
or U8284 (N_8284,N_4743,N_2333);
and U8285 (N_8285,N_3660,N_2930);
and U8286 (N_8286,N_4415,N_3598);
nor U8287 (N_8287,N_3469,N_3162);
and U8288 (N_8288,N_2571,N_1549);
and U8289 (N_8289,N_2888,N_4918);
and U8290 (N_8290,N_2414,N_1182);
nor U8291 (N_8291,N_2618,N_3501);
nand U8292 (N_8292,N_4579,N_723);
or U8293 (N_8293,N_587,N_1824);
xnor U8294 (N_8294,N_3445,N_3675);
nand U8295 (N_8295,N_1643,N_3601);
and U8296 (N_8296,N_4102,N_1179);
and U8297 (N_8297,N_3580,N_4853);
and U8298 (N_8298,N_2501,N_1445);
nor U8299 (N_8299,N_4340,N_2343);
nand U8300 (N_8300,N_1168,N_2036);
or U8301 (N_8301,N_2764,N_2679);
and U8302 (N_8302,N_2853,N_4240);
and U8303 (N_8303,N_1784,N_3348);
and U8304 (N_8304,N_1643,N_645);
or U8305 (N_8305,N_3997,N_1205);
and U8306 (N_8306,N_3132,N_4524);
or U8307 (N_8307,N_3616,N_3192);
or U8308 (N_8308,N_716,N_1640);
nor U8309 (N_8309,N_527,N_2433);
and U8310 (N_8310,N_2995,N_2610);
and U8311 (N_8311,N_2376,N_4947);
nor U8312 (N_8312,N_165,N_2287);
nand U8313 (N_8313,N_751,N_2922);
and U8314 (N_8314,N_2006,N_844);
or U8315 (N_8315,N_4179,N_527);
nand U8316 (N_8316,N_2902,N_1777);
nand U8317 (N_8317,N_4908,N_3860);
nor U8318 (N_8318,N_310,N_2968);
or U8319 (N_8319,N_187,N_2149);
nor U8320 (N_8320,N_3379,N_212);
nand U8321 (N_8321,N_1827,N_352);
and U8322 (N_8322,N_2074,N_1553);
nand U8323 (N_8323,N_1904,N_4249);
nor U8324 (N_8324,N_3082,N_4476);
nand U8325 (N_8325,N_1062,N_3417);
nand U8326 (N_8326,N_4314,N_2504);
or U8327 (N_8327,N_3341,N_2420);
nor U8328 (N_8328,N_3940,N_2475);
nand U8329 (N_8329,N_4352,N_3098);
nand U8330 (N_8330,N_4281,N_1822);
and U8331 (N_8331,N_534,N_3044);
nand U8332 (N_8332,N_1811,N_790);
and U8333 (N_8333,N_3962,N_1731);
nand U8334 (N_8334,N_2504,N_1351);
nor U8335 (N_8335,N_3903,N_70);
or U8336 (N_8336,N_1847,N_444);
nand U8337 (N_8337,N_2896,N_2892);
nor U8338 (N_8338,N_1881,N_2589);
and U8339 (N_8339,N_2675,N_4698);
nand U8340 (N_8340,N_545,N_3214);
and U8341 (N_8341,N_2917,N_1501);
nor U8342 (N_8342,N_2171,N_3709);
xor U8343 (N_8343,N_2893,N_2419);
nand U8344 (N_8344,N_728,N_3615);
nor U8345 (N_8345,N_222,N_3998);
nor U8346 (N_8346,N_2527,N_2970);
nand U8347 (N_8347,N_2281,N_4717);
or U8348 (N_8348,N_1693,N_3833);
and U8349 (N_8349,N_3957,N_872);
and U8350 (N_8350,N_4786,N_1889);
xnor U8351 (N_8351,N_716,N_387);
nand U8352 (N_8352,N_989,N_3262);
nor U8353 (N_8353,N_2816,N_3836);
and U8354 (N_8354,N_1814,N_1944);
or U8355 (N_8355,N_4773,N_4581);
or U8356 (N_8356,N_2009,N_1955);
and U8357 (N_8357,N_297,N_3169);
or U8358 (N_8358,N_1951,N_3042);
or U8359 (N_8359,N_4134,N_3369);
or U8360 (N_8360,N_1610,N_4140);
and U8361 (N_8361,N_3349,N_2212);
and U8362 (N_8362,N_701,N_312);
nor U8363 (N_8363,N_3267,N_2536);
nand U8364 (N_8364,N_3193,N_3018);
nand U8365 (N_8365,N_578,N_3970);
nor U8366 (N_8366,N_1636,N_4165);
nand U8367 (N_8367,N_4208,N_608);
nor U8368 (N_8368,N_2742,N_3134);
or U8369 (N_8369,N_4232,N_3050);
nor U8370 (N_8370,N_1531,N_3760);
or U8371 (N_8371,N_1980,N_4207);
and U8372 (N_8372,N_3045,N_1521);
and U8373 (N_8373,N_4266,N_4136);
nor U8374 (N_8374,N_3033,N_49);
or U8375 (N_8375,N_3383,N_309);
nor U8376 (N_8376,N_2811,N_2329);
or U8377 (N_8377,N_2258,N_4907);
and U8378 (N_8378,N_2049,N_2988);
nand U8379 (N_8379,N_3087,N_3608);
nor U8380 (N_8380,N_4431,N_2064);
nand U8381 (N_8381,N_1808,N_975);
nand U8382 (N_8382,N_873,N_3582);
nand U8383 (N_8383,N_3990,N_1174);
or U8384 (N_8384,N_3706,N_4361);
or U8385 (N_8385,N_2144,N_4418);
or U8386 (N_8386,N_580,N_1060);
and U8387 (N_8387,N_3862,N_4745);
nand U8388 (N_8388,N_2129,N_436);
nor U8389 (N_8389,N_4844,N_2419);
nor U8390 (N_8390,N_512,N_1971);
xor U8391 (N_8391,N_1324,N_3192);
or U8392 (N_8392,N_4146,N_315);
nor U8393 (N_8393,N_1853,N_1494);
nand U8394 (N_8394,N_3095,N_1227);
nor U8395 (N_8395,N_2424,N_2227);
nor U8396 (N_8396,N_2734,N_4018);
nand U8397 (N_8397,N_4862,N_4110);
nand U8398 (N_8398,N_748,N_1937);
or U8399 (N_8399,N_944,N_1867);
nand U8400 (N_8400,N_3454,N_4069);
nor U8401 (N_8401,N_919,N_3340);
or U8402 (N_8402,N_4351,N_2398);
nand U8403 (N_8403,N_4554,N_1506);
or U8404 (N_8404,N_4038,N_1083);
and U8405 (N_8405,N_4140,N_2931);
nor U8406 (N_8406,N_349,N_491);
nor U8407 (N_8407,N_1253,N_2013);
nand U8408 (N_8408,N_3003,N_1532);
or U8409 (N_8409,N_1389,N_4877);
nor U8410 (N_8410,N_342,N_657);
or U8411 (N_8411,N_1957,N_3059);
and U8412 (N_8412,N_2960,N_143);
or U8413 (N_8413,N_186,N_1193);
nor U8414 (N_8414,N_4070,N_1178);
nor U8415 (N_8415,N_699,N_152);
nand U8416 (N_8416,N_981,N_3702);
or U8417 (N_8417,N_3112,N_3687);
and U8418 (N_8418,N_1364,N_2722);
or U8419 (N_8419,N_1283,N_929);
xnor U8420 (N_8420,N_3866,N_1869);
or U8421 (N_8421,N_1472,N_2522);
xnor U8422 (N_8422,N_1253,N_4607);
nand U8423 (N_8423,N_1253,N_4117);
nor U8424 (N_8424,N_4772,N_627);
or U8425 (N_8425,N_1492,N_1460);
and U8426 (N_8426,N_597,N_76);
nor U8427 (N_8427,N_3081,N_3397);
nand U8428 (N_8428,N_2751,N_4394);
or U8429 (N_8429,N_184,N_4800);
nand U8430 (N_8430,N_950,N_2937);
or U8431 (N_8431,N_1684,N_2073);
nand U8432 (N_8432,N_2568,N_1861);
and U8433 (N_8433,N_688,N_4812);
or U8434 (N_8434,N_4596,N_4820);
nor U8435 (N_8435,N_1115,N_1104);
or U8436 (N_8436,N_1806,N_1449);
or U8437 (N_8437,N_1726,N_1450);
nor U8438 (N_8438,N_304,N_3537);
and U8439 (N_8439,N_1274,N_532);
or U8440 (N_8440,N_1914,N_2901);
and U8441 (N_8441,N_126,N_537);
nand U8442 (N_8442,N_2663,N_441);
nor U8443 (N_8443,N_3270,N_929);
or U8444 (N_8444,N_4165,N_4128);
or U8445 (N_8445,N_3589,N_172);
or U8446 (N_8446,N_2997,N_4873);
or U8447 (N_8447,N_529,N_2711);
nand U8448 (N_8448,N_2990,N_3275);
nor U8449 (N_8449,N_3543,N_493);
nor U8450 (N_8450,N_3198,N_1312);
and U8451 (N_8451,N_1290,N_4192);
and U8452 (N_8452,N_4450,N_2530);
or U8453 (N_8453,N_4341,N_1563);
nor U8454 (N_8454,N_3835,N_635);
nor U8455 (N_8455,N_4739,N_3926);
nand U8456 (N_8456,N_615,N_4908);
and U8457 (N_8457,N_4405,N_2448);
and U8458 (N_8458,N_3612,N_493);
nor U8459 (N_8459,N_3521,N_314);
nand U8460 (N_8460,N_4460,N_2747);
and U8461 (N_8461,N_2623,N_3995);
or U8462 (N_8462,N_2759,N_2478);
nor U8463 (N_8463,N_2104,N_2802);
nand U8464 (N_8464,N_1401,N_1675);
nand U8465 (N_8465,N_1896,N_454);
or U8466 (N_8466,N_1071,N_3930);
nor U8467 (N_8467,N_563,N_3846);
nor U8468 (N_8468,N_426,N_4195);
and U8469 (N_8469,N_4480,N_3288);
or U8470 (N_8470,N_3118,N_3854);
and U8471 (N_8471,N_2380,N_919);
or U8472 (N_8472,N_1594,N_3159);
or U8473 (N_8473,N_3068,N_1960);
nand U8474 (N_8474,N_4748,N_186);
nor U8475 (N_8475,N_3907,N_3546);
nor U8476 (N_8476,N_3968,N_4417);
nand U8477 (N_8477,N_848,N_2006);
nor U8478 (N_8478,N_2204,N_2630);
or U8479 (N_8479,N_1550,N_2887);
nand U8480 (N_8480,N_2710,N_2352);
nor U8481 (N_8481,N_306,N_4132);
xnor U8482 (N_8482,N_3458,N_2520);
or U8483 (N_8483,N_4661,N_3499);
or U8484 (N_8484,N_4434,N_3986);
and U8485 (N_8485,N_1993,N_4883);
nand U8486 (N_8486,N_3836,N_4656);
nand U8487 (N_8487,N_4344,N_934);
and U8488 (N_8488,N_3922,N_4003);
or U8489 (N_8489,N_725,N_184);
or U8490 (N_8490,N_4083,N_3173);
nor U8491 (N_8491,N_4451,N_3524);
nor U8492 (N_8492,N_1308,N_3076);
or U8493 (N_8493,N_683,N_88);
and U8494 (N_8494,N_4329,N_4770);
and U8495 (N_8495,N_2621,N_113);
nor U8496 (N_8496,N_78,N_2742);
nand U8497 (N_8497,N_3280,N_4364);
nor U8498 (N_8498,N_4671,N_861);
or U8499 (N_8499,N_3407,N_1170);
or U8500 (N_8500,N_3643,N_352);
nor U8501 (N_8501,N_3266,N_2640);
nor U8502 (N_8502,N_1012,N_3570);
and U8503 (N_8503,N_1202,N_1792);
nor U8504 (N_8504,N_2716,N_999);
or U8505 (N_8505,N_3993,N_104);
or U8506 (N_8506,N_2670,N_3797);
nor U8507 (N_8507,N_882,N_3569);
or U8508 (N_8508,N_4748,N_2400);
and U8509 (N_8509,N_3818,N_1860);
or U8510 (N_8510,N_2600,N_972);
or U8511 (N_8511,N_1969,N_17);
nor U8512 (N_8512,N_2511,N_4611);
nor U8513 (N_8513,N_3309,N_3826);
nand U8514 (N_8514,N_3077,N_2318);
or U8515 (N_8515,N_3545,N_3409);
and U8516 (N_8516,N_3388,N_3399);
and U8517 (N_8517,N_497,N_3995);
and U8518 (N_8518,N_2670,N_3466);
and U8519 (N_8519,N_3412,N_4138);
nand U8520 (N_8520,N_426,N_1824);
nor U8521 (N_8521,N_1848,N_352);
nand U8522 (N_8522,N_1251,N_2001);
nor U8523 (N_8523,N_1363,N_4770);
and U8524 (N_8524,N_1080,N_4475);
and U8525 (N_8525,N_169,N_938);
nor U8526 (N_8526,N_913,N_2930);
nor U8527 (N_8527,N_740,N_3012);
nor U8528 (N_8528,N_681,N_4062);
and U8529 (N_8529,N_954,N_567);
and U8530 (N_8530,N_3025,N_3318);
or U8531 (N_8531,N_648,N_1328);
nor U8532 (N_8532,N_2710,N_263);
and U8533 (N_8533,N_3295,N_2298);
nor U8534 (N_8534,N_905,N_1194);
and U8535 (N_8535,N_4400,N_2636);
nor U8536 (N_8536,N_1680,N_3374);
or U8537 (N_8537,N_160,N_3260);
or U8538 (N_8538,N_2854,N_1513);
or U8539 (N_8539,N_99,N_3832);
or U8540 (N_8540,N_1775,N_2490);
or U8541 (N_8541,N_1894,N_2616);
or U8542 (N_8542,N_1244,N_4210);
and U8543 (N_8543,N_758,N_2314);
and U8544 (N_8544,N_3490,N_258);
nor U8545 (N_8545,N_2710,N_3646);
nand U8546 (N_8546,N_459,N_1962);
and U8547 (N_8547,N_320,N_3269);
nor U8548 (N_8548,N_3647,N_3771);
nand U8549 (N_8549,N_4778,N_2126);
or U8550 (N_8550,N_2931,N_4706);
nor U8551 (N_8551,N_1588,N_329);
and U8552 (N_8552,N_2269,N_360);
nor U8553 (N_8553,N_4377,N_1203);
or U8554 (N_8554,N_3830,N_3579);
xnor U8555 (N_8555,N_4017,N_186);
and U8556 (N_8556,N_2005,N_1474);
and U8557 (N_8557,N_4589,N_4966);
nand U8558 (N_8558,N_4854,N_3699);
or U8559 (N_8559,N_4483,N_57);
nand U8560 (N_8560,N_998,N_2351);
or U8561 (N_8561,N_876,N_2496);
or U8562 (N_8562,N_4300,N_2364);
nor U8563 (N_8563,N_1991,N_3430);
nand U8564 (N_8564,N_4908,N_3540);
or U8565 (N_8565,N_1549,N_4622);
nand U8566 (N_8566,N_3097,N_553);
and U8567 (N_8567,N_4696,N_1179);
or U8568 (N_8568,N_3792,N_1678);
nand U8569 (N_8569,N_575,N_2505);
xnor U8570 (N_8570,N_2301,N_278);
or U8571 (N_8571,N_4478,N_3066);
or U8572 (N_8572,N_2224,N_2508);
nand U8573 (N_8573,N_3167,N_3136);
nor U8574 (N_8574,N_4283,N_521);
and U8575 (N_8575,N_780,N_1252);
or U8576 (N_8576,N_900,N_3436);
nor U8577 (N_8577,N_1559,N_1156);
nand U8578 (N_8578,N_78,N_762);
and U8579 (N_8579,N_1013,N_506);
nand U8580 (N_8580,N_3386,N_303);
nand U8581 (N_8581,N_4352,N_2455);
or U8582 (N_8582,N_1858,N_485);
nor U8583 (N_8583,N_4816,N_4954);
and U8584 (N_8584,N_504,N_3358);
nand U8585 (N_8585,N_4994,N_1078);
and U8586 (N_8586,N_4077,N_4377);
nor U8587 (N_8587,N_4113,N_2029);
nand U8588 (N_8588,N_1136,N_2170);
xnor U8589 (N_8589,N_3775,N_2860);
nor U8590 (N_8590,N_858,N_1351);
and U8591 (N_8591,N_4262,N_2807);
nor U8592 (N_8592,N_457,N_3221);
and U8593 (N_8593,N_3950,N_1895);
and U8594 (N_8594,N_1376,N_3821);
and U8595 (N_8595,N_1472,N_3419);
and U8596 (N_8596,N_3101,N_842);
or U8597 (N_8597,N_2293,N_266);
nor U8598 (N_8598,N_1324,N_3390);
or U8599 (N_8599,N_1979,N_3062);
nand U8600 (N_8600,N_4041,N_156);
and U8601 (N_8601,N_1325,N_4277);
nor U8602 (N_8602,N_1918,N_1437);
and U8603 (N_8603,N_2017,N_4419);
nand U8604 (N_8604,N_583,N_4192);
nand U8605 (N_8605,N_1808,N_1898);
xor U8606 (N_8606,N_2244,N_923);
or U8607 (N_8607,N_2754,N_1944);
and U8608 (N_8608,N_4738,N_2456);
and U8609 (N_8609,N_3234,N_1107);
nor U8610 (N_8610,N_3492,N_1609);
and U8611 (N_8611,N_2007,N_2364);
or U8612 (N_8612,N_1425,N_1458);
and U8613 (N_8613,N_3144,N_4084);
or U8614 (N_8614,N_532,N_1775);
nor U8615 (N_8615,N_1283,N_4752);
nor U8616 (N_8616,N_3932,N_2533);
nand U8617 (N_8617,N_3960,N_4900);
or U8618 (N_8618,N_4151,N_3913);
nor U8619 (N_8619,N_2675,N_4019);
nor U8620 (N_8620,N_1847,N_304);
nor U8621 (N_8621,N_1170,N_2898);
or U8622 (N_8622,N_404,N_3712);
nor U8623 (N_8623,N_1748,N_684);
nor U8624 (N_8624,N_4034,N_202);
nand U8625 (N_8625,N_30,N_1777);
nand U8626 (N_8626,N_4522,N_3621);
nor U8627 (N_8627,N_3326,N_1676);
or U8628 (N_8628,N_3303,N_1947);
nand U8629 (N_8629,N_1258,N_1845);
nand U8630 (N_8630,N_258,N_2316);
nor U8631 (N_8631,N_3425,N_1338);
nand U8632 (N_8632,N_4679,N_1980);
and U8633 (N_8633,N_4278,N_4308);
and U8634 (N_8634,N_4069,N_2833);
and U8635 (N_8635,N_4574,N_2619);
and U8636 (N_8636,N_1592,N_1);
and U8637 (N_8637,N_1561,N_2338);
nand U8638 (N_8638,N_3811,N_1964);
nor U8639 (N_8639,N_4388,N_820);
nor U8640 (N_8640,N_4863,N_2443);
nor U8641 (N_8641,N_4076,N_747);
or U8642 (N_8642,N_3932,N_1434);
nor U8643 (N_8643,N_4652,N_4811);
and U8644 (N_8644,N_2555,N_4905);
nor U8645 (N_8645,N_4569,N_4536);
nand U8646 (N_8646,N_585,N_1566);
nand U8647 (N_8647,N_2837,N_20);
and U8648 (N_8648,N_3948,N_966);
nor U8649 (N_8649,N_1060,N_2403);
nor U8650 (N_8650,N_430,N_3574);
or U8651 (N_8651,N_4703,N_1751);
or U8652 (N_8652,N_4337,N_1186);
and U8653 (N_8653,N_4570,N_631);
and U8654 (N_8654,N_4036,N_4635);
and U8655 (N_8655,N_1225,N_4104);
nor U8656 (N_8656,N_3490,N_4789);
or U8657 (N_8657,N_4208,N_797);
and U8658 (N_8658,N_4551,N_2466);
nand U8659 (N_8659,N_3542,N_2750);
nor U8660 (N_8660,N_3891,N_1288);
nand U8661 (N_8661,N_3483,N_3566);
or U8662 (N_8662,N_2056,N_1278);
nand U8663 (N_8663,N_3796,N_4905);
and U8664 (N_8664,N_2674,N_1927);
nand U8665 (N_8665,N_1646,N_967);
nor U8666 (N_8666,N_1213,N_57);
nor U8667 (N_8667,N_1150,N_2271);
or U8668 (N_8668,N_259,N_2309);
nand U8669 (N_8669,N_431,N_3085);
or U8670 (N_8670,N_289,N_1527);
or U8671 (N_8671,N_1600,N_2711);
or U8672 (N_8672,N_4278,N_4084);
and U8673 (N_8673,N_3488,N_906);
nand U8674 (N_8674,N_4162,N_3269);
nand U8675 (N_8675,N_904,N_4893);
nand U8676 (N_8676,N_4935,N_1433);
nor U8677 (N_8677,N_2983,N_2729);
nand U8678 (N_8678,N_2115,N_4158);
nor U8679 (N_8679,N_828,N_1997);
and U8680 (N_8680,N_2947,N_3953);
or U8681 (N_8681,N_1333,N_311);
nand U8682 (N_8682,N_2118,N_2375);
nand U8683 (N_8683,N_2927,N_1889);
and U8684 (N_8684,N_526,N_1886);
or U8685 (N_8685,N_2933,N_2383);
nand U8686 (N_8686,N_1889,N_3811);
nor U8687 (N_8687,N_856,N_1114);
nand U8688 (N_8688,N_3793,N_4352);
nand U8689 (N_8689,N_2984,N_3535);
or U8690 (N_8690,N_1484,N_4074);
and U8691 (N_8691,N_4990,N_177);
nand U8692 (N_8692,N_4863,N_4685);
or U8693 (N_8693,N_1310,N_2420);
or U8694 (N_8694,N_4690,N_2009);
nand U8695 (N_8695,N_2154,N_4075);
and U8696 (N_8696,N_1049,N_436);
nor U8697 (N_8697,N_4606,N_1828);
or U8698 (N_8698,N_4945,N_1898);
or U8699 (N_8699,N_2415,N_290);
and U8700 (N_8700,N_1564,N_3931);
or U8701 (N_8701,N_3642,N_3301);
nand U8702 (N_8702,N_2702,N_780);
or U8703 (N_8703,N_2081,N_4194);
nand U8704 (N_8704,N_3006,N_2388);
or U8705 (N_8705,N_337,N_4246);
nor U8706 (N_8706,N_1016,N_699);
or U8707 (N_8707,N_3421,N_1774);
nor U8708 (N_8708,N_328,N_3892);
nor U8709 (N_8709,N_438,N_433);
nand U8710 (N_8710,N_3093,N_4533);
nor U8711 (N_8711,N_2520,N_884);
and U8712 (N_8712,N_3771,N_2589);
nand U8713 (N_8713,N_44,N_4919);
xor U8714 (N_8714,N_806,N_4420);
nand U8715 (N_8715,N_1895,N_2662);
nand U8716 (N_8716,N_2653,N_4909);
nor U8717 (N_8717,N_1799,N_3761);
nand U8718 (N_8718,N_804,N_437);
nand U8719 (N_8719,N_1536,N_4966);
and U8720 (N_8720,N_1461,N_3597);
nor U8721 (N_8721,N_823,N_2237);
and U8722 (N_8722,N_1648,N_2999);
and U8723 (N_8723,N_3556,N_1102);
nor U8724 (N_8724,N_3664,N_3222);
nand U8725 (N_8725,N_4944,N_2063);
or U8726 (N_8726,N_3881,N_4417);
or U8727 (N_8727,N_4018,N_3614);
and U8728 (N_8728,N_1198,N_2449);
nor U8729 (N_8729,N_2781,N_2254);
nand U8730 (N_8730,N_940,N_4201);
xnor U8731 (N_8731,N_2533,N_4375);
nor U8732 (N_8732,N_724,N_821);
or U8733 (N_8733,N_1983,N_439);
nor U8734 (N_8734,N_1745,N_2918);
nor U8735 (N_8735,N_1022,N_1396);
nor U8736 (N_8736,N_2084,N_3078);
nand U8737 (N_8737,N_2757,N_883);
xnor U8738 (N_8738,N_1300,N_1959);
and U8739 (N_8739,N_2176,N_3128);
and U8740 (N_8740,N_1533,N_2144);
or U8741 (N_8741,N_2516,N_91);
or U8742 (N_8742,N_4926,N_717);
and U8743 (N_8743,N_3885,N_3325);
or U8744 (N_8744,N_2004,N_1608);
and U8745 (N_8745,N_3408,N_1703);
nor U8746 (N_8746,N_1848,N_2498);
and U8747 (N_8747,N_2956,N_1093);
nand U8748 (N_8748,N_1148,N_2071);
or U8749 (N_8749,N_4173,N_128);
or U8750 (N_8750,N_2925,N_1423);
nand U8751 (N_8751,N_86,N_1281);
nor U8752 (N_8752,N_605,N_2309);
and U8753 (N_8753,N_8,N_1642);
or U8754 (N_8754,N_3246,N_1406);
and U8755 (N_8755,N_3173,N_741);
nand U8756 (N_8756,N_3080,N_3708);
or U8757 (N_8757,N_604,N_1416);
nor U8758 (N_8758,N_2752,N_461);
or U8759 (N_8759,N_3095,N_806);
nor U8760 (N_8760,N_422,N_1053);
nor U8761 (N_8761,N_1936,N_1);
or U8762 (N_8762,N_3778,N_4311);
nand U8763 (N_8763,N_1467,N_3947);
xnor U8764 (N_8764,N_2952,N_1114);
or U8765 (N_8765,N_1213,N_1627);
and U8766 (N_8766,N_3917,N_4335);
nand U8767 (N_8767,N_2886,N_4754);
nor U8768 (N_8768,N_1339,N_2330);
nor U8769 (N_8769,N_3444,N_654);
nand U8770 (N_8770,N_2201,N_3004);
nand U8771 (N_8771,N_2598,N_963);
or U8772 (N_8772,N_4548,N_473);
nor U8773 (N_8773,N_2189,N_1868);
and U8774 (N_8774,N_3076,N_4058);
and U8775 (N_8775,N_1681,N_2087);
nor U8776 (N_8776,N_2173,N_1327);
nand U8777 (N_8777,N_1755,N_4580);
nand U8778 (N_8778,N_1083,N_4404);
nor U8779 (N_8779,N_4050,N_1962);
nor U8780 (N_8780,N_1210,N_4095);
and U8781 (N_8781,N_2527,N_964);
or U8782 (N_8782,N_4938,N_2109);
nor U8783 (N_8783,N_3916,N_3425);
nor U8784 (N_8784,N_62,N_3688);
nand U8785 (N_8785,N_3366,N_2895);
xor U8786 (N_8786,N_4508,N_3273);
and U8787 (N_8787,N_3469,N_3053);
or U8788 (N_8788,N_4166,N_3372);
or U8789 (N_8789,N_4013,N_2191);
nor U8790 (N_8790,N_2940,N_2687);
and U8791 (N_8791,N_3349,N_3843);
nor U8792 (N_8792,N_2959,N_2736);
and U8793 (N_8793,N_2723,N_611);
and U8794 (N_8794,N_2473,N_3478);
nor U8795 (N_8795,N_2950,N_4592);
nand U8796 (N_8796,N_217,N_519);
nand U8797 (N_8797,N_2709,N_887);
or U8798 (N_8798,N_4756,N_3021);
or U8799 (N_8799,N_283,N_3032);
nor U8800 (N_8800,N_3875,N_3799);
and U8801 (N_8801,N_3758,N_4920);
and U8802 (N_8802,N_1128,N_3232);
or U8803 (N_8803,N_836,N_10);
or U8804 (N_8804,N_2306,N_1484);
and U8805 (N_8805,N_4993,N_1758);
nand U8806 (N_8806,N_4408,N_1408);
and U8807 (N_8807,N_3705,N_14);
nor U8808 (N_8808,N_2161,N_1736);
or U8809 (N_8809,N_3842,N_3087);
and U8810 (N_8810,N_1439,N_1870);
or U8811 (N_8811,N_4698,N_3705);
nor U8812 (N_8812,N_852,N_201);
and U8813 (N_8813,N_1633,N_2757);
nor U8814 (N_8814,N_3754,N_3522);
or U8815 (N_8815,N_2675,N_3119);
nor U8816 (N_8816,N_4026,N_4592);
and U8817 (N_8817,N_4274,N_108);
nand U8818 (N_8818,N_4385,N_4183);
nand U8819 (N_8819,N_1489,N_4977);
xor U8820 (N_8820,N_2202,N_2164);
or U8821 (N_8821,N_2558,N_719);
nor U8822 (N_8822,N_4492,N_2393);
nor U8823 (N_8823,N_991,N_118);
and U8824 (N_8824,N_60,N_4881);
and U8825 (N_8825,N_1861,N_2827);
and U8826 (N_8826,N_3293,N_4747);
and U8827 (N_8827,N_397,N_45);
or U8828 (N_8828,N_74,N_1032);
or U8829 (N_8829,N_1306,N_4219);
nand U8830 (N_8830,N_88,N_4940);
nor U8831 (N_8831,N_925,N_346);
nor U8832 (N_8832,N_108,N_2164);
and U8833 (N_8833,N_986,N_4470);
and U8834 (N_8834,N_2886,N_289);
nand U8835 (N_8835,N_1976,N_2825);
nor U8836 (N_8836,N_1024,N_4961);
or U8837 (N_8837,N_1942,N_3612);
nor U8838 (N_8838,N_3614,N_3447);
or U8839 (N_8839,N_482,N_2679);
or U8840 (N_8840,N_1586,N_1040);
or U8841 (N_8841,N_1560,N_1767);
nand U8842 (N_8842,N_2409,N_1722);
and U8843 (N_8843,N_1091,N_61);
and U8844 (N_8844,N_3217,N_2079);
nor U8845 (N_8845,N_3520,N_4999);
nand U8846 (N_8846,N_576,N_2638);
nand U8847 (N_8847,N_3400,N_1766);
or U8848 (N_8848,N_3633,N_3020);
nand U8849 (N_8849,N_2799,N_112);
and U8850 (N_8850,N_1395,N_4845);
nand U8851 (N_8851,N_328,N_4595);
nand U8852 (N_8852,N_4445,N_4547);
and U8853 (N_8853,N_2406,N_900);
and U8854 (N_8854,N_1818,N_614);
nor U8855 (N_8855,N_3811,N_3546);
and U8856 (N_8856,N_3711,N_967);
or U8857 (N_8857,N_3625,N_3796);
and U8858 (N_8858,N_2006,N_3001);
nor U8859 (N_8859,N_3753,N_1505);
and U8860 (N_8860,N_3861,N_501);
or U8861 (N_8861,N_3279,N_3110);
and U8862 (N_8862,N_2236,N_2462);
nand U8863 (N_8863,N_2116,N_1721);
or U8864 (N_8864,N_810,N_2852);
nand U8865 (N_8865,N_1322,N_726);
nor U8866 (N_8866,N_1916,N_3788);
nand U8867 (N_8867,N_2587,N_2077);
nor U8868 (N_8868,N_1872,N_1531);
and U8869 (N_8869,N_3797,N_4556);
or U8870 (N_8870,N_2751,N_3461);
nor U8871 (N_8871,N_4,N_3100);
nand U8872 (N_8872,N_2640,N_4726);
nor U8873 (N_8873,N_2977,N_741);
or U8874 (N_8874,N_1722,N_1101);
nor U8875 (N_8875,N_3511,N_428);
or U8876 (N_8876,N_2058,N_1006);
nor U8877 (N_8877,N_995,N_15);
nor U8878 (N_8878,N_3558,N_4279);
nor U8879 (N_8879,N_3472,N_1289);
or U8880 (N_8880,N_544,N_3274);
or U8881 (N_8881,N_470,N_10);
or U8882 (N_8882,N_4459,N_820);
or U8883 (N_8883,N_2649,N_672);
or U8884 (N_8884,N_1885,N_2611);
nand U8885 (N_8885,N_4700,N_3696);
nand U8886 (N_8886,N_601,N_4476);
and U8887 (N_8887,N_888,N_2029);
and U8888 (N_8888,N_1540,N_867);
nand U8889 (N_8889,N_343,N_2049);
nand U8890 (N_8890,N_454,N_4003);
nand U8891 (N_8891,N_3930,N_1774);
and U8892 (N_8892,N_4904,N_4342);
and U8893 (N_8893,N_4984,N_4693);
or U8894 (N_8894,N_557,N_2740);
nand U8895 (N_8895,N_2948,N_2706);
nor U8896 (N_8896,N_459,N_2692);
and U8897 (N_8897,N_3959,N_608);
nand U8898 (N_8898,N_2724,N_2677);
nor U8899 (N_8899,N_2737,N_19);
xor U8900 (N_8900,N_2042,N_3164);
nor U8901 (N_8901,N_4860,N_3385);
nand U8902 (N_8902,N_4243,N_1362);
nand U8903 (N_8903,N_2795,N_3178);
nand U8904 (N_8904,N_1002,N_4945);
xor U8905 (N_8905,N_2989,N_4465);
and U8906 (N_8906,N_2635,N_3237);
nand U8907 (N_8907,N_4111,N_2375);
nor U8908 (N_8908,N_1562,N_3991);
nand U8909 (N_8909,N_353,N_3456);
and U8910 (N_8910,N_643,N_828);
or U8911 (N_8911,N_4395,N_4195);
or U8912 (N_8912,N_442,N_1317);
nand U8913 (N_8913,N_2367,N_254);
xnor U8914 (N_8914,N_10,N_4355);
xor U8915 (N_8915,N_4968,N_2473);
nor U8916 (N_8916,N_1901,N_1554);
or U8917 (N_8917,N_351,N_1148);
or U8918 (N_8918,N_224,N_4701);
nand U8919 (N_8919,N_4591,N_2239);
and U8920 (N_8920,N_3933,N_3453);
and U8921 (N_8921,N_4717,N_117);
nor U8922 (N_8922,N_1858,N_2248);
nor U8923 (N_8923,N_545,N_1604);
or U8924 (N_8924,N_4915,N_4198);
nor U8925 (N_8925,N_2510,N_4961);
nand U8926 (N_8926,N_3632,N_4029);
nand U8927 (N_8927,N_2998,N_80);
or U8928 (N_8928,N_395,N_3741);
or U8929 (N_8929,N_4990,N_1836);
nand U8930 (N_8930,N_606,N_4773);
or U8931 (N_8931,N_1215,N_3782);
and U8932 (N_8932,N_1499,N_1048);
nor U8933 (N_8933,N_4178,N_3703);
nand U8934 (N_8934,N_788,N_1688);
and U8935 (N_8935,N_1970,N_3637);
nor U8936 (N_8936,N_571,N_4248);
or U8937 (N_8937,N_4853,N_4667);
or U8938 (N_8938,N_1162,N_4696);
nand U8939 (N_8939,N_4372,N_786);
nor U8940 (N_8940,N_4945,N_2778);
xnor U8941 (N_8941,N_1996,N_4622);
nand U8942 (N_8942,N_3536,N_3596);
xnor U8943 (N_8943,N_1465,N_3251);
nor U8944 (N_8944,N_314,N_4276);
nor U8945 (N_8945,N_3475,N_1103);
and U8946 (N_8946,N_1873,N_2006);
nor U8947 (N_8947,N_3385,N_2174);
nor U8948 (N_8948,N_1752,N_1253);
or U8949 (N_8949,N_3566,N_4533);
and U8950 (N_8950,N_4175,N_2472);
and U8951 (N_8951,N_1061,N_2260);
nand U8952 (N_8952,N_4396,N_2454);
nand U8953 (N_8953,N_2344,N_4105);
nand U8954 (N_8954,N_4923,N_2654);
nand U8955 (N_8955,N_4428,N_4880);
and U8956 (N_8956,N_2439,N_3907);
nand U8957 (N_8957,N_2594,N_867);
and U8958 (N_8958,N_2792,N_1096);
nand U8959 (N_8959,N_4965,N_3256);
xor U8960 (N_8960,N_772,N_1518);
nor U8961 (N_8961,N_746,N_350);
or U8962 (N_8962,N_2334,N_3084);
nor U8963 (N_8963,N_4495,N_4857);
nand U8964 (N_8964,N_4653,N_1189);
or U8965 (N_8965,N_2293,N_2787);
nor U8966 (N_8966,N_3950,N_808);
or U8967 (N_8967,N_4596,N_761);
or U8968 (N_8968,N_894,N_3663);
nand U8969 (N_8969,N_543,N_2244);
nor U8970 (N_8970,N_1947,N_1204);
nand U8971 (N_8971,N_3002,N_1113);
nor U8972 (N_8972,N_1465,N_805);
and U8973 (N_8973,N_421,N_4959);
or U8974 (N_8974,N_3674,N_3957);
nor U8975 (N_8975,N_4417,N_3138);
nor U8976 (N_8976,N_3568,N_3107);
nand U8977 (N_8977,N_4675,N_1580);
and U8978 (N_8978,N_1338,N_425);
or U8979 (N_8979,N_836,N_1490);
or U8980 (N_8980,N_3610,N_1866);
and U8981 (N_8981,N_412,N_4747);
and U8982 (N_8982,N_2855,N_3297);
or U8983 (N_8983,N_2371,N_3399);
or U8984 (N_8984,N_2245,N_749);
or U8985 (N_8985,N_2051,N_136);
or U8986 (N_8986,N_4739,N_3685);
and U8987 (N_8987,N_223,N_1826);
nor U8988 (N_8988,N_3293,N_4349);
nand U8989 (N_8989,N_3750,N_54);
or U8990 (N_8990,N_1442,N_3629);
nor U8991 (N_8991,N_32,N_3120);
and U8992 (N_8992,N_4414,N_529);
or U8993 (N_8993,N_4478,N_2547);
and U8994 (N_8994,N_4437,N_943);
or U8995 (N_8995,N_1364,N_2960);
or U8996 (N_8996,N_2665,N_703);
or U8997 (N_8997,N_4008,N_2344);
nand U8998 (N_8998,N_4183,N_3982);
nand U8999 (N_8999,N_3816,N_4953);
nor U9000 (N_9000,N_2597,N_2008);
nand U9001 (N_9001,N_2070,N_3195);
and U9002 (N_9002,N_4336,N_3066);
or U9003 (N_9003,N_306,N_1516);
and U9004 (N_9004,N_396,N_2763);
nor U9005 (N_9005,N_3183,N_992);
nor U9006 (N_9006,N_3330,N_3408);
or U9007 (N_9007,N_1788,N_4746);
nand U9008 (N_9008,N_1433,N_1537);
or U9009 (N_9009,N_430,N_4183);
nand U9010 (N_9010,N_6,N_4929);
xor U9011 (N_9011,N_4526,N_3728);
and U9012 (N_9012,N_2305,N_4591);
and U9013 (N_9013,N_4565,N_1082);
and U9014 (N_9014,N_3350,N_3309);
nand U9015 (N_9015,N_2925,N_2291);
or U9016 (N_9016,N_977,N_3522);
or U9017 (N_9017,N_3519,N_1360);
and U9018 (N_9018,N_2103,N_2591);
nand U9019 (N_9019,N_3659,N_2441);
and U9020 (N_9020,N_2369,N_1778);
nor U9021 (N_9021,N_1292,N_1488);
nand U9022 (N_9022,N_3197,N_2296);
or U9023 (N_9023,N_4999,N_951);
nand U9024 (N_9024,N_1034,N_3491);
and U9025 (N_9025,N_4322,N_3377);
nand U9026 (N_9026,N_4620,N_3547);
and U9027 (N_9027,N_153,N_4335);
nand U9028 (N_9028,N_3598,N_2543);
and U9029 (N_9029,N_668,N_2830);
or U9030 (N_9030,N_4588,N_3052);
nand U9031 (N_9031,N_2892,N_1152);
and U9032 (N_9032,N_850,N_523);
nand U9033 (N_9033,N_4708,N_2838);
or U9034 (N_9034,N_2580,N_2503);
or U9035 (N_9035,N_3507,N_3007);
nand U9036 (N_9036,N_4508,N_4852);
nor U9037 (N_9037,N_1337,N_2673);
nor U9038 (N_9038,N_1507,N_3922);
nor U9039 (N_9039,N_1961,N_1301);
nor U9040 (N_9040,N_3179,N_1523);
nor U9041 (N_9041,N_1277,N_637);
nand U9042 (N_9042,N_373,N_3360);
nor U9043 (N_9043,N_28,N_2115);
nand U9044 (N_9044,N_3227,N_4495);
nand U9045 (N_9045,N_2310,N_1729);
and U9046 (N_9046,N_2682,N_4777);
or U9047 (N_9047,N_1884,N_1442);
nand U9048 (N_9048,N_1388,N_955);
or U9049 (N_9049,N_3415,N_2846);
nor U9050 (N_9050,N_2384,N_2688);
nand U9051 (N_9051,N_2526,N_700);
and U9052 (N_9052,N_954,N_449);
nor U9053 (N_9053,N_1012,N_768);
nand U9054 (N_9054,N_1597,N_1912);
nor U9055 (N_9055,N_3809,N_45);
and U9056 (N_9056,N_1949,N_4158);
nand U9057 (N_9057,N_263,N_1893);
nand U9058 (N_9058,N_3770,N_3900);
nand U9059 (N_9059,N_1822,N_85);
or U9060 (N_9060,N_855,N_787);
nand U9061 (N_9061,N_4225,N_403);
or U9062 (N_9062,N_4757,N_3145);
and U9063 (N_9063,N_3397,N_1026);
nand U9064 (N_9064,N_4393,N_920);
and U9065 (N_9065,N_741,N_2660);
and U9066 (N_9066,N_4469,N_2172);
nor U9067 (N_9067,N_1237,N_635);
and U9068 (N_9068,N_3471,N_4528);
nor U9069 (N_9069,N_4614,N_3331);
nand U9070 (N_9070,N_55,N_16);
and U9071 (N_9071,N_572,N_1803);
and U9072 (N_9072,N_1619,N_2353);
and U9073 (N_9073,N_3423,N_1387);
nor U9074 (N_9074,N_943,N_1211);
or U9075 (N_9075,N_1388,N_4889);
nand U9076 (N_9076,N_374,N_2720);
or U9077 (N_9077,N_2705,N_4786);
and U9078 (N_9078,N_613,N_2525);
nand U9079 (N_9079,N_1993,N_835);
nand U9080 (N_9080,N_4001,N_2594);
nor U9081 (N_9081,N_2687,N_921);
nor U9082 (N_9082,N_15,N_579);
nand U9083 (N_9083,N_1179,N_3632);
or U9084 (N_9084,N_4067,N_699);
and U9085 (N_9085,N_2759,N_3498);
and U9086 (N_9086,N_3332,N_4750);
nand U9087 (N_9087,N_2126,N_4265);
and U9088 (N_9088,N_3249,N_2515);
nand U9089 (N_9089,N_98,N_3506);
nor U9090 (N_9090,N_2902,N_4582);
or U9091 (N_9091,N_72,N_4565);
nor U9092 (N_9092,N_3336,N_4623);
nor U9093 (N_9093,N_3345,N_1114);
and U9094 (N_9094,N_3968,N_1706);
or U9095 (N_9095,N_716,N_4952);
nor U9096 (N_9096,N_3503,N_4276);
or U9097 (N_9097,N_2046,N_4564);
and U9098 (N_9098,N_4055,N_173);
or U9099 (N_9099,N_4169,N_750);
and U9100 (N_9100,N_4781,N_3624);
nand U9101 (N_9101,N_1795,N_1930);
or U9102 (N_9102,N_136,N_3847);
nand U9103 (N_9103,N_3823,N_861);
nor U9104 (N_9104,N_2644,N_559);
nand U9105 (N_9105,N_341,N_3439);
or U9106 (N_9106,N_443,N_701);
and U9107 (N_9107,N_2750,N_2439);
and U9108 (N_9108,N_352,N_699);
nor U9109 (N_9109,N_4065,N_2690);
nor U9110 (N_9110,N_182,N_4184);
or U9111 (N_9111,N_476,N_2894);
nor U9112 (N_9112,N_2112,N_1239);
nor U9113 (N_9113,N_4425,N_2066);
or U9114 (N_9114,N_2480,N_4529);
and U9115 (N_9115,N_3727,N_3359);
nor U9116 (N_9116,N_2472,N_4172);
nor U9117 (N_9117,N_4858,N_165);
nor U9118 (N_9118,N_2245,N_4672);
xnor U9119 (N_9119,N_535,N_3370);
or U9120 (N_9120,N_1017,N_4744);
or U9121 (N_9121,N_1956,N_3751);
or U9122 (N_9122,N_1445,N_2796);
or U9123 (N_9123,N_2387,N_1614);
and U9124 (N_9124,N_4715,N_3241);
nand U9125 (N_9125,N_11,N_1125);
nand U9126 (N_9126,N_1431,N_3034);
or U9127 (N_9127,N_4660,N_2529);
nand U9128 (N_9128,N_2256,N_221);
nand U9129 (N_9129,N_1514,N_1586);
or U9130 (N_9130,N_4518,N_1863);
nand U9131 (N_9131,N_636,N_1405);
nand U9132 (N_9132,N_48,N_349);
nand U9133 (N_9133,N_97,N_3754);
or U9134 (N_9134,N_3956,N_2379);
and U9135 (N_9135,N_4729,N_1998);
nand U9136 (N_9136,N_3288,N_2406);
and U9137 (N_9137,N_3926,N_2973);
nor U9138 (N_9138,N_2151,N_3490);
nand U9139 (N_9139,N_1187,N_2310);
or U9140 (N_9140,N_2033,N_2255);
or U9141 (N_9141,N_2624,N_4579);
xnor U9142 (N_9142,N_4107,N_1784);
and U9143 (N_9143,N_3019,N_3041);
and U9144 (N_9144,N_871,N_3383);
nor U9145 (N_9145,N_1058,N_1456);
nand U9146 (N_9146,N_2545,N_2367);
nor U9147 (N_9147,N_146,N_3238);
nor U9148 (N_9148,N_2003,N_1746);
nor U9149 (N_9149,N_4243,N_3503);
and U9150 (N_9150,N_2448,N_3534);
and U9151 (N_9151,N_153,N_4980);
and U9152 (N_9152,N_1721,N_776);
or U9153 (N_9153,N_835,N_2368);
xnor U9154 (N_9154,N_4086,N_3740);
xnor U9155 (N_9155,N_1024,N_4053);
and U9156 (N_9156,N_4305,N_3352);
and U9157 (N_9157,N_971,N_1583);
nor U9158 (N_9158,N_3273,N_714);
nor U9159 (N_9159,N_2727,N_4864);
or U9160 (N_9160,N_1652,N_1472);
and U9161 (N_9161,N_3721,N_1615);
nand U9162 (N_9162,N_4759,N_3399);
nand U9163 (N_9163,N_3767,N_2722);
and U9164 (N_9164,N_2522,N_684);
nor U9165 (N_9165,N_3344,N_516);
and U9166 (N_9166,N_4303,N_2358);
and U9167 (N_9167,N_2069,N_1690);
or U9168 (N_9168,N_154,N_3365);
nor U9169 (N_9169,N_1354,N_3115);
xnor U9170 (N_9170,N_154,N_3726);
or U9171 (N_9171,N_273,N_1215);
nor U9172 (N_9172,N_3625,N_1125);
nand U9173 (N_9173,N_1209,N_4379);
or U9174 (N_9174,N_1049,N_1155);
or U9175 (N_9175,N_4438,N_1501);
nand U9176 (N_9176,N_1320,N_3157);
nand U9177 (N_9177,N_152,N_3155);
and U9178 (N_9178,N_546,N_4757);
nor U9179 (N_9179,N_3774,N_1824);
nand U9180 (N_9180,N_1520,N_527);
nand U9181 (N_9181,N_1259,N_2115);
and U9182 (N_9182,N_521,N_2295);
nor U9183 (N_9183,N_1671,N_608);
or U9184 (N_9184,N_4173,N_4886);
and U9185 (N_9185,N_4381,N_1802);
nor U9186 (N_9186,N_664,N_3968);
and U9187 (N_9187,N_4023,N_1404);
and U9188 (N_9188,N_434,N_459);
nand U9189 (N_9189,N_623,N_3846);
nand U9190 (N_9190,N_4528,N_1847);
nor U9191 (N_9191,N_80,N_171);
or U9192 (N_9192,N_1906,N_1810);
nand U9193 (N_9193,N_1611,N_1523);
nor U9194 (N_9194,N_4126,N_682);
and U9195 (N_9195,N_3020,N_3718);
and U9196 (N_9196,N_3690,N_1161);
and U9197 (N_9197,N_4479,N_3588);
nand U9198 (N_9198,N_4301,N_2029);
nand U9199 (N_9199,N_3288,N_605);
nor U9200 (N_9200,N_2486,N_4789);
nor U9201 (N_9201,N_4491,N_1466);
or U9202 (N_9202,N_4121,N_3324);
or U9203 (N_9203,N_4635,N_125);
nor U9204 (N_9204,N_2186,N_2406);
nand U9205 (N_9205,N_1333,N_1567);
nand U9206 (N_9206,N_974,N_4956);
nand U9207 (N_9207,N_3968,N_2608);
or U9208 (N_9208,N_3363,N_858);
nand U9209 (N_9209,N_3837,N_4569);
nand U9210 (N_9210,N_408,N_2011);
nor U9211 (N_9211,N_3402,N_2133);
or U9212 (N_9212,N_21,N_1941);
nand U9213 (N_9213,N_3371,N_1820);
nor U9214 (N_9214,N_4579,N_4247);
and U9215 (N_9215,N_2977,N_134);
nand U9216 (N_9216,N_4428,N_4918);
or U9217 (N_9217,N_2892,N_3211);
nor U9218 (N_9218,N_1803,N_978);
nor U9219 (N_9219,N_688,N_4624);
nor U9220 (N_9220,N_3250,N_3077);
nand U9221 (N_9221,N_1527,N_4580);
nand U9222 (N_9222,N_4504,N_2356);
and U9223 (N_9223,N_89,N_2406);
and U9224 (N_9224,N_1766,N_1459);
nand U9225 (N_9225,N_2737,N_4476);
nor U9226 (N_9226,N_3355,N_140);
or U9227 (N_9227,N_1385,N_4610);
and U9228 (N_9228,N_1410,N_3455);
xor U9229 (N_9229,N_3458,N_316);
or U9230 (N_9230,N_4363,N_3373);
or U9231 (N_9231,N_486,N_1152);
nor U9232 (N_9232,N_1838,N_208);
or U9233 (N_9233,N_559,N_14);
or U9234 (N_9234,N_679,N_1092);
nor U9235 (N_9235,N_166,N_2698);
nand U9236 (N_9236,N_4666,N_2985);
nand U9237 (N_9237,N_2902,N_3986);
or U9238 (N_9238,N_2961,N_1797);
or U9239 (N_9239,N_264,N_3928);
and U9240 (N_9240,N_1330,N_4401);
and U9241 (N_9241,N_4339,N_4952);
or U9242 (N_9242,N_3581,N_4240);
nor U9243 (N_9243,N_286,N_1575);
xor U9244 (N_9244,N_4220,N_2136);
or U9245 (N_9245,N_1875,N_4632);
xnor U9246 (N_9246,N_248,N_3821);
nor U9247 (N_9247,N_429,N_727);
or U9248 (N_9248,N_4644,N_4842);
nor U9249 (N_9249,N_3852,N_3822);
and U9250 (N_9250,N_3175,N_1273);
nor U9251 (N_9251,N_773,N_659);
or U9252 (N_9252,N_396,N_3540);
or U9253 (N_9253,N_1197,N_1905);
and U9254 (N_9254,N_2099,N_4665);
or U9255 (N_9255,N_3202,N_691);
nand U9256 (N_9256,N_1466,N_2053);
nand U9257 (N_9257,N_4634,N_1213);
and U9258 (N_9258,N_1335,N_2644);
and U9259 (N_9259,N_2329,N_4476);
and U9260 (N_9260,N_4392,N_3868);
and U9261 (N_9261,N_1290,N_1875);
nand U9262 (N_9262,N_3387,N_3255);
and U9263 (N_9263,N_2393,N_3675);
nand U9264 (N_9264,N_4790,N_711);
and U9265 (N_9265,N_342,N_4407);
and U9266 (N_9266,N_17,N_2519);
or U9267 (N_9267,N_2709,N_739);
and U9268 (N_9268,N_1111,N_2273);
nand U9269 (N_9269,N_1355,N_1072);
and U9270 (N_9270,N_2188,N_1082);
and U9271 (N_9271,N_1427,N_1102);
nand U9272 (N_9272,N_4358,N_3038);
or U9273 (N_9273,N_3020,N_224);
nor U9274 (N_9274,N_3320,N_4143);
nor U9275 (N_9275,N_739,N_3082);
nand U9276 (N_9276,N_267,N_707);
xor U9277 (N_9277,N_4103,N_3331);
or U9278 (N_9278,N_1691,N_604);
or U9279 (N_9279,N_2528,N_3608);
nor U9280 (N_9280,N_4705,N_846);
nor U9281 (N_9281,N_4850,N_60);
or U9282 (N_9282,N_4529,N_4843);
and U9283 (N_9283,N_3475,N_3462);
nor U9284 (N_9284,N_357,N_3571);
nand U9285 (N_9285,N_1171,N_1120);
or U9286 (N_9286,N_3254,N_3179);
nor U9287 (N_9287,N_4810,N_1599);
nand U9288 (N_9288,N_2269,N_1264);
nor U9289 (N_9289,N_1542,N_2909);
or U9290 (N_9290,N_2644,N_1472);
or U9291 (N_9291,N_4613,N_2556);
or U9292 (N_9292,N_60,N_4373);
xnor U9293 (N_9293,N_123,N_3429);
and U9294 (N_9294,N_1186,N_3996);
and U9295 (N_9295,N_489,N_4561);
nand U9296 (N_9296,N_1711,N_1732);
nor U9297 (N_9297,N_259,N_740);
nor U9298 (N_9298,N_3432,N_145);
xnor U9299 (N_9299,N_3705,N_4489);
nand U9300 (N_9300,N_2876,N_2854);
nand U9301 (N_9301,N_1554,N_2799);
or U9302 (N_9302,N_4418,N_3405);
nor U9303 (N_9303,N_508,N_3946);
or U9304 (N_9304,N_1614,N_3336);
and U9305 (N_9305,N_4553,N_1021);
nand U9306 (N_9306,N_250,N_4338);
nor U9307 (N_9307,N_3062,N_4095);
nand U9308 (N_9308,N_384,N_4536);
and U9309 (N_9309,N_4257,N_1887);
nand U9310 (N_9310,N_3862,N_4784);
and U9311 (N_9311,N_2202,N_3034);
or U9312 (N_9312,N_3138,N_2950);
nand U9313 (N_9313,N_2205,N_3770);
nor U9314 (N_9314,N_3842,N_675);
and U9315 (N_9315,N_1065,N_3932);
or U9316 (N_9316,N_119,N_3719);
nand U9317 (N_9317,N_1564,N_648);
nor U9318 (N_9318,N_3623,N_2823);
and U9319 (N_9319,N_2710,N_957);
nor U9320 (N_9320,N_2773,N_4130);
or U9321 (N_9321,N_4908,N_1220);
and U9322 (N_9322,N_751,N_3635);
and U9323 (N_9323,N_272,N_2284);
or U9324 (N_9324,N_2160,N_1450);
nor U9325 (N_9325,N_3195,N_834);
nor U9326 (N_9326,N_3900,N_2439);
nand U9327 (N_9327,N_2966,N_842);
nand U9328 (N_9328,N_513,N_4350);
nor U9329 (N_9329,N_4450,N_1647);
and U9330 (N_9330,N_1486,N_2634);
and U9331 (N_9331,N_24,N_4283);
or U9332 (N_9332,N_2025,N_2190);
nand U9333 (N_9333,N_2102,N_1423);
and U9334 (N_9334,N_4818,N_4086);
nor U9335 (N_9335,N_2934,N_3206);
or U9336 (N_9336,N_2307,N_2824);
nand U9337 (N_9337,N_4084,N_217);
nand U9338 (N_9338,N_1650,N_4853);
nor U9339 (N_9339,N_862,N_2538);
nor U9340 (N_9340,N_122,N_1480);
nor U9341 (N_9341,N_474,N_2284);
and U9342 (N_9342,N_714,N_970);
nor U9343 (N_9343,N_3982,N_112);
nor U9344 (N_9344,N_32,N_4598);
or U9345 (N_9345,N_2201,N_4947);
and U9346 (N_9346,N_4271,N_2449);
nor U9347 (N_9347,N_1538,N_950);
or U9348 (N_9348,N_670,N_4100);
and U9349 (N_9349,N_2587,N_4907);
or U9350 (N_9350,N_519,N_3978);
or U9351 (N_9351,N_1772,N_1280);
or U9352 (N_9352,N_3483,N_3639);
nor U9353 (N_9353,N_4359,N_3357);
nor U9354 (N_9354,N_662,N_2204);
and U9355 (N_9355,N_1728,N_1183);
nand U9356 (N_9356,N_1986,N_1260);
and U9357 (N_9357,N_4607,N_2773);
and U9358 (N_9358,N_3257,N_1780);
and U9359 (N_9359,N_2004,N_3765);
and U9360 (N_9360,N_2041,N_4563);
nor U9361 (N_9361,N_2885,N_1578);
nor U9362 (N_9362,N_4648,N_3698);
nand U9363 (N_9363,N_814,N_3218);
nor U9364 (N_9364,N_1981,N_713);
nor U9365 (N_9365,N_4166,N_4733);
or U9366 (N_9366,N_2292,N_2220);
nand U9367 (N_9367,N_2265,N_4430);
xnor U9368 (N_9368,N_1732,N_1516);
nor U9369 (N_9369,N_1472,N_1343);
or U9370 (N_9370,N_2590,N_2875);
nand U9371 (N_9371,N_2354,N_604);
or U9372 (N_9372,N_4398,N_796);
nor U9373 (N_9373,N_409,N_1662);
and U9374 (N_9374,N_2862,N_3135);
or U9375 (N_9375,N_3951,N_2689);
nor U9376 (N_9376,N_466,N_2342);
xor U9377 (N_9377,N_4084,N_751);
and U9378 (N_9378,N_3319,N_4503);
and U9379 (N_9379,N_1056,N_721);
and U9380 (N_9380,N_4770,N_3680);
nor U9381 (N_9381,N_3573,N_4142);
nand U9382 (N_9382,N_130,N_1951);
and U9383 (N_9383,N_2184,N_2849);
nor U9384 (N_9384,N_2144,N_1911);
or U9385 (N_9385,N_4786,N_3504);
or U9386 (N_9386,N_3062,N_631);
or U9387 (N_9387,N_1209,N_811);
nand U9388 (N_9388,N_3293,N_2065);
nor U9389 (N_9389,N_4334,N_4239);
or U9390 (N_9390,N_1775,N_4512);
nand U9391 (N_9391,N_4787,N_968);
or U9392 (N_9392,N_900,N_721);
or U9393 (N_9393,N_637,N_4717);
or U9394 (N_9394,N_2591,N_72);
nor U9395 (N_9395,N_140,N_2908);
nor U9396 (N_9396,N_1941,N_254);
or U9397 (N_9397,N_2831,N_3253);
nor U9398 (N_9398,N_4240,N_4352);
nand U9399 (N_9399,N_169,N_3340);
and U9400 (N_9400,N_3852,N_3752);
nand U9401 (N_9401,N_1140,N_4942);
and U9402 (N_9402,N_1552,N_292);
nand U9403 (N_9403,N_3453,N_212);
nor U9404 (N_9404,N_3320,N_2006);
and U9405 (N_9405,N_394,N_821);
or U9406 (N_9406,N_484,N_3741);
nand U9407 (N_9407,N_3709,N_1220);
and U9408 (N_9408,N_4638,N_491);
nand U9409 (N_9409,N_2849,N_913);
nand U9410 (N_9410,N_4914,N_3081);
and U9411 (N_9411,N_3181,N_2940);
nand U9412 (N_9412,N_483,N_2531);
or U9413 (N_9413,N_2731,N_2453);
or U9414 (N_9414,N_4841,N_2364);
nand U9415 (N_9415,N_3043,N_2553);
and U9416 (N_9416,N_4567,N_147);
and U9417 (N_9417,N_3045,N_1958);
nand U9418 (N_9418,N_1716,N_3943);
nor U9419 (N_9419,N_113,N_3123);
and U9420 (N_9420,N_2014,N_4474);
nor U9421 (N_9421,N_1525,N_234);
or U9422 (N_9422,N_800,N_480);
nor U9423 (N_9423,N_2539,N_2464);
and U9424 (N_9424,N_420,N_3628);
or U9425 (N_9425,N_3165,N_2050);
nor U9426 (N_9426,N_3,N_3382);
or U9427 (N_9427,N_2611,N_3882);
or U9428 (N_9428,N_4900,N_2850);
and U9429 (N_9429,N_733,N_4978);
nor U9430 (N_9430,N_1785,N_4384);
or U9431 (N_9431,N_1658,N_1771);
nand U9432 (N_9432,N_1555,N_4369);
nand U9433 (N_9433,N_408,N_1534);
nor U9434 (N_9434,N_2328,N_3747);
xor U9435 (N_9435,N_49,N_3705);
or U9436 (N_9436,N_1253,N_627);
or U9437 (N_9437,N_2345,N_1183);
nor U9438 (N_9438,N_4608,N_1449);
and U9439 (N_9439,N_1281,N_3314);
nand U9440 (N_9440,N_3758,N_4883);
nor U9441 (N_9441,N_1288,N_270);
nor U9442 (N_9442,N_2951,N_2470);
or U9443 (N_9443,N_4433,N_2989);
nand U9444 (N_9444,N_3225,N_4830);
and U9445 (N_9445,N_4391,N_155);
nand U9446 (N_9446,N_3729,N_4461);
nand U9447 (N_9447,N_1565,N_532);
nor U9448 (N_9448,N_2190,N_4411);
nand U9449 (N_9449,N_3121,N_2408);
nor U9450 (N_9450,N_2595,N_4654);
nand U9451 (N_9451,N_995,N_2728);
or U9452 (N_9452,N_514,N_1409);
nor U9453 (N_9453,N_277,N_4388);
or U9454 (N_9454,N_1341,N_321);
and U9455 (N_9455,N_3013,N_4851);
nor U9456 (N_9456,N_1408,N_1983);
nor U9457 (N_9457,N_3620,N_1570);
and U9458 (N_9458,N_1728,N_1217);
and U9459 (N_9459,N_3780,N_3288);
or U9460 (N_9460,N_2518,N_1731);
and U9461 (N_9461,N_2153,N_361);
or U9462 (N_9462,N_3266,N_4678);
and U9463 (N_9463,N_2901,N_3587);
and U9464 (N_9464,N_862,N_9);
and U9465 (N_9465,N_3529,N_2732);
nor U9466 (N_9466,N_554,N_2250);
or U9467 (N_9467,N_3199,N_3545);
and U9468 (N_9468,N_3186,N_3459);
nand U9469 (N_9469,N_3858,N_3750);
nand U9470 (N_9470,N_3724,N_2657);
or U9471 (N_9471,N_847,N_2212);
nand U9472 (N_9472,N_823,N_4513);
or U9473 (N_9473,N_4707,N_1890);
and U9474 (N_9474,N_3041,N_2560);
nand U9475 (N_9475,N_2229,N_3323);
and U9476 (N_9476,N_153,N_2420);
nor U9477 (N_9477,N_3880,N_2088);
and U9478 (N_9478,N_927,N_313);
or U9479 (N_9479,N_1916,N_4322);
or U9480 (N_9480,N_4911,N_503);
nand U9481 (N_9481,N_3076,N_76);
xnor U9482 (N_9482,N_2484,N_4643);
or U9483 (N_9483,N_3112,N_1053);
xor U9484 (N_9484,N_3993,N_251);
nand U9485 (N_9485,N_4450,N_1314);
or U9486 (N_9486,N_315,N_3285);
and U9487 (N_9487,N_1346,N_1320);
nand U9488 (N_9488,N_2790,N_869);
or U9489 (N_9489,N_2661,N_3103);
nor U9490 (N_9490,N_4680,N_1929);
nor U9491 (N_9491,N_3871,N_1460);
or U9492 (N_9492,N_4186,N_3394);
nand U9493 (N_9493,N_1399,N_4656);
and U9494 (N_9494,N_1565,N_1101);
or U9495 (N_9495,N_631,N_4136);
or U9496 (N_9496,N_2795,N_3248);
nor U9497 (N_9497,N_1968,N_4349);
xor U9498 (N_9498,N_2727,N_1512);
nor U9499 (N_9499,N_3592,N_1773);
or U9500 (N_9500,N_1241,N_2051);
nor U9501 (N_9501,N_2449,N_73);
nand U9502 (N_9502,N_80,N_2341);
or U9503 (N_9503,N_3039,N_2625);
or U9504 (N_9504,N_3584,N_2589);
nand U9505 (N_9505,N_1516,N_4999);
nand U9506 (N_9506,N_4657,N_4684);
and U9507 (N_9507,N_3258,N_331);
or U9508 (N_9508,N_162,N_4042);
and U9509 (N_9509,N_2080,N_2271);
nand U9510 (N_9510,N_403,N_3577);
nand U9511 (N_9511,N_1652,N_128);
xor U9512 (N_9512,N_4056,N_4941);
nor U9513 (N_9513,N_3245,N_537);
or U9514 (N_9514,N_1910,N_410);
nor U9515 (N_9515,N_1560,N_1848);
nor U9516 (N_9516,N_601,N_4153);
or U9517 (N_9517,N_290,N_4444);
and U9518 (N_9518,N_640,N_2695);
and U9519 (N_9519,N_935,N_439);
and U9520 (N_9520,N_1709,N_3590);
or U9521 (N_9521,N_4053,N_3085);
or U9522 (N_9522,N_2930,N_191);
nand U9523 (N_9523,N_4659,N_4222);
and U9524 (N_9524,N_1168,N_3098);
nor U9525 (N_9525,N_4182,N_4226);
or U9526 (N_9526,N_1449,N_3872);
nor U9527 (N_9527,N_1265,N_4669);
and U9528 (N_9528,N_3818,N_4222);
or U9529 (N_9529,N_3182,N_4897);
or U9530 (N_9530,N_1065,N_2789);
and U9531 (N_9531,N_150,N_2987);
nor U9532 (N_9532,N_1827,N_3999);
nor U9533 (N_9533,N_1398,N_1199);
nor U9534 (N_9534,N_3884,N_4987);
or U9535 (N_9535,N_134,N_2996);
nor U9536 (N_9536,N_3386,N_2820);
nand U9537 (N_9537,N_4199,N_3984);
and U9538 (N_9538,N_181,N_3432);
nand U9539 (N_9539,N_4498,N_681);
nand U9540 (N_9540,N_4810,N_4163);
nor U9541 (N_9541,N_235,N_3266);
or U9542 (N_9542,N_4758,N_1597);
nand U9543 (N_9543,N_2384,N_1813);
nor U9544 (N_9544,N_3566,N_4356);
nand U9545 (N_9545,N_2989,N_1181);
nor U9546 (N_9546,N_2766,N_4865);
or U9547 (N_9547,N_12,N_660);
and U9548 (N_9548,N_4610,N_1683);
and U9549 (N_9549,N_2341,N_1746);
or U9550 (N_9550,N_2585,N_800);
nand U9551 (N_9551,N_4000,N_3711);
or U9552 (N_9552,N_4351,N_1854);
and U9553 (N_9553,N_3796,N_137);
and U9554 (N_9554,N_1225,N_3047);
nor U9555 (N_9555,N_4550,N_3008);
or U9556 (N_9556,N_864,N_3568);
nand U9557 (N_9557,N_3451,N_924);
nor U9558 (N_9558,N_1369,N_2585);
or U9559 (N_9559,N_2064,N_3796);
or U9560 (N_9560,N_4814,N_2903);
nand U9561 (N_9561,N_1737,N_400);
nand U9562 (N_9562,N_1962,N_3625);
and U9563 (N_9563,N_2350,N_2812);
and U9564 (N_9564,N_2652,N_3942);
nor U9565 (N_9565,N_2565,N_4257);
nor U9566 (N_9566,N_1001,N_2965);
or U9567 (N_9567,N_1281,N_3997);
nand U9568 (N_9568,N_755,N_4611);
nand U9569 (N_9569,N_3523,N_480);
and U9570 (N_9570,N_1260,N_311);
nand U9571 (N_9571,N_3609,N_3119);
and U9572 (N_9572,N_2168,N_2915);
or U9573 (N_9573,N_376,N_446);
and U9574 (N_9574,N_2709,N_541);
and U9575 (N_9575,N_3580,N_3813);
or U9576 (N_9576,N_1178,N_2665);
and U9577 (N_9577,N_1004,N_1593);
nor U9578 (N_9578,N_953,N_3401);
and U9579 (N_9579,N_2266,N_2922);
xnor U9580 (N_9580,N_0,N_1959);
nor U9581 (N_9581,N_4319,N_91);
and U9582 (N_9582,N_644,N_54);
and U9583 (N_9583,N_3134,N_1615);
nand U9584 (N_9584,N_281,N_1473);
or U9585 (N_9585,N_740,N_158);
nand U9586 (N_9586,N_4376,N_2781);
nand U9587 (N_9587,N_3307,N_2224);
and U9588 (N_9588,N_3149,N_3528);
and U9589 (N_9589,N_3954,N_1716);
nand U9590 (N_9590,N_268,N_495);
and U9591 (N_9591,N_3302,N_1276);
and U9592 (N_9592,N_4506,N_4635);
nand U9593 (N_9593,N_759,N_4536);
and U9594 (N_9594,N_3530,N_2593);
and U9595 (N_9595,N_4488,N_107);
nor U9596 (N_9596,N_3407,N_1169);
nand U9597 (N_9597,N_2292,N_943);
nor U9598 (N_9598,N_1872,N_4761);
or U9599 (N_9599,N_1452,N_3217);
and U9600 (N_9600,N_1088,N_3642);
nor U9601 (N_9601,N_393,N_2233);
and U9602 (N_9602,N_2252,N_3908);
nor U9603 (N_9603,N_4534,N_3977);
xor U9604 (N_9604,N_2748,N_4135);
nand U9605 (N_9605,N_1985,N_3089);
and U9606 (N_9606,N_2752,N_4310);
or U9607 (N_9607,N_3206,N_605);
and U9608 (N_9608,N_2014,N_600);
and U9609 (N_9609,N_1736,N_4068);
and U9610 (N_9610,N_3822,N_4527);
nor U9611 (N_9611,N_3768,N_3409);
nand U9612 (N_9612,N_1306,N_2654);
or U9613 (N_9613,N_2441,N_328);
and U9614 (N_9614,N_3257,N_4125);
nand U9615 (N_9615,N_4085,N_893);
nand U9616 (N_9616,N_2336,N_2690);
or U9617 (N_9617,N_3679,N_4070);
nor U9618 (N_9618,N_4973,N_1678);
nor U9619 (N_9619,N_4686,N_1423);
nor U9620 (N_9620,N_2176,N_1794);
nand U9621 (N_9621,N_47,N_1369);
and U9622 (N_9622,N_1375,N_4030);
or U9623 (N_9623,N_3061,N_3389);
xnor U9624 (N_9624,N_4062,N_4615);
nand U9625 (N_9625,N_2065,N_244);
nand U9626 (N_9626,N_1895,N_1365);
and U9627 (N_9627,N_1578,N_719);
nor U9628 (N_9628,N_1327,N_1526);
and U9629 (N_9629,N_1833,N_4402);
or U9630 (N_9630,N_1335,N_3010);
and U9631 (N_9631,N_4851,N_1744);
and U9632 (N_9632,N_834,N_870);
or U9633 (N_9633,N_409,N_1099);
and U9634 (N_9634,N_3269,N_2700);
nand U9635 (N_9635,N_4767,N_4472);
nor U9636 (N_9636,N_1455,N_4464);
xor U9637 (N_9637,N_522,N_1353);
or U9638 (N_9638,N_2528,N_1107);
and U9639 (N_9639,N_246,N_777);
or U9640 (N_9640,N_3322,N_3483);
nand U9641 (N_9641,N_2209,N_1056);
nor U9642 (N_9642,N_428,N_2960);
and U9643 (N_9643,N_2774,N_491);
nor U9644 (N_9644,N_1969,N_4005);
nand U9645 (N_9645,N_3865,N_2758);
nor U9646 (N_9646,N_4157,N_3638);
nor U9647 (N_9647,N_4075,N_1489);
nand U9648 (N_9648,N_2937,N_782);
and U9649 (N_9649,N_2540,N_1587);
nand U9650 (N_9650,N_2089,N_3893);
and U9651 (N_9651,N_1906,N_4239);
and U9652 (N_9652,N_4055,N_65);
or U9653 (N_9653,N_2228,N_3020);
nand U9654 (N_9654,N_2989,N_3823);
nand U9655 (N_9655,N_4137,N_743);
and U9656 (N_9656,N_3398,N_765);
or U9657 (N_9657,N_1715,N_3524);
or U9658 (N_9658,N_2252,N_93);
and U9659 (N_9659,N_4954,N_3431);
or U9660 (N_9660,N_3464,N_1027);
and U9661 (N_9661,N_451,N_2904);
or U9662 (N_9662,N_2668,N_4807);
nor U9663 (N_9663,N_2984,N_404);
and U9664 (N_9664,N_2856,N_3070);
nand U9665 (N_9665,N_4466,N_2520);
nor U9666 (N_9666,N_1325,N_930);
nand U9667 (N_9667,N_3991,N_3595);
nor U9668 (N_9668,N_891,N_286);
or U9669 (N_9669,N_847,N_3676);
xnor U9670 (N_9670,N_4380,N_2142);
and U9671 (N_9671,N_2809,N_3691);
xnor U9672 (N_9672,N_797,N_2818);
or U9673 (N_9673,N_4318,N_4354);
nand U9674 (N_9674,N_2528,N_1236);
nand U9675 (N_9675,N_1195,N_3941);
and U9676 (N_9676,N_3052,N_1377);
and U9677 (N_9677,N_1469,N_4601);
and U9678 (N_9678,N_2309,N_3083);
or U9679 (N_9679,N_4112,N_2209);
or U9680 (N_9680,N_3836,N_2049);
or U9681 (N_9681,N_4014,N_3373);
and U9682 (N_9682,N_4915,N_1097);
nand U9683 (N_9683,N_1023,N_961);
or U9684 (N_9684,N_4662,N_1407);
or U9685 (N_9685,N_531,N_973);
nor U9686 (N_9686,N_3702,N_2861);
or U9687 (N_9687,N_4389,N_2295);
and U9688 (N_9688,N_2936,N_2625);
nor U9689 (N_9689,N_3570,N_4998);
nor U9690 (N_9690,N_1269,N_1026);
nor U9691 (N_9691,N_2386,N_1668);
nand U9692 (N_9692,N_4412,N_2055);
and U9693 (N_9693,N_2445,N_3303);
and U9694 (N_9694,N_1655,N_4914);
nor U9695 (N_9695,N_4971,N_1148);
nor U9696 (N_9696,N_276,N_1309);
and U9697 (N_9697,N_182,N_3667);
nand U9698 (N_9698,N_578,N_1992);
or U9699 (N_9699,N_1770,N_216);
nand U9700 (N_9700,N_3193,N_1178);
and U9701 (N_9701,N_3957,N_4674);
nor U9702 (N_9702,N_2719,N_2584);
and U9703 (N_9703,N_1644,N_2113);
and U9704 (N_9704,N_1419,N_370);
and U9705 (N_9705,N_186,N_3599);
or U9706 (N_9706,N_2588,N_1872);
or U9707 (N_9707,N_2789,N_2004);
or U9708 (N_9708,N_137,N_525);
xnor U9709 (N_9709,N_4440,N_2386);
xnor U9710 (N_9710,N_937,N_3129);
nand U9711 (N_9711,N_398,N_487);
or U9712 (N_9712,N_4166,N_3830);
nand U9713 (N_9713,N_4224,N_4449);
xor U9714 (N_9714,N_1571,N_4152);
xnor U9715 (N_9715,N_1196,N_4261);
nor U9716 (N_9716,N_3548,N_554);
and U9717 (N_9717,N_4638,N_287);
or U9718 (N_9718,N_3135,N_3685);
xnor U9719 (N_9719,N_3151,N_3191);
and U9720 (N_9720,N_2462,N_1997);
nor U9721 (N_9721,N_3365,N_2406);
or U9722 (N_9722,N_4190,N_19);
or U9723 (N_9723,N_2794,N_389);
nand U9724 (N_9724,N_3490,N_1098);
nor U9725 (N_9725,N_4854,N_2330);
or U9726 (N_9726,N_3404,N_1354);
nand U9727 (N_9727,N_2161,N_2671);
nand U9728 (N_9728,N_4878,N_4872);
and U9729 (N_9729,N_773,N_2246);
and U9730 (N_9730,N_310,N_4174);
nor U9731 (N_9731,N_1227,N_4339);
nand U9732 (N_9732,N_917,N_3427);
nand U9733 (N_9733,N_4441,N_4957);
or U9734 (N_9734,N_993,N_1648);
and U9735 (N_9735,N_166,N_1917);
or U9736 (N_9736,N_3766,N_4233);
xnor U9737 (N_9737,N_4972,N_1796);
nand U9738 (N_9738,N_4849,N_908);
nand U9739 (N_9739,N_661,N_1848);
and U9740 (N_9740,N_3181,N_762);
and U9741 (N_9741,N_2588,N_598);
and U9742 (N_9742,N_2677,N_4079);
nand U9743 (N_9743,N_4221,N_1520);
nor U9744 (N_9744,N_1130,N_2309);
and U9745 (N_9745,N_2961,N_4509);
nand U9746 (N_9746,N_4774,N_722);
or U9747 (N_9747,N_1459,N_1062);
or U9748 (N_9748,N_3759,N_2995);
nor U9749 (N_9749,N_938,N_3477);
nand U9750 (N_9750,N_1688,N_1226);
and U9751 (N_9751,N_3594,N_4380);
nand U9752 (N_9752,N_2969,N_3760);
or U9753 (N_9753,N_3279,N_3579);
or U9754 (N_9754,N_324,N_1725);
nor U9755 (N_9755,N_4726,N_1338);
nand U9756 (N_9756,N_45,N_4971);
nor U9757 (N_9757,N_1027,N_432);
nor U9758 (N_9758,N_4479,N_4269);
and U9759 (N_9759,N_12,N_3820);
nor U9760 (N_9760,N_2917,N_2728);
and U9761 (N_9761,N_3828,N_3417);
or U9762 (N_9762,N_2563,N_3993);
or U9763 (N_9763,N_2453,N_1214);
nor U9764 (N_9764,N_2865,N_3115);
nor U9765 (N_9765,N_1803,N_3800);
nor U9766 (N_9766,N_109,N_2868);
or U9767 (N_9767,N_4705,N_4031);
and U9768 (N_9768,N_4331,N_4264);
or U9769 (N_9769,N_2947,N_4273);
nor U9770 (N_9770,N_52,N_2591);
nand U9771 (N_9771,N_1854,N_2634);
or U9772 (N_9772,N_3314,N_3162);
nor U9773 (N_9773,N_2091,N_2253);
nand U9774 (N_9774,N_3945,N_789);
or U9775 (N_9775,N_3344,N_2371);
nor U9776 (N_9776,N_3339,N_1674);
xnor U9777 (N_9777,N_1930,N_2218);
nor U9778 (N_9778,N_1164,N_680);
nor U9779 (N_9779,N_4118,N_2210);
nor U9780 (N_9780,N_3161,N_4261);
nand U9781 (N_9781,N_74,N_1530);
and U9782 (N_9782,N_543,N_190);
or U9783 (N_9783,N_2306,N_295);
nand U9784 (N_9784,N_1657,N_4241);
nor U9785 (N_9785,N_13,N_4084);
or U9786 (N_9786,N_3445,N_4838);
nand U9787 (N_9787,N_4551,N_4297);
nand U9788 (N_9788,N_2952,N_3092);
and U9789 (N_9789,N_243,N_228);
nor U9790 (N_9790,N_1447,N_3211);
or U9791 (N_9791,N_197,N_2391);
or U9792 (N_9792,N_2000,N_4958);
and U9793 (N_9793,N_733,N_2167);
or U9794 (N_9794,N_265,N_4034);
and U9795 (N_9795,N_763,N_849);
and U9796 (N_9796,N_2609,N_2021);
nand U9797 (N_9797,N_913,N_2086);
nor U9798 (N_9798,N_3128,N_2944);
nand U9799 (N_9799,N_4939,N_1068);
nand U9800 (N_9800,N_3020,N_3116);
nor U9801 (N_9801,N_475,N_1390);
or U9802 (N_9802,N_690,N_3006);
nor U9803 (N_9803,N_62,N_566);
nand U9804 (N_9804,N_782,N_779);
nand U9805 (N_9805,N_1418,N_302);
nand U9806 (N_9806,N_446,N_921);
and U9807 (N_9807,N_965,N_2733);
or U9808 (N_9808,N_2631,N_2157);
nand U9809 (N_9809,N_2579,N_1865);
and U9810 (N_9810,N_3176,N_1051);
nor U9811 (N_9811,N_4641,N_1866);
and U9812 (N_9812,N_3080,N_3644);
or U9813 (N_9813,N_3617,N_297);
xor U9814 (N_9814,N_2582,N_1818);
or U9815 (N_9815,N_4449,N_3545);
or U9816 (N_9816,N_3699,N_3899);
nor U9817 (N_9817,N_703,N_2002);
nand U9818 (N_9818,N_2157,N_3567);
or U9819 (N_9819,N_3795,N_2684);
or U9820 (N_9820,N_4006,N_1033);
or U9821 (N_9821,N_304,N_811);
nor U9822 (N_9822,N_4741,N_1455);
and U9823 (N_9823,N_682,N_2906);
and U9824 (N_9824,N_800,N_971);
nand U9825 (N_9825,N_4263,N_3311);
or U9826 (N_9826,N_1711,N_325);
nand U9827 (N_9827,N_243,N_2034);
and U9828 (N_9828,N_43,N_2385);
nand U9829 (N_9829,N_849,N_972);
nor U9830 (N_9830,N_2023,N_3561);
nor U9831 (N_9831,N_1200,N_4771);
and U9832 (N_9832,N_2724,N_345);
nand U9833 (N_9833,N_4443,N_4913);
and U9834 (N_9834,N_1592,N_279);
and U9835 (N_9835,N_2746,N_1002);
and U9836 (N_9836,N_4433,N_1318);
or U9837 (N_9837,N_2521,N_1722);
nand U9838 (N_9838,N_2817,N_3712);
and U9839 (N_9839,N_255,N_2107);
nand U9840 (N_9840,N_588,N_1373);
nor U9841 (N_9841,N_1252,N_4549);
and U9842 (N_9842,N_3383,N_1533);
nor U9843 (N_9843,N_2271,N_4319);
nand U9844 (N_9844,N_2501,N_1029);
nor U9845 (N_9845,N_601,N_2672);
or U9846 (N_9846,N_2230,N_3741);
or U9847 (N_9847,N_1178,N_2900);
or U9848 (N_9848,N_2423,N_3541);
nand U9849 (N_9849,N_4322,N_3066);
nor U9850 (N_9850,N_1532,N_4651);
or U9851 (N_9851,N_1878,N_4088);
nor U9852 (N_9852,N_4198,N_2909);
nor U9853 (N_9853,N_4316,N_4932);
nand U9854 (N_9854,N_4182,N_2359);
and U9855 (N_9855,N_3379,N_4927);
nor U9856 (N_9856,N_3314,N_1019);
or U9857 (N_9857,N_1612,N_3480);
nor U9858 (N_9858,N_3100,N_4089);
nand U9859 (N_9859,N_992,N_3041);
or U9860 (N_9860,N_4314,N_326);
nor U9861 (N_9861,N_1982,N_3875);
nor U9862 (N_9862,N_1056,N_3237);
nand U9863 (N_9863,N_84,N_2611);
nand U9864 (N_9864,N_4161,N_2296);
and U9865 (N_9865,N_4099,N_691);
nand U9866 (N_9866,N_206,N_2000);
or U9867 (N_9867,N_4318,N_3591);
nand U9868 (N_9868,N_1140,N_1409);
nand U9869 (N_9869,N_2410,N_334);
and U9870 (N_9870,N_3456,N_3799);
and U9871 (N_9871,N_2292,N_4342);
and U9872 (N_9872,N_3610,N_270);
nand U9873 (N_9873,N_3319,N_4113);
and U9874 (N_9874,N_2364,N_3701);
and U9875 (N_9875,N_1900,N_3310);
or U9876 (N_9876,N_2181,N_4207);
nand U9877 (N_9877,N_3414,N_2952);
or U9878 (N_9878,N_1734,N_212);
and U9879 (N_9879,N_397,N_3319);
nor U9880 (N_9880,N_2970,N_1012);
and U9881 (N_9881,N_2206,N_2887);
and U9882 (N_9882,N_3267,N_3161);
nor U9883 (N_9883,N_1430,N_4570);
nor U9884 (N_9884,N_1606,N_4893);
nand U9885 (N_9885,N_4979,N_287);
nor U9886 (N_9886,N_4112,N_1504);
or U9887 (N_9887,N_2127,N_968);
or U9888 (N_9888,N_2676,N_4358);
and U9889 (N_9889,N_3977,N_361);
and U9890 (N_9890,N_2955,N_47);
nand U9891 (N_9891,N_1116,N_4968);
and U9892 (N_9892,N_2193,N_2681);
nor U9893 (N_9893,N_543,N_2093);
nand U9894 (N_9894,N_3345,N_4302);
and U9895 (N_9895,N_1138,N_3018);
nor U9896 (N_9896,N_3314,N_184);
nand U9897 (N_9897,N_3905,N_3104);
or U9898 (N_9898,N_478,N_4610);
or U9899 (N_9899,N_4975,N_1866);
nand U9900 (N_9900,N_3297,N_111);
nor U9901 (N_9901,N_1654,N_4522);
and U9902 (N_9902,N_4903,N_4292);
and U9903 (N_9903,N_3250,N_4343);
and U9904 (N_9904,N_1996,N_3788);
nand U9905 (N_9905,N_2754,N_1455);
nor U9906 (N_9906,N_1773,N_4181);
or U9907 (N_9907,N_3890,N_4486);
and U9908 (N_9908,N_3276,N_4032);
and U9909 (N_9909,N_133,N_3578);
nor U9910 (N_9910,N_3036,N_3707);
or U9911 (N_9911,N_4744,N_4932);
or U9912 (N_9912,N_692,N_1894);
or U9913 (N_9913,N_1756,N_1806);
and U9914 (N_9914,N_1463,N_129);
nor U9915 (N_9915,N_2000,N_2726);
and U9916 (N_9916,N_1321,N_2605);
or U9917 (N_9917,N_469,N_1727);
nor U9918 (N_9918,N_3976,N_4889);
and U9919 (N_9919,N_3350,N_1090);
or U9920 (N_9920,N_4580,N_1936);
nand U9921 (N_9921,N_3724,N_2971);
nand U9922 (N_9922,N_375,N_3714);
nor U9923 (N_9923,N_1471,N_324);
nand U9924 (N_9924,N_3635,N_4378);
or U9925 (N_9925,N_3770,N_3001);
xor U9926 (N_9926,N_3961,N_1246);
and U9927 (N_9927,N_4789,N_3947);
or U9928 (N_9928,N_342,N_4447);
xor U9929 (N_9929,N_1680,N_841);
nand U9930 (N_9930,N_278,N_3095);
nor U9931 (N_9931,N_2414,N_222);
xor U9932 (N_9932,N_2167,N_3837);
and U9933 (N_9933,N_1648,N_303);
nand U9934 (N_9934,N_2268,N_4027);
and U9935 (N_9935,N_2122,N_1533);
nand U9936 (N_9936,N_3410,N_1114);
nand U9937 (N_9937,N_686,N_2175);
nor U9938 (N_9938,N_1625,N_3107);
nand U9939 (N_9939,N_149,N_2853);
nand U9940 (N_9940,N_1941,N_1702);
or U9941 (N_9941,N_511,N_2095);
or U9942 (N_9942,N_3718,N_4335);
and U9943 (N_9943,N_3078,N_2489);
or U9944 (N_9944,N_1420,N_2137);
nor U9945 (N_9945,N_4954,N_2053);
or U9946 (N_9946,N_1288,N_1133);
nor U9947 (N_9947,N_1561,N_248);
nand U9948 (N_9948,N_4473,N_756);
nor U9949 (N_9949,N_4771,N_612);
or U9950 (N_9950,N_3439,N_1590);
or U9951 (N_9951,N_1973,N_793);
and U9952 (N_9952,N_3263,N_1598);
nand U9953 (N_9953,N_670,N_1678);
and U9954 (N_9954,N_4370,N_3909);
or U9955 (N_9955,N_139,N_2068);
nor U9956 (N_9956,N_414,N_3186);
and U9957 (N_9957,N_4799,N_2646);
nor U9958 (N_9958,N_4835,N_3040);
and U9959 (N_9959,N_3841,N_1263);
nand U9960 (N_9960,N_1831,N_4547);
nand U9961 (N_9961,N_2517,N_4564);
nand U9962 (N_9962,N_2683,N_2354);
nand U9963 (N_9963,N_2444,N_2677);
nor U9964 (N_9964,N_4073,N_3886);
nand U9965 (N_9965,N_3770,N_784);
xor U9966 (N_9966,N_1376,N_2939);
nor U9967 (N_9967,N_1532,N_3086);
xnor U9968 (N_9968,N_4216,N_1263);
or U9969 (N_9969,N_4214,N_2304);
and U9970 (N_9970,N_1902,N_2893);
and U9971 (N_9971,N_3322,N_3687);
nor U9972 (N_9972,N_3948,N_1152);
or U9973 (N_9973,N_1907,N_1942);
xnor U9974 (N_9974,N_2681,N_1849);
nand U9975 (N_9975,N_4698,N_3946);
or U9976 (N_9976,N_4857,N_1933);
nor U9977 (N_9977,N_3500,N_1123);
nand U9978 (N_9978,N_3152,N_1391);
nand U9979 (N_9979,N_3352,N_4885);
nand U9980 (N_9980,N_4207,N_1334);
nor U9981 (N_9981,N_4095,N_4383);
and U9982 (N_9982,N_3355,N_4893);
nand U9983 (N_9983,N_2500,N_4862);
and U9984 (N_9984,N_4729,N_1127);
nor U9985 (N_9985,N_2549,N_3429);
or U9986 (N_9986,N_2764,N_3626);
and U9987 (N_9987,N_1932,N_620);
and U9988 (N_9988,N_4024,N_3979);
nand U9989 (N_9989,N_597,N_1211);
or U9990 (N_9990,N_2574,N_3738);
or U9991 (N_9991,N_409,N_116);
nand U9992 (N_9992,N_3129,N_3109);
nand U9993 (N_9993,N_4838,N_717);
or U9994 (N_9994,N_2825,N_3056);
or U9995 (N_9995,N_4657,N_4588);
nor U9996 (N_9996,N_2296,N_2574);
nand U9997 (N_9997,N_972,N_2334);
and U9998 (N_9998,N_910,N_338);
nor U9999 (N_9999,N_3928,N_170);
or UO_0 (O_0,N_7479,N_5781);
nor UO_1 (O_1,N_5479,N_7718);
and UO_2 (O_2,N_5219,N_5466);
or UO_3 (O_3,N_9642,N_7351);
or UO_4 (O_4,N_6538,N_7085);
and UO_5 (O_5,N_6750,N_8441);
nor UO_6 (O_6,N_5365,N_6063);
nand UO_7 (O_7,N_6268,N_5569);
or UO_8 (O_8,N_9296,N_9837);
or UO_9 (O_9,N_5658,N_9881);
and UO_10 (O_10,N_8170,N_7816);
and UO_11 (O_11,N_7248,N_7174);
or UO_12 (O_12,N_6500,N_7165);
nand UO_13 (O_13,N_6235,N_9127);
nand UO_14 (O_14,N_8014,N_8943);
nand UO_15 (O_15,N_9740,N_5156);
and UO_16 (O_16,N_7742,N_9324);
or UO_17 (O_17,N_8904,N_8204);
or UO_18 (O_18,N_8201,N_9871);
nor UO_19 (O_19,N_8109,N_7975);
nor UO_20 (O_20,N_8474,N_6737);
nand UO_21 (O_21,N_9336,N_5670);
nor UO_22 (O_22,N_9057,N_9408);
nor UO_23 (O_23,N_5933,N_9147);
nand UO_24 (O_24,N_8467,N_7626);
nand UO_25 (O_25,N_7497,N_5847);
and UO_26 (O_26,N_7612,N_5359);
nand UO_27 (O_27,N_5362,N_5572);
nor UO_28 (O_28,N_7772,N_9510);
and UO_29 (O_29,N_5061,N_7394);
nor UO_30 (O_30,N_9527,N_9067);
or UO_31 (O_31,N_9678,N_7199);
or UO_32 (O_32,N_8333,N_8780);
or UO_33 (O_33,N_7989,N_9679);
nand UO_34 (O_34,N_7131,N_9716);
or UO_35 (O_35,N_8125,N_7910);
and UO_36 (O_36,N_7766,N_5643);
nor UO_37 (O_37,N_6592,N_9850);
nand UO_38 (O_38,N_8625,N_8387);
nand UO_39 (O_39,N_5964,N_7378);
and UO_40 (O_40,N_6212,N_6545);
nor UO_41 (O_41,N_5216,N_9557);
or UO_42 (O_42,N_7948,N_7689);
nor UO_43 (O_43,N_7927,N_8172);
and UO_44 (O_44,N_8838,N_7080);
nor UO_45 (O_45,N_9455,N_7643);
or UO_46 (O_46,N_9741,N_5307);
nand UO_47 (O_47,N_5026,N_6007);
nand UO_48 (O_48,N_8071,N_6362);
nand UO_49 (O_49,N_6757,N_5058);
nor UO_50 (O_50,N_5371,N_7933);
nor UO_51 (O_51,N_6780,N_7542);
nor UO_52 (O_52,N_5203,N_5095);
and UO_53 (O_53,N_8468,N_5722);
nand UO_54 (O_54,N_6800,N_7760);
and UO_55 (O_55,N_5090,N_6252);
nand UO_56 (O_56,N_5806,N_9235);
and UO_57 (O_57,N_9795,N_6760);
or UO_58 (O_58,N_6176,N_9236);
or UO_59 (O_59,N_8583,N_8935);
or UO_60 (O_60,N_8034,N_8844);
and UO_61 (O_61,N_5837,N_5169);
nor UO_62 (O_62,N_7840,N_6261);
nand UO_63 (O_63,N_5733,N_9356);
and UO_64 (O_64,N_8248,N_7860);
xnor UO_65 (O_65,N_6919,N_7453);
or UO_66 (O_66,N_9401,N_8191);
and UO_67 (O_67,N_8531,N_9903);
and UO_68 (O_68,N_6018,N_7337);
or UO_69 (O_69,N_5689,N_7220);
nand UO_70 (O_70,N_5303,N_8492);
nand UO_71 (O_71,N_6094,N_7460);
nor UO_72 (O_72,N_5653,N_6483);
nor UO_73 (O_73,N_7030,N_9593);
nand UO_74 (O_74,N_5690,N_8603);
and UO_75 (O_75,N_6150,N_9253);
nand UO_76 (O_76,N_8540,N_8792);
or UO_77 (O_77,N_6840,N_5279);
nor UO_78 (O_78,N_8427,N_7743);
nand UO_79 (O_79,N_6367,N_5502);
and UO_80 (O_80,N_9766,N_6103);
nand UO_81 (O_81,N_9524,N_6621);
nor UO_82 (O_82,N_8135,N_8178);
nand UO_83 (O_83,N_6651,N_8321);
nor UO_84 (O_84,N_9694,N_7599);
nand UO_85 (O_85,N_9874,N_9828);
nor UO_86 (O_86,N_5002,N_5474);
nand UO_87 (O_87,N_7804,N_6182);
nand UO_88 (O_88,N_7924,N_8083);
nor UO_89 (O_89,N_7365,N_8054);
nand UO_90 (O_90,N_7427,N_8395);
and UO_91 (O_91,N_9586,N_8657);
nand UO_92 (O_92,N_8070,N_9106);
and UO_93 (O_93,N_7702,N_5958);
nor UO_94 (O_94,N_7719,N_8401);
and UO_95 (O_95,N_8377,N_6655);
nand UO_96 (O_96,N_5411,N_8850);
and UO_97 (O_97,N_9998,N_5185);
and UO_98 (O_98,N_8629,N_6769);
and UO_99 (O_99,N_8475,N_7455);
nor UO_100 (O_100,N_6186,N_7155);
nor UO_101 (O_101,N_6220,N_6251);
nor UO_102 (O_102,N_8899,N_8330);
or UO_103 (O_103,N_5776,N_8458);
nand UO_104 (O_104,N_5092,N_7143);
nor UO_105 (O_105,N_7906,N_5327);
nand UO_106 (O_106,N_6696,N_6831);
or UO_107 (O_107,N_6819,N_5969);
nor UO_108 (O_108,N_8013,N_6353);
nor UO_109 (O_109,N_9706,N_5387);
and UO_110 (O_110,N_5779,N_6626);
and UO_111 (O_111,N_7069,N_7728);
nor UO_112 (O_112,N_8922,N_8591);
nor UO_113 (O_113,N_9447,N_7587);
nor UO_114 (O_114,N_5119,N_6173);
nand UO_115 (O_115,N_9051,N_9457);
or UO_116 (O_116,N_8337,N_5178);
nor UO_117 (O_117,N_6991,N_8880);
nor UO_118 (O_118,N_8534,N_9569);
nor UO_119 (O_119,N_5443,N_7466);
nor UO_120 (O_120,N_6127,N_7622);
and UO_121 (O_121,N_5903,N_8686);
nand UO_122 (O_122,N_9878,N_5591);
nand UO_123 (O_123,N_5366,N_9392);
and UO_124 (O_124,N_5065,N_7683);
or UO_125 (O_125,N_7234,N_7524);
nand UO_126 (O_126,N_6658,N_8350);
nand UO_127 (O_127,N_7281,N_9574);
and UO_128 (O_128,N_8815,N_5114);
nand UO_129 (O_129,N_5323,N_5580);
nor UO_130 (O_130,N_9971,N_6882);
nor UO_131 (O_131,N_7959,N_5107);
and UO_132 (O_132,N_7389,N_7151);
nor UO_133 (O_133,N_8845,N_6188);
nor UO_134 (O_134,N_9717,N_5336);
xor UO_135 (O_135,N_9161,N_5313);
or UO_136 (O_136,N_6908,N_9768);
xnor UO_137 (O_137,N_9399,N_8003);
nor UO_138 (O_138,N_6472,N_5745);
nor UO_139 (O_139,N_6590,N_9108);
nor UO_140 (O_140,N_7516,N_6948);
nor UO_141 (O_141,N_7409,N_5145);
and UO_142 (O_142,N_8498,N_9341);
xor UO_143 (O_143,N_7846,N_8897);
and UO_144 (O_144,N_9544,N_5438);
nor UO_145 (O_145,N_6710,N_8763);
or UO_146 (O_146,N_5924,N_7486);
nor UO_147 (O_147,N_9503,N_8554);
xnor UO_148 (O_148,N_8536,N_5310);
or UO_149 (O_149,N_6872,N_9267);
nor UO_150 (O_150,N_9536,N_7392);
nand UO_151 (O_151,N_6042,N_8995);
xor UO_152 (O_152,N_9489,N_7700);
nor UO_153 (O_153,N_9529,N_9495);
and UO_154 (O_154,N_7709,N_5423);
nand UO_155 (O_155,N_5814,N_6891);
nor UO_156 (O_156,N_8101,N_6324);
and UO_157 (O_157,N_9224,N_8920);
or UO_158 (O_158,N_6321,N_8903);
and UO_159 (O_159,N_7041,N_6735);
nor UO_160 (O_160,N_6053,N_6951);
or UO_161 (O_161,N_5351,N_5442);
nand UO_162 (O_162,N_9686,N_6743);
and UO_163 (O_163,N_6070,N_6000);
nor UO_164 (O_164,N_9938,N_7917);
and UO_165 (O_165,N_7915,N_5631);
nand UO_166 (O_166,N_5281,N_8209);
and UO_167 (O_167,N_9985,N_9330);
nand UO_168 (O_168,N_7062,N_8579);
and UO_169 (O_169,N_8038,N_5570);
nand UO_170 (O_170,N_7211,N_8478);
nand UO_171 (O_171,N_7834,N_8386);
and UO_172 (O_172,N_7032,N_7480);
or UO_173 (O_173,N_8994,N_5153);
nand UO_174 (O_174,N_5714,N_6405);
nor UO_175 (O_175,N_5273,N_9266);
nor UO_176 (O_176,N_8491,N_5163);
and UO_177 (O_177,N_5356,N_5805);
nor UO_178 (O_178,N_9910,N_7271);
or UO_179 (O_179,N_9928,N_7302);
nand UO_180 (O_180,N_6269,N_7472);
and UO_181 (O_181,N_8449,N_8433);
nand UO_182 (O_182,N_8050,N_7641);
nand UO_183 (O_183,N_8108,N_5031);
nor UO_184 (O_184,N_7146,N_6529);
and UO_185 (O_185,N_5704,N_8339);
or UO_186 (O_186,N_9261,N_7735);
or UO_187 (O_187,N_5605,N_6947);
nor UO_188 (O_188,N_9037,N_6377);
nor UO_189 (O_189,N_5982,N_9228);
or UO_190 (O_190,N_5735,N_6154);
nor UO_191 (O_191,N_5651,N_9939);
xnor UO_192 (O_192,N_5575,N_9595);
or UO_193 (O_193,N_7417,N_5025);
or UO_194 (O_194,N_9786,N_6921);
nand UO_195 (O_195,N_8161,N_8102);
nand UO_196 (O_196,N_9525,N_8722);
nand UO_197 (O_197,N_8821,N_9827);
and UO_198 (O_198,N_7613,N_5050);
and UO_199 (O_199,N_7078,N_8368);
and UO_200 (O_200,N_7693,N_5046);
nand UO_201 (O_201,N_9386,N_7525);
nand UO_202 (O_202,N_7185,N_7849);
or UO_203 (O_203,N_9930,N_7190);
or UO_204 (O_204,N_5737,N_7968);
or UO_205 (O_205,N_7096,N_8932);
nor UO_206 (O_206,N_9745,N_7025);
nor UO_207 (O_207,N_7859,N_5463);
nand UO_208 (O_208,N_9916,N_9785);
nor UO_209 (O_209,N_9986,N_6850);
xnor UO_210 (O_210,N_7082,N_9722);
nor UO_211 (O_211,N_6732,N_8493);
nand UO_212 (O_212,N_6709,N_8879);
nor UO_213 (O_213,N_9240,N_7355);
and UO_214 (O_214,N_6668,N_9777);
nor UO_215 (O_215,N_9379,N_7379);
and UO_216 (O_216,N_5942,N_8504);
xnor UO_217 (O_217,N_7255,N_7822);
nor UO_218 (O_218,N_5346,N_8187);
and UO_219 (O_219,N_6312,N_5673);
or UO_220 (O_220,N_8304,N_5703);
nor UO_221 (O_221,N_9382,N_7784);
or UO_222 (O_222,N_9007,N_6841);
and UO_223 (O_223,N_6851,N_5786);
or UO_224 (O_224,N_6184,N_7420);
or UO_225 (O_225,N_6790,N_7873);
nand UO_226 (O_226,N_6979,N_9921);
nand UO_227 (O_227,N_8749,N_6010);
or UO_228 (O_228,N_5915,N_9223);
nand UO_229 (O_229,N_9444,N_6749);
nand UO_230 (O_230,N_9549,N_5309);
and UO_231 (O_231,N_5836,N_7692);
nor UO_232 (O_232,N_5455,N_8481);
nor UO_233 (O_233,N_5268,N_6469);
nand UO_234 (O_234,N_5447,N_7419);
nor UO_235 (O_235,N_5376,N_8026);
nor UO_236 (O_236,N_7803,N_8760);
and UO_237 (O_237,N_7006,N_8260);
or UO_238 (O_238,N_6953,N_5978);
or UO_239 (O_239,N_5030,N_9798);
and UO_240 (O_240,N_7909,N_6443);
and UO_241 (O_241,N_8887,N_7869);
and UO_242 (O_242,N_9825,N_8335);
nor UO_243 (O_243,N_7245,N_6016);
or UO_244 (O_244,N_8354,N_8244);
nor UO_245 (O_245,N_6835,N_6166);
nor UO_246 (O_246,N_6167,N_7888);
nand UO_247 (O_247,N_6195,N_8099);
nand UO_248 (O_248,N_7157,N_6807);
nand UO_249 (O_249,N_8403,N_5707);
and UO_250 (O_250,N_7598,N_7176);
and UO_251 (O_251,N_6153,N_7246);
and UO_252 (O_252,N_7467,N_7218);
nand UO_253 (O_253,N_5028,N_8207);
nor UO_254 (O_254,N_8518,N_5062);
nor UO_255 (O_255,N_7299,N_8343);
nor UO_256 (O_256,N_8596,N_9990);
or UO_257 (O_257,N_6510,N_9947);
nor UO_258 (O_258,N_9661,N_9538);
and UO_259 (O_259,N_9935,N_6243);
nor UO_260 (O_260,N_6684,N_8284);
and UO_261 (O_261,N_5968,N_8598);
or UO_262 (O_262,N_7729,N_9258);
nand UO_263 (O_263,N_6532,N_5518);
nor UO_264 (O_264,N_8707,N_8486);
and UO_265 (O_265,N_5330,N_6722);
nor UO_266 (O_266,N_7748,N_5769);
xnor UO_267 (O_267,N_5419,N_5235);
nor UO_268 (O_268,N_6899,N_7962);
and UO_269 (O_269,N_9855,N_5338);
or UO_270 (O_270,N_6145,N_5688);
and UO_271 (O_271,N_9961,N_5602);
nor UO_272 (O_272,N_9136,N_6878);
nor UO_273 (O_273,N_9133,N_7077);
and UO_274 (O_274,N_6803,N_8262);
and UO_275 (O_275,N_8764,N_9426);
and UO_276 (O_276,N_6904,N_9934);
or UO_277 (O_277,N_8348,N_9188);
or UO_278 (O_278,N_7847,N_8236);
and UO_279 (O_279,N_7903,N_8927);
and UO_280 (O_280,N_6004,N_9863);
or UO_281 (O_281,N_6326,N_6620);
and UO_282 (O_282,N_8575,N_8770);
and UO_283 (O_283,N_5041,N_9395);
or UO_284 (O_284,N_9388,N_8389);
nor UO_285 (O_285,N_5223,N_6833);
and UO_286 (O_286,N_9018,N_6060);
or UO_287 (O_287,N_6989,N_7415);
nand UO_288 (O_288,N_9323,N_8325);
and UO_289 (O_289,N_6230,N_7960);
and UO_290 (O_290,N_5398,N_9482);
and UO_291 (O_291,N_8664,N_5908);
and UO_292 (O_292,N_7684,N_9911);
nand UO_293 (O_293,N_9400,N_7442);
nor UO_294 (O_294,N_7835,N_8599);
nor UO_295 (O_295,N_9300,N_6172);
nand UO_296 (O_296,N_9669,N_5794);
xnor UO_297 (O_297,N_9187,N_9234);
or UO_298 (O_298,N_6128,N_5173);
or UO_299 (O_299,N_9427,N_6298);
nor UO_300 (O_300,N_8173,N_5788);
nand UO_301 (O_301,N_6075,N_8302);
and UO_302 (O_302,N_5824,N_6662);
nand UO_303 (O_303,N_6605,N_7276);
or UO_304 (O_304,N_9282,N_8222);
nor UO_305 (O_305,N_9782,N_8517);
nor UO_306 (O_306,N_7652,N_6864);
nand UO_307 (O_307,N_6748,N_7750);
nand UO_308 (O_308,N_9492,N_7054);
nor UO_309 (O_309,N_5742,N_6496);
nor UO_310 (O_310,N_7004,N_7123);
nor UO_311 (O_311,N_7076,N_8698);
nor UO_312 (O_312,N_7242,N_8681);
and UO_313 (O_313,N_6858,N_6234);
or UO_314 (O_314,N_9584,N_6700);
and UO_315 (O_315,N_7349,N_5057);
and UO_316 (O_316,N_8048,N_7861);
nand UO_317 (O_317,N_7899,N_7391);
or UO_318 (O_318,N_7940,N_9734);
and UO_319 (O_319,N_9963,N_6633);
or UO_320 (O_320,N_8081,N_6586);
or UO_321 (O_321,N_8870,N_7440);
nor UO_322 (O_322,N_7883,N_6600);
nand UO_323 (O_323,N_5654,N_6178);
nand UO_324 (O_324,N_5304,N_5981);
or UO_325 (O_325,N_6236,N_7459);
nand UO_326 (O_326,N_5453,N_6536);
or UO_327 (O_327,N_6995,N_6565);
or UO_328 (O_328,N_6986,N_7588);
nor UO_329 (O_329,N_5427,N_6521);
nand UO_330 (O_330,N_6577,N_6418);
or UO_331 (O_331,N_6376,N_6849);
nand UO_332 (O_332,N_5679,N_8211);
nor UO_333 (O_333,N_7843,N_5392);
nand UO_334 (O_334,N_9824,N_9648);
and UO_335 (O_335,N_6993,N_6466);
and UO_336 (O_336,N_5881,N_9045);
nand UO_337 (O_337,N_9391,N_8342);
or UO_338 (O_338,N_5731,N_6115);
nor UO_339 (O_339,N_9890,N_7550);
nand UO_340 (O_340,N_9080,N_7801);
xnor UO_341 (O_341,N_9124,N_9338);
xor UO_342 (O_342,N_9583,N_6135);
or UO_343 (O_343,N_6387,N_8736);
and UO_344 (O_344,N_6058,N_6628);
nor UO_345 (O_345,N_6718,N_5947);
and UO_346 (O_346,N_7753,N_5233);
nand UO_347 (O_347,N_5245,N_6008);
nand UO_348 (O_348,N_5839,N_7039);
nor UO_349 (O_349,N_6960,N_7485);
and UO_350 (O_350,N_5301,N_9636);
nor UO_351 (O_351,N_8516,N_6049);
nor UO_352 (O_352,N_6752,N_7519);
nor UO_353 (O_353,N_9672,N_7708);
nor UO_354 (O_354,N_7536,N_6451);
or UO_355 (O_355,N_8167,N_5540);
nand UO_356 (O_356,N_6400,N_8501);
nor UO_357 (O_357,N_7053,N_8298);
and UO_358 (O_358,N_7400,N_9475);
nand UO_359 (O_359,N_8131,N_8238);
or UO_360 (O_360,N_7582,N_7602);
and UO_361 (O_361,N_5483,N_9857);
nor UO_362 (O_362,N_8232,N_9275);
nor UO_363 (O_363,N_5094,N_9005);
nand UO_364 (O_364,N_6608,N_8273);
nor UO_365 (O_365,N_7217,N_7705);
and UO_366 (O_366,N_6231,N_5285);
or UO_367 (O_367,N_9281,N_9621);
or UO_368 (O_368,N_8500,N_8265);
nand UO_369 (O_369,N_9831,N_5949);
and UO_370 (O_370,N_5300,N_8926);
and UO_371 (O_371,N_8743,N_8062);
nor UO_372 (O_372,N_7528,N_7716);
or UO_373 (O_373,N_5812,N_7955);
nand UO_374 (O_374,N_7125,N_8307);
or UO_375 (O_375,N_9152,N_9171);
nor UO_376 (O_376,N_5260,N_9058);
nand UO_377 (O_377,N_7347,N_9695);
nand UO_378 (O_378,N_7396,N_9848);
and UO_379 (O_379,N_6978,N_9762);
or UO_380 (O_380,N_8233,N_6740);
and UO_381 (O_381,N_5807,N_8606);
xnor UO_382 (O_382,N_9978,N_7807);
nor UO_383 (O_383,N_9480,N_9950);
nor UO_384 (O_384,N_8317,N_8004);
and UO_385 (O_385,N_8503,N_8957);
or UO_386 (O_386,N_9897,N_5750);
and UO_387 (O_387,N_5516,N_6778);
nand UO_388 (O_388,N_8509,N_9446);
or UO_389 (O_389,N_9919,N_8221);
and UO_390 (O_390,N_8185,N_9571);
nor UO_391 (O_391,N_9436,N_6028);
nor UO_392 (O_392,N_5087,N_5638);
nand UO_393 (O_393,N_6366,N_9693);
nand UO_394 (O_394,N_9699,N_7159);
and UO_395 (O_395,N_6068,N_6892);
nor UO_396 (O_396,N_6552,N_5868);
nand UO_397 (O_397,N_8746,N_7904);
nor UO_398 (O_398,N_5842,N_5409);
and UO_399 (O_399,N_8414,N_9579);
or UO_400 (O_400,N_5914,N_5866);
and UO_401 (O_401,N_9092,N_9239);
and UO_402 (O_402,N_5543,N_5925);
nand UO_403 (O_403,N_8608,N_9748);
or UO_404 (O_404,N_6436,N_8645);
nand UO_405 (O_405,N_5258,N_6909);
and UO_406 (O_406,N_5831,N_6467);
nor UO_407 (O_407,N_5636,N_5149);
nand UO_408 (O_408,N_9882,N_6185);
and UO_409 (O_409,N_8460,N_8600);
or UO_410 (O_410,N_5402,N_5410);
or UO_411 (O_411,N_8507,N_7788);
nor UO_412 (O_412,N_9737,N_8544);
nand UO_413 (O_413,N_8067,N_8510);
or UO_414 (O_414,N_6885,N_9488);
and UO_415 (O_415,N_6123,N_9813);
xnor UO_416 (O_416,N_8824,N_5302);
or UO_417 (O_417,N_6373,N_9011);
and UO_418 (O_418,N_7926,N_8437);
nand UO_419 (O_419,N_9074,N_8465);
nor UO_420 (O_420,N_9359,N_7776);
nor UO_421 (O_421,N_5103,N_5311);
nor UO_422 (O_422,N_9575,N_7891);
nor UO_423 (O_423,N_8662,N_8020);
and UO_424 (O_424,N_7227,N_9470);
or UO_425 (O_425,N_7414,N_6265);
nand UO_426 (O_426,N_5197,N_9808);
nor UO_427 (O_427,N_8093,N_8310);
or UO_428 (O_428,N_5488,N_9906);
or UO_429 (O_429,N_8963,N_6980);
and UO_430 (O_430,N_7979,N_8812);
nor UO_431 (O_431,N_7061,N_5512);
nand UO_432 (O_432,N_9702,N_6002);
nand UO_433 (O_433,N_5927,N_7311);
nor UO_434 (O_434,N_8079,N_6071);
or UO_435 (O_435,N_8594,N_9806);
or UO_436 (O_436,N_9344,N_6283);
nand UO_437 (O_437,N_5193,N_8773);
and UO_438 (O_438,N_6598,N_6407);
nor UO_439 (O_439,N_5497,N_5622);
xor UO_440 (O_440,N_6571,N_8419);
or UO_441 (O_441,N_9019,N_8968);
and UO_442 (O_442,N_6964,N_7896);
nor UO_443 (O_443,N_8382,N_7639);
nand UO_444 (O_444,N_5860,N_9351);
nor UO_445 (O_445,N_8863,N_7688);
nor UO_446 (O_446,N_6097,N_5125);
and UO_447 (O_447,N_7818,N_8529);
nand UO_448 (O_448,N_6119,N_5270);
and UO_449 (O_449,N_6755,N_5291);
and UO_450 (O_450,N_7008,N_5343);
xor UO_451 (O_451,N_7059,N_6320);
or UO_452 (O_452,N_7865,N_6292);
nand UO_453 (O_453,N_9826,N_6454);
or UO_454 (O_454,N_8858,N_5504);
nand UO_455 (O_455,N_7286,N_7385);
nor UO_456 (O_456,N_5526,N_9499);
or UO_457 (O_457,N_7775,N_6660);
or UO_458 (O_458,N_8356,N_6022);
or UO_459 (O_459,N_9555,N_7471);
nor UO_460 (O_460,N_7318,N_9190);
nand UO_461 (O_461,N_8946,N_6224);
nand UO_462 (O_462,N_6828,N_9464);
and UO_463 (O_463,N_8929,N_7722);
and UO_464 (O_464,N_8000,N_6138);
nand UO_465 (O_465,N_8789,N_8388);
nand UO_466 (O_466,N_7504,N_7293);
or UO_467 (O_467,N_7274,N_8230);
nand UO_468 (O_468,N_8872,N_6168);
nand UO_469 (O_469,N_6524,N_7045);
and UO_470 (O_470,N_5054,N_7509);
nand UO_471 (O_471,N_8533,N_7540);
or UO_472 (O_472,N_6548,N_7239);
nand UO_473 (O_473,N_9794,N_6064);
nor UO_474 (O_474,N_7791,N_9200);
or UO_475 (O_475,N_7254,N_8697);
and UO_476 (O_476,N_5720,N_6393);
and UO_477 (O_477,N_5530,N_7879);
nand UO_478 (O_478,N_7231,N_6546);
or UO_479 (O_479,N_7312,N_5727);
xor UO_480 (O_480,N_5462,N_9157);
nand UO_481 (O_481,N_7488,N_9783);
and UO_482 (O_482,N_8912,N_7543);
nand UO_483 (O_483,N_5320,N_8561);
or UO_484 (O_484,N_7514,N_8188);
or UO_485 (O_485,N_5762,N_7922);
nand UO_486 (O_486,N_9908,N_7866);
and UO_487 (O_487,N_5840,N_9015);
nand UO_488 (O_488,N_9967,N_6907);
nor UO_489 (O_489,N_6200,N_9039);
nand UO_490 (O_490,N_7135,N_5599);
and UO_491 (O_491,N_9884,N_5862);
or UO_492 (O_492,N_8801,N_7247);
or UO_493 (O_493,N_7002,N_5215);
or UO_494 (O_494,N_8918,N_9770);
and UO_495 (O_495,N_9632,N_9888);
nand UO_496 (O_496,N_5275,N_9264);
nand UO_497 (O_497,N_6044,N_5715);
or UO_498 (O_498,N_7695,N_8261);
nor UO_499 (O_499,N_6675,N_9673);
and UO_500 (O_500,N_9325,N_8549);
nor UO_501 (O_501,N_5926,N_8836);
nand UO_502 (O_502,N_7289,N_7821);
and UO_503 (O_503,N_9010,N_8398);
nand UO_504 (O_504,N_6187,N_5086);
or UO_505 (O_505,N_7342,N_8977);
or UO_506 (O_506,N_6464,N_7916);
or UO_507 (O_507,N_8630,N_9833);
nand UO_508 (O_508,N_8118,N_9515);
nor UO_509 (O_509,N_5147,N_5113);
or UO_510 (O_510,N_7785,N_6842);
or UO_511 (O_511,N_5692,N_5017);
or UO_512 (O_512,N_8691,N_6194);
and UO_513 (O_513,N_9319,N_8309);
or UO_514 (O_514,N_8751,N_5976);
and UO_515 (O_515,N_8426,N_5435);
or UO_516 (O_516,N_9635,N_7011);
and UO_517 (O_517,N_5630,N_6193);
nand UO_518 (O_518,N_7428,N_7901);
nand UO_519 (O_519,N_5736,N_6276);
or UO_520 (O_520,N_6616,N_5980);
nor UO_521 (O_521,N_9626,N_7957);
or UO_522 (O_522,N_8163,N_5222);
or UO_523 (O_523,N_5916,N_8349);
and UO_524 (O_524,N_5133,N_9417);
nand UO_525 (O_525,N_6879,N_9799);
or UO_526 (O_526,N_5471,N_8060);
or UO_527 (O_527,N_8277,N_6202);
or UO_528 (O_528,N_5446,N_6477);
nor UO_529 (O_529,N_5904,N_9690);
or UO_530 (O_530,N_9212,N_6862);
and UO_531 (O_531,N_5637,N_8737);
nor UO_532 (O_532,N_7995,N_7137);
nor UO_533 (O_533,N_8699,N_8524);
nand UO_534 (O_534,N_8962,N_5545);
and UO_535 (O_535,N_5508,N_6039);
xor UO_536 (O_536,N_6015,N_9478);
nor UO_537 (O_537,N_6293,N_7184);
nor UO_538 (O_538,N_7738,N_5213);
nor UO_539 (O_539,N_8953,N_5850);
nand UO_540 (O_540,N_5700,N_5909);
and UO_541 (O_541,N_9842,N_5406);
and UO_542 (O_542,N_9056,N_6659);
nand UO_543 (O_543,N_6706,N_9425);
xnor UO_544 (O_544,N_7352,N_5091);
nand UO_545 (O_545,N_6595,N_6383);
nand UO_546 (O_546,N_6361,N_6666);
or UO_547 (O_547,N_6412,N_8842);
nor UO_548 (O_548,N_7303,N_8959);
nand UO_549 (O_549,N_6487,N_9383);
nand UO_550 (O_550,N_6967,N_9951);
or UO_551 (O_551,N_9229,N_9969);
and UO_552 (O_552,N_7767,N_6332);
nand UO_553 (O_553,N_5131,N_7993);
nand UO_554 (O_554,N_8854,N_9864);
or UO_555 (O_555,N_5896,N_6080);
or UO_556 (O_556,N_9629,N_8750);
nor UO_557 (O_557,N_6987,N_7589);
nand UO_558 (O_558,N_7597,N_7370);
or UO_559 (O_559,N_5457,N_6035);
or UO_560 (O_560,N_6961,N_5767);
nand UO_561 (O_561,N_7042,N_9624);
or UO_562 (O_562,N_7628,N_7701);
and UO_563 (O_563,N_8216,N_9608);
and UO_564 (O_564,N_8406,N_5385);
and UO_565 (O_565,N_7777,N_7279);
and UO_566 (O_566,N_9840,N_7196);
or UO_567 (O_567,N_7258,N_8329);
nor UO_568 (O_568,N_7670,N_6797);
or UO_569 (O_569,N_6815,N_9968);
or UO_570 (O_570,N_9820,N_7696);
nand UO_571 (O_571,N_8646,N_7983);
nor UO_572 (O_572,N_7224,N_8948);
and UO_573 (O_573,N_8641,N_5616);
or UO_574 (O_574,N_8281,N_9250);
nand UO_575 (O_575,N_9994,N_5424);
and UO_576 (O_576,N_6653,N_7014);
nand UO_577 (O_577,N_9120,N_6429);
nor UO_578 (O_578,N_7723,N_5361);
and UO_579 (O_579,N_9548,N_6300);
nand UO_580 (O_580,N_5272,N_5897);
or UO_581 (O_581,N_5695,N_6284);
or UO_582 (O_582,N_7291,N_9830);
nor UO_583 (O_583,N_6478,N_8119);
nand UO_584 (O_584,N_5752,N_6131);
nand UO_585 (O_585,N_6430,N_7783);
nor UO_586 (O_586,N_6537,N_9533);
and UO_587 (O_587,N_7358,N_9742);
and UO_588 (O_588,N_7878,N_8619);
nand UO_589 (O_589,N_9099,N_9029);
nand UO_590 (O_590,N_8694,N_5010);
and UO_591 (O_591,N_9668,N_8642);
xor UO_592 (O_592,N_9345,N_8381);
nor UO_593 (O_593,N_7408,N_5822);
or UO_594 (O_594,N_9651,N_9249);
and UO_595 (O_595,N_6504,N_7075);
and UO_596 (O_596,N_7424,N_7994);
and UO_597 (O_597,N_6799,N_6488);
and UO_598 (O_598,N_5347,N_6409);
or UO_599 (O_599,N_7026,N_9363);
and UO_600 (O_600,N_6204,N_8860);
nor UO_601 (O_601,N_5972,N_9765);
or UO_602 (O_602,N_8982,N_8623);
nor UO_603 (O_603,N_9043,N_7021);
nand UO_604 (O_604,N_7285,N_9339);
xor UO_605 (O_605,N_6981,N_5774);
or UO_606 (O_606,N_9090,N_8058);
nand UO_607 (O_607,N_7828,N_9764);
and UO_608 (O_608,N_7063,N_7381);
nor UO_609 (O_609,N_7897,N_6245);
and UO_610 (O_610,N_8373,N_7961);
or UO_611 (O_611,N_9176,N_8018);
nand UO_612 (O_612,N_8429,N_8894);
or UO_613 (O_613,N_5873,N_9754);
nor UO_614 (O_614,N_6343,N_5019);
nand UO_615 (O_615,N_7235,N_5883);
nand UO_616 (O_616,N_9634,N_8584);
nor UO_617 (O_617,N_9290,N_6455);
nor UO_618 (O_618,N_6848,N_7898);
nand UO_619 (O_619,N_5209,N_6870);
nand UO_620 (O_620,N_5698,N_9691);
or UO_621 (O_621,N_8011,N_9219);
or UO_622 (O_622,N_9035,N_5819);
and UO_623 (O_623,N_7206,N_9150);
or UO_624 (O_624,N_9366,N_8526);
or UO_625 (O_625,N_9895,N_6491);
nand UO_626 (O_626,N_8757,N_5290);
or UO_627 (O_627,N_5564,N_5136);
and UO_628 (O_628,N_8618,N_8066);
and UO_629 (O_629,N_8794,N_6108);
nand UO_630 (O_630,N_6578,N_8105);
nand UO_631 (O_631,N_7619,N_5627);
and UO_632 (O_632,N_8915,N_8296);
nand UO_633 (O_633,N_6638,N_7028);
nor UO_634 (O_634,N_7508,N_8859);
nor UO_635 (O_635,N_5228,N_5390);
xnor UO_636 (O_636,N_5282,N_7786);
nor UO_637 (O_637,N_5117,N_8190);
and UO_638 (O_638,N_7102,N_7664);
nor UO_639 (O_639,N_8001,N_6539);
nand UO_640 (O_640,N_6378,N_6730);
or UO_641 (O_641,N_5729,N_8939);
nand UO_642 (O_642,N_6012,N_7833);
nand UO_643 (O_643,N_8519,N_8825);
and UO_644 (O_644,N_9853,N_9546);
or UO_645 (O_645,N_9553,N_8010);
nand UO_646 (O_646,N_7473,N_5533);
nand UO_647 (O_647,N_6770,N_9110);
and UO_648 (O_648,N_5170,N_5557);
and UO_649 (O_649,N_7880,N_5001);
or UO_650 (O_650,N_6228,N_7380);
nor UO_651 (O_651,N_8171,N_9834);
and UO_652 (O_652,N_9310,N_7761);
or UO_653 (O_653,N_9076,N_9027);
or UO_654 (O_654,N_8647,N_7928);
nand UO_655 (O_655,N_5901,N_6936);
nand UO_656 (O_656,N_7614,N_6177);
nand UO_657 (O_657,N_6604,N_7774);
and UO_658 (O_658,N_5221,N_8287);
nor UO_659 (O_659,N_7104,N_5566);
or UO_660 (O_660,N_9252,N_8499);
nor UO_661 (O_661,N_7747,N_8046);
and UO_662 (O_662,N_7087,N_5967);
nor UO_663 (O_663,N_9936,N_6191);
and UO_664 (O_664,N_9195,N_7344);
nand UO_665 (O_665,N_8759,N_6253);
and UO_666 (O_666,N_8404,N_9711);
xnor UO_667 (O_667,N_5146,N_7094);
nor UO_668 (O_668,N_6549,N_7017);
and UO_669 (O_669,N_9450,N_6762);
nor UO_670 (O_670,N_9453,N_6346);
nand UO_671 (O_671,N_6408,N_6746);
nor UO_672 (O_672,N_6096,N_8420);
nor UO_673 (O_673,N_6787,N_8890);
nand UO_674 (O_674,N_5397,N_7566);
nand UO_675 (O_675,N_7889,N_5439);
nor UO_676 (O_676,N_5952,N_5921);
and UO_677 (O_677,N_5261,N_9490);
nor UO_678 (O_678,N_7958,N_9746);
nand UO_679 (O_679,N_7168,N_5608);
nand UO_680 (O_680,N_5761,N_9956);
and UO_681 (O_681,N_5399,N_6745);
nor UO_682 (O_682,N_7923,N_7464);
or UO_683 (O_683,N_6143,N_5263);
nand UO_684 (O_684,N_6394,N_7034);
or UO_685 (O_685,N_9960,N_8754);
nor UO_686 (O_686,N_6619,N_9174);
and UO_687 (O_687,N_5276,N_6726);
or UO_688 (O_688,N_7606,N_5864);
or UO_689 (O_689,N_6218,N_8272);
nor UO_690 (O_690,N_6020,N_9342);
xnor UO_691 (O_691,N_6246,N_8654);
nand UO_692 (O_692,N_8807,N_6385);
or UO_693 (O_693,N_8434,N_7164);
nor UO_694 (O_694,N_7309,N_7790);
nor UO_695 (O_695,N_6676,N_5499);
or UO_696 (O_696,N_7499,N_8814);
or UO_697 (O_697,N_8040,N_7058);
and UO_698 (O_698,N_9819,N_6079);
and UO_699 (O_699,N_5996,N_7787);
and UO_700 (O_700,N_6581,N_9774);
nor UO_701 (O_701,N_9512,N_7779);
nand UO_702 (O_702,N_5537,N_7117);
and UO_703 (O_703,N_7230,N_8074);
and UO_704 (O_704,N_7863,N_9031);
or UO_705 (O_705,N_5751,N_6369);
and UO_706 (O_706,N_6727,N_5013);
nor UO_707 (O_707,N_9591,N_9940);
or UO_708 (O_708,N_6943,N_7313);
or UO_709 (O_709,N_5623,N_7445);
or UO_710 (O_710,N_8649,N_7477);
or UO_711 (O_711,N_9689,N_5870);
nand UO_712 (O_712,N_7163,N_8114);
nor UO_713 (O_713,N_8856,N_7084);
or UO_714 (O_714,N_6895,N_7936);
or UO_715 (O_715,N_6796,N_6687);
nand UO_716 (O_716,N_6975,N_5452);
and UO_717 (O_717,N_6855,N_7260);
nand UO_718 (O_718,N_6032,N_8791);
nand UO_719 (O_719,N_5386,N_5256);
nand UO_720 (O_720,N_8984,N_8886);
nand UO_721 (O_721,N_8196,N_9862);
or UO_722 (O_722,N_8515,N_7666);
or UO_723 (O_723,N_5437,N_9182);
or UO_724 (O_724,N_8883,N_7534);
nor UO_725 (O_725,N_9348,N_6519);
or UO_726 (O_726,N_7435,N_9451);
or UO_727 (O_727,N_6933,N_6527);
and UO_728 (O_728,N_8955,N_8059);
and UO_729 (O_729,N_7226,N_7844);
nand UO_730 (O_730,N_6765,N_8587);
or UO_731 (O_731,N_9047,N_7908);
nor UO_732 (O_732,N_5852,N_6043);
and UO_733 (O_733,N_8182,N_9973);
or UO_734 (O_734,N_5994,N_6055);
and UO_735 (O_735,N_9924,N_6716);
nand UO_736 (O_736,N_9053,N_5764);
or UO_737 (O_737,N_7574,N_5887);
nand UO_738 (O_738,N_8487,N_9977);
nand UO_739 (O_739,N_5249,N_7511);
nor UO_740 (O_740,N_8987,N_5848);
nor UO_741 (O_741,N_8711,N_7895);
nor UO_742 (O_742,N_9160,N_6683);
and UO_743 (O_743,N_6389,N_6470);
or UO_744 (O_744,N_6679,N_9471);
or UO_745 (O_745,N_8667,N_7086);
nor UO_746 (O_746,N_8226,N_5478);
xnor UO_747 (O_747,N_6615,N_9859);
nand UO_748 (O_748,N_7364,N_5826);
and UO_749 (O_749,N_6823,N_8084);
nor UO_750 (O_750,N_5238,N_7448);
nor UO_751 (O_751,N_5845,N_7280);
and UO_752 (O_752,N_7642,N_8862);
nand UO_753 (O_753,N_7618,N_7621);
nor UO_754 (O_754,N_9173,N_9154);
and UO_755 (O_755,N_9927,N_6084);
nand UO_756 (O_756,N_6494,N_7854);
nor UO_757 (O_757,N_8966,N_5183);
and UO_758 (O_758,N_8710,N_9413);
and UO_759 (O_759,N_8762,N_9721);
and UO_760 (O_760,N_9036,N_5162);
and UO_761 (O_761,N_7433,N_5963);
nor UO_762 (O_762,N_9999,N_9719);
nand UO_763 (O_763,N_6927,N_8921);
nand UO_764 (O_764,N_6768,N_8885);
and UO_765 (O_765,N_8930,N_7403);
or UO_766 (O_766,N_9081,N_5049);
or UO_767 (O_767,N_6190,N_5861);
or UO_768 (O_768,N_5267,N_6338);
nand UO_769 (O_769,N_6416,N_9284);
nor UO_770 (O_770,N_6413,N_7977);
and UO_771 (O_771,N_8477,N_5237);
xnor UO_772 (O_772,N_7421,N_9790);
nand UO_773 (O_773,N_7690,N_9793);
xnor UO_774 (O_774,N_9899,N_8152);
nand UO_775 (O_775,N_8165,N_9017);
xnor UO_776 (O_776,N_5407,N_5755);
nand UO_777 (O_777,N_8878,N_8496);
nand UO_778 (O_778,N_7806,N_7182);
nor UO_779 (O_779,N_5710,N_9487);
nand UO_780 (O_780,N_5625,N_9659);
nand UO_781 (O_781,N_5642,N_9012);
and UO_782 (O_782,N_5364,N_5568);
nand UO_783 (O_783,N_5266,N_5043);
and UO_784 (O_784,N_7676,N_8829);
nor UO_785 (O_785,N_5024,N_8376);
or UO_786 (O_786,N_6763,N_5022);
nor UO_787 (O_787,N_6325,N_7031);
or UO_788 (O_788,N_6355,N_6392);
and UO_789 (O_789,N_8572,N_6985);
and UO_790 (O_790,N_8148,N_6814);
nor UO_791 (O_791,N_9972,N_9491);
and UO_792 (O_792,N_7204,N_8364);
and UO_793 (O_793,N_5900,N_7659);
nor UO_794 (O_794,N_6052,N_6460);
nor UO_795 (O_795,N_9272,N_8910);
xnor UO_796 (O_796,N_8347,N_5573);
and UO_797 (O_797,N_9771,N_8696);
nand UO_798 (O_798,N_6379,N_6714);
nand UO_799 (O_799,N_5167,N_7141);
nor UO_800 (O_800,N_9333,N_8089);
or UO_801 (O_801,N_9415,N_5771);
or UO_802 (O_802,N_7605,N_7138);
nand UO_803 (O_803,N_9743,N_5691);
nor UO_804 (O_804,N_9430,N_7815);
nand UO_805 (O_805,N_9414,N_9759);
xnor UO_806 (O_806,N_5417,N_7564);
xor UO_807 (O_807,N_6724,N_7097);
nand UO_808 (O_808,N_9909,N_9653);
nor UO_809 (O_809,N_6583,N_9736);
or UO_810 (O_810,N_8411,N_6213);
or UO_811 (O_811,N_8344,N_6161);
nor UO_812 (O_812,N_6345,N_5274);
and UO_813 (O_813,N_7810,N_8494);
nor UO_814 (O_814,N_9616,N_6445);
xnor UO_815 (O_815,N_6526,N_6913);
nor UO_816 (O_816,N_8944,N_8315);
nand UO_817 (O_817,N_6384,N_5498);
nand UO_818 (O_818,N_9428,N_5763);
and UO_819 (O_819,N_5708,N_8362);
and UO_820 (O_820,N_9605,N_5538);
nand UO_821 (O_821,N_7046,N_6057);
or UO_822 (O_822,N_6845,N_9688);
and UO_823 (O_823,N_8162,N_8206);
and UO_824 (O_824,N_7653,N_8928);
and UO_825 (O_825,N_9657,N_8571);
nand UO_826 (O_826,N_8229,N_9159);
nand UO_827 (O_827,N_6811,N_9886);
nand UO_828 (O_828,N_7491,N_5973);
or UO_829 (O_829,N_6589,N_9677);
or UO_830 (O_830,N_7057,N_6189);
and UO_831 (O_831,N_7167,N_9685);
nor UO_832 (O_832,N_5059,N_9445);
and UO_833 (O_833,N_5859,N_5155);
or UO_834 (O_834,N_6742,N_9778);
nand UO_835 (O_835,N_5201,N_8463);
nor UO_836 (O_836,N_5084,N_6836);
or UO_837 (O_837,N_8095,N_7233);
nand UO_838 (O_838,N_6474,N_9809);
nor UO_839 (O_839,N_5529,N_5808);
nor UO_840 (O_840,N_5869,N_7560);
and UO_841 (O_841,N_7237,N_6133);
nand UO_842 (O_842,N_6697,N_9481);
and UO_843 (O_843,N_5319,N_7241);
nor UO_844 (O_844,N_6827,N_6125);
or UO_845 (O_845,N_8525,N_5646);
or UO_846 (O_846,N_8905,N_7029);
nor UO_847 (O_847,N_5828,N_5950);
xor UO_848 (O_848,N_6279,N_5418);
xor UO_849 (O_849,N_8940,N_7538);
nand UO_850 (O_850,N_8790,N_9587);
and UO_851 (O_851,N_5659,N_9603);
nand UO_852 (O_852,N_9214,N_6505);
or UO_853 (O_853,N_9231,N_7278);
nor UO_854 (O_854,N_8157,N_9023);
and UO_855 (O_855,N_5148,N_5492);
xnor UO_856 (O_856,N_5560,N_8612);
and UO_857 (O_857,N_8924,N_7809);
nor UO_858 (O_858,N_8739,N_6903);
and UO_859 (O_859,N_6497,N_5322);
nand UO_860 (O_860,N_7022,N_5181);
or UO_861 (O_861,N_8268,N_9164);
nand UO_862 (O_862,N_6219,N_9286);
nor UO_863 (O_863,N_8769,N_7305);
or UO_864 (O_864,N_7991,N_8950);
nand UO_865 (O_865,N_8126,N_7413);
and UO_866 (O_866,N_7813,N_9869);
nor UO_867 (O_867,N_9542,N_9705);
nand UO_868 (O_868,N_8416,N_6447);
nor UO_869 (O_869,N_7823,N_5798);
or UO_870 (O_870,N_9558,N_6535);
nand UO_871 (O_871,N_7608,N_9262);
xor UO_872 (O_872,N_6082,N_9181);
or UO_873 (O_873,N_8747,N_9726);
and UO_874 (O_874,N_5759,N_9680);
nand UO_875 (O_875,N_7740,N_9100);
or UO_876 (O_876,N_8631,N_8249);
nand UO_877 (O_877,N_7782,N_6117);
nand UO_878 (O_878,N_5171,N_7065);
nor UO_879 (O_879,N_9925,N_9216);
nand UO_880 (O_880,N_8846,N_9597);
and UO_881 (O_881,N_6607,N_8061);
xnor UO_882 (O_882,N_8080,N_8259);
or UO_883 (O_883,N_7484,N_7572);
nand UO_884 (O_884,N_7555,N_9140);
nand UO_885 (O_885,N_5680,N_9069);
or UO_886 (O_886,N_9552,N_9507);
nand UO_887 (O_887,N_8193,N_9025);
nand UO_888 (O_888,N_6613,N_8720);
and UO_889 (O_889,N_8923,N_6813);
nor UO_890 (O_890,N_5598,N_8250);
or UO_891 (O_891,N_5085,N_6533);
and UO_892 (O_892,N_7988,N_8563);
and UO_893 (O_893,N_6169,N_5490);
or UO_894 (O_894,N_8611,N_8613);
or UO_895 (O_895,N_7631,N_9804);
nor UO_896 (O_896,N_8512,N_8402);
and UO_897 (O_897,N_7269,N_6818);
nor UO_898 (O_898,N_5000,N_8956);
and UO_899 (O_899,N_8351,N_9180);
or UO_900 (O_900,N_9612,N_7067);
nand UO_901 (O_901,N_9233,N_8604);
and UO_902 (O_902,N_7153,N_7892);
nor UO_903 (O_903,N_5415,N_8900);
and UO_904 (O_904,N_6512,N_8107);
nand UO_905 (O_905,N_7110,N_6794);
nor UO_906 (O_906,N_8378,N_5231);
nor UO_907 (O_907,N_6492,N_9952);
nand UO_908 (O_908,N_6421,N_5886);
or UO_909 (O_909,N_9165,N_7900);
nand UO_910 (O_910,N_7426,N_7853);
and UO_911 (O_911,N_9729,N_9008);
nor UO_912 (O_912,N_7294,N_8151);
or UO_913 (O_913,N_6217,N_6834);
nor UO_914 (O_914,N_7156,N_9949);
or UO_915 (O_915,N_7829,N_8719);
and UO_916 (O_916,N_9305,N_7663);
nor UO_917 (O_917,N_9024,N_5048);
and UO_918 (O_918,N_7338,N_5192);
nor UO_919 (O_919,N_5393,N_8785);
nand UO_920 (O_920,N_9995,N_9221);
nor UO_921 (O_921,N_7283,N_9509);
nand UO_922 (O_922,N_8889,N_6557);
nor UO_923 (O_923,N_9751,N_9326);
or UO_924 (O_924,N_7320,N_8258);
nand UO_925 (O_925,N_9331,N_5944);
or UO_926 (O_926,N_9572,N_6624);
nand UO_927 (O_927,N_8012,N_8092);
xor UO_928 (O_928,N_5038,N_9155);
and UO_929 (O_929,N_6594,N_7502);
and UO_930 (O_930,N_8576,N_6422);
or UO_931 (O_931,N_5552,N_6100);
or UO_932 (O_932,N_8136,N_7114);
nor UO_933 (O_933,N_9420,N_6208);
and UO_934 (O_934,N_8146,N_5464);
nand UO_935 (O_935,N_6337,N_7444);
nand UO_936 (O_936,N_6398,N_6210);
or UO_937 (O_937,N_7671,N_7319);
and UO_938 (O_938,N_6341,N_9532);
and UO_939 (O_939,N_9792,N_7567);
or UO_940 (O_940,N_5389,N_8235);
or UO_941 (O_941,N_6597,N_9932);
nor UO_942 (O_942,N_8993,N_5649);
nor UO_943 (O_943,N_6249,N_5230);
nand UO_944 (O_944,N_8902,N_5823);
nor UO_945 (O_945,N_7321,N_6632);
nand UO_946 (O_946,N_8695,N_8617);
and UO_947 (O_947,N_8578,N_7256);
nor UO_948 (O_948,N_8875,N_5988);
or UO_949 (O_949,N_5542,N_6956);
nand UO_950 (O_950,N_8314,N_6342);
or UO_951 (O_951,N_9385,N_5957);
or UO_952 (O_952,N_7044,N_9343);
or UO_953 (O_953,N_9393,N_7950);
and UO_954 (O_954,N_7270,N_7257);
nand UO_955 (O_955,N_6806,N_9523);
and UO_956 (O_956,N_5208,N_5905);
nor UO_957 (O_957,N_5053,N_5528);
or UO_958 (O_958,N_8180,N_6997);
nor UO_959 (O_959,N_7954,N_6286);
nand UO_960 (O_960,N_5706,N_8881);
or UO_961 (O_961,N_7655,N_6639);
nand UO_962 (O_962,N_6810,N_6520);
and UO_963 (O_963,N_6650,N_5684);
nand UO_964 (O_964,N_8580,N_8816);
nand UO_965 (O_965,N_8721,N_7580);
nand UO_966 (O_966,N_9779,N_5430);
xor UO_967 (O_967,N_6289,N_5713);
or UO_968 (O_968,N_8044,N_9992);
xnor UO_969 (O_969,N_5874,N_7064);
nor UO_970 (O_970,N_8145,N_9472);
nor UO_971 (O_971,N_6759,N_6873);
nand UO_972 (O_972,N_7098,N_6452);
nand UO_973 (O_973,N_9601,N_6574);
and UO_974 (O_974,N_9192,N_8545);
nand UO_975 (O_975,N_7223,N_9189);
xnor UO_976 (O_976,N_8552,N_8511);
or UO_977 (O_977,N_5610,N_7188);
nand UO_978 (O_978,N_9184,N_7912);
or UO_979 (O_979,N_5626,N_5717);
xor UO_980 (O_980,N_9404,N_6782);
nor UO_981 (O_981,N_8896,N_9274);
or UO_982 (O_982,N_8774,N_9520);
and UO_983 (O_983,N_9596,N_8031);
nor UO_984 (O_984,N_8473,N_5491);
and UO_985 (O_985,N_6940,N_8819);
nor UO_986 (O_986,N_7811,N_8855);
or UO_987 (O_987,N_8508,N_5394);
nor UO_988 (O_988,N_7714,N_6209);
nand UO_989 (O_989,N_5246,N_8194);
or UO_990 (O_990,N_9666,N_9304);
or UO_991 (O_991,N_6902,N_7634);
or UO_992 (O_992,N_5433,N_8756);
nor UO_993 (O_993,N_9438,N_5550);
nand UO_994 (O_994,N_7366,N_8958);
nor UO_995 (O_995,N_9957,N_5184);
and UO_996 (O_996,N_5895,N_8275);
or UO_997 (O_997,N_5645,N_5685);
xnor UO_998 (O_998,N_8015,N_5199);
nor UO_999 (O_999,N_8784,N_9983);
or UO_1000 (O_1000,N_8007,N_9530);
and UO_1001 (O_1001,N_5531,N_9646);
or UO_1002 (O_1002,N_5655,N_8289);
xor UO_1003 (O_1003,N_8039,N_9620);
nand UO_1004 (O_1004,N_9295,N_8882);
nand UO_1005 (O_1005,N_7841,N_8143);
nor UO_1006 (O_1006,N_5635,N_5785);
nand UO_1007 (O_1007,N_8384,N_6174);
and UO_1008 (O_1008,N_8199,N_7343);
and UO_1009 (O_1009,N_5678,N_9013);
nand UO_1010 (O_1010,N_7331,N_8919);
nand UO_1011 (O_1011,N_9357,N_9215);
or UO_1012 (O_1012,N_6725,N_9676);
and UO_1013 (O_1013,N_5998,N_9815);
and UO_1014 (O_1014,N_7544,N_8551);
and UO_1015 (O_1015,N_5207,N_7978);
nor UO_1016 (O_1016,N_6334,N_6226);
nand UO_1017 (O_1017,N_8482,N_9454);
nor UO_1018 (O_1018,N_6297,N_9637);
nor UO_1019 (O_1019,N_5579,N_7939);
and UO_1020 (O_1020,N_7450,N_7604);
nor UO_1021 (O_1021,N_8833,N_5269);
or UO_1022 (O_1022,N_6736,N_5414);
and UO_1023 (O_1023,N_5953,N_8911);
nand UO_1024 (O_1024,N_7192,N_5565);
nor UO_1025 (O_1025,N_7795,N_9054);
or UO_1026 (O_1026,N_5844,N_5003);
nand UO_1027 (O_1027,N_7585,N_7298);
nand UO_1028 (O_1028,N_8665,N_6523);
and UO_1029 (O_1029,N_9803,N_9614);
nand UO_1030 (O_1030,N_6352,N_8391);
or UO_1031 (O_1031,N_9276,N_7986);
or UO_1032 (O_1032,N_7475,N_8693);
nor UO_1033 (O_1033,N_5624,N_6259);
or UO_1034 (O_1034,N_5851,N_9700);
nand UO_1035 (O_1035,N_5581,N_6083);
or UO_1036 (O_1036,N_5791,N_6427);
nand UO_1037 (O_1037,N_8738,N_5449);
and UO_1038 (O_1038,N_6232,N_5039);
nor UO_1039 (O_1039,N_5214,N_5396);
nor UO_1040 (O_1040,N_7697,N_7452);
or UO_1041 (O_1041,N_9675,N_5429);
and UO_1042 (O_1042,N_9647,N_9125);
or UO_1043 (O_1043,N_5254,N_9193);
xnor UO_1044 (O_1044,N_5158,N_7733);
nor UO_1045 (O_1045,N_7329,N_8979);
and UO_1046 (O_1046,N_9230,N_9113);
nor UO_1047 (O_1047,N_8115,N_9543);
and UO_1048 (O_1048,N_7999,N_7682);
or UO_1049 (O_1049,N_8992,N_5948);
or UO_1050 (O_1050,N_6920,N_8834);
nand UO_1051 (O_1051,N_6086,N_9814);
and UO_1052 (O_1052,N_6654,N_7051);
nand UO_1053 (O_1053,N_7264,N_9241);
or UO_1054 (O_1054,N_9365,N_5018);
or UO_1055 (O_1055,N_6046,N_8295);
and UO_1056 (O_1056,N_8941,N_9724);
nand UO_1057 (O_1057,N_7197,N_7099);
xnor UO_1058 (O_1058,N_7794,N_8840);
or UO_1059 (O_1059,N_9800,N_5465);
and UO_1060 (O_1060,N_7920,N_8077);
nand UO_1061 (O_1061,N_7855,N_9104);
nand UO_1062 (O_1062,N_8017,N_5820);
nor UO_1063 (O_1063,N_6237,N_7857);
or UO_1064 (O_1064,N_5756,N_8786);
or UO_1065 (O_1065,N_7814,N_8176);
and UO_1066 (O_1066,N_9486,N_5639);
nand UO_1067 (O_1067,N_5753,N_8380);
and UO_1068 (O_1068,N_5012,N_6006);
and UO_1069 (O_1069,N_8539,N_5448);
nand UO_1070 (O_1070,N_7633,N_7931);
and UO_1071 (O_1071,N_6110,N_9892);
or UO_1072 (O_1072,N_8045,N_6444);
or UO_1073 (O_1073,N_9433,N_8852);
and UO_1074 (O_1074,N_5308,N_6005);
nand UO_1075 (O_1075,N_5015,N_6465);
and UO_1076 (O_1076,N_9511,N_9052);
nand UO_1077 (O_1077,N_8964,N_5189);
and UO_1078 (O_1078,N_9362,N_8189);
xor UO_1079 (O_1079,N_8297,N_7465);
or UO_1080 (O_1080,N_6816,N_5793);
or UO_1081 (O_1081,N_8352,N_5681);
or UO_1082 (O_1082,N_5127,N_8431);
or UO_1083 (O_1083,N_6753,N_9880);
nand UO_1084 (O_1084,N_6973,N_6785);
or UO_1085 (O_1085,N_7976,N_5358);
and UO_1086 (O_1086,N_7951,N_9369);
or UO_1087 (O_1087,N_6065,N_6801);
or UO_1088 (O_1088,N_8705,N_6518);
nor UO_1089 (O_1089,N_9317,N_7679);
and UO_1090 (O_1090,N_7103,N_8672);
nand UO_1091 (O_1091,N_7650,N_8771);
and UO_1092 (O_1092,N_5797,N_6148);
nand UO_1093 (O_1093,N_6889,N_8868);
nand UO_1094 (O_1094,N_8768,N_8869);
and UO_1095 (O_1095,N_9761,N_8202);
and UO_1096 (O_1096,N_9371,N_8085);
and UO_1097 (O_1097,N_8971,N_8758);
nand UO_1098 (O_1098,N_9713,N_7941);
xnor UO_1099 (O_1099,N_6969,N_9308);
nand UO_1100 (O_1100,N_8983,N_8022);
nor UO_1101 (O_1101,N_9243,N_9026);
nand UO_1102 (O_1102,N_7015,N_6731);
or UO_1103 (O_1103,N_5129,N_8213);
nand UO_1104 (O_1104,N_6678,N_6331);
nor UO_1105 (O_1105,N_6381,N_5126);
or UO_1106 (O_1106,N_9148,N_9199);
nand UO_1107 (O_1107,N_6554,N_9149);
nor UO_1108 (O_1108,N_5289,N_6550);
nor UO_1109 (O_1109,N_5954,N_9364);
or UO_1110 (O_1110,N_5441,N_8644);
nor UO_1111 (O_1111,N_5965,N_9655);
nor UO_1112 (O_1112,N_7734,N_8301);
and UO_1113 (O_1113,N_5687,N_5782);
and UO_1114 (O_1114,N_6397,N_9554);
or UO_1115 (O_1115,N_5140,N_8748);
or UO_1116 (O_1116,N_7559,N_8588);
nand UO_1117 (O_1117,N_5534,N_5589);
nor UO_1118 (O_1118,N_6506,N_6307);
nor UO_1119 (O_1119,N_6798,N_9476);
nand UO_1120 (O_1120,N_8615,N_6875);
and UO_1121 (O_1121,N_7685,N_5749);
or UO_1122 (O_1122,N_7756,N_8357);
and UO_1123 (O_1123,N_6837,N_6772);
and UO_1124 (O_1124,N_7093,N_8655);
and UO_1125 (O_1125,N_5348,N_8361);
nor UO_1126 (O_1126,N_6102,N_6033);
and UO_1127 (O_1127,N_8817,N_8985);
nand UO_1128 (O_1128,N_7677,N_5381);
nand UO_1129 (O_1129,N_8292,N_7867);
and UO_1130 (O_1130,N_9517,N_6846);
nand UO_1131 (O_1131,N_9321,N_5422);
nor UO_1132 (O_1132,N_6641,N_5034);
and UO_1133 (O_1133,N_8142,N_7992);
and UO_1134 (O_1134,N_7170,N_7535);
nand UO_1135 (O_1135,N_6609,N_7539);
nor UO_1136 (O_1136,N_9618,N_8810);
nor UO_1137 (O_1137,N_9550,N_8088);
and UO_1138 (O_1138,N_6313,N_9135);
or UO_1139 (O_1139,N_6304,N_8322);
nor UO_1140 (O_1140,N_7703,N_5335);
and UO_1141 (O_1141,N_9434,N_6734);
xor UO_1142 (O_1142,N_6702,N_6541);
nor UO_1143 (O_1143,N_6146,N_5374);
nand UO_1144 (O_1144,N_7356,N_6922);
and UO_1145 (O_1145,N_9622,N_9107);
or UO_1146 (O_1146,N_5813,N_9521);
or UO_1147 (O_1147,N_9623,N_7249);
or UO_1148 (O_1148,N_8514,N_7244);
and UO_1149 (O_1149,N_6114,N_9625);
or UO_1150 (O_1150,N_6829,N_7969);
and UO_1151 (O_1151,N_6553,N_5477);
nor UO_1152 (O_1152,N_9513,N_6348);
nand UO_1153 (O_1153,N_5548,N_6781);
xor UO_1154 (O_1154,N_6992,N_9287);
or UO_1155 (O_1155,N_5456,N_6432);
nand UO_1156 (O_1156,N_6534,N_5596);
nor UO_1157 (O_1157,N_8933,N_6674);
nor UO_1158 (O_1158,N_8568,N_6134);
nand UO_1159 (O_1159,N_6998,N_8082);
or UO_1160 (O_1160,N_9089,N_9059);
nand UO_1161 (O_1161,N_6808,N_8895);
or UO_1162 (O_1162,N_9256,N_6031);
or UO_1163 (O_1163,N_8479,N_5367);
or UO_1164 (O_1164,N_7503,N_6915);
xnor UO_1165 (O_1165,N_9979,N_7020);
nand UO_1166 (O_1166,N_5176,N_7133);
nor UO_1167 (O_1167,N_9209,N_7354);
and UO_1168 (O_1168,N_6719,N_7627);
and UO_1169 (O_1169,N_8744,N_5029);
nand UO_1170 (O_1170,N_6977,N_8166);
nand UO_1171 (O_1171,N_9749,N_7259);
and UO_1172 (O_1172,N_7175,N_6540);
nor UO_1173 (O_1173,N_6363,N_6972);
or UO_1174 (O_1174,N_8288,N_5014);
nor UO_1175 (O_1175,N_7405,N_7095);
nand UO_1176 (O_1176,N_7225,N_5876);
and UO_1177 (O_1177,N_7265,N_7662);
nand UO_1178 (O_1178,N_6489,N_9372);
nand UO_1179 (O_1179,N_9559,N_6847);
and UO_1180 (O_1180,N_9303,N_5739);
nand UO_1181 (O_1181,N_6789,N_6233);
and UO_1182 (O_1182,N_7638,N_8505);
and UO_1183 (O_1183,N_6860,N_8443);
nand UO_1184 (O_1184,N_8214,N_6744);
or UO_1185 (O_1185,N_9041,N_7746);
nor UO_1186 (O_1186,N_6485,N_5938);
and UO_1187 (O_1187,N_8121,N_5412);
and UO_1188 (O_1188,N_5072,N_8565);
nor UO_1189 (O_1189,N_5940,N_8198);
nor UO_1190 (O_1190,N_6906,N_7706);
or UO_1191 (O_1191,N_9163,N_7987);
nor UO_1192 (O_1192,N_8675,N_6777);
or UO_1193 (O_1193,N_9671,N_8715);
and UO_1194 (O_1194,N_6901,N_6996);
or UO_1195 (O_1195,N_7106,N_8684);
nor UO_1196 (O_1196,N_5721,N_7617);
nor UO_1197 (O_1197,N_5683,N_6579);
or UO_1198 (O_1198,N_6517,N_7864);
or UO_1199 (O_1199,N_8724,N_9918);
nand UO_1200 (O_1200,N_7837,N_6137);
and UO_1201 (O_1201,N_6333,N_7765);
and UO_1202 (O_1202,N_9946,N_7429);
nor UO_1203 (O_1203,N_7667,N_8636);
or UO_1204 (O_1204,N_9914,N_7698);
nand UO_1205 (O_1205,N_5137,N_5760);
or UO_1206 (O_1206,N_7050,N_9788);
nor UO_1207 (O_1207,N_6074,N_6866);
or UO_1208 (O_1208,N_6036,N_8577);
and UO_1209 (O_1209,N_6360,N_5612);
nor UO_1210 (O_1210,N_9714,N_7570);
or UO_1211 (O_1211,N_8220,N_7369);
and UO_1212 (O_1212,N_7070,N_5487);
or UO_1213 (O_1213,N_6617,N_8803);
nor UO_1214 (O_1214,N_6471,N_9139);
xnor UO_1215 (O_1215,N_9656,N_7781);
nor UO_1216 (O_1216,N_9844,N_5554);
nor UO_1217 (O_1217,N_8150,N_5283);
and UO_1218 (O_1218,N_5986,N_6101);
or UO_1219 (O_1219,N_8632,N_5164);
or UO_1220 (O_1220,N_6575,N_6225);
nor UO_1221 (O_1221,N_9941,N_7720);
nand UO_1222 (O_1222,N_5006,N_6897);
nor UO_1223 (O_1223,N_7425,N_8444);
and UO_1224 (O_1224,N_8712,N_7552);
nand UO_1225 (O_1225,N_9065,N_6404);
nor UO_1226 (O_1226,N_5920,N_5741);
and UO_1227 (O_1227,N_5317,N_5326);
and UO_1228 (O_1228,N_7100,N_8428);
nor UO_1229 (O_1229,N_6336,N_5878);
and UO_1230 (O_1230,N_9311,N_6411);
nor UO_1231 (O_1231,N_5699,N_5804);
and UO_1232 (O_1232,N_7970,N_9177);
and UO_1233 (O_1233,N_9337,N_5525);
nor UO_1234 (O_1234,N_9298,N_7515);
or UO_1235 (O_1235,N_6824,N_7101);
and UO_1236 (O_1236,N_7527,N_9701);
nor UO_1237 (O_1237,N_8787,N_9867);
and UO_1238 (O_1238,N_7219,N_9227);
nand UO_1239 (O_1239,N_5773,N_7586);
and UO_1240 (O_1240,N_9461,N_5519);
and UO_1241 (O_1241,N_8346,N_6203);
nand UO_1242 (O_1242,N_5083,N_6266);
nand UO_1243 (O_1243,N_8436,N_9185);
nor UO_1244 (O_1244,N_6025,N_9854);
and UO_1245 (O_1245,N_8800,N_9708);
or UO_1246 (O_1246,N_6844,N_6952);
nand UO_1247 (O_1247,N_7526,N_8123);
nor UO_1248 (O_1248,N_6156,N_6514);
nand UO_1249 (O_1249,N_7494,N_9738);
nor UO_1250 (O_1250,N_5251,N_7562);
nor UO_1251 (O_1251,N_7193,N_5360);
nor UO_1252 (O_1252,N_7949,N_6832);
nand UO_1253 (O_1253,N_9506,N_6019);
nand UO_1254 (O_1254,N_8442,N_9358);
nor UO_1255 (O_1255,N_6707,N_7322);
and UO_1256 (O_1256,N_6547,N_8138);
and UO_1257 (O_1257,N_6106,N_6723);
xor UO_1258 (O_1258,N_6865,N_9000);
nor UO_1259 (O_1259,N_8614,N_6314);
nand UO_1260 (O_1260,N_6382,N_6155);
nand UO_1261 (O_1261,N_8931,N_6295);
nor UO_1262 (O_1262,N_6694,N_7334);
nor UO_1263 (O_1263,N_9320,N_5618);
or UO_1264 (O_1264,N_6239,N_5342);
nor UO_1265 (O_1265,N_9265,N_7072);
nor UO_1266 (O_1266,N_5517,N_5838);
and UO_1267 (O_1267,N_7827,N_7200);
or UO_1268 (O_1268,N_9283,N_6351);
nor UO_1269 (O_1269,N_5278,N_8909);
nor UO_1270 (O_1270,N_6040,N_8778);
nor UO_1271 (O_1271,N_9374,N_8907);
or UO_1272 (O_1272,N_6165,N_8586);
and UO_1273 (O_1273,N_9218,N_5867);
nand UO_1274 (O_1274,N_7282,N_6925);
nand UO_1275 (O_1275,N_9641,N_6739);
and UO_1276 (O_1276,N_5211,N_7884);
nand UO_1277 (O_1277,N_7744,N_7645);
nor UO_1278 (O_1278,N_7411,N_5191);
nand UO_1279 (O_1279,N_7549,N_7496);
nand UO_1280 (O_1280,N_6729,N_8184);
and UO_1281 (O_1281,N_7868,N_9327);
nand UO_1282 (O_1282,N_5872,N_9516);
or UO_1283 (O_1283,N_7541,N_5493);
or UO_1284 (O_1284,N_9072,N_5108);
or UO_1285 (O_1285,N_8804,N_5509);
nor UO_1286 (O_1286,N_5527,N_7717);
or UO_1287 (O_1287,N_9332,N_8124);
nor UO_1288 (O_1288,N_9562,N_6260);
nor UO_1289 (O_1289,N_8965,N_8374);
nor UO_1290 (O_1290,N_9780,N_9119);
xor UO_1291 (O_1291,N_8831,N_8393);
nor UO_1292 (O_1292,N_7517,N_8418);
nand UO_1293 (O_1293,N_8610,N_5112);
or UO_1294 (O_1294,N_6087,N_8397);
or UO_1295 (O_1295,N_8409,N_6254);
nor UO_1296 (O_1296,N_8917,N_8306);
and UO_1297 (O_1297,N_5809,N_6671);
or UO_1298 (O_1298,N_5619,N_8947);
and UO_1299 (O_1299,N_7872,N_9551);
nor UO_1300 (O_1300,N_7359,N_6301);
nand UO_1301 (O_1301,N_8435,N_9463);
nand UO_1302 (O_1302,N_6690,N_5174);
and UO_1303 (O_1303,N_6170,N_5040);
and UO_1304 (O_1304,N_6446,N_9079);
or UO_1305 (O_1305,N_8490,N_7681);
or UO_1306 (O_1306,N_5350,N_7142);
nor UO_1307 (O_1307,N_5522,N_7561);
and UO_1308 (O_1308,N_9064,N_6564);
nand UO_1309 (O_1309,N_7412,N_8820);
nand UO_1310 (O_1310,N_7615,N_6380);
or UO_1311 (O_1311,N_7956,N_9075);
and UO_1312 (O_1312,N_5594,N_8472);
nor UO_1313 (O_1313,N_6560,N_6930);
nor UO_1314 (O_1314,N_9913,N_6403);
or UO_1315 (O_1315,N_6458,N_5521);
and UO_1316 (O_1316,N_6109,N_9412);
or UO_1317 (O_1317,N_9807,N_9739);
and UO_1318 (O_1318,N_5816,N_6113);
nor UO_1319 (O_1319,N_5467,N_9370);
and UO_1320 (O_1320,N_6867,N_7522);
and UO_1321 (O_1321,N_6843,N_5660);
and UO_1322 (O_1322,N_9818,N_7796);
and UO_1323 (O_1323,N_6942,N_9592);
or UO_1324 (O_1324,N_7764,N_8635);
or UO_1325 (O_1325,N_9334,N_8471);
nor UO_1326 (O_1326,N_5151,N_5983);
nor UO_1327 (O_1327,N_6029,N_8832);
or UO_1328 (O_1328,N_8345,N_7974);
nor UO_1329 (O_1329,N_9613,N_7376);
nand UO_1330 (O_1330,N_8841,N_9439);
and UO_1331 (O_1331,N_7942,N_9964);
and UO_1332 (O_1332,N_7482,N_6473);
nand UO_1333 (O_1333,N_9791,N_9922);
nor UO_1334 (O_1334,N_9627,N_7401);
or UO_1335 (O_1335,N_5033,N_6486);
xor UO_1336 (O_1336,N_6588,N_5532);
xor UO_1337 (O_1337,N_8906,N_9522);
nand UO_1338 (O_1338,N_9836,N_9926);
and UO_1339 (O_1339,N_5899,N_6401);
xor UO_1340 (O_1340,N_8626,N_5956);
nor UO_1341 (O_1341,N_9429,N_9095);
nand UO_1342 (O_1342,N_7672,N_6515);
nand UO_1343 (O_1343,N_8308,N_8952);
nor UO_1344 (O_1344,N_8874,N_5379);
or UO_1345 (O_1345,N_5445,N_7292);
and UO_1346 (O_1346,N_6375,N_6272);
and UO_1347 (O_1347,N_8936,N_7451);
nand UO_1348 (O_1348,N_5669,N_5607);
nand UO_1349 (O_1349,N_8723,N_6437);
nand UO_1350 (O_1350,N_5454,N_9203);
nand UO_1351 (O_1351,N_9084,N_8975);
nand UO_1352 (O_1352,N_7967,N_6971);
nor UO_1353 (O_1353,N_5971,N_7441);
or UO_1354 (O_1354,N_6157,N_8538);
nand UO_1355 (O_1355,N_5055,N_6868);
nor UO_1356 (O_1356,N_5640,N_5037);
and UO_1357 (O_1357,N_5370,N_5459);
nand UO_1358 (O_1358,N_8311,N_5765);
or UO_1359 (O_1359,N_5656,N_6792);
nand UO_1360 (O_1360,N_8658,N_6501);
and UO_1361 (O_1361,N_9437,N_5472);
nor UO_1362 (O_1362,N_6910,N_5470);
nor UO_1363 (O_1363,N_8055,N_8669);
or UO_1364 (O_1364,N_6622,N_7739);
nor UO_1365 (O_1365,N_7205,N_5186);
nand UO_1366 (O_1366,N_7074,N_6222);
or UO_1367 (O_1367,N_9109,N_6001);
or UO_1368 (O_1368,N_8865,N_8628);
nor UO_1369 (O_1369,N_7530,N_6490);
nor UO_1370 (O_1370,N_6839,N_7877);
or UO_1371 (O_1371,N_6207,N_9169);
and UO_1372 (O_1372,N_7115,N_5632);
or UO_1373 (O_1373,N_8278,N_9640);
nor UO_1374 (O_1374,N_9394,N_7687);
or UO_1375 (O_1375,N_8464,N_9839);
nor UO_1376 (O_1376,N_8643,N_7548);
and UO_1377 (O_1377,N_8799,N_9823);
nor UO_1378 (O_1378,N_6646,N_9315);
or UO_1379 (O_1379,N_6963,N_7140);
nor UO_1380 (O_1380,N_9752,N_8781);
nor UO_1381 (O_1381,N_8876,N_5941);
and UO_1382 (O_1382,N_7371,N_8455);
nor UO_1383 (O_1383,N_9111,N_6795);
nor UO_1384 (O_1384,N_7649,N_9560);
xnor UO_1385 (O_1385,N_7187,N_8558);
nand UO_1386 (O_1386,N_7092,N_8637);
or UO_1387 (O_1387,N_5875,N_8359);
or UO_1388 (O_1388,N_6302,N_8363);
nor UO_1389 (O_1389,N_6120,N_5224);
and UO_1390 (O_1390,N_8566,N_5984);
nand UO_1391 (O_1391,N_8019,N_6747);
nor UO_1392 (O_1392,N_5507,N_8513);
nand UO_1393 (O_1393,N_5475,N_5559);
nand UO_1394 (O_1394,N_5501,N_5758);
and UO_1395 (O_1395,N_7007,N_8285);
nand UO_1396 (O_1396,N_9033,N_6073);
nor UO_1397 (O_1397,N_5265,N_8485);
nor UO_1398 (O_1398,N_6738,N_5500);
nor UO_1399 (O_1399,N_6965,N_6423);
nand UO_1400 (O_1400,N_7112,N_5206);
xnor UO_1401 (O_1401,N_6582,N_5481);
nand UO_1402 (O_1402,N_7132,N_7483);
nand UO_1403 (O_1403,N_5469,N_8217);
nand UO_1404 (O_1404,N_9683,N_9817);
nor UO_1405 (O_1405,N_7363,N_9811);
nand UO_1406 (O_1406,N_9086,N_5023);
nor UO_1407 (O_1407,N_5344,N_7789);
or UO_1408 (O_1408,N_7757,N_5187);
or UO_1409 (O_1409,N_9094,N_5168);
nor UO_1410 (O_1410,N_8375,N_9898);
nor UO_1411 (O_1411,N_7436,N_5052);
nor UO_1412 (O_1412,N_5110,N_8777);
nand UO_1413 (O_1413,N_7126,N_9953);
nand UO_1414 (O_1414,N_8430,N_9526);
or UO_1415 (O_1415,N_9763,N_8652);
and UO_1416 (O_1416,N_9367,N_7998);
and UO_1417 (O_1417,N_9715,N_5600);
and UO_1418 (O_1418,N_8035,N_9942);
nand UO_1419 (O_1419,N_5434,N_5604);
and UO_1420 (O_1420,N_7172,N_8267);
or UO_1421 (O_1421,N_8680,N_6774);
nor UO_1422 (O_1422,N_6406,N_6092);
or UO_1423 (O_1423,N_5889,N_8274);
or UO_1424 (O_1424,N_5225,N_8372);
or UO_1425 (O_1425,N_7935,N_6652);
nor UO_1426 (O_1426,N_6152,N_7551);
nor UO_1427 (O_1427,N_6069,N_7710);
or UO_1428 (O_1428,N_9494,N_9496);
and UO_1429 (O_1429,N_9649,N_5440);
xor UO_1430 (O_1430,N_9902,N_9205);
or UO_1431 (O_1431,N_8299,N_7554);
and UO_1432 (O_1432,N_8864,N_8385);
and UO_1433 (O_1433,N_9984,N_6453);
or UO_1434 (O_1434,N_5830,N_5891);
nor UO_1435 (O_1435,N_9912,N_6349);
and UO_1436 (O_1436,N_6227,N_9847);
nor UO_1437 (O_1437,N_8231,N_5154);
or UO_1438 (O_1438,N_8280,N_9540);
and UO_1439 (O_1439,N_9508,N_5250);
or UO_1440 (O_1440,N_8383,N_5293);
and UO_1441 (O_1441,N_6435,N_7997);
nor UO_1442 (O_1442,N_8271,N_9829);
nand UO_1443 (O_1443,N_6262,N_7147);
nand UO_1444 (O_1444,N_6893,N_9633);
nor UO_1445 (O_1445,N_8164,N_9087);
nor UO_1446 (O_1446,N_9747,N_9993);
nor UO_1447 (O_1447,N_9889,N_8797);
nand UO_1448 (O_1448,N_5716,N_7158);
nand UO_1449 (O_1449,N_7402,N_7755);
nand UO_1450 (O_1450,N_7797,N_8676);
and UO_1451 (O_1451,N_8326,N_5321);
nand UO_1452 (O_1452,N_5666,N_5738);
or UO_1453 (O_1453,N_5601,N_5671);
nor UO_1454 (O_1454,N_7930,N_5295);
nor UO_1455 (O_1455,N_6728,N_9469);
nand UO_1456 (O_1456,N_6838,N_8153);
nand UO_1457 (O_1457,N_8761,N_9226);
or UO_1458 (O_1458,N_6681,N_9531);
nand UO_1459 (O_1459,N_8530,N_5020);
and UO_1460 (O_1460,N_6580,N_8597);
and UO_1461 (O_1461,N_7297,N_9458);
nor UO_1462 (O_1462,N_8122,N_7593);
nand UO_1463 (O_1463,N_9872,N_9879);
nand UO_1464 (O_1464,N_6098,N_5800);
or UO_1465 (O_1465,N_8282,N_6764);
nand UO_1466 (O_1466,N_5436,N_5506);
nand UO_1467 (O_1467,N_9202,N_7636);
or UO_1468 (O_1468,N_5614,N_7838);
nor UO_1469 (O_1469,N_6280,N_9534);
nor UO_1470 (O_1470,N_5633,N_6791);
nor UO_1471 (O_1471,N_7079,N_8253);
and UO_1472 (O_1472,N_5296,N_8400);
nor UO_1473 (O_1473,N_9197,N_6130);
nand UO_1474 (O_1474,N_5705,N_9483);
or UO_1475 (O_1475,N_7339,N_9222);
or UO_1476 (O_1476,N_5586,N_8767);
and UO_1477 (O_1477,N_7771,N_8564);
or UO_1478 (O_1478,N_5451,N_8497);
nand UO_1479 (O_1479,N_9418,N_5740);
and UO_1480 (O_1480,N_5489,N_6081);
and UO_1481 (O_1481,N_8266,N_5832);
and UO_1482 (O_1482,N_8892,N_8448);
and UO_1483 (O_1483,N_7902,N_5582);
or UO_1484 (O_1484,N_6809,N_6704);
nand UO_1485 (O_1485,N_9528,N_5352);
and UO_1486 (O_1486,N_6093,N_7323);
nand UO_1487 (O_1487,N_9568,N_6459);
or UO_1488 (O_1488,N_6244,N_8252);
and UO_1489 (O_1489,N_8257,N_6691);
nor UO_1490 (O_1490,N_6277,N_9225);
or UO_1491 (O_1491,N_9931,N_8366);
nor UO_1492 (O_1492,N_7802,N_9206);
nand UO_1493 (O_1493,N_6368,N_9462);
or UO_1494 (O_1494,N_9755,N_7468);
or UO_1495 (O_1495,N_9144,N_9146);
nor UO_1496 (O_1496,N_6318,N_6285);
or UO_1497 (O_1497,N_5743,N_5959);
and UO_1498 (O_1498,N_9046,N_7623);
nor UO_1499 (O_1499,N_7272,N_7673);
endmodule